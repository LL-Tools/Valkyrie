

module b17_C_SARLock_k_64_10 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, U355, U356, U357, U358, 
        U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, 
        U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, 
        U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, 
        U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, 
        U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, 
        U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, 
        U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, 
        U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9911, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
         n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
         n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
         n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
         n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
         n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
         n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
         n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
         n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
         n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
         n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
         n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812,
         n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
         n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
         n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
         n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
         n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
         n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
         n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
         n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108,
         n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
         n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
         n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
         n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
         n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
         n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
         n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
         n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
         n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931;

  INV_X1 U11030 ( .A(n14758), .ZN(n14899) );
  AND2_X1 U11031 ( .A1(n9976), .A2(n9975), .ZN(n15288) );
  NAND2_X1 U11033 ( .A1(n12653), .A2(n12651), .ZN(n15846) );
  INV_X1 U11034 ( .A(n18215), .ZN(n17209) );
  BUF_X2 U11036 ( .A(n12718), .Z(n17125) );
  AND2_X1 U11037 ( .A1(n10375), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10440) );
  INV_X1 U11038 ( .A(n16984), .ZN(n17108) );
  CLKBUF_X1 U11040 ( .A(n12381), .Z(n12476) );
  BUF_X1 U11041 ( .A(n11475), .Z(n20076) );
  CLKBUF_X2 U11042 ( .A(n11362), .Z(n12435) );
  INV_X1 U11043 ( .A(n11553), .ZN(n11518) );
  NAND3_X1 U11044 ( .A1(n13145), .A2(n10277), .A3(n10096), .ZN(n11249) );
  BUF_X2 U11045 ( .A(n11415), .Z(n12486) );
  AND2_X2 U11046 ( .A1(n14053), .A2(n10528), .ZN(n10235) );
  AND2_X1 U11047 ( .A1(n13640), .A2(n13435), .ZN(n11386) );
  AND2_X1 U11048 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11328) );
  CLKBUF_X1 U11049 ( .A(n19908), .Z(n9585) );
  NOR2_X1 U11050 ( .A1(n14106), .A2(n14096), .ZN(n19908) );
  NOR2_X1 U11051 ( .A1(n10577), .A2(n10576), .ZN(n10111) );
  AND2_X1 U11054 ( .A1(n11465), .A2(n12000), .ZN(n11495) );
  AND2_X2 U11055 ( .A1(n14053), .A2(n10528), .ZN(n9587) );
  XNOR2_X1 U11056 ( .A(n10577), .B(n10576), .ZN(n10752) );
  AOI21_X1 U11057 ( .B1(n10254), .B2(n10275), .A(n10233), .ZN(n10970) );
  AND4_X1 U11059 ( .A1(n11366), .A2(n11365), .A3(n11364), .A4(n11363), .ZN(
        n11377) );
  INV_X1 U11060 ( .A(n12987), .ZN(n11178) );
  AND2_X1 U11061 ( .A1(n9586), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10418) );
  AND2_X1 U11062 ( .A1(n10375), .A2(n15811), .ZN(n10434) );
  NAND2_X1 U11063 ( .A1(n10261), .A2(n10297), .ZN(n10327) );
  INV_X1 U11064 ( .A(n17147), .ZN(n14469) );
  NAND2_X1 U11065 ( .A1(n9756), .A2(n11492), .ZN(n11546) );
  NOR2_X1 U11066 ( .A1(n10867), .A2(n10085), .ZN(n10084) );
  CLKBUF_X2 U11067 ( .A(n10323), .Z(n10784) );
  NAND2_X1 U11068 ( .A1(n10094), .A2(n9798), .ZN(n10641) );
  INV_X1 U11069 ( .A(n12870), .ZN(n10350) );
  OR2_X2 U11070 ( .A1(n15855), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12600) );
  NOR3_X1 U11071 ( .A1(n18207), .A2(n12649), .A3(n12661), .ZN(n12667) );
  INV_X1 U11072 ( .A(n14469), .ZN(n17109) );
  INV_X1 U11073 ( .A(n9635), .ZN(n17142) );
  AND4_X1 U11074 ( .A1(n11390), .A2(n11389), .A3(n11388), .A4(n11387), .ZN(
        n11402) );
  NAND2_X1 U11075 ( .A1(n10631), .A2(n10168), .ZN(n10890) );
  OR2_X1 U11076 ( .A1(n10647), .A2(n10646), .ZN(n10662) );
  AND2_X1 U11077 ( .A1(n10631), .A2(n10616), .ZN(n10630) );
  OAI21_X1 U11078 ( .B1(n14542), .B2(n14543), .A(n10905), .ZN(n10911) );
  NAND2_X1 U11079 ( .A1(n10874), .A2(n15494), .ZN(n15489) );
  NAND2_X1 U11080 ( .A1(n10569), .A2(n10568), .ZN(n14079) );
  INV_X1 U11081 ( .A(n18658), .ZN(n18634) );
  BUF_X2 U11082 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n16322) );
  INV_X1 U11083 ( .A(n18225), .ZN(n16928) );
  NOR2_X1 U11084 ( .A1(n12611), .A2(n12610), .ZN(n17353) );
  INV_X1 U11085 ( .A(n14278), .ZN(n14276) );
  AOI211_X1 U11086 ( .C1(n20717), .C2(n19980), .A(n19946), .B(n19945), .ZN(
        n19953) );
  OAI21_X1 U11087 ( .B1(n14572), .B2(n14573), .A(n9608), .ZN(n14889) );
  INV_X1 U11088 ( .A(n17151), .ZN(n12605) );
  XNOR2_X1 U11089 ( .A(n11546), .B(n11506), .ZN(n12014) );
  NAND2_X2 U11091 ( .A1(n10613), .A2(n9621), .ZN(n10094) );
  NOR2_X2 U11092 ( .A1(n15133), .A2(n11764), .ZN(n11765) );
  NAND2_X2 U11093 ( .A1(n15489), .A2(n15488), .ZN(n15490) );
  OAI21_X2 U11095 ( .B1(n13523), .B2(n13524), .A(n12868), .ZN(n13538) );
  AND2_X1 U11096 ( .A1(n14053), .A2(n10528), .ZN(n9586) );
  INV_X4 U11098 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10528) );
  AOI21_X2 U11099 ( .B1(n14967), .B2(n11760), .A(n11759), .ZN(n15132) );
  AND2_X4 U11100 ( .A1(n14128), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10225) );
  NOR2_X4 U11101 ( .A1(n16905), .A2(n12561), .ZN(n17147) );
  AND2_X4 U11104 ( .A1(n13297), .A2(n19839), .ZN(n11308) );
  INV_X2 U11105 ( .A(n10364), .ZN(n13297) );
  NOR2_X1 U11106 ( .A1(n12568), .A2(n12567), .ZN(n12716) );
  INV_X4 U11107 ( .A(n12600), .ZN(n14458) );
  NAND2_X1 U11108 ( .A1(n10854), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15481) );
  CLKBUF_X2 U11109 ( .A(n11753), .Z(n15136) );
  AND2_X1 U11110 ( .A1(n12800), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17488) );
  NOR2_X1 U11111 ( .A1(n12800), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17487) );
  INV_X2 U11112 ( .A(n19983), .ZN(n19958) );
  INV_X1 U11113 ( .A(n10752), .ZN(n9589) );
  OAI21_X1 U11114 ( .B1(n10552), .B2(n9760), .A(n10744), .ZN(n13816) );
  NOR3_X1 U11115 ( .A1(n17529), .A2(n17537), .A3(n17898), .ZN(n12796) );
  CLKBUF_X1 U11116 ( .A(n13680), .Z(n9595) );
  INV_X2 U11117 ( .A(n17848), .ZN(n17837) );
  OR2_X1 U11118 ( .A1(n10357), .A2(n12860), .ZN(n10359) );
  OR2_X1 U11119 ( .A1(n12373), .A2(n12372), .ZN(n12412) );
  AND2_X1 U11120 ( .A1(n12860), .A2(n15792), .ZN(n10349) );
  AND2_X1 U11121 ( .A1(n10338), .A2(n13541), .ZN(n19239) );
  NOR2_X1 U11122 ( .A1(n18901), .A2(n18903), .ZN(n18902) );
  INV_X2 U11123 ( .A(n18626), .ZN(n17918) );
  AND2_X1 U11124 ( .A1(n11546), .A2(n11545), .ZN(n11598) );
  NAND2_X2 U11125 ( .A1(n18635), .A2(n18634), .ZN(n18078) );
  INV_X2 U11126 ( .A(n18633), .ZN(n18635) );
  AOI21_X1 U11127 ( .B1(n12656), .B2(n12650), .A(n13255), .ZN(n12668) );
  NAND2_X1 U11128 ( .A1(n10630), .A2(n10629), .ZN(n10633) );
  NAND2_X1 U11129 ( .A1(n17418), .A2(n15847), .ZN(n13255) );
  NOR3_X2 U11130 ( .A1(n17353), .A2(n18215), .A3(n15846), .ZN(n17416) );
  AND3_X1 U11131 ( .A1(n13430), .A2(n11478), .A3(n11971), .ZN(n11494) );
  NOR2_X1 U11133 ( .A1(n18185), .A2(n16928), .ZN(n12656) );
  AND2_X1 U11134 ( .A1(n10962), .A2(n19831), .ZN(n16363) );
  NAND2_X1 U11135 ( .A1(n11537), .A2(n15926), .ZN(n14111) );
  INV_X1 U11136 ( .A(n20061), .ZN(n11537) );
  NAND2_X1 U11137 ( .A1(n11479), .A2(n9842), .ZN(n11487) );
  INV_X4 U11138 ( .A(n10038), .ZN(n11054) );
  NAND2_X1 U11140 ( .A1(n9795), .A2(n10168), .ZN(n10254) );
  NAND2_X1 U11141 ( .A1(n13196), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13193) );
  INV_X2 U11142 ( .A(n10217), .ZN(n10264) );
  NAND2_X2 U11143 ( .A1(n9797), .A2(n9796), .ZN(n13298) );
  INV_X2 U11144 ( .A(n9604), .ZN(n17116) );
  BUF_X2 U11146 ( .A(n12599), .Z(n17159) );
  BUF_X2 U11148 ( .A(n10241), .Z(n13133) );
  CLKBUF_X2 U11149 ( .A(n11412), .Z(n12484) );
  CLKBUF_X2 U11150 ( .A(n10374), .Z(n13129) );
  AND2_X2 U11151 ( .A1(n13638), .A2(n13436), .ZN(n11362) );
  NOR2_X4 U11152 ( .A1(n12567), .A2(n12563), .ZN(n17151) );
  BUF_X4 U11153 ( .A(n10202), .Z(n9590) );
  NOR2_X2 U11155 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13436) );
  NAND2_X1 U11156 ( .A1(n12463), .A2(n12462), .ZN(n14877) );
  NAND2_X1 U11157 ( .A1(n9608), .A2(n12461), .ZN(n12462) );
  XNOR2_X1 U11158 ( .A(n12542), .B(n12541), .ZN(n14489) );
  AOI21_X1 U11159 ( .B1(n11301), .B2(n16271), .A(n9778), .ZN(n10013) );
  AOI21_X1 U11160 ( .B1(n15582), .B2(n11010), .A(n14541), .ZN(n15571) );
  NAND2_X1 U11161 ( .A1(n11769), .A2(n15136), .ZN(n14911) );
  CLKBUF_X1 U11162 ( .A(n15453), .Z(n15461) );
  OR2_X1 U11163 ( .A1(n15293), .A2(n15295), .ZN(n9980) );
  CLKBUF_X1 U11164 ( .A(n15746), .Z(n15747) );
  XNOR2_X1 U11165 ( .A(n13070), .B(n10134), .ZN(n15293) );
  OR2_X1 U11166 ( .A1(n14949), .A2(n11767), .ZN(n11768) );
  NAND2_X1 U11167 ( .A1(n15299), .A2(n10130), .ZN(n13070) );
  NOR2_X1 U11168 ( .A1(n16049), .A2(n9845), .ZN(n14979) );
  OR2_X1 U11169 ( .A1(n14968), .A2(n14980), .ZN(n15133) );
  OAI22_X1 U11170 ( .A1(n14079), .A2(n14078), .B1(n10572), .B2(n14199), .ZN(
        n14190) );
  NAND2_X1 U11171 ( .A1(n11702), .A2(n11701), .ZN(n14141) );
  NOR2_X1 U11172 ( .A1(n15312), .A2(n15231), .ZN(n15233) );
  AND2_X1 U11173 ( .A1(n16033), .A2(n16037), .ZN(n11760) );
  OR2_X1 U11174 ( .A1(n14343), .A2(n14342), .ZN(n9763) );
  INV_X1 U11175 ( .A(n17216), .ZN(n17211) );
  OR2_X1 U11176 ( .A1(n15136), .A2(n11917), .ZN(n16037) );
  NAND2_X1 U11177 ( .A1(n9589), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14192) );
  AND2_X1 U11178 ( .A1(n10760), .A2(n10110), .ZN(n10758) );
  OR2_X1 U11179 ( .A1(n10760), .A2(n10628), .ZN(n10766) );
  NAND2_X1 U11180 ( .A1(n11292), .A2(n11247), .ZN(n11305) );
  NAND2_X1 U11181 ( .A1(n11731), .A2(n11743), .ZN(n11753) );
  OR2_X1 U11182 ( .A1(n10111), .A2(n10753), .ZN(n10110) );
  NOR2_X1 U11183 ( .A1(n15679), .A2(n11268), .ZN(n15651) );
  NAND2_X1 U11184 ( .A1(n9758), .A2(n11657), .ZN(n13768) );
  OR2_X1 U11185 ( .A1(n17520), .A2(n12797), .ZN(n12798) );
  NAND2_X1 U11186 ( .A1(n9831), .A2(n9664), .ZN(n15679) );
  INV_X1 U11187 ( .A(n15683), .ZN(n9831) );
  AND2_X1 U11188 ( .A1(n15218), .A2(n9949), .ZN(n15197) );
  NOR2_X1 U11189 ( .A1(n14136), .A2(n14137), .ZN(n14174) );
  XNOR2_X1 U11190 ( .A(n14099), .B(n14098), .ZN(n14492) );
  OR2_X1 U11191 ( .A1(n16267), .A2(n11266), .ZN(n15683) );
  OR2_X1 U11192 ( .A1(n13956), .A2(n14070), .ZN(n14136) );
  OR2_X1 U11193 ( .A1(n14097), .A2(n20877), .ZN(n14099) );
  AND2_X1 U11194 ( .A1(n13534), .A2(n13533), .ZN(n13740) );
  AND2_X1 U11195 ( .A1(n10609), .A2(n10608), .ZN(n10753) );
  NAND2_X1 U11196 ( .A1(n10502), .A2(n10501), .ZN(n10576) );
  NOR2_X1 U11197 ( .A1(n16299), .A2(n11263), .ZN(n15783) );
  AND2_X1 U11198 ( .A1(n11618), .A2(n12125), .ZN(n9995) );
  AND4_X1 U11199 ( .A1(n10344), .A2(n10343), .A3(n10342), .A4(n10341), .ZN(
        n10363) );
  OR2_X1 U11200 ( .A1(n16155), .A2(n10628), .ZN(n10884) );
  XNOR2_X1 U11201 ( .A(n13461), .B(n11568), .ZN(n13689) );
  AND2_X1 U11202 ( .A1(n12879), .A2(n13579), .ZN(n13539) );
  NOR2_X2 U11203 ( .A1(n12531), .A2(n20053), .ZN(n12532) );
  NAND2_X1 U11204 ( .A1(n11650), .A2(n11649), .ZN(n20211) );
  INV_X1 U11205 ( .A(n10587), .ZN(n19269) );
  NAND2_X1 U11206 ( .A1(n13462), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13461) );
  OR2_X1 U11207 ( .A1(n18914), .A2(n10684), .ZN(n15527) );
  NAND2_X1 U11208 ( .A1(n10349), .A2(n10352), .ZN(n19547) );
  NAND2_X1 U11209 ( .A1(n9609), .A2(n10352), .ZN(n10474) );
  OAI22_X1 U11210 ( .A1(n10339), .A2(n19359), .B1(n19576), .B2(n10369), .ZN(
        n10340) );
  NOR2_X2 U11211 ( .A1(n10095), .A2(n10358), .ZN(n10482) );
  OR2_X1 U11212 ( .A1(n15263), .A2(n10628), .ZN(n10694) );
  NAND2_X1 U11213 ( .A1(n18842), .A2(n16538), .ZN(n17848) );
  AND2_X1 U11214 ( .A1(n9834), .A2(n9832), .ZN(n13827) );
  NAND2_X1 U11215 ( .A1(n10350), .A2(n9610), .ZN(n19576) );
  AOI22_X1 U11216 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19239), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10342) );
  NAND2_X1 U11217 ( .A1(n9610), .A2(n13541), .ZN(n10579) );
  OAI21_X1 U11218 ( .B1(n12013), .B2(n11813), .A(n11539), .ZN(n13462) );
  NAND2_X1 U11219 ( .A1(n9609), .A2(n9643), .ZN(n19330) );
  NAND2_X1 U11220 ( .A1(n10349), .A2(n9643), .ZN(n10587) );
  AND2_X1 U11221 ( .A1(n10335), .A2(n10350), .ZN(n10468) );
  AND2_X1 U11222 ( .A1(n10683), .A2(n10685), .ZN(n10691) );
  NAND2_X1 U11223 ( .A1(n12875), .A2(n12874), .ZN(n12881) );
  AND2_X1 U11224 ( .A1(n10330), .A2(n13541), .ZN(n19179) );
  AND2_X1 U11225 ( .A1(n10698), .A2(n10697), .ZN(n18904) );
  AND2_X1 U11226 ( .A1(n10068), .A2(n10069), .ZN(n17671) );
  NAND2_X1 U11227 ( .A1(n9850), .A2(n11531), .ZN(n11573) );
  OR2_X1 U11228 ( .A1(n12870), .A2(n12869), .ZN(n12875) );
  NAND2_X1 U11229 ( .A1(n11258), .A2(n11033), .ZN(n19128) );
  NAND2_X1 U11230 ( .A1(n11548), .A2(n11547), .ZN(n20502) );
  INV_X1 U11231 ( .A(n15792), .ZN(n10358) );
  AND2_X1 U11232 ( .A1(n11008), .A2(n13220), .ZN(n11258) );
  AND2_X1 U11233 ( .A1(n10677), .A2(n9683), .ZN(n10702) );
  CLKBUF_X1 U11234 ( .A(n12014), .Z(n9594) );
  AND2_X1 U11235 ( .A1(n18912), .A2(n18911), .ZN(n18921) );
  NOR2_X2 U11236 ( .A1(n18078), .A2(n18654), .ZN(n18120) );
  OAI21_X2 U11237 ( .B1(n13963), .B2(n12869), .A(n12866), .ZN(n13968) );
  AOI21_X2 U11238 ( .B1(n15963), .B2(n15962), .A(n18839), .ZN(n17202) );
  NOR2_X2 U11239 ( .A1(n19150), .A2(n19363), .ZN(n19151) );
  NOR2_X2 U11240 ( .A1(n14283), .A2(n19363), .ZN(n14284) );
  NOR2_X2 U11241 ( .A1(n19065), .A2(n19363), .ZN(n14299) );
  OR2_X1 U11242 ( .A1(n17765), .A2(n18094), .ZN(n17763) );
  NAND2_X1 U11243 ( .A1(n11584), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9756) );
  NAND2_X1 U11244 ( .A1(n10313), .A2(n10312), .ZN(n10333) );
  XNOR2_X1 U11245 ( .A(n10781), .B(n10782), .ZN(n10778) );
  INV_X2 U11246 ( .A(n17354), .ZN(n17397) );
  NAND2_X1 U11247 ( .A1(n10329), .A2(n10328), .ZN(n10782) );
  NAND2_X1 U11248 ( .A1(n10326), .A2(n10325), .ZN(n10781) );
  NAND3_X1 U11249 ( .A1(n10299), .A2(n10298), .A3(n10123), .ZN(n10310) );
  NOR2_X1 U11250 ( .A1(n11067), .A2(n11066), .ZN(n11073) );
  AND2_X1 U11251 ( .A1(n10728), .A2(n11013), .ZN(n10979) );
  AND2_X1 U11252 ( .A1(n10122), .A2(n10293), .ZN(n10299) );
  OR2_X1 U11253 ( .A1(n10292), .A2(n13325), .ZN(n10122) );
  CLKBUF_X1 U11254 ( .A(n12515), .Z(n13431) );
  OR2_X1 U11255 ( .A1(n10562), .A2(n10563), .ZN(n10545) );
  AND2_X1 U11256 ( .A1(n11020), .A2(n19833), .ZN(n11032) );
  INV_X1 U11257 ( .A(n10547), .ZN(n9894) );
  INV_X4 U11258 ( .A(n10936), .ZN(n10940) );
  AND2_X1 U11259 ( .A1(n10234), .A2(n10269), .ZN(n10288) );
  OR2_X1 U11260 ( .A1(n10466), .A2(n10465), .ZN(n11081) );
  NAND2_X1 U11261 ( .A1(n11495), .A2(n11466), .ZN(n9754) );
  AND2_X1 U11262 ( .A1(n11380), .A2(n11379), .ZN(n11421) );
  NAND2_X1 U11263 ( .A1(n10098), .A2(n13221), .ZN(n13145) );
  OR2_X1 U11264 ( .A1(n11481), .A2(n11483), .ZN(n11466) );
  OR2_X1 U11265 ( .A1(n11055), .A2(n11054), .ZN(n11077) );
  NAND2_X2 U11266 ( .A1(n15926), .A2(n20061), .ZN(n11496) );
  NAND3_X1 U11267 ( .A1(n12638), .A2(n12637), .A3(n12636), .ZN(n18215) );
  OR2_X1 U11268 ( .A1(n10451), .A2(n10450), .ZN(n10734) );
  INV_X2 U11269 ( .A(n18193), .ZN(n18842) );
  NAND3_X1 U11270 ( .A1(n12701), .A2(n12700), .A3(n12699), .ZN(n12813) );
  NAND2_X2 U11271 ( .A1(n9638), .A2(n9753), .ZN(n20061) );
  NAND2_X1 U11272 ( .A1(n10168), .A2(n13298), .ZN(n11060) );
  INV_X1 U11273 ( .A(n13221), .ZN(n19833) );
  NAND2_X1 U11274 ( .A1(n11475), .A2(n9858), .ZN(n11938) );
  NAND2_X1 U11275 ( .A1(n10364), .A2(n19839), .ZN(n11055) );
  NAND4_X2 U11276 ( .A1(n9784), .A2(n9641), .A3(n12617), .A4(n12612), .ZN(
        n18225) );
  CLKBUF_X1 U11277 ( .A(n11476), .Z(n12464) );
  OR2_X1 U11278 ( .A1(n10500), .A2(n10499), .ZN(n11086) );
  OR2_X1 U11279 ( .A1(n10382), .A2(n10381), .ZN(n10537) );
  CLKBUF_X1 U11280 ( .A(n10233), .Z(n19167) );
  AND2_X1 U11281 ( .A1(n10364), .A2(n10274), .ZN(n19831) );
  AOI211_X1 U11282 ( .C1(n17116), .C2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A(
        n12698), .B(n12697), .ZN(n12699) );
  AND4_X1 U11283 ( .A1(n10511), .A2(n10510), .A3(n10509), .A4(n10508), .ZN(
        n10523) );
  CLKBUF_X1 U11284 ( .A(n11536), .Z(n20093) );
  INV_X2 U11285 ( .A(n13121), .ZN(n10364) );
  AND2_X1 U11286 ( .A1(n9959), .A2(n9961), .ZN(n9955) );
  NOR2_X1 U11287 ( .A1(n12737), .A2(n12736), .ZN(n17335) );
  NAND4_X2 U11288 ( .A1(n11463), .A2(n11462), .A3(n11461), .A4(n11460), .ZN(
        n11475) );
  AND4_X1 U11289 ( .A1(n10507), .A2(n10506), .A3(n10505), .A4(n10504), .ZN(
        n10524) );
  AND3_X1 U11290 ( .A1(n10143), .A2(n11417), .A3(n11416), .ZN(n11418) );
  OR2_X2 U11291 ( .A1(n11356), .A2(n11355), .ZN(n11477) );
  NAND2_X1 U11292 ( .A1(n9961), .A2(n9960), .ZN(n19154) );
  NAND2_X1 U11293 ( .A1(n10232), .A2(n10231), .ZN(n13121) );
  NOR2_X1 U11294 ( .A1(n9616), .A2(n9650), .ZN(n9753) );
  AND4_X1 U11295 ( .A1(n11430), .A2(n11429), .A3(n11428), .A4(n11427), .ZN(
        n11440) );
  AND4_X1 U11296 ( .A1(n11395), .A2(n11394), .A3(n11393), .A4(n11392), .ZN(
        n11401) );
  NAND3_X1 U11297 ( .A1(n10167), .A2(n10166), .A3(n10132), .ZN(n9796) );
  NAND2_X1 U11298 ( .A1(n10200), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9958) );
  NAND3_X1 U11299 ( .A1(n10162), .A2(n10131), .A3(n10161), .ZN(n9797) );
  NAND2_X1 U11300 ( .A1(n10133), .A2(n10172), .ZN(n9961) );
  AND4_X1 U11301 ( .A1(n11325), .A2(n11324), .A3(n11323), .A4(n11322), .ZN(
        n11334) );
  AND4_X1 U11302 ( .A1(n11332), .A2(n11331), .A3(n11330), .A4(n11329), .ZN(
        n11333) );
  AND4_X1 U11303 ( .A1(n11361), .A2(n11360), .A3(n11359), .A4(n11358), .ZN(
        n11378) );
  AND4_X1 U11304 ( .A1(n11451), .A2(n11450), .A3(n11449), .A4(n11448), .ZN(
        n11462) );
  INV_X2 U11305 ( .A(n16984), .ZN(n17144) );
  AND4_X1 U11306 ( .A1(n10199), .A2(n10198), .A3(n10197), .A4(n10196), .ZN(
        n10200) );
  NAND2_X2 U11307 ( .A1(n18786), .A2(n18718), .ZN(n18768) );
  INV_X1 U11308 ( .A(n12600), .ZN(n17126) );
  INV_X2 U11309 ( .A(n18725), .ZN(n9591) );
  AOI22_X1 U11310 ( .A1(n11362), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11335), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11338) );
  AND4_X1 U11311 ( .A1(n11374), .A2(n11373), .A3(n11372), .A4(n11371), .ZN(
        n11375) );
  AND3_X1 U11312 ( .A1(n10238), .A2(n10237), .A3(n10236), .ZN(n10239) );
  BUF_X2 U11313 ( .A(n11345), .Z(n12289) );
  AND2_X2 U11314 ( .A1(n13129), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10426) );
  INV_X2 U11315 ( .A(n16523), .ZN(U215) );
  NAND2_X2 U11316 ( .A1(n19858), .A2(n19740), .ZN(n19779) );
  NAND2_X2 U11317 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19858), .ZN(n19780) );
  BUF_X2 U11318 ( .A(n11406), .Z(n12359) );
  BUF_X2 U11319 ( .A(n11391), .Z(n12395) );
  BUF_X2 U11320 ( .A(n11386), .Z(n12485) );
  INV_X2 U11321 ( .A(n20740), .ZN(n20017) );
  OR2_X2 U11322 ( .A1(n13464), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16134) );
  INV_X2 U11323 ( .A(n11519), .ZN(n9593) );
  INV_X2 U11324 ( .A(n16527), .ZN(n16529) );
  CLKBUF_X2 U11325 ( .A(n10225), .Z(n9596) );
  AND2_X2 U11326 ( .A1(n13002), .A2(n15811), .ZN(n10445) );
  NAND2_X1 U11327 ( .A1(n9791), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15855) );
  INV_X2 U11328 ( .A(n18661), .ZN(n18650) );
  CLKBUF_X2 U11329 ( .A(n11415), .Z(n12422) );
  AND2_X2 U11330 ( .A1(n11326), .A2(n11328), .ZN(n11517) );
  NAND2_X1 U11331 ( .A1(n18798), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12567) );
  NAND2_X1 U11332 ( .A1(n18821), .A2(n12565), .ZN(n16905) );
  NOR2_X1 U11333 ( .A1(n12565), .A2(n18821), .ZN(n18661) );
  AND2_X1 U11334 ( .A1(n9839), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13640) );
  AND2_X2 U11335 ( .A1(n11328), .A2(n13435), .ZN(n11407) );
  AND2_X1 U11337 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14054) );
  NAND2_X1 U11338 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13203) );
  INV_X1 U11339 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15811) );
  NAND2_X1 U11340 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12564) );
  INV_X1 U11341 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18798) );
  NOR2_X2 U11342 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11327) );
  NAND2_X1 U11343 ( .A1(n20717), .A2(n20744), .ZN(n11650) );
  AOI21_X2 U11344 ( .B1(n11562), .B2(n20744), .A(n10127), .ZN(n12004) );
  NAND2_X2 U11345 ( .A1(n10327), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n9764) );
  INV_X2 U11346 ( .A(n13207), .ZN(n9951) );
  XNOR2_X1 U11347 ( .A(n12007), .B(n12006), .ZN(n13680) );
  NAND2_X2 U11348 ( .A1(n10314), .A2(n10345), .ZN(n10332) );
  AND2_X2 U11349 ( .A1(n10316), .A2(n10319), .ZN(n10314) );
  NAND4_X2 U11350 ( .A1(n10280), .A2(n10268), .A3(n9765), .A4(n9764), .ZN(
        n10316) );
  NOR2_X2 U11352 ( .A1(n11249), .A2(n10972), .ZN(n11049) );
  AND2_X1 U11353 ( .A1(n14128), .A2(n10528), .ZN(n9597) );
  AND2_X1 U11354 ( .A1(n11032), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9598) );
  AND2_X4 U11355 ( .A1(n11032), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9599) );
  AND2_X2 U11356 ( .A1(n11032), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10926) );
  INV_X1 U11357 ( .A(n10364), .ZN(n9600) );
  INV_X1 U11358 ( .A(n13297), .ZN(n10383) );
  AND2_X2 U11359 ( .A1(n9596), .A2(n15811), .ZN(n10503) );
  AND2_X1 U11360 ( .A1(n14128), .A2(n10528), .ZN(n10202) );
  AND2_X1 U11361 ( .A1(n20061), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11532) );
  OR2_X1 U11362 ( .A1(n11483), .A2(n20744), .ZN(n11637) );
  AOI21_X1 U11363 ( .B1(n11807), .B2(n11806), .A(n11797), .ZN(n11801) );
  AOI21_X1 U11364 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19803), .A(
        n10541), .ZN(n10710) );
  AND2_X1 U11365 ( .A1(n15460), .A2(n15455), .ZN(n10892) );
  NAND2_X1 U11366 ( .A1(n11060), .A2(n11025), .ZN(n9777) );
  INV_X1 U11367 ( .A(n11837), .ZN(n11824) );
  INV_X1 U11368 ( .A(n11572), .ZN(n9852) );
  INV_X1 U11369 ( .A(n11651), .ZN(n9854) );
  INV_X1 U11370 ( .A(n11814), .ZN(n11847) );
  AND2_X1 U11371 ( .A1(n10527), .A2(n10526), .ZN(n10533) );
  OR2_X1 U11372 ( .A1(n10982), .A2(n10711), .ZN(n10527) );
  AND2_X1 U11373 ( .A1(n10539), .A2(n10538), .ZN(n10541) );
  NOR3_X1 U11374 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n11798), .A3(
        n11802), .ZN(n11818) );
  NAND2_X1 U11375 ( .A1(n11970), .A2(n11484), .ZN(n11783) );
  INV_X1 U11376 ( .A(n14224), .ZN(n10001) );
  NAND2_X1 U11377 ( .A1(n14573), .A2(n10012), .ZN(n10011) );
  INV_X1 U11378 ( .A(n14588), .ZN(n10012) );
  NAND2_X1 U11379 ( .A1(n14378), .A2(n14733), .ZN(n9998) );
  XNOR2_X1 U11380 ( .A(n11731), .B(n11730), .ZN(n12064) );
  INV_X1 U11381 ( .A(n12035), .ZN(n12499) );
  OR2_X1 U11382 ( .A1(n12000), .A2(n12409), .ZN(n12453) );
  OR2_X1 U11383 ( .A1(n11960), .A2(n11914), .ZN(n11959) );
  CLKBUF_X1 U11384 ( .A(n11537), .Z(n14092) );
  NAND2_X1 U11385 ( .A1(n11532), .A2(n11483), .ZN(n11814) );
  OR2_X1 U11386 ( .A1(n11968), .A2(n11938), .ZN(n13430) );
  NOR2_X1 U11387 ( .A1(n11814), .A2(n11813), .ZN(n11841) );
  NAND2_X1 U11388 ( .A1(n11850), .A2(n9751), .ZN(n9750) );
  NAND2_X1 U11389 ( .A1(n20744), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n9751) );
  AND4_X1 U11390 ( .A1(n11459), .A2(n11458), .A3(n11457), .A4(n11456), .ZN(
        n11460) );
  AND4_X1 U11391 ( .A1(n11446), .A2(n11445), .A3(n11444), .A4(n11443), .ZN(
        n11463) );
  AND4_X1 U11392 ( .A1(n11455), .A2(n11454), .A3(n11453), .A4(n11452), .ZN(
        n11461) );
  INV_X1 U11393 ( .A(n15476), .ZN(n10089) );
  NOR2_X1 U11394 ( .A1(n15475), .A2(n10091), .ZN(n10090) );
  INV_X1 U11395 ( .A(n10878), .ZN(n10091) );
  AND2_X1 U11396 ( .A1(n15517), .A2(n9815), .ZN(n9812) );
  INV_X1 U11397 ( .A(n10640), .ZN(n10088) );
  OR2_X1 U11398 ( .A1(n13919), .A2(n10628), .ZN(n10645) );
  AND2_X1 U11399 ( .A1(n10099), .A2(n10097), .ZN(n10096) );
  AND2_X1 U11400 ( .A1(n10252), .A2(n11021), .ZN(n10277) );
  OAI21_X1 U11401 ( .B1(n10274), .B2(n10275), .A(n19154), .ZN(n10097) );
  AND2_X1 U11402 ( .A1(n10214), .A2(n10531), .ZN(n10265) );
  NAND2_X1 U11403 ( .A1(n9836), .A2(n9835), .ZN(n11001) );
  NAND2_X1 U11404 ( .A1(n13325), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n9835) );
  OAI21_X1 U11405 ( .B1(n10998), .B2(n10999), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n9836) );
  AND2_X1 U11406 ( .A1(n12864), .A2(n9963), .ZN(n9962) );
  NAND2_X1 U11407 ( .A1(n12862), .A2(n12869), .ZN(n9963) );
  INV_X1 U11408 ( .A(n12690), .ZN(n16984) );
  NOR2_X1 U11409 ( .A1(n18650), .A2(n12566), .ZN(n12717) );
  NOR2_X1 U11410 ( .A1(n12628), .A2(n12627), .ZN(n12671) );
  NOR2_X1 U11411 ( .A1(n15846), .A2(n18645), .ZN(n15848) );
  OR2_X1 U11412 ( .A1(n14112), .A2(n14092), .ZN(n14106) );
  OR2_X1 U11414 ( .A1(n11987), .A2(n13290), .ZN(n16098) );
  INV_X1 U11415 ( .A(n10274), .ZN(n19846) );
  AND2_X1 U11416 ( .A1(n11286), .A2(n9689), .ZN(n13180) );
  INV_X1 U11417 ( .A(n13181), .ZN(n10053) );
  AND2_X1 U11418 ( .A1(n13565), .A2(n13563), .ZN(n13564) );
  NAND2_X1 U11419 ( .A1(n13126), .A2(n9973), .ZN(n9972) );
  NAND2_X1 U11420 ( .A1(n9981), .A2(n9978), .ZN(n9977) );
  NAND2_X1 U11421 ( .A1(n13071), .A2(n9981), .ZN(n9974) );
  INV_X1 U11422 ( .A(n10628), .ZN(n11094) );
  AOI21_X1 U11423 ( .B1(n13181), .B2(n15176), .A(n13180), .ZN(n15419) );
  AOI21_X1 U11424 ( .B1(n9812), .B2(n9810), .A(n9809), .ZN(n9808) );
  INV_X1 U11425 ( .A(n10856), .ZN(n9810) );
  INV_X1 U11426 ( .A(n10859), .ZN(n9809) );
  INV_X1 U11427 ( .A(n9812), .ZN(n9811) );
  INV_X1 U11428 ( .A(n16182), .ZN(n9825) );
  INV_X1 U11429 ( .A(n10727), .ZN(n11013) );
  INV_X1 U11430 ( .A(n15869), .ZN(n18627) );
  OAI221_X1 U11431 ( .B1(n15853), .B2(n17416), .C1(n15853), .C2(n18193), .A(
        n15849), .ZN(n15963) );
  AOI21_X1 U11432 ( .B1(n17626), .B2(n12837), .A(n12788), .ZN(n12789) );
  NAND2_X1 U11433 ( .A1(n11825), .A2(n9734), .ZN(n11830) );
  OR2_X1 U11434 ( .A1(n11826), .A2(n11836), .ZN(n9734) );
  AND2_X1 U11435 ( .A1(n9733), .A2(n9732), .ZN(n11831) );
  NAND2_X1 U11436 ( .A1(n11827), .A2(n11828), .ZN(n9733) );
  NAND2_X1 U11437 ( .A1(n11847), .A2(n11829), .ZN(n9732) );
  NAND2_X1 U11439 ( .A1(n10388), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10389) );
  AOI22_X1 U11440 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19179), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10393) );
  NAND2_X1 U11441 ( .A1(n10248), .A2(n10247), .ZN(n10290) );
  NAND2_X1 U11442 ( .A1(n11796), .A2(n11795), .ZN(n11807) );
  AND2_X1 U11443 ( .A1(n20211), .A2(n11668), .ZN(n9853) );
  AND4_X1 U11444 ( .A1(n11339), .A2(n11338), .A3(n11337), .A4(n11336), .ZN(
        n11344) );
  NAND2_X1 U11445 ( .A1(n9849), .A2(n9848), .ZN(n11581) );
  AOI21_X1 U11446 ( .B1(n9851), .B2(n11530), .A(n11742), .ZN(n9848) );
  AOI21_X1 U11447 ( .B1(n11531), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n9852), 
        .ZN(n9851) );
  CLKBUF_X1 U11448 ( .A(n11543), .Z(n11592) );
  NAND2_X1 U11449 ( .A1(n11536), .A2(n11476), .ZN(n11422) );
  NAND2_X1 U11450 ( .A1(n11638), .A2(n11637), .ZN(n11837) );
  NAND2_X1 U11451 ( .A1(n9728), .A2(n9727), .ZN(n9726) );
  INV_X1 U11452 ( .A(n11844), .ZN(n9727) );
  NAND2_X1 U11453 ( .A1(n9735), .A2(n9729), .ZN(n9728) );
  AOI21_X1 U11454 ( .B1(n10533), .B2(n10530), .A(n10529), .ZN(n10539) );
  AND2_X1 U11455 ( .A1(n10528), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10529) );
  XNOR2_X1 U11456 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10538) );
  NOR2_X1 U11457 ( .A1(n10687), .A2(n9900), .ZN(n9899) );
  INV_X1 U11458 ( .A(n10676), .ZN(n9900) );
  INV_X1 U11459 ( .A(n11086), .ZN(n10546) );
  OAI21_X1 U11460 ( .B1(n10278), .B2(n16363), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10279) );
  NAND2_X1 U11461 ( .A1(n10350), .A2(n13963), .ZN(n10357) );
  AND2_X1 U11462 ( .A1(n10375), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10175) );
  NOR2_X1 U11463 ( .A1(n12564), .A2(n16905), .ZN(n12691) );
  NAND2_X1 U11464 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18637), .ZN(
        n12674) );
  OR2_X1 U11465 ( .A1(n13285), .A2(n20741), .ZN(n12513) );
  INV_X1 U11466 ( .A(n12496), .ZN(n12450) );
  NOR2_X1 U11467 ( .A1(n10004), .A2(n14695), .ZN(n10003) );
  INV_X1 U11468 ( .A(n10006), .ZN(n10004) );
  NOR2_X1 U11469 ( .A1(n11787), .A2(n20744), .ZN(n12496) );
  NOR2_X1 U11470 ( .A1(n14787), .A2(n9997), .ZN(n9996) );
  INV_X1 U11471 ( .A(n14734), .ZN(n9997) );
  AND2_X1 U11472 ( .A1(n12519), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12036) );
  NAND2_X1 U11473 ( .A1(n9880), .A2(n14637), .ZN(n9879) );
  INV_X1 U11474 ( .A(n14661), .ZN(n9880) );
  NAND2_X1 U11475 ( .A1(n14943), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11769) );
  NAND2_X1 U11476 ( .A1(n15001), .A2(n11765), .ZN(n9856) );
  NAND2_X1 U11477 ( .A1(n11766), .A2(n11765), .ZN(n9857) );
  NAND2_X1 U11478 ( .A1(n9870), .A2(n14697), .ZN(n9869) );
  INV_X1 U11479 ( .A(n14779), .ZN(n9870) );
  NAND2_X1 U11480 ( .A1(n14979), .A2(n11756), .ZN(n14967) );
  INV_X1 U11481 ( .A(n11959), .ZN(n11946) );
  NAND2_X1 U11482 ( .A1(n15131), .A2(n11755), .ZN(n9847) );
  NOR2_X1 U11483 ( .A1(n9872), .A2(n14336), .ZN(n9871) );
  INV_X1 U11484 ( .A(n14214), .ZN(n9872) );
  OR2_X1 U11485 ( .A1(n11516), .A2(n11515), .ZN(n11745) );
  INV_X1 U11486 ( .A(n12465), .ZN(n11471) );
  INV_X1 U11487 ( .A(n14111), .ZN(n11470) );
  NAND2_X1 U11488 ( .A1(n12464), .A2(n11745), .ZN(n11534) );
  XNOR2_X1 U11489 ( .A(n11581), .B(n11579), .ZN(n12005) );
  INV_X1 U11490 ( .A(n13429), .ZN(n11562) );
  XNOR2_X1 U11491 ( .A(n11615), .B(n11614), .ZN(n11616) );
  OAI22_X1 U11492 ( .A1(n13475), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11622), 
        .B2(n11637), .ZN(n11615) );
  NAND2_X1 U11493 ( .A1(n11591), .A2(n11590), .ZN(n11599) );
  INV_X1 U11494 ( .A(n11589), .ZN(n11590) );
  NAND2_X1 U11495 ( .A1(n11632), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11591) );
  OAI21_X1 U11496 ( .B1(n20071), .B2(n13464), .A(n11588), .ZN(n11589) );
  CLKBUF_X1 U11498 ( .A(n11500), .Z(n11501) );
  NAND2_X1 U11499 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n9944) );
  AND2_X1 U11500 ( .A1(n13736), .A2(n9890), .ZN(n9889) );
  NOR2_X1 U11501 ( .A1(n10545), .A2(n9893), .ZN(n10622) );
  NAND2_X1 U11502 ( .A1(n10571), .A2(n9894), .ZN(n9893) );
  INV_X1 U11503 ( .A(n13566), .ZN(n10049) );
  OR2_X1 U11504 ( .A1(n13055), .A2(n13056), .ZN(n10130) );
  INV_X1 U11505 ( .A(n15214), .ZN(n10028) );
  NOR2_X1 U11506 ( .A1(n15235), .A2(n10030), .ZN(n10029) );
  INV_X1 U11507 ( .A(n15382), .ZN(n10030) );
  AND2_X1 U11508 ( .A1(n15270), .A2(n15661), .ZN(n10033) );
  NOR2_X1 U11509 ( .A1(n11114), .A2(n10026), .ZN(n10025) );
  INV_X1 U11510 ( .A(n14350), .ZN(n10026) );
  NOR2_X1 U11511 ( .A1(n15432), .A2(n9928), .ZN(n9927) );
  OR2_X1 U11512 ( .A1(n9944), .A2(n15542), .ZN(n9943) );
  AND2_X1 U11513 ( .A1(n10763), .A2(n9763), .ZN(n9761) );
  AND4_X1 U11514 ( .A1(n10520), .A2(n10519), .A3(n10518), .A4(n10517), .ZN(
        n10521) );
  NOR2_X2 U11515 ( .A1(n11305), .A2(n15180), .ZN(n13169) );
  NOR2_X1 U11516 ( .A1(n10018), .A2(n15733), .ZN(n10017) );
  INV_X1 U11517 ( .A(n14241), .ZN(n10018) );
  INV_X1 U11518 ( .A(n14039), .ZN(n10019) );
  INV_X1 U11519 ( .A(n13743), .ZN(n10046) );
  INV_X1 U11520 ( .A(n13605), .ZN(n10045) );
  NOR2_X1 U11521 ( .A1(n12884), .A2(n14302), .ZN(n12867) );
  INV_X1 U11522 ( .A(n10972), .ZN(n11027) );
  INV_X1 U11523 ( .A(n19816), .ZN(n19268) );
  NAND2_X1 U11524 ( .A1(n10183), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9956) );
  NOR2_X1 U11525 ( .A1(n16928), .A2(n12652), .ZN(n12651) );
  NAND2_X1 U11526 ( .A1(n16876), .A2(n17474), .ZN(n9911) );
  AND2_X1 U11529 ( .A1(n12719), .A2(n10058), .ZN(n10057) );
  NAND2_X1 U11530 ( .A1(n17763), .A2(n9640), .ZN(n12784) );
  AND2_X1 U11531 ( .A1(n12776), .A2(n12803), .ZN(n12777) );
  INV_X1 U11532 ( .A(n12739), .ZN(n10065) );
  AND2_X1 U11533 ( .A1(n17812), .A2(n10065), .ZN(n10063) );
  XNOR2_X1 U11534 ( .A(n12813), .B(n12811), .ZN(n12726) );
  CLKBUF_X1 U11535 ( .A(n11788), .Z(n11789) );
  AND2_X1 U11536 ( .A1(n20738), .A2(n14090), .ZN(n19972) );
  NAND2_X1 U11537 ( .A1(n19942), .A2(n19948), .ZN(n19888) );
  OR2_X1 U11538 ( .A1(n19972), .A2(n12409), .ZN(n14112) );
  AND3_X1 U11539 ( .A1(n11494), .A2(n11503), .A3(n10124), .ZN(n11505) );
  INV_X1 U11540 ( .A(n12453), .ZN(n12539) );
  INV_X1 U11541 ( .A(n12110), .ZN(n12538) );
  OAI22_X1 U11542 ( .A1(n12512), .A2(n12513), .B1(n15936), .B2(n13286), .ZN(
        n13447) );
  AND2_X1 U11543 ( .A1(n10000), .A2(n14334), .ZN(n9999) );
  NOR2_X1 U11544 ( .A1(n10009), .A2(n12461), .ZN(n10008) );
  OR2_X1 U11545 ( .A1(n10011), .A2(n10010), .ZN(n10009) );
  INV_X1 U11546 ( .A(n14601), .ZN(n10010) );
  NOR2_X1 U11547 ( .A1(n12302), .A2(n12301), .ZN(n12303) );
  OR2_X1 U11548 ( .A1(n12284), .A2(n14832), .ZN(n12302) );
  AND2_X1 U11549 ( .A1(n12033), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12045) );
  NAND2_X1 U11550 ( .A1(n9875), .A2(n9877), .ZN(n9874) );
  AND2_X1 U11551 ( .A1(n14574), .A2(n12468), .ZN(n9877) );
  AND2_X1 U11552 ( .A1(n14591), .A2(n14574), .ZN(n14576) );
  NOR2_X1 U11553 ( .A1(n14616), .A2(n9873), .ZN(n14591) );
  INV_X1 U11554 ( .A(n9875), .ZN(n9873) );
  OR2_X1 U11555 ( .A1(n14626), .A2(n14614), .ZN(n14616) );
  NOR2_X1 U11556 ( .A1(n14616), .A2(n14602), .ZN(n14604) );
  NOR2_X1 U11557 ( .A1(n9739), .A2(n16071), .ZN(n9738) );
  INV_X1 U11558 ( .A(n15088), .ZN(n9739) );
  OR2_X1 U11559 ( .A1(n9659), .A2(n14670), .ZN(n14672) );
  AND2_X1 U11560 ( .A1(n11928), .A2(n11927), .ZN(n14683) );
  NOR3_X1 U11561 ( .A1(n14780), .A2(n14713), .A3(n14779), .ZN(n14712) );
  OR2_X1 U11562 ( .A1(n14791), .A2(n14726), .ZN(n14780) );
  AND2_X1 U11563 ( .A1(n16132), .A2(n11902), .ZN(n14215) );
  NAND2_X1 U11564 ( .A1(n14558), .A2(n20744), .ZN(n13464) );
  NAND2_X1 U11565 ( .A1(n9865), .A2(n9862), .ZN(n9861) );
  OR2_X1 U11566 ( .A1(n11960), .A2(n9864), .ZN(n9865) );
  INV_X1 U11567 ( .A(n9863), .ZN(n9862) );
  OAI22_X1 U11568 ( .A1(n13404), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n11956), .B2(P1_EBX_REG_1__SCAN_IN), .ZN(n9863) );
  NOR2_X1 U11570 ( .A1(n9721), .A2(n9601), .ZN(n11987) );
  AOI21_X1 U11571 ( .B1(n11852), .B2(n9722), .A(n19862), .ZN(n9721) );
  NAND2_X1 U11572 ( .A1(n11597), .A2(n20502), .ZN(n13429) );
  AND4_X1 U11573 ( .A1(n11399), .A2(n11398), .A3(n11397), .A4(n11396), .ZN(
        n11400) );
  AND4_X1 U11574 ( .A1(n11385), .A2(n11384), .A3(n11383), .A4(n11382), .ZN(
        n11403) );
  OR2_X1 U11575 ( .A1(n9595), .A2(n12013), .ZN(n20505) );
  AND2_X1 U11576 ( .A1(n20394), .A2(n20216), .ZN(n20543) );
  OR2_X1 U11577 ( .A1(n11999), .A2(n20058), .ZN(n20580) );
  NAND2_X1 U11578 ( .A1(n9748), .A2(n11851), .ZN(n13444) );
  NAND2_X1 U11579 ( .A1(n11848), .A2(n9749), .ZN(n9748) );
  AOI21_X1 U11580 ( .B1(n9752), .B2(n9662), .A(n9750), .ZN(n9749) );
  INV_X2 U11581 ( .A(n11475), .ZN(n15926) );
  AOI221_X1 U11582 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10710), 
        .C1(n15860), .C2(n10710), .A(n10709), .ZN(n10999) );
  INV_X1 U11583 ( .A(n9947), .ZN(n9946) );
  OAI21_X1 U11584 ( .B1(n9951), .B2(n9948), .A(n9950), .ZN(n9947) );
  NOR2_X1 U11585 ( .A1(n15204), .A2(n10893), .ZN(n10901) );
  NAND2_X1 U11586 ( .A1(n15224), .A2(n15202), .ZN(n15204) );
  NOR2_X1 U11587 ( .A1(n9634), .A2(n9896), .ZN(n15203) );
  NAND2_X1 U11588 ( .A1(n15301), .A2(n9897), .ZN(n9896) );
  NOR2_X1 U11589 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(P2_EBX_REG_26__SCAN_IN), 
        .ZN(n9897) );
  NOR2_X2 U11590 ( .A1(n10662), .A2(n10661), .ZN(n10672) );
  OAI22_X1 U11591 ( .A1(n13186), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n13325), 
        .B2(n10855), .ZN(n13207) );
  AND2_X1 U11592 ( .A1(n12887), .A2(n13564), .ZN(n12888) );
  AND2_X1 U11593 ( .A1(n12886), .A2(n13571), .ZN(n13563) );
  NAND2_X1 U11594 ( .A1(n10322), .A2(n10321), .ZN(n10779) );
  NAND2_X1 U11595 ( .A1(n9801), .A2(n9803), .ZN(n9800) );
  INV_X1 U11596 ( .A(n11307), .ZN(n11309) );
  AND2_X1 U11597 ( .A1(n9988), .A2(n9986), .ZN(n9985) );
  INV_X1 U11598 ( .A(n15320), .ZN(n9986) );
  NOR2_X1 U11599 ( .A1(n10023), .A2(n11085), .ZN(n10022) );
  INV_X1 U11600 ( .A(n13822), .ZN(n10023) );
  INV_X1 U11601 ( .A(n18863), .ZN(n13220) );
  NAND2_X1 U11602 ( .A1(n10274), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13324) );
  NAND2_X1 U11603 ( .A1(n16340), .A2(n13297), .ZN(n13322) );
  AND2_X1 U11604 ( .A1(n9611), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9934) );
  INV_X1 U11605 ( .A(n13714), .ZN(n10796) );
  NAND2_X1 U11606 ( .A1(n10039), .A2(n13583), .ZN(n13715) );
  AOI21_X1 U11607 ( .B1(n10957), .B2(n10897), .A(n9882), .ZN(n10898) );
  OAI21_X1 U11608 ( .B1(n9885), .B2(n9884), .A(n9883), .ZN(n9882) );
  NAND2_X1 U11609 ( .A1(n10866), .A2(n10087), .ZN(n10080) );
  OR2_X1 U11610 ( .A1(n10081), .A2(n10084), .ZN(n10079) );
  OR2_X1 U11611 ( .A1(n10873), .A2(n15640), .ZN(n15494) );
  NAND2_X1 U11612 ( .A1(n10083), .A2(n10084), .ZN(n10078) );
  AND2_X1 U11613 ( .A1(n10101), .A2(n10112), .ZN(n9776) );
  AND2_X1 U11614 ( .A1(n10102), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10101) );
  INV_X1 U11615 ( .A(n10102), .ZN(n10100) );
  NAND2_X1 U11616 ( .A1(n15539), .A2(n10856), .ZN(n9813) );
  AND2_X1 U11617 ( .A1(n9816), .A2(n15527), .ZN(n9815) );
  NAND2_X1 U11618 ( .A1(n15540), .A2(n10856), .ZN(n9816) );
  NAND2_X1 U11619 ( .A1(n10019), .A2(n10016), .ZN(n15718) );
  AND2_X1 U11620 ( .A1(n10017), .A2(n15716), .ZN(n10016) );
  NAND2_X1 U11621 ( .A1(n9671), .A2(n10857), .ZN(n9821) );
  OAI21_X1 U11622 ( .B1(n9825), .B2(n9820), .A(n9818), .ZN(n15548) );
  INV_X1 U11623 ( .A(n9821), .ZN(n9820) );
  AOI21_X1 U11624 ( .B1(n9823), .B2(n9821), .A(n9819), .ZN(n9818) );
  INV_X1 U11625 ( .A(n15549), .ZN(n9819) );
  NAND2_X1 U11626 ( .A1(n10019), .A2(n10017), .ZN(n14242) );
  NAND2_X1 U11627 ( .A1(n10086), .A2(n15742), .ZN(n16182) );
  AND2_X1 U11628 ( .A1(n15761), .A2(n10092), .ZN(n9798) );
  NAND3_X1 U11629 ( .A1(n10757), .A2(n10756), .A3(n10755), .ZN(n14313) );
  NAND2_X1 U11630 ( .A1(n14313), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14312) );
  NOR2_X1 U11631 ( .A1(n19128), .A2(n19126), .ZN(n9833) );
  AND2_X1 U11632 ( .A1(n11016), .A2(n11015), .ZN(n16334) );
  XNOR2_X1 U11633 ( .A(n13968), .B(n12867), .ZN(n13384) );
  NAND2_X1 U11634 ( .A1(n19795), .A2(n18986), .ZN(n19327) );
  INV_X1 U11635 ( .A(n10579), .ZN(n19300) );
  NOR2_X1 U11636 ( .A1(n19796), .A2(n19327), .ZN(n19332) );
  NAND2_X1 U11637 ( .A1(n19795), .A2(n19825), .ZN(n19367) );
  NOR2_X1 U11638 ( .A1(n19795), .A2(n19825), .ZN(n19611) );
  OR2_X1 U11639 ( .A1(n19795), .A2(n18986), .ZN(n19584) );
  AOI21_X2 U11640 ( .B1(n16359), .B2(n14273), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19662) );
  INV_X1 U11641 ( .A(n19662), .ZN(n19363) );
  NOR2_X1 U11642 ( .A1(n13257), .A2(n13256), .ZN(n18622) );
  NOR2_X1 U11643 ( .A1(n16610), .A2(n16611), .ZN(n16609) );
  INV_X1 U11645 ( .A(n17533), .ZN(n9921) );
  NOR2_X1 U11646 ( .A1(n16653), .A2(n17540), .ZN(n16652) );
  NOR2_X1 U11647 ( .A1(n17007), .A2(n16982), .ZN(n15820) );
  AOI21_X1 U11648 ( .B1(n15848), .B2(n18627), .A(n9790), .ZN(n15961) );
  AND2_X1 U11649 ( .A1(n14482), .A2(n14481), .ZN(n9790) );
  NOR2_X1 U11650 ( .A1(n17575), .A2(n17574), .ZN(n17551) );
  NOR2_X1 U11651 ( .A1(n17613), .A2(n17612), .ZN(n17587) );
  NOR2_X1 U11652 ( .A1(n17678), .A2(n9902), .ZN(n17634) );
  NAND2_X1 U11653 ( .A1(n17656), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9902) );
  NAND3_X1 U11654 ( .A1(n17746), .A2(n17718), .A3(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17678) );
  INV_X1 U11655 ( .A(n17521), .ZN(n17529) );
  NOR2_X1 U11656 ( .A1(n12793), .A2(n12792), .ZN(n17619) );
  NAND2_X1 U11657 ( .A1(n17672), .A2(n12783), .ZN(n12793) );
  NAND2_X1 U11658 ( .A1(n9715), .A2(n17672), .ZN(n17626) );
  NOR2_X1 U11659 ( .A1(n9717), .A2(n9716), .ZN(n9715) );
  INV_X1 U11660 ( .A(n12783), .ZN(n9716) );
  OR2_X1 U11661 ( .A1(n17689), .A2(n17627), .ZN(n17672) );
  NAND2_X1 U11662 ( .A1(n17624), .A2(n17627), .ZN(n10069) );
  NAND2_X1 U11663 ( .A1(n10068), .A2(n17624), .ZN(n17750) );
  NAND2_X1 U11664 ( .A1(n9718), .A2(n17784), .ZN(n17775) );
  OAI21_X1 U11665 ( .B1(n17783), .B2(n17785), .A(n17786), .ZN(n9718) );
  NOR2_X1 U11666 ( .A1(n18624), .A2(n15872), .ZN(n15870) );
  INV_X1 U11667 ( .A(n18622), .ZN(n15865) );
  NOR2_X1 U11668 ( .A1(n12588), .A2(n12587), .ZN(n15862) );
  NOR2_X1 U11669 ( .A1(n17813), .A2(n17812), .ZN(n17811) );
  INV_X1 U11670 ( .A(n12671), .ZN(n18219) );
  AOI22_X1 U11671 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12576) );
  AOI22_X1 U11672 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12703), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12577) );
  NOR2_X1 U11673 ( .A1(n18688), .A2(n18690), .ZN(n18679) );
  INV_X1 U11674 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20499) );
  CLKBUF_X1 U11675 ( .A(n13429), .Z(n20537) );
  CLKBUF_X1 U11676 ( .A(n13475), .Z(n13476) );
  NAND2_X1 U11677 ( .A1(n10979), .A2(n10729), .ZN(n18865) );
  NAND2_X1 U11678 ( .A1(n15176), .A2(n15175), .ZN(n15573) );
  AND2_X1 U11679 ( .A1(n15316), .A2(n10252), .ZN(n15342) );
  INV_X1 U11680 ( .A(n9969), .ZN(n9968) );
  OAI22_X1 U11681 ( .A1(n15277), .A2(n9972), .B1(n13126), .B2(n9973), .ZN(
        n9969) );
  AND2_X1 U11682 ( .A1(n13378), .A2(n14276), .ZN(n19011) );
  AND2_X1 U11683 ( .A1(n16265), .A2(n19814), .ZN(n19117) );
  AND2_X1 U11684 ( .A1(n16265), .A2(n13308), .ZN(n16255) );
  AND2_X2 U11685 ( .A1(n10348), .A2(n10332), .ZN(n15792) );
  NOR2_X2 U11686 ( .A1(n18865), .A2(n10383), .ZN(n19121) );
  INV_X1 U11687 ( .A(n9780), .ZN(n9779) );
  OAI21_X1 U11688 ( .B1(n19004), .B2(n19143), .A(n10014), .ZN(n9780) );
  OR2_X1 U11689 ( .A1(n15276), .A2(n19138), .ZN(n10014) );
  NAND2_X1 U11690 ( .A1(n9770), .A2(n10855), .ZN(n9767) );
  NAND2_X1 U11691 ( .A1(n9769), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9768) );
  AOI21_X1 U11692 ( .B1(n15419), .B2(n16302), .A(n15420), .ZN(n9837) );
  INV_X1 U11693 ( .A(n9885), .ZN(n10959) );
  NAND2_X1 U11694 ( .A1(n11010), .A2(n11012), .ZN(n12855) );
  OR2_X1 U11695 ( .A1(n11011), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11012) );
  NAND2_X1 U11696 ( .A1(n9806), .A2(n9804), .ZN(n10707) );
  AOI21_X1 U11697 ( .B1(n9613), .B2(n9811), .A(n9805), .ZN(n9804) );
  INV_X1 U11698 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19828) );
  OR2_X1 U11699 ( .A1(n19804), .A2(n19816), .ZN(n19796) );
  NAND2_X1 U11700 ( .A1(n13537), .A2(n13540), .ZN(n19795) );
  OR2_X1 U11701 ( .A1(n13538), .A2(n13539), .ZN(n13540) );
  INV_X1 U11702 ( .A(n16917), .ZN(n16878) );
  INV_X1 U11703 ( .A(n16881), .ZN(n16916) );
  NAND2_X1 U11705 ( .A1(n18632), .A2(n17202), .ZN(n17350) );
  OR2_X1 U11706 ( .A1(n12843), .A2(n12842), .ZN(n12844) );
  NOR2_X1 U11707 ( .A1(n16407), .A2(n9712), .ZN(n9711) );
  OAI21_X1 U11708 ( .B1(n16405), .B2(n16406), .A(n9713), .ZN(n9712) );
  NOR2_X2 U11709 ( .A1(n17847), .A2(n17321), .ZN(n17738) );
  NAND2_X1 U11710 ( .A1(n12802), .A2(n16379), .ZN(n15952) );
  OR2_X1 U11711 ( .A1(n12801), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12802) );
  XNOR2_X1 U11712 ( .A(n9714), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16404) );
  AOI21_X1 U11713 ( .B1(n15874), .B2(n15873), .A(n16426), .ZN(n9714) );
  NAND2_X1 U11714 ( .A1(n9759), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11816) );
  NAND2_X1 U11715 ( .A1(n9731), .A2(n9730), .ZN(n9729) );
  NAND2_X1 U11716 ( .A1(n11849), .A2(n11829), .ZN(n9730) );
  NAND2_X1 U11717 ( .A1(n11830), .A2(n11831), .ZN(n9731) );
  NAND2_X1 U11718 ( .A1(n11833), .A2(n11832), .ZN(n9735) );
  AND4_X1 U11719 ( .A1(n10473), .A2(n10472), .A3(n10471), .A4(n10470), .ZN(
        n10486) );
  INV_X1 U11720 ( .A(n11819), .ZN(n11809) );
  NAND2_X1 U11721 ( .A1(n11474), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11543) );
  OR2_X1 U11722 ( .A1(n11716), .A2(n11715), .ZN(n11732) );
  OR2_X1 U11723 ( .A1(n11693), .A2(n11692), .ZN(n11721) );
  OR2_X1 U11724 ( .A1(n11667), .A2(n11666), .ZN(n11676) );
  OR2_X1 U11725 ( .A1(n11560), .A2(n11559), .ZN(n11620) );
  INV_X1 U11726 ( .A(n9754), .ZN(n11970) );
  AOI21_X1 U11727 ( .B1(n14092), .B2(n11968), .A(n9841), .ZN(n11969) );
  OR2_X1 U11728 ( .A1(n11648), .A2(n11647), .ZN(n11672) );
  NOR2_X1 U11729 ( .A1(n10252), .A2(n10038), .ZN(n10037) );
  NAND2_X1 U11730 ( .A1(n10323), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9765) );
  NAND2_X1 U11731 ( .A1(n10677), .A2(n10676), .ZN(n10688) );
  AOI22_X1 U11732 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19239), .B1(
        n10469), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10392) );
  NAND2_X1 U11733 ( .A1(n9598), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10293) );
  NAND2_X1 U11734 ( .A1(n10260), .A2(n10259), .ZN(n10297) );
  NAND2_X1 U11735 ( .A1(n10251), .A2(n10214), .ZN(n10215) );
  AOI21_X1 U11736 ( .B1(n9587), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n10178), .ZN(n10179) );
  AND2_X1 U11737 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10178) );
  NAND2_X1 U11738 ( .A1(n15828), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10058) );
  NOR2_X1 U11739 ( .A1(n17328), .A2(n12763), .ZN(n12776) );
  NOR2_X1 U11740 ( .A1(n12546), .A2(n12674), .ZN(n12547) );
  NAND2_X1 U11741 ( .A1(n18215), .A2(n18219), .ZN(n12661) );
  AND2_X1 U11742 ( .A1(n10001), .A2(n14327), .ZN(n10000) );
  CLKBUF_X1 U11743 ( .A(n11481), .Z(n11482) );
  NOR2_X1 U11744 ( .A1(n12220), .A2(n14700), .ZN(n12250) );
  NOR2_X1 U11745 ( .A1(n14777), .A2(n10007), .ZN(n10006) );
  INV_X1 U11746 ( .A(n14709), .ZN(n10007) );
  NOR2_X1 U11747 ( .A1(n9876), .A2(n14602), .ZN(n9875) );
  INV_X1 U11748 ( .A(n14589), .ZN(n9876) );
  NAND2_X1 U11749 ( .A1(n14911), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11771) );
  NAND2_X1 U11750 ( .A1(n11875), .A2(n11938), .ZN(n11956) );
  INV_X1 U11751 ( .A(n13453), .ZN(n9723) );
  INV_X1 U11752 ( .A(n11853), .ZN(n9724) );
  NAND2_X1 U11753 ( .A1(n11583), .A2(n11582), .ZN(n11617) );
  OR2_X1 U11754 ( .A1(n11581), .A2(n11580), .ZN(n11582) );
  INV_X1 U11756 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9839) );
  AND2_X1 U11757 ( .A1(n11601), .A2(n11600), .ZN(n11631) );
  AND4_X1 U11758 ( .A1(n11426), .A2(n11425), .A3(n11424), .A4(n11423), .ZN(
        n11441) );
  AND2_X1 U11759 ( .A1(n20424), .A2(n11587), .ZN(n20071) );
  CLKBUF_X1 U11760 ( .A(n11784), .Z(n11785) );
  AND2_X1 U11761 ( .A1(n13457), .A2(n13456), .ZN(n13665) );
  INV_X1 U11762 ( .A(n11849), .ZN(n9752) );
  NAND2_X1 U11763 ( .A1(n9726), .A2(n9725), .ZN(n11845) );
  AND2_X1 U11764 ( .A1(n11843), .A2(n11842), .ZN(n9725) );
  AOI21_X1 U11765 ( .B1(n11801), .B2(n11800), .A(n11799), .ZN(n11815) );
  NOR2_X1 U11766 ( .A1(n10193), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10195) );
  NAND2_X1 U11767 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19828), .ZN(
        n10711) );
  AND3_X1 U11768 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10710), .A3(
        n15860), .ZN(n10723) );
  OR2_X1 U11769 ( .A1(n10541), .A2(n10540), .ZN(n10991) );
  NAND2_X1 U11771 ( .A1(n9949), .A2(n13215), .ZN(n9950) );
  INV_X1 U11772 ( .A(n15443), .ZN(n9948) );
  INV_X1 U11773 ( .A(n9951), .ZN(n9949) );
  NAND2_X1 U11774 ( .A1(n10677), .A2(n9691), .ZN(n10871) );
  NAND2_X1 U11775 ( .A1(n10677), .A2(n9899), .ZN(n10696) );
  NAND2_X1 U11776 ( .A1(n10672), .A2(n14074), .ZN(n10675) );
  NAND2_X1 U11777 ( .A1(n9891), .A2(n9889), .ZN(n10642) );
  AND2_X1 U11778 ( .A1(n10056), .A2(n10055), .ZN(n10054) );
  INV_X1 U11779 ( .A(n15174), .ZN(n10055) );
  AND2_X1 U11780 ( .A1(n11287), .A2(n11046), .ZN(n10056) );
  OR2_X1 U11781 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10717), .ZN(
        n11180) );
  NOR2_X1 U11782 ( .A1(n10052), .A2(n13572), .ZN(n10051) );
  INV_X1 U11783 ( .A(n13727), .ZN(n10052) );
  INV_X1 U11784 ( .A(n13697), .ZN(n10050) );
  OR2_X1 U11785 ( .A1(n10308), .A2(n10307), .ZN(n10315) );
  NAND2_X1 U11786 ( .A1(n10332), .A2(n10316), .ZN(n9801) );
  AND2_X1 U11787 ( .A1(n10159), .A2(n10158), .ZN(n10162) );
  INV_X1 U11788 ( .A(n15295), .ZN(n9978) );
  NOR3_X1 U11789 ( .A1(n9989), .A2(n13035), .A3(n15307), .ZN(n13036) );
  AND2_X1 U11790 ( .A1(n12902), .A2(n9699), .ZN(n9982) );
  AND2_X1 U11791 ( .A1(n10022), .A2(n13997), .ZN(n10021) );
  NOR2_X1 U11792 ( .A1(n10269), .A2(n10972), .ZN(n11020) );
  NOR2_X1 U11793 ( .A1(n10841), .A2(n9936), .ZN(n9935) );
  INV_X1 U11794 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n9936) );
  INV_X1 U11795 ( .A(n15266), .ZN(n10042) );
  NOR2_X1 U11796 ( .A1(n9665), .A2(n9930), .ZN(n9929) );
  INV_X1 U11797 ( .A(n9932), .ZN(n9930) );
  NOR2_X1 U11798 ( .A1(n16227), .A2(n9933), .ZN(n9932) );
  INV_X1 U11799 ( .A(n13198), .ZN(n9931) );
  AND2_X1 U11800 ( .A1(n13582), .A2(n13613), .ZN(n10039) );
  AND2_X1 U11801 ( .A1(n10939), .A2(n10938), .ZN(n13181) );
  NOR2_X1 U11802 ( .A1(n15582), .A2(n11275), .ZN(n10109) );
  INV_X1 U11803 ( .A(n11043), .ZN(n9884) );
  NAND2_X1 U11804 ( .A1(n9773), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9772) );
  INV_X1 U11805 ( .A(n10103), .ZN(n9773) );
  NAND2_X1 U11806 ( .A1(n10104), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10103) );
  INV_X1 U11807 ( .A(n10105), .ZN(n10104) );
  OR2_X1 U11808 ( .A1(n10106), .A2(n15464), .ZN(n10105) );
  NAND2_X1 U11809 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10106) );
  AND2_X1 U11810 ( .A1(n10113), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10112) );
  NOR2_X1 U11811 ( .A1(n10772), .A2(n15698), .ZN(n10102) );
  NAND2_X1 U11812 ( .A1(n10771), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10772) );
  INV_X1 U11813 ( .A(n11230), .ZN(n11303) );
  INV_X1 U11814 ( .A(n11308), .ZN(n11302) );
  NOR2_X1 U11815 ( .A1(n10658), .A2(n9827), .ZN(n9826) );
  NOR2_X1 U11816 ( .A1(n10651), .A2(n16180), .ZN(n9827) );
  AND2_X1 U11817 ( .A1(n15731), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10113) );
  AND2_X1 U11818 ( .A1(n10093), .A2(n16213), .ZN(n10092) );
  AND2_X1 U11819 ( .A1(n10626), .A2(n9692), .ZN(n10093) );
  NAND2_X1 U11820 ( .A1(n10111), .A2(n10753), .ZN(n10760) );
  NAND2_X1 U11821 ( .A1(n9760), .A2(n10552), .ZN(n10744) );
  NAND2_X1 U11822 ( .A1(n9643), .A2(n10337), .ZN(n10095) );
  NAND2_X1 U11823 ( .A1(n13541), .A2(n10335), .ZN(n19359) );
  NOR2_X1 U11824 ( .A1(n9612), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9829) );
  NAND2_X1 U11825 ( .A1(n10188), .A2(n10192), .ZN(n9957) );
  AOI21_X1 U11826 ( .B1(n9590), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A(n10175), .ZN(n10177) );
  AND2_X1 U11827 ( .A1(n10375), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10203) );
  NAND3_X1 U11828 ( .A1(n19793), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19662), 
        .ZN(n14277) );
  AND2_X1 U11829 ( .A1(n12860), .A2(n10336), .ZN(n10335) );
  AOI21_X1 U11830 ( .B1(n17209), .B2(n12662), .A(n18200), .ZN(n12653) );
  NAND2_X1 U11831 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n12565), .ZN(
        n12563) );
  NAND2_X1 U11832 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18821), .ZN(
        n12568) );
  NOR2_X1 U11833 ( .A1(n12568), .A2(n12561), .ZN(n12599) );
  NAND2_X1 U11834 ( .A1(n18798), .A2(n18808), .ZN(n12566) );
  OR2_X1 U11835 ( .A1(n16905), .A2(n12567), .ZN(n12704) );
  NOR2_X1 U11836 ( .A1(n12566), .A2(n12563), .ZN(n12718) );
  INV_X1 U11837 ( .A(n12691), .ZN(n14457) );
  NAND2_X1 U11838 ( .A1(n12670), .A2(n16531), .ZN(n15847) );
  NOR2_X1 U11839 ( .A1(n17470), .A2(n17471), .ZN(n9924) );
  AND2_X1 U11840 ( .A1(n17476), .A2(n12799), .ZN(n10060) );
  NAND2_X1 U11841 ( .A1(n17488), .A2(n9687), .ZN(n16380) );
  INV_X1 U11842 ( .A(n17969), .ZN(n17850) );
  NOR2_X1 U11843 ( .A1(n17773), .A2(n12775), .ZN(n12779) );
  AND2_X1 U11844 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12774), .ZN(
        n12775) );
  INV_X1 U11845 ( .A(n12668), .ZN(n13254) );
  NOR2_X1 U11846 ( .A1(n12598), .A2(n12597), .ZN(n12652) );
  NOR2_X1 U11847 ( .A1(n12648), .A2(n12647), .ZN(n12657) );
  AND2_X1 U11848 ( .A1(n12174), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12190) );
  INV_X1 U11849 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n14364) );
  INV_X1 U11850 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19893) );
  NOR3_X1 U11851 ( .A1(n14672), .A2(n9675), .A3(n14661), .ZN(n14651) );
  OR2_X1 U11852 ( .A1(n13444), .A2(n13290), .ZN(n13454) );
  AND3_X1 U11853 ( .A1(n12079), .A2(n12078), .A3(n12077), .ZN(n14224) );
  AND2_X1 U11854 ( .A1(n13419), .A2(n13418), .ZN(n19998) );
  AOI22_X1 U11855 ( .A1(n12501), .A2(n12500), .B1(n14533), .B2(n12499), .ZN(
        n12536) );
  OR2_X1 U11856 ( .A1(n12457), .A2(n12456), .ZN(n14097) );
  AOI21_X1 U11857 ( .B1(n12499), .B2(n14578), .A(n12434), .ZN(n14573) );
  AOI21_X1 U11858 ( .B1(n12499), .B2(n14902), .A(n12393), .ZN(n14601) );
  NAND2_X1 U11859 ( .A1(n12371), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12373) );
  OAI22_X1 U11860 ( .A1(n12376), .A2(n12375), .B1(n12035), .B2(n14916), .ZN(
        n14613) );
  CLKBUF_X1 U11861 ( .A(n14611), .Z(n14612) );
  NAND2_X1 U11862 ( .A1(n12329), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12370) );
  NOR2_X1 U11863 ( .A1(n12298), .A2(n14956), .ZN(n12268) );
  AND2_X1 U11864 ( .A1(n12250), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12251) );
  NAND2_X1 U11865 ( .A1(n12251), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12298) );
  CLKBUF_X1 U11866 ( .A(n14644), .Z(n14645) );
  AND2_X1 U11867 ( .A1(n10003), .A2(n12235), .ZN(n10002) );
  OR2_X1 U11868 ( .A1(n12204), .A2(n14972), .ZN(n12220) );
  INV_X1 U11869 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14700) );
  NAND2_X1 U11870 ( .A1(n12190), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12204) );
  AND2_X1 U11871 ( .A1(n12157), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12174) );
  CLKBUF_X1 U11872 ( .A(n14723), .Z(n14724) );
  AND2_X1 U11873 ( .A1(n12142), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12157) );
  NOR2_X1 U11874 ( .A1(n12139), .A2(n15991), .ZN(n12142) );
  XNOR2_X1 U11875 ( .A(n14333), .B(n12126), .ZN(n14380) );
  NOR2_X1 U11876 ( .A1(n12095), .A2(n14364), .ZN(n12109) );
  NAND2_X1 U11877 ( .A1(n12091), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12095) );
  NOR2_X1 U11878 ( .A1(n12058), .A2(n19893), .ZN(n12091) );
  AOI21_X1 U11879 ( .B1(n12064), .B2(n12125), .A(n12063), .ZN(n14163) );
  AOI21_X1 U11880 ( .B1(n12057), .B2(n12125), .A(n12056), .ZN(n14066) );
  NAND2_X1 U11881 ( .A1(n12054), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12058) );
  AND2_X1 U11882 ( .A1(n12045), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12054) );
  NAND2_X1 U11883 ( .A1(n12053), .A2(n12052), .ZN(n13842) );
  AOI21_X1 U11884 ( .B1(n12043), .B2(n12125), .A(n12042), .ZN(n13805) );
  CLKBUF_X1 U11885 ( .A(n13778), .Z(n13779) );
  CLKBUF_X1 U11886 ( .A(n13803), .Z(n13804) );
  AND2_X1 U11887 ( .A1(n13444), .A2(n13280), .ZN(n13463) );
  OR2_X1 U11888 ( .A1(n9879), .A2(n14627), .ZN(n9878) );
  NOR2_X1 U11889 ( .A1(n15940), .A2(n9738), .ZN(n15076) );
  AND2_X1 U11890 ( .A1(n14961), .A2(n9700), .ZN(n9855) );
  NOR2_X1 U11891 ( .A1(n14672), .A2(n14661), .ZN(n15946) );
  OAI21_X1 U11892 ( .B1(n16092), .B2(n9747), .A(n9746), .ZN(n15096) );
  AND2_X1 U11893 ( .A1(n15118), .A2(n11989), .ZN(n9747) );
  AOI21_X1 U11894 ( .B1(n15121), .B2(n9690), .A(n15119), .ZN(n9746) );
  AND2_X1 U11895 ( .A1(n11931), .A2(n11930), .ZN(n14670) );
  OR3_X1 U11896 ( .A1(n14713), .A2(n9869), .A3(n9868), .ZN(n9867) );
  INV_X1 U11897 ( .A(n14683), .ZN(n9868) );
  NOR3_X1 U11898 ( .A1(n14780), .A2(n14713), .A3(n9869), .ZN(n14699) );
  AND2_X1 U11899 ( .A1(n14981), .A2(n11758), .ZN(n16033) );
  AND2_X1 U11900 ( .A1(n11920), .A2(n11919), .ZN(n14779) );
  NAND2_X1 U11901 ( .A1(n9847), .A2(n9846), .ZN(n9845) );
  OR2_X1 U11902 ( .A1(n11753), .A2(n16089), .ZN(n14981) );
  INV_X1 U11903 ( .A(n9847), .ZN(n14992) );
  NAND2_X1 U11904 ( .A1(n14215), .A2(n9666), .ZN(n14791) );
  AND2_X1 U11905 ( .A1(n14215), .A2(n9628), .ZN(n14789) );
  NAND2_X1 U11906 ( .A1(n14215), .A2(n9871), .ZN(n14382) );
  NAND2_X1 U11907 ( .A1(n14215), .A2(n14214), .ZN(n14335) );
  NOR2_X1 U11908 ( .A1(n16128), .A2(n11893), .ZN(n16132) );
  OR2_X1 U11909 ( .A1(n13772), .A2(n13771), .ZN(n16128) );
  NAND2_X1 U11910 ( .A1(n11628), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11629) );
  NOR2_X1 U11911 ( .A1(n9861), .A2(n9860), .ZN(n13549) );
  NOR2_X1 U11912 ( .A1(n13403), .A2(n11914), .ZN(n9860) );
  XNOR2_X1 U11913 ( .A(n11628), .B(n13554), .ZN(n13545) );
  INV_X1 U11914 ( .A(n13547), .ZN(n15119) );
  INV_X1 U11915 ( .A(n16098), .ZN(n15121) );
  NOR2_X1 U11916 ( .A1(n11987), .A2(n11980), .ZN(n13550) );
  NAND2_X2 U11917 ( .A1(n11879), .A2(n11938), .ZN(n13404) );
  OAI211_X1 U11918 ( .C1(n11814), .C2(n11535), .A(n11534), .B(n11533), .ZN(
        n11572) );
  INV_X1 U11919 ( .A(n12004), .ZN(n12007) );
  INV_X1 U11920 ( .A(n12005), .ZN(n12006) );
  NAND2_X1 U11921 ( .A1(n11636), .A2(n11635), .ZN(n20212) );
  CLKBUF_X1 U11923 ( .A(n11786), .Z(n11787) );
  CLKBUF_X1 U11924 ( .A(n13436), .Z(n13663) );
  INV_X1 U11925 ( .A(n20305), .ZN(n20714) );
  AND4_X1 U11926 ( .A1(n11370), .A2(n11369), .A3(n11368), .A4(n11367), .ZN(
        n11376) );
  AND3_X1 U11927 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20744), .A3(n20060), 
        .ZN(n20104) );
  INV_X1 U11928 ( .A(n11598), .ZN(n11547) );
  INV_X1 U11929 ( .A(n20580), .ZN(n20534) );
  AOI21_X1 U11930 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20499), .A(n20114), 
        .ZN(n20581) );
  AND2_X1 U11931 ( .A1(n14094), .A2(n14093), .ZN(n15925) );
  CLKBUF_X1 U11932 ( .A(n11866), .Z(n15927) );
  NAND2_X1 U11933 ( .A1(n10526), .A2(n10525), .ZN(n10982) );
  INV_X1 U11934 ( .A(n13176), .ZN(n16339) );
  INV_X1 U11935 ( .A(n15522), .ZN(n9953) );
  OR2_X1 U11936 ( .A1(n18921), .A2(n9951), .ZN(n9954) );
  AOI21_X1 U11937 ( .B1(n10890), .B2(n9888), .A(n9685), .ZN(n9886) );
  INV_X1 U11938 ( .A(n9889), .ZN(n9888) );
  NAND2_X1 U11939 ( .A1(n10642), .A2(n10890), .ZN(n13849) );
  OR2_X1 U11940 ( .A1(n10545), .A2(n9895), .ZN(n10548) );
  NAND2_X1 U11941 ( .A1(n18987), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18974) );
  AND2_X1 U11942 ( .A1(n12888), .A2(n9679), .ZN(n9992) );
  NOR2_X1 U11943 ( .A1(n13697), .A2(n10047), .ZN(n13735) );
  NAND2_X1 U11944 ( .A1(n9614), .A2(n10048), .ZN(n10047) );
  INV_X1 U11945 ( .A(n13733), .ZN(n10048) );
  AND2_X1 U11946 ( .A1(n10811), .A2(n10810), .ZN(n13566) );
  NAND2_X1 U11947 ( .A1(n10050), .A2(n10051), .ZN(n13726) );
  NOR2_X1 U11948 ( .A1(n13697), .A2(n13572), .ZN(n13728) );
  CLKBUF_X1 U11949 ( .A(n13561), .Z(n13562) );
  INV_X1 U11950 ( .A(n13144), .ZN(n9973) );
  NOR2_X1 U11951 ( .A1(n9971), .A2(n9973), .ZN(n9970) );
  INV_X1 U11952 ( .A(n15277), .ZN(n9971) );
  AND2_X2 U11953 ( .A1(n15247), .A2(n9688), .ZN(n11292) );
  INV_X1 U11954 ( .A(n11290), .ZN(n10027) );
  NAND2_X1 U11955 ( .A1(n9619), .A2(n9980), .ZN(n9976) );
  NAND2_X1 U11956 ( .A1(n15247), .A2(n9680), .ZN(n15216) );
  NAND2_X1 U11957 ( .A1(n15247), .A2(n10029), .ZN(n15237) );
  NAND2_X1 U11958 ( .A1(n9983), .A2(n9684), .ZN(n9987) );
  INV_X1 U11959 ( .A(n15325), .ZN(n9990) );
  AND2_X1 U11960 ( .A1(n10033), .A2(n10032), .ZN(n10031) );
  CLKBUF_X1 U11961 ( .A(n15323), .Z(n15324) );
  OR2_X1 U11962 ( .A1(n12955), .A2(n12954), .ZN(n15340) );
  OR2_X1 U11963 ( .A1(n12929), .A2(n12928), .ZN(n14170) );
  NAND2_X1 U11964 ( .A1(n10252), .A2(n11054), .ZN(n13161) );
  AND2_X1 U11965 ( .A1(n10025), .A2(n15778), .ZN(n10024) );
  NAND2_X1 U11966 ( .A1(n14351), .A2(n14350), .ZN(n14352) );
  OR2_X1 U11967 ( .A1(n16337), .A2(n13228), .ZN(n13275) );
  OR2_X1 U11968 ( .A1(n13227), .A2(n18863), .ZN(n13228) );
  INV_X1 U11969 ( .A(n13160), .ZN(n14278) );
  AND2_X1 U11970 ( .A1(n12849), .A2(n9695), .ZN(n10945) );
  NOR2_X1 U11971 ( .A1(n10954), .A2(n10953), .ZN(n11284) );
  OR2_X1 U11972 ( .A1(n15244), .A2(n15245), .ZN(n15310) );
  OR2_X1 U11973 ( .A1(n15310), .A2(n15309), .ZN(n15312) );
  AND2_X1 U11974 ( .A1(n14174), .A2(n10040), .ZN(n15337) );
  AND2_X1 U11975 ( .A1(n9660), .A2(n10041), .ZN(n10040) );
  INV_X1 U11976 ( .A(n15335), .ZN(n10041) );
  NAND2_X1 U11977 ( .A1(n14174), .A2(n9660), .ZN(n15336) );
  NAND2_X1 U11978 ( .A1(n9942), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9941) );
  INV_X1 U11979 ( .A(n9943), .ZN(n9942) );
  INV_X1 U11980 ( .A(n10112), .ZN(n9774) );
  INV_X1 U11981 ( .A(n15746), .ZN(n9775) );
  AND2_X1 U11982 ( .A1(n10821), .A2(n10820), .ZN(n13743) );
  NOR2_X1 U11983 ( .A1(n13605), .A2(n13743), .ZN(n13837) );
  OR2_X1 U11984 ( .A1(n10762), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9622) );
  INV_X1 U11985 ( .A(n13717), .ZN(n10801) );
  NAND2_X1 U11986 ( .A1(n10801), .A2(n10136), .ZN(n13697) );
  INV_X1 U11987 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18973) );
  AND2_X1 U11988 ( .A1(n10795), .A2(n10794), .ZN(n13714) );
  AND2_X1 U11989 ( .A1(n10783), .A2(n10117), .ZN(n13583) );
  INV_X1 U11990 ( .A(n14544), .ZN(n10904) );
  INV_X1 U11991 ( .A(n9770), .ZN(n9769) );
  NAND2_X1 U11992 ( .A1(n9771), .A2(n10107), .ZN(n9770) );
  NOR2_X1 U11993 ( .A1(n10108), .A2(n11311), .ZN(n10107) );
  INV_X1 U11994 ( .A(n9772), .ZN(n9771) );
  INV_X1 U11995 ( .A(n10109), .ZN(n10108) );
  NAND2_X1 U11996 ( .A1(n15193), .A2(n11094), .ZN(n9885) );
  OR3_X1 U11997 ( .A1(n15243), .A2(n10628), .A3(n15464), .ZN(n15459) );
  AND2_X1 U11998 ( .A1(n15337), .A2(n10845), .ZN(n15328) );
  INV_X1 U11999 ( .A(n15503), .ZN(n9805) );
  AND2_X1 U12000 ( .A1(n9661), .A2(n10044), .ZN(n10043) );
  INV_X1 U12001 ( .A(n13959), .ZN(n10044) );
  NAND2_X1 U12002 ( .A1(n10045), .A2(n9661), .ZN(n13958) );
  OR2_X1 U12003 ( .A1(n14253), .A2(n10666), .ZN(n15560) );
  AND2_X1 U12004 ( .A1(n9824), .A2(n9826), .ZN(n15563) );
  NAND2_X1 U12005 ( .A1(n9825), .A2(n16179), .ZN(n9824) );
  NAND2_X1 U12006 ( .A1(n10094), .A2(n10092), .ZN(n15760) );
  AND2_X1 U12007 ( .A1(n10094), .A2(n10093), .ZN(n16211) );
  OR2_X1 U12008 ( .A1(n14197), .A2(n11260), .ZN(n11261) );
  NAND2_X1 U12009 ( .A1(n9799), .A2(n10628), .ZN(n13811) );
  INV_X1 U12010 ( .A(n13816), .ZN(n9799) );
  INV_X1 U12011 ( .A(n10310), .ZN(n10313) );
  INV_X1 U12012 ( .A(n10311), .ZN(n10312) );
  AOI211_X1 U12013 ( .C1(n13305), .C2(n11224), .A(n11068), .B(n11053), .ZN(
        n13379) );
  NOR2_X1 U12014 ( .A1(n10038), .A2(n18988), .ZN(n10036) );
  NAND2_X1 U12015 ( .A1(n12860), .A2(n12859), .ZN(n9965) );
  OAI22_X1 U12016 ( .A1(n13383), .A2(n13384), .B1(n12867), .B2(n13968), .ZN(
        n13524) );
  AND3_X1 U12017 ( .A1(n11031), .A2(n11030), .A3(n11029), .ZN(n15801) );
  NAND2_X1 U12018 ( .A1(n11001), .A2(n11000), .ZN(n16340) );
  NAND2_X1 U12019 ( .A1(n10263), .A2(n19846), .ZN(n10965) );
  AND2_X1 U12020 ( .A1(n19804), .A2(n19268), .ZN(n19790) );
  OR2_X1 U12021 ( .A1(n10388), .A2(n19485), .ZN(n19492) );
  INV_X1 U12022 ( .A(n19547), .ZN(n19541) );
  NOR2_X2 U12023 ( .A1(n14278), .A2(n14277), .ZN(n19170) );
  NOR2_X2 U12024 ( .A1(n14276), .A2(n14277), .ZN(n19171) );
  INV_X1 U12025 ( .A(n19170), .ZN(n19162) );
  INV_X1 U12026 ( .A(n19171), .ZN(n19164) );
  NOR2_X1 U12027 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19840) );
  INV_X1 U12028 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19848) );
  NOR2_X1 U12029 ( .A1(n18185), .A2(n18842), .ZN(n12670) );
  OR2_X1 U12030 ( .A1(n15853), .A2(n13255), .ZN(n18621) );
  INV_X1 U12031 ( .A(n9909), .ZN(n9908) );
  OAI21_X1 U12032 ( .B1(n9919), .B2(n17497), .A(n9911), .ZN(n9909) );
  OR2_X1 U12033 ( .A1(n16673), .A2(n9905), .ZN(n9903) );
  OR2_X1 U12034 ( .A1(n17566), .A2(n17576), .ZN(n9905) );
  OR2_X1 U12035 ( .A1(n16876), .A2(n17566), .ZN(n9904) );
  OR2_X1 U12036 ( .A1(n16673), .A2(n17576), .ZN(n9906) );
  NOR2_X1 U12037 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16702), .ZN(n16694) );
  INV_X1 U12038 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16751) );
  INV_X1 U12039 ( .A(n13259), .ZN(n13260) );
  NOR2_X1 U12040 ( .A1(n18855), .A2(n17353), .ZN(n13259) );
  NAND4_X1 U12041 ( .A1(n18122), .A2(n18855), .A3(n18694), .A4(n18685), .ZN(
        n16807) );
  NAND2_X1 U12042 ( .A1(n17141), .A2(n9631), .ZN(n15835) );
  NOR2_X1 U12043 ( .A1(n17094), .A2(n9782), .ZN(n9781) );
  INV_X1 U12044 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n9782) );
  OR2_X1 U12045 ( .A1(n15961), .A2(n9788), .ZN(n17171) );
  NAND2_X1 U12046 ( .A1(n9789), .A2(n18185), .ZN(n9788) );
  INV_X1 U12047 ( .A(n14483), .ZN(n9789) );
  INV_X1 U12048 ( .A(n12723), .ZN(n10059) );
  NOR2_X1 U12049 ( .A1(n18219), .A2(n17209), .ZN(n18632) );
  AOI21_X1 U12050 ( .B1(n15847), .B2(n18681), .A(n18840), .ZN(n17352) );
  INV_X1 U12051 ( .A(n17416), .ZN(n17418) );
  INV_X1 U12052 ( .A(n17417), .ZN(n17415) );
  AND2_X1 U12053 ( .A1(n17512), .A2(n9923), .ZN(n16398) );
  AND2_X1 U12054 ( .A1(n9602), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9923) );
  NAND2_X1 U12055 ( .A1(n17512), .A2(n9602), .ZN(n12841) );
  NAND2_X1 U12056 ( .A1(n16408), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9713) );
  NOR2_X1 U12057 ( .A1(n17543), .A2(n17514), .ZN(n17512) );
  INV_X1 U12058 ( .A(n16772), .ZN(n17718) );
  INV_X1 U12059 ( .A(n18046), .ZN(n17712) );
  NOR2_X1 U12060 ( .A1(n17772), .A2(n17777), .ZN(n17746) );
  NOR2_X1 U12061 ( .A1(n17832), .A2(n12714), .ZN(n9720) );
  XOR2_X1 U12062 ( .A(n12813), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n17834) );
  OAI21_X1 U12063 ( .B1(n16377), .B2(n17627), .A(n16380), .ZN(n12801) );
  NAND2_X1 U12064 ( .A1(n12801), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16379) );
  NAND2_X1 U12065 ( .A1(n17488), .A2(n17627), .ZN(n15874) );
  INV_X1 U12066 ( .A(n17858), .ZN(n17475) );
  INV_X1 U12067 ( .A(n15874), .ZN(n16429) );
  NOR2_X1 U12068 ( .A1(n17499), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17498) );
  INV_X1 U12069 ( .A(n16430), .ZN(n17860) );
  NOR2_X1 U12070 ( .A1(n17893), .A2(n17535), .ZN(n17519) );
  NAND2_X1 U12071 ( .A1(n12837), .A2(n17993), .ZN(n17894) );
  NOR2_X1 U12072 ( .A1(n17627), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17606) );
  NOR2_X1 U12073 ( .A1(n17663), .A2(n17650), .ZN(n17913) );
  INV_X1 U12074 ( .A(n17686), .ZN(n18025) );
  AND2_X1 U12075 ( .A1(n12785), .A2(n9698), .ZN(n17689) );
  OAI21_X2 U12076 ( .B1(n18644), .B2(n13254), .A(n18643), .ZN(n18633) );
  NAND2_X1 U12077 ( .A1(n18842), .A2(n18120), .ZN(n18626) );
  INV_X1 U12078 ( .A(n17711), .ZN(n18044) );
  NOR2_X1 U12079 ( .A1(n17702), .A2(n20851), .ZN(n18046) );
  NOR2_X1 U12080 ( .A1(n17752), .A2(n20851), .ZN(n17751) );
  AOI21_X1 U12081 ( .B1(n10063), .B2(n9642), .A(n10062), .ZN(n10061) );
  NOR2_X1 U12082 ( .A1(n10067), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10062) );
  NOR2_X1 U12083 ( .A1(n18081), .A2(n15872), .ZN(n18623) );
  INV_X1 U12084 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18637) );
  INV_X1 U12085 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18638) );
  NAND2_X1 U12086 ( .A1(n18854), .A2(n15848), .ZN(n18648) );
  INV_X1 U12087 ( .A(n12564), .ZN(n9791) );
  NOR2_X1 U12088 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18184), .ZN(n18535) );
  INV_X1 U12089 ( .A(n18535), .ZN(n18376) );
  AOI22_X1 U12090 ( .A1(n18627), .A2(n17918), .B1(n18120), .B2(n15870), .ZN(
        n18630) );
  INV_X1 U12091 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n15851) );
  AND2_X1 U12092 ( .A1(n18786), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18725) );
  AND2_X1 U12093 ( .A1(n19888), .A2(n14503), .ZN(n15968) );
  INV_X1 U12094 ( .A(n9585), .ZN(n19944) );
  INV_X1 U12095 ( .A(n19903), .ZN(n19899) );
  NAND2_X1 U12096 ( .A1(n14095), .A2(n15925), .ZN(n19942) );
  INV_X1 U12097 ( .A(n14106), .ZN(n14095) );
  OR3_X1 U12098 ( .A1(n19972), .A2(n14100), .A3(n16149), .ZN(n19983) );
  NOR2_X2 U12099 ( .A1(n14106), .A2(n14105), .ZN(n19971) );
  AND2_X1 U12100 ( .A1(n14113), .A2(n19903), .ZN(n19976) );
  INV_X1 U12101 ( .A(n14836), .ZN(n14857) );
  NAND2_X1 U12102 ( .A1(n12518), .A2(n13280), .ZN(n14861) );
  OR2_X1 U12103 ( .A1(n13447), .A2(n12517), .ZN(n12518) );
  INV_X2 U12104 ( .A(n14861), .ZN(n14867) );
  XNOR2_X1 U12105 ( .A(n12537), .B(n12536), .ZN(n14540) );
  INV_X1 U12106 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14956) );
  INV_X1 U12107 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14972) );
  NAND2_X1 U12108 ( .A1(n13463), .A2(n15920), .ZN(n19869) );
  NAND2_X1 U12109 ( .A1(n20718), .A2(n13460), .ZN(n20055) );
  OAI211_X1 U12110 ( .C1(n11775), .C2(n15131), .A(n10129), .B(n11781), .ZN(
        n14494) );
  AND2_X1 U12111 ( .A1(n15009), .A2(n11997), .ZN(n9743) );
  NAND2_X1 U12112 ( .A1(n11998), .A2(n9742), .ZN(n9741) );
  INV_X1 U12113 ( .A(n14490), .ZN(n9742) );
  NAND2_X1 U12114 ( .A1(n14514), .A2(n16119), .ZN(n11998) );
  OR2_X1 U12115 ( .A1(n14576), .A2(n14575), .ZN(n15036) );
  OR2_X1 U12116 ( .A1(n14591), .A2(n14590), .ZN(n15041) );
  NOR3_X1 U12117 ( .A1(n15940), .A2(n9738), .A3(n9736), .ZN(n15056) );
  NAND2_X1 U12118 ( .A1(n11992), .A2(n11991), .ZN(n9736) );
  NOR3_X1 U12119 ( .A1(n15940), .A2(n9738), .A3(n9737), .ZN(n15065) );
  NOR2_X1 U12120 ( .A1(n15096), .A2(n15113), .ZN(n15111) );
  NAND2_X1 U12121 ( .A1(n11750), .A2(n11749), .ZN(n14211) );
  CLKBUF_X1 U12122 ( .A(n14146), .Z(n14149) );
  CLKBUF_X1 U12123 ( .A(n13792), .Z(n13794) );
  XNOR2_X1 U12124 ( .A(n9861), .B(n13403), .ZN(n13536) );
  INV_X1 U12125 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20386) );
  OR2_X1 U12126 ( .A1(n13673), .A2(n20216), .ZN(n20725) );
  NOR2_X1 U12127 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14558) );
  CLKBUF_X1 U12128 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n20708) );
  CLKBUF_X1 U12129 ( .A(n12511), .Z(n12512) );
  OAI211_X1 U12130 ( .C1(n20073), .C2(n20070), .A(n20391), .B(n20068), .ZN(
        n20109) );
  INV_X1 U12131 ( .A(n20230), .ZN(n20235) );
  NAND2_X1 U12132 ( .A1(n20714), .A2(n20533), .ZN(n20319) );
  OAI211_X1 U12133 ( .C1(n20353), .C2(n20338), .A(n20391), .B(n20337), .ZN(
        n20356) );
  OAI211_X1 U12134 ( .C1(n20460), .C2(n12409), .A(n20543), .B(n20459), .ZN(
        n20495) );
  OAI211_X1 U12135 ( .C1(n20566), .C2(n20544), .A(n20543), .B(n20542), .ZN(
        n20568) );
  INV_X1 U12136 ( .A(n20455), .ZN(n20578) );
  INV_X1 U12137 ( .A(n20467), .ZN(n20588) );
  INV_X1 U12138 ( .A(n20471), .ZN(n20594) );
  INV_X1 U12139 ( .A(n20475), .ZN(n20599) );
  INV_X1 U12140 ( .A(n20479), .ZN(n20605) );
  INV_X1 U12141 ( .A(n20483), .ZN(n20611) );
  INV_X1 U12142 ( .A(n20487), .ZN(n20617) );
  NOR2_X1 U12143 ( .A1(n20499), .A2(n20579), .ZN(n20625) );
  NAND2_X1 U12144 ( .A1(n20534), .A2(n20533), .ZN(n20632) );
  INV_X1 U12145 ( .A(n20621), .ZN(n20628) );
  INV_X1 U12146 ( .A(n20492), .ZN(n20626) );
  INV_X1 U12147 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16149) );
  NAND2_X1 U12148 ( .A1(n16149), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20634) );
  NAND2_X1 U12149 ( .A1(n16350), .A2(n13220), .ZN(n19841) );
  INV_X1 U12150 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19791) );
  INV_X1 U12151 ( .A(n10254), .ZN(n10255) );
  INV_X1 U12152 ( .A(n10253), .ZN(n10256) );
  OR2_X1 U12153 ( .A1(n15203), .A2(n10891), .ZN(n15224) );
  AND2_X1 U12154 ( .A1(n9954), .A2(n9953), .ZN(n15261) );
  OR3_X1 U12155 ( .A1(n19841), .A2(n19844), .A3(n16360), .ZN(n18989) );
  INV_X1 U12156 ( .A(n18974), .ZN(n19000) );
  INV_X1 U12157 ( .A(n18978), .ZN(n18999) );
  XNOR2_X1 U12158 ( .A(n13180), .B(n10944), .ZN(n15276) );
  OR2_X1 U12159 ( .A1(n11045), .A2(n11288), .ZN(n15440) );
  CLKBUF_X1 U12160 ( .A(n13953), .Z(n13954) );
  OR2_X1 U12161 ( .A1(n11206), .A2(n11205), .ZN(n13836) );
  OR2_X1 U12162 ( .A1(n11173), .A2(n11172), .ZN(n13609) );
  OR2_X1 U12163 ( .A1(n11160), .A2(n11159), .ZN(n13732) );
  OR2_X1 U12164 ( .A1(n11143), .A2(n11142), .ZN(n13565) );
  OR2_X1 U12165 ( .A1(n11127), .A2(n11126), .ZN(n13721) );
  OR2_X1 U12166 ( .A1(n11110), .A2(n11109), .ZN(n13722) );
  CLKBUF_X1 U12167 ( .A(n10337), .Z(n19139) );
  CLKBUF_X1 U12168 ( .A(n13618), .Z(n15347) );
  NAND2_X1 U12169 ( .A1(n13301), .A2(n13300), .ZN(n18986) );
  INV_X1 U12170 ( .A(n15342), .ZN(n15350) );
  INV_X1 U12171 ( .A(n14242), .ZN(n15715) );
  INV_X1 U12172 ( .A(n15410), .ZN(n19009) );
  AND2_X1 U12173 ( .A1(n13823), .A2(n10022), .ZN(n13996) );
  NOR2_X1 U12174 ( .A1(n13149), .A2(n19056), .ZN(n19048) );
  OR2_X1 U12175 ( .A1(n13378), .A2(n19009), .ZN(n19033) );
  INV_X1 U12176 ( .A(n15385), .ZN(n19056) );
  INV_X1 U12177 ( .A(n19033), .ZN(n19064) );
  NAND2_X1 U12178 ( .A1(n19104), .A2(n19843), .ZN(n19071) );
  INV_X2 U12179 ( .A(n19071), .ZN(n19102) );
  INV_X2 U12180 ( .A(n13532), .ZN(n19109) );
  AND2_X1 U12181 ( .A1(n13276), .A2(n9600), .ZN(n19107) );
  AOI21_X1 U12182 ( .B1(n15432), .B2(n12850), .A(n13217), .ZN(n15435) );
  INV_X1 U12183 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15542) );
  INV_X1 U12184 ( .A(n19121), .ZN(n16258) );
  NAND2_X1 U12185 ( .A1(n18865), .A2(n10775), .ZN(n16265) );
  INV_X1 U12186 ( .A(n19117), .ZN(n16247) );
  OR2_X1 U12187 ( .A1(n15618), .A2(n15619), .ZN(n15610) );
  NAND2_X1 U12188 ( .A1(n15490), .A2(n10878), .ZN(n15478) );
  NAND2_X1 U12189 ( .A1(n10078), .A2(n10077), .ZN(n15495) );
  AOI21_X1 U12190 ( .B1(n10084), .B2(n10082), .A(n10081), .ZN(n10077) );
  OR2_X1 U12191 ( .A1(n15677), .A2(n11042), .ZN(n15654) );
  NAND2_X1 U12192 ( .A1(n9807), .A2(n9808), .ZN(n15505) );
  OR2_X1 U12193 ( .A1(n15539), .A2(n9811), .ZN(n9807) );
  NAND2_X1 U12194 ( .A1(n9813), .A2(n9815), .ZN(n15515) );
  NAND2_X1 U12195 ( .A1(n9814), .A2(n10856), .ZN(n15530) );
  OR2_X1 U12196 ( .A1(n15539), .A2(n15540), .ZN(n9814) );
  NAND2_X1 U12197 ( .A1(n9817), .A2(n9821), .ZN(n15550) );
  NAND2_X1 U12198 ( .A1(n9825), .A2(n9822), .ZN(n9817) );
  NAND2_X1 U12199 ( .A1(n15783), .A2(n11265), .ZN(n16267) );
  AOI21_X1 U12200 ( .B1(n16182), .B2(n16180), .A(n10651), .ZN(n15730) );
  NAND2_X1 U12201 ( .A1(n10641), .A2(n10640), .ZN(n15745) );
  NOR2_X1 U12202 ( .A1(n11037), .A2(n11261), .ZN(n16310) );
  NAND2_X1 U12203 ( .A1(n14312), .A2(n10763), .ZN(n14345) );
  NAND2_X1 U12204 ( .A1(n11259), .A2(n19127), .ZN(n9834) );
  NAND2_X2 U12205 ( .A1(n10333), .A2(n10345), .ZN(n13963) );
  INV_X1 U12206 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19822) );
  INV_X1 U12207 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19803) );
  INV_X1 U12208 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16330) );
  XNOR2_X1 U12209 ( .A(n13383), .B(n13385), .ZN(n19816) );
  NAND2_X1 U12210 ( .A1(n16340), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16359) );
  CLKBUF_X1 U12211 ( .A(n10965), .Z(n10966) );
  NOR2_X1 U12212 ( .A1(n19420), .A2(n19367), .ZN(n19229) );
  NOR2_X1 U12213 ( .A1(n19367), .A2(n19481), .ZN(n19286) );
  AND2_X1 U12214 ( .A1(n19299), .A2(n19298), .ZN(n19309) );
  INV_X1 U12215 ( .A(n19337), .ZN(n19355) );
  NOR2_X2 U12216 ( .A1(n19545), .A2(n19583), .ZN(n19601) );
  INV_X1 U12217 ( .A(n19702), .ZN(n19600) );
  INV_X1 U12218 ( .A(n19601), .ZN(n19609) );
  INV_X1 U12219 ( .A(n19684), .ZN(n19632) );
  INV_X1 U12220 ( .A(n19690), .ZN(n19636) );
  NOR2_X2 U12221 ( .A1(n19584), .A2(n19583), .ZN(n19649) );
  OAI22_X1 U12222 ( .A1(n19165), .A2(n19164), .B1(n19163), .B2(n19162), .ZN(
        n19650) );
  INV_X1 U12223 ( .A(n19625), .ZN(n19665) );
  INV_X1 U12224 ( .A(n19489), .ZN(n19657) );
  INV_X1 U12225 ( .A(n19629), .ZN(n19670) );
  INV_X1 U12226 ( .A(n19499), .ZN(n19669) );
  OAI22_X1 U12227 ( .A1(n20843), .A2(n19164), .B1(n18212), .B2(n19162), .ZN(
        n19693) );
  OAI22_X1 U12228 ( .A1(n16459), .A2(n19164), .B1(n20902), .B2(n19162), .ZN(
        n19699) );
  INV_X1 U12229 ( .A(n19526), .ZN(n19697) );
  NOR2_X2 U12230 ( .A1(n19584), .A2(n19796), .ZN(n19708) );
  INV_X1 U12231 ( .A(n19655), .ZN(n19707) );
  INV_X1 U12232 ( .A(n19650), .ZN(n19713) );
  NAND2_X1 U12233 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19714), .ZN(n18863) );
  NOR2_X1 U12234 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n13325), .ZN(n19714) );
  AND2_X1 U12235 ( .A1(n16371), .A2(n16370), .ZN(n19719) );
  NOR2_X1 U12236 ( .A1(n12670), .A2(n12669), .ZN(n18854) );
  NAND2_X1 U12237 ( .A1(n18621), .A2(n17415), .ZN(n18855) );
  INV_X1 U12238 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18688) );
  INV_X1 U12239 ( .A(n16537), .ZN(n16531) );
  NAND2_X1 U12240 ( .A1(n18679), .A2(n15865), .ZN(n17417) );
  NOR2_X1 U12241 ( .A1(n18630), .A2(n18839), .ZN(n16538) );
  INV_X1 U12242 ( .A(n9915), .ZN(n16601) );
  NOR2_X1 U12243 ( .A1(n16909), .A2(n16568), .ZN(n16614) );
  NOR2_X1 U12244 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16659), .ZN(n16631) );
  INV_X1 U12245 ( .A(n9918), .ZN(n9917) );
  OAI22_X1 U12246 ( .A1(n9919), .A2(n16566), .B1(n9919), .B2(n9921), .ZN(n9918) );
  INV_X1 U12247 ( .A(n9922), .ZN(n16646) );
  NAND2_X1 U12248 ( .A1(n9920), .A2(n16876), .ZN(n9922) );
  AND3_X1 U12249 ( .A1(n9903), .A2(n9904), .A3(n16876), .ZN(n13252) );
  NAND2_X1 U12250 ( .A1(n9903), .A2(n9904), .ZN(n16664) );
  NOR2_X1 U12251 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16823), .ZN(n16805) );
  NOR4_X1 U12252 ( .A1(n16643), .A2(n14485), .A3(n16979), .A4(n14484), .ZN(
        n16927) );
  AOI21_X1 U12253 ( .B1(n16956), .B2(n9633), .A(n17198), .ZN(n16932) );
  AND2_X1 U12254 ( .A1(n16956), .A2(P3_EBX_REG_24__SCAN_IN), .ZN(n16948) );
  NOR3_X1 U12255 ( .A1(n16950), .A2(n16949), .A3(n16968), .ZN(n16956) );
  INV_X1 U12256 ( .A(n15820), .ZN(n16995) );
  NAND2_X1 U12257 ( .A1(n17019), .A2(P3_EBX_REG_19__SCAN_IN), .ZN(n17007) );
  NOR3_X1 U12258 ( .A1(n17036), .A2(n17020), .A3(n9787), .ZN(n17019) );
  NAND2_X1 U12259 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_17__SCAN_IN), 
        .ZN(n9787) );
  NOR2_X1 U12260 ( .A1(n15835), .A2(n16761), .ZN(n17080) );
  NAND2_X1 U12261 ( .A1(n17141), .A2(P3_EBX_REG_10__SCAN_IN), .ZN(n17120) );
  NOR2_X1 U12262 ( .A1(n17123), .A2(n17163), .ZN(n17141) );
  NAND2_X1 U12263 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17170), .ZN(n17163) );
  INV_X1 U12264 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n20813) );
  NOR2_X1 U12265 ( .A1(n17167), .A2(n17166), .ZN(n17170) );
  NOR2_X1 U12266 ( .A1(n17171), .A2(n17172), .ZN(n17176) );
  INV_X1 U12267 ( .A(n17171), .ZN(n17201) );
  INV_X1 U12268 ( .A(n17238), .ZN(n17234) );
  NAND2_X1 U12269 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17234), .ZN(n17233) );
  NOR3_X1 U12270 ( .A1(n17283), .A2(n17248), .A3(n17206), .ZN(n17244) );
  INV_X1 U12271 ( .A(n17286), .ZN(n17274) );
  NAND2_X1 U12272 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17287), .ZN(n17283) );
  INV_X1 U12273 ( .A(n17256), .ZN(n17282) );
  NOR3_X1 U12274 ( .A1(n17399), .A2(n17401), .A3(n17324), .ZN(n17323) );
  INV_X1 U12275 ( .A(n15879), .ZN(n17321) );
  NAND2_X1 U12276 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17333), .ZN(n17324) );
  AND2_X1 U12277 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17337), .ZN(n17333) );
  NOR2_X1 U12278 ( .A1(n17407), .A2(n17334), .ZN(n17337) );
  NOR3_X1 U12279 ( .A1(n17440), .A2(n17414), .A3(n17292), .ZN(n17338) );
  NOR2_X1 U12280 ( .A1(n17440), .A2(n17346), .ZN(n17344) );
  AOI211_X1 U12282 ( .C1(n17152), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n12710), .B(n12709), .ZN(n12711) );
  OR3_X1 U12283 ( .A1(n15961), .A2(n18185), .A3(n18193), .ZN(n15962) );
  INV_X1 U12284 ( .A(n17350), .ZN(n17317) );
  NOR2_X1 U12285 ( .A1(n18632), .A2(n20931), .ZN(n17348) );
  NAND2_X1 U12286 ( .A1(n18835), .A2(n17413), .ZN(n17354) );
  OAI211_X1 U12287 ( .C1(n18843), .C2(n18842), .A(n17416), .B(n17415), .ZN(
        n17460) );
  INV_X1 U12288 ( .A(n17430), .ZN(n17462) );
  INV_X1 U12290 ( .A(n17462), .ZN(n17464) );
  NAND2_X1 U12291 ( .A1(n17512), .A2(n9681), .ZN(n17492) );
  NAND2_X1 U12292 ( .A1(n17587), .A2(n9669), .ZN(n17575) );
  NAND2_X1 U12293 ( .A1(n17634), .A2(n9670), .ZN(n17613) );
  INV_X1 U12294 ( .A(n17696), .ZN(n17649) );
  NOR2_X1 U12295 ( .A1(n17804), .A2(n17805), .ZN(n17782) );
  NOR2_X2 U12296 ( .A1(n18376), .A2(n18532), .ZN(n18568) );
  INV_X1 U12297 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17805) );
  INV_X1 U12298 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18801) );
  INV_X1 U12299 ( .A(n17833), .ZN(n17847) );
  NOR2_X1 U12300 ( .A1(n10076), .A2(n10075), .ZN(n10074) );
  INV_X1 U12301 ( .A(n16412), .ZN(n10075) );
  INV_X1 U12302 ( .A(n15955), .ZN(n10076) );
  OR2_X1 U12303 ( .A1(n15954), .A2(n15953), .ZN(n10073) );
  NAND2_X1 U12304 ( .A1(n17536), .A2(n12794), .ZN(n17530) );
  NOR2_X1 U12305 ( .A1(n12785), .A2(n10069), .ZN(n17742) );
  OAI221_X2 U12306 ( .B1(n15871), .B2(n15870), .C1(n15871), .C2(n18219), .A(
        n18679), .ZN(n18154) );
  NAND2_X1 U12307 ( .A1(n9630), .A2(n17801), .ZN(n17800) );
  INV_X1 U12308 ( .A(n18156), .ZN(n18119) );
  INV_X1 U12309 ( .A(n18648), .ZN(n18654) );
  NOR2_X1 U12310 ( .A1(n18165), .A2(n18162), .ZN(n18156) );
  INV_X1 U12311 ( .A(n18154), .ZN(n18162) );
  INV_X1 U12312 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18670) );
  INV_X1 U12313 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18665) );
  INV_X2 U12314 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18821) );
  NOR2_X1 U12315 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18794), .ZN(
        n18815) );
  AND2_X1 U12316 ( .A1(n12529), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20053)
         );
  OAI22_X1 U12318 ( .A1(n9859), .A2(n19985), .B1(n19997), .B2(n14756), .ZN(
        P1_U2841) );
  INV_X1 U12319 ( .A(n14514), .ZN(n9859) );
  OAI21_X1 U12320 ( .B1(n14877), .B2(n19992), .A(n12472), .ZN(P1_U2843) );
  AND2_X1 U12321 ( .A1(n12471), .A2(n12470), .ZN(n12472) );
  OR2_X1 U12322 ( .A1(n15019), .A2(n19985), .ZN(n12471) );
  NAND2_X1 U12323 ( .A1(n9745), .A2(n9740), .ZN(P1_U3000) );
  AOI211_X1 U12324 ( .C1(n15015), .C2(n9744), .A(n9743), .B(n9741), .ZN(n9740)
         );
  NAND2_X1 U12325 ( .A1(n14494), .A2(n16122), .ZN(n9745) );
  NOR2_X1 U12326 ( .A1(n11994), .A2(n13442), .ZN(n9744) );
  OR2_X1 U12327 ( .A1(n15179), .A2(n15165), .ZN(n15188) );
  NAND2_X1 U12328 ( .A1(n15178), .A2(n18984), .ZN(n15179) );
  AND2_X1 U12329 ( .A1(n13183), .A2(n10118), .ZN(n13184) );
  NAND2_X1 U12330 ( .A1(n13179), .A2(n13149), .ZN(n13175) );
  INV_X1 U12331 ( .A(n12856), .ZN(n12857) );
  OAI21_X1 U12332 ( .B1(n15660), .B2(n16256), .A(n10849), .ZN(n10850) );
  NAND2_X1 U12333 ( .A1(n11318), .A2(n9779), .ZN(n9778) );
  NAND2_X1 U12334 ( .A1(n9838), .A2(n9648), .ZN(n14552) );
  OR2_X1 U12335 ( .A1(n14550), .A2(n14549), .ZN(n9838) );
  OAI211_X1 U12336 ( .C1(n15582), .C2(n11276), .A(n15586), .B(n15585), .ZN(
        n15587) );
  OR2_X1 U12337 ( .A1(n16595), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9901) );
  AOI21_X1 U12338 ( .B1(n12845), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n12844), .ZN(n12846) );
  INV_X1 U12339 ( .A(n9710), .ZN(n16409) );
  OAI21_X1 U12340 ( .B1(n16404), .B2(n17756), .A(n9711), .ZN(n9710) );
  OAI21_X1 U12341 ( .B1(n15952), .B2(n18091), .A(n10070), .ZN(P3_U2832) );
  INV_X1 U12342 ( .A(n10071), .ZN(n10070) );
  OAI211_X1 U12343 ( .C1(n20799), .C2(n10074), .A(n10073), .B(n10072), .ZN(
        n10071) );
  NAND2_X1 U12344 ( .A1(n18165), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n10072) );
  NOR2_X2 U12345 ( .A1(n12566), .A2(n16905), .ZN(n12689) );
  AND3_X1 U12346 ( .A1(n11857), .A2(n13463), .A3(n9842), .ZN(n9601) );
  NAND2_X1 U12347 ( .A1(n10005), .A2(n10006), .ZN(n14694) );
  AND2_X1 U12348 ( .A1(n9624), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9602) );
  AND2_X1 U12349 ( .A1(n9632), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n9603) );
  OR2_X1 U12351 ( .A1(n18650), .A2(n12564), .ZN(n9604) );
  NOR2_X1 U12352 ( .A1(n11994), .A2(n9645), .ZN(n9605) );
  NOR2_X1 U12353 ( .A1(n15481), .A2(n10105), .ZN(n15448) );
  NOR2_X1 U12354 ( .A1(n15481), .A2(n10876), .ZN(n15471) );
  AND2_X1 U12355 ( .A1(n10005), .A2(n10003), .ZN(n9606) );
  AND2_X1 U12356 ( .A1(n10128), .A2(n10034), .ZN(n9607) );
  OR2_X1 U12357 ( .A1(n14587), .A2(n10011), .ZN(n9608) );
  AND2_X1 U12358 ( .A1(n12860), .A2(n10358), .ZN(n9609) );
  AND2_X1 U12359 ( .A1(n12860), .A2(n10331), .ZN(n9610) );
  INV_X1 U12360 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13984) );
  AND2_X1 U12361 ( .A1(n9935), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9611) );
  AND2_X1 U12362 ( .A1(n9597), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n9612)
         );
  AND2_X1 U12363 ( .A1(n9808), .A2(n15502), .ZN(n9613) );
  AND2_X1 U12364 ( .A1(n10051), .A2(n10049), .ZN(n9614) );
  NOR2_X1 U12365 ( .A1(n15304), .A2(n15306), .ZN(n15305) );
  INV_X1 U12366 ( .A(n10087), .ZN(n10082) );
  NOR2_X1 U12367 ( .A1(n15743), .A2(n10088), .ZN(n10087) );
  AND2_X1 U12368 ( .A1(n9652), .A2(n11749), .ZN(n9615) );
  NAND4_X1 U12369 ( .A1(n11434), .A2(n11433), .A3(n11432), .A4(n11431), .ZN(
        n9616) );
  NAND2_X1 U12370 ( .A1(n12881), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n9617) );
  NAND2_X1 U12371 ( .A1(n9952), .A2(n15189), .ZN(n9618) );
  AND2_X1 U12372 ( .A1(n9979), .A2(n13089), .ZN(n9619) );
  AND3_X1 U12373 ( .A1(n12720), .A2(n12721), .A3(n10057), .ZN(n9620) );
  AND2_X1 U12374 ( .A1(n10612), .A2(n9667), .ZN(n9621) );
  NAND2_X1 U12375 ( .A1(n9931), .A2(n9932), .ZN(n13197) );
  NOR2_X1 U12376 ( .A1(n13193), .A2(n9943), .ZN(n13208) );
  NAND2_X1 U12377 ( .A1(n13190), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10777) );
  NOR2_X1 U12378 ( .A1(n13193), .A2(n14244), .ZN(n13194) );
  AND4_X1 U12379 ( .A1(n9940), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9623) );
  NAND2_X1 U12380 ( .A1(n9991), .A2(n9617), .ZN(n13561) );
  AND2_X1 U12381 ( .A1(n9681), .A2(n9924), .ZN(n9624) );
  AND2_X1 U12382 ( .A1(n9982), .A2(n14170), .ZN(n9625) );
  NAND2_X1 U12383 ( .A1(n12903), .A2(n9982), .ZN(n9626) );
  OR3_X1 U12384 ( .A1(n14672), .A2(n9675), .A3(n9879), .ZN(n9627) );
  AND2_X1 U12385 ( .A1(n9871), .A2(n9663), .ZN(n9628) );
  AND2_X1 U12386 ( .A1(n9625), .A2(n15346), .ZN(n9629) );
  NAND2_X1 U12387 ( .A1(n12849), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12850) );
  NOR2_X1 U12388 ( .A1(n17811), .A2(n12739), .ZN(n9630) );
  NAND2_X1 U12389 ( .A1(n13190), .A2(n9611), .ZN(n13188) );
  INV_X1 U12390 ( .A(n17474), .ZN(n9914) );
  AND2_X1 U12391 ( .A1(n9781), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n9631) );
  AND2_X1 U12392 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .ZN(n9632) );
  AND2_X1 U12393 ( .A1(n9603), .A2(n15821), .ZN(n9633) );
  AND2_X1 U12394 ( .A1(n9590), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10427) );
  OR2_X1 U12395 ( .A1(n10880), .A2(n10879), .ZN(n9634) );
  NAND2_X1 U12396 ( .A1(n10770), .A2(n10769), .ZN(n15506) );
  OR2_X1 U12397 ( .A1(n12564), .A2(n12563), .ZN(n9635) );
  AND2_X1 U12398 ( .A1(n16956), .A2(n9603), .ZN(n9636) );
  INV_X2 U12399 ( .A(n11753), .ZN(n15941) );
  NOR2_X1 U12400 ( .A1(n14587), .A2(n14588), .ZN(n14572) );
  AND2_X1 U12401 ( .A1(n10338), .A2(n10350), .ZN(n10388) );
  AND2_X1 U12402 ( .A1(n16956), .A2(n9632), .ZN(n9637) );
  AND2_X1 U12403 ( .A1(n11440), .A2(n11441), .ZN(n9638) );
  NOR2_X1 U12404 ( .A1(n15552), .A2(n10100), .ZN(n10773) );
  INV_X1 U12405 ( .A(n11350), .ZN(n12273) );
  NAND2_X1 U12406 ( .A1(n15247), .A2(n15382), .ZN(n15234) );
  OR2_X1 U12407 ( .A1(n15481), .A2(n10106), .ZN(n15463) );
  AND2_X1 U12408 ( .A1(n11595), .A2(n11594), .ZN(n9639) );
  OR2_X1 U12409 ( .A1(n12779), .A2(n12778), .ZN(n9640) );
  AND2_X1 U12410 ( .A1(n14600), .A2(n10008), .ZN(n12537) );
  AND4_X1 U12411 ( .A1(n12616), .A2(n12615), .A3(n12614), .A4(n12613), .ZN(
        n9641) );
  NOR2_X1 U12412 ( .A1(n14723), .A2(n14777), .ZN(n14708) );
  AND2_X1 U12413 ( .A1(n15747), .A2(n10113), .ZN(n15726) );
  NAND2_X1 U12414 ( .A1(n15747), .A2(n15731), .ZN(n15748) );
  OR2_X1 U12415 ( .A1(n17801), .A2(n10066), .ZN(n9642) );
  NAND2_X1 U12416 ( .A1(n11344), .A2(n10144), .ZN(n11381) );
  AND2_X1 U12417 ( .A1(n10330), .A2(n10350), .ZN(n10469) );
  INV_X1 U12418 ( .A(n13091), .ZN(n9975) );
  NAND2_X1 U12419 ( .A1(n10094), .A2(n10626), .ZN(n15784) );
  NAND2_X1 U12420 ( .A1(n11381), .A2(n12000), .ZN(n11472) );
  NOR2_X1 U12421 ( .A1(n15481), .A2(n9772), .ZN(n11011) );
  NOR2_X1 U12422 ( .A1(n10274), .A2(n13121), .ZN(n10276) );
  AND2_X1 U12423 ( .A1(n12870), .A2(n13963), .ZN(n9643) );
  NOR2_X1 U12424 ( .A1(n15305), .A2(n13036), .ZN(n13055) );
  OR2_X1 U12425 ( .A1(n15447), .A2(n19137), .ZN(n9644) );
  OR2_X1 U12426 ( .A1(n15481), .A2(n10103), .ZN(n11281) );
  AND2_X1 U12427 ( .A1(n15056), .A2(n11995), .ZN(n9645) );
  NOR2_X1 U12428 ( .A1(n14634), .A2(n14635), .ZN(n14624) );
  OR3_X1 U12429 ( .A1(n9634), .A2(P2_EBX_REG_25__SCAN_IN), .A3(
        P2_EBX_REG_24__SCAN_IN), .ZN(n9646) );
  INV_X1 U12430 ( .A(n9980), .ZN(n15294) );
  NAND2_X1 U12431 ( .A1(n9994), .A2(n12110), .ZN(n12019) );
  NAND2_X1 U12432 ( .A1(n16231), .A2(n10768), .ZN(n15746) );
  INV_X1 U12433 ( .A(n10956), .ZN(n9883) );
  AND2_X1 U12434 ( .A1(n10758), .A2(n14192), .ZN(n9647) );
  AND2_X1 U12435 ( .A1(n10120), .A2(n9837), .ZN(n9648) );
  AND2_X1 U12436 ( .A1(n16098), .A2(n16092), .ZN(n16071) );
  OR2_X1 U12437 ( .A1(n12855), .A2(n19137), .ZN(n9649) );
  NAND2_X1 U12438 ( .A1(n15746), .A2(n9776), .ZN(n10853) );
  NAND4_X1 U12439 ( .A1(n11439), .A2(n11438), .A3(n11437), .A4(n11436), .ZN(
        n9650) );
  NOR2_X1 U12440 ( .A1(n13379), .A2(n9607), .ZN(n11064) );
  OR2_X1 U12441 ( .A1(n15196), .A2(n9951), .ZN(n9952) );
  AND2_X1 U12442 ( .A1(n15233), .A2(n15213), .ZN(n11286) );
  NAND2_X2 U12443 ( .A1(n11418), .A2(n10146), .ZN(n9858) );
  AND3_X1 U12444 ( .A1(n9957), .A2(n9958), .A3(n9960), .ZN(n9651) );
  OR2_X1 U12445 ( .A1(n15131), .A2(n11751), .ZN(n9652) );
  NOR2_X1 U12446 ( .A1(n11534), .A2(n20744), .ZN(n11742) );
  NAND2_X1 U12447 ( .A1(n9998), .A2(n14734), .ZN(n14736) );
  NAND2_X1 U12448 ( .A1(n10285), .A2(n10279), .ZN(n10323) );
  AND2_X1 U12449 ( .A1(n10244), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9653) );
  AND2_X1 U12450 ( .A1(n12725), .A2(n12724), .ZN(n9654) );
  OR2_X1 U12451 ( .A1(n10633), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n9655) );
  INV_X1 U12452 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10192) );
  INV_X2 U12453 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20744) );
  INV_X1 U12454 ( .A(n10251), .ZN(n11021) );
  AND2_X1 U12455 ( .A1(n9915), .A2(n9914), .ZN(n9656) );
  INV_X1 U12456 ( .A(n10309), .ZN(n9803) );
  AND2_X1 U12457 ( .A1(n10315), .A2(n10320), .ZN(n10309) );
  NAND2_X1 U12458 ( .A1(n11096), .A2(n11095), .ZN(n14351) );
  OR2_X1 U12459 ( .A1(n14616), .A2(n9874), .ZN(n9657) );
  NOR2_X1 U12460 ( .A1(n15395), .A2(n15394), .ZN(n15248) );
  INV_X1 U12461 ( .A(n12862), .ZN(n9964) );
  INV_X1 U12462 ( .A(n11477), .ZN(n11563) );
  INV_X1 U12463 ( .A(n11477), .ZN(n9842) );
  NOR2_X1 U12464 ( .A1(n13195), .A2(n16189), .ZN(n13196) );
  NOR2_X1 U12465 ( .A1(n13200), .A2(n18973), .ZN(n13201) );
  NOR2_X1 U12466 ( .A1(n13203), .A2(n13984), .ZN(n13204) );
  NOR2_X1 U12467 ( .A1(n13198), .A2(n16227), .ZN(n13199) );
  INV_X1 U12468 ( .A(n11536), .ZN(n9759) );
  NAND2_X1 U12469 ( .A1(n17618), .A2(n17743), .ZN(n17536) );
  AND3_X1 U12470 ( .A1(n12065), .A2(n14065), .A3(n10001), .ZN(n14225) );
  AND2_X1 U12471 ( .A1(n12903), .A2(n9629), .ZN(n15339) );
  AND3_X1 U12472 ( .A1(n12065), .A2(n14065), .A3(n10000), .ZN(n14326) );
  AND2_X1 U12473 ( .A1(n14351), .A2(n10025), .ZN(n13868) );
  NAND2_X1 U12474 ( .A1(n14065), .A2(n12065), .ZN(n14164) );
  INV_X1 U12475 ( .A(n11487), .ZN(n9841) );
  NOR2_X1 U12476 ( .A1(n14039), .A2(n15733), .ZN(n14240) );
  INV_X1 U12477 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11321) );
  NAND2_X1 U12478 ( .A1(n14174), .A2(n14173), .ZN(n14172) );
  NAND2_X1 U12479 ( .A1(n15879), .A2(n12777), .ZN(n17743) );
  INV_X1 U12480 ( .A(n17743), .ZN(n17627) );
  NOR2_X1 U12481 ( .A1(n15247), .A2(n15250), .ZN(n9658) );
  OR2_X1 U12482 ( .A1(n14780), .A2(n9867), .ZN(n9659) );
  AND2_X1 U12483 ( .A1(n14173), .A2(n10042), .ZN(n9660) );
  AND2_X1 U12484 ( .A1(n10046), .A2(n13838), .ZN(n9661) );
  BUF_X1 U12485 ( .A(n12870), .Z(n13541) );
  NAND2_X1 U12486 ( .A1(n9755), .A2(n11727), .ZN(n16061) );
  AND2_X1 U12487 ( .A1(n15269), .A2(n15270), .ZN(n15268) );
  OAI21_X1 U12488 ( .B1(n15792), .B2(n12869), .A(n12865), .ZN(n13383) );
  NAND2_X1 U12489 ( .A1(n11501), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12188) );
  INV_X1 U12490 ( .A(n12188), .ZN(n12125) );
  AND2_X1 U12491 ( .A1(n14255), .A2(n11234), .ZN(n15269) );
  NAND2_X1 U12492 ( .A1(n15269), .A2(n10033), .ZN(n15401) );
  NOR2_X1 U12493 ( .A1(n15718), .A2(n14256), .ZN(n14255) );
  AND2_X1 U12494 ( .A1(n15318), .A2(n13017), .ZN(n15304) );
  AND2_X1 U12495 ( .A1(n11847), .A2(n11818), .ZN(n9662) );
  AND2_X1 U12496 ( .A1(n14739), .A2(n14740), .ZN(n9663) );
  OR2_X1 U12497 ( .A1(n15766), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9664) );
  OR2_X1 U12498 ( .A1(n13917), .A2(n16206), .ZN(n9665) );
  AND2_X1 U12499 ( .A1(n9628), .A2(n14788), .ZN(n9666) );
  AND2_X1 U12500 ( .A1(n16235), .A2(n16233), .ZN(n9667) );
  AND3_X1 U12501 ( .A1(n11165), .A2(n11164), .A3(n11163), .ZN(n9668) );
  OR2_X1 U12502 ( .A1(n10433), .A2(n10432), .ZN(n10731) );
  INV_X1 U12503 ( .A(n11991), .ZN(n9737) );
  AND2_X1 U12504 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9669) );
  AND2_X1 U12505 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n9670) );
  INV_X1 U12506 ( .A(n9846), .ZN(n16045) );
  NAND2_X1 U12507 ( .A1(n15131), .A2(n11762), .ZN(n9846) );
  INV_X1 U12508 ( .A(n9823), .ZN(n9822) );
  NAND2_X1 U12509 ( .A1(n10857), .A2(n16179), .ZN(n9823) );
  NAND2_X1 U12510 ( .A1(n9826), .A2(n15560), .ZN(n9671) );
  NOR2_X1 U12511 ( .A1(n12864), .A2(n9964), .ZN(n9672) );
  AND2_X1 U12512 ( .A1(n9922), .A2(n9921), .ZN(n9673) );
  AND2_X1 U12513 ( .A1(n9992), .A2(n13836), .ZN(n9674) );
  INV_X1 U12514 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16264) );
  OR2_X1 U12515 ( .A1(n14647), .A2(n15945), .ZN(n9675) );
  INV_X1 U12517 ( .A(n19133), .ZN(n16300) );
  NAND2_X1 U12518 ( .A1(n11258), .A2(n11014), .ZN(n19137) );
  AND2_X1 U12519 ( .A1(n13562), .A2(n9992), .ZN(n13746) );
  NAND2_X1 U12520 ( .A1(n13823), .A2(n13822), .ZN(n13824) );
  INV_X1 U12521 ( .A(n13033), .ZN(n9989) );
  AND2_X1 U12522 ( .A1(n13191), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13190) );
  NAND2_X1 U12523 ( .A1(n13562), .A2(n12888), .ZN(n13608) );
  AND2_X1 U12524 ( .A1(n12903), .A2(n9625), .ZN(n9676) );
  AND2_X1 U12525 ( .A1(n12903), .A2(n12902), .ZN(n9677) );
  OR2_X1 U12526 ( .A1(n14780), .A2(n14779), .ZN(n9678) );
  OR2_X1 U12527 ( .A1(n11191), .A2(n11190), .ZN(n9679) );
  NOR2_X1 U12528 ( .A1(n13193), .A2(n9941), .ZN(n13191) );
  AND2_X1 U12529 ( .A1(n10029), .A2(n10028), .ZN(n9680) );
  AND2_X1 U12530 ( .A1(n17511), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9681) );
  AND2_X1 U12531 ( .A1(n13190), .A2(n9934), .ZN(n13189) );
  INV_X1 U12532 ( .A(n19862), .ZN(n13280) );
  OR2_X1 U12533 ( .A1(n11987), .A2(n11869), .ZN(n16136) );
  INV_X1 U12534 ( .A(n16136), .ZN(n16119) );
  NAND2_X1 U12535 ( .A1(n10050), .A2(n9614), .ZN(n9682) );
  NOR2_X1 U12536 ( .A1(n12784), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12785) );
  INV_X1 U12537 ( .A(n12785), .ZN(n10068) );
  AND2_X1 U12538 ( .A1(n9899), .A2(n9898), .ZN(n9683) );
  AND2_X1 U12539 ( .A1(n13033), .A2(n9990), .ZN(n9684) );
  AND2_X1 U12540 ( .A1(n11054), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n9685) );
  AOI21_X1 U12541 ( .B1(n18921), .B2(n9953), .A(n9951), .ZN(n18901) );
  NOR2_X1 U12542 ( .A1(n13880), .A2(n11147), .ZN(n13844) );
  AND2_X1 U12543 ( .A1(n18225), .A2(n17201), .ZN(n17198) );
  INV_X2 U12544 ( .A(n17198), .ZN(n17192) );
  AND2_X1 U12545 ( .A1(n13561), .A2(n9674), .ZN(n9686) );
  AND2_X1 U12546 ( .A1(n17627), .A2(n15950), .ZN(n9687) );
  NAND2_X1 U12547 ( .A1(n10064), .A2(n10061), .ZN(n17783) );
  INV_X1 U12548 ( .A(n13089), .ZN(n9981) );
  AND2_X1 U12549 ( .A1(n9680), .A2(n10027), .ZN(n9688) );
  AND2_X1 U12550 ( .A1(n10054), .A2(n10053), .ZN(n9689) );
  OR2_X1 U12551 ( .A1(n15144), .A2(n11988), .ZN(n9690) );
  NOR3_X1 U12552 ( .A1(n14672), .A2(n9675), .A3(n9878), .ZN(n9881) );
  NAND2_X1 U12553 ( .A1(n17141), .A2(n9781), .ZN(n9783) );
  AND2_X1 U12554 ( .A1(n9683), .A2(n15333), .ZN(n9691) );
  NAND2_X1 U12555 ( .A1(n10637), .A2(n15788), .ZN(n9692) );
  INV_X1 U12556 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n9933) );
  INV_X1 U12557 ( .A(n15742), .ZN(n10085) );
  AND2_X1 U12558 ( .A1(n13583), .A2(n13582), .ZN(n9693) );
  AND2_X1 U12559 ( .A1(n13190), .A2(n9935), .ZN(n9694) );
  AND2_X1 U12560 ( .A1(n9927), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9695) );
  OR2_X1 U12561 ( .A1(n13193), .A2(n9944), .ZN(n9696) );
  AND2_X1 U12562 ( .A1(n9906), .A2(n16876), .ZN(n9697) );
  NAND2_X1 U12563 ( .A1(n12849), .A2(n9927), .ZN(n13216) );
  NAND2_X1 U12564 ( .A1(n10774), .A2(n10383), .ZN(n16256) );
  INV_X1 U12565 ( .A(n16256), .ZN(n19118) );
  NOR2_X1 U12566 ( .A1(n13210), .A2(n15467), .ZN(n13212) );
  INV_X1 U12567 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n9866) );
  INV_X1 U12568 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10066) );
  INV_X1 U12569 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n9937) );
  INV_X1 U12570 ( .A(n15402), .ZN(n10032) );
  INV_X1 U12571 ( .A(n11501), .ZN(n9843) );
  AND3_X1 U12572 ( .A1(n18019), .A2(n12781), .A3(n12780), .ZN(n9698) );
  INV_X1 U12573 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n9898) );
  NAND2_X1 U12574 ( .A1(n17512), .A2(n9624), .ZN(n9926) );
  INV_X1 U12575 ( .A(n11257), .ZN(n19113) );
  INV_X1 U12576 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n9928) );
  OR2_X1 U12577 ( .A1(n12916), .A2(n12915), .ZN(n9699) );
  NOR2_X2 U12578 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14128) );
  NOR2_X1 U12579 ( .A1(n15104), .A2(n15113), .ZN(n9700) );
  INV_X1 U12580 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9925) );
  INV_X1 U12581 ( .A(n13488), .ZN(n9844) );
  AND2_X1 U12582 ( .A1(n13637), .A2(n13636), .ZN(n9701) );
  INV_X1 U12583 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n9864) );
  INV_X1 U12584 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n9890) );
  INV_X1 U12585 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9840) );
  OAI221_X1 U12586 ( .B1(n20234), .B2(n20338), .C1(n20234), .C2(n20217), .A(
        n20543), .ZN(n20236) );
  INV_X1 U12587 ( .A(n20513), .ZN(n9702) );
  INV_X1 U12588 ( .A(n9702), .ZN(n9703) );
  INV_X1 U12589 ( .A(n20622), .ZN(n9704) );
  INV_X1 U12590 ( .A(n9704), .ZN(n9705) );
  INV_X1 U12591 ( .A(n20526), .ZN(n9706) );
  INV_X1 U12592 ( .A(n9706), .ZN(n9707) );
  INV_X1 U12593 ( .A(n20633), .ZN(n9708) );
  INV_X1 U12594 ( .A(n9708), .ZN(n9709) );
  AOI22_X2 U12595 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20102), .B1(DATAI_23_), 
        .B2(n20103), .ZN(n20571) );
  AOI22_X2 U12596 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20102), .B1(DATAI_18_), 
        .B2(n20103), .ZN(n20597) );
  AOI22_X2 U12597 ( .A1(DATAI_21_), .A2(n20103), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20102), .ZN(n20615) );
  NOR2_X2 U12598 ( .A1(n20055), .A2(n20054), .ZN(n20102) );
  NOR2_X2 U12599 ( .A1(n18194), .A2(n18285), .ZN(n18575) );
  INV_X1 U12600 ( .A(n18568), .ZN(n18285) );
  AOI22_X2 U12601 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20102), .B1(DATAI_27_), 
        .B2(n20103), .ZN(n20517) );
  NOR2_X2 U12602 ( .A1(n20053), .A2(n20055), .ZN(n20103) );
  INV_X1 U12603 ( .A(n12790), .ZN(n9717) );
  NOR2_X1 U12604 ( .A1(n17775), .A2(n17774), .ZN(n17773) );
  NOR2_X1 U12605 ( .A1(n17823), .A2(n9719), .ZN(n18141) );
  AND2_X1 U12606 ( .A1(n17824), .A2(n9720), .ZN(n9719) );
  NOR2_X1 U12607 ( .A1(n9720), .A2(n17824), .ZN(n17823) );
  NAND3_X1 U12608 ( .A1(n12794), .A2(n17535), .A3(n17536), .ZN(n17521) );
  NOR2_X1 U12609 ( .A1(n9724), .A2(n9723), .ZN(n9722) );
  NAND3_X1 U12610 ( .A1(n9753), .A2(n9638), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11638) );
  NOR2_X2 U12611 ( .A1(n9754), .A2(n11480), .ZN(n11784) );
  NAND2_X1 U12612 ( .A1(n16061), .A2(n16063), .ZN(n11740) );
  NAND2_X1 U12613 ( .A1(n14141), .A2(n14140), .ZN(n9755) );
  NAND2_X2 U12614 ( .A1(n11543), .A2(n9757), .ZN(n11584) );
  AOI21_X2 U12615 ( .B1(n11491), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11490), 
        .ZN(n9757) );
  NAND2_X1 U12616 ( .A1(n13768), .A2(n13767), .ZN(n11683) );
  NAND2_X1 U12617 ( .A1(n13702), .A2(n13703), .ZN(n9758) );
  NAND2_X1 U12618 ( .A1(n11630), .A2(n11629), .ZN(n13702) );
  OAI21_X2 U12619 ( .B1(n15942), .B2(n11937), .A(n15131), .ZN(n14943) );
  NAND2_X1 U12620 ( .A1(n11381), .A2(n9759), .ZN(n11465) );
  NAND2_X2 U12621 ( .A1(n15153), .A2(n11752), .ZN(n15001) );
  NAND2_X2 U12622 ( .A1(n11750), .A2(n9615), .ZN(n15153) );
  XNOR2_X2 U12623 ( .A(n11573), .B(n11572), .ZN(n12013) );
  NAND2_X2 U12624 ( .A1(n10385), .A2(n10384), .ZN(n9760) );
  NAND2_X1 U12625 ( .A1(n14312), .A2(n9761), .ZN(n9762) );
  NAND2_X1 U12626 ( .A1(n9622), .A2(n9762), .ZN(n16228) );
  INV_X1 U12627 ( .A(n16228), .ZN(n10765) );
  NAND2_X1 U12628 ( .A1(n10280), .A2(n9765), .ZN(n10281) );
  NAND2_X1 U12629 ( .A1(n9764), .A2(n10268), .ZN(n10282) );
  NAND2_X1 U12630 ( .A1(n15481), .A2(n10855), .ZN(n9766) );
  OAI211_X1 U12631 ( .C1(n15481), .C2(n9768), .A(n9767), .B(n9766), .ZN(n11300) );
  NOR2_X2 U12632 ( .A1(n9775), .A2(n9774), .ZN(n10770) );
  INV_X1 U12633 ( .A(n10770), .ZN(n15552) );
  INV_X1 U12634 ( .A(n10853), .ZN(n10854) );
  NAND4_X1 U12635 ( .A1(n10216), .A2(n10264), .A3(n10254), .A4(n9777), .ZN(
        n10219) );
  INV_X1 U12636 ( .A(n9783), .ZN(n17093) );
  AOI211_X1 U12637 ( .C1(n17150), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n9786), .B(n9785), .ZN(n9784) );
  NOR2_X1 U12638 ( .A1(n12578), .A2(n20813), .ZN(n9785) );
  INV_X1 U12639 ( .A(n12618), .ZN(n9786) );
  INV_X2 U12640 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12565) );
  NAND2_X2 U12642 ( .A1(n9794), .A2(n9793), .ZN(n10531) );
  NAND4_X1 U12643 ( .A1(n10152), .A2(n10150), .A3(n10151), .A4(n10149), .ZN(
        n9793) );
  NAND4_X1 U12644 ( .A1(n10157), .A2(n10155), .A3(n10156), .A4(n10154), .ZN(
        n9794) );
  INV_X1 U12645 ( .A(n13298), .ZN(n9795) );
  NAND2_X2 U12646 ( .A1(n9802), .A2(n9800), .ZN(n10337) );
  NAND3_X1 U12647 ( .A1(n10309), .A2(n10316), .A3(n10332), .ZN(n9802) );
  INV_X2 U12648 ( .A(n10337), .ZN(n12860) );
  NAND2_X1 U12649 ( .A1(n15539), .A2(n9613), .ZN(n9806) );
  NAND2_X2 U12650 ( .A1(n13121), .A2(n10274), .ZN(n13221) );
  AND2_X2 U12651 ( .A1(n9830), .A2(n9828), .ZN(n10274) );
  NAND3_X1 U12652 ( .A1(n10239), .A2(n10240), .A3(n9829), .ZN(n9828) );
  NAND4_X1 U12653 ( .A1(n10245), .A2(n10243), .A3(n10242), .A4(n9653), .ZN(
        n9830) );
  NOR2_X1 U12654 ( .A1(n19130), .A2(n9833), .ZN(n9832) );
  AND2_X2 U12655 ( .A1(n11326), .A2(n13640), .ZN(n11391) );
  AND2_X2 U12656 ( .A1(n9840), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11326) );
  NAND2_X1 U12657 ( .A1(n9841), .A2(n9759), .ZN(n12465) );
  OR2_X1 U12658 ( .A1(n11487), .A2(n9843), .ZN(n11967) );
  OR2_X1 U12659 ( .A1(n11487), .A2(n9701), .ZN(n13651) );
  NOR2_X1 U12660 ( .A1(n11487), .A2(n9844), .ZN(n13483) );
  NAND2_X1 U12661 ( .A1(n12014), .A2(n9851), .ZN(n9849) );
  NAND2_X1 U12662 ( .A1(n12014), .A2(n20744), .ZN(n9850) );
  NAND3_X1 U12663 ( .A1(n11731), .A2(n12057), .A3(n11741), .ZN(n11725) );
  NAND2_X1 U12664 ( .A1(n9853), .A2(n9854), .ZN(n11703) );
  NAND2_X1 U12665 ( .A1(n9854), .A2(n20211), .ZN(n11670) );
  OAI21_X1 U12666 ( .B1(n15001), .B2(n11766), .A(n11765), .ZN(n14949) );
  NAND3_X1 U12667 ( .A1(n9857), .A2(n9856), .A3(n14961), .ZN(n14948) );
  NAND3_X1 U12668 ( .A1(n9857), .A2(n9856), .A3(n9855), .ZN(n15942) );
  INV_X1 U12669 ( .A(n9858), .ZN(n11479) );
  NAND2_X1 U12670 ( .A1(n11563), .A2(n9858), .ZN(n11480) );
  NAND2_X1 U12671 ( .A1(n11786), .A2(n9858), .ZN(n11420) );
  NAND2_X1 U12672 ( .A1(n14092), .A2(n9858), .ZN(n11623) );
  NAND2_X1 U12673 ( .A1(n20104), .A2(n9858), .ZN(n20475) );
  INV_X1 U12674 ( .A(n9881), .ZN(n14626) );
  NAND2_X1 U12675 ( .A1(n10633), .A2(n10890), .ZN(n9887) );
  NAND2_X1 U12676 ( .A1(n9887), .A2(n9886), .ZN(n10647) );
  INV_X1 U12677 ( .A(n10633), .ZN(n9891) );
  NAND3_X1 U12678 ( .A1(n10615), .A2(n9894), .A3(n10571), .ZN(n9892) );
  NOR2_X4 U12679 ( .A1(n10545), .A2(n9892), .ZN(n10631) );
  INV_X1 U12680 ( .A(n10571), .ZN(n9895) );
  INV_X1 U12681 ( .A(n10545), .ZN(n10570) );
  NOR2_X1 U12682 ( .A1(n9634), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10885) );
  NAND3_X1 U12683 ( .A1(n16588), .A2(n16587), .A3(n9901), .ZN(P3_U2641) );
  INV_X1 U12684 ( .A(n9906), .ZN(n16672) );
  NAND2_X1 U12685 ( .A1(n9907), .A2(n9908), .ZN(n16590) );
  NAND2_X1 U12686 ( .A1(n16610), .A2(n16876), .ZN(n9907) );
  NAND2_X1 U12687 ( .A1(n9913), .A2(n16876), .ZN(n9915) );
  INV_X1 U12688 ( .A(n16609), .ZN(n9913) );
  NAND2_X1 U12689 ( .A1(n9916), .A2(n9917), .ZN(n16633) );
  NAND2_X1 U12690 ( .A1(n16653), .A2(n16876), .ZN(n9916) );
  INV_X1 U12691 ( .A(n16652), .ZN(n9920) );
  INV_X1 U12692 ( .A(n9926), .ZN(n16397) );
  NAND2_X1 U12693 ( .A1(n9931), .A2(n9929), .ZN(n13195) );
  NAND2_X1 U12694 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n9939) );
  NAND3_X1 U12695 ( .A1(n9940), .A2(n9938), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13200) );
  NOR2_X1 U12696 ( .A1(n16264), .A2(n9939), .ZN(n9938) );
  INV_X1 U12697 ( .A(n13203), .ZN(n9940) );
  NAND3_X1 U12698 ( .A1(n9940), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13202) );
  NAND2_X1 U12699 ( .A1(n15197), .A2(n9949), .ZN(n9945) );
  NOR2_X1 U12700 ( .A1(n15197), .A2(n15443), .ZN(n15196) );
  NAND2_X1 U12701 ( .A1(n9945), .A2(n9946), .ZN(n15177) );
  INV_X1 U12702 ( .A(n9954), .ZN(n15260) );
  NAND2_X1 U12703 ( .A1(n10195), .A2(n10194), .ZN(n9959) );
  NAND3_X1 U12704 ( .A1(n10141), .A2(n10135), .A3(n10177), .ZN(n9960) );
  INV_X2 U12705 ( .A(n10233), .ZN(n10252) );
  NAND2_X2 U12706 ( .A1(n9959), .A2(n9958), .ZN(n10233) );
  NAND2_X1 U12707 ( .A1(n9956), .A2(n9957), .ZN(n10217) );
  NAND4_X2 U12708 ( .A1(n9651), .A2(n9956), .A3(n10251), .A4(n9955), .ZN(
        n10253) );
  OAI21_X2 U12709 ( .B1(n12860), .B2(n9964), .A(n9962), .ZN(n12868) );
  NAND2_X1 U12710 ( .A1(n9965), .A2(n9672), .ZN(n9966) );
  NAND2_X1 U12711 ( .A1(n12868), .A2(n9966), .ZN(n13523) );
  NAND2_X1 U12712 ( .A1(n15278), .A2(n9970), .ZN(n9967) );
  NAND2_X1 U12713 ( .A1(n15278), .A2(n15277), .ZN(n15279) );
  OAI211_X1 U12714 ( .C1(n15278), .C2(n9972), .A(n9967), .B(n9968), .ZN(n13179) );
  OAI21_X1 U12715 ( .B1(n15293), .B2(n9977), .A(n9974), .ZN(n13091) );
  INV_X1 U12716 ( .A(n13071), .ZN(n9979) );
  NAND3_X1 U12717 ( .A1(n9987), .A2(n9985), .A3(n9984), .ZN(n15318) );
  NAND2_X1 U12718 ( .A1(n15323), .A2(n9989), .ZN(n9984) );
  INV_X1 U12719 ( .A(n15323), .ZN(n9983) );
  NAND3_X1 U12720 ( .A1(n9987), .A2(n9988), .A3(n9984), .ZN(n15317) );
  NOR2_X1 U12721 ( .A1(n15323), .A2(n15325), .ZN(n13016) );
  NAND2_X1 U12722 ( .A1(n9989), .A2(n15325), .ZN(n9988) );
  INV_X1 U12723 ( .A(n13577), .ZN(n9991) );
  AND2_X2 U12724 ( .A1(n9993), .A2(n11328), .ZN(n11345) );
  AND2_X2 U12725 ( .A1(n9993), .A2(n11327), .ZN(n11435) );
  AND2_X2 U12726 ( .A1(n13638), .A2(n9993), .ZN(n11406) );
  AND2_X2 U12727 ( .A1(n13640), .A2(n9993), .ZN(n11412) );
  AND2_X2 U12728 ( .A1(n11320), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9993) );
  XNOR2_X2 U12729 ( .A(n12019), .B(n12020), .ZN(n13739) );
  NAND2_X1 U12730 ( .A1(n9995), .A2(n11651), .ZN(n9994) );
  NAND2_X1 U12731 ( .A1(n11651), .A2(n11618), .ZN(n11999) );
  NAND2_X1 U12732 ( .A1(n13739), .A2(n13740), .ZN(n12023) );
  NAND2_X1 U12733 ( .A1(n9998), .A2(n9996), .ZN(n14721) );
  NAND3_X1 U12734 ( .A1(n12065), .A2(n9999), .A3(n14065), .ZN(n14333) );
  INV_X1 U12735 ( .A(n14723), .ZN(n10005) );
  NAND2_X1 U12736 ( .A1(n10005), .A2(n10002), .ZN(n14668) );
  NAND2_X1 U12737 ( .A1(n14600), .A2(n14601), .ZN(n14587) );
  NAND2_X1 U12738 ( .A1(n10015), .A2(n10013), .ZN(P2_U3015) );
  NAND2_X1 U12739 ( .A1(n11319), .A2(n16300), .ZN(n10015) );
  NAND2_X1 U12740 ( .A1(n10020), .A2(n11092), .ZN(n13892) );
  NAND2_X1 U12741 ( .A1(n13823), .A2(n10021), .ZN(n10020) );
  NAND2_X1 U12742 ( .A1(n14351), .A2(n10024), .ZN(n13880) );
  NAND2_X1 U12743 ( .A1(n15269), .A2(n10031), .ZN(n15395) );
  INV_X1 U12744 ( .A(n11055), .ZN(n10035) );
  NAND3_X1 U12745 ( .A1(n10035), .A2(n10036), .A3(n10252), .ZN(n10034) );
  OR2_X2 U12746 ( .A1(n13161), .A2(n11055), .ZN(n11307) );
  INV_X1 U12747 ( .A(n10531), .ZN(n10038) );
  NAND3_X1 U12748 ( .A1(n10251), .A2(n10037), .A3(n10214), .ZN(n10269) );
  NAND3_X1 U12749 ( .A1(n10039), .A2(n13583), .A3(n10796), .ZN(n13717) );
  NAND2_X1 U12750 ( .A1(n10045), .A2(n10043), .ZN(n13956) );
  NAND2_X1 U12751 ( .A1(n11286), .A2(n10054), .ZN(n15176) );
  NAND2_X1 U12752 ( .A1(n11286), .A2(n10056), .ZN(n11044) );
  AND2_X1 U12753 ( .A1(n11286), .A2(n11287), .ZN(n11045) );
  NAND4_X1 U12754 ( .A1(n12722), .A2(n10059), .A3(n9654), .A4(n9620), .ZN(
        n12811) );
  NAND2_X1 U12755 ( .A1(n17487), .A2(n17476), .ZN(n15873) );
  NAND2_X1 U12756 ( .A1(n17487), .A2(n10060), .ZN(n16377) );
  NAND3_X1 U12757 ( .A1(n17813), .A2(n10065), .A3(n9642), .ZN(n10064) );
  INV_X1 U12758 ( .A(n17801), .ZN(n10067) );
  INV_X1 U12759 ( .A(n10866), .ZN(n10081) );
  NAND2_X1 U12760 ( .A1(n10641), .A2(n10087), .ZN(n10086) );
  INV_X1 U12761 ( .A(n10641), .ZN(n10083) );
  OAI211_X1 U12762 ( .C1(n10083), .C2(n10080), .A(n15493), .B(n10079), .ZN(
        n10874) );
  AOI21_X2 U12763 ( .B1(n15490), .B2(n10090), .A(n10089), .ZN(n15453) );
  AND2_X2 U12764 ( .A1(n15453), .A2(n10892), .ZN(n10957) );
  NAND2_X1 U12765 ( .A1(n10613), .A2(n10612), .ZN(n14340) );
  NOR2_X2 U12766 ( .A1(n10095), .A2(n15792), .ZN(n10481) );
  INV_X1 U12767 ( .A(n10276), .ZN(n10098) );
  NAND2_X2 U12768 ( .A1(n13298), .A2(n10531), .ZN(n10275) );
  INV_X1 U12769 ( .A(n11060), .ZN(n13148) );
  NAND2_X1 U12770 ( .A1(n11025), .A2(n11060), .ZN(n10099) );
  AND2_X1 U12771 ( .A1(n11011), .A2(n10109), .ZN(n14541) );
  NAND2_X1 U12772 ( .A1(n11011), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11010) );
  AND2_X1 U12773 ( .A1(n10217), .A2(n19149), .ZN(n19674) );
  INV_X1 U12774 ( .A(n10531), .ZN(n10168) );
  NAND2_X1 U12775 ( .A1(n11617), .A2(n11616), .ZN(n11618) );
  OR2_X2 U12776 ( .A1(n11617), .A2(n11616), .ZN(n11651) );
  NAND2_X1 U12777 ( .A1(n15177), .A2(n15435), .ZN(n15178) );
  XNOR2_X1 U12778 ( .A(n10961), .B(n10960), .ZN(n12848) );
  AND2_X1 U12779 ( .A1(n10374), .A2(n15811), .ZN(n10444) );
  AOI22_X1 U12780 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9597), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10156) );
  AOI22_X2 U12781 ( .A1(n11048), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19840), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10268) );
  AOI22_X1 U12782 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11337) );
  NAND2_X1 U12783 ( .A1(n13168), .A2(n13171), .ZN(n14548) );
  AND2_X4 U12785 ( .A1(n11321), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13638) );
  NAND2_X1 U12786 ( .A1(n13169), .A2(n13170), .ZN(n13168) );
  OR2_X1 U12787 ( .A1(n13170), .A2(n13169), .ZN(n13171) );
  INV_X1 U12788 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14135) );
  NAND2_X1 U12789 ( .A1(n19822), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10526) );
  AND2_X1 U12790 ( .A1(n10337), .A2(n10336), .ZN(n10338) );
  AND2_X1 U12791 ( .A1(n10337), .A2(n10331), .ZN(n10330) );
  INV_X1 U12792 ( .A(n14196), .ZN(n10751) );
  INV_X1 U12793 ( .A(n10758), .ZN(n10750) );
  NAND2_X1 U12794 ( .A1(n11060), .A2(n11021), .ZN(n10967) );
  OAI21_X1 U12795 ( .B1(n14540), .B2(n19992), .A(n12510), .ZN(P1_U2842) );
  XNOR2_X1 U12796 ( .A(n11064), .B(n11065), .ZN(n13757) );
  NAND2_X1 U12797 ( .A1(n14489), .A2(n12543), .ZN(n12544) );
  AND2_X1 U12798 ( .A1(n13207), .A2(n18923), .ZN(n10114) );
  INV_X1 U12799 ( .A(n13212), .ZN(n13214) );
  AND4_X1 U12800 ( .A1(n10585), .A2(n10584), .A3(n10583), .A4(n10582), .ZN(
        n10115) );
  AND2_X1 U12801 ( .A1(n11258), .A2(n11252), .ZN(n16298) );
  INV_X1 U12802 ( .A(n16298), .ZN(n19143) );
  INV_X1 U12803 ( .A(n15572), .ZN(n11276) );
  AND4_X1 U12804 ( .A1(n15579), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15581), .A4(n10855), .ZN(n10116) );
  AND2_X2 U12805 ( .A1(n12467), .A2(n13280), .ZN(n19997) );
  INV_X1 U12806 ( .A(n19997), .ZN(n12469) );
  INV_X1 U12807 ( .A(n19985), .ZN(n12508) );
  OR2_X1 U12808 ( .A1(n10782), .A2(n10781), .ZN(n10117) );
  OR2_X1 U12809 ( .A1(n15316), .A2(n13182), .ZN(n10118) );
  AND2_X1 U12810 ( .A1(n11967), .A2(n11502), .ZN(n10119) );
  OR2_X1 U12811 ( .A1(n14548), .A2(n19143), .ZN(n10120) );
  NOR3_X1 U12812 ( .A1(n16368), .A2(n19848), .A3(n10302), .ZN(n10121) );
  AND4_X1 U12813 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        n10123) );
  AND2_X1 U12814 ( .A1(n11879), .A2(n10119), .ZN(n10124) );
  NAND2_X2 U12815 ( .A1(n14867), .A2(n13619), .ZN(n14869) );
  NOR3_X1 U12816 ( .A1(n9595), .A2(n20573), .A3(n20742), .ZN(n10125) );
  NOR2_X1 U12817 ( .A1(n9595), .A2(n20059), .ZN(n10126) );
  AND2_X1 U12818 ( .A1(n11561), .A2(n11620), .ZN(n10127) );
  AND2_X1 U12819 ( .A1(n11058), .A2(n11057), .ZN(n10128) );
  OR2_X1 U12820 ( .A1(n14872), .A2(n11780), .ZN(n10129) );
  INV_X1 U12821 ( .A(n10357), .ZN(n10352) );
  INV_X1 U12822 ( .A(n20573), .ZN(n20718) );
  NAND2_X1 U12823 ( .A1(n12409), .A2(n20338), .ZN(n20573) );
  INV_X1 U12824 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12799) );
  INV_X1 U12825 ( .A(n15316), .ZN(n13618) );
  INV_X1 U12826 ( .A(n11787), .ZN(n13478) );
  INV_X1 U12827 ( .A(n15012), .ZN(n12509) );
  INV_X1 U12828 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12781) );
  INV_X1 U12829 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11803) );
  INV_X1 U12830 ( .A(n15475), .ZN(n10883) );
  AND2_X1 U12831 ( .A1(n10160), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10131) );
  INV_X1 U12832 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12780) );
  INV_X1 U12833 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16206) );
  INV_X1 U12834 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19813) );
  AND2_X1 U12835 ( .A1(n10165), .A2(n10192), .ZN(n10132) );
  AND4_X1 U12836 ( .A1(n10171), .A2(n10170), .A3(n10192), .A4(n10169), .ZN(
        n10133) );
  AND2_X1 U12837 ( .A1(n13069), .A2(n13087), .ZN(n10134) );
  INV_X1 U12838 ( .A(n19060), .ZN(n13149) );
  INV_X1 U12839 ( .A(n19717), .ZN(n18984) );
  AND2_X1 U12840 ( .A1(n10176), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10135) );
  NAND2_X1 U12841 ( .A1(n10800), .A2(n10799), .ZN(n10136) );
  OR2_X1 U12842 ( .A1(n12968), .A2(n12967), .ZN(n10137) );
  OR2_X1 U12843 ( .A1(n17743), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10138) );
  AND3_X1 U12844 ( .A1(n10209), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10208), .ZN(n10139) );
  NOR2_X1 U12845 ( .A1(n15521), .A2(n15520), .ZN(n10140) );
  INV_X1 U12846 ( .A(n18995), .ZN(n13236) );
  INV_X1 U12847 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13474) );
  CLKBUF_X3 U12848 ( .A(n12717), .Z(n17148) );
  AND2_X1 U12849 ( .A1(n10174), .A2(n10173), .ZN(n10141) );
  XOR2_X1 U12850 ( .A(n10906), .B(n10902), .Z(n10142) );
  INV_X1 U12851 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20338) );
  INV_X1 U12852 ( .A(n10784), .ZN(n10943) );
  INV_X1 U12853 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n13325) );
  AND2_X1 U12854 ( .A1(n11414), .A2(n11413), .ZN(n10143) );
  AND4_X1 U12855 ( .A1(n11343), .A2(n11342), .A3(n11341), .A4(n11340), .ZN(
        n10144) );
  AND2_X1 U12856 ( .A1(n14668), .A2(n14669), .ZN(n10145) );
  AND4_X1 U12857 ( .A1(n11411), .A2(n11410), .A3(n11409), .A4(n11408), .ZN(
        n10146) );
  INV_X1 U12858 ( .A(n11854), .ZN(n11855) );
  OR2_X1 U12859 ( .A1(n11496), .A2(n12464), .ZN(n11478) );
  INV_X1 U12860 ( .A(n19359), .ZN(n10578) );
  AND2_X1 U12861 ( .A1(n11536), .A2(n11381), .ZN(n11357) );
  INV_X1 U12862 ( .A(n13637), .ZN(n11335) );
  OR2_X1 U12863 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n11803), .ZN(
        n11794) );
  NAND2_X1 U12864 ( .A1(n10269), .A2(n19154), .ZN(n10247) );
  NAND2_X1 U12865 ( .A1(n11422), .A2(n11477), .ZN(n11379) );
  INV_X1 U12866 ( .A(n11419), .ZN(n11404) );
  AND3_X1 U12867 ( .A1(n11578), .A2(n11577), .A3(n11576), .ZN(n11579) );
  INV_X1 U12868 ( .A(n11483), .ZN(n11476) );
  INV_X1 U12869 ( .A(n11530), .ZN(n11531) );
  AND2_X1 U12870 ( .A1(n13070), .A2(n10134), .ZN(n13071) );
  NAND2_X1 U12871 ( .A1(n13016), .A2(n13033), .ZN(n13017) );
  NAND2_X1 U12872 ( .A1(n10376), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10236) );
  INV_X1 U12873 ( .A(n11056), .ZN(n11058) );
  AOI21_X1 U12874 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18638), .A(
        n12547), .ZN(n12552) );
  INV_X1 U12875 ( .A(n11669), .ZN(n11668) );
  INV_X1 U12876 ( .A(n12327), .ZN(n12328) );
  INV_X1 U12877 ( .A(n14660), .ZN(n12301) );
  NOR2_X1 U12878 ( .A1(n10607), .A2(n10606), .ZN(n11090) );
  INV_X1 U12879 ( .A(n19154), .ZN(n11025) );
  AND2_X1 U12880 ( .A1(n10201), .A2(n10192), .ZN(n10206) );
  AOI21_X1 U12881 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n18670), .A(
        n12548), .ZN(n12549) );
  NOR2_X1 U12882 ( .A1(n12561), .A2(n12563), .ZN(n12690) );
  INV_X1 U12883 ( .A(n14722), .ZN(n12172) );
  INV_X1 U12884 ( .A(n12370), .ZN(n12371) );
  AND2_X1 U12885 ( .A1(n12328), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12329) );
  INV_X1 U12886 ( .A(n14682), .ZN(n12235) );
  OR2_X1 U12887 ( .A1(n14333), .A2(n12127), .ZN(n14733) );
  OR2_X1 U12888 ( .A1(n11529), .A2(n11528), .ZN(n11619) );
  NAND2_X1 U12889 ( .A1(n11854), .A2(n11875), .ZN(n12514) );
  AND2_X1 U12890 ( .A1(n10164), .A2(n10163), .ZN(n10167) );
  AND2_X1 U12891 ( .A1(n13086), .A2(n13085), .ZN(n13088) );
  INV_X1 U12892 ( .A(n15698), .ZN(n10769) );
  AND2_X1 U12893 ( .A1(n15204), .A2(n11094), .ZN(n10955) );
  INV_X1 U12894 ( .A(n10926), .ZN(n10934) );
  AND4_X1 U12895 ( .A1(n10524), .A2(n10523), .A3(n10522), .A4(n10521), .ZN(
        n10628) );
  INV_X1 U12896 ( .A(n16229), .ZN(n10764) );
  OAI21_X1 U12897 ( .B1(n13298), .B2(n13325), .A(n19839), .ZN(n12873) );
  NAND2_X1 U12898 ( .A1(n17743), .A2(n12782), .ZN(n12783) );
  NOR2_X1 U12899 ( .A1(n17331), .A2(n12821), .ZN(n12805) );
  INV_X1 U12900 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n20845) );
  AND2_X1 U12901 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n12024), .ZN(
        n12033) );
  OR2_X1 U12902 ( .A1(n12414), .A2(n14592), .ZN(n12454) );
  OR2_X1 U12903 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n12035) );
  NAND2_X1 U12904 ( .A1(n12109), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12139) );
  NAND2_X1 U12905 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12025) );
  OAI21_X1 U12906 ( .B1(n20748), .B2(n13672), .A(n20705), .ZN(n20060) );
  INV_X1 U12907 ( .A(n10142), .ZN(n13237) );
  AND2_X1 U12908 ( .A1(n10815), .A2(n10814), .ZN(n13733) );
  NAND2_X1 U12909 ( .A1(n10957), .A2(n10955), .ZN(n10952) );
  NOR2_X1 U12910 ( .A1(n15610), .A2(n11273), .ZN(n15579) );
  OR2_X1 U12911 ( .A1(n15891), .A2(n10628), .ZN(n10873) );
  INV_X1 U12912 ( .A(n14255), .ZN(n15685) );
  NAND2_X1 U12913 ( .A1(n10610), .A2(n13895), .ZN(n10611) );
  INV_X2 U12914 ( .A(n11077), .ZN(n11224) );
  NOR2_X1 U12915 ( .A1(n17844), .A2(n17803), .ZN(n17577) );
  NOR2_X1 U12916 ( .A1(n18025), .A2(n18000), .ZN(n17664) );
  NOR2_X1 U12917 ( .A1(n15879), .A2(n16428), .ZN(n18026) );
  NOR2_X1 U12918 ( .A1(n12823), .A2(n17788), .ZN(n12825) );
  INV_X1 U12919 ( .A(n9635), .ZN(n15823) );
  AND2_X1 U12920 ( .A1(n11854), .A2(n20061), .ZN(n11866) );
  OR2_X1 U12921 ( .A1(n14599), .A2(n14508), .ZN(n14532) );
  OR2_X1 U12922 ( .A1(n19942), .A2(n14501), .ZN(n14696) );
  INV_X1 U12923 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15991) );
  OR2_X1 U12924 ( .A1(n19972), .A2(n14563), .ZN(n19918) );
  OR2_X1 U12925 ( .A1(n19972), .A2(n20338), .ZN(n19975) );
  INV_X1 U12926 ( .A(n14834), .ZN(n14855) );
  INV_X1 U12927 ( .A(n11760), .ZN(n14968) );
  OR2_X1 U12928 ( .A1(n11778), .A2(n15941), .ZN(n11781) );
  AND2_X1 U12929 ( .A1(n11941), .A2(n11940), .ZN(n15945) );
  NOR2_X1 U12930 ( .A1(n15097), .A2(n13550), .ZN(n16092) );
  NAND2_X1 U12931 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n13444), .ZN(n20705) );
  OR2_X1 U12932 ( .A1(n11999), .A2(n20211), .ZN(n20305) );
  AND2_X1 U12933 ( .A1(n20536), .A2(n20216), .ZN(n20391) );
  NAND2_X1 U12934 ( .A1(n20744), .A2(n20060), .ZN(n20114) );
  NOR2_X1 U12935 ( .A1(n16337), .A2(n16336), .ZN(n16350) );
  AND2_X1 U12936 ( .A1(n10805), .A2(n10804), .ZN(n13572) );
  NAND2_X1 U12937 ( .A1(n12881), .A2(n12878), .ZN(n13579) );
  NAND2_X1 U12938 ( .A1(n13103), .A2(n13102), .ZN(n15283) );
  NAND2_X1 U12939 ( .A1(n19041), .A2(n13162), .ZN(n15410) );
  AND2_X1 U12940 ( .A1(n19041), .A2(n13150), .ZN(n13378) );
  OAI21_X1 U12941 ( .B1(n13159), .B2(n13158), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13160) );
  AND2_X1 U12942 ( .A1(n11317), .A2(n11316), .ZN(n11318) );
  INV_X1 U12943 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11275) );
  AND2_X1 U12944 ( .A1(n10975), .A2(n10974), .ZN(n11016) );
  INV_X1 U12945 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14051) );
  INV_X1 U12946 ( .A(n19395), .ZN(n19392) );
  AND2_X1 U12947 ( .A1(n19359), .A2(n19358), .ZN(n19364) );
  NAND2_X1 U12948 ( .A1(n19804), .A2(n19816), .ZN(n19420) );
  OR2_X1 U12949 ( .A1(n19804), .A2(n19268), .ZN(n19583) );
  INV_X1 U12950 ( .A(n19166), .ZN(n19149) );
  NOR2_X1 U12951 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16684), .ZN(n16674) );
  NOR2_X1 U12952 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16734), .ZN(n16716) );
  NOR2_X1 U12953 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16853), .ZN(n16834) );
  INV_X1 U12954 ( .A(n16869), .ZN(n16909) );
  AND2_X1 U12955 ( .A1(n17649), .A2(n16581), .ZN(n12842) );
  INV_X1 U12956 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17574) );
  NOR2_X1 U12957 ( .A1(n17712), .A2(n18003), .ZN(n17686) );
  NOR2_X1 U12958 ( .A1(n17627), .A2(n12784), .ZN(n17702) );
  INV_X1 U12959 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17777) );
  INV_X1 U12960 ( .A(n17577), .ZN(n17500) );
  INV_X1 U12961 ( .A(n17914), .ZN(n17993) );
  INV_X1 U12962 ( .A(n17670), .ZN(n18003) );
  INV_X1 U12963 ( .A(n18026), .ZN(n18045) );
  NOR2_X1 U12964 ( .A1(n18095), .A2(n17770), .ZN(n17769) );
  NOR2_X1 U12965 ( .A1(n17823), .A2(n12727), .ZN(n17813) );
  INV_X1 U12966 ( .A(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n20795) );
  AOI211_X1 U12967 ( .C1(n17132), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n12635), .B(n12634), .ZN(n12636) );
  AOI21_X1 U12968 ( .B1(n12839), .B2(n18173), .A(n18815), .ZN(n18184) );
  OR2_X1 U12969 ( .A1(n20634), .A2(n20744), .ZN(n19862) );
  OR2_X1 U12970 ( .A1(n15968), .A2(n14505), .ZN(n14640) );
  NOR2_X1 U12971 ( .A1(n20672), .A2(n14696), .ZN(n14692) );
  INV_X1 U12972 ( .A(n19975), .ZN(n19959) );
  NOR2_X1 U12973 ( .A1(n19997), .A2(n12506), .ZN(n12507) );
  INV_X1 U12974 ( .A(n14065), .ZN(n14166) );
  INV_X1 U12975 ( .A(n13588), .ZN(n20037) );
  INV_X1 U12976 ( .A(n13596), .ZN(n20026) );
  NAND2_X1 U12977 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12268), .ZN(
        n12327) );
  INV_X1 U12978 ( .A(n16069), .ZN(n16055) );
  INV_X1 U12979 ( .A(n19869), .ZN(n16065) );
  NOR2_X1 U12980 ( .A1(n16090), .A2(n16089), .ZN(n15138) );
  NOR2_X1 U12981 ( .A1(n11987), .A2(n13643), .ZN(n15097) );
  INV_X1 U12982 ( .A(n16134), .ZN(n16118) );
  NOR2_X2 U12983 ( .A1(n11987), .A2(n11865), .ZN(n16122) );
  INV_X1 U12984 ( .A(n20114), .ZN(n20216) );
  OAI22_X1 U12985 ( .A1(n20073), .A2(n20072), .B1(n20394), .B2(n20213), .ZN(
        n20108) );
  INV_X1 U12986 ( .A(n20167), .ZN(n20138) );
  OAI22_X1 U12987 ( .A1(n20145), .A2(n20144), .B1(n20394), .B2(n20272), .ZN(
        n20169) );
  NAND2_X1 U12988 ( .A1(n20719), .A2(n11999), .ZN(n20175) );
  INV_X1 U12989 ( .A(n20265), .ZN(n20254) );
  OAI22_X1 U12990 ( .A1(n20274), .A2(n20273), .B1(n20272), .B2(n20536), .ZN(
        n20297) );
  NOR2_X1 U12991 ( .A1(n20499), .A2(n20303), .ZN(n20324) );
  INV_X1 U12992 ( .A(n20330), .ZN(n20355) );
  INV_X1 U12993 ( .A(n20423), .ZN(n20380) );
  OAI22_X1 U12994 ( .A1(n20396), .A2(n20395), .B1(n20394), .B2(n20535), .ZN(
        n20419) );
  OAI22_X1 U12995 ( .A1(n20464), .A2(n20463), .B1(n20462), .B2(n20536), .ZN(
        n20494) );
  OR2_X1 U12996 ( .A1(n20719), .A2(n20331), .ZN(n20432) );
  OAI21_X1 U12997 ( .B1(n20504), .B2(n20503), .A(n20581), .ZN(n20529) );
  NOR2_X2 U12998 ( .A1(n20580), .A2(n20505), .ZN(n20567) );
  INV_X1 U12999 ( .A(n16145), .ZN(n13672) );
  AND2_X1 U13000 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_1__SCAN_IN), 
        .ZN(n20646) );
  INV_X1 U13001 ( .A(n20695), .ZN(n20689) );
  NAND2_X1 U13002 ( .A1(n13239), .A2(n13238), .ZN(n13240) );
  INV_X1 U13003 ( .A(n18951), .ZN(n18987) );
  NOR2_X1 U13004 ( .A1(n9951), .A2(n13206), .ZN(n18922) );
  AND2_X1 U13005 ( .A1(n19841), .A2(n13226), .ZN(n18951) );
  INV_X1 U13006 ( .A(n18989), .ZN(n18954) );
  OR2_X1 U13007 ( .A1(n11223), .A2(n11222), .ZN(n13955) );
  INV_X1 U13008 ( .A(n13384), .ZN(n13385) );
  OR2_X1 U13009 ( .A1(n12942), .A2(n12941), .ZN(n15346) );
  AND2_X1 U13010 ( .A1(n13378), .A2(n14278), .ZN(n19010) );
  INV_X1 U13011 ( .A(n19041), .ZN(n19055) );
  OAI21_X1 U13012 ( .B1(n12855), .B2(n16256), .A(n12854), .ZN(n12856) );
  INV_X1 U13013 ( .A(n16265), .ZN(n19114) );
  INV_X1 U13014 ( .A(n19138), .ZN(n16302) );
  AND2_X1 U13015 ( .A1(n15789), .A2(n11040), .ZN(n16268) );
  AND2_X1 U13016 ( .A1(n16310), .A2(n16308), .ZN(n15789) );
  INV_X1 U13017 ( .A(n19137), .ZN(n16271) );
  INV_X1 U13018 ( .A(n15766), .ZN(n15797) );
  INV_X1 U13019 ( .A(n18986), .ZN(n19825) );
  OAI21_X1 U13020 ( .B1(n14282), .B2(n14281), .A(n14280), .ZN(n19172) );
  INV_X1 U13021 ( .A(n19263), .ZN(n19249) );
  INV_X1 U13022 ( .A(n19273), .ZN(n19291) );
  INV_X1 U13023 ( .A(n19309), .ZN(n19323) );
  AND2_X1 U13024 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19361), .ZN(
        n19395) );
  INV_X1 U13025 ( .A(n19419), .ZN(n19411) );
  OAI21_X1 U13026 ( .B1(n19428), .B2(n19427), .A(n19426), .ZN(n19445) );
  INV_X1 U13027 ( .A(n19474), .ZN(n19536) );
  INV_X1 U13028 ( .A(n19790), .ZN(n19481) );
  INV_X1 U13029 ( .A(n19597), .ZN(n19606) );
  OAI21_X1 U13030 ( .B1(n19622), .B2(n19621), .A(n19620), .ZN(n19651) );
  INV_X1 U13031 ( .A(n19521), .ZN(n19691) );
  INV_X1 U13032 ( .A(n19796), .ZN(n19610) );
  NOR2_X1 U13033 ( .A1(n10302), .A2(n19848), .ZN(n14270) );
  INV_X1 U13034 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19740) );
  INV_X1 U13035 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19722) );
  NOR2_X1 U13036 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16621), .ZN(n16620) );
  NOR2_X1 U13037 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16665), .ZN(n16660) );
  NOR2_X1 U13038 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16758), .ZN(n16739) );
  NOR2_X1 U13039 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16779), .ZN(n16762) );
  NOR2_X1 U13040 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16801), .ZN(n16789) );
  NOR2_X2 U13041 ( .A1(n18794), .A2(n16919), .ZN(n16879) );
  NOR2_X2 U13042 ( .A1(n18680), .A2(n13260), .ZN(n16869) );
  INV_X1 U13043 ( .A(n16807), .ZN(n16919) );
  INV_X1 U13044 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17123) );
  NOR2_X1 U13045 ( .A1(n17362), .A2(n17233), .ZN(n17228) );
  NOR2_X1 U13046 ( .A1(n18225), .A2(n17243), .ZN(n17239) );
  NOR3_X1 U13047 ( .A1(n18225), .A2(n17283), .A3(n17421), .ZN(n17275) );
  AND2_X1 U13048 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17323), .ZN(n17312) );
  NAND3_X1 U13049 ( .A1(n12687), .A2(n12686), .A3(n12685), .ZN(n15879) );
  NOR2_X1 U13050 ( .A1(n17465), .A2(n18842), .ZN(n17466) );
  NOR2_X1 U13051 ( .A1(n17969), .A2(n17741), .ZN(n17620) );
  NOR2_X1 U13052 ( .A1(n12835), .A2(n17751), .ZN(n17711) );
  AOI21_X1 U13053 ( .B1(n15851), .B2(n18838), .A(n16538), .ZN(n17803) );
  NOR2_X1 U13054 ( .A1(n17535), .A2(n17894), .ZN(n17510) );
  INV_X1 U13055 ( .A(n18120), .ZN(n18081) );
  INV_X1 U13056 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18000) );
  NOR2_X2 U13057 ( .A1(n18169), .A2(n17321), .ZN(n18072) );
  NAND2_X1 U13058 ( .A1(n12668), .A2(n13253), .ZN(n18658) );
  INV_X1 U13059 ( .A(n18171), .ZN(n18152) );
  INV_X1 U13060 ( .A(n18282), .ZN(n20755) );
  INV_X1 U13061 ( .A(n20761), .ZN(n18346) );
  INV_X1 U13062 ( .A(n18369), .ZN(n18371) );
  INV_X1 U13063 ( .A(n15862), .ZN(n18200) );
  INV_X1 U13064 ( .A(n18445), .ZN(n18447) );
  INV_X1 U13065 ( .A(n17353), .ZN(n18185) );
  INV_X1 U13066 ( .A(n12657), .ZN(n18207) );
  INV_X1 U13067 ( .A(n18540), .ZN(n18557) );
  INV_X1 U13068 ( .A(n18579), .ZN(n18614) );
  INV_X1 U13069 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18705) );
  NAND2_X1 U13070 ( .A1(n15927), .A2(n13463), .ZN(n14564) );
  AND2_X1 U13071 ( .A1(n14562), .A2(n14564), .ZN(n20738) );
  INV_X1 U13072 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20742) );
  OR2_X1 U13073 ( .A1(n14621), .A2(n14506), .ZN(n14599) );
  OR3_X1 U13074 ( .A1(n19972), .A2(n16149), .A3(n14492), .ZN(n19903) );
  INV_X1 U13075 ( .A(n19971), .ZN(n19968) );
  NAND2_X1 U13076 ( .A1(n19997), .A2(n14525), .ZN(n19985) );
  OR2_X1 U13077 ( .A1(n13740), .A2(n13535), .ZN(n19977) );
  OR2_X1 U13078 ( .A1(n14861), .A2(n13619), .ZN(n14866) );
  INV_X1 U13079 ( .A(n19998), .ZN(n20019) );
  NOR2_X1 U13080 ( .A1(n14564), .A2(n13388), .ZN(n13596) );
  OR2_X1 U13081 ( .A1(n16060), .A2(n13785), .ZN(n16069) );
  OR2_X1 U13082 ( .A1(n15051), .A2(n11993), .ZN(n15046) );
  INV_X1 U13083 ( .A(n16122), .ZN(n16137) );
  INV_X1 U13084 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20727) );
  NAND2_X1 U13085 ( .A1(n20057), .A2(n10126), .ZN(n20136) );
  OR2_X1 U13086 ( .A1(n20175), .A2(n20505), .ZN(n20167) );
  OR2_X1 U13087 ( .A1(n20175), .A2(n20385), .ZN(n20205) );
  OR2_X1 U13088 ( .A1(n20175), .A2(n20431), .ZN(n20230) );
  NAND2_X1 U13089 ( .A1(n20714), .A2(n10126), .ZN(n20265) );
  NAND2_X1 U13090 ( .A1(n20714), .A2(n20243), .ZN(n20301) );
  NAND2_X1 U13091 ( .A1(n20714), .A2(n20308), .ZN(n20330) );
  NAND2_X1 U13092 ( .A1(n20332), .A2(n10126), .ZN(n20384) );
  OR2_X1 U13093 ( .A1(n20432), .A2(n20505), .ZN(n20423) );
  OR2_X1 U13094 ( .A1(n20432), .A2(n20385), .ZN(n20448) );
  OR2_X1 U13095 ( .A1(n20432), .A2(n20431), .ZN(n20498) );
  NAND2_X1 U13096 ( .A1(n20534), .A2(n10126), .ZN(n20532) );
  NAND2_X1 U13097 ( .A1(n20534), .A2(n20308), .ZN(n20621) );
  INV_X1 U13098 ( .A(n20704), .ZN(n20637) );
  INV_X1 U13099 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20650) );
  INV_X1 U13100 ( .A(n20675), .ZN(n20752) );
  NOR2_X1 U13101 ( .A1(n13241), .A2(n13240), .ZN(n13242) );
  OR3_X1 U13102 ( .A1(n13224), .A2(n13223), .A3(n13229), .ZN(n18995) );
  OR2_X1 U13103 ( .A1(n13224), .A2(n13222), .ZN(n18978) );
  AND2_X1 U13104 ( .A1(n13178), .A2(n13220), .ZN(n15316) );
  XNOR2_X1 U13105 ( .A(n13524), .B(n13523), .ZN(n19804) );
  AND2_X1 U13106 ( .A1(n13147), .A2(n13220), .ZN(n19041) );
  NAND2_X1 U13107 ( .A1(n19041), .A2(n13148), .ZN(n19060) );
  OR2_X1 U13108 ( .A1(n19104), .A2(n13324), .ZN(n19067) );
  NAND2_X1 U13109 ( .A1(n13323), .A2(n19845), .ZN(n19104) );
  OR2_X1 U13110 ( .A1(n13275), .A2(n13297), .ZN(n13532) );
  OAI21_X1 U13111 ( .B1(n11283), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11282), .ZN(n15447) );
  INV_X1 U13112 ( .A(n10850), .ZN(n10851) );
  INV_X1 U13113 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16189) );
  INV_X1 U13114 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16227) );
  INV_X1 U13115 ( .A(n16255), .ZN(n19125) );
  NOR2_X1 U13116 ( .A1(n11278), .A2(n11277), .ZN(n11279) );
  NAND2_X1 U13117 ( .A1(n11258), .A2(n11009), .ZN(n19133) );
  INV_X1 U13118 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15860) );
  AOI211_X2 U13119 ( .C1(n14275), .C2(n14281), .A(n14274), .B(n19363), .ZN(
        n19176) );
  INV_X1 U13120 ( .A(n19229), .ZN(n19218) );
  OR2_X1 U13121 ( .A1(n19327), .A2(n19481), .ZN(n19263) );
  INV_X1 U13122 ( .A(n19286), .ZN(n19294) );
  INV_X1 U13123 ( .A(n19332), .ZN(n19389) );
  OR2_X1 U13124 ( .A1(n19796), .A2(n19367), .ZN(n19419) );
  NAND2_X1 U13125 ( .A1(n19611), .A2(n19422), .ZN(n19449) );
  OR2_X1 U13126 ( .A1(n19584), .A2(n19481), .ZN(n19571) );
  AND2_X1 U13127 ( .A1(n19579), .A2(n19578), .ZN(n19597) );
  INV_X1 U13128 ( .A(n19699), .ZN(n19604) );
  INV_X1 U13129 ( .A(n19693), .ZN(n19643) );
  NAND2_X1 U13130 ( .A1(n19611), .A2(n19610), .ZN(n19712) );
  INV_X2 U13131 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19839) );
  INV_X1 U13132 ( .A(n19789), .ZN(n19720) );
  OR2_X1 U13133 ( .A1(n19722), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n19859) );
  INV_X1 U13134 ( .A(n18780), .ZN(n18851) );
  INV_X1 U13135 ( .A(n16879), .ZN(n16907) );
  AND2_X1 U13136 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17301), .ZN(n17304) );
  NOR2_X1 U13137 ( .A1(n12762), .A2(n12761), .ZN(n17328) );
  INV_X1 U13138 ( .A(n17348), .ZN(n17343) );
  OR2_X1 U13139 ( .A1(n17413), .A2(n17353), .ZN(n17381) );
  NAND2_X1 U13140 ( .A1(n17415), .A2(n17352), .ZN(n17413) );
  INV_X1 U13141 ( .A(n17466), .ZN(n17458) );
  NAND3_X1 U13142 ( .A1(n18841), .A2(n17843), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n17696) );
  AOI22_X1 U13143 ( .A1(n18044), .A2(n17837), .B1(n17753), .B2(n18046), .ZN(
        n17741) );
  INV_X1 U13144 ( .A(n17738), .ZN(n17756) );
  INV_X1 U13145 ( .A(n17803), .ZN(n17843) );
  OR2_X1 U13146 ( .A1(n17931), .A2(n17930), .ZN(n17957) );
  INV_X1 U13147 ( .A(n18122), .ZN(n18153) );
  INV_X1 U13148 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18042) );
  INV_X1 U13149 ( .A(n18072), .ZN(n18091) );
  NAND2_X1 U13150 ( .A1(n18162), .A2(n18623), .ZN(n18169) );
  INV_X1 U13151 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18631) );
  INV_X1 U13152 ( .A(n18599), .ZN(n20762) );
  INV_X1 U13153 ( .A(n18679), .ZN(n18839) );
  INV_X1 U13154 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18794) );
  INV_X1 U13155 ( .A(n18702), .ZN(n18790) );
  INV_X1 U13156 ( .A(n18851), .ZN(n18786) );
  INV_X1 U13157 ( .A(n18851), .ZN(n18850) );
  NOR2_X1 U13158 ( .A1(n18705), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18780) );
  NOR2_X1 U13159 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13248), .ZN(n16525)
         );
  INV_X1 U13160 ( .A(n16491), .ZN(n16494) );
  NAND2_X1 U13161 ( .A1(n12847), .A2(n12846), .ZN(P3_U2800) );
  INV_X2 U13162 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13965) );
  AND2_X4 U13163 ( .A1(n14054), .A2(n13965), .ZN(n10376) );
  AOI22_X1 U13164 ( .A1(n9597), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10147) );
  AND2_X1 U13165 ( .A1(n10147), .A2(n15811), .ZN(n10152) );
  AND2_X2 U13166 ( .A1(n14135), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10148) );
  AND2_X4 U13167 ( .A1(n10148), .A2(n16322), .ZN(n10374) );
  AND2_X4 U13168 ( .A1(n10148), .A2(n10528), .ZN(n10241) );
  AOI22_X1 U13169 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10241), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10151) );
  AND2_X4 U13170 ( .A1(n14053), .A2(n16322), .ZN(n13002) );
  AOI22_X1 U13171 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10150) );
  AND3_X4 U13172 ( .A1(n10528), .A2(n13965), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10375) );
  AOI22_X1 U13173 ( .A1(n10225), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10149) );
  AOI22_X1 U13174 ( .A1(n10241), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10153) );
  AND2_X1 U13175 ( .A1(n10153), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10157) );
  AOI22_X1 U13176 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10235), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U13177 ( .A1(n10225), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10154) );
  AOI22_X1 U13178 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10159) );
  AOI22_X1 U13179 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10235), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10158) );
  AOI22_X1 U13180 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10161) );
  AOI22_X1 U13181 ( .A1(n10241), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10225), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10160) );
  AOI22_X1 U13182 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10164) );
  AOI22_X1 U13183 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10235), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U13184 ( .A1(n10241), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10225), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10165) );
  AOI22_X1 U13185 ( .A1(n9597), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10166) );
  AOI22_X1 U13186 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U13187 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10241), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10171) );
  AOI22_X1 U13188 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10170) );
  AOI22_X1 U13189 ( .A1(n10225), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10169) );
  AOI22_X1 U13190 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10241), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U13191 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10235), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10173) );
  AOI22_X1 U13192 ( .A1(n10225), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U13193 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10241), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10182) );
  AOI22_X1 U13194 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10181) );
  AOI22_X1 U13195 ( .A1(n10225), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10180) );
  NAND4_X1 U13196 ( .A1(n10182), .A2(n10181), .A3(n10180), .A4(n10179), .ZN(
        n10183) );
  AOI22_X1 U13197 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9586), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U13198 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10241), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10186) );
  AOI22_X1 U13199 ( .A1(n10225), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10185) );
  AOI22_X1 U13200 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10184) );
  NAND4_X1 U13201 ( .A1(n10187), .A2(n10186), .A3(n10185), .A4(n10184), .ZN(
        n10188) );
  AOI22_X1 U13202 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10241), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10191) );
  AOI22_X1 U13203 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9586), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U13204 ( .A1(n10225), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10189) );
  NAND3_X1 U13205 ( .A1(n10191), .A2(n10190), .A3(n10189), .ZN(n10193) );
  AOI22_X1 U13206 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10194) );
  AOI22_X1 U13207 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10241), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10199) );
  AOI22_X1 U13208 ( .A1(n10225), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10198) );
  AOI22_X1 U13209 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10235), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10197) );
  AOI22_X1 U13210 ( .A1(n9597), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U13211 ( .A1(n10225), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10207) );
  AOI22_X1 U13212 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10241), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10201) );
  AOI22_X1 U13213 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n10235), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10205) );
  AOI21_X1 U13214 ( .B1(n9590), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A(n10203), .ZN(n10204) );
  NAND4_X1 U13215 ( .A1(n10207), .A2(n10206), .A3(n10205), .A4(n10204), .ZN(
        n10213) );
  AOI22_X1 U13216 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10235), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10209) );
  AOI22_X1 U13217 ( .A1(n10225), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10208) );
  AOI22_X1 U13218 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10241), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10211) );
  AOI22_X1 U13219 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10210) );
  NAND3_X1 U13220 ( .A1(n10139), .A2(n10211), .A3(n10210), .ZN(n10212) );
  NAND2_X2 U13221 ( .A1(n10213), .A2(n10212), .ZN(n10251) );
  INV_X2 U13222 ( .A(n13298), .ZN(n10214) );
  OAI21_X1 U13223 ( .B1(n10233), .B2(n10251), .A(n10215), .ZN(n10216) );
  AND4_X1 U13224 ( .A1(n10217), .A2(n10251), .A3(n19154), .A4(n10214), .ZN(
        n10218) );
  NAND2_X1 U13225 ( .A1(n10218), .A2(n10970), .ZN(n10262) );
  NAND2_X1 U13226 ( .A1(n10219), .A2(n10262), .ZN(n11017) );
  AOI22_X1 U13227 ( .A1(n9597), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10223) );
  AOI22_X1 U13228 ( .A1(n10225), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10222) );
  AOI22_X1 U13229 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10241), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10221) );
  AOI22_X1 U13230 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10220) );
  NAND4_X1 U13231 ( .A1(n10223), .A2(n10222), .A3(n10221), .A4(n10220), .ZN(
        n10224) );
  NAND2_X1 U13232 ( .A1(n10224), .A2(n10192), .ZN(n10232) );
  AOI22_X1 U13233 ( .A1(n9597), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10229) );
  AOI22_X1 U13234 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10241), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10228) );
  AOI22_X1 U13235 ( .A1(n10225), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10227) );
  AOI22_X1 U13236 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10226) );
  NAND4_X1 U13237 ( .A1(n10229), .A2(n10228), .A3(n10227), .A4(n10226), .ZN(
        n10230) );
  NAND2_X1 U13238 ( .A1(n10230), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10231) );
  NOR2_X1 U13239 ( .A1(n13148), .A2(n9600), .ZN(n10234) );
  NAND2_X1 U13240 ( .A1(n11017), .A2(n10288), .ZN(n10246) );
  AOI22_X1 U13241 ( .A1(n10241), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10225), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10240) );
  AOI22_X1 U13242 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10238) );
  AOI22_X1 U13243 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10237) );
  AOI22_X1 U13244 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9597), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10245) );
  AOI22_X1 U13245 ( .A1(n10241), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10244) );
  AOI22_X1 U13246 ( .A1(n10225), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10243) );
  AOI22_X1 U13247 ( .A1(n13002), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10242) );
  NAND2_X1 U13248 ( .A1(n10246), .A2(n19846), .ZN(n10291) );
  NAND3_X1 U13249 ( .A1(n10251), .A2(n10254), .A3(n10275), .ZN(n10971) );
  NAND3_X1 U13250 ( .A1(n10971), .A2(n10967), .A3(n10252), .ZN(n11018) );
  NAND2_X1 U13251 ( .A1(n11018), .A2(n11025), .ZN(n10248) );
  NAND2_X1 U13252 ( .A1(n10290), .A2(n19833), .ZN(n10249) );
  NAND2_X1 U13253 ( .A1(n10291), .A2(n10249), .ZN(n10250) );
  NAND2_X1 U13254 ( .A1(n10250), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10261) );
  NOR2_X4 U13255 ( .A1(n10253), .A2(n10275), .ZN(n10962) );
  INV_X1 U13256 ( .A(n10962), .ZN(n10258) );
  NAND2_X1 U13257 ( .A1(n10256), .A2(n10255), .ZN(n10727) );
  NAND3_X1 U13258 ( .A1(n10727), .A2(n10264), .A3(n9600), .ZN(n10257) );
  NAND2_X1 U13259 ( .A1(n10258), .A2(n10257), .ZN(n11250) );
  INV_X1 U13260 ( .A(n11250), .ZN(n10260) );
  INV_X1 U13261 ( .A(n13324), .ZN(n10259) );
  INV_X1 U13262 ( .A(n10262), .ZN(n10263) );
  NAND4_X1 U13263 ( .A1(n10276), .A2(n10265), .A3(n11027), .A4(n10252), .ZN(
        n10266) );
  NAND2_X1 U13264 ( .A1(n10965), .A2(n10266), .ZN(n10278) );
  NAND2_X1 U13265 ( .A1(n10962), .A2(n10274), .ZN(n13227) );
  INV_X1 U13266 ( .A(n13227), .ZN(n10267) );
  OR2_X2 U13267 ( .A1(n10278), .A2(n10267), .ZN(n11048) );
  NOR2_X2 U13268 ( .A1(n10364), .A2(n13324), .ZN(n10270) );
  NAND2_X4 U13269 ( .A1(n10962), .A2(n10270), .ZN(n10936) );
  INV_X1 U13270 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10272) );
  INV_X2 U13271 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n10302) );
  INV_X1 U13272 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10271) );
  OAI22_X1 U13273 ( .A1(n10936), .A2(n10272), .B1(n10302), .B2(n10271), .ZN(
        n10273) );
  AOI21_X1 U13274 ( .B1(n9598), .B2(P2_EBX_REG_1__SCAN_IN), .A(n10273), .ZN(
        n10280) );
  NAND2_X1 U13275 ( .A1(n11049), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10285) );
  NAND2_X1 U13276 ( .A1(n10282), .A2(n10281), .ZN(n10319) );
  AND3_X1 U13277 ( .A1(n11027), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n19833), 
        .ZN(n10283) );
  OAI22_X1 U13278 ( .A1(n10327), .A2(n10283), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n10926), .ZN(n10287) );
  NAND2_X1 U13279 ( .A1(n19840), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10284) );
  AND2_X1 U13280 ( .A1(n10285), .A2(n10284), .ZN(n10286) );
  NAND2_X1 U13281 ( .A1(n10287), .A2(n10286), .ZN(n10311) );
  INV_X1 U13282 ( .A(n10288), .ZN(n10289) );
  NAND2_X1 U13283 ( .A1(n10290), .A2(n10289), .ZN(n11026) );
  AND2_X1 U13284 ( .A1(n10291), .A2(n11026), .ZN(n10292) );
  NAND2_X1 U13285 ( .A1(n10323), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10298) );
  INV_X1 U13286 ( .A(n19840), .ZN(n10296) );
  NAND2_X1 U13287 ( .A1(n10940), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10295) );
  NAND2_X1 U13288 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10294) );
  NAND2_X2 U13289 ( .A1(n10311), .A2(n10310), .ZN(n10345) );
  NAND2_X1 U13290 ( .A1(n10327), .A2(n16322), .ZN(n10301) );
  AOI21_X1 U13291 ( .B1(n13325), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10300) );
  NAND2_X1 U13292 ( .A1(n10301), .A2(n10300), .ZN(n10308) );
  NAND2_X1 U13293 ( .A1(n10323), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10306) );
  INV_X1 U13294 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n13397) );
  INV_X1 U13295 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10303) );
  OAI22_X1 U13296 ( .A1(n10936), .A2(n13397), .B1(n10302), .B2(n10303), .ZN(
        n10304) );
  AOI21_X1 U13297 ( .B1(n9599), .B2(P2_EBX_REG_2__SCAN_IN), .A(n10304), .ZN(
        n10305) );
  NAND2_X1 U13298 ( .A1(n10306), .A2(n10305), .ZN(n10307) );
  NAND2_X1 U13299 ( .A1(n10308), .A2(n10307), .ZN(n10320) );
  NOR2_X1 U13300 ( .A1(n13963), .A2(n10314), .ZN(n10331) );
  INV_X1 U13301 ( .A(n10320), .ZN(n10317) );
  OAI21_X1 U13302 ( .B1(n10317), .B2(n10316), .A(n10315), .ZN(n10318) );
  INV_X1 U13303 ( .A(n10318), .ZN(n10322) );
  NAND3_X1 U13304 ( .A1(n10345), .A2(n10320), .A3(n10319), .ZN(n10321) );
  NAND2_X1 U13305 ( .A1(n10323), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10326) );
  INV_X1 U13306 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13817) );
  OAI22_X1 U13307 ( .A1(n10936), .A2(n13817), .B1(n10302), .B2(n13984), .ZN(
        n10324) );
  AOI21_X1 U13308 ( .B1(n10926), .B2(P2_EBX_REG_3__SCAN_IN), .A(n10324), .ZN(
        n10325) );
  NAND2_X1 U13309 ( .A1(n10327), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10329) );
  NAND2_X1 U13310 ( .A1(n19840), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10328) );
  XNOR2_X2 U13311 ( .A(n10779), .B(n10778), .ZN(n12870) );
  AOI22_X1 U13312 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19179), .B1(
        n10469), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10344) );
  INV_X1 U13313 ( .A(n10333), .ZN(n10334) );
  NOR2_X1 U13314 ( .A1(n10332), .A2(n10334), .ZN(n10336) );
  AOI22_X1 U13315 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19300), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10343) );
  INV_X1 U13316 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10339) );
  INV_X1 U13317 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10369) );
  INV_X1 U13318 ( .A(n10340), .ZN(n10341) );
  INV_X1 U13319 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10351) );
  INV_X1 U13320 ( .A(n10314), .ZN(n10347) );
  INV_X1 U13321 ( .A(n10345), .ZN(n10346) );
  NAND2_X1 U13322 ( .A1(n10347), .A2(n10346), .ZN(n10348) );
  INV_X1 U13323 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11150) );
  OAI22_X1 U13324 ( .A1(n10351), .A2(n10587), .B1(n10474), .B2(n11150), .ZN(
        n10356) );
  INV_X1 U13325 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10354) );
  INV_X1 U13326 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10353) );
  OAI22_X1 U13327 ( .A1(n10354), .A2(n19330), .B1(n19547), .B2(n10353), .ZN(
        n10355) );
  NOR2_X1 U13328 ( .A1(n10356), .A2(n10355), .ZN(n10362) );
  NOR2_X2 U13329 ( .A1(n10359), .A2(n15792), .ZN(n19454) );
  AOI22_X1 U13330 ( .A1(n19454), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10481), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10361) );
  NOR2_X2 U13331 ( .A1(n10359), .A2(n10358), .ZN(n19396) );
  AOI22_X1 U13332 ( .A1(n19396), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10360) );
  NAND4_X1 U13333 ( .A1(n10363), .A2(n10362), .A3(n10361), .A4(n10360), .ZN(
        n10365) );
  NAND2_X1 U13334 ( .A1(n10365), .A2(n13297), .ZN(n10385) );
  AND2_X2 U13335 ( .A1(n13133), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10460) );
  AOI22_X1 U13336 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10503), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10373) );
  AND2_X2 U13337 ( .A1(n9590), .A2(n15811), .ZN(n10491) );
  AOI22_X1 U13338 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10372) );
  NAND2_X2 U13339 ( .A1(n9596), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12987) );
  NAND2_X1 U13340 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10368) );
  NAND3_X1 U13341 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n16322), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10717) );
  INV_X1 U13342 ( .A(n10717), .ZN(n10366) );
  AND2_X2 U13343 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10366), .ZN(
        n12983) );
  INV_X2 U13344 ( .A(n11180), .ZN(n12982) );
  AOI22_X1 U13345 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__3__SCAN_IN), .B2(n12982), .ZN(n10367) );
  OAI211_X1 U13346 ( .C1(n12987), .C2(n10369), .A(n10368), .B(n10367), .ZN(
        n10370) );
  INV_X1 U13347 ( .A(n10370), .ZN(n10371) );
  NAND3_X1 U13348 ( .A1(n10373), .A2(n10372), .A3(n10371), .ZN(n10382) );
  AND2_X2 U13349 ( .A1(n13133), .A2(n15811), .ZN(n10411) );
  AOI22_X1 U13350 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U13351 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__3__SCAN_IN), .B2(n10434), .ZN(n10379) );
  AND2_X2 U13352 ( .A1(n10376), .A2(n15811), .ZN(n10410) );
  AOI22_X1 U13353 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10410), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10378) );
  AND2_X2 U13354 ( .A1(n10235), .A2(n15811), .ZN(n10516) );
  AOI22_X1 U13355 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10516), .B1(
        n10445), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10377) );
  NAND4_X1 U13356 ( .A1(n10380), .A2(n10379), .A3(n10378), .A4(n10377), .ZN(
        n10381) );
  NAND2_X1 U13357 ( .A1(n10537), .A2(n10364), .ZN(n10384) );
  INV_X1 U13358 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10386) );
  INV_X1 U13359 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10421) );
  OAI22_X1 U13360 ( .A1(n10386), .A2(n10579), .B1(n19576), .B2(n10421), .ZN(
        n10387) );
  INV_X1 U13361 ( .A(n10387), .ZN(n10391) );
  NAND2_X1 U13362 ( .A1(n19269), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10390) );
  NAND3_X1 U13363 ( .A1(n10391), .A2(n10390), .A3(n10389), .ZN(n10395) );
  NAND2_X1 U13364 ( .A1(n10393), .A2(n10392), .ZN(n10394) );
  NOR2_X1 U13365 ( .A1(n10395), .A2(n10394), .ZN(n10405) );
  INV_X1 U13366 ( .A(n10482), .ZN(n10398) );
  INV_X1 U13367 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14302) );
  AOI21_X1 U13368 ( .B1(n10578), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n10383), .ZN(n10397) );
  NAND2_X1 U13369 ( .A1(n19541), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10396) );
  OAI211_X1 U13370 ( .C1(n10398), .C2(n14302), .A(n10397), .B(n10396), .ZN(
        n10399) );
  INV_X1 U13371 ( .A(n10399), .ZN(n10404) );
  AOI22_X1 U13372 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10481), .B1(
        n19396), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10403) );
  INV_X1 U13373 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10400) );
  INV_X1 U13374 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11117) );
  OAI22_X1 U13375 ( .A1(n10400), .A2(n19330), .B1(n10474), .B2(n11117), .ZN(
        n10401) );
  AOI21_X1 U13376 ( .B1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n19454), .A(
        n10401), .ZN(n10402) );
  NAND4_X1 U13377 ( .A1(n10405), .A2(n10404), .A3(n10403), .A4(n10402), .ZN(
        n10452) );
  AOI22_X1 U13378 ( .A1(n11178), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10409) );
  AOI22_X1 U13379 ( .A1(n10503), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12983), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10408) );
  AOI22_X1 U13380 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10407) );
  AOI22_X1 U13381 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10406) );
  NAND4_X1 U13382 ( .A1(n10409), .A2(n10408), .A3(n10407), .A4(n10406), .ZN(
        n10417) );
  AOI22_X1 U13383 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10415) );
  AOI22_X1 U13384 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10414) );
  AOI22_X1 U13385 ( .A1(n10410), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12982), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10413) );
  AOI22_X1 U13386 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10445), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10412) );
  NAND4_X1 U13387 ( .A1(n10415), .A2(n10414), .A3(n10413), .A4(n10412), .ZN(
        n10416) );
  NOR2_X1 U13388 ( .A1(n10417), .A2(n10416), .ZN(n10553) );
  INV_X1 U13389 ( .A(n10553), .ZN(n13305) );
  AOI22_X1 U13390 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10503), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10425) );
  NAND2_X1 U13391 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10420) );
  AOI22_X1 U13392 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n12982), .ZN(n10419) );
  OAI211_X1 U13393 ( .C1(n12987), .C2(n10421), .A(n10420), .B(n10419), .ZN(
        n10422) );
  INV_X1 U13394 ( .A(n10422), .ZN(n10424) );
  AOI22_X1 U13395 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n10434), .ZN(n10423) );
  NAND3_X1 U13396 ( .A1(n10425), .A2(n10424), .A3(n10423), .ZN(n10433) );
  AOI22_X1 U13397 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10431) );
  AOI22_X1 U13398 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10430) );
  AOI22_X1 U13399 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10410), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10429) );
  AOI22_X1 U13400 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10516), .B1(
        n10445), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10428) );
  NAND4_X1 U13401 ( .A1(n10431), .A2(n10430), .A3(n10429), .A4(n10428), .ZN(
        n10432) );
  NAND2_X1 U13402 ( .A1(n13305), .A2(n10731), .ZN(n10733) );
  AOI22_X1 U13403 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__2__SCAN_IN), .B2(n10434), .ZN(n10443) );
  INV_X1 U13404 ( .A(n10503), .ZN(n10438) );
  INV_X1 U13405 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10437) );
  NAND2_X1 U13406 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10436) );
  AOI22_X1 U13407 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__2__SCAN_IN), .B2(n12982), .ZN(n10435) );
  OAI211_X1 U13408 ( .C1(n10438), .C2(n10437), .A(n10436), .B(n10435), .ZN(
        n10439) );
  INV_X1 U13409 ( .A(n10439), .ZN(n10442) );
  AOI22_X1 U13410 ( .A1(n10491), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10441) );
  NAND3_X1 U13411 ( .A1(n10443), .A2(n10442), .A3(n10441), .ZN(n10451) );
  AOI22_X1 U13412 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10444), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10449) );
  AOI22_X1 U13413 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11178), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10448) );
  AOI22_X1 U13414 ( .A1(n10427), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10410), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10447) );
  AOI22_X1 U13415 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10516), .B1(
        n10445), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10446) );
  NAND4_X1 U13416 ( .A1(n10449), .A2(n10448), .A3(n10447), .A4(n10446), .ZN(
        n10450) );
  INV_X1 U13417 ( .A(n10734), .ZN(n11070) );
  OAI21_X1 U13418 ( .B1(n10733), .B2(n13297), .A(n11070), .ZN(n10737) );
  AND2_X2 U13419 ( .A1(n10452), .A2(n10737), .ZN(n10552) );
  AOI22_X1 U13420 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10491), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10459) );
  INV_X1 U13421 ( .A(n10426), .ZN(n10718) );
  INV_X1 U13422 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10455) );
  AOI22_X1 U13423 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__4__SCAN_IN), .B2(n12982), .ZN(n10454) );
  NAND2_X1 U13424 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10453) );
  OAI211_X1 U13425 ( .C1(n10718), .C2(n10455), .A(n10454), .B(n10453), .ZN(
        n10456) );
  INV_X1 U13426 ( .A(n10456), .ZN(n10458) );
  AOI22_X1 U13427 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_11__4__SCAN_IN), .B2(n10440), .ZN(n10457) );
  NAND3_X1 U13428 ( .A1(n10459), .A2(n10458), .A3(n10457), .ZN(n10466) );
  AOI22_X1 U13429 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11178), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10464) );
  AOI22_X1 U13430 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10503), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10463) );
  AOI22_X1 U13431 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10410), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10462) );
  AOI22_X1 U13432 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10516), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10461) );
  NAND4_X1 U13433 ( .A1(n10464), .A2(n10463), .A3(n10462), .A4(n10461), .ZN(
        n10465) );
  INV_X1 U13434 ( .A(n19576), .ZN(n10467) );
  AOI22_X1 U13435 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n10578), .B1(
        n10467), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10473) );
  AOI22_X1 U13436 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19300), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U13437 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19179), .B1(
        n10469), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10471) );
  AOI22_X1 U13438 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19239), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10470) );
  INV_X1 U13439 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10476) );
  INV_X1 U13440 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10475) );
  OAI22_X1 U13441 ( .A1(n10476), .A2(n10587), .B1(n10474), .B2(n10475), .ZN(
        n10480) );
  INV_X1 U13442 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10478) );
  INV_X1 U13443 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10477) );
  OAI22_X1 U13444 ( .A1(n10478), .A2(n19330), .B1(n19547), .B2(n10477), .ZN(
        n10479) );
  NOR2_X1 U13445 ( .A1(n10480), .A2(n10479), .ZN(n10485) );
  AOI22_X1 U13446 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n10481), .B1(
        n19454), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10484) );
  AOI22_X1 U13447 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n10482), .B1(
        n19396), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10483) );
  NAND4_X1 U13448 ( .A1(n10486), .A2(n10485), .A3(n10484), .A4(n10483), .ZN(
        n10502) );
  AOI22_X1 U13449 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10460), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10490) );
  AOI22_X1 U13450 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10503), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10489) );
  AOI22_X1 U13451 ( .A1(n10410), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13452 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10487) );
  NAND4_X1 U13453 ( .A1(n10490), .A2(n10489), .A3(n10488), .A4(n10487), .ZN(
        n10500) );
  AOI22_X1 U13454 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10498) );
  AOI22_X1 U13455 ( .A1(n11178), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10497) );
  INV_X1 U13456 ( .A(n12983), .ZN(n10493) );
  INV_X1 U13457 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14295) );
  NAND2_X1 U13458 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n12982), .ZN(
        n10492) );
  OAI21_X1 U13459 ( .B1(n10493), .B2(n14295), .A(n10492), .ZN(n10494) );
  AOI21_X1 U13460 ( .B1(n10434), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n10494), .ZN(n10496) );
  NAND2_X1 U13461 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10495) );
  NAND4_X1 U13462 ( .A1(n10498), .A2(n10497), .A3(n10496), .A4(n10495), .ZN(
        n10499) );
  NAND2_X1 U13463 ( .A1(n10546), .A2(n10383), .ZN(n10501) );
  NAND2_X1 U13464 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10507) );
  NAND2_X1 U13465 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10506) );
  NAND2_X1 U13466 ( .A1(n10503), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10505) );
  NAND2_X1 U13467 ( .A1(n10434), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10504) );
  NAND2_X1 U13468 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10511) );
  NAND2_X1 U13469 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10510) );
  NAND2_X1 U13470 ( .A1(n10491), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10509) );
  NAND2_X1 U13471 ( .A1(n10427), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10508) );
  INV_X1 U13472 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10514) );
  NAND2_X1 U13473 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10513) );
  AOI22_X1 U13474 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n12982), .ZN(n10512) );
  OAI211_X1 U13475 ( .C1(n12987), .C2(n10514), .A(n10513), .B(n10512), .ZN(
        n10515) );
  INV_X1 U13476 ( .A(n10515), .ZN(n10522) );
  NAND2_X1 U13477 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10520) );
  NAND2_X1 U13478 ( .A1(n10516), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10519) );
  NAND2_X1 U13479 ( .A1(n10410), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10518) );
  NAND2_X1 U13480 ( .A1(n10440), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10517) );
  NAND2_X1 U13481 ( .A1(n9589), .A2(n10628), .ZN(n10551) );
  NAND2_X1 U13482 ( .A1(n14135), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10525) );
  NAND2_X1 U13483 ( .A1(n16322), .A2(n19813), .ZN(n10530) );
  INV_X1 U13484 ( .A(n10723), .ZN(n10997) );
  MUX2_X1 U13485 ( .A(n11081), .B(n10997), .S(n13221), .Z(n10532) );
  INV_X1 U13486 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n13585) );
  MUX2_X1 U13487 ( .A(n10532), .B(n13585), .S(n11054), .Z(n10571) );
  MUX2_X1 U13488 ( .A(n19813), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        n16322), .Z(n10535) );
  INV_X1 U13489 ( .A(n10535), .ZN(n10534) );
  MUX2_X1 U13490 ( .A(n10535), .B(n10534), .S(n10533), .Z(n10708) );
  INV_X1 U13491 ( .A(n10708), .ZN(n10981) );
  MUX2_X1 U13492 ( .A(n10734), .B(n10981), .S(n13221), .Z(n10720) );
  INV_X1 U13493 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n14014) );
  MUX2_X1 U13494 ( .A(n10720), .B(n14014), .S(n11054), .Z(n10558) );
  NOR2_X1 U13495 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n10536) );
  MUX2_X1 U13496 ( .A(n10731), .B(n10536), .S(n11054), .Z(n10557) );
  NAND2_X1 U13497 ( .A1(n10558), .A2(n10557), .ZN(n10562) );
  INV_X1 U13498 ( .A(n10537), .ZN(n11076) );
  NOR2_X1 U13499 ( .A1(n10539), .A2(n10538), .ZN(n10540) );
  MUX2_X1 U13500 ( .A(n11076), .B(n10991), .S(n13221), .Z(n10542) );
  INV_X1 U13501 ( .A(n10542), .ZN(n10544) );
  NAND2_X1 U13502 ( .A1(n11054), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10543) );
  OAI21_X1 U13503 ( .B1(n10544), .B2(n11054), .A(n10543), .ZN(n10563) );
  MUX2_X1 U13504 ( .A(n10546), .B(P2_EBX_REG_5__SCAN_IN), .S(n11054), .Z(
        n10547) );
  INV_X1 U13505 ( .A(n10622), .ZN(n10550) );
  NAND2_X1 U13506 ( .A1(n10548), .A2(n10547), .ZN(n10549) );
  NAND2_X1 U13507 ( .A1(n10550), .A2(n10549), .ZN(n13999) );
  NAND2_X1 U13508 ( .A1(n10551), .A2(n13999), .ZN(n10573) );
  INV_X1 U13509 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14200) );
  XNOR2_X1 U13510 ( .A(n10573), .B(n14200), .ZN(n14189) );
  OAI21_X1 U13511 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19828), .A(
        n10711), .ZN(n10983) );
  MUX2_X1 U13512 ( .A(n10553), .B(n10983), .S(n13221), .Z(n10722) );
  INV_X1 U13513 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n10554) );
  MUX2_X1 U13514 ( .A(n10722), .B(n10554), .S(n11054), .Z(n18994) );
  INV_X1 U13515 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13304) );
  NOR2_X1 U13516 ( .A1(n18994), .A2(n13304), .ZN(n13345) );
  AND3_X1 U13517 ( .A1(n11054), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n10555) );
  NOR2_X1 U13518 ( .A1(n10557), .A2(n10555), .ZN(n14181) );
  NAND2_X1 U13519 ( .A1(n13345), .A2(n14181), .ZN(n10556) );
  NOR2_X1 U13520 ( .A1(n13345), .A2(n14181), .ZN(n13344) );
  AOI21_X1 U13521 ( .B1(n14051), .B2(n10556), .A(n13344), .ZN(n13394) );
  OAI21_X1 U13522 ( .B1(n10558), .B2(n10557), .A(n10562), .ZN(n14017) );
  XNOR2_X1 U13523 ( .A(n14017), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13393) );
  NAND2_X1 U13524 ( .A1(n13394), .A2(n13393), .ZN(n10561) );
  INV_X1 U13525 ( .A(n14017), .ZN(n10559) );
  NAND2_X1 U13526 ( .A1(n10559), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10560) );
  NAND2_X1 U13527 ( .A1(n10561), .A2(n10560), .ZN(n13812) );
  INV_X1 U13528 ( .A(n10562), .ZN(n10565) );
  INV_X1 U13529 ( .A(n10563), .ZN(n10564) );
  NOR2_X1 U13530 ( .A1(n10565), .A2(n10564), .ZN(n10566) );
  NOR2_X1 U13531 ( .A1(n10566), .A2(n10570), .ZN(n13988) );
  AOI21_X1 U13532 ( .B1(n13812), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n13988), .ZN(n10567) );
  NAND2_X1 U13533 ( .A1(n13811), .A2(n10567), .ZN(n10569) );
  OR2_X1 U13534 ( .A1(n13812), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10568) );
  XNOR2_X1 U13535 ( .A(n10571), .B(n10545), .ZN(n13910) );
  XNOR2_X1 U13536 ( .A(n13910), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14078) );
  INV_X1 U13537 ( .A(n13910), .ZN(n10572) );
  INV_X1 U13538 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14199) );
  NAND2_X1 U13539 ( .A1(n14189), .A2(n14190), .ZN(n10575) );
  NAND2_X1 U13540 ( .A1(n10573), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10574) );
  NAND2_X1 U13541 ( .A1(n10575), .A2(n10574), .ZN(n14314) );
  AOI22_X1 U13542 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10578), .B1(
        n10468), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10585) );
  AOI22_X1 U13543 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19179), .B1(
        n10388), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10584) );
  AOI22_X1 U13544 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19239), .B1(
        n10469), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10583) );
  INV_X1 U13545 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10580) );
  INV_X1 U13546 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10601) );
  OAI22_X1 U13547 ( .A1(n10580), .A2(n10579), .B1(n19576), .B2(n10601), .ZN(
        n10581) );
  INV_X1 U13548 ( .A(n10581), .ZN(n10582) );
  INV_X1 U13549 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10588) );
  INV_X1 U13550 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10586) );
  OAI22_X1 U13551 ( .A1(n10588), .A2(n19330), .B1(n10587), .B2(n10586), .ZN(
        n10591) );
  INV_X1 U13552 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10589) );
  INV_X1 U13553 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11196) );
  OAI22_X1 U13554 ( .A1(n10589), .A2(n19547), .B1(n10474), .B2(n11196), .ZN(
        n10590) );
  NOR2_X1 U13555 ( .A1(n10591), .A2(n10590), .ZN(n10594) );
  AOI22_X1 U13556 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19454), .B1(
        n19396), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U13557 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10481), .B1(
        n10482), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10592) );
  NAND4_X1 U13558 ( .A1(n10115), .A2(n10594), .A3(n10593), .A4(n10592), .ZN(
        n10609) );
  AOI22_X1 U13559 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10598) );
  AOI22_X1 U13560 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10597) );
  AOI22_X1 U13561 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10410), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10596) );
  AOI22_X1 U13562 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10516), .B1(
        n10445), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10595) );
  NAND4_X1 U13563 ( .A1(n10598), .A2(n10597), .A3(n10596), .A4(n10595), .ZN(
        n10607) );
  AOI22_X1 U13564 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10503), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10605) );
  NAND2_X1 U13565 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10600) );
  AOI22_X1 U13566 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__6__SCAN_IN), .B2(n12982), .ZN(n10599) );
  OAI211_X1 U13567 ( .C1(n12987), .C2(n10601), .A(n10600), .B(n10599), .ZN(
        n10602) );
  INV_X1 U13568 ( .A(n10602), .ZN(n10604) );
  AOI22_X1 U13569 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n10434), .ZN(n10603) );
  NAND3_X1 U13570 ( .A1(n10605), .A2(n10604), .A3(n10603), .ZN(n10606) );
  NAND2_X1 U13571 ( .A1(n11090), .A2(n10364), .ZN(n10608) );
  NAND2_X1 U13572 ( .A1(n10758), .A2(n10628), .ZN(n10610) );
  MUX2_X1 U13573 ( .A(n11090), .B(P2_EBX_REG_6__SCAN_IN), .S(n11054), .Z(
        n10614) );
  INV_X1 U13574 ( .A(n10614), .ZN(n10621) );
  XNOR2_X1 U13575 ( .A(n10622), .B(n10621), .ZN(n13895) );
  INV_X1 U13576 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11037) );
  XNOR2_X1 U13577 ( .A(n10611), .B(n11037), .ZN(n14315) );
  NAND2_X1 U13578 ( .A1(n14314), .A2(n14315), .ZN(n10613) );
  NAND2_X1 U13579 ( .A1(n10611), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10612) );
  MUX2_X1 U13580 ( .A(n10628), .B(P2_EBX_REG_7__SCAN_IN), .S(n11054), .Z(
        n10619) );
  NOR2_X1 U13581 ( .A1(n10614), .A2(n10619), .ZN(n10615) );
  NAND2_X1 U13582 ( .A1(n11054), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10616) );
  NOR2_X1 U13583 ( .A1(n10631), .A2(n10616), .ZN(n10617) );
  NOR2_X1 U13584 ( .A1(n10630), .A2(n10617), .ZN(n13874) );
  AND2_X1 U13585 ( .A1(n11094), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10618) );
  NAND2_X1 U13586 ( .A1(n13874), .A2(n10618), .ZN(n16235) );
  INV_X1 U13587 ( .A(n10619), .ZN(n10620) );
  AOI21_X1 U13588 ( .B1(n10622), .B2(n10621), .A(n10620), .ZN(n10623) );
  NOR2_X1 U13589 ( .A1(n10623), .A2(n10631), .ZN(n18976) );
  NAND2_X1 U13590 ( .A1(n18976), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16233) );
  NAND2_X1 U13591 ( .A1(n13874), .A2(n11094), .ZN(n10624) );
  INV_X1 U13592 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11038) );
  NAND2_X1 U13593 ( .A1(n10624), .A2(n11038), .ZN(n16236) );
  INV_X1 U13594 ( .A(n18976), .ZN(n10625) );
  INV_X1 U13595 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n14342) );
  NAND2_X1 U13596 ( .A1(n10625), .A2(n14342), .ZN(n16232) );
  AND2_X1 U13597 ( .A1(n16236), .A2(n16232), .ZN(n10626) );
  AND2_X1 U13598 ( .A1(n11054), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10627) );
  XNOR2_X1 U13599 ( .A(n10630), .B(n10627), .ZN(n18962) );
  NAND2_X1 U13600 ( .A1(n18962), .A2(n11094), .ZN(n10637) );
  INV_X1 U13601 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15788) );
  INV_X1 U13602 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10629) );
  NAND3_X1 U13603 ( .A1(n10633), .A2(n11054), .A3(P2_EBX_REG_10__SCAN_IN), 
        .ZN(n10632) );
  OAI211_X1 U13604 ( .C1(n10633), .C2(P2_EBX_REG_10__SCAN_IN), .A(n10890), .B(
        n10632), .ZN(n13884) );
  INV_X1 U13605 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15768) );
  OAI21_X1 U13606 ( .B1(n13884), .B2(n10628), .A(n15768), .ZN(n16213) );
  INV_X1 U13607 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13736) );
  AND2_X1 U13608 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n9655), .ZN(n10634) );
  NAND2_X1 U13609 ( .A1(n11054), .A2(n10634), .ZN(n13850) );
  NAND2_X1 U13610 ( .A1(n13850), .A2(n11094), .ZN(n10635) );
  OR2_X1 U13611 ( .A1(n13849), .A2(n10635), .ZN(n10639) );
  INV_X1 U13612 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15767) );
  NAND2_X1 U13613 ( .A1(n10639), .A2(n15767), .ZN(n15761) );
  NAND2_X1 U13614 ( .A1(n11094), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10636) );
  OR2_X1 U13615 ( .A1(n13884), .A2(n10636), .ZN(n16212) );
  INV_X1 U13616 ( .A(n10637), .ZN(n10638) );
  NAND2_X1 U13617 ( .A1(n10638), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16209) );
  NAND2_X1 U13618 ( .A1(n16212), .A2(n16209), .ZN(n15758) );
  NOR2_X1 U13619 ( .A1(n10639), .A2(n15767), .ZN(n15763) );
  NOR2_X1 U13620 ( .A1(n15758), .A2(n15763), .ZN(n10640) );
  NAND2_X1 U13621 ( .A1(n9685), .A2(n10642), .ZN(n10643) );
  NAND2_X1 U13622 ( .A1(n10647), .A2(n10643), .ZN(n13919) );
  INV_X1 U13623 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10644) );
  NOR2_X1 U13624 ( .A1(n10645), .A2(n10644), .ZN(n15743) );
  NAND2_X1 U13625 ( .A1(n10645), .A2(n10644), .ZN(n15742) );
  AND2_X1 U13626 ( .A1(n11054), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10646) );
  NAND2_X1 U13627 ( .A1(n10647), .A2(n10646), .ZN(n10648) );
  AND2_X1 U13628 ( .A1(n10662), .A2(n10648), .ZN(n14033) );
  NAND2_X1 U13629 ( .A1(n14033), .A2(n11094), .ZN(n10650) );
  INV_X1 U13630 ( .A(n10650), .ZN(n10649) );
  NAND2_X1 U13631 ( .A1(n10649), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16180) );
  INV_X1 U13632 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16276) );
  NAND2_X1 U13633 ( .A1(n10650), .A2(n16276), .ZN(n16179) );
  INV_X1 U13634 ( .A(n16179), .ZN(n10651) );
  NAND2_X1 U13635 ( .A1(n10662), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10652) );
  MUX2_X1 U13636 ( .A(n10652), .B(n10662), .S(n10038), .Z(n10653) );
  INV_X1 U13637 ( .A(n10653), .ZN(n10656) );
  INV_X1 U13638 ( .A(n10662), .ZN(n10654) );
  INV_X1 U13639 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n10659) );
  NAND2_X1 U13640 ( .A1(n10654), .A2(n10659), .ZN(n10663) );
  INV_X1 U13641 ( .A(n10663), .ZN(n10655) );
  NOR2_X1 U13642 ( .A1(n10656), .A2(n10655), .ZN(n18947) );
  NAND2_X1 U13643 ( .A1(n18947), .A2(n11094), .ZN(n10669) );
  INV_X1 U13644 ( .A(n10669), .ZN(n10657) );
  NAND2_X1 U13645 ( .A1(n10657), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15727) );
  INV_X1 U13646 ( .A(n15727), .ZN(n10658) );
  INV_X1 U13647 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n14249) );
  NAND2_X1 U13648 ( .A1(n10659), .A2(n14249), .ZN(n10660) );
  AND2_X1 U13649 ( .A1(n11054), .A2(n10660), .ZN(n10661) );
  INV_X1 U13650 ( .A(n10672), .ZN(n10665) );
  NAND3_X1 U13651 ( .A1(n10663), .A2(P2_EBX_REG_15__SCAN_IN), .A3(n11054), 
        .ZN(n10664) );
  NAND2_X1 U13652 ( .A1(n10665), .A2(n10664), .ZN(n14253) );
  NAND2_X1 U13653 ( .A1(n11094), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10666) );
  OR2_X1 U13654 ( .A1(n14253), .A2(n10628), .ZN(n10668) );
  INV_X1 U13655 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10667) );
  NAND2_X1 U13656 ( .A1(n10668), .A2(n10667), .ZN(n15561) );
  AND2_X1 U13657 ( .A1(n15561), .A2(n16179), .ZN(n10670) );
  INV_X1 U13658 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15736) );
  NAND2_X1 U13659 ( .A1(n10669), .A2(n15736), .ZN(n15728) );
  AND2_X1 U13660 ( .A1(n10670), .A2(n15728), .ZN(n10857) );
  NAND2_X1 U13661 ( .A1(n11054), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10671) );
  INV_X1 U13662 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n14074) );
  OAI211_X1 U13663 ( .C1(n10672), .C2(n10671), .A(n10890), .B(n10675), .ZN(
        n18937) );
  OR2_X1 U13664 ( .A1(n18937), .A2(n10628), .ZN(n10673) );
  XNOR2_X1 U13665 ( .A(n10673), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15549) );
  NAND2_X1 U13666 ( .A1(n11094), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10674) );
  OR2_X1 U13667 ( .A1(n18937), .A2(n10674), .ZN(n10861) );
  NAND2_X1 U13668 ( .A1(n15548), .A2(n10861), .ZN(n15539) );
  NAND2_X2 U13669 ( .A1(n10675), .A2(n10890), .ZN(n10677) );
  NAND2_X1 U13670 ( .A1(n11054), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10676) );
  OR2_X1 U13671 ( .A1(n10677), .A2(n10676), .ZN(n10678) );
  AND2_X1 U13672 ( .A1(n10688), .A2(n10678), .ZN(n10680) );
  NAND2_X1 U13673 ( .A1(n10680), .A2(n11094), .ZN(n10679) );
  INV_X1 U13674 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15702) );
  NAND2_X1 U13675 ( .A1(n10679), .A2(n15702), .ZN(n10856) );
  INV_X1 U13676 ( .A(n10680), .ZN(n18925) );
  NAND2_X1 U13677 ( .A1(n11094), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10681) );
  OR2_X1 U13678 ( .A1(n18925), .A2(n10681), .ZN(n10862) );
  NAND2_X1 U13679 ( .A1(n10856), .A2(n10862), .ZN(n15540) );
  NAND2_X1 U13680 ( .A1(n10688), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10682) );
  MUX2_X1 U13681 ( .A(n10688), .B(n10682), .S(n11054), .Z(n10683) );
  OR2_X1 U13682 ( .A1(n10688), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10685) );
  INV_X1 U13683 ( .A(n10691), .ZN(n18914) );
  NAND2_X1 U13684 ( .A1(n11094), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10684) );
  NAND3_X1 U13685 ( .A1(n10685), .A2(P2_EBX_REG_19__SCAN_IN), .A3(n11054), 
        .ZN(n10689) );
  INV_X1 U13686 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n15348) );
  INV_X1 U13687 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n14178) );
  NAND2_X1 U13688 ( .A1(n15348), .A2(n14178), .ZN(n10686) );
  AND2_X1 U13689 ( .A1(n11054), .A2(n10686), .ZN(n10687) );
  NAND2_X1 U13690 ( .A1(n10689), .A2(n10696), .ZN(n15263) );
  INV_X1 U13691 ( .A(n10694), .ZN(n10690) );
  NAND2_X1 U13692 ( .A1(n10690), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15517) );
  NAND2_X1 U13693 ( .A1(n10691), .A2(n11094), .ZN(n10692) );
  INV_X1 U13694 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15688) );
  NAND2_X1 U13695 ( .A1(n10692), .A2(n15688), .ZN(n15528) );
  INV_X1 U13696 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10693) );
  NAND2_X1 U13697 ( .A1(n10694), .A2(n10693), .ZN(n15516) );
  AND2_X1 U13698 ( .A1(n15528), .A2(n15516), .ZN(n10859) );
  INV_X1 U13699 ( .A(n10702), .ZN(n10698) );
  NAND2_X1 U13700 ( .A1(n10696), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10695) );
  MUX2_X1 U13701 ( .A(n10696), .B(n10695), .S(n11054), .Z(n10697) );
  NAND2_X1 U13702 ( .A1(n18904), .A2(n11094), .ZN(n10699) );
  INV_X1 U13703 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15508) );
  NAND2_X1 U13704 ( .A1(n10699), .A2(n15508), .ZN(n15502) );
  INV_X1 U13705 ( .A(n10699), .ZN(n10700) );
  NAND2_X1 U13706 ( .A1(n10700), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15503) );
  INV_X1 U13707 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n15333) );
  NAND2_X1 U13708 ( .A1(n10871), .A2(n10890), .ZN(n10868) );
  NAND2_X1 U13709 ( .A1(n11054), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10701) );
  NOR2_X1 U13710 ( .A1(n10702), .A2(n10701), .ZN(n10703) );
  OR2_X1 U13711 ( .A1(n10868), .A2(n10703), .ZN(n18889) );
  OR2_X1 U13712 ( .A1(n18889), .A2(n10628), .ZN(n10704) );
  INV_X1 U13713 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11269) );
  NAND2_X1 U13714 ( .A1(n10704), .A2(n11269), .ZN(n10860) );
  NAND2_X1 U13715 ( .A1(n11094), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10705) );
  OR2_X1 U13716 ( .A1(n18889), .A2(n10705), .ZN(n10864) );
  NAND2_X1 U13717 ( .A1(n10860), .A2(n10864), .ZN(n10706) );
  XNOR2_X1 U13718 ( .A(n10707), .B(n10706), .ZN(n15650) );
  NOR3_X1 U13719 ( .A1(n10991), .A2(n10723), .A3(n10708), .ZN(n10713) );
  INV_X1 U13720 ( .A(n10713), .ZN(n10716) );
  NOR2_X1 U13721 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16330), .ZN(
        n10709) );
  INV_X1 U13722 ( .A(n10711), .ZN(n10712) );
  XNOR2_X1 U13723 ( .A(n10982), .B(n10712), .ZN(n10984) );
  AND2_X1 U13724 ( .A1(n10984), .A2(n10713), .ZN(n10714) );
  OR2_X1 U13725 ( .A1(n10999), .A2(n10714), .ZN(n16337) );
  INV_X1 U13726 ( .A(n16337), .ZN(n10715) );
  OAI21_X1 U13727 ( .B1(n10983), .B2(n10716), .A(n10715), .ZN(n10719) );
  AND2_X1 U13728 ( .A1(n15860), .A2(n10717), .ZN(n16343) );
  AOI21_X1 U13729 ( .B1(n10718), .B2(n16343), .A(P2_FLUSH_REG_SCAN_IN), .ZN(
        n16368) );
  MUX2_X1 U13730 ( .A(n10719), .B(n16368), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n19834) );
  INV_X1 U13731 ( .A(n10999), .ZN(n10726) );
  INV_X1 U13732 ( .A(n10720), .ZN(n10721) );
  OAI21_X1 U13733 ( .B1(n10722), .B2(n10982), .A(n10721), .ZN(n10724) );
  NOR2_X1 U13734 ( .A1(n10723), .A2(n10991), .ZN(n10995) );
  NAND2_X1 U13735 ( .A1(n10724), .A2(n10995), .ZN(n10725) );
  NAND2_X1 U13736 ( .A1(n10726), .A2(n10725), .ZN(n19832) );
  INV_X1 U13737 ( .A(n19831), .ZN(n19844) );
  OAI22_X1 U13738 ( .A1(n19834), .A2(n10364), .B1(n19832), .B2(n19844), .ZN(
        n10728) );
  NOR2_X1 U13739 ( .A1(n19846), .A2(n18863), .ZN(n10729) );
  NAND2_X1 U13740 ( .A1(n15650), .A2(n19121), .ZN(n10852) );
  INV_X1 U13741 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11034) );
  NOR2_X1 U13742 ( .A1(n13305), .A2(n13304), .ZN(n13303) );
  INV_X1 U13743 ( .A(n10731), .ZN(n11063) );
  NAND2_X1 U13744 ( .A1(n13303), .A2(n10731), .ZN(n10732) );
  NOR2_X1 U13745 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13305), .ZN(
        n10730) );
  XNOR2_X1 U13746 ( .A(n10731), .B(n10730), .ZN(n13348) );
  NAND2_X1 U13747 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13348), .ZN(
        n13347) );
  NAND2_X1 U13748 ( .A1(n10732), .A2(n13347), .ZN(n10738) );
  XNOR2_X1 U13749 ( .A(n11034), .B(n10738), .ZN(n13396) );
  INV_X1 U13750 ( .A(n10733), .ZN(n10735) );
  NAND2_X1 U13751 ( .A1(n10735), .A2(n10734), .ZN(n10736) );
  NAND2_X1 U13752 ( .A1(n10737), .A2(n10736), .ZN(n13395) );
  NAND2_X1 U13753 ( .A1(n13396), .A2(n13395), .ZN(n10740) );
  NAND2_X1 U13754 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10738), .ZN(
        n10739) );
  NAND2_X1 U13755 ( .A1(n10740), .A2(n10739), .ZN(n10741) );
  XNOR2_X1 U13756 ( .A(n10741), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13815) );
  NAND2_X1 U13757 ( .A1(n10741), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10742) );
  OAI21_X2 U13758 ( .B1(n13816), .B2(n13815), .A(n10742), .ZN(n10746) );
  INV_X1 U13759 ( .A(n11081), .ZN(n10743) );
  XNOR2_X1 U13760 ( .A(n10744), .B(n10743), .ZN(n10747) );
  INV_X1 U13761 ( .A(n10747), .ZN(n10745) );
  NAND2_X1 U13762 ( .A1(n10746), .A2(n10745), .ZN(n14075) );
  NAND2_X1 U13763 ( .A1(n14075), .A2(n14199), .ZN(n10749) );
  INV_X1 U13764 ( .A(n10746), .ZN(n10748) );
  NAND2_X1 U13765 ( .A1(n10748), .A2(n10747), .ZN(n14076) );
  AND2_X2 U13766 ( .A1(n10749), .A2(n14076), .ZN(n14194) );
  NAND2_X1 U13767 ( .A1(n10752), .A2(n14200), .ZN(n14191) );
  NAND2_X2 U13768 ( .A1(n14194), .A2(n14191), .ZN(n14196) );
  NAND2_X1 U13769 ( .A1(n10751), .A2(n10750), .ZN(n10757) );
  NAND2_X1 U13770 ( .A1(n14196), .A2(n9647), .ZN(n10756) );
  INV_X1 U13771 ( .A(n14192), .ZN(n14195) );
  INV_X1 U13772 ( .A(n10753), .ZN(n10754) );
  NAND2_X1 U13773 ( .A1(n14195), .A2(n10754), .ZN(n10755) );
  NAND2_X1 U13774 ( .A1(n14196), .A2(n14192), .ZN(n10759) );
  NAND2_X1 U13775 ( .A1(n10759), .A2(n10758), .ZN(n10763) );
  NAND2_X1 U13776 ( .A1(n10760), .A2(n10628), .ZN(n10761) );
  NAND2_X1 U13777 ( .A1(n10766), .A2(n10761), .ZN(n14343) );
  INV_X1 U13778 ( .A(n14343), .ZN(n10762) );
  XNOR2_X1 U13779 ( .A(n10766), .B(n11038), .ZN(n16229) );
  NAND2_X1 U13780 ( .A1(n10765), .A2(n10764), .ZN(n16231) );
  INV_X1 U13781 ( .A(n10766), .ZN(n10767) );
  NAND2_X1 U13782 ( .A1(n10767), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10768) );
  AND3_X1 U13783 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15734) );
  AND2_X1 U13784 ( .A1(n15734), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15731) );
  NAND2_X1 U13785 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15698) );
  AND2_X1 U13786 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11267) );
  INV_X1 U13787 ( .A(n11267), .ZN(n11042) );
  NOR2_X1 U13788 ( .A1(n11042), .A2(n15688), .ZN(n10771) );
  OAI21_X1 U13789 ( .B1(n10773), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n10853), .ZN(n15660) );
  INV_X1 U13790 ( .A(n18865), .ZN(n10774) );
  NOR2_X2 U13791 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19793) );
  NAND2_X1 U13792 ( .A1(n10302), .A2(n19839), .ZN(n15857) );
  INV_X1 U13793 ( .A(n15857), .ZN(n19792) );
  OR2_X1 U13794 ( .A1(n19793), .A2(n19792), .ZN(n19824) );
  NAND2_X1 U13795 ( .A1(n19824), .A2(n13325), .ZN(n10775) );
  NAND2_X1 U13796 ( .A1(n13325), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12869) );
  NAND2_X1 U13797 ( .A1(n19791), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10776) );
  NAND2_X1 U13798 ( .A1(n12869), .A2(n10776), .ZN(n13308) );
  NAND2_X1 U13799 ( .A1(n13201), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13198) );
  INV_X1 U13800 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n14244) );
  INV_X1 U13801 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10841) );
  AOI21_X1 U13802 ( .B1(n10777), .B2(n10841), .A(n9694), .ZN(n18887) );
  NOR2_X1 U13803 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n15857), .ZN(n13267) );
  NAND2_X1 U13804 ( .A1(n13267), .A2(n13325), .ZN(n11257) );
  OR2_X1 U13805 ( .A1(n15534), .A2(n19763), .ZN(n15653) );
  OAI21_X1 U13806 ( .B1(n16265), .B2(n10841), .A(n15653), .ZN(n10848) );
  INV_X1 U13807 ( .A(n10778), .ZN(n10780) );
  NAND2_X1 U13808 ( .A1(n10780), .A2(n10779), .ZN(n10783) );
  NAND2_X1 U13809 ( .A1(n10784), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10788) );
  INV_X1 U13810 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11084) );
  INV_X1 U13811 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10785) );
  OAI22_X1 U13812 ( .A1(n10936), .A2(n11084), .B1(n10302), .B2(n10785), .ZN(
        n10786) );
  AOI21_X1 U13813 ( .B1(n10926), .B2(P2_EBX_REG_4__SCAN_IN), .A(n10786), .ZN(
        n10787) );
  NAND2_X1 U13814 ( .A1(n10788), .A2(n10787), .ZN(n13582) );
  NAND2_X1 U13815 ( .A1(n10784), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10791) );
  INV_X1 U13816 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n11089) );
  OAI22_X1 U13817 ( .A1(n10936), .A2(n11089), .B1(n10302), .B2(n16264), .ZN(
        n10789) );
  AOI21_X1 U13818 ( .B1(n10926), .B2(P2_EBX_REG_5__SCAN_IN), .A(n10789), .ZN(
        n10790) );
  NAND2_X1 U13819 ( .A1(n10791), .A2(n10790), .ZN(n13613) );
  NAND2_X1 U13820 ( .A1(n10784), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10795) );
  INV_X1 U13821 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n14317) );
  INV_X1 U13822 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10792) );
  OAI22_X1 U13823 ( .A1(n10936), .A2(n14317), .B1(n10302), .B2(n10792), .ZN(
        n10793) );
  AOI21_X1 U13824 ( .B1(n9599), .B2(P2_EBX_REG_6__SCAN_IN), .A(n10793), .ZN(
        n10794) );
  NAND2_X1 U13825 ( .A1(n10784), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10800) );
  INV_X1 U13826 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n10797) );
  OAI22_X1 U13827 ( .A1(n10936), .A2(n10797), .B1(n10302), .B2(n18973), .ZN(
        n10798) );
  AOI21_X1 U13828 ( .B1(n9599), .B2(P2_EBX_REG_7__SCAN_IN), .A(n10798), .ZN(
        n10799) );
  NAND2_X1 U13829 ( .A1(n10784), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10805) );
  INV_X1 U13830 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n11113) );
  INV_X1 U13831 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10802) );
  OAI22_X1 U13832 ( .A1(n10936), .A2(n11113), .B1(n10302), .B2(n10802), .ZN(
        n10803) );
  AOI21_X1 U13833 ( .B1(n9599), .B2(P2_EBX_REG_8__SCAN_IN), .A(n10803), .ZN(
        n10804) );
  NAND2_X1 U13834 ( .A1(n10784), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10808) );
  INV_X1 U13835 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n11130) );
  OAI22_X1 U13836 ( .A1(n10936), .A2(n11130), .B1(n10302), .B2(n16227), .ZN(
        n10806) );
  AOI21_X1 U13837 ( .B1(n9599), .B2(P2_EBX_REG_9__SCAN_IN), .A(n10806), .ZN(
        n10807) );
  NAND2_X1 U13838 ( .A1(n10808), .A2(n10807), .ZN(n13727) );
  NAND2_X1 U13839 ( .A1(n10784), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10811) );
  INV_X1 U13840 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n11146) );
  OAI22_X1 U13841 ( .A1(n10936), .A2(n11146), .B1(n10302), .B2(n9933), .ZN(
        n10809) );
  AOI21_X1 U13842 ( .B1(n10926), .B2(P2_EBX_REG_10__SCAN_IN), .A(n10809), .ZN(
        n10810) );
  NAND2_X1 U13843 ( .A1(n10784), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10815) );
  INV_X1 U13844 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n10812) );
  OAI22_X1 U13845 ( .A1(n10936), .A2(n10812), .B1(n10302), .B2(n16206), .ZN(
        n10813) );
  AOI21_X1 U13846 ( .B1(n9599), .B2(P2_EBX_REG_11__SCAN_IN), .A(n10813), .ZN(
        n10814) );
  NAND2_X1 U13847 ( .A1(n10784), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10818) );
  INV_X1 U13848 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n11176) );
  OAI22_X1 U13849 ( .A1(n10936), .A2(n11176), .B1(n10302), .B2(n13917), .ZN(
        n10816) );
  AOI21_X1 U13850 ( .B1(n9599), .B2(P2_EBX_REG_12__SCAN_IN), .A(n10816), .ZN(
        n10817) );
  NAND2_X1 U13851 ( .A1(n10818), .A2(n10817), .ZN(n13604) );
  NAND2_X1 U13852 ( .A1(n13735), .A2(n13604), .ZN(n13605) );
  NAND2_X1 U13853 ( .A1(n10784), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10821) );
  INV_X1 U13854 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n14042) );
  OAI22_X1 U13855 ( .A1(n10936), .A2(n14042), .B1(n10302), .B2(n16189), .ZN(
        n10819) );
  AOI21_X1 U13856 ( .B1(n10926), .B2(P2_EBX_REG_13__SCAN_IN), .A(n10819), .ZN(
        n10820) );
  NAND2_X1 U13857 ( .A1(n10784), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10825) );
  INV_X1 U13858 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n11209) );
  INV_X1 U13859 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10822) );
  OAI22_X1 U13860 ( .A1(n10936), .A2(n11209), .B1(n10302), .B2(n10822), .ZN(
        n10823) );
  AOI21_X1 U13861 ( .B1(n9599), .B2(P2_EBX_REG_14__SCAN_IN), .A(n10823), .ZN(
        n10824) );
  NAND2_X1 U13862 ( .A1(n10825), .A2(n10824), .ZN(n13838) );
  AOI22_X1 U13863 ( .A1(n10940), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n10826) );
  OAI21_X1 U13864 ( .B1(n10934), .B2(n14249), .A(n10826), .ZN(n10827) );
  AOI21_X1 U13865 ( .B1(n10784), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n10827), .ZN(n13959) );
  AOI22_X1 U13866 ( .A1(n10940), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n10828) );
  OAI21_X1 U13867 ( .B1(n10934), .B2(n14074), .A(n10828), .ZN(n10829) );
  AOI21_X1 U13868 ( .B1(n10784), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n10829), .ZN(n14070) );
  INV_X1 U13869 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n10831) );
  AOI22_X1 U13870 ( .A1(n10940), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n10830) );
  OAI21_X1 U13871 ( .B1(n10934), .B2(n10831), .A(n10830), .ZN(n10832) );
  AOI21_X1 U13872 ( .B1(n10784), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10832), .ZN(n14137) );
  NAND2_X1 U13873 ( .A1(n10784), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10836) );
  INV_X1 U13874 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15533) );
  INV_X1 U13875 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10833) );
  OAI22_X1 U13876 ( .A1(n10936), .A2(n15533), .B1(n10302), .B2(n10833), .ZN(
        n10834) );
  AOI21_X1 U13877 ( .B1(n10926), .B2(P2_EBX_REG_18__SCAN_IN), .A(n10834), .ZN(
        n10835) );
  NAND2_X1 U13878 ( .A1(n10836), .A2(n10835), .ZN(n14173) );
  AOI22_X1 U13879 ( .A1(n10940), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n10837) );
  OAI21_X1 U13880 ( .B1(n10934), .B2(n15348), .A(n10837), .ZN(n10838) );
  AOI21_X1 U13881 ( .B1(n10784), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n10838), .ZN(n15266) );
  AOI22_X1 U13882 ( .A1(n10940), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n10839) );
  OAI21_X1 U13883 ( .B1(n10934), .B2(n9898), .A(n10839), .ZN(n10840) );
  AOI21_X1 U13884 ( .B1(n10784), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n10840), .ZN(n15335) );
  NAND2_X1 U13885 ( .A1(n10784), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10844) );
  OAI22_X1 U13886 ( .A1(n10936), .A2(n19763), .B1(n10302), .B2(n10841), .ZN(
        n10842) );
  AOI21_X1 U13887 ( .B1(n9599), .B2(P2_EBX_REG_21__SCAN_IN), .A(n10842), .ZN(
        n10843) );
  NAND2_X1 U13888 ( .A1(n10844), .A2(n10843), .ZN(n10845) );
  NOR2_X1 U13889 ( .A1(n15337), .A2(n10845), .ZN(n10846) );
  OR2_X1 U13890 ( .A1(n15328), .A2(n10846), .ZN(n18892) );
  AND2_X1 U13891 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19814) );
  NOR2_X1 U13892 ( .A1(n18892), .A2(n16247), .ZN(n10847) );
  AOI211_X1 U13893 ( .C1(n16255), .C2(n18887), .A(n10848), .B(n10847), .ZN(
        n10849) );
  NAND2_X1 U13894 ( .A1(n10852), .A2(n10851), .ZN(P2_U2993) );
  INV_X1 U13895 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15640) );
  INV_X1 U13896 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10876) );
  INV_X1 U13897 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15464) );
  INV_X1 U13898 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11289) );
  INV_X1 U13899 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15582) );
  INV_X1 U13900 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10855) );
  NAND2_X1 U13901 ( .A1(n11301), .A2(n19118), .ZN(n10951) );
  AND3_X1 U13902 ( .A1(n10857), .A2(n10856), .A3(n15549), .ZN(n10858) );
  NAND4_X1 U13903 ( .A1(n10860), .A2(n10859), .A3(n10858), .A4(n15502), .ZN(
        n10867) );
  AND3_X1 U13904 ( .A1(n10861), .A2(n15560), .A3(n16180), .ZN(n10863) );
  AND4_X1 U13905 ( .A1(n15517), .A2(n10863), .A3(n15727), .A4(n10862), .ZN(
        n10865) );
  AND4_X1 U13906 ( .A1(n15503), .A2(n10865), .A3(n15527), .A4(n10864), .ZN(
        n10866) );
  NAND2_X1 U13907 ( .A1(n11054), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10869) );
  NAND2_X1 U13908 ( .A1(n10868), .A2(n10869), .ZN(n10880) );
  INV_X1 U13909 ( .A(n10869), .ZN(n10870) );
  NAND2_X1 U13910 ( .A1(n10871), .A2(n10870), .ZN(n10872) );
  NAND2_X1 U13911 ( .A1(n10880), .A2(n10872), .ZN(n15891) );
  NAND2_X1 U13912 ( .A1(n10873), .A2(n15640), .ZN(n15493) );
  AND2_X1 U13913 ( .A1(n11054), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10879) );
  INV_X1 U13914 ( .A(n10879), .ZN(n10875) );
  XNOR2_X1 U13915 ( .A(n10880), .B(n10875), .ZN(n15258) );
  NAND2_X1 U13916 ( .A1(n15258), .A2(n11094), .ZN(n10877) );
  XNOR2_X1 U13917 ( .A(n10877), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15488) );
  OR2_X1 U13918 ( .A1(n10877), .A2(n10876), .ZN(n10878) );
  NAND3_X1 U13919 ( .A1(n9634), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n11054), .ZN(
        n10881) );
  NAND2_X1 U13920 ( .A1(n10881), .A2(n10890), .ZN(n10882) );
  OR2_X1 U13921 ( .A1(n10885), .A2(n10882), .ZN(n16155) );
  INV_X1 U13922 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15619) );
  NOR2_X1 U13923 ( .A1(n10884), .A2(n15619), .ZN(n15475) );
  NAND2_X1 U13924 ( .A1(n10884), .A2(n15619), .ZN(n15476) );
  INV_X1 U13925 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15301) );
  NOR2_X1 U13926 ( .A1(n10885), .A2(n15301), .ZN(n10886) );
  NAND2_X1 U13927 ( .A1(n11054), .A2(n10886), .ZN(n10887) );
  AND2_X1 U13928 ( .A1(n10890), .A2(n10887), .ZN(n10888) );
  NAND2_X1 U13929 ( .A1(n9646), .A2(n10888), .ZN(n15243) );
  OR2_X1 U13930 ( .A1(n15243), .A2(n10628), .ZN(n10889) );
  NAND2_X1 U13931 ( .A1(n10889), .A2(n15464), .ZN(n15460) );
  INV_X1 U13932 ( .A(n10890), .ZN(n10891) );
  OR2_X1 U13933 ( .A1(n15224), .A2(n10628), .ZN(n10894) );
  XNOR2_X1 U13934 ( .A(n10894), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15455) );
  NAND2_X1 U13935 ( .A1(n11054), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15202) );
  NAND2_X1 U13936 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15583) );
  INV_X1 U13937 ( .A(n15583), .ZN(n10897) );
  AND2_X1 U13938 ( .A1(n11054), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10893) );
  AOI21_X1 U13939 ( .B1(n10893), .B2(n15204), .A(n10901), .ZN(n15193) );
  NAND2_X1 U13940 ( .A1(n11275), .A2(n11289), .ZN(n11043) );
  INV_X1 U13941 ( .A(n10894), .ZN(n10895) );
  NAND2_X1 U13942 ( .A1(n10895), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10896) );
  NAND2_X1 U13943 ( .A1(n15459), .A2(n10896), .ZN(n10956) );
  NAND2_X1 U13944 ( .A1(n10952), .A2(n10898), .ZN(n15428) );
  NAND2_X1 U13945 ( .A1(n11054), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10900) );
  XOR2_X1 U13946 ( .A(n10900), .B(n10901), .Z(n15186) );
  INV_X1 U13947 ( .A(n15186), .ZN(n10899) );
  OAI21_X1 U13948 ( .B1(n10899), .B2(n10628), .A(n15582), .ZN(n15430) );
  NAND2_X1 U13949 ( .A1(n15428), .A2(n15430), .ZN(n14542) );
  NAND2_X1 U13950 ( .A1(n10901), .A2(n10900), .ZN(n10906) );
  NAND2_X1 U13951 ( .A1(n11054), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10902) );
  AOI21_X1 U13952 ( .B1(n13237), .B2(n11094), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14543) );
  INV_X1 U13953 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11311) );
  OR3_X1 U13954 ( .A1(n10142), .A2(n10628), .A3(n11311), .ZN(n14544) );
  NAND3_X1 U13955 ( .A1(n15186), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11094), .ZN(n15429) );
  INV_X1 U13956 ( .A(n15429), .ZN(n10903) );
  NOR2_X1 U13957 ( .A1(n10904), .A2(n10903), .ZN(n10905) );
  INV_X1 U13958 ( .A(n15224), .ZN(n10908) );
  NOR2_X1 U13959 ( .A1(n10906), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10907) );
  MUX2_X1 U13960 ( .A(n10908), .B(n10907), .S(n11054), .Z(n15171) );
  NAND2_X1 U13961 ( .A1(n15171), .A2(n11094), .ZN(n10909) );
  XOR2_X1 U13962 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n10909), .Z(
        n10910) );
  XNOR2_X1 U13963 ( .A(n10911), .B(n10910), .ZN(n11319) );
  NAND2_X1 U13964 ( .A1(n11319), .A2(n19121), .ZN(n10950) );
  NAND2_X1 U13965 ( .A1(n10784), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10914) );
  INV_X1 U13966 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19765) );
  OAI22_X1 U13967 ( .A1(n10936), .A2(n19765), .B1(n10302), .B2(n9937), .ZN(
        n10912) );
  AOI21_X1 U13968 ( .B1(n9599), .B2(P2_EBX_REG_22__SCAN_IN), .A(n10912), .ZN(
        n10913) );
  NAND2_X1 U13969 ( .A1(n10914), .A2(n10913), .ZN(n15327) );
  NAND2_X1 U13970 ( .A1(n15328), .A2(n15327), .ZN(n15244) );
  INV_X1 U13971 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10916) );
  AOI22_X1 U13972 ( .A1(n10940), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n10915) );
  OAI21_X1 U13973 ( .B1(n10934), .B2(n10916), .A(n10915), .ZN(n10917) );
  AOI21_X1 U13974 ( .B1(n10784), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n10917), .ZN(n15245) );
  INV_X1 U13975 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n15315) );
  AOI22_X1 U13976 ( .A1(n10940), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n10918) );
  OAI21_X1 U13977 ( .B1(n10934), .B2(n15315), .A(n10918), .ZN(n10919) );
  AOI21_X1 U13978 ( .B1(n10784), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n10919), .ZN(n15309) );
  AOI22_X1 U13979 ( .A1(n10940), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n10920) );
  OAI21_X1 U13980 ( .B1(n10934), .B2(n15301), .A(n10920), .ZN(n10921) );
  AOI21_X1 U13981 ( .B1(n10784), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n10921), .ZN(n15231) );
  NAND2_X1 U13982 ( .A1(n10784), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10924) );
  INV_X1 U13983 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n15223) );
  INV_X1 U13984 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15449) );
  OAI22_X1 U13985 ( .A1(n10936), .A2(n15223), .B1(n10302), .B2(n15449), .ZN(
        n10922) );
  AOI21_X1 U13986 ( .B1(n9599), .B2(P2_EBX_REG_26__SCAN_IN), .A(n10922), .ZN(
        n10923) );
  NAND2_X1 U13987 ( .A1(n10924), .A2(n10923), .ZN(n15213) );
  NAND2_X1 U13988 ( .A1(n10784), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10928) );
  INV_X1 U13989 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19775) );
  INV_X1 U13990 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15439) );
  OAI22_X1 U13991 ( .A1(n10936), .A2(n19775), .B1(n10302), .B2(n15439), .ZN(
        n10925) );
  AOI21_X1 U13992 ( .B1(n9599), .B2(P2_EBX_REG_27__SCAN_IN), .A(n10925), .ZN(
        n10927) );
  NAND2_X1 U13993 ( .A1(n10928), .A2(n10927), .ZN(n11287) );
  NAND2_X1 U13994 ( .A1(n10784), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10931) );
  INV_X1 U13995 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19776) );
  OAI22_X1 U13996 ( .A1(n10936), .A2(n19776), .B1(n10302), .B2(n9928), .ZN(
        n10929) );
  AOI21_X1 U13997 ( .B1(n10926), .B2(P2_EBX_REG_28__SCAN_IN), .A(n10929), .ZN(
        n10930) );
  NAND2_X1 U13998 ( .A1(n10931), .A2(n10930), .ZN(n11046) );
  INV_X1 U13999 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n10933) );
  AOI22_X1 U14000 ( .A1(n10940), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n10932) );
  OAI21_X1 U14001 ( .B1(n10934), .B2(n10933), .A(n10932), .ZN(n10935) );
  AOI21_X1 U14002 ( .B1(n10784), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n10935), .ZN(n15174) );
  NAND2_X1 U14003 ( .A1(n10784), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10939) );
  INV_X1 U14004 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n14551) );
  INV_X1 U14005 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13234) );
  OAI22_X1 U14006 ( .A1(n10936), .A2(n14551), .B1(n10302), .B2(n13234), .ZN(
        n10937) );
  AOI21_X1 U14007 ( .B1(n10926), .B2(P2_EBX_REG_30__SCAN_IN), .A(n10937), .ZN(
        n10938) );
  AOI22_X1 U14008 ( .A1(n10940), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n10942) );
  NAND2_X1 U14009 ( .A1(n9599), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n10941) );
  OAI211_X1 U14010 ( .C1(n10943), .C2(n10855), .A(n10942), .B(n10941), .ZN(
        n10944) );
  NOR2_X1 U14011 ( .A1(n15276), .A2(n16247), .ZN(n10948) );
  INV_X1 U14012 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15484) );
  NAND2_X1 U14013 ( .A1(n13189), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13210) );
  INV_X1 U14014 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15467) );
  NAND2_X1 U14015 ( .A1(n13212), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13187) );
  INV_X1 U14016 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15432) );
  XNOR2_X1 U14017 ( .A(n10945), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13186) );
  NAND2_X1 U14018 ( .A1(n19113), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n11316) );
  NAND2_X1 U14019 ( .A1(n19114), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10946) );
  OAI211_X1 U14020 ( .C1(n19125), .C2(n13186), .A(n11316), .B(n10946), .ZN(
        n10947) );
  NOR2_X1 U14021 ( .A1(n10948), .A2(n10947), .ZN(n10949) );
  NAND3_X1 U14022 ( .A1(n10951), .A2(n10950), .A3(n10949), .ZN(P2_U2983) );
  OAI21_X1 U14023 ( .B1(n10957), .B2(n10955), .A(n9883), .ZN(n10954) );
  INV_X1 U14024 ( .A(n10952), .ZN(n10953) );
  NAND2_X1 U14025 ( .A1(n11284), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11285) );
  OAI21_X1 U14026 ( .B1(n10957), .B2(n10956), .A(n10955), .ZN(n10958) );
  NAND2_X1 U14027 ( .A1(n11285), .A2(n10958), .ZN(n10961) );
  XNOR2_X1 U14028 ( .A(n10959), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10960) );
  MUX2_X1 U14029 ( .A(n10962), .B(n10217), .S(n10383), .Z(n10963) );
  INV_X1 U14030 ( .A(READY21_REG_SCAN_IN), .ZN(n20830) );
  INV_X1 U14031 ( .A(READY12_REG_SCAN_IN), .ZN(n20849) );
  NOR2_X1 U14032 ( .A1(n20830), .A2(n20849), .ZN(n19849) );
  INV_X1 U14033 ( .A(n19849), .ZN(n19721) );
  NAND2_X1 U14034 ( .A1(n10963), .A2(n19721), .ZN(n10977) );
  NOR2_X1 U14035 ( .A1(n19722), .A2(n19740), .ZN(n19731) );
  NOR2_X1 U14036 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19733) );
  NOR3_X1 U14037 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19731), .A3(n19733), 
        .ZN(n19845) );
  NAND2_X1 U14038 ( .A1(n19721), .A2(n19845), .ZN(n13970) );
  INV_X1 U14039 ( .A(n13970), .ZN(n16347) );
  NAND2_X1 U14040 ( .A1(n10962), .A2(n16347), .ZN(n10964) );
  OR2_X1 U14041 ( .A1(n16337), .A2(n10964), .ZN(n10976) );
  NAND2_X1 U14042 ( .A1(n10967), .A2(n10264), .ZN(n10968) );
  NAND2_X1 U14043 ( .A1(n10966), .A2(n10968), .ZN(n10975) );
  NOR2_X1 U14044 ( .A1(n10251), .A2(n13297), .ZN(n11015) );
  OAI21_X1 U14045 ( .B1(n11015), .B2(n10274), .A(n10252), .ZN(n10969) );
  NAND2_X1 U14046 ( .A1(n10969), .A2(n10264), .ZN(n10973) );
  OR2_X1 U14047 ( .A1(n19844), .A2(n10970), .ZN(n11019) );
  AND4_X1 U14048 ( .A1(n10973), .A2(n11019), .A3(n10972), .A4(n10971), .ZN(
        n10974) );
  AND2_X1 U14049 ( .A1(n10976), .A2(n11016), .ZN(n13974) );
  OAI21_X1 U14050 ( .B1(n16337), .B2(n10977), .A(n13974), .ZN(n10978) );
  NOR2_X1 U14051 ( .A1(n10979), .A2(n10978), .ZN(n11007) );
  NAND2_X1 U14052 ( .A1(n13324), .A2(n13297), .ZN(n10980) );
  MUX2_X1 U14053 ( .A(n10980), .B(n13221), .S(n10981), .Z(n10990) );
  NAND2_X1 U14054 ( .A1(n10276), .A2(n10981), .ZN(n10988) );
  OAI21_X1 U14055 ( .B1(n10983), .B2(n10982), .A(n19833), .ZN(n10987) );
  INV_X1 U14056 ( .A(n10983), .ZN(n10985) );
  OAI211_X1 U14057 ( .C1(n13297), .C2(n10985), .A(n19846), .B(n10984), .ZN(
        n10986) );
  NAND3_X1 U14058 ( .A1(n10988), .A2(n10987), .A3(n10986), .ZN(n10989) );
  NAND2_X1 U14059 ( .A1(n10990), .A2(n10989), .ZN(n10993) );
  INV_X1 U14060 ( .A(n10991), .ZN(n10992) );
  NAND2_X1 U14061 ( .A1(n10993), .A2(n10992), .ZN(n10994) );
  OAI21_X1 U14062 ( .B1(n10995), .B2(n19833), .A(n10994), .ZN(n10996) );
  OAI21_X1 U14063 ( .B1(n13221), .B2(n10997), .A(n10996), .ZN(n10998) );
  NAND2_X1 U14064 ( .A1(n10999), .A2(n10259), .ZN(n11000) );
  INV_X1 U14065 ( .A(n11001), .ZN(n11002) );
  NAND2_X1 U14066 ( .A1(n13322), .A2(n11002), .ZN(n11003) );
  OAI21_X1 U14067 ( .B1(n19846), .B2(n16340), .A(n11003), .ZN(n11004) );
  NAND2_X1 U14068 ( .A1(n11004), .A2(n11021), .ZN(n11006) );
  INV_X1 U14069 ( .A(n13322), .ZN(n13972) );
  NAND3_X1 U14070 ( .A1(n13972), .A2(n10217), .A3(n16347), .ZN(n11005) );
  NAND3_X1 U14071 ( .A1(n11007), .A2(n11006), .A3(n11005), .ZN(n11008) );
  AND2_X1 U14072 ( .A1(n11013), .A2(n19833), .ZN(n11009) );
  NAND2_X1 U14073 ( .A1(n12848), .A2(n16300), .ZN(n11280) );
  AND2_X1 U14074 ( .A1(n11013), .A2(n19831), .ZN(n11014) );
  NAND2_X1 U14075 ( .A1(n11258), .A2(n16334), .ZN(n19147) );
  NAND2_X1 U14076 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15796) );
  AND2_X1 U14077 ( .A1(n11034), .A2(n15796), .ZN(n19127) );
  MUX2_X1 U14078 ( .A(n11017), .B(n10264), .S(n10274), .Z(n11031) );
  NAND2_X1 U14079 ( .A1(n11018), .A2(n13297), .ZN(n13964) );
  NAND2_X1 U14080 ( .A1(n13964), .A2(n11019), .ZN(n11024) );
  NAND2_X1 U14081 ( .A1(n11020), .A2(n10276), .ZN(n13146) );
  INV_X1 U14082 ( .A(n13145), .ZN(n13274) );
  OAI21_X1 U14083 ( .B1(n11027), .B2(n11021), .A(n13274), .ZN(n11022) );
  NAND2_X1 U14084 ( .A1(n13146), .A2(n11022), .ZN(n11023) );
  AOI21_X1 U14085 ( .B1(n11025), .B2(n11024), .A(n11023), .ZN(n11030) );
  INV_X1 U14086 ( .A(n11026), .ZN(n11028) );
  NAND2_X1 U14087 ( .A1(n11028), .A2(n11027), .ZN(n11029) );
  INV_X1 U14088 ( .A(n11032), .ZN(n13177) );
  NAND2_X1 U14089 ( .A1(n15801), .A2(n13177), .ZN(n11033) );
  NOR2_X1 U14090 ( .A1(n11034), .A2(n15796), .ZN(n19126) );
  INV_X1 U14091 ( .A(n19126), .ZN(n11035) );
  OR2_X1 U14092 ( .A1(n19128), .A2(n11035), .ZN(n11036) );
  OAI21_X1 U14093 ( .B1(n19147), .B2(n19127), .A(n11036), .ZN(n13826) );
  NAND2_X1 U14094 ( .A1(n13826), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14197) );
  NOR2_X1 U14095 ( .A1(n14200), .A2(n14199), .ZN(n14198) );
  INV_X1 U14096 ( .A(n14198), .ZN(n11260) );
  NOR2_X1 U14097 ( .A1(n14342), .A2(n11038), .ZN(n16308) );
  AND2_X1 U14098 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11039) );
  NAND2_X1 U14099 ( .A1(n15731), .A2(n11039), .ZN(n11264) );
  INV_X1 U14100 ( .A(n11264), .ZN(n11040) );
  INV_X1 U14101 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15713) );
  NOR3_X1 U14102 ( .A1(n15702), .A2(n10667), .A3(n15713), .ZN(n15689) );
  AND2_X1 U14103 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15689), .ZN(
        n11041) );
  NAND2_X1 U14104 ( .A1(n16268), .A2(n11041), .ZN(n15677) );
  NOR2_X1 U14105 ( .A1(n15654), .A2(n11269), .ZN(n15641) );
  AND2_X1 U14106 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11271) );
  NAND2_X1 U14107 ( .A1(n15641), .A2(n11271), .ZN(n15618) );
  NAND2_X1 U14108 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11273) );
  NAND3_X1 U14109 ( .A1(n15579), .A2(n15583), .A3(n11043), .ZN(n11256) );
  OR2_X1 U14110 ( .A1(n11045), .A2(n11046), .ZN(n11047) );
  NAND2_X1 U14111 ( .A1(n11044), .A2(n11047), .ZN(n15287) );
  INV_X1 U14112 ( .A(n15287), .ZN(n11254) );
  NAND2_X1 U14113 ( .A1(n11048), .A2(n10383), .ZN(n11051) );
  INV_X1 U14114 ( .A(n11049), .ZN(n11050) );
  NAND2_X1 U14115 ( .A1(n11051), .A2(n11050), .ZN(n11052) );
  NAND2_X1 U14116 ( .A1(n11258), .A2(n11052), .ZN(n19138) );
  AND2_X1 U14117 ( .A1(n13148), .A2(n11308), .ZN(n11068) );
  MUX2_X1 U14118 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n19167), .S(
        n19839), .Z(n11053) );
  INV_X1 U14119 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18988) );
  OAI21_X1 U14120 ( .B1(n10383), .B2(n13304), .A(n19839), .ZN(n11056) );
  NAND2_X1 U14121 ( .A1(n19167), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n11057) );
  AND2_X2 U14122 ( .A1(n19167), .A2(n19839), .ZN(n11230) );
  AOI22_X1 U14123 ( .A1(n11230), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11308), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11059) );
  OAI21_X1 U14124 ( .B1(n11307), .B2(n10272), .A(n11059), .ZN(n11065) );
  NAND2_X1 U14125 ( .A1(n11060), .A2(n10252), .ZN(n11061) );
  MUX2_X1 U14126 ( .A(n19822), .B(n11061), .S(n19839), .Z(n11062) );
  OAI21_X1 U14127 ( .B1(n11063), .B2(n11077), .A(n11062), .ZN(n13756) );
  NOR2_X1 U14128 ( .A1(n13757), .A2(n13756), .ZN(n11067) );
  NOR2_X1 U14129 ( .A1(n11064), .A2(n11065), .ZN(n11066) );
  AOI21_X1 U14130 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(
        P2_STATE2_REG_3__SCAN_IN), .A(n11068), .ZN(n11069) );
  OAI21_X1 U14131 ( .B1(n11070), .B2(n11077), .A(n11069), .ZN(n11072) );
  XNOR2_X1 U14132 ( .A(n11073), .B(n11072), .ZN(n13752) );
  AOI22_X1 U14133 ( .A1(n11230), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11308), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11071) );
  OAI21_X1 U14134 ( .B1(n11307), .B2(n13397), .A(n11071), .ZN(n13751) );
  NOR2_X1 U14135 ( .A1(n13752), .A2(n13751), .ZN(n13753) );
  NOR2_X1 U14136 ( .A1(n11073), .A2(n11072), .ZN(n11074) );
  NOR2_X2 U14137 ( .A1(n13753), .A2(n11074), .ZN(n13823) );
  NAND2_X1 U14138 ( .A1(n11230), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11075) );
  OAI21_X1 U14139 ( .B1(n11077), .B2(n11076), .A(n11075), .ZN(n11078) );
  INV_X1 U14140 ( .A(n11078), .ZN(n11080) );
  AOI22_X1 U14141 ( .A1(n11308), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11079) );
  OAI211_X1 U14142 ( .C1(n11307), .C2(n13817), .A(n11080), .B(n11079), .ZN(
        n13822) );
  AOI22_X1 U14143 ( .A1(n11230), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11308), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11083) );
  NAND2_X1 U14144 ( .A1(n11224), .A2(n11081), .ZN(n11082) );
  OAI211_X1 U14145 ( .C1(n11307), .C2(n11084), .A(n11083), .B(n11082), .ZN(
        n13904) );
  INV_X1 U14146 ( .A(n13904), .ZN(n11085) );
  AOI22_X1 U14147 ( .A1(n11230), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11308), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11088) );
  NAND2_X1 U14148 ( .A1(n11224), .A2(n11086), .ZN(n11087) );
  OAI211_X1 U14149 ( .C1(n11307), .C2(n11089), .A(n11088), .B(n11087), .ZN(
        n13997) );
  INV_X1 U14150 ( .A(n11090), .ZN(n11091) );
  NAND2_X1 U14151 ( .A1(n11224), .A2(n11091), .ZN(n11092) );
  AOI22_X1 U14152 ( .A1(n11230), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11308), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11093) );
  OAI21_X1 U14153 ( .B1(n11307), .B2(n14317), .A(n11093), .ZN(n13893) );
  NAND2_X1 U14154 ( .A1(n13892), .A2(n13893), .ZN(n11096) );
  NAND2_X1 U14155 ( .A1(n11224), .A2(n11094), .ZN(n11095) );
  AOI22_X1 U14156 ( .A1(n11230), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11308), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11097) );
  OAI21_X1 U14157 ( .B1(n11307), .B2(n10797), .A(n11097), .ZN(n14350) );
  AOI22_X1 U14158 ( .A1(n11230), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11308), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11112) );
  AOI22_X1 U14159 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10503), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11104) );
  INV_X1 U14160 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11100) );
  NAND2_X1 U14161 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11099) );
  AOI22_X1 U14162 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12982), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11098) );
  OAI211_X1 U14163 ( .C1(n12987), .C2(n11100), .A(n11099), .B(n11098), .ZN(
        n11101) );
  INV_X1 U14164 ( .A(n11101), .ZN(n11103) );
  AOI22_X1 U14165 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11102) );
  NAND3_X1 U14166 ( .A1(n11104), .A2(n11103), .A3(n11102), .ZN(n11110) );
  AOI22_X1 U14167 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11108) );
  AOI22_X1 U14168 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11107) );
  AOI22_X1 U14169 ( .A1(n10410), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11106) );
  AOI22_X1 U14170 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11105) );
  NAND4_X1 U14171 ( .A1(n11108), .A2(n11107), .A3(n11106), .A4(n11105), .ZN(
        n11109) );
  NAND2_X1 U14172 ( .A1(n11224), .A2(n13722), .ZN(n11111) );
  OAI211_X1 U14173 ( .C1(n11307), .C2(n11113), .A(n11112), .B(n11111), .ZN(
        n13867) );
  INV_X1 U14174 ( .A(n13867), .ZN(n11114) );
  AOI22_X1 U14175 ( .A1(n11230), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11308), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11129) );
  AOI22_X1 U14176 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10503), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11121) );
  NAND2_X1 U14177 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11116) );
  AOI22_X1 U14178 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n12982), .ZN(n11115) );
  OAI211_X1 U14179 ( .C1(n12987), .C2(n11117), .A(n11116), .B(n11115), .ZN(
        n11118) );
  INV_X1 U14180 ( .A(n11118), .ZN(n11120) );
  AOI22_X1 U14181 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n10434), .ZN(n11119) );
  NAND3_X1 U14182 ( .A1(n11121), .A2(n11120), .A3(n11119), .ZN(n11127) );
  AOI22_X1 U14183 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11125) );
  AOI22_X1 U14184 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11124) );
  AOI22_X1 U14185 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10410), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11123) );
  AOI22_X1 U14186 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10516), .B1(
        n10445), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11122) );
  NAND4_X1 U14187 ( .A1(n11125), .A2(n11124), .A3(n11123), .A4(n11122), .ZN(
        n11126) );
  NAND2_X1 U14188 ( .A1(n11224), .A2(n13721), .ZN(n11128) );
  OAI211_X1 U14189 ( .C1(n11307), .C2(n11130), .A(n11129), .B(n11128), .ZN(
        n15778) );
  AOI22_X1 U14190 ( .A1(n11230), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11308), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11145) );
  AOI22_X1 U14191 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11137) );
  INV_X1 U14192 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11133) );
  NAND2_X1 U14193 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11132) );
  AOI22_X1 U14194 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n12982), .ZN(n11131) );
  OAI211_X1 U14195 ( .C1(n12987), .C2(n11133), .A(n11132), .B(n11131), .ZN(
        n11134) );
  INV_X1 U14196 ( .A(n11134), .ZN(n11136) );
  AOI22_X1 U14197 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__2__SCAN_IN), .B2(n10440), .ZN(n11135) );
  NAND3_X1 U14198 ( .A1(n11137), .A2(n11136), .A3(n11135), .ZN(n11143) );
  AOI22_X1 U14199 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10503), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11141) );
  AOI22_X1 U14200 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__2__SCAN_IN), .B2(n10434), .ZN(n11140) );
  AOI22_X1 U14201 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10410), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11139) );
  AOI22_X1 U14202 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10516), .B1(
        n10418), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11138) );
  NAND4_X1 U14203 ( .A1(n11141), .A2(n11140), .A3(n11139), .A4(n11138), .ZN(
        n11142) );
  NAND2_X1 U14204 ( .A1(n11224), .A2(n13565), .ZN(n11144) );
  OAI211_X1 U14205 ( .C1(n11307), .C2(n11146), .A(n11145), .B(n11144), .ZN(
        n13882) );
  INV_X1 U14206 ( .A(n13882), .ZN(n11147) );
  AOI22_X1 U14207 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10503), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11154) );
  NAND2_X1 U14208 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11149) );
  AOI22_X1 U14209 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n12982), .ZN(n11148) );
  OAI211_X1 U14210 ( .C1(n12987), .C2(n11150), .A(n11149), .B(n11148), .ZN(
        n11151) );
  INV_X1 U14211 ( .A(n11151), .ZN(n11153) );
  AOI22_X1 U14212 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__3__SCAN_IN), .B2(n10434), .ZN(n11152) );
  NAND3_X1 U14213 ( .A1(n11154), .A2(n11153), .A3(n11152), .ZN(n11160) );
  AOI22_X1 U14214 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11158) );
  AOI22_X1 U14215 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11157) );
  AOI22_X1 U14216 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10410), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11156) );
  AOI22_X1 U14217 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10516), .B1(
        n10445), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11155) );
  NAND4_X1 U14218 ( .A1(n11158), .A2(n11157), .A3(n11156), .A4(n11155), .ZN(
        n11159) );
  AOI22_X1 U14219 ( .A1(n11309), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n11224), 
        .B2(n13732), .ZN(n11162) );
  AOI22_X1 U14220 ( .A1(n11230), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11308), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11161) );
  NAND2_X1 U14221 ( .A1(n11162), .A2(n11161), .ZN(n13846) );
  NAND2_X1 U14222 ( .A1(n13844), .A2(n13846), .ZN(n13845) );
  AOI22_X1 U14223 ( .A1(n11230), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11308), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11175) );
  AOI22_X1 U14224 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10460), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11167) );
  NAND2_X1 U14225 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11165) );
  NAND2_X1 U14226 ( .A1(n10434), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11164) );
  AOI22_X1 U14227 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12982), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11163) );
  AOI22_X1 U14228 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10491), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11166) );
  NAND3_X1 U14229 ( .A1(n11167), .A2(n9668), .A3(n11166), .ZN(n11173) );
  AOI22_X1 U14230 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11178), .B1(
        n10444), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11171) );
  AOI22_X1 U14231 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10503), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11170) );
  AOI22_X1 U14232 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n10410), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11169) );
  AOI22_X1 U14233 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10516), .B1(
        n10445), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11168) );
  NAND4_X1 U14234 ( .A1(n11171), .A2(n11170), .A3(n11169), .A4(n11168), .ZN(
        n11172) );
  NAND2_X1 U14235 ( .A1(n11224), .A2(n13609), .ZN(n11174) );
  OAI211_X1 U14236 ( .C1(n11307), .C2(n11176), .A(n11175), .B(n11174), .ZN(
        n11177) );
  INV_X1 U14237 ( .A(n11177), .ZN(n13913) );
  AOI22_X1 U14239 ( .A1(n11230), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11308), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11193) );
  AOI22_X1 U14240 ( .A1(n11178), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10444), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11185) );
  NAND2_X1 U14241 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11179) );
  OAI21_X1 U14242 ( .B1(n14295), .B2(n11180), .A(n11179), .ZN(n11181) );
  AOI21_X1 U14243 ( .B1(n10503), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n11181), .ZN(n11184) );
  AOI22_X1 U14244 ( .A1(n10491), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11183) );
  NAND2_X1 U14245 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11182) );
  NAND4_X1 U14246 ( .A1(n11185), .A2(n11184), .A3(n11183), .A4(n11182), .ZN(
        n11191) );
  AOI22_X1 U14247 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11189) );
  AOI22_X1 U14248 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11188) );
  AOI22_X1 U14249 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10410), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11187) );
  AOI22_X1 U14250 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11186) );
  NAND4_X1 U14251 ( .A1(n11189), .A2(n11188), .A3(n11187), .A4(n11186), .ZN(
        n11190) );
  NAND2_X1 U14252 ( .A1(n11224), .A2(n9679), .ZN(n11192) );
  OAI211_X1 U14253 ( .C1(n11307), .C2(n14042), .A(n11193), .B(n11192), .ZN(
        n14038) );
  NAND2_X1 U14254 ( .A1(n14037), .A2(n14038), .ZN(n14039) );
  AOI22_X1 U14255 ( .A1(n11230), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11308), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11208) );
  AOI22_X1 U14256 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10503), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11200) );
  NAND2_X1 U14257 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11195) );
  AOI22_X1 U14258 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n12982), .ZN(n11194) );
  OAI211_X1 U14259 ( .C1(n12987), .C2(n11196), .A(n11195), .B(n11194), .ZN(
        n11197) );
  INV_X1 U14260 ( .A(n11197), .ZN(n11199) );
  AOI22_X1 U14261 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__6__SCAN_IN), .B2(n10434), .ZN(n11198) );
  NAND3_X1 U14262 ( .A1(n11200), .A2(n11199), .A3(n11198), .ZN(n11206) );
  AOI22_X1 U14263 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11204) );
  AOI22_X1 U14264 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11203) );
  AOI22_X1 U14265 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n10410), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11202) );
  AOI22_X1 U14266 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10516), .B1(
        n10445), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11201) );
  NAND4_X1 U14267 ( .A1(n11204), .A2(n11203), .A3(n11202), .A4(n11201), .ZN(
        n11205) );
  NAND2_X1 U14268 ( .A1(n11224), .A2(n13836), .ZN(n11207) );
  OAI211_X1 U14269 ( .C1(n11307), .C2(n11209), .A(n11208), .B(n11207), .ZN(
        n11210) );
  INV_X1 U14270 ( .A(n11210), .ZN(n15733) );
  INV_X1 U14271 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n11227) );
  AOI22_X1 U14272 ( .A1(n11230), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11308), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11226) );
  AOI22_X1 U14273 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10503), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11217) );
  AOI22_X1 U14274 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11216) );
  INV_X1 U14275 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11213) );
  NAND2_X1 U14276 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11212) );
  AOI22_X1 U14277 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n12982), .ZN(n11211) );
  OAI211_X1 U14278 ( .C1(n12987), .C2(n11213), .A(n11212), .B(n11211), .ZN(
        n11214) );
  INV_X1 U14279 ( .A(n11214), .ZN(n11215) );
  NAND3_X1 U14280 ( .A1(n11217), .A2(n11216), .A3(n11215), .ZN(n11223) );
  AOI22_X1 U14281 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11221) );
  AOI22_X1 U14282 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n10434), .ZN(n11220) );
  AOI22_X1 U14283 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10410), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11219) );
  AOI22_X1 U14284 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10516), .B1(
        n10445), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11218) );
  NAND4_X1 U14285 ( .A1(n11221), .A2(n11220), .A3(n11219), .A4(n11218), .ZN(
        n11222) );
  NAND2_X1 U14286 ( .A1(n11224), .A2(n13955), .ZN(n11225) );
  OAI211_X1 U14287 ( .C1(n11307), .C2(n11227), .A(n11226), .B(n11225), .ZN(
        n14241) );
  INV_X1 U14288 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n11229) );
  AOI22_X1 U14289 ( .A1(n11230), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11308), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11228) );
  OAI21_X1 U14290 ( .B1(n11307), .B2(n11229), .A(n11228), .ZN(n15716) );
  INV_X1 U14291 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14254) );
  OAI22_X1 U14292 ( .A1(n11303), .A2(n14254), .B1(n11302), .B2(n15702), .ZN(
        n11231) );
  AOI21_X1 U14293 ( .B1(n11309), .B2(P2_REIP_REG_17__SCAN_IN), .A(n11231), 
        .ZN(n14256) );
  INV_X1 U14294 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n11232) );
  OAI22_X1 U14295 ( .A1(n11303), .A2(n11232), .B1(n11302), .B2(n15688), .ZN(
        n11233) );
  AOI21_X1 U14296 ( .B1(n11309), .B2(P2_REIP_REG_18__SCAN_IN), .A(n11233), 
        .ZN(n15684) );
  INV_X1 U14297 ( .A(n15684), .ZN(n11234) );
  INV_X1 U14298 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19760) );
  AOI22_X1 U14299 ( .A1(n11230), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11308), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11235) );
  OAI21_X1 U14300 ( .B1(n11307), .B2(n19760), .A(n11235), .ZN(n15270) );
  INV_X1 U14301 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n15509) );
  AOI22_X1 U14302 ( .A1(n11230), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11308), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11236) );
  OAI21_X1 U14303 ( .B1(n11307), .B2(n15509), .A(n11236), .ZN(n15661) );
  INV_X1 U14304 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15403) );
  OAI22_X1 U14305 ( .A1(n11303), .A2(n15403), .B1(n11302), .B2(n11269), .ZN(
        n11237) );
  AOI21_X1 U14306 ( .B1(n11309), .B2(P2_REIP_REG_21__SCAN_IN), .A(n11237), 
        .ZN(n15402) );
  INV_X1 U14307 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n11238) );
  OAI22_X1 U14308 ( .A1(n11303), .A2(n11238), .B1(n11302), .B2(n15640), .ZN(
        n11239) );
  AOI21_X1 U14309 ( .B1(n11309), .B2(P2_REIP_REG_22__SCAN_IN), .A(n11239), 
        .ZN(n15394) );
  INV_X1 U14310 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19767) );
  AOI22_X1 U14311 ( .A1(n11230), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11308), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11240) );
  OAI21_X1 U14312 ( .B1(n11307), .B2(n19767), .A(n11240), .ZN(n15249) );
  AND2_X2 U14313 ( .A1(n15248), .A2(n15249), .ZN(n15247) );
  INV_X1 U14314 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19769) );
  AOI22_X1 U14315 ( .A1(n11230), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11308), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11241) );
  OAI21_X1 U14316 ( .B1(n11307), .B2(n19769), .A(n11241), .ZN(n15382) );
  INV_X1 U14317 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n15376) );
  OAI22_X1 U14318 ( .A1(n11303), .A2(n15376), .B1(n11302), .B2(n15464), .ZN(
        n11242) );
  AOI21_X1 U14319 ( .B1(n11309), .B2(P2_REIP_REG_25__SCAN_IN), .A(n11242), 
        .ZN(n15235) );
  INV_X1 U14320 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n15370) );
  INV_X1 U14321 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11243) );
  OAI22_X1 U14322 ( .A1(n11303), .A2(n15370), .B1(n11302), .B2(n11243), .ZN(
        n11244) );
  AOI21_X1 U14323 ( .B1(n11309), .B2(P2_REIP_REG_26__SCAN_IN), .A(n11244), 
        .ZN(n15214) );
  INV_X1 U14324 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n20882) );
  OAI22_X1 U14325 ( .A1(n11303), .A2(n20882), .B1(n11302), .B2(n11289), .ZN(
        n11245) );
  AOI21_X1 U14326 ( .B1(n11309), .B2(P2_REIP_REG_27__SCAN_IN), .A(n11245), 
        .ZN(n11290) );
  AOI22_X1 U14327 ( .A1(n11230), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11308), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11246) );
  OAI21_X1 U14328 ( .B1(n11307), .B2(n19776), .A(n11246), .ZN(n11247) );
  OR2_X1 U14329 ( .A1(n11292), .A2(n11247), .ZN(n11248) );
  NAND2_X1 U14330 ( .A1(n11305), .A2(n11248), .ZN(n15360) );
  AND2_X1 U14331 ( .A1(n10966), .A2(n13227), .ZN(n16336) );
  INV_X1 U14332 ( .A(n11249), .ZN(n11251) );
  NAND2_X1 U14333 ( .A1(n11251), .A2(n11250), .ZN(n13176) );
  OAI21_X1 U14334 ( .B1(n16336), .B2(n10364), .A(n13176), .ZN(n11252) );
  OR2_X1 U14335 ( .A1(n15534), .A2(n19776), .ZN(n12851) );
  OAI21_X1 U14336 ( .B1(n15360), .B2(n19143), .A(n12851), .ZN(n11253) );
  AOI21_X1 U14337 ( .B1(n11254), .B2(n16302), .A(n11253), .ZN(n11255) );
  NAND2_X1 U14338 ( .A1(n11256), .A2(n11255), .ZN(n11278) );
  AND2_X2 U14339 ( .A1(n19147), .A2(n19128), .ZN(n15766) );
  INV_X1 U14340 ( .A(n19147), .ZN(n11259) );
  INV_X1 U14341 ( .A(n11257), .ZN(n16279) );
  NOR2_X1 U14342 ( .A1(n11258), .A2(n16279), .ZN(n19130) );
  OAI21_X1 U14343 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15766), .A(
        n13827), .ZN(n14203) );
  AOI21_X1 U14344 ( .B1(n15797), .B2(n11260), .A(n14203), .ZN(n14316) );
  NOR2_X1 U14345 ( .A1(n11261), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14321) );
  INV_X1 U14346 ( .A(n14321), .ZN(n11262) );
  NAND2_X1 U14347 ( .A1(n14316), .A2(n11262), .ZN(n16299) );
  NOR2_X1 U14348 ( .A1(n15766), .A2(n16308), .ZN(n11263) );
  NAND2_X1 U14349 ( .A1(n15797), .A2(n11264), .ZN(n11265) );
  NOR2_X1 U14350 ( .A1(n15766), .A2(n15689), .ZN(n11266) );
  NOR2_X1 U14351 ( .A1(n15766), .A2(n11267), .ZN(n11268) );
  NAND2_X1 U14352 ( .A1(n15797), .A2(n11269), .ZN(n11270) );
  NAND2_X1 U14353 ( .A1(n15651), .A2(n11270), .ZN(n15646) );
  OAI21_X1 U14354 ( .B1(n15766), .B2(n11271), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11272) );
  OR2_X1 U14355 ( .A1(n15646), .A2(n11272), .ZN(n15616) );
  NAND2_X1 U14356 ( .A1(n15651), .A2(n15766), .ZN(n11313) );
  NAND2_X1 U14357 ( .A1(n15616), .A2(n11313), .ZN(n15591) );
  NAND2_X1 U14358 ( .A1(n11313), .A2(n11273), .ZN(n11274) );
  NAND2_X1 U14359 ( .A1(n15591), .A2(n11274), .ZN(n15572) );
  NOR2_X1 U14360 ( .A1(n11276), .A2(n11275), .ZN(n11277) );
  NAND3_X1 U14361 ( .A1(n11280), .A2(n9649), .A3(n11279), .ZN(P2_U3018) );
  INV_X1 U14362 ( .A(n11281), .ZN(n11283) );
  INV_X1 U14363 ( .A(n11011), .ZN(n11282) );
  OR2_X1 U14364 ( .A1(n11284), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15444) );
  NAND3_X1 U14365 ( .A1(n15444), .A2(n11285), .A3(n16300), .ZN(n11299) );
  NOR2_X1 U14366 ( .A1(n11286), .A2(n11287), .ZN(n11288) );
  NAND2_X1 U14367 ( .A1(n15579), .A2(n11289), .ZN(n11295) );
  AND2_X1 U14368 ( .A1(n15216), .A2(n11290), .ZN(n11291) );
  NOR2_X1 U14369 ( .A1(n11292), .A2(n11291), .ZN(n15365) );
  OR2_X1 U14370 ( .A1(n15534), .A2(n19775), .ZN(n15438) );
  INV_X1 U14371 ( .A(n15438), .ZN(n11293) );
  AOI21_X1 U14372 ( .B1(n15365), .B2(n16298), .A(n11293), .ZN(n11294) );
  OAI211_X1 U14373 ( .C1(n15440), .C2(n19138), .A(n11295), .B(n11294), .ZN(
        n11296) );
  INV_X1 U14374 ( .A(n11296), .ZN(n11298) );
  NAND2_X1 U14375 ( .A1(n15572), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11297) );
  NAND4_X1 U14376 ( .A1(n9644), .A2(n11299), .A3(n11298), .A4(n11297), .ZN(
        P2_U3019) );
  INV_X1 U14377 ( .A(n11300), .ZN(n11301) );
  INV_X1 U14378 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n15352) );
  OAI22_X1 U14379 ( .A1(n11303), .A2(n15352), .B1(n11302), .B2(n15582), .ZN(
        n11304) );
  AOI21_X1 U14380 ( .B1(n11309), .B2(P2_REIP_REG_29__SCAN_IN), .A(n11304), 
        .ZN(n15180) );
  AOI22_X1 U14381 ( .A1(n11230), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11308), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11306) );
  OAI21_X1 U14382 ( .B1(n11307), .B2(n14551), .A(n11306), .ZN(n13170) );
  AOI222_X1 U14383 ( .A1(n11309), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n11308), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C1(n11230), .C2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n11310) );
  XNOR2_X2 U14384 ( .A(n13168), .B(n11310), .ZN(n19004) );
  NOR2_X1 U14385 ( .A1(n15582), .A2(n15583), .ZN(n15581) );
  INV_X1 U14386 ( .A(n15581), .ZN(n11312) );
  AOI211_X1 U14387 ( .C1(n11313), .C2(n11312), .A(n11311), .B(n15572), .ZN(
        n14550) );
  INV_X1 U14388 ( .A(n11313), .ZN(n11314) );
  NOR3_X1 U14389 ( .A1(n14550), .A2(n11314), .A3(n10855), .ZN(n11315) );
  NOR2_X1 U14390 ( .A1(n11315), .A2(n10116), .ZN(n11317) );
  INV_X1 U14391 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11320) );
  AOI22_X1 U14392 ( .A1(n11386), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11435), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14393 ( .A1(n11362), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11335), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11324) );
  AND2_X2 U14394 ( .A1(n13640), .A2(n13436), .ZN(n12342) );
  AND2_X4 U14395 ( .A1(n11327), .A2(n13435), .ZN(n12290) );
  AOI22_X1 U14396 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11323) );
  AOI22_X1 U14397 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11345), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11322) );
  NAND2_X2 U14398 ( .A1(n13638), .A2(n11326), .ZN(n11350) );
  INV_X2 U14399 ( .A(n11350), .ZN(n11710) );
  AOI22_X1 U14400 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11412), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11332) );
  AND2_X2 U14401 ( .A1(n11326), .A2(n11327), .ZN(n11447) );
  AOI22_X1 U14402 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11447), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U14404 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11554), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11330) );
  AND2_X2 U14405 ( .A1(n13436), .A2(n11327), .ZN(n11415) );
  AOI22_X1 U14406 ( .A1(n11415), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11407), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11329) );
  NAND2_X2 U14407 ( .A1(n11334), .A2(n11333), .ZN(n11536) );
  AOI22_X1 U14408 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11345), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11339) );
  AOI22_X1 U14409 ( .A1(n11386), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11435), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U14410 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11447), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14411 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11412), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U14412 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11554), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11341) );
  AOI22_X1 U14413 ( .A1(n11415), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11407), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11340) );
  BUF_X4 U14414 ( .A(n11345), .Z(n12477) );
  AOI22_X1 U14415 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11349) );
  INV_X2 U14416 ( .A(n13637), .ZN(n12381) );
  AOI22_X1 U14417 ( .A1(n11362), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12381), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11348) );
  AOI22_X1 U14418 ( .A1(n11386), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11435), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11347) );
  AOI22_X1 U14419 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11346) );
  NAND4_X1 U14420 ( .A1(n11349), .A2(n11348), .A3(n11347), .A4(n11346), .ZN(
        n11356) );
  AOI22_X1 U14421 ( .A1(n12273), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11412), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11354) );
  AOI22_X1 U14422 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11447), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14423 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11554), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U14424 ( .A1(n12422), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11407), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11351) );
  NAND4_X1 U14425 ( .A1(n11354), .A2(n11353), .A3(n11352), .A4(n11351), .ZN(
        n11355) );
  NAND2_X1 U14426 ( .A1(n11357), .A2(n11563), .ZN(n11380) );
  NAND2_X1 U14427 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11361) );
  NAND2_X1 U14428 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11360) );
  NAND2_X1 U14429 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11359) );
  NAND2_X1 U14430 ( .A1(n11554), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11358) );
  NAND2_X1 U14431 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11366) );
  NAND2_X1 U14432 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11365) );
  NAND2_X1 U14433 ( .A1(n11362), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11364) );
  NAND2_X1 U14434 ( .A1(n11345), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11363) );
  NAND2_X1 U14435 ( .A1(n11447), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11370) );
  NAND2_X1 U14436 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11369) );
  NAND2_X1 U14437 ( .A1(n11415), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11368) );
  NAND2_X1 U14438 ( .A1(n11407), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11367) );
  NAND2_X1 U14439 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11374) );
  NAND2_X1 U14440 ( .A1(n11386), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11373) );
  NAND2_X1 U14441 ( .A1(n11435), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11372) );
  NAND2_X1 U14442 ( .A1(n12290), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11371) );
  INV_X1 U14443 ( .A(n11381), .ZN(n11500) );
  NAND2_X1 U14444 ( .A1(n11536), .A2(n11500), .ZN(n11481) );
  INV_X1 U14445 ( .A(n11481), .ZN(n11405) );
  NAND2_X1 U14446 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11385) );
  NAND2_X1 U14447 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11384) );
  NAND2_X1 U14448 ( .A1(n11447), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11383) );
  NAND2_X1 U14449 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11382) );
  NAND2_X1 U14450 ( .A1(n12381), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11390) );
  NAND2_X1 U14451 ( .A1(n11386), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11389) );
  NAND2_X1 U14452 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11388) );
  NAND2_X1 U14453 ( .A1(n12290), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11387) );
  NAND2_X1 U14454 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11395) );
  NAND2_X1 U14455 ( .A1(n11362), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11394) );
  BUF_X4 U14456 ( .A(n11435), .Z(n12436) );
  NAND2_X1 U14457 ( .A1(n12436), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11393) );
  NAND2_X1 U14458 ( .A1(n11345), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11392) );
  NAND2_X1 U14459 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11399) );
  NAND2_X1 U14460 ( .A1(n11407), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11398) );
  NAND2_X1 U14461 ( .A1(n11415), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11397) );
  NAND2_X1 U14462 ( .A1(n11554), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11396) );
  NAND4_X4 U14463 ( .A1(n11403), .A2(n11402), .A3(n11401), .A4(n11400), .ZN(
        n12000) );
  NAND2_X1 U14464 ( .A1(n11483), .A2(n12000), .ZN(n11419) );
  NAND2_X1 U14465 ( .A1(n11405), .A2(n11404), .ZN(n11786) );
  AOI22_X1 U14466 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11407), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11411) );
  AOI22_X1 U14467 ( .A1(n11386), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11435), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14468 ( .A1(n11362), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11447), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11409) );
  AOI22_X1 U14469 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11408) );
  AOI22_X1 U14470 ( .A1(n12273), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11412), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U14471 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11554), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11413) );
  AOI22_X1 U14472 ( .A1(n12381), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U14473 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11416) );
  NAND2_X1 U14474 ( .A1(n11419), .A2(n11472), .ZN(n11467) );
  AND3_X2 U14475 ( .A1(n11421), .A2(n11420), .A3(n11467), .ZN(n11486) );
  NAND2_X1 U14476 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11426) );
  NAND2_X1 U14477 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11425) );
  NAND2_X1 U14478 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11424) );
  NAND2_X1 U14479 ( .A1(n11554), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11423) );
  NAND2_X1 U14480 ( .A1(n12381), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11430) );
  NAND2_X1 U14481 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11429) );
  NAND2_X1 U14482 ( .A1(n11362), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11428) );
  NAND2_X1 U14483 ( .A1(n12289), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11427) );
  NAND2_X1 U14484 ( .A1(n11447), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11434) );
  NAND2_X1 U14485 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11433) );
  NAND2_X1 U14486 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11432) );
  NAND2_X1 U14487 ( .A1(n11407), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11431) );
  NAND2_X1 U14488 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11439) );
  NAND2_X1 U14489 ( .A1(n11386), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11438) );
  BUF_X4 U14490 ( .A(n11435), .Z(n12394) );
  NAND2_X1 U14491 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11437) );
  NAND2_X1 U14492 ( .A1(n12290), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11436) );
  NOR2_X1 U14493 ( .A1(n11968), .A2(n20061), .ZN(n11442) );
  NAND2_X1 U14494 ( .A1(n11486), .A2(n11442), .ZN(n11788) );
  INV_X1 U14495 ( .A(n11788), .ZN(n11464) );
  NAND2_X1 U14496 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11446) );
  NAND2_X1 U14497 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11445) );
  NAND2_X1 U14498 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11444) );
  NAND2_X1 U14499 ( .A1(n11415), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11443) );
  NAND2_X1 U14500 ( .A1(n11335), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11451) );
  BUF_X4 U14501 ( .A(n11447), .Z(n12475) );
  NAND2_X1 U14502 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11450) );
  NAND2_X1 U14503 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11449) );
  NAND2_X1 U14504 ( .A1(n12290), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11448) );
  NAND2_X1 U14505 ( .A1(n11386), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11455) );
  NAND2_X1 U14506 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11454) );
  NAND2_X1 U14507 ( .A1(n12289), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11453) );
  NAND2_X1 U14508 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11452) );
  NAND2_X1 U14509 ( .A1(n11362), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11459) );
  NAND2_X1 U14510 ( .A1(n11406), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11458) );
  NAND2_X1 U14511 ( .A1(n11407), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11457) );
  NAND2_X1 U14512 ( .A1(n11554), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11456) );
  NAND2_X1 U14513 ( .A1(n11464), .A2(n15926), .ZN(n12511) );
  INV_X1 U14514 ( .A(n11467), .ZN(n11468) );
  AND2_X2 U14515 ( .A1(n11784), .A2(n11468), .ZN(n11854) );
  NAND2_X1 U14516 ( .A1(n20061), .A2(n11475), .ZN(n11894) );
  AND2_X2 U14517 ( .A1(n12511), .A2(n12514), .ZN(n11864) );
  NOR2_X1 U14518 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n11469) );
  NOR2_X1 U14519 ( .A1(n20646), .A2(n11469), .ZN(n11791) );
  NAND2_X1 U14520 ( .A1(n11866), .A2(n11791), .ZN(n11473) );
  NAND2_X1 U14521 ( .A1(n11471), .A2(n11470), .ZN(n12515) );
  OR2_X2 U14522 ( .A1(n12515), .A2(n11472), .ZN(n11867) );
  NAND3_X1 U14523 ( .A1(n11864), .A2(n11473), .A3(n11867), .ZN(n11474) );
  NAND2_X1 U14524 ( .A1(n11477), .A2(n20061), .ZN(n11971) );
  NAND2_X1 U14525 ( .A1(n11479), .A2(n20061), .ZN(n11879) );
  NAND2_X1 U14526 ( .A1(n13404), .A2(n11480), .ZN(n11972) );
  NAND2_X1 U14527 ( .A1(n11482), .A2(n11483), .ZN(n11484) );
  INV_X1 U14528 ( .A(n11783), .ZN(n11485) );
  NAND3_X1 U14529 ( .A1(n11494), .A2(n11972), .A3(n11485), .ZN(n11491) );
  INV_X1 U14530 ( .A(n11486), .ZN(n11493) );
  NAND2_X1 U14531 ( .A1(n11487), .A2(n15926), .ZN(n11488) );
  INV_X1 U14532 ( .A(n11638), .ZN(n11575) );
  OAI21_X1 U14533 ( .B1(n11493), .B2(n11488), .A(n11575), .ZN(n11489) );
  INV_X1 U14534 ( .A(n11489), .ZN(n11490) );
  INV_X1 U14535 ( .A(n20634), .ZN(n15932) );
  MUX2_X1 U14536 ( .A(n15932), .B(n13464), .S(n20499), .Z(n11492) );
  NAND2_X1 U14537 ( .A1(n11493), .A2(n11470), .ZN(n11975) );
  INV_X1 U14538 ( .A(n11495), .ZN(n11498) );
  NAND2_X1 U14539 ( .A1(n11482), .A2(n20061), .ZN(n11497) );
  NAND2_X1 U14540 ( .A1(n11537), .A2(n20076), .ZN(n14091) );
  NAND2_X1 U14541 ( .A1(n11496), .A2(n14091), .ZN(n13477) );
  OAI21_X1 U14542 ( .B1(n11498), .B2(n11497), .A(n13477), .ZN(n11503) );
  NAND2_X1 U14543 ( .A1(n14558), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19865) );
  INV_X1 U14544 ( .A(n19865), .ZN(n11502) );
  NAND2_X1 U14545 ( .A1(n11783), .A2(n20076), .ZN(n11504) );
  NAND3_X1 U14546 ( .A1(n11975), .A2(n11505), .A3(n11504), .ZN(n11545) );
  INV_X1 U14547 ( .A(n11545), .ZN(n11506) );
  AOI22_X1 U14548 ( .A1(n12273), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U14549 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11509) );
  INV_X1 U14550 ( .A(n11554), .ZN(n11519) );
  AOI22_X1 U14551 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n11518), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11508) );
  AOI22_X1 U14552 ( .A1(n12422), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11507) );
  NAND4_X1 U14553 ( .A1(n11510), .A2(n11509), .A3(n11508), .A4(n11507), .ZN(
        n11516) );
  AOI22_X1 U14554 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12435), .B1(
        n12381), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11514) );
  INV_X1 U14555 ( .A(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n20883) );
  AOI22_X1 U14556 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11513) );
  AOI22_X1 U14557 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n12485), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14558 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n12479), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11511) );
  NAND4_X1 U14559 ( .A1(n11514), .A2(n11513), .A3(n11512), .A4(n11511), .ZN(
        n11515) );
  NOR2_X1 U14560 ( .A1(n11637), .A2(n11745), .ZN(n11574) );
  INV_X1 U14561 ( .A(n11517), .ZN(n11553) );
  AOI22_X1 U14562 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11518), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U14563 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11522) );
  AOI22_X1 U14564 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11521) );
  AOI22_X1 U14565 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11520) );
  NAND4_X1 U14566 ( .A1(n11523), .A2(n11522), .A3(n11521), .A4(n11520), .ZN(
        n11529) );
  AOI22_X1 U14567 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U14568 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14569 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12478), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11525) );
  INV_X1 U14570 ( .A(n11350), .ZN(n12441) );
  AOI22_X1 U14571 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11524) );
  NAND4_X1 U14572 ( .A1(n11527), .A2(n11526), .A3(n11525), .A4(n11524), .ZN(
        n11528) );
  MUX2_X1 U14573 ( .A(n11742), .B(n11574), .S(n11619), .Z(n11530) );
  INV_X1 U14574 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11535) );
  INV_X1 U14575 ( .A(n11532), .ZN(n11821) );
  OAI21_X1 U14576 ( .B1(n11619), .B2(n20744), .A(n11821), .ZN(n11533) );
  NAND2_X1 U14577 ( .A1(n20093), .A2(n20076), .ZN(n11813) );
  OAI21_X1 U14578 ( .B1(n11496), .B2(n11619), .A(n11623), .ZN(n11538) );
  INV_X1 U14579 ( .A(n11538), .ZN(n11539) );
  NAND2_X1 U14580 ( .A1(n11584), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11542) );
  NAND2_X1 U14581 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11586) );
  OAI21_X1 U14582 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n11586), .ZN(n20393) );
  NAND2_X1 U14583 ( .A1(n20634), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11593) );
  OAI21_X1 U14584 ( .B1(n13464), .B2(n20393), .A(n11593), .ZN(n11540) );
  INV_X1 U14585 ( .A(n11540), .ZN(n11541) );
  NAND2_X1 U14586 ( .A1(n11542), .A2(n11541), .ZN(n11544) );
  XNOR2_X2 U14587 ( .A(n11544), .B(n11592), .ZN(n20176) );
  NAND2_X1 U14588 ( .A1(n20176), .A2(n11598), .ZN(n11597) );
  INV_X1 U14589 ( .A(n20176), .ZN(n11548) );
  INV_X1 U14590 ( .A(n11637), .ZN(n11561) );
  AOI22_X1 U14591 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11552) );
  AOI22_X1 U14592 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12435), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U14593 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11550) );
  AOI22_X1 U14594 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11549) );
  NAND4_X1 U14595 ( .A1(n11552), .A2(n11551), .A3(n11550), .A4(n11549), .ZN(
        n11560) );
  AOI22_X1 U14596 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11558) );
  AOI22_X1 U14597 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12479), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U14598 ( .A1(n11518), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U14599 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12478), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11555) );
  NAND4_X1 U14600 ( .A1(n11558), .A2(n11557), .A3(n11556), .A4(n11555), .ZN(
        n11559) );
  NAND2_X1 U14601 ( .A1(n12004), .A2(n20076), .ZN(n11567) );
  XNOR2_X1 U14602 ( .A(n11620), .B(n11619), .ZN(n11564) );
  OAI211_X1 U14603 ( .C1(n11564), .C2(n11496), .A(n9842), .B(n20093), .ZN(
        n11565) );
  INV_X1 U14604 ( .A(n11565), .ZN(n11566) );
  NAND2_X1 U14605 ( .A1(n11567), .A2(n11566), .ZN(n11568) );
  NAND2_X1 U14606 ( .A1(n13689), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11571) );
  INV_X1 U14607 ( .A(n11568), .ZN(n11569) );
  OR2_X1 U14608 ( .A1(n13461), .A2(n11569), .ZN(n11570) );
  NAND2_X1 U14609 ( .A1(n11571), .A2(n11570), .ZN(n11628) );
  INV_X1 U14610 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13554) );
  NAND2_X1 U14611 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11578) );
  INV_X1 U14612 ( .A(n11574), .ZN(n11577) );
  NAND2_X1 U14613 ( .A1(n11575), .A2(n11620), .ZN(n11576) );
  NAND2_X1 U14614 ( .A1(n12005), .A2(n12004), .ZN(n11583) );
  INV_X1 U14615 ( .A(n11579), .ZN(n11580) );
  INV_X1 U14616 ( .A(n11586), .ZN(n11585) );
  NAND2_X1 U14617 ( .A1(n11585), .A2(n11803), .ZN(n20424) );
  NAND2_X1 U14618 ( .A1(n11586), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11587) );
  NAND2_X1 U14619 ( .A1(n20634), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11588) );
  INV_X1 U14620 ( .A(n11592), .ZN(n11595) );
  NAND2_X1 U14621 ( .A1(n11593), .A2(n11792), .ZN(n11594) );
  NOR2_X1 U14622 ( .A1(n11599), .A2(n9639), .ZN(n11596) );
  NAND2_X1 U14623 ( .A1(n11597), .A2(n11596), .ZN(n11602) );
  NAND3_X1 U14624 ( .A1(n20176), .A2(n11599), .A3(n11598), .ZN(n11601) );
  NAND2_X1 U14625 ( .A1(n11599), .A2(n9639), .ZN(n11600) );
  NAND2_X1 U14626 ( .A1(n11602), .A2(n11631), .ZN(n13475) );
  AOI22_X1 U14627 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11606) );
  AOI22_X1 U14628 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U14629 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14630 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12478), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11603) );
  NAND4_X1 U14631 ( .A1(n11606), .A2(n11605), .A3(n11604), .A4(n11603), .ZN(
        n11612) );
  AOI22_X1 U14632 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U14633 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U14634 ( .A1(n11518), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11608) );
  AOI22_X1 U14635 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11607) );
  NAND4_X1 U14636 ( .A1(n11610), .A2(n11609), .A3(n11608), .A4(n11607), .ZN(
        n11611) );
  NOR2_X1 U14637 ( .A1(n11612), .A2(n11611), .ZN(n11622) );
  INV_X1 U14638 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11613) );
  OAI22_X1 U14639 ( .A1(n11814), .A2(n11613), .B1(n11622), .B2(n11638), .ZN(
        n11614) );
  OR2_X1 U14640 ( .A1(n11999), .A2(n11813), .ZN(n11627) );
  NAND2_X1 U14641 ( .A1(n11620), .A2(n11619), .ZN(n11621) );
  NAND2_X1 U14642 ( .A1(n11621), .A2(n11622), .ZN(n11673) );
  OAI21_X1 U14643 ( .B1(n11622), .B2(n11621), .A(n11673), .ZN(n11625) );
  INV_X1 U14644 ( .A(n11496), .ZN(n20743) );
  INV_X1 U14645 ( .A(n11623), .ZN(n11624) );
  AOI21_X1 U14646 ( .B1(n11625), .B2(n20743), .A(n11624), .ZN(n11626) );
  NAND2_X1 U14647 ( .A1(n11627), .A2(n11626), .ZN(n13544) );
  NAND2_X1 U14648 ( .A1(n13545), .A2(n13544), .ZN(n11630) );
  NAND2_X1 U14649 ( .A1(n11632), .A2(n20708), .ZN(n11636) );
  INV_X1 U14650 ( .A(n13464), .ZN(n11634) );
  NAND3_X1 U14651 ( .A1(n20727), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20303) );
  INV_X1 U14652 ( .A(n20324), .ZN(n11633) );
  NAND3_X1 U14653 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20579) );
  AOI21_X1 U14654 ( .B1(n20727), .B2(n11633), .A(n20625), .ZN(n20333) );
  AOI22_X1 U14655 ( .A1(n11634), .A2(n20333), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20634), .ZN(n11635) );
  XNOR2_X2 U14656 ( .A(n13470), .B(n20212), .ZN(n20717) );
  AOI22_X1 U14657 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11642) );
  AOI22_X1 U14658 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12381), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11641) );
  AOI22_X1 U14659 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12479), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11640) );
  AOI22_X1 U14660 ( .A1(n11518), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11639) );
  NAND4_X1 U14661 ( .A1(n11642), .A2(n11641), .A3(n11640), .A4(n11639), .ZN(
        n11648) );
  AOI22_X1 U14662 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14663 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14664 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14665 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12478), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11643) );
  NAND4_X1 U14666 ( .A1(n11646), .A2(n11645), .A3(n11644), .A4(n11643), .ZN(
        n11647) );
  AOI22_X1 U14667 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11837), .B2(n11672), .ZN(n11649) );
  INV_X1 U14668 ( .A(n20211), .ZN(n20058) );
  NAND2_X1 U14669 ( .A1(n11651), .A2(n20058), .ZN(n11652) );
  NAND2_X1 U14670 ( .A1(n11670), .A2(n11652), .ZN(n20056) );
  INV_X1 U14671 ( .A(n11672), .ZN(n11653) );
  XNOR2_X1 U14672 ( .A(n11673), .B(n11653), .ZN(n11654) );
  NAND2_X1 U14673 ( .A1(n11654), .A2(n20743), .ZN(n11655) );
  OAI21_X1 U14674 ( .B1(n20056), .B2(n11813), .A(n11655), .ZN(n11656) );
  INV_X1 U14675 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11880) );
  XNOR2_X1 U14676 ( .A(n11656), .B(n11880), .ZN(n13703) );
  NAND2_X1 U14677 ( .A1(n11656), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11657) );
  AOI22_X1 U14678 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11661) );
  INV_X1 U14679 ( .A(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n20862) );
  AOI22_X1 U14680 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U14681 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14682 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12478), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11658) );
  NAND4_X1 U14683 ( .A1(n11661), .A2(n11660), .A3(n11659), .A4(n11658), .ZN(
        n11667) );
  AOI22_X1 U14684 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11665) );
  AOI22_X1 U14685 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11664) );
  AOI22_X1 U14686 ( .A1(n11518), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11663) );
  AOI22_X1 U14687 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11662) );
  NAND4_X1 U14688 ( .A1(n11665), .A2(n11664), .A3(n11663), .A4(n11662), .ZN(
        n11666) );
  AOI22_X1 U14689 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11837), .B2(n11676), .ZN(n11669) );
  NAND2_X1 U14690 ( .A1(n11670), .A2(n11669), .ZN(n11671) );
  AND2_X1 U14691 ( .A1(n11703), .A2(n11671), .ZN(n12043) );
  INV_X1 U14692 ( .A(n11813), .ZN(n11741) );
  NAND2_X1 U14693 ( .A1(n12043), .A2(n11741), .ZN(n11679) );
  NAND2_X1 U14694 ( .A1(n11673), .A2(n11672), .ZN(n11675) );
  INV_X1 U14695 ( .A(n11675), .ZN(n11677) );
  INV_X1 U14696 ( .A(n11676), .ZN(n11674) );
  NOR2_X1 U14697 ( .A1(n11675), .A2(n11674), .ZN(n11722) );
  INV_X1 U14698 ( .A(n11722), .ZN(n11696) );
  OAI211_X1 U14699 ( .C1(n11677), .C2(n11676), .A(n20743), .B(n11696), .ZN(
        n11678) );
  NAND2_X1 U14700 ( .A1(n11679), .A2(n11678), .ZN(n11681) );
  INV_X1 U14701 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11680) );
  XNOR2_X1 U14702 ( .A(n11681), .B(n11680), .ZN(n13767) );
  NAND2_X1 U14703 ( .A1(n11681), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11682) );
  NAND2_X1 U14704 ( .A1(n11683), .A2(n11682), .ZN(n13792) );
  INV_X1 U14705 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14706 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U14707 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11686) );
  AOI22_X1 U14708 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11685) );
  AOI22_X1 U14709 ( .A1(n11518), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11684) );
  NAND4_X1 U14710 ( .A1(n11687), .A2(n11686), .A3(n11685), .A4(n11684), .ZN(
        n11693) );
  AOI22_X1 U14711 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11691) );
  AOI22_X1 U14712 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U14713 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U14714 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12478), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11688) );
  NAND4_X1 U14715 ( .A1(n11691), .A2(n11690), .A3(n11689), .A4(n11688), .ZN(
        n11692) );
  NAND2_X1 U14716 ( .A1(n11837), .A2(n11721), .ZN(n11694) );
  OAI21_X1 U14717 ( .B1(n11814), .B2(n11695), .A(n11694), .ZN(n11704) );
  XNOR2_X1 U14718 ( .A(n11703), .B(n11704), .ZN(n12044) );
  NAND2_X1 U14719 ( .A1(n12044), .A2(n11741), .ZN(n11699) );
  XNOR2_X1 U14720 ( .A(n11696), .B(n11721), .ZN(n11697) );
  NAND2_X1 U14721 ( .A1(n11697), .A2(n20743), .ZN(n11698) );
  NAND2_X1 U14722 ( .A1(n11699), .A2(n11698), .ZN(n11700) );
  INV_X1 U14723 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n20852) );
  XNOR2_X1 U14724 ( .A(n11700), .B(n20852), .ZN(n13793) );
  NAND2_X1 U14725 ( .A1(n13792), .A2(n13793), .ZN(n11702) );
  NAND2_X1 U14726 ( .A1(n11700), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11701) );
  INV_X1 U14727 ( .A(n11703), .ZN(n11705) );
  NAND2_X1 U14728 ( .A1(n11705), .A2(n11704), .ZN(n11720) );
  INV_X1 U14729 ( .A(n11720), .ZN(n11718) );
  AOI22_X1 U14730 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U14731 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U14732 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11707) );
  AOI22_X1 U14733 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12478), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11706) );
  NAND4_X1 U14734 ( .A1(n11709), .A2(n11708), .A3(n11707), .A4(n11706), .ZN(
        n11716) );
  AOI22_X1 U14735 ( .A1(n11710), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U14736 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U14737 ( .A1(n11518), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U14738 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11711) );
  NAND4_X1 U14739 ( .A1(n11714), .A2(n11713), .A3(n11712), .A4(n11711), .ZN(
        n11715) );
  AOI22_X1 U14740 ( .A1(n11847), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11837), .B2(n11732), .ZN(n11719) );
  INV_X1 U14741 ( .A(n11719), .ZN(n11717) );
  NAND2_X1 U14742 ( .A1(n11718), .A2(n11717), .ZN(n11731) );
  NAND2_X1 U14743 ( .A1(n11720), .A2(n11719), .ZN(n12057) );
  NAND2_X1 U14744 ( .A1(n11722), .A2(n11721), .ZN(n11733) );
  XNOR2_X1 U14745 ( .A(n11733), .B(n11732), .ZN(n11723) );
  NAND2_X1 U14746 ( .A1(n11723), .A2(n20743), .ZN(n11724) );
  NAND2_X1 U14747 ( .A1(n11725), .A2(n11724), .ZN(n11726) );
  INV_X1 U14748 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16142) );
  XNOR2_X1 U14749 ( .A(n11726), .B(n16142), .ZN(n14140) );
  NAND2_X1 U14750 ( .A1(n11726), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11727) );
  INV_X1 U14751 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11729) );
  NAND2_X1 U14752 ( .A1(n11837), .A2(n11745), .ZN(n11728) );
  OAI21_X1 U14753 ( .B1(n11814), .B2(n11729), .A(n11728), .ZN(n11730) );
  NAND2_X1 U14754 ( .A1(n12064), .A2(n11741), .ZN(n11738) );
  INV_X1 U14755 ( .A(n11732), .ZN(n11734) );
  NOR2_X1 U14756 ( .A1(n11734), .A2(n11733), .ZN(n11744) );
  INV_X1 U14757 ( .A(n11744), .ZN(n11735) );
  XNOR2_X1 U14758 ( .A(n11745), .B(n11735), .ZN(n11736) );
  NAND2_X1 U14759 ( .A1(n20743), .A2(n11736), .ZN(n11737) );
  NAND2_X1 U14760 ( .A1(n11738), .A2(n11737), .ZN(n11739) );
  OR2_X1 U14761 ( .A1(n11739), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16063) );
  NAND2_X1 U14762 ( .A1(n11739), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16062) );
  NAND2_X1 U14763 ( .A1(n11740), .A2(n16062), .ZN(n14146) );
  AND2_X1 U14764 ( .A1(n11742), .A2(n11741), .ZN(n11743) );
  INV_X4 U14765 ( .A(n15941), .ZN(n15131) );
  NAND2_X1 U14766 ( .A1(n11745), .A2(n11744), .ZN(n11746) );
  OR2_X1 U14767 ( .A1(n11496), .A2(n11746), .ZN(n11747) );
  NAND2_X1 U14768 ( .A1(n15131), .A2(n11747), .ZN(n14147) );
  OR2_X1 U14769 ( .A1(n14147), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11748) );
  NAND2_X1 U14770 ( .A1(n14146), .A2(n11748), .ZN(n11750) );
  NAND2_X1 U14771 ( .A1(n14147), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11749) );
  INV_X1 U14772 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11751) );
  NAND2_X1 U14773 ( .A1(n15131), .A2(n11751), .ZN(n11752) );
  INV_X1 U14774 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16089) );
  NAND2_X1 U14775 ( .A1(n15131), .A2(n16089), .ZN(n11754) );
  NAND2_X1 U14776 ( .A1(n14981), .A2(n11754), .ZN(n16049) );
  INV_X1 U14777 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11762) );
  NAND2_X1 U14778 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11755) );
  INV_X1 U14779 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11757) );
  NAND2_X1 U14780 ( .A1(n15131), .A2(n11757), .ZN(n11756) );
  OR2_X1 U14781 ( .A1(n11753), .A2(n11757), .ZN(n11758) );
  INV_X1 U14782 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11917) );
  XNOR2_X1 U14783 ( .A(n15136), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14970) );
  NAND2_X1 U14784 ( .A1(n15131), .A2(n11917), .ZN(n16036) );
  NAND2_X1 U14785 ( .A1(n14970), .A2(n16036), .ZN(n11759) );
  OAI21_X1 U14786 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n15941), .A(
        n15132), .ZN(n11766) );
  NOR2_X1 U14787 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11761) );
  OR2_X1 U14788 ( .A1(n15136), .A2(n11761), .ZN(n14993) );
  OR2_X1 U14789 ( .A1(n15136), .A2(n11762), .ZN(n14991) );
  NAND2_X1 U14790 ( .A1(n14993), .A2(n14991), .ZN(n14980) );
  NOR2_X1 U14791 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11763) );
  NOR2_X1 U14792 ( .A1(n15131), .A2(n11763), .ZN(n11764) );
  XNOR2_X1 U14793 ( .A(n15136), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14961) );
  INV_X1 U14794 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15104) );
  INV_X1 U14795 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15113) );
  INV_X1 U14796 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11937) );
  NOR2_X1 U14797 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14950) );
  NAND3_X1 U14798 ( .A1(n14950), .A2(n15104), .A3(n11937), .ZN(n11767) );
  NAND2_X1 U14799 ( .A1(n11768), .A2(n15941), .ZN(n14942) );
  AND2_X2 U14800 ( .A1(n11769), .A2(n14942), .ZN(n14932) );
  NOR3_X1 U14801 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14879) );
  NAND2_X1 U14802 ( .A1(n14932), .A2(n14879), .ZN(n14906) );
  INV_X1 U14803 ( .A(n11771), .ZN(n11770) );
  NOR2_X1 U14804 ( .A1(n14906), .A2(n11770), .ZN(n14891) );
  NOR2_X1 U14805 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15030) );
  NAND2_X1 U14806 ( .A1(n14891), .A2(n15030), .ZN(n14517) );
  AND2_X1 U14807 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11984) );
  NAND2_X1 U14808 ( .A1(n11984), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14878) );
  NOR2_X2 U14809 ( .A1(n11771), .A2(n14878), .ZN(n14890) );
  NAND2_X1 U14810 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15032) );
  INV_X1 U14811 ( .A(n15032), .ZN(n11772) );
  AND2_X2 U14812 ( .A1(n14890), .A2(n11772), .ZN(n11776) );
  AOI21_X2 U14813 ( .B1(n14517), .B2(n15941), .A(n11776), .ZN(n14872) );
  INV_X1 U14814 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15010) );
  INV_X1 U14815 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15020) );
  NAND2_X1 U14816 ( .A1(n15010), .A2(n15020), .ZN(n11773) );
  NOR2_X1 U14817 ( .A1(n11773), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11774) );
  NAND2_X1 U14818 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11777) );
  NOR2_X1 U14819 ( .A1(n11777), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11997) );
  MUX2_X1 U14820 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11997), .S(
        n15131), .Z(n11779) );
  AOI22_X1 U14821 ( .A1(n14872), .A2(n11774), .B1(n11779), .B2(n11773), .ZN(
        n11775) );
  INV_X1 U14822 ( .A(n11776), .ZN(n14518) );
  OAI21_X1 U14823 ( .B1(n14518), .B2(n11777), .A(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11778) );
  INV_X1 U14824 ( .A(n11779), .ZN(n11780) );
  NOR2_X1 U14825 ( .A1(n11482), .A2(n20076), .ZN(n11782) );
  OAI21_X1 U14826 ( .B1(n11783), .B2(n11782), .A(n20061), .ZN(n11977) );
  NAND2_X1 U14827 ( .A1(n11787), .A2(n14092), .ZN(n11859) );
  NAND3_X1 U14828 ( .A1(n11977), .A2(n11785), .A3(n11859), .ZN(n11790) );
  NAND2_X1 U14829 ( .A1(n11790), .A2(n11789), .ZN(n13453) );
  NAND2_X1 U14830 ( .A1(n11791), .A2(n20650), .ZN(n15956) );
  INV_X1 U14831 ( .A(n15956), .ZN(n13418) );
  MUX2_X1 U14832 ( .A(n20386), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11810) );
  NAND2_X1 U14833 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20499), .ZN(
        n11819) );
  NAND2_X1 U14834 ( .A1(n11810), .A2(n11809), .ZN(n11808) );
  INV_X1 U14835 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11792) );
  INV_X1 U14836 ( .A(n11792), .ZN(n13648) );
  NAND2_X1 U14837 ( .A1(n13648), .A2(n20386), .ZN(n11793) );
  NAND2_X1 U14838 ( .A1(n11808), .A2(n11793), .ZN(n11805) );
  NAND2_X1 U14839 ( .A1(n11805), .A2(n11794), .ZN(n11796) );
  NAND2_X1 U14840 ( .A1(n11803), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11795) );
  XNOR2_X1 U14841 ( .A(n20708), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11806) );
  NOR2_X1 U14842 ( .A1(n11321), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11797) );
  INV_X1 U14843 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n11798) );
  NAND2_X1 U14844 ( .A1(n11798), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11800) );
  NOR2_X1 U14845 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n11798), .ZN(
        n11799) );
  INV_X1 U14846 ( .A(n11801), .ZN(n11802) );
  MUX2_X1 U14847 ( .A(n11803), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11804) );
  XNOR2_X1 U14848 ( .A(n11805), .B(n11804), .ZN(n11835) );
  XNOR2_X1 U14849 ( .A(n11807), .B(n11806), .ZN(n11840) );
  OAI21_X1 U14850 ( .B1(n11810), .B2(n11809), .A(n11808), .ZN(n11829) );
  NOR4_X1 U14851 ( .A1(n11818), .A2(n11835), .A3(n11840), .A4(n11829), .ZN(
        n11811) );
  OR2_X1 U14852 ( .A1(n11815), .A2(n11811), .ZN(n13285) );
  NAND2_X1 U14853 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20647) );
  INV_X1 U14854 ( .A(n20647), .ZN(n20741) );
  INV_X1 U14855 ( .A(n12513), .ZN(n11812) );
  OAI211_X1 U14856 ( .C1(n15926), .C2(n13418), .A(n11812), .B(n11477), .ZN(
        n11853) );
  NAND2_X1 U14857 ( .A1(n11841), .A2(n11815), .ZN(n11851) );
  NAND2_X1 U14858 ( .A1(n11815), .A2(n11837), .ZN(n11850) );
  NAND2_X1 U14859 ( .A1(n11824), .A2(n11816), .ZN(n11827) );
  INV_X1 U14860 ( .A(n11827), .ZN(n11817) );
  NAND2_X1 U14861 ( .A1(n11817), .A2(n20076), .ZN(n11849) );
  INV_X1 U14862 ( .A(n11818), .ZN(n11846) );
  OAI21_X1 U14863 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20499), .A(
        n11819), .ZN(n11823) );
  INV_X1 U14864 ( .A(n11823), .ZN(n11820) );
  OAI21_X1 U14865 ( .B1(n11968), .B2(n11821), .A(n11820), .ZN(n11826) );
  NAND2_X1 U14866 ( .A1(n15926), .A2(n20093), .ZN(n11828) );
  NAND2_X1 U14867 ( .A1(n14111), .A2(n11828), .ZN(n11836) );
  INV_X1 U14868 ( .A(n11841), .ZN(n11822) );
  OAI21_X1 U14869 ( .B1(n11824), .B2(n11823), .A(n11822), .ZN(n11825) );
  INV_X1 U14870 ( .A(n11830), .ZN(n11833) );
  INV_X1 U14871 ( .A(n11831), .ZN(n11832) );
  INV_X1 U14872 ( .A(n11835), .ZN(n11839) );
  AOI21_X1 U14873 ( .B1(n11839), .B2(n11837), .A(n11836), .ZN(n11834) );
  NOR2_X1 U14874 ( .A1(n11834), .A2(n11840), .ZN(n11838) );
  AOI21_X1 U14875 ( .B1(n11847), .B2(n11835), .A(n11838), .ZN(n11844) );
  NAND4_X1 U14876 ( .A1(n11839), .A2(n11838), .A3(n11837), .A4(n11836), .ZN(
        n11843) );
  NAND2_X1 U14877 ( .A1(n11841), .A2(n11840), .ZN(n11842) );
  OAI21_X1 U14878 ( .B1(n11847), .B2(n11846), .A(n11845), .ZN(n11848) );
  OR3_X1 U14879 ( .A1(n11787), .A2(n13444), .A3(n15926), .ZN(n11852) );
  NAND2_X1 U14880 ( .A1(n15926), .A2(n15956), .ZN(n14094) );
  NAND2_X1 U14881 ( .A1(n14094), .A2(n20647), .ZN(n11856) );
  OAI211_X1 U14882 ( .C1(n11855), .C2(n11856), .A(n20061), .B(n11472), .ZN(
        n11857) );
  INV_X1 U14883 ( .A(n11968), .ZN(n11858) );
  AND2_X1 U14884 ( .A1(n11859), .A2(n11858), .ZN(n11860) );
  AND2_X1 U14885 ( .A1(n11785), .A2(n11860), .ZN(n15920) );
  NOR2_X1 U14886 ( .A1(n14111), .A2(n11480), .ZN(n11861) );
  NAND2_X1 U14887 ( .A1(n13478), .A2(n11861), .ZN(n13286) );
  OAI21_X1 U14888 ( .B1(n11867), .B2(n12464), .A(n13286), .ZN(n11862) );
  NOR2_X1 U14889 ( .A1(n15920), .A2(n11862), .ZN(n11863) );
  AND2_X1 U14890 ( .A1(n11864), .A2(n11863), .ZN(n11865) );
  NOR2_X1 U14891 ( .A1(n11867), .A2(n11483), .ZN(n11868) );
  AOI21_X1 U14892 ( .B1(n15927), .B2(n15926), .A(n11868), .ZN(n11869) );
  NAND2_X1 U14893 ( .A1(n13404), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n11871) );
  NAND2_X1 U14894 ( .A1(n11914), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11870) );
  AND2_X1 U14895 ( .A1(n11871), .A2(n11870), .ZN(n12504) );
  INV_X1 U14896 ( .A(n11894), .ZN(n11875) );
  INV_X1 U14897 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n11872) );
  OR2_X1 U14898 ( .A1(n11879), .A2(n11872), .ZN(n11874) );
  INV_X1 U14899 ( .A(n11938), .ZN(n13281) );
  NAND2_X1 U14900 ( .A1(n13281), .A2(n11872), .ZN(n11873) );
  NAND2_X1 U14901 ( .A1(n11874), .A2(n11873), .ZN(n13403) );
  OR2_X1 U14902 ( .A1(n13404), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11878) );
  INV_X1 U14903 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n11876) );
  MUX2_X1 U14904 ( .A(n11960), .B(n11956), .S(n11876), .Z(n11877) );
  AND2_X1 U14905 ( .A1(n11878), .A2(n11877), .ZN(n13548) );
  AND2_X1 U14906 ( .A1(n13549), .A2(n13548), .ZN(n13708) );
  NAND2_X1 U14907 ( .A1(n11499), .A2(n11880), .ZN(n11881) );
  OAI211_X1 U14908 ( .C1(n11914), .C2(P1_EBX_REG_3__SCAN_IN), .A(n11881), .B(
        n11960), .ZN(n11882) );
  OAI21_X1 U14909 ( .B1(P1_EBX_REG_3__SCAN_IN), .B2(n11959), .A(n11882), .ZN(
        n13707) );
  NAND2_X1 U14910 ( .A1(n13708), .A2(n13707), .ZN(n13772) );
  OR2_X1 U14911 ( .A1(n11956), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n11885) );
  NAND2_X1 U14912 ( .A1(n11960), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11883) );
  OAI211_X1 U14913 ( .C1(n11914), .C2(P1_EBX_REG_4__SCAN_IN), .A(n11499), .B(
        n11883), .ZN(n11884) );
  NAND2_X1 U14914 ( .A1(n11885), .A2(n11884), .ZN(n13771) );
  OR2_X1 U14915 ( .A1(n11956), .A2(P1_EBX_REG_6__SCAN_IN), .ZN(n11888) );
  NAND2_X1 U14916 ( .A1(n11960), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11886) );
  OAI211_X1 U14917 ( .C1(n11914), .C2(P1_EBX_REG_6__SCAN_IN), .A(n11499), .B(
        n11886), .ZN(n11887) );
  AND2_X1 U14918 ( .A1(n11888), .A2(n11887), .ZN(n16129) );
  NAND2_X1 U14919 ( .A1(n11960), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11889) );
  NAND2_X1 U14920 ( .A1(n11499), .A2(n11889), .ZN(n11891) );
  OR2_X1 U14921 ( .A1(n11914), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n11890) );
  NAND2_X1 U14922 ( .A1(n11891), .A2(n11890), .ZN(n11892) );
  OAI21_X1 U14923 ( .B1(n11959), .B2(P1_EBX_REG_5__SCAN_IN), .A(n11892), .ZN(
        n16130) );
  NAND2_X1 U14924 ( .A1(n16129), .A2(n16130), .ZN(n11893) );
  OR2_X1 U14925 ( .A1(n11956), .A2(P1_EBX_REG_8__SCAN_IN), .ZN(n11897) );
  NAND2_X1 U14926 ( .A1(n11960), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11895) );
  OAI211_X1 U14927 ( .C1(n11914), .C2(P1_EBX_REG_8__SCAN_IN), .A(n11499), .B(
        n11895), .ZN(n11896) );
  AND2_X1 U14928 ( .A1(n11897), .A2(n11896), .ZN(n14158) );
  NAND2_X1 U14929 ( .A1(n11960), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11898) );
  NAND2_X1 U14930 ( .A1(n11499), .A2(n11898), .ZN(n11900) );
  OR2_X1 U14931 ( .A1(n11914), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n11899) );
  NAND2_X1 U14932 ( .A1(n11900), .A2(n11899), .ZN(n11901) );
  OAI21_X1 U14933 ( .B1(n11959), .B2(P1_EBX_REG_7__SCAN_IN), .A(n11901), .ZN(
        n14167) );
  AND2_X1 U14934 ( .A1(n14158), .A2(n14167), .ZN(n11902) );
  NAND2_X1 U14935 ( .A1(n11960), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11903) );
  NAND2_X1 U14936 ( .A1(n11499), .A2(n11903), .ZN(n11905) );
  OR2_X1 U14937 ( .A1(n11914), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n11904) );
  NAND2_X1 U14938 ( .A1(n11905), .A2(n11904), .ZN(n11906) );
  OAI21_X1 U14939 ( .B1(n11959), .B2(P1_EBX_REG_9__SCAN_IN), .A(n11906), .ZN(
        n14214) );
  MUX2_X1 U14940 ( .A(n11956), .B(n11960), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n11907) );
  OAI21_X1 U14941 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n13404), .A(
        n11907), .ZN(n14336) );
  MUX2_X1 U14942 ( .A(n11956), .B(n11960), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n11909) );
  OR2_X1 U14943 ( .A1(n13404), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11908) );
  AND2_X1 U14944 ( .A1(n11909), .A2(n11908), .ZN(n14739) );
  INV_X1 U14945 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n20800) );
  NAND2_X1 U14946 ( .A1(n11499), .A2(n20800), .ZN(n11911) );
  OR2_X1 U14947 ( .A1(n11914), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n11910) );
  NAND3_X1 U14948 ( .A1(n11911), .A2(n11910), .A3(n11960), .ZN(n11912) );
  OAI21_X1 U14949 ( .B1(n11959), .B2(P1_EBX_REG_11__SCAN_IN), .A(n11912), .ZN(
        n14740) );
  NAND2_X1 U14950 ( .A1(n11499), .A2(n16089), .ZN(n11913) );
  OAI211_X1 U14951 ( .C1(n11914), .C2(P1_EBX_REG_13__SCAN_IN), .A(n11913), .B(
        n11960), .ZN(n11915) );
  OAI21_X1 U14952 ( .B1(P1_EBX_REG_13__SCAN_IN), .B2(n11959), .A(n11915), .ZN(
        n14788) );
  MUX2_X1 U14953 ( .A(n11956), .B(n11938), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n11916) );
  OAI21_X1 U14954 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n13404), .A(
        n11916), .ZN(n14726) );
  INV_X1 U14955 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14782) );
  NAND2_X1 U14956 ( .A1(n11946), .A2(n14782), .ZN(n11920) );
  NAND2_X1 U14957 ( .A1(n11499), .A2(n11917), .ZN(n11918) );
  OAI211_X1 U14958 ( .C1(n11914), .C2(P1_EBX_REG_15__SCAN_IN), .A(n11918), .B(
        n11960), .ZN(n11919) );
  MUX2_X1 U14959 ( .A(n11956), .B(n11960), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n11922) );
  OR2_X1 U14960 ( .A1(n13404), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11921) );
  NAND2_X1 U14961 ( .A1(n11922), .A2(n11921), .ZN(n14713) );
  INV_X1 U14962 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11923) );
  NAND2_X1 U14963 ( .A1(n11499), .A2(n11923), .ZN(n11924) );
  OAI211_X1 U14964 ( .C1(n11914), .C2(P1_EBX_REG_17__SCAN_IN), .A(n11924), .B(
        n11960), .ZN(n11925) );
  OAI21_X1 U14965 ( .B1(P1_EBX_REG_17__SCAN_IN), .B2(n11959), .A(n11925), .ZN(
        n14697) );
  OR2_X1 U14966 ( .A1(n11956), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n11928) );
  NAND2_X1 U14967 ( .A1(n11960), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11926) );
  OAI211_X1 U14968 ( .C1(n11914), .C2(P1_EBX_REG_18__SCAN_IN), .A(n11499), .B(
        n11926), .ZN(n11927) );
  INV_X1 U14969 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14770) );
  NAND2_X1 U14970 ( .A1(n11946), .A2(n14770), .ZN(n11931) );
  NAND2_X1 U14971 ( .A1(n11499), .A2(n15113), .ZN(n11929) );
  OAI211_X1 U14972 ( .C1(n11914), .C2(P1_EBX_REG_19__SCAN_IN), .A(n11929), .B(
        n11938), .ZN(n11930) );
  OR2_X1 U14973 ( .A1(n11956), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n11934) );
  NAND2_X1 U14974 ( .A1(n11960), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11932) );
  OAI211_X1 U14975 ( .C1(n11914), .C2(P1_EBX_REG_20__SCAN_IN), .A(n11499), .B(
        n11932), .ZN(n11933) );
  NAND2_X1 U14976 ( .A1(n11934), .A2(n11933), .ZN(n14661) );
  MUX2_X1 U14977 ( .A(n11956), .B(n11960), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n11936) );
  OR2_X1 U14978 ( .A1(n13404), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11935) );
  NAND2_X1 U14979 ( .A1(n11936), .A2(n11935), .ZN(n14647) );
  INV_X1 U14980 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n16016) );
  NAND2_X1 U14981 ( .A1(n11946), .A2(n16016), .ZN(n11941) );
  NAND2_X1 U14982 ( .A1(n11499), .A2(n11937), .ZN(n11939) );
  OAI211_X1 U14983 ( .C1(n11914), .C2(P1_EBX_REG_21__SCAN_IN), .A(n11939), .B(
        n11938), .ZN(n11940) );
  INV_X1 U14984 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15077) );
  NAND2_X1 U14985 ( .A1(n11499), .A2(n15077), .ZN(n11942) );
  OAI211_X1 U14986 ( .C1(n11914), .C2(P1_EBX_REG_23__SCAN_IN), .A(n11942), .B(
        n11960), .ZN(n11943) );
  OAI21_X1 U14987 ( .B1(P1_EBX_REG_23__SCAN_IN), .B2(n11959), .A(n11943), .ZN(
        n14637) );
  MUX2_X1 U14988 ( .A(n11956), .B(n11960), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n11945) );
  OR2_X1 U14989 ( .A1(n13404), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11944) );
  NAND2_X1 U14990 ( .A1(n11945), .A2(n11944), .ZN(n14627) );
  INV_X1 U14991 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14762) );
  NAND2_X1 U14992 ( .A1(n11946), .A2(n14762), .ZN(n11949) );
  INV_X1 U14993 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15060) );
  NAND2_X1 U14994 ( .A1(n11499), .A2(n15060), .ZN(n11947) );
  OAI211_X1 U14995 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n11914), .A(n11947), .B(
        n11960), .ZN(n11948) );
  AND2_X1 U14996 ( .A1(n11949), .A2(n11948), .ZN(n14614) );
  MUX2_X1 U14997 ( .A(n11956), .B(n11960), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n11951) );
  OR2_X1 U14998 ( .A1(n13404), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11950) );
  NAND2_X1 U14999 ( .A1(n11951), .A2(n11950), .ZN(n14602) );
  NAND2_X1 U15000 ( .A1(n11960), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11952) );
  NAND2_X1 U15001 ( .A1(n11499), .A2(n11952), .ZN(n11954) );
  OR2_X1 U15002 ( .A1(n11914), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n11953) );
  NAND2_X1 U15003 ( .A1(n11954), .A2(n11953), .ZN(n11955) );
  OAI21_X1 U15004 ( .B1(n11959), .B2(P1_EBX_REG_27__SCAN_IN), .A(n11955), .ZN(
        n14589) );
  MUX2_X1 U15005 ( .A(n11956), .B(n11960), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n11958) );
  OR2_X1 U15006 ( .A1(n13404), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11957) );
  AND2_X1 U15007 ( .A1(n11958), .A2(n11957), .ZN(n14574) );
  OAI22_X1 U15008 ( .A1(n13404), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        P1_EBX_REG_29__SCAN_IN), .B2(n11914), .ZN(n12502) );
  OAI22_X1 U15009 ( .A1(n12502), .A2(n13281), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n11959), .ZN(n12468) );
  MUX2_X1 U15010 ( .A(n12504), .B(n11960), .S(n9657), .Z(n11963) );
  NOR2_X1 U15011 ( .A1(n9657), .A2(n12504), .ZN(n11962) );
  AOI22_X1 U15012 ( .A1(n13404), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n11914), .ZN(n11961) );
  MUX2_X1 U15013 ( .A(n11963), .B(n11962), .S(n11961), .Z(n14514) );
  NAND2_X1 U15014 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15088) );
  NAND4_X1 U15015 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15123) );
  INV_X1 U15016 ( .A(n15123), .ZN(n15122) );
  NAND2_X1 U15017 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15122), .ZN(
        n11988) );
  INV_X1 U15018 ( .A(n11988), .ZN(n11989) );
  OR2_X1 U15019 ( .A1(n11789), .A2(n15926), .ZN(n13643) );
  NOR2_X1 U15020 ( .A1(n13554), .A2(n9866), .ZN(n13796) );
  NOR2_X1 U15021 ( .A1(n11680), .A2(n11880), .ZN(n13797) );
  NAND2_X1 U15022 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13797), .ZN(
        n11965) );
  INV_X1 U15023 ( .A(n11965), .ZN(n14153) );
  NAND2_X1 U15024 ( .A1(n13796), .A2(n14153), .ZN(n16095) );
  INV_X1 U15025 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14155) );
  INV_X1 U15026 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n14154) );
  NOR3_X1 U15027 ( .A1(n14155), .A2(n14154), .A3(n16142), .ZN(n14213) );
  NAND3_X1 U15028 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n14213), .ZN(n16094) );
  NOR2_X1 U15029 ( .A1(n20800), .A2(n16094), .ZN(n16105) );
  NAND2_X1 U15030 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16105), .ZN(
        n11966) );
  NOR2_X1 U15031 ( .A1(n16095), .A2(n11966), .ZN(n11983) );
  NOR2_X1 U15032 ( .A1(n11480), .A2(n11914), .ZN(n11964) );
  NAND2_X1 U15033 ( .A1(n13478), .A2(n11964), .ZN(n13290) );
  AOI21_X1 U15034 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13706) );
  NOR2_X1 U15035 ( .A1(n13706), .A2(n11965), .ZN(n14212) );
  INV_X1 U15036 ( .A(n14212), .ZN(n13795) );
  NOR2_X1 U15037 ( .A1(n11966), .A2(n13795), .ZN(n11986) );
  INV_X1 U15038 ( .A(n11986), .ZN(n11982) );
  INV_X1 U15039 ( .A(n11983), .ZN(n11985) );
  INV_X1 U15040 ( .A(n13430), .ZN(n11979) );
  INV_X1 U15041 ( .A(n11967), .ZN(n11978) );
  NAND2_X1 U15042 ( .A1(n11970), .A2(n11969), .ZN(n11974) );
  NAND2_X1 U15043 ( .A1(n11972), .A2(n11971), .ZN(n11973) );
  AOI21_X1 U15044 ( .B1(n11974), .B2(n20076), .A(n11973), .ZN(n11976) );
  NAND3_X1 U15045 ( .A1(n11977), .A2(n11976), .A3(n11975), .ZN(n13433) );
  AOI211_X1 U15046 ( .C1(n11979), .C2(n14092), .A(n11978), .B(n13433), .ZN(
        n11980) );
  NAND2_X1 U15047 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n13550), .ZN(
        n11981) );
  OAI22_X1 U15048 ( .A1(n16098), .A2(n11982), .B1(n11985), .B2(n11981), .ZN(
        n15095) );
  AOI21_X1 U15049 ( .B1(n15097), .B2(n11983), .A(n15095), .ZN(n16090) );
  NAND2_X1 U15050 ( .A1(n11989), .A2(n15138), .ZN(n15112) );
  NOR2_X1 U15051 ( .A1(n15113), .A2(n15112), .ZN(n15105) );
  NAND2_X1 U15052 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15105), .ZN(
        n15949) );
  NOR2_X1 U15053 ( .A1(n15088), .A2(n15949), .ZN(n15074) );
  NAND2_X1 U15054 ( .A1(n15074), .A2(n11984), .ZN(n15051) );
  NAND2_X1 U15055 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11993) );
  NOR2_X1 U15056 ( .A1(n15046), .A2(n15032), .ZN(n15009) );
  INV_X1 U15057 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20696) );
  NOR2_X1 U15058 ( .A1(n16134), .A2(n20696), .ZN(n14490) );
  INV_X1 U15059 ( .A(n16071), .ZN(n11990) );
  NOR2_X1 U15060 ( .A1(n16089), .A2(n11985), .ZN(n15118) );
  NAND2_X1 U15061 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n11986), .ZN(
        n15144) );
  INV_X1 U15062 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13552) );
  AOI22_X1 U15063 ( .A1(n16134), .A2(n11987), .B1(n13552), .B2(n13550), .ZN(
        n13547) );
  NOR2_X1 U15064 ( .A1(n11990), .A2(n15119), .ZN(n14219) );
  AOI21_X1 U15065 ( .B1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n15111), .A(
        n14219), .ZN(n15940) );
  AND2_X1 U15066 ( .A1(n16071), .A2(n15076), .ZN(n11994) );
  INV_X1 U15067 ( .A(n11994), .ZN(n11996) );
  INV_X1 U15068 ( .A(n14878), .ZN(n14903) );
  OR2_X1 U15069 ( .A1(n16071), .A2(n14903), .ZN(n11992) );
  OR2_X1 U15070 ( .A1(n16098), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11991) );
  INV_X1 U15071 ( .A(n11993), .ZN(n11995) );
  AOI21_X1 U15072 ( .B1(n15032), .B2(n11996), .A(n9605), .ZN(n15021) );
  OAI211_X1 U15073 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16071), .A(
        n15021), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15015) );
  INV_X2 U15074 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n12409) );
  NAND2_X1 U15075 ( .A1(n12409), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12110) );
  INV_X1 U15076 ( .A(n11472), .ZN(n12519) );
  INV_X1 U15077 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n12002) );
  OAI21_X1 U15078 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12025), .ZN(n19956) );
  AOI22_X1 U15079 ( .A1(n12538), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n12499), .B2(n19956), .ZN(n12001) );
  OAI21_X1 U15080 ( .B1(n12453), .B2(n12002), .A(n12001), .ZN(n12003) );
  AOI21_X1 U15081 ( .B1(n12036), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12003), .ZN(n12020) );
  NAND2_X1 U15082 ( .A1(n13680), .A2(n12125), .ZN(n12012) );
  INV_X1 U15083 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n12009) );
  INV_X1 U15084 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12008) );
  OAI22_X1 U15085 ( .A1(n12453), .A2(n12009), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n12008), .ZN(n12010) );
  AOI21_X1 U15086 ( .B1(n12036), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n12010), .ZN(n12011) );
  NAND2_X1 U15087 ( .A1(n12012), .A2(n12011), .ZN(n13534) );
  AOI21_X1 U15088 ( .B1(n12013), .B2(n11501), .A(n12409), .ZN(n13408) );
  NAND2_X1 U15089 ( .A1(n9594), .A2(n12125), .ZN(n12018) );
  INV_X1 U15090 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n12015) );
  INV_X1 U15091 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14101) );
  OAI22_X1 U15092 ( .A1(n12453), .A2(n12015), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14101), .ZN(n12016) );
  AOI21_X1 U15093 ( .B1(n12036), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12016), .ZN(n12017) );
  NAND2_X1 U15094 ( .A1(n12018), .A2(n12017), .ZN(n13407) );
  MUX2_X1 U15095 ( .A(n12499), .B(n13408), .S(n13407), .Z(n13533) );
  INV_X1 U15096 ( .A(n12020), .ZN(n12021) );
  NAND2_X1 U15097 ( .A1(n12019), .A2(n12021), .ZN(n12022) );
  NAND2_X1 U15098 ( .A1(n12023), .A2(n12022), .ZN(n13777) );
  OR2_X1 U15099 ( .A1(n20056), .A2(n12188), .ZN(n12032) );
  INV_X1 U15100 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n12029) );
  INV_X1 U15101 ( .A(n12025), .ZN(n12024) );
  INV_X1 U15102 ( .A(n12033), .ZN(n12027) );
  INV_X1 U15103 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n19943) );
  NAND2_X1 U15104 ( .A1(n19943), .A2(n12025), .ZN(n12026) );
  NAND2_X1 U15105 ( .A1(n12027), .A2(n12026), .ZN(n19949) );
  AOI22_X1 U15106 ( .A1(n19949), .A2(n12499), .B1(n12538), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12028) );
  OAI21_X1 U15107 ( .B1(n12453), .B2(n12029), .A(n12028), .ZN(n12030) );
  AOI21_X1 U15108 ( .B1(n12036), .B2(n20708), .A(n12030), .ZN(n12031) );
  NAND2_X1 U15109 ( .A1(n12032), .A2(n12031), .ZN(n13780) );
  NAND2_X1 U15110 ( .A1(n13777), .A2(n13780), .ZN(n13778) );
  NOR2_X1 U15111 ( .A1(n12033), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12034) );
  NOR2_X1 U15112 ( .A1(n12045), .A2(n12034), .ZN(n14004) );
  INV_X1 U15113 ( .A(n12036), .ZN(n12039) );
  INV_X1 U15114 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13664) );
  NAND2_X1 U15115 ( .A1(n12409), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12038) );
  NAND2_X1 U15116 ( .A1(n12539), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12037) );
  OAI211_X1 U15117 ( .C1(n12039), .C2(n13664), .A(n12038), .B(n12037), .ZN(
        n12040) );
  NAND2_X1 U15118 ( .A1(n12040), .A2(n12035), .ZN(n12041) );
  OAI21_X1 U15119 ( .B1(n14004), .B2(n12035), .A(n12041), .ZN(n12042) );
  NOR2_X2 U15120 ( .A1(n13778), .A2(n13805), .ZN(n13803) );
  NAND2_X1 U15121 ( .A1(n12044), .A2(n12125), .ZN(n12053) );
  INV_X1 U15122 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n12050) );
  INV_X1 U15123 ( .A(n12054), .ZN(n12048) );
  INV_X1 U15124 ( .A(n12045), .ZN(n12046) );
  INV_X1 U15125 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19920) );
  NAND2_X1 U15126 ( .A1(n12046), .A2(n19920), .ZN(n12047) );
  NAND2_X1 U15127 ( .A1(n12048), .A2(n12047), .ZN(n19929) );
  AOI22_X1 U15128 ( .A1(n19929), .A2(n12499), .B1(n12538), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12049) );
  OAI21_X1 U15129 ( .B1(n12453), .B2(n12050), .A(n12049), .ZN(n12051) );
  INV_X1 U15130 ( .A(n12051), .ZN(n12052) );
  NAND2_X1 U15131 ( .A1(n13803), .A2(n13842), .ZN(n13841) );
  INV_X1 U15132 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n14068) );
  OAI21_X1 U15133 ( .B1(n12054), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n12058), .ZN(n19916) );
  AOI22_X1 U15134 ( .A1(n19916), .A2(n12499), .B1(n12538), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12055) );
  OAI21_X1 U15135 ( .B1(n12453), .B2(n14068), .A(n12055), .ZN(n12056) );
  NOR2_X2 U15136 ( .A1(n13841), .A2(n14066), .ZN(n14065) );
  INV_X1 U15137 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n12062) );
  INV_X1 U15138 ( .A(n12058), .ZN(n12060) );
  INV_X1 U15139 ( .A(n12091), .ZN(n12059) );
  OAI21_X1 U15140 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n12060), .A(
        n12059), .ZN(n19902) );
  AOI22_X1 U15141 ( .A1(n12499), .A2(n19902), .B1(n12538), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12061) );
  OAI21_X1 U15142 ( .B1(n12453), .B2(n12062), .A(n12061), .ZN(n12063) );
  INV_X1 U15143 ( .A(n14163), .ZN(n12065) );
  NAND2_X1 U15144 ( .A1(n12539), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15145 ( .A1(n12273), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15146 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11518), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U15147 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12381), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12067) );
  AOI22_X1 U15148 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12066) );
  NAND4_X1 U15149 ( .A1(n12069), .A2(n12068), .A3(n12067), .A4(n12066), .ZN(
        n12075) );
  AOI22_X1 U15150 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12342), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12073) );
  AOI22_X1 U15151 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12072) );
  AOI22_X1 U15152 ( .A1(n11362), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U15153 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12070) );
  NAND4_X1 U15154 ( .A1(n12073), .A2(n12072), .A3(n12071), .A4(n12070), .ZN(
        n12074) );
  NOR2_X1 U15155 ( .A1(n12075), .A2(n12074), .ZN(n12076) );
  OR2_X1 U15156 ( .A1(n12188), .A2(n12076), .ZN(n12078) );
  XOR2_X1 U15157 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n12091), .Z(n14308) );
  INV_X1 U15158 ( .A(n14308), .ZN(n14227) );
  AOI22_X1 U15159 ( .A1(n12538), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n12499), .B2(n14227), .ZN(n12077) );
  INV_X1 U15160 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n14332) );
  AOI22_X1 U15161 ( .A1(n12273), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U15162 ( .A1(n11362), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U15163 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12479), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12081) );
  AOI22_X1 U15164 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12080) );
  NAND4_X1 U15165 ( .A1(n12083), .A2(n12082), .A3(n12081), .A4(n12080), .ZN(
        n12089) );
  AOI22_X1 U15166 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12436), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12087) );
  AOI22_X1 U15167 ( .A1(n11518), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12086) );
  AOI22_X1 U15168 ( .A1(n12289), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12085) );
  AOI22_X1 U15169 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12084) );
  NAND4_X1 U15170 ( .A1(n12087), .A2(n12086), .A3(n12085), .A4(n12084), .ZN(
        n12088) );
  NOR2_X1 U15171 ( .A1(n12089), .A2(n12088), .ZN(n12090) );
  OR2_X1 U15172 ( .A1(n12188), .A2(n12090), .ZN(n12094) );
  INV_X1 U15173 ( .A(n12095), .ZN(n12092) );
  XNOR2_X1 U15174 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n12092), .ZN(
        n14373) );
  AOI22_X1 U15175 ( .A1(n12499), .A2(n14373), .B1(n12538), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12093) );
  OAI211_X1 U15176 ( .C1(n12453), .C2(n14332), .A(n12094), .B(n12093), .ZN(
        n14327) );
  XOR2_X1 U15177 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B(n12109), .Z(
        n16054) );
  AOI22_X1 U15178 ( .A1(n12273), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11518), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12099) );
  AOI22_X1 U15179 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U15180 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U15181 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12096) );
  NAND4_X1 U15182 ( .A1(n12099), .A2(n12098), .A3(n12097), .A4(n12096), .ZN(
        n12105) );
  AOI22_X1 U15183 ( .A1(n11362), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12381), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12103) );
  AOI22_X1 U15184 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U15185 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U15186 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12100) );
  NAND4_X1 U15187 ( .A1(n12103), .A2(n12102), .A3(n12101), .A4(n12100), .ZN(
        n12104) );
  OR2_X1 U15188 ( .A1(n12105), .A2(n12104), .ZN(n12106) );
  AOI22_X1 U15189 ( .A1(n12125), .A2(n12106), .B1(n12538), .B2(
        P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12108) );
  NAND2_X1 U15190 ( .A1(n12539), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12107) );
  OAI211_X1 U15191 ( .C1(n16054), .C2(n12035), .A(n12108), .B(n12107), .ZN(
        n14334) );
  XNOR2_X1 U15192 ( .A(n12139), .B(n15991), .ZN(n15993) );
  NAND2_X1 U15193 ( .A1(n15993), .A2(n12499), .ZN(n12113) );
  INV_X1 U15194 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20005) );
  OAI22_X1 U15195 ( .A1(n12453), .A2(n20005), .B1(n12110), .B2(n15991), .ZN(
        n12111) );
  INV_X1 U15196 ( .A(n12111), .ZN(n12112) );
  NAND2_X1 U15197 ( .A1(n12113), .A2(n12112), .ZN(n12126) );
  AOI22_X1 U15198 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12485), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12117) );
  AOI22_X1 U15199 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12116) );
  AOI22_X1 U15200 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12436), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U15201 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12114) );
  NAND4_X1 U15202 ( .A1(n12117), .A2(n12116), .A3(n12115), .A4(n12114), .ZN(
        n12123) );
  AOI22_X1 U15203 ( .A1(n11518), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12381), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12121) );
  AOI22_X1 U15204 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12120) );
  AOI22_X1 U15205 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U15206 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12118) );
  NAND4_X1 U15207 ( .A1(n12121), .A2(n12120), .A3(n12119), .A4(n12118), .ZN(
        n12122) );
  OR2_X1 U15208 ( .A1(n12123), .A2(n12122), .ZN(n12124) );
  AND2_X1 U15209 ( .A1(n12125), .A2(n12124), .ZN(n14379) );
  NAND2_X1 U15210 ( .A1(n14380), .A2(n14379), .ZN(n14378) );
  INV_X1 U15211 ( .A(n12126), .ZN(n12127) );
  INV_X1 U15212 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14868) );
  AOI22_X1 U15213 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U15214 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12381), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12130) );
  AOI22_X1 U15215 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U15216 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12128) );
  NAND4_X1 U15217 ( .A1(n12131), .A2(n12130), .A3(n12129), .A4(n12128), .ZN(
        n12137) );
  AOI22_X1 U15218 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12479), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12135) );
  AOI22_X1 U15219 ( .A1(n11518), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U15220 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15221 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12132) );
  NAND4_X1 U15222 ( .A1(n12135), .A2(n12134), .A3(n12133), .A4(n12132), .ZN(
        n12136) );
  NOR2_X1 U15223 ( .A1(n12137), .A2(n12136), .ZN(n12138) );
  OR2_X1 U15224 ( .A1(n12188), .A2(n12138), .ZN(n12141) );
  XNOR2_X1 U15225 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12142), .ZN(
        n14997) );
  AOI22_X1 U15226 ( .A1(n12499), .A2(n14997), .B1(n12538), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12140) );
  OAI211_X1 U15227 ( .C1(n12453), .C2(n14868), .A(n12141), .B(n12140), .ZN(
        n14734) );
  XOR2_X1 U15228 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12157), .Z(
        n16050) );
  INV_X1 U15229 ( .A(n16050), .ZN(n15989) );
  AOI22_X1 U15230 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11412), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U15231 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12145) );
  AOI22_X1 U15232 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12381), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12144) );
  AOI22_X1 U15233 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12143) );
  NAND4_X1 U15234 ( .A1(n12146), .A2(n12145), .A3(n12144), .A4(n12143), .ZN(
        n12152) );
  AOI22_X1 U15235 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12479), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U15236 ( .A1(n11518), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U15237 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15238 ( .A1(n12422), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12147) );
  NAND4_X1 U15239 ( .A1(n12150), .A2(n12149), .A3(n12148), .A4(n12147), .ZN(
        n12151) );
  NOR2_X1 U15240 ( .A1(n12152), .A2(n12151), .ZN(n12155) );
  NAND2_X1 U15241 ( .A1(n12539), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12154) );
  NAND2_X1 U15242 ( .A1(n12538), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12153) );
  OAI211_X1 U15243 ( .C1(n12188), .C2(n12155), .A(n12154), .B(n12153), .ZN(
        n12156) );
  AOI21_X1 U15244 ( .B1(n15989), .B2(n12499), .A(n12156), .ZN(n14787) );
  INV_X1 U15245 ( .A(n14721), .ZN(n12173) );
  XNOR2_X1 U15246 ( .A(n12174), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14987) );
  AOI22_X1 U15247 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12161) );
  AOI22_X1 U15248 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12485), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12160) );
  AOI22_X1 U15249 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15250 ( .A1(n12422), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11407), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12158) );
  NAND4_X1 U15251 ( .A1(n12161), .A2(n12160), .A3(n12159), .A4(n12158), .ZN(
        n12167) );
  AOI22_X1 U15252 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11517), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12165) );
  AOI22_X1 U15253 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12359), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U15254 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12436), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12163) );
  AOI22_X1 U15255 ( .A1(n12289), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12162) );
  NAND4_X1 U15256 ( .A1(n12165), .A2(n12164), .A3(n12163), .A4(n12162), .ZN(
        n12166) );
  NOR2_X1 U15257 ( .A1(n12167), .A2(n12166), .ZN(n12170) );
  NAND2_X1 U15258 ( .A1(n12539), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12169) );
  NAND2_X1 U15259 ( .A1(n12538), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12168) );
  OAI211_X1 U15260 ( .C1(n12188), .C2(n12170), .A(n12169), .B(n12168), .ZN(
        n12171) );
  AOI21_X1 U15261 ( .B1(n14987), .B2(n12499), .A(n12171), .ZN(n14722) );
  NAND2_X1 U15262 ( .A1(n12173), .A2(n12172), .ZN(n14723) );
  XOR2_X1 U15263 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n12190), .Z(
        n15972) );
  INV_X1 U15264 ( .A(n15972), .ZN(n16040) );
  AOI22_X1 U15265 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12475), .B1(
        n12381), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U15266 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n12479), .B1(
        n12436), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12177) );
  AOI22_X1 U15267 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11407), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12176) );
  AOI22_X1 U15268 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12175) );
  NAND4_X1 U15269 ( .A1(n12178), .A2(n12177), .A3(n12176), .A4(n12175), .ZN(
        n12184) );
  AOI22_X1 U15270 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12435), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12182) );
  AOI22_X1 U15271 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n12485), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15272 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n11518), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15273 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12179) );
  NAND4_X1 U15274 ( .A1(n12182), .A2(n12181), .A3(n12180), .A4(n12179), .ZN(
        n12183) );
  NOR2_X1 U15275 ( .A1(n12184), .A2(n12183), .ZN(n12187) );
  NAND2_X1 U15276 ( .A1(n12539), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12186) );
  NAND2_X1 U15277 ( .A1(n12538), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12185) );
  OAI211_X1 U15278 ( .C1(n12188), .C2(n12187), .A(n12186), .B(n12185), .ZN(
        n12189) );
  AOI21_X1 U15279 ( .B1(n16040), .B2(n12499), .A(n12189), .ZN(n14777) );
  XNOR2_X1 U15280 ( .A(n12204), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14977) );
  AOI21_X1 U15281 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14972), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12191) );
  AOI21_X1 U15282 ( .B1(n12539), .B2(P1_EAX_REG_16__SCAN_IN), .A(n12191), .ZN(
        n12203) );
  AOI22_X1 U15283 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11412), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15284 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12436), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15285 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11407), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U15286 ( .A1(n12289), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12192) );
  NAND4_X1 U15287 ( .A1(n12195), .A2(n12194), .A3(n12193), .A4(n12192), .ZN(
        n12201) );
  AOI22_X1 U15288 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U15289 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12381), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U15290 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12479), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12197) );
  AOI22_X1 U15291 ( .A1(n11518), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12196) );
  NAND4_X1 U15292 ( .A1(n12199), .A2(n12198), .A3(n12197), .A4(n12196), .ZN(
        n12200) );
  OAI21_X1 U15293 ( .B1(n12201), .B2(n12200), .A(n12496), .ZN(n12202) );
  AOI22_X1 U15294 ( .A1(n14977), .A2(n12499), .B1(n12203), .B2(n12202), .ZN(
        n14709) );
  XOR2_X1 U15295 ( .A(n14700), .B(n12220), .Z(n16028) );
  INV_X1 U15296 ( .A(n16028), .ZN(n12219) );
  AOI22_X1 U15297 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11412), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U15298 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U15299 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U15300 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12436), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12205) );
  NAND4_X1 U15301 ( .A1(n12208), .A2(n12207), .A3(n12206), .A4(n12205), .ZN(
        n12214) );
  AOI22_X1 U15302 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15303 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12211) );
  AOI22_X1 U15304 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15305 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11407), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12209) );
  NAND4_X1 U15306 ( .A1(n12212), .A2(n12211), .A3(n12210), .A4(n12209), .ZN(
        n12213) );
  NOR2_X1 U15307 ( .A1(n12214), .A2(n12213), .ZN(n12217) );
  NAND2_X1 U15308 ( .A1(n12539), .A2(P1_EAX_REG_17__SCAN_IN), .ZN(n12216) );
  NAND2_X1 U15309 ( .A1(n12538), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12215) );
  OAI211_X1 U15310 ( .C1(n12450), .C2(n12217), .A(n12216), .B(n12215), .ZN(
        n12218) );
  AOI21_X1 U15311 ( .B1(n12219), .B2(n12499), .A(n12218), .ZN(n14695) );
  XNOR2_X1 U15312 ( .A(n12250), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14684) );
  AOI22_X1 U15313 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15314 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12223) );
  AOI22_X1 U15315 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12222) );
  AOI22_X1 U15316 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12221) );
  NAND4_X1 U15317 ( .A1(n12224), .A2(n12223), .A3(n12222), .A4(n12221), .ZN(
        n12230) );
  AOI22_X1 U15318 ( .A1(n12273), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11412), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15319 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15320 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12436), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15321 ( .A1(n12422), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11407), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12225) );
  NAND4_X1 U15322 ( .A1(n12228), .A2(n12227), .A3(n12226), .A4(n12225), .ZN(
        n12229) );
  OAI21_X1 U15323 ( .B1(n12230), .B2(n12229), .A(n12496), .ZN(n12233) );
  INV_X1 U15324 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14847) );
  INV_X1 U15325 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14960) );
  OAI22_X1 U15326 ( .A1(n12453), .A2(n14847), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14960), .ZN(n12231) );
  INV_X1 U15327 ( .A(n12231), .ZN(n12232) );
  AOI21_X1 U15328 ( .B1(n12233), .B2(n12232), .A(n12499), .ZN(n12234) );
  AOI21_X1 U15329 ( .B1(n14684), .B2(n12499), .A(n12234), .ZN(n14682) );
  AOI22_X1 U15330 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11518), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12239) );
  AOI22_X1 U15331 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12381), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12238) );
  AOI22_X1 U15332 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11407), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12237) );
  AOI22_X1 U15333 ( .A1(n12289), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12236) );
  NAND4_X1 U15334 ( .A1(n12239), .A2(n12238), .A3(n12237), .A4(n12236), .ZN(
        n12245) );
  AOI22_X1 U15335 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12479), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12243) );
  AOI22_X1 U15336 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12436), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12242) );
  AOI22_X1 U15337 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12241) );
  AOI22_X1 U15338 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12240) );
  NAND4_X1 U15339 ( .A1(n12243), .A2(n12242), .A3(n12241), .A4(n12240), .ZN(
        n12244) );
  NOR2_X1 U15340 ( .A1(n12245), .A2(n12244), .ZN(n12249) );
  INV_X1 U15341 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14843) );
  NAND2_X1 U15342 ( .A1(n12409), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12246) );
  OAI211_X1 U15343 ( .C1(n12453), .C2(n14843), .A(n12035), .B(n12246), .ZN(
        n12247) );
  INV_X1 U15344 ( .A(n12247), .ZN(n12248) );
  OAI21_X1 U15345 ( .B1(n12450), .B2(n12249), .A(n12248), .ZN(n12253) );
  OAI21_X1 U15346 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n12251), .A(
        n12298), .ZN(n16027) );
  OR2_X1 U15347 ( .A1(n12035), .A2(n16027), .ZN(n12252) );
  NAND2_X1 U15348 ( .A1(n12253), .A2(n12252), .ZN(n14669) );
  NOR2_X2 U15349 ( .A1(n14668), .A2(n14669), .ZN(n14644) );
  AOI22_X1 U15350 ( .A1(n11362), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12257) );
  AOI22_X1 U15351 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12479), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12256) );
  AOI22_X1 U15352 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U15353 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12254) );
  NAND4_X1 U15354 ( .A1(n12257), .A2(n12256), .A3(n12255), .A4(n12254), .ZN(
        n12263) );
  AOI22_X1 U15355 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12381), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12261) );
  AOI22_X1 U15356 ( .A1(n12273), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12260) );
  AOI22_X1 U15357 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12259) );
  AOI22_X1 U15358 ( .A1(n12289), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12258) );
  NAND4_X1 U15359 ( .A1(n12261), .A2(n12260), .A3(n12259), .A4(n12258), .ZN(
        n12262) );
  OAI21_X1 U15360 ( .B1(n12263), .B2(n12262), .A(n12496), .ZN(n12267) );
  INV_X1 U15361 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14826) );
  NAND2_X1 U15362 ( .A1(n12409), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12264) );
  OAI211_X1 U15363 ( .C1(n12453), .C2(n14826), .A(n12035), .B(n12264), .ZN(
        n12265) );
  INV_X1 U15364 ( .A(n12265), .ZN(n12266) );
  XNOR2_X1 U15365 ( .A(n12327), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14941) );
  AOI22_X1 U15366 ( .A1(n12267), .A2(n12266), .B1(n12499), .B2(n14941), .ZN(
        n14646) );
  INV_X1 U15367 ( .A(n14646), .ZN(n12284) );
  OAI21_X1 U15368 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n12268), .A(
        n12327), .ZN(n16021) );
  AOI22_X1 U15369 ( .A1(n11412), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11517), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15370 ( .A1(n11391), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12359), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12271) );
  AOI22_X1 U15371 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U15372 ( .A1(n12289), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12269) );
  NAND4_X1 U15373 ( .A1(n12272), .A2(n12271), .A3(n12270), .A4(n12269), .ZN(
        n12279) );
  AOI22_X1 U15374 ( .A1(n11362), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12277) );
  AOI22_X1 U15375 ( .A1(n12476), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12485), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U15376 ( .A1(n12273), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12275) );
  AOI22_X1 U15377 ( .A1(n12422), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12274) );
  NAND4_X1 U15378 ( .A1(n12277), .A2(n12276), .A3(n12275), .A4(n12274), .ZN(
        n12278) );
  OAI21_X1 U15379 ( .B1(n12279), .B2(n12278), .A(n12496), .ZN(n12282) );
  NAND2_X1 U15380 ( .A1(n12539), .A2(P1_EAX_REG_21__SCAN_IN), .ZN(n12281) );
  NAND2_X1 U15381 ( .A1(n12409), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12280) );
  NAND4_X1 U15382 ( .A1(n12282), .A2(n12035), .A3(n12281), .A4(n12280), .ZN(
        n12283) );
  OAI21_X1 U15383 ( .B1(n12035), .B2(n16021), .A(n12283), .ZN(n14832) );
  AOI22_X1 U15384 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11518), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12288) );
  AOI22_X1 U15385 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12287) );
  AOI22_X1 U15386 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12436), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12286) );
  AOI22_X1 U15387 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11407), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12285) );
  NAND4_X1 U15388 ( .A1(n12288), .A2(n12287), .A3(n12286), .A4(n12285), .ZN(
        n12296) );
  AOI22_X1 U15389 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12289), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12294) );
  AOI22_X1 U15390 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U15391 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12292) );
  AOI22_X1 U15392 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12290), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12291) );
  NAND4_X1 U15393 ( .A1(n12294), .A2(n12293), .A3(n12292), .A4(n12291), .ZN(
        n12295) );
  OAI21_X1 U15394 ( .B1(n12296), .B2(n12295), .A(n12496), .ZN(n12300) );
  AOI21_X1 U15395 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14956), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12297) );
  AOI21_X1 U15396 ( .B1(n12539), .B2(P1_EAX_REG_20__SCAN_IN), .A(n12297), .ZN(
        n12299) );
  XNOR2_X1 U15397 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n12298), .ZN(
        n14954) );
  AOI22_X1 U15398 ( .A1(n12300), .A2(n12299), .B1(n12499), .B2(n14954), .ZN(
        n14660) );
  NAND2_X1 U15399 ( .A1(n14644), .A2(n12303), .ZN(n14634) );
  AOI22_X1 U15400 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12307) );
  AOI22_X1 U15401 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U15402 ( .A1(n11518), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12305) );
  AOI22_X1 U15403 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12478), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12304) );
  NAND4_X1 U15404 ( .A1(n12307), .A2(n12306), .A3(n12305), .A4(n12304), .ZN(
        n12313) );
  AOI22_X1 U15405 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12311) );
  AOI22_X1 U15406 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12310) );
  AOI22_X1 U15407 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U15408 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12308) );
  NAND4_X1 U15409 ( .A1(n12311), .A2(n12310), .A3(n12309), .A4(n12308), .ZN(
        n12312) );
  NOR2_X1 U15410 ( .A1(n12313), .A2(n12312), .ZN(n12336) );
  AOI22_X1 U15411 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12435), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12318) );
  AOI22_X1 U15412 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n12485), .B1(
        n12479), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12317) );
  AOI22_X1 U15413 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12316) );
  AOI22_X1 U15414 ( .A1(n12314), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12315) );
  NAND4_X1 U15415 ( .A1(n12318), .A2(n12317), .A3(n12316), .A4(n12315), .ZN(
        n12324) );
  AOI22_X1 U15416 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n12484), .B1(
        n11518), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12322) );
  AOI22_X1 U15417 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12475), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12321) );
  AOI22_X1 U15418 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12320) );
  AOI22_X1 U15419 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12394), .B1(
        n12478), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12319) );
  NAND4_X1 U15420 ( .A1(n12322), .A2(n12321), .A3(n12320), .A4(n12319), .ZN(
        n12323) );
  NOR2_X1 U15421 ( .A1(n12324), .A2(n12323), .ZN(n12335) );
  XNOR2_X1 U15422 ( .A(n12336), .B(n12335), .ZN(n12325) );
  NOR2_X1 U15423 ( .A1(n12450), .A2(n12325), .ZN(n12333) );
  INV_X1 U15424 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14822) );
  NAND2_X1 U15425 ( .A1(n12409), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12326) );
  OAI211_X1 U15426 ( .C1(n12453), .C2(n14822), .A(n12035), .B(n12326), .ZN(
        n12332) );
  INV_X1 U15427 ( .A(n12329), .ZN(n12330) );
  INV_X1 U15428 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14636) );
  NAND2_X1 U15429 ( .A1(n12330), .A2(n14636), .ZN(n12331) );
  NAND2_X1 U15430 ( .A1(n12370), .A2(n12331), .ZN(n14934) );
  OAI22_X1 U15431 ( .A1(n12333), .A2(n12332), .B1(n12035), .B2(n14934), .ZN(
        n14635) );
  XNOR2_X1 U15432 ( .A(n12370), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14924) );
  INV_X1 U15433 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12334) );
  AOI21_X1 U15434 ( .B1(n12334), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12353) );
  NOR2_X1 U15435 ( .A1(n12336), .A2(n12335), .ZN(n12367) );
  INV_X1 U15436 ( .A(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12337) );
  NOR2_X1 U15437 ( .A1(n11350), .A2(n12337), .ZN(n12341) );
  INV_X1 U15438 ( .A(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12339) );
  INV_X1 U15439 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12338) );
  OAI22_X1 U15440 ( .A1(n11553), .A2(n12339), .B1(n11519), .B2(n12338), .ZN(
        n12340) );
  AOI211_X1 U15441 ( .C1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .C2(n12484), .A(
        n12341), .B(n12340), .ZN(n12350) );
  AOI22_X1 U15442 ( .A1(n12422), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12349) );
  AOI22_X1 U15443 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12348) );
  AOI22_X1 U15444 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12346) );
  AOI22_X1 U15445 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12345) );
  AOI22_X1 U15446 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12344) );
  AOI22_X1 U15447 ( .A1(n12342), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12478), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12343) );
  AND4_X1 U15448 ( .A1(n12346), .A2(n12345), .A3(n12344), .A4(n12343), .ZN(
        n12347) );
  NAND4_X1 U15449 ( .A1(n12350), .A2(n12349), .A3(n12348), .A4(n12347), .ZN(
        n12366) );
  XNOR2_X1 U15450 ( .A(n12367), .B(n12366), .ZN(n12351) );
  NOR2_X1 U15451 ( .A1(n12351), .A2(n12450), .ZN(n12352) );
  AOI211_X1 U15452 ( .C1(n12539), .C2(P1_EAX_REG_24__SCAN_IN), .A(n12353), .B(
        n12352), .ZN(n12354) );
  AOI21_X1 U15453 ( .B1(n12499), .B2(n14924), .A(n12354), .ZN(n14625) );
  NAND2_X1 U15454 ( .A1(n14624), .A2(n14625), .ZN(n14611) );
  AOI22_X1 U15455 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U15456 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12357) );
  AOI22_X1 U15457 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12479), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12356) );
  AOI22_X1 U15458 ( .A1(n11518), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12355) );
  NAND4_X1 U15459 ( .A1(n12358), .A2(n12357), .A3(n12356), .A4(n12355), .ZN(
        n12365) );
  AOI22_X1 U15460 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12435), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12363) );
  AOI22_X1 U15461 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12362) );
  AOI22_X1 U15462 ( .A1(n12422), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U15463 ( .A1(n12394), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12478), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12360) );
  NAND4_X1 U15464 ( .A1(n12363), .A2(n12362), .A3(n12361), .A4(n12360), .ZN(
        n12364) );
  NOR2_X1 U15465 ( .A1(n12365), .A2(n12364), .ZN(n12389) );
  NAND2_X1 U15466 ( .A1(n12367), .A2(n12366), .ZN(n12388) );
  XNOR2_X1 U15467 ( .A(n12389), .B(n12388), .ZN(n12368) );
  NOR2_X1 U15468 ( .A1(n12368), .A2(n12450), .ZN(n12376) );
  INV_X1 U15469 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14814) );
  NAND2_X1 U15470 ( .A1(n12409), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12369) );
  OAI211_X1 U15471 ( .C1(n12453), .C2(n14814), .A(n12035), .B(n12369), .ZN(
        n12375) );
  INV_X1 U15472 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12372) );
  NAND2_X1 U15473 ( .A1(n12373), .A2(n12372), .ZN(n12374) );
  NAND2_X1 U15474 ( .A1(n12412), .A2(n12374), .ZN(n14916) );
  NOR2_X2 U15475 ( .A1(n14611), .A2(n14613), .ZN(n14600) );
  XNOR2_X1 U15476 ( .A(n12412), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14902) );
  AOI22_X1 U15477 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12380) );
  INV_X1 U15478 ( .A(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n20870) );
  AOI22_X1 U15479 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12379) );
  AOI22_X1 U15480 ( .A1(n11518), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12378) );
  AOI22_X1 U15481 ( .A1(n12422), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12377) );
  NAND4_X1 U15482 ( .A1(n12380), .A2(n12379), .A3(n12378), .A4(n12377), .ZN(
        n12387) );
  AOI22_X1 U15483 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12381), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12385) );
  AOI22_X1 U15484 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12384) );
  AOI22_X1 U15485 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12383) );
  AOI22_X1 U15486 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12478), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12382) );
  NAND4_X1 U15487 ( .A1(n12385), .A2(n12384), .A3(n12383), .A4(n12382), .ZN(
        n12386) );
  OR2_X1 U15488 ( .A1(n12387), .A2(n12386), .ZN(n12406) );
  NOR2_X1 U15489 ( .A1(n12389), .A2(n12388), .ZN(n12407) );
  XOR2_X1 U15490 ( .A(n12406), .B(n12407), .Z(n12392) );
  INV_X1 U15491 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14810) );
  NAND2_X1 U15492 ( .A1(n12409), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12390) );
  OAI211_X1 U15493 ( .C1(n12453), .C2(n14810), .A(n12035), .B(n12390), .ZN(
        n12391) );
  AOI21_X1 U15494 ( .B1(n12392), .B2(n12496), .A(n12391), .ZN(n12393) );
  AOI22_X1 U15495 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12399) );
  AOI22_X1 U15496 ( .A1(n11517), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12398) );
  AOI22_X1 U15497 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12478), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12397) );
  AOI22_X1 U15498 ( .A1(n12422), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12396) );
  NAND4_X1 U15499 ( .A1(n12399), .A2(n12398), .A3(n12397), .A4(n12396), .ZN(
        n12405) );
  AOI22_X1 U15500 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12403) );
  AOI22_X1 U15501 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12402) );
  AOI22_X1 U15502 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12401) );
  AOI22_X1 U15503 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12400) );
  NAND4_X1 U15504 ( .A1(n12403), .A2(n12402), .A3(n12401), .A4(n12400), .ZN(
        n12404) );
  NOR2_X1 U15505 ( .A1(n12405), .A2(n12404), .ZN(n12430) );
  NAND2_X1 U15506 ( .A1(n12407), .A2(n12406), .ZN(n12429) );
  XNOR2_X1 U15507 ( .A(n12430), .B(n12429), .ZN(n12408) );
  NOR2_X1 U15508 ( .A1(n12408), .A2(n12450), .ZN(n12417) );
  INV_X1 U15509 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n12411) );
  NAND2_X1 U15510 ( .A1(n12409), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12410) );
  OAI211_X1 U15511 ( .C1(n12453), .C2(n12411), .A(n12035), .B(n12410), .ZN(
        n12416) );
  INV_X1 U15512 ( .A(n12412), .ZN(n12413) );
  NAND2_X1 U15513 ( .A1(n12413), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12414) );
  INV_X1 U15514 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14592) );
  NAND2_X1 U15515 ( .A1(n12414), .A2(n14592), .ZN(n12415) );
  NAND2_X1 U15516 ( .A1(n12454), .A2(n12415), .ZN(n14896) );
  OAI22_X1 U15517 ( .A1(n12417), .A2(n12416), .B1(n12035), .B2(n14896), .ZN(
        n14588) );
  XNOR2_X1 U15518 ( .A(n12454), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14578) );
  AOI22_X1 U15519 ( .A1(n11362), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12421) );
  AOI22_X1 U15520 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12420) );
  AOI22_X1 U15521 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12419) );
  AOI22_X1 U15522 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12478), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12418) );
  NAND4_X1 U15523 ( .A1(n12421), .A2(n12420), .A3(n12419), .A4(n12418), .ZN(
        n12428) );
  AOI22_X1 U15524 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12426) );
  AOI22_X1 U15525 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12425) );
  AOI22_X1 U15526 ( .A1(n11518), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9593), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12424) );
  AOI22_X1 U15527 ( .A1(n12422), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12423) );
  NAND4_X1 U15528 ( .A1(n12426), .A2(n12425), .A3(n12424), .A4(n12423), .ZN(
        n12427) );
  OR2_X1 U15529 ( .A1(n12428), .A2(n12427), .ZN(n12448) );
  NOR2_X1 U15530 ( .A1(n12430), .A2(n12429), .ZN(n12449) );
  XOR2_X1 U15531 ( .A(n12448), .B(n12449), .Z(n12433) );
  INV_X1 U15532 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14802) );
  NAND2_X1 U15533 ( .A1(n12409), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12431) );
  OAI211_X1 U15534 ( .C1(n12453), .C2(n14802), .A(n12035), .B(n12431), .ZN(
        n12432) );
  AOI21_X1 U15535 ( .B1(n12433), .B2(n12496), .A(n12432), .ZN(n12434) );
  AOI22_X1 U15536 ( .A1(n12435), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12440) );
  AOI22_X1 U15537 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12436), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12439) );
  AOI22_X1 U15538 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U15539 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12478), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12437) );
  NAND4_X1 U15540 ( .A1(n12440), .A2(n12439), .A3(n12438), .A4(n12437), .ZN(
        n12447) );
  AOI22_X1 U15541 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12445) );
  AOI22_X1 U15542 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12444) );
  AOI22_X1 U15543 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12443) );
  AOI22_X1 U15544 ( .A1(n11518), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12442) );
  NAND4_X1 U15545 ( .A1(n12445), .A2(n12444), .A3(n12443), .A4(n12442), .ZN(
        n12446) );
  NOR2_X1 U15546 ( .A1(n12447), .A2(n12446), .ZN(n12474) );
  NAND2_X1 U15547 ( .A1(n12449), .A2(n12448), .ZN(n12473) );
  XNOR2_X1 U15548 ( .A(n12474), .B(n12473), .ZN(n12451) );
  NOR2_X1 U15549 ( .A1(n12451), .A2(n12450), .ZN(n12460) );
  INV_X1 U15550 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14797) );
  NAND2_X1 U15551 ( .A1(n12409), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12452) );
  OAI211_X1 U15552 ( .C1(n12453), .C2(n14797), .A(n12035), .B(n12452), .ZN(
        n12459) );
  INV_X1 U15553 ( .A(n12454), .ZN(n12455) );
  NAND2_X1 U15554 ( .A1(n12455), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12457) );
  INV_X1 U15555 ( .A(n12457), .ZN(n12458) );
  INV_X1 U15556 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12456) );
  OAI21_X1 U15557 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n12458), .A(
        n14097), .ZN(n14874) );
  OAI22_X1 U15558 ( .A1(n12460), .A2(n12459), .B1(n12035), .B2(n14874), .ZN(
        n12461) );
  INV_X1 U15559 ( .A(n12537), .ZN(n12463) );
  INV_X1 U15560 ( .A(n12000), .ZN(n14525) );
  NAND3_X1 U15561 ( .A1(n14525), .A2(n12464), .A3(n9843), .ZN(n12516) );
  OR3_X1 U15562 ( .A1(n12516), .A2(n12465), .A3(n11914), .ZN(n12466) );
  NAND2_X1 U15563 ( .A1(n13454), .A2(n12466), .ZN(n12467) );
  NAND2_X2 U15564 ( .A1(n19997), .A2(n12000), .ZN(n19992) );
  OAI21_X1 U15565 ( .B1(n14576), .B2(n12468), .A(n9657), .ZN(n15019) );
  NAND2_X1 U15566 ( .A1(n12469), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n12470) );
  NOR2_X1 U15567 ( .A1(n12474), .A2(n12473), .ZN(n12495) );
  AOI22_X1 U15568 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12475), .B1(
        n11517), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12483) );
  AOI22_X1 U15569 ( .A1(n11362), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12476), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12482) );
  AOI22_X1 U15570 ( .A1(n12395), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12477), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12481) );
  AOI22_X1 U15571 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12478), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12480) );
  NAND4_X1 U15572 ( .A1(n12483), .A2(n12482), .A3(n12481), .A4(n12480), .ZN(
        n12493) );
  AOI22_X1 U15573 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n12441), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12491) );
  AOI22_X1 U15574 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n12485), .B1(
        n12394), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12490) );
  AOI22_X1 U15575 ( .A1(n12359), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12486), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12489) );
  AOI22_X1 U15576 ( .A1(n9593), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12487), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12488) );
  NAND4_X1 U15577 ( .A1(n12491), .A2(n12490), .A3(n12489), .A4(n12488), .ZN(
        n12492) );
  NOR2_X1 U15578 ( .A1(n12493), .A2(n12492), .ZN(n12494) );
  XNOR2_X1 U15579 ( .A(n12495), .B(n12494), .ZN(n12497) );
  NAND2_X1 U15580 ( .A1(n12497), .A2(n12496), .ZN(n12501) );
  INV_X1 U15581 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n20877) );
  NOR2_X1 U15582 ( .A1(n20877), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12498) );
  AOI211_X1 U15583 ( .C1(n12539), .C2(P1_EAX_REG_30__SCAN_IN), .A(n12498), .B(
        n12499), .ZN(n12500) );
  XNOR2_X1 U15584 ( .A(n14097), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14533) );
  INV_X1 U15585 ( .A(n12502), .ZN(n12503) );
  AOI22_X1 U15586 ( .A1(n9657), .A2(n13281), .B1(n12503), .B2(n14576), .ZN(
        n12505) );
  XNOR2_X1 U15587 ( .A(n12505), .B(n12504), .ZN(n15012) );
  INV_X1 U15588 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n12506) );
  AOI21_X1 U15589 ( .B1(n12509), .B2(n12508), .A(n12507), .ZN(n12510) );
  INV_X1 U15590 ( .A(n13444), .ZN(n15936) );
  NAND2_X1 U15591 ( .A1(n13444), .A2(n20647), .ZN(n13448) );
  OAI22_X1 U15592 ( .A1(n12514), .A2(n13448), .B1(n13431), .B2(n12516), .ZN(
        n12517) );
  NAND2_X1 U15593 ( .A1(n14867), .A2(n12519), .ZN(n12531) );
  INV_X1 U15594 ( .A(n12531), .ZN(n12530) );
  NOR4_X1 U15595 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_ADDRESS_REG_15__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_13__SCAN_IN), .ZN(n12523) );
  NOR4_X1 U15596 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(
        P1_ADDRESS_REG_19__SCAN_IN), .A3(P1_ADDRESS_REG_18__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n12522) );
  NOR4_X1 U15597 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12521) );
  NOR4_X1 U15598 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(
        P1_ADDRESS_REG_11__SCAN_IN), .A3(P1_ADDRESS_REG_10__SCAN_IN), .A4(
        P1_ADDRESS_REG_9__SCAN_IN), .ZN(n12520) );
  AND4_X1 U15599 ( .A1(n12523), .A2(n12522), .A3(n12521), .A4(n12520), .ZN(
        n12528) );
  NOR4_X1 U15600 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_6__SCAN_IN), .ZN(n12526) );
  NOR4_X1 U15601 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(
        P1_ADDRESS_REG_23__SCAN_IN), .A3(P1_ADDRESS_REG_22__SCAN_IN), .A4(
        P1_ADDRESS_REG_21__SCAN_IN), .ZN(n12525) );
  NOR4_X1 U15602 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(
        P1_ADDRESS_REG_27__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_25__SCAN_IN), .ZN(n12524) );
  INV_X1 U15603 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20656) );
  AND4_X1 U15604 ( .A1(n12526), .A2(n12525), .A3(n12524), .A4(n20656), .ZN(
        n12527) );
  NAND2_X1 U15605 ( .A1(n12528), .A2(n12527), .ZN(n12529) );
  NAND2_X1 U15606 ( .A1(n12530), .A2(n20053), .ZN(n14836) );
  INV_X1 U15607 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19165) );
  NOR2_X1 U15608 ( .A1(n14836), .A2(n19165), .ZN(n12535) );
  AOI22_X1 U15609 ( .A1(n12532), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14861), .ZN(n12533) );
  INV_X1 U15610 ( .A(n12533), .ZN(n12534) );
  NOR2_X1 U15611 ( .A1(n12535), .A2(n12534), .ZN(n12545) );
  NAND2_X1 U15612 ( .A1(n12537), .A2(n12536), .ZN(n12542) );
  AOI22_X1 U15613 ( .A1(n12539), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n12538), .ZN(n12540) );
  INV_X1 U15614 ( .A(n12540), .ZN(n12541) );
  AND2_X1 U15615 ( .A1(n14867), .A2(n14525), .ZN(n12543) );
  NAND2_X1 U15616 ( .A1(n12545), .A2(n12544), .ZN(P1_U2873) );
  OAI21_X1 U15617 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18637), .A(
        n12674), .ZN(n12676) );
  OAI22_X1 U15618 ( .A1(n12565), .A2(n18638), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12675) );
  INV_X1 U15619 ( .A(n12675), .ZN(n12546) );
  OR2_X1 U15620 ( .A1(n12676), .A2(n12546), .ZN(n12560) );
  OAI22_X1 U15621 ( .A1(n18808), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18670), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12551) );
  NOR2_X1 U15622 ( .A1(n12552), .A2(n12551), .ZN(n12548) );
  NOR2_X1 U15623 ( .A1(n12549), .A2(n18798), .ZN(n12554) );
  NAND2_X1 U15624 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18631), .ZN(
        n12550) );
  AOI22_X1 U15625 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18631), .B1(
        n12549), .B2(n18798), .ZN(n12553) );
  OAI22_X1 U15626 ( .A1(n12554), .A2(n12550), .B1(n12553), .B2(n18665), .ZN(
        n12559) );
  XNOR2_X1 U15627 ( .A(n12552), .B(n12551), .ZN(n12557) );
  OAI21_X1 U15628 ( .B1(n18665), .B2(n12554), .A(n12553), .ZN(n12555) );
  OAI21_X1 U15629 ( .B1(n18631), .B2(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n12555), .ZN(n12556) );
  INV_X1 U15630 ( .A(n12556), .ZN(n12672) );
  OAI21_X1 U15631 ( .B1(n12557), .B2(n12559), .A(n12672), .ZN(n12558) );
  INV_X1 U15632 ( .A(n12558), .ZN(n13257) );
  OAI21_X1 U15633 ( .B1(n12560), .B2(n12559), .A(n13257), .ZN(n15869) );
  NOR2_X2 U15634 ( .A1(n18650), .A2(n12561), .ZN(n12703) );
  INV_X4 U15635 ( .A(n12704), .ZN(n17150) );
  AOI22_X1 U15636 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12562) );
  OAI21_X1 U15637 ( .B1(n12605), .B2(n20845), .A(n12562), .ZN(n12574) );
  AOI22_X1 U15639 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17132), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12572) );
  NOR2_X2 U15640 ( .A1(n18650), .A2(n12567), .ZN(n12692) );
  AOI22_X1 U15641 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12571) );
  NOR2_X1 U15642 ( .A1(n12566), .A2(n12568), .ZN(n12677) );
  AOI22_X1 U15643 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12570) );
  INV_X1 U15644 ( .A(n12689), .ZN(n12578) );
  AOI22_X1 U15645 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12569) );
  NAND4_X1 U15646 ( .A1(n12572), .A2(n12571), .A3(n12570), .A4(n12569), .ZN(
        n12573) );
  AOI211_X2 U15647 ( .C1(n17142), .C2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n12574), .B(n12573), .ZN(n12575) );
  NAND3_X2 U15648 ( .A1(n12577), .A2(n12576), .A3(n12575), .ZN(n18193) );
  AOI22_X1 U15649 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17142), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12582) );
  AOI22_X1 U15650 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12581) );
  INV_X2 U15651 ( .A(n12578), .ZN(n17143) );
  AOI22_X1 U15652 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12580) );
  AOI22_X1 U15653 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12579) );
  NAND4_X1 U15654 ( .A1(n12582), .A2(n12581), .A3(n12580), .A4(n12579), .ZN(
        n12588) );
  INV_X4 U15655 ( .A(n12742), .ZN(n17149) );
  AOI22_X1 U15656 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12586) );
  AOI22_X1 U15657 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U15658 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12584) );
  AOI22_X1 U15659 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12583) );
  NAND4_X1 U15660 ( .A1(n12586), .A2(n12585), .A3(n12584), .A4(n12583), .ZN(
        n12587) );
  AOI22_X1 U15661 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12592) );
  AOI22_X1 U15662 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U15663 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12590) );
  AOI22_X1 U15664 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12589) );
  NAND4_X1 U15665 ( .A1(n12592), .A2(n12591), .A3(n12590), .A4(n12589), .ZN(
        n12598) );
  AOI22_X1 U15666 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12596) );
  AOI22_X1 U15667 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12595) );
  AOI22_X1 U15668 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12594) );
  AOI22_X1 U15669 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12593) );
  NAND4_X1 U15670 ( .A1(n12596), .A2(n12595), .A3(n12594), .A4(n12593), .ZN(
        n12597) );
  NAND2_X1 U15671 ( .A1(n15862), .A2(n12652), .ZN(n18644) );
  AOI22_X1 U15672 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12604) );
  AOI22_X1 U15673 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12603) );
  AOI22_X1 U15674 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17142), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12602) );
  AOI22_X1 U15675 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12601) );
  NAND4_X1 U15676 ( .A1(n12604), .A2(n12603), .A3(n12602), .A4(n12601), .ZN(
        n12611) );
  INV_X2 U15677 ( .A(n12605), .ZN(n17127) );
  AOI22_X1 U15678 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17127), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12609) );
  AOI22_X1 U15679 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12608) );
  AOI22_X1 U15680 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12607) );
  AOI22_X1 U15681 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12606) );
  NAND4_X1 U15682 ( .A1(n12609), .A2(n12608), .A3(n12607), .A4(n12606), .ZN(
        n12610) );
  AOI22_X1 U15683 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n17127), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12618) );
  AOI22_X1 U15684 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n17147), .ZN(n12617) );
  AOI22_X1 U15685 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n14458), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17037), .ZN(n12612) );
  AOI22_X1 U15686 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17149), .ZN(n12616) );
  AOI22_X1 U15687 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17108), .ZN(n12615) );
  AOI22_X1 U15688 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n17125), .B1(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n15823), .ZN(n12614) );
  INV_X2 U15689 ( .A(n9604), .ZN(n17133) );
  AOI22_X1 U15690 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12613) );
  AOI22_X1 U15691 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17127), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12622) );
  AOI22_X1 U15692 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12621) );
  AOI22_X1 U15693 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17142), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12620) );
  AOI22_X1 U15694 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12619) );
  NAND4_X1 U15695 ( .A1(n12622), .A2(n12621), .A3(n12620), .A4(n12619), .ZN(
        n12628) );
  AOI22_X1 U15696 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12626) );
  AOI22_X1 U15697 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12625) );
  AOI22_X1 U15698 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12624) );
  AOI22_X1 U15699 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12623) );
  NAND4_X1 U15700 ( .A1(n12626), .A2(n12625), .A3(n12624), .A4(n12623), .ZN(
        n12627) );
  AOI22_X1 U15701 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12638) );
  AOI22_X1 U15702 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12637) );
  INV_X1 U15703 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17178) );
  AOI22_X1 U15704 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12629) );
  OAI21_X1 U15705 ( .B1(n12578), .B2(n17178), .A(n12629), .ZN(n12635) );
  AOI22_X1 U15706 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12633) );
  AOI22_X1 U15707 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17127), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12632) );
  AOI22_X1 U15708 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12631) );
  AOI22_X1 U15709 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12630) );
  NAND4_X1 U15710 ( .A1(n12633), .A2(n12632), .A3(n12631), .A4(n12630), .ZN(
        n12634) );
  NOR3_X1 U15711 ( .A1(n12671), .A2(n18215), .A3(n18644), .ZN(n14482) );
  AND2_X1 U15712 ( .A1(n18842), .A2(n14482), .ZN(n12650) );
  AOI22_X1 U15713 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12642) );
  AOI22_X1 U15714 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12641) );
  AOI22_X1 U15715 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12640) );
  AOI22_X1 U15716 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12639) );
  NAND4_X1 U15717 ( .A1(n12642), .A2(n12641), .A3(n12640), .A4(n12639), .ZN(
        n12648) );
  AOI22_X1 U15718 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12646) );
  AOI22_X1 U15719 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12645) );
  AOI22_X1 U15720 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17142), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12644) );
  AOI22_X1 U15721 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17127), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12643) );
  NAND4_X1 U15722 ( .A1(n12646), .A2(n12645), .A3(n12644), .A4(n12643), .ZN(
        n12647) );
  NAND2_X1 U15723 ( .A1(n12657), .A2(n12671), .ZN(n12662) );
  NAND2_X1 U15724 ( .A1(n12652), .A2(n12656), .ZN(n12649) );
  NAND2_X1 U15725 ( .A1(n12667), .A2(n18200), .ZN(n16537) );
  NOR3_X1 U15726 ( .A1(n18842), .A2(n12651), .A3(n13255), .ZN(n12665) );
  INV_X1 U15727 ( .A(n12652), .ZN(n18204) );
  NOR2_X1 U15728 ( .A1(n18193), .A2(n17353), .ZN(n12669) );
  OAI21_X1 U15729 ( .B1(n16928), .B2(n18632), .A(n12669), .ZN(n15843) );
  AOI21_X1 U15730 ( .B1(n12653), .B2(n15843), .A(n12652), .ZN(n12654) );
  INV_X1 U15731 ( .A(n12654), .ZN(n12655) );
  OAI21_X1 U15732 ( .B1(n12656), .B2(n18204), .A(n12655), .ZN(n12664) );
  AOI21_X1 U15733 ( .B1(n15862), .B2(n17353), .A(n18632), .ZN(n12663) );
  OR2_X1 U15734 ( .A1(n18200), .A2(n12670), .ZN(n12659) );
  AOI21_X1 U15735 ( .B1(n18225), .B2(n12661), .A(n12657), .ZN(n12658) );
  AOI21_X1 U15736 ( .B1(n12661), .B2(n12659), .A(n12658), .ZN(n12660) );
  OAI221_X1 U15737 ( .B1(n12663), .B2(n12662), .C1(n12663), .C2(n12661), .A(
        n12660), .ZN(n15844) );
  NOR3_X1 U15738 ( .A1(n12665), .A2(n12664), .A3(n15844), .ZN(n18643) );
  INV_X1 U15739 ( .A(n15844), .ZN(n12666) );
  NAND2_X1 U15740 ( .A1(n12667), .A2(n12666), .ZN(n13253) );
  NAND2_X1 U15741 ( .A1(n12671), .A2(n18207), .ZN(n18645) );
  OAI21_X1 U15742 ( .B1(n12675), .B2(n12674), .A(n12672), .ZN(n12673) );
  AOI21_X1 U15743 ( .B1(n12675), .B2(n12674), .A(n12673), .ZN(n13256) );
  AOI21_X1 U15744 ( .B1(n13256), .B2(n12676), .A(n13257), .ZN(n18624) );
  NAND2_X1 U15745 ( .A1(n15862), .A2(n18193), .ZN(n15872) );
  NAND2_X1 U15746 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18801), .ZN(n18690) );
  NAND2_X1 U15747 ( .A1(n18679), .A2(n18193), .ZN(n14483) );
  NOR2_X2 U15748 ( .A1(n18630), .A2(n14483), .ZN(n17833) );
  AOI22_X1 U15749 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15823), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12687) );
  AOI22_X1 U15750 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12686) );
  BUF_X1 U15751 ( .A(n17148), .Z(n17045) );
  AOI22_X1 U15752 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12678) );
  OAI21_X1 U15753 ( .B1(n9604), .B2(n20813), .A(n12678), .ZN(n12684) );
  AOI22_X1 U15754 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12682) );
  AOI22_X1 U15755 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12681) );
  AOI22_X1 U15756 ( .A1(n17127), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12680) );
  AOI22_X1 U15757 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12679) );
  NAND4_X1 U15758 ( .A1(n12682), .A2(n12681), .A3(n12680), .A4(n12679), .ZN(
        n12683) );
  AOI211_X1 U15759 ( .C1(n17045), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n12684), .B(n12683), .ZN(n12685) );
  AOI22_X1 U15760 ( .A1(n12716), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12701) );
  AOI22_X1 U15761 ( .A1(n15823), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12703), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12700) );
  AOI22_X1 U15762 ( .A1(n17147), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12718), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12688) );
  OAI21_X1 U15763 ( .B1(n12704), .B2(n20845), .A(n12688), .ZN(n12698) );
  AOI22_X1 U15764 ( .A1(n12677), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12696) );
  AOI22_X1 U15765 ( .A1(n12717), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12689), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12695) );
  AOI22_X1 U15766 ( .A1(n12691), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12690), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12694) );
  AOI22_X1 U15767 ( .A1(n12692), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17126), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12693) );
  NAND4_X1 U15768 ( .A1(n12696), .A2(n12695), .A3(n12694), .A4(n12693), .ZN(
        n12697) );
  INV_X1 U15769 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18802) );
  NOR2_X1 U15770 ( .A1(n12813), .A2(n18802), .ZN(n12714) );
  AOI22_X1 U15771 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12713) );
  AOI22_X1 U15772 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n15823), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12712) );
  INV_X1 U15773 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17146) );
  AOI22_X1 U15774 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12702) );
  OAI21_X1 U15775 ( .B1(n9604), .B2(n17146), .A(n12702), .ZN(n12710) );
  AOI22_X1 U15776 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12703), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12708) );
  AOI22_X1 U15777 ( .A1(n12689), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12707) );
  AOI22_X1 U15778 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12692), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12706) );
  AOI22_X1 U15779 ( .A1(n12718), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12705) );
  NAND4_X1 U15780 ( .A1(n12708), .A2(n12707), .A3(n12706), .A4(n12705), .ZN(
        n12709) );
  NAND3_X1 U15781 ( .A1(n12713), .A2(n12712), .A3(n12711), .ZN(n17842) );
  NAND2_X1 U15782 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17842), .ZN(
        n17841) );
  NOR2_X1 U15783 ( .A1(n17841), .A2(n17834), .ZN(n17832) );
  AOI22_X1 U15784 ( .A1(n12691), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12703), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12725) );
  AOI22_X1 U15785 ( .A1(n12689), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12692), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12724) );
  INV_X1 U15786 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17191) );
  AOI22_X1 U15787 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12715) );
  OAI21_X1 U15788 ( .B1(n9604), .B2(n17191), .A(n12715), .ZN(n12723) );
  AOI22_X1 U15789 ( .A1(n15823), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12722) );
  AOI22_X1 U15790 ( .A1(n12717), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12721) );
  AOI22_X1 U15791 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12720) );
  AOI22_X1 U15792 ( .A1(n12677), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12718), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12719) );
  XOR2_X1 U15793 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12726), .Z(
        n17824) );
  INV_X1 U15794 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18135) );
  NOR2_X1 U15795 ( .A1(n18135), .A2(n12726), .ZN(n12727) );
  INV_X1 U15796 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18118) );
  NAND2_X1 U15797 ( .A1(n12813), .A2(n12811), .ZN(n12740) );
  AOI22_X1 U15798 ( .A1(n15823), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12731) );
  AOI22_X1 U15799 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17127), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12730) );
  AOI22_X1 U15800 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12729) );
  AOI22_X1 U15801 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12728) );
  NAND4_X1 U15802 ( .A1(n12731), .A2(n12730), .A3(n12729), .A4(n12728), .ZN(
        n12737) );
  AOI22_X1 U15803 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12692), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12735) );
  AOI22_X1 U15804 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12734) );
  AOI22_X1 U15805 ( .A1(n12689), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12733) );
  AOI22_X1 U15806 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12703), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12732) );
  NAND4_X1 U15807 ( .A1(n12735), .A2(n12734), .A3(n12733), .A4(n12732), .ZN(
        n12736) );
  INV_X1 U15808 ( .A(n17335), .ZN(n12809) );
  XNOR2_X1 U15809 ( .A(n12740), .B(n12809), .ZN(n12738) );
  XOR2_X1 U15810 ( .A(n18118), .B(n12738), .Z(n17812) );
  AND2_X1 U15811 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12738), .ZN(
        n12739) );
  NOR2_X1 U15812 ( .A1(n17335), .A2(n12740), .ZN(n12752) );
  AOI22_X1 U15813 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12692), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U15814 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15823), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12750) );
  AOI22_X1 U15815 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12741) );
  OAI21_X1 U15816 ( .B1(n12742), .B2(n20795), .A(n12741), .ZN(n12748) );
  AOI22_X1 U15817 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12746) );
  AOI22_X1 U15818 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12745) );
  AOI22_X1 U15819 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12744) );
  AOI22_X1 U15820 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12743) );
  NAND4_X1 U15821 ( .A1(n12746), .A2(n12745), .A3(n12744), .A4(n12743), .ZN(
        n12747) );
  AOI211_X1 U15822 ( .C1(n17152), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n12748), .B(n12747), .ZN(n12749) );
  NAND3_X1 U15823 ( .A1(n12751), .A2(n12750), .A3(n12749), .ZN(n12804) );
  XNOR2_X1 U15824 ( .A(n12752), .B(n12804), .ZN(n17801) );
  NAND2_X1 U15825 ( .A1(n12752), .A2(n12804), .ZN(n12763) );
  AOI22_X1 U15826 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U15827 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U15828 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12754) );
  AOI22_X1 U15829 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12753) );
  NAND4_X1 U15830 ( .A1(n12756), .A2(n12755), .A3(n12754), .A4(n12753), .ZN(
        n12762) );
  AOI22_X1 U15831 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U15832 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12759) );
  AOI22_X1 U15833 ( .A1(n15823), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12758) );
  AOI22_X1 U15834 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12757) );
  NAND4_X1 U15835 ( .A1(n12760), .A2(n12759), .A3(n12758), .A4(n12757), .ZN(
        n12761) );
  XNOR2_X1 U15836 ( .A(n12763), .B(n17328), .ZN(n17785) );
  NAND2_X1 U15837 ( .A1(n17783), .A2(n17785), .ZN(n17784) );
  INV_X1 U15838 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18095) );
  AOI22_X1 U15839 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12773) );
  AOI22_X1 U15840 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12772) );
  INV_X1 U15841 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17174) );
  AOI22_X1 U15842 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12764) );
  OAI21_X1 U15843 ( .B1(n9604), .B2(n17174), .A(n12764), .ZN(n12770) );
  AOI22_X1 U15844 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12768) );
  AOI22_X1 U15845 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12767) );
  AOI22_X1 U15846 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12766) );
  AOI22_X1 U15847 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12765) );
  NAND4_X1 U15848 ( .A1(n12768), .A2(n12767), .A3(n12766), .A4(n12765), .ZN(
        n12769) );
  AOI211_X1 U15849 ( .C1(n17152), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n12770), .B(n12769), .ZN(n12771) );
  NAND3_X1 U15850 ( .A1(n12773), .A2(n12772), .A3(n12771), .ZN(n12803) );
  XOR2_X1 U15851 ( .A(n12776), .B(n12803), .Z(n12774) );
  XOR2_X1 U15852 ( .A(n18095), .B(n12774), .Z(n17774) );
  OAI21_X1 U15853 ( .B1(n12777), .B2(n15879), .A(n17743), .ZN(n12778) );
  XNOR2_X1 U15854 ( .A(n12779), .B(n12778), .ZN(n17765) );
  INV_X1 U15855 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18094) );
  INV_X1 U15856 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18005) );
  INV_X1 U15857 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17650) );
  NAND4_X1 U15858 ( .A1(n18005), .A2(n18042), .A3(n18000), .A4(n17650), .ZN(
        n12782) );
  NOR2_X1 U15859 ( .A1(n12781), .A2(n12780), .ZN(n18051) );
  NAND2_X1 U15860 ( .A1(n18051), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18036) );
  NOR2_X1 U15861 ( .A1(n18036), .A2(n18042), .ZN(n17670) );
  NOR3_X1 U15862 ( .A1(n18005), .A2(n18003), .A3(n18000), .ZN(n17987) );
  NAND2_X1 U15863 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17987), .ZN(
        n17969) );
  NAND2_X1 U15864 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n12784), .ZN(
        n17624) );
  NAND2_X1 U15865 ( .A1(n17850), .A2(n17671), .ZN(n12790) );
  NAND2_X1 U15866 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17609) );
  NAND2_X1 U15867 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17921) );
  INV_X1 U15868 ( .A(n17921), .ZN(n17937) );
  NAND3_X1 U15869 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n17937), .ZN(n17911) );
  INV_X1 U15870 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17929) );
  NOR2_X1 U15871 ( .A1(n17911), .A2(n17929), .ZN(n17878) );
  INV_X1 U15872 ( .A(n17878), .ZN(n17867) );
  NOR2_X1 U15873 ( .A1(n17609), .A2(n17867), .ZN(n15876) );
  INV_X1 U15874 ( .A(n15876), .ZN(n12786) );
  INV_X1 U15875 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17898) );
  NOR2_X1 U15876 ( .A1(n12786), .A2(n17898), .ZN(n12837) );
  INV_X1 U15877 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n20876) );
  NAND2_X1 U15878 ( .A1(n17606), .A2(n20876), .ZN(n12787) );
  NOR2_X1 U15879 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n12787), .ZN(
        n17569) );
  INV_X1 U15880 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17932) );
  NAND2_X1 U15881 ( .A1(n17569), .A2(n17932), .ZN(n17556) );
  NOR3_X1 U15882 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17556), .ZN(n12788) );
  INV_X1 U15883 ( .A(n12789), .ZN(n12794) );
  INV_X1 U15884 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17982) );
  AOI22_X1 U15885 ( .A1(n12790), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n17982), .B2(n17627), .ZN(n12791) );
  INV_X1 U15886 ( .A(n12791), .ZN(n12792) );
  INV_X1 U15887 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17964) );
  NAND2_X1 U15888 ( .A1(n17619), .A2(n17964), .ZN(n17618) );
  INV_X1 U15889 ( .A(n17609), .ZN(n17963) );
  NAND2_X1 U15890 ( .A1(n17963), .A2(n17626), .ZN(n17567) );
  NAND2_X1 U15891 ( .A1(n17536), .A2(n17567), .ZN(n17568) );
  NAND2_X1 U15892 ( .A1(n17878), .A2(n17568), .ZN(n17537) );
  INV_X1 U15893 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17880) );
  NAND2_X1 U15894 ( .A1(n17743), .A2(n17521), .ZN(n12795) );
  OAI211_X1 U15895 ( .C1(n12796), .C2(n17880), .A(n12795), .B(n10138), .ZN(
        n17499) );
  NOR2_X1 U15896 ( .A1(n12796), .A2(n17743), .ZN(n17520) );
  INV_X1 U15897 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17875) );
  NOR2_X1 U15898 ( .A1(n17880), .A2(n17875), .ZN(n12838) );
  INV_X1 U15899 ( .A(n12838), .ZN(n17854) );
  AND2_X1 U15900 ( .A1(n17627), .A2(n17854), .ZN(n12797) );
  NOR2_X2 U15901 ( .A1(n17498), .A2(n12798), .ZN(n12800) );
  INV_X1 U15902 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17476) );
  NAND2_X1 U15903 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16431) );
  NOR2_X1 U15904 ( .A1(n16431), .A2(n12799), .ZN(n15950) );
  INV_X1 U15905 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n20799) );
  NAND2_X1 U15906 ( .A1(n15950), .A2(n20799), .ZN(n15953) );
  INV_X1 U15907 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17535) );
  NOR2_X1 U15908 ( .A1(n17898), .A2(n17535), .ZN(n17879) );
  INV_X1 U15909 ( .A(n17879), .ZN(n17876) );
  NOR2_X1 U15910 ( .A1(n17854), .A2(n17876), .ZN(n17849) );
  INV_X1 U15911 ( .A(n12803), .ZN(n17325) );
  INV_X1 U15912 ( .A(n12804), .ZN(n17331) );
  INV_X1 U15913 ( .A(n12811), .ZN(n17340) );
  NAND2_X1 U15914 ( .A1(n12813), .A2(n17842), .ZN(n12810) );
  NAND2_X1 U15915 ( .A1(n17340), .A2(n12810), .ZN(n12808) );
  NAND2_X1 U15916 ( .A1(n12809), .A2(n12808), .ZN(n12821) );
  INV_X1 U15917 ( .A(n17328), .ZN(n12806) );
  NAND2_X1 U15918 ( .A1(n12805), .A2(n12806), .ZN(n12824) );
  NOR2_X1 U15919 ( .A1(n17325), .A2(n12824), .ZN(n12828) );
  NAND2_X1 U15920 ( .A1(n12828), .A2(n15879), .ZN(n12829) );
  XOR2_X1 U15921 ( .A(n12806), .B(n12805), .Z(n12807) );
  AND2_X1 U15922 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n12807), .ZN(
        n12823) );
  INV_X1 U15923 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17786) );
  XOR2_X1 U15924 ( .A(n17786), .B(n12807), .Z(n17790) );
  XOR2_X1 U15925 ( .A(n12809), .B(n12808), .Z(n12819) );
  AND2_X1 U15926 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12819), .ZN(
        n12820) );
  XNOR2_X1 U15927 ( .A(n12811), .B(n12810), .ZN(n12812) );
  NOR2_X1 U15928 ( .A1(n12812), .A2(n18135), .ZN(n12818) );
  XOR2_X1 U15929 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12812), .Z(
        n17826) );
  INV_X1 U15930 ( .A(n12813), .ZN(n17351) );
  INV_X1 U15931 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18818) );
  NOR2_X1 U15932 ( .A1(n17351), .A2(n18818), .ZN(n12816) );
  INV_X1 U15933 ( .A(n17842), .ZN(n12815) );
  NAND3_X1 U15934 ( .A1(n12815), .A2(n17351), .A3(n18818), .ZN(n12814) );
  OAI221_X1 U15935 ( .B1(n12816), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n12815), .C2(n17351), .A(n12814), .ZN(n17825) );
  NOR2_X1 U15936 ( .A1(n17826), .A2(n17825), .ZN(n12817) );
  NOR2_X1 U15937 ( .A1(n12818), .A2(n12817), .ZN(n17816) );
  XOR2_X1 U15938 ( .A(n18118), .B(n12819), .Z(n17815) );
  NOR2_X1 U15939 ( .A1(n17816), .A2(n17815), .ZN(n17814) );
  NOR2_X1 U15940 ( .A1(n12820), .A2(n17814), .ZN(n17797) );
  XNOR2_X1 U15941 ( .A(n17331), .B(n12821), .ZN(n17798) );
  NOR2_X1 U15942 ( .A1(n17797), .A2(n17798), .ZN(n12822) );
  NAND2_X1 U15943 ( .A1(n17797), .A2(n17798), .ZN(n17796) );
  OAI21_X1 U15944 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n12822), .A(
        n17796), .ZN(n17789) );
  NOR2_X1 U15945 ( .A1(n17790), .A2(n17789), .ZN(n17788) );
  XNOR2_X1 U15946 ( .A(n17325), .B(n12824), .ZN(n12826) );
  NOR2_X1 U15947 ( .A1(n12825), .A2(n12826), .ZN(n12827) );
  XNOR2_X1 U15948 ( .A(n12826), .B(n12825), .ZN(n17770) );
  NOR2_X1 U15949 ( .A1(n12827), .A2(n17769), .ZN(n12830) );
  XOR2_X1 U15950 ( .A(n17321), .B(n12828), .Z(n12831) );
  NAND2_X1 U15951 ( .A1(n12830), .A2(n12831), .ZN(n17757) );
  NAND2_X1 U15952 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17757), .ZN(
        n12833) );
  NOR2_X1 U15953 ( .A1(n12829), .A2(n12833), .ZN(n12835) );
  INV_X1 U15954 ( .A(n12829), .ZN(n12834) );
  OR2_X1 U15955 ( .A1(n12831), .A2(n12830), .ZN(n17758) );
  OAI21_X1 U15956 ( .B1(n12834), .B2(n12833), .A(n17758), .ZN(n12832) );
  AOI21_X1 U15957 ( .B1(n12834), .B2(n12833), .A(n12832), .ZN(n17752) );
  INV_X1 U15958 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n20851) );
  NAND2_X1 U15959 ( .A1(n17321), .A2(n17833), .ZN(n17685) );
  INV_X2 U15960 ( .A(n17685), .ZN(n17753) );
  NAND2_X1 U15961 ( .A1(n15876), .A2(n17620), .ZN(n17548) );
  INV_X1 U15962 ( .A(n17548), .ZN(n17506) );
  NAND2_X1 U15963 ( .A1(n17849), .A2(n17506), .ZN(n17491) );
  OAI22_X1 U15964 ( .A1(n17756), .A2(n15952), .B1(n15953), .B2(n17491), .ZN(
        n12836) );
  INV_X1 U15965 ( .A(n12836), .ZN(n12847) );
  NAND2_X1 U15966 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17664), .ZN(
        n17663) );
  NAND2_X1 U15967 ( .A1(n17913), .A2(n12837), .ZN(n17893) );
  NAND2_X1 U15968 ( .A1(n17519), .A2(n12838), .ZN(n17858) );
  NAND2_X1 U15969 ( .A1(n17475), .A2(n15950), .ZN(n16391) );
  NAND2_X1 U15970 ( .A1(n17753), .A2(n16391), .ZN(n16405) );
  NAND2_X1 U15971 ( .A1(n18044), .A2(n17850), .ZN(n17914) );
  NAND2_X1 U15972 ( .A1(n12838), .A2(n17510), .ZN(n16430) );
  NAND2_X1 U15973 ( .A1(n15950), .A2(n17860), .ZN(n16393) );
  NAND2_X1 U15974 ( .A1(n17837), .A2(n16393), .ZN(n16411) );
  NAND2_X1 U15975 ( .A1(n16405), .A2(n16411), .ZN(n12845) );
  INV_X1 U15976 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17612) );
  NAND2_X1 U15977 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17804) );
  NAND2_X1 U15978 ( .A1(n17782), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17772) );
  NAND2_X1 U15979 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17745) );
  INV_X1 U15980 ( .A(n17745), .ZN(n17732) );
  NAND2_X1 U15981 ( .A1(n17732), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17730) );
  INV_X1 U15982 ( .A(n17730), .ZN(n17716) );
  NAND2_X1 U15983 ( .A1(n17716), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16772) );
  INV_X1 U15984 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17691) );
  NOR2_X1 U15985 ( .A1(n17691), .A2(n16751), .ZN(n17656) );
  INV_X1 U15986 ( .A(n17656), .ZN(n17680) );
  NAND3_X1 U15987 ( .A1(n17551), .A2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17543) );
  INV_X1 U15988 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17514) );
  NAND2_X1 U15989 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16561) );
  INV_X1 U15990 ( .A(n16561), .ZN(n17511) );
  INV_X1 U15991 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17470) );
  INV_X1 U15992 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17471) );
  NAND2_X1 U15993 ( .A1(n15851), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17844) );
  AOI21_X1 U15994 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18838)
         );
  NOR2_X1 U15995 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18845) );
  INV_X1 U15996 ( .A(n18845), .ZN(n12839) );
  NAND2_X1 U15997 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n18173) );
  NAND3_X1 U15998 ( .A1(n18688), .A2(n18794), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18532) );
  AOI21_X1 U15999 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17577), .A(
        n18568), .ZN(n17679) );
  OR2_X1 U16000 ( .A1(n12841), .A2(n17679), .ZN(n16389) );
  INV_X1 U16001 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16582) );
  NOR2_X1 U16002 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17500), .ZN(
        n16400) );
  NAND2_X1 U16003 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16397), .ZN(
        n16399) );
  INV_X1 U16004 ( .A(n16399), .ZN(n16559) );
  NAND2_X1 U16005 ( .A1(n18568), .A2(n12841), .ZN(n16403) );
  OAI211_X1 U16006 ( .C1(n16559), .C2(n17844), .A(n17843), .B(n16403), .ZN(
        n16408) );
  NOR2_X1 U16007 ( .A1(n16400), .A2(n16408), .ZN(n16387) );
  NAND2_X1 U16008 ( .A1(n18801), .A2(n18794), .ZN(n18853) );
  INV_X1 U16009 ( .A(n18853), .ZN(n18817) );
  NAND3_X2 U16010 ( .A1(n18817), .A2(n18688), .A3(n15851), .ZN(n18122) );
  NAND2_X1 U16011 ( .A1(n18153), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n12840) );
  OAI221_X1 U16012 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16389), .C1(
        n16582), .C2(n16387), .A(n12840), .ZN(n12843) );
  INV_X1 U16013 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18841) );
  INV_X1 U16014 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16912) );
  XNOR2_X1 U16015 ( .A(n16582), .B(n16398), .ZN(n16581) );
  NAND2_X1 U16016 ( .A1(n12848), .A2(n19121), .ZN(n12858) );
  OAI21_X1 U16017 ( .B1(n12849), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n12850), .ZN(n15189) );
  INV_X1 U16018 ( .A(n15189), .ZN(n13215) );
  OAI21_X1 U16019 ( .B1(n16265), .B2(n9928), .A(n12851), .ZN(n12853) );
  NOR2_X1 U16020 ( .A1(n15287), .A2(n16247), .ZN(n12852) );
  AOI211_X1 U16021 ( .C1(n16255), .C2(n13215), .A(n12853), .B(n12852), .ZN(
        n12854) );
  NAND2_X1 U16022 ( .A1(n12858), .A2(n12857), .ZN(P2_U2986) );
  INV_X1 U16023 ( .A(n12869), .ZN(n12859) );
  NAND2_X1 U16024 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19482) );
  NAND2_X1 U16025 ( .A1(n19482), .A2(n19813), .ZN(n12861) );
  NOR2_X1 U16026 ( .A1(n19813), .A2(n19822), .ZN(n19612) );
  NAND2_X1 U16027 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19612), .ZN(
        n14268) );
  AND2_X1 U16028 ( .A1(n12861), .A2(n14268), .ZN(n19264) );
  AOI22_X1 U16029 ( .A1(n12873), .A2(n16322), .B1(n19793), .B2(n19264), .ZN(
        n12862) );
  NAND3_X1 U16030 ( .A1(n13298), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13297), 
        .ZN(n12884) );
  INV_X1 U16031 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12863) );
  NOR2_X1 U16032 ( .A1(n12884), .A2(n12863), .ZN(n12864) );
  XNOR2_X1 U16033 ( .A(n19822), .B(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19265) );
  AND2_X1 U16034 ( .A1(n19265), .A2(n19793), .ZN(n19450) );
  AOI21_X1 U16035 ( .B1(n12873), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19450), .ZN(n12865) );
  AOI22_X1 U16036 ( .A1(n12873), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19793), .B2(n19828), .ZN(n12866) );
  NAND2_X1 U16037 ( .A1(n19612), .A2(n19803), .ZN(n19328) );
  INV_X1 U16038 ( .A(n19328), .ZN(n19361) );
  NAND2_X1 U16039 ( .A1(n14268), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12871) );
  NAND2_X1 U16040 ( .A1(n19392), .A2(n12871), .ZN(n12872) );
  AND2_X1 U16041 ( .A1(n12872), .A2(n19793), .ZN(n19540) );
  AOI21_X1 U16042 ( .B1(n12873), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19540), .ZN(n12874) );
  INV_X1 U16043 ( .A(n12881), .ZN(n12876) );
  INV_X1 U16044 ( .A(n12884), .ZN(n13087) );
  NAND2_X1 U16045 ( .A1(n13087), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12877) );
  NAND2_X1 U16046 ( .A1(n12876), .A2(n12877), .ZN(n12879) );
  INV_X1 U16047 ( .A(n12877), .ZN(n12878) );
  NAND2_X1 U16048 ( .A1(n13538), .A2(n13539), .ZN(n13537) );
  NAND2_X1 U16049 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n10214), .ZN(
        n12880) );
  NAND2_X1 U16050 ( .A1(n13537), .A2(n12880), .ZN(n13577) );
  AND2_X1 U16051 ( .A1(n13609), .A2(n13732), .ZN(n12887) );
  AND2_X1 U16052 ( .A1(n13722), .A2(n13721), .ZN(n12886) );
  NAND2_X1 U16053 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12882) );
  NOR2_X1 U16054 ( .A1(n12882), .A2(n14295), .ZN(n12885) );
  INV_X1 U16055 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12883) );
  NOR2_X1 U16056 ( .A1(n12884), .A2(n12883), .ZN(n13580) );
  AND2_X1 U16057 ( .A1(n12885), .A2(n13580), .ZN(n13571) );
  NAND2_X1 U16058 ( .A1(n9686), .A2(n13955), .ZN(n13953) );
  INV_X1 U16059 ( .A(n13953), .ZN(n12903) );
  AOI22_X1 U16060 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12892) );
  AOI22_X1 U16061 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12891) );
  AOI22_X1 U16062 ( .A1(n10410), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12890) );
  AOI22_X1 U16063 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12889) );
  NAND4_X1 U16064 ( .A1(n12892), .A2(n12891), .A3(n12890), .A4(n12889), .ZN(
        n12901) );
  AOI22_X1 U16065 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10503), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12899) );
  INV_X1 U16066 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12895) );
  NAND2_X1 U16067 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12894) );
  AOI22_X1 U16068 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12982), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12893) );
  OAI211_X1 U16069 ( .C1(n12987), .C2(n12895), .A(n12894), .B(n12893), .ZN(
        n12896) );
  INV_X1 U16070 ( .A(n12896), .ZN(n12898) );
  AOI22_X1 U16071 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12897) );
  NAND3_X1 U16072 ( .A1(n12899), .A2(n12898), .A3(n12897), .ZN(n12900) );
  NOR2_X1 U16073 ( .A1(n12901), .A2(n12900), .ZN(n14069) );
  INV_X1 U16074 ( .A(n14069), .ZN(n12902) );
  AOI22_X1 U16075 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12907) );
  AOI22_X1 U16076 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12906) );
  AOI22_X1 U16077 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n10410), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12905) );
  AOI22_X1 U16078 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10516), .B1(
        n10445), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12904) );
  NAND4_X1 U16079 ( .A1(n12907), .A2(n12906), .A3(n12905), .A4(n12904), .ZN(
        n12916) );
  AOI22_X1 U16080 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10503), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12914) );
  INV_X1 U16081 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12910) );
  NAND2_X1 U16082 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12909) );
  AOI22_X1 U16083 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n12982), .ZN(n12908) );
  OAI211_X1 U16084 ( .C1(n12987), .C2(n12910), .A(n12909), .B(n12908), .ZN(
        n12911) );
  INV_X1 U16085 ( .A(n12911), .ZN(n12913) );
  AOI22_X1 U16086 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n10434), .ZN(n12912) );
  NAND3_X1 U16087 ( .A1(n12914), .A2(n12913), .A3(n12912), .ZN(n12915) );
  AOI22_X1 U16088 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10503), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12923) );
  INV_X1 U16089 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12919) );
  NAND2_X1 U16090 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12918) );
  AOI22_X1 U16091 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n12982), .ZN(n12917) );
  OAI211_X1 U16092 ( .C1(n12987), .C2(n12919), .A(n12918), .B(n12917), .ZN(
        n12920) );
  INV_X1 U16093 ( .A(n12920), .ZN(n12922) );
  AOI22_X1 U16094 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__2__SCAN_IN), .B2(n10434), .ZN(n12921) );
  NAND3_X1 U16095 ( .A1(n12923), .A2(n12922), .A3(n12921), .ZN(n12929) );
  AOI22_X1 U16096 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12927) );
  AOI22_X1 U16097 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12926) );
  AOI22_X1 U16098 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n10410), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12925) );
  AOI22_X1 U16099 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10516), .B1(
        n10445), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12924) );
  NAND4_X1 U16100 ( .A1(n12927), .A2(n12926), .A3(n12925), .A4(n12924), .ZN(
        n12928) );
  AOI22_X1 U16101 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10503), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12936) );
  INV_X1 U16102 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12932) );
  NAND2_X1 U16103 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12931) );
  AOI22_X1 U16104 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n12982), .ZN(n12930) );
  OAI211_X1 U16105 ( .C1(n12987), .C2(n12932), .A(n12931), .B(n12930), .ZN(
        n12933) );
  INV_X1 U16106 ( .A(n12933), .ZN(n12935) );
  AOI22_X1 U16107 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__3__SCAN_IN), .B2(n10434), .ZN(n12934) );
  NAND3_X1 U16108 ( .A1(n12936), .A2(n12935), .A3(n12934), .ZN(n12942) );
  AOI22_X1 U16109 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12940) );
  AOI22_X1 U16110 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12939) );
  AOI22_X1 U16111 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n10410), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12938) );
  AOI22_X1 U16112 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10516), .B1(
        n10445), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12937) );
  NAND4_X1 U16113 ( .A1(n12940), .A2(n12939), .A3(n12938), .A4(n12937), .ZN(
        n12941) );
  AOI22_X1 U16114 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10503), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12949) );
  INV_X1 U16115 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12945) );
  NAND2_X1 U16116 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12944) );
  AOI22_X1 U16117 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n12982), .ZN(n12943) );
  OAI211_X1 U16118 ( .C1(n12987), .C2(n12945), .A(n12944), .B(n12943), .ZN(
        n12946) );
  INV_X1 U16119 ( .A(n12946), .ZN(n12948) );
  AOI22_X1 U16120 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__4__SCAN_IN), .B2(n10434), .ZN(n12947) );
  NAND3_X1 U16121 ( .A1(n12949), .A2(n12948), .A3(n12947), .ZN(n12955) );
  AOI22_X1 U16122 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12953) );
  AOI22_X1 U16123 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12952) );
  AOI22_X1 U16124 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n10410), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12951) );
  AOI22_X1 U16125 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10516), .B1(
        n10445), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12950) );
  NAND4_X1 U16126 ( .A1(n12953), .A2(n12952), .A3(n12951), .A4(n12950), .ZN(
        n12954) );
  NAND2_X1 U16127 ( .A1(n15339), .A2(n15340), .ZN(n15331) );
  AOI22_X1 U16128 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12959) );
  AOI22_X1 U16129 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12958) );
  AOI22_X1 U16130 ( .A1(n10410), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12957) );
  AOI22_X1 U16131 ( .A1(n10445), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10516), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12956) );
  NAND4_X1 U16132 ( .A1(n12959), .A2(n12958), .A3(n12957), .A4(n12956), .ZN(
        n12968) );
  AOI22_X1 U16133 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10503), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12966) );
  INV_X1 U16134 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12962) );
  NAND2_X1 U16135 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12961) );
  AOI22_X1 U16136 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12982), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12960) );
  OAI211_X1 U16137 ( .C1(n12987), .C2(n12962), .A(n12961), .B(n12960), .ZN(
        n12963) );
  INV_X1 U16138 ( .A(n12963), .ZN(n12965) );
  AOI22_X1 U16139 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10434), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12964) );
  NAND3_X1 U16140 ( .A1(n12966), .A2(n12965), .A3(n12964), .ZN(n12967) );
  NAND2_X1 U16141 ( .A1(n15332), .A2(n10137), .ZN(n15323) );
  AOI22_X1 U16142 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12972) );
  AOI22_X1 U16143 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12971) );
  AOI22_X1 U16144 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10410), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12970) );
  AOI22_X1 U16145 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n10516), .B1(
        n10445), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12969) );
  NAND4_X1 U16146 ( .A1(n12972), .A2(n12971), .A3(n12970), .A4(n12969), .ZN(
        n12981) );
  AOI22_X1 U16147 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10503), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12979) );
  INV_X1 U16148 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12975) );
  NAND2_X1 U16149 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12974) );
  AOI22_X1 U16150 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n12982), .ZN(n12973) );
  OAI211_X1 U16151 ( .C1(n12987), .C2(n12975), .A(n12974), .B(n12973), .ZN(
        n12976) );
  INV_X1 U16152 ( .A(n12976), .ZN(n12978) );
  AOI22_X1 U16153 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__6__SCAN_IN), .B2(n10434), .ZN(n12977) );
  NAND3_X1 U16154 ( .A1(n12979), .A2(n12978), .A3(n12977), .ZN(n12980) );
  NOR2_X1 U16155 ( .A1(n12981), .A2(n12980), .ZN(n15325) );
  AOI22_X1 U16156 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10491), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12991) );
  AOI22_X1 U16157 ( .A1(n10411), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10427), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12990) );
  INV_X1 U16158 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12986) );
  NAND2_X1 U16159 ( .A1(n10418), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12985) );
  AOI22_X1 U16160 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n12982), .ZN(n12984) );
  OAI211_X1 U16161 ( .C1(n12987), .C2(n12986), .A(n12985), .B(n12984), .ZN(
        n12988) );
  INV_X1 U16162 ( .A(n12988), .ZN(n12989) );
  NAND3_X1 U16163 ( .A1(n12991), .A2(n12990), .A3(n12989), .ZN(n12997) );
  AOI22_X1 U16164 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10503), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12995) );
  AOI22_X1 U16165 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n10434), .ZN(n12994) );
  AOI22_X1 U16166 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n10410), .B1(
        n10440), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12993) );
  AOI22_X1 U16167 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10516), .B1(
        n10445), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12992) );
  NAND4_X1 U16168 ( .A1(n12995), .A2(n12994), .A3(n12993), .A4(n12992), .ZN(
        n12996) );
  OR2_X1 U16169 ( .A1(n12997), .A2(n12996), .ZN(n13019) );
  NAND2_X1 U16170 ( .A1(n13133), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n13001) );
  NAND2_X1 U16171 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n13000) );
  NAND2_X1 U16172 ( .A1(n10375), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12999) );
  NAND2_X1 U16173 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12998) );
  AND4_X1 U16174 ( .A1(n13001), .A2(n13000), .A3(n12999), .A4(n12998), .ZN(
        n13005) );
  AOI22_X1 U16175 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13004) );
  INV_X1 U16176 ( .A(n13002), .ZN(n15802) );
  INV_X1 U16177 ( .A(n15802), .ZN(n13137) );
  AOI22_X1 U16178 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13003) );
  XNOR2_X1 U16179 ( .A(n16322), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13134) );
  NAND4_X1 U16180 ( .A1(n13005), .A2(n13004), .A3(n13003), .A4(n13134), .ZN(
        n13014) );
  NAND2_X1 U16181 ( .A1(n13133), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13009) );
  NAND2_X1 U16182 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13008) );
  NAND2_X1 U16183 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n13007) );
  NAND2_X1 U16184 ( .A1(n10375), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13006) );
  AND4_X1 U16185 ( .A1(n13009), .A2(n13008), .A3(n13007), .A4(n13006), .ZN(
        n13012) );
  INV_X1 U16186 ( .A(n13134), .ZN(n13131) );
  AOI22_X1 U16187 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13011) );
  AOI22_X1 U16188 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10235), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13010) );
  NAND4_X1 U16189 ( .A1(n13012), .A2(n13131), .A3(n13011), .A4(n13010), .ZN(
        n13013) );
  NAND2_X1 U16190 ( .A1(n13014), .A2(n13013), .ZN(n13035) );
  NOR2_X1 U16191 ( .A1(n10364), .A2(n13035), .ZN(n13015) );
  XOR2_X1 U16192 ( .A(n13019), .B(n13015), .Z(n13033) );
  INV_X1 U16193 ( .A(n13035), .ZN(n13018) );
  NAND2_X1 U16194 ( .A1(n10364), .A2(n13018), .ZN(n15320) );
  NAND2_X1 U16195 ( .A1(n13019), .A2(n13018), .ZN(n13038) );
  AOI22_X1 U16196 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10235), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13021) );
  AOI22_X1 U16197 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13020) );
  AND2_X1 U16198 ( .A1(n13021), .A2(n13020), .ZN(n13024) );
  AOI22_X1 U16199 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13023) );
  AOI22_X1 U16200 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13022) );
  NAND4_X1 U16201 ( .A1(n13024), .A2(n13023), .A3(n13022), .A4(n13134), .ZN(
        n13031) );
  AOI22_X1 U16202 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10235), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13026) );
  AOI22_X1 U16203 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13025) );
  AND2_X1 U16204 ( .A1(n13026), .A2(n13025), .ZN(n13029) );
  AOI22_X1 U16205 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13028) );
  AOI22_X1 U16206 ( .A1(n13129), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13027) );
  NAND4_X1 U16207 ( .A1(n13029), .A2(n13131), .A3(n13028), .A4(n13027), .ZN(
        n13030) );
  NAND2_X1 U16208 ( .A1(n13031), .A2(n13030), .ZN(n13037) );
  XOR2_X1 U16209 ( .A(n13038), .B(n13037), .Z(n13032) );
  NAND2_X1 U16210 ( .A1(n13032), .A2(n13087), .ZN(n15306) );
  INV_X1 U16211 ( .A(n13037), .ZN(n13034) );
  NAND2_X1 U16212 ( .A1(n10383), .A2(n13034), .ZN(n15307) );
  NOR2_X1 U16213 ( .A1(n13038), .A2(n13037), .ZN(n13051) );
  AOI22_X1 U16214 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13040) );
  AOI22_X1 U16215 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13039) );
  AND2_X1 U16216 ( .A1(n13040), .A2(n13039), .ZN(n13043) );
  AOI22_X1 U16217 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13042) );
  AOI22_X1 U16218 ( .A1(n13129), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13041) );
  NAND4_X1 U16219 ( .A1(n13043), .A2(n13042), .A3(n13041), .A4(n13134), .ZN(
        n13050) );
  AOI22_X1 U16220 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13045) );
  AOI22_X1 U16221 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13044) );
  AND2_X1 U16222 ( .A1(n13045), .A2(n13044), .ZN(n13048) );
  AOI22_X1 U16223 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13047) );
  AOI22_X1 U16224 ( .A1(n13129), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13046) );
  NAND4_X1 U16225 ( .A1(n13048), .A2(n13131), .A3(n13047), .A4(n13046), .ZN(
        n13049) );
  AND2_X1 U16226 ( .A1(n13050), .A2(n13049), .ZN(n13053) );
  NAND2_X1 U16227 ( .A1(n13051), .A2(n13053), .ZN(n13084) );
  OAI211_X1 U16228 ( .C1(n13051), .C2(n13053), .A(n13084), .B(n13087), .ZN(
        n13056) );
  INV_X1 U16229 ( .A(n13056), .ZN(n13052) );
  XNOR2_X1 U16230 ( .A(n13055), .B(n13052), .ZN(n15298) );
  INV_X1 U16231 ( .A(n13053), .ZN(n13054) );
  NOR2_X1 U16232 ( .A1(n9600), .A2(n13054), .ZN(n15300) );
  NAND2_X1 U16233 ( .A1(n15298), .A2(n15300), .ZN(n15299) );
  AOI22_X1 U16234 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9586), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13058) );
  AOI22_X1 U16235 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13057) );
  AND2_X1 U16236 ( .A1(n13058), .A2(n13057), .ZN(n13061) );
  AOI22_X1 U16237 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13060) );
  AOI22_X1 U16238 ( .A1(n13129), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13059) );
  NAND4_X1 U16239 ( .A1(n13061), .A2(n13060), .A3(n13059), .A4(n13134), .ZN(
        n13068) );
  AOI22_X1 U16240 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13063) );
  AOI22_X1 U16241 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13062) );
  AND2_X1 U16242 ( .A1(n13063), .A2(n13062), .ZN(n13066) );
  AOI22_X1 U16243 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13065) );
  AOI22_X1 U16244 ( .A1(n13129), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13064) );
  NAND4_X1 U16245 ( .A1(n13066), .A2(n13131), .A3(n13065), .A4(n13064), .ZN(
        n13067) );
  AND2_X1 U16246 ( .A1(n13068), .A2(n13067), .ZN(n13085) );
  XNOR2_X1 U16247 ( .A(n13084), .B(n13085), .ZN(n13069) );
  NAND2_X1 U16248 ( .A1(n10364), .A2(n13085), .ZN(n15295) );
  INV_X1 U16249 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n20803) );
  AOI22_X1 U16250 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13073) );
  AOI22_X1 U16251 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13072) );
  AND2_X1 U16252 ( .A1(n13073), .A2(n13072), .ZN(n13076) );
  AOI22_X1 U16253 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13075) );
  AOI22_X1 U16254 ( .A1(n13129), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13074) );
  NAND4_X1 U16255 ( .A1(n13076), .A2(n13075), .A3(n13074), .A4(n13134), .ZN(
        n13083) );
  AOI22_X1 U16256 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10235), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13078) );
  AOI22_X1 U16257 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13077) );
  AND2_X1 U16258 ( .A1(n13078), .A2(n13077), .ZN(n13081) );
  AOI22_X1 U16259 ( .A1(n13133), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13080) );
  AOI22_X1 U16260 ( .A1(n13129), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9590), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13079) );
  NAND4_X1 U16261 ( .A1(n13081), .A2(n13131), .A3(n13080), .A4(n13079), .ZN(
        n13082) );
  AND2_X1 U16262 ( .A1(n13083), .A2(n13082), .ZN(n13090) );
  INV_X1 U16263 ( .A(n13084), .ZN(n13086) );
  NAND2_X1 U16264 ( .A1(n13088), .A2(n13090), .ZN(n15282) );
  OAI211_X1 U16265 ( .C1(n13090), .C2(n13088), .A(n13087), .B(n15282), .ZN(
        n13089) );
  AND2_X1 U16266 ( .A1(n10383), .A2(n13090), .ZN(n15290) );
  NAND2_X1 U16267 ( .A1(n15288), .A2(n15290), .ZN(n15289) );
  AOI22_X1 U16268 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9586), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13093) );
  AOI22_X1 U16269 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13092) );
  AND2_X1 U16270 ( .A1(n13093), .A2(n13092), .ZN(n13096) );
  AOI22_X1 U16271 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13095) );
  AOI22_X1 U16272 ( .A1(n13129), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13094) );
  NAND4_X1 U16273 ( .A1(n13096), .A2(n13095), .A3(n13094), .A4(n13134), .ZN(
        n13103) );
  AOI22_X1 U16274 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10235), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13098) );
  AOI22_X1 U16275 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13097) );
  AND2_X1 U16276 ( .A1(n13098), .A2(n13097), .ZN(n13101) );
  AOI22_X1 U16277 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13100) );
  AOI22_X1 U16278 ( .A1(n13129), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13099) );
  NAND4_X1 U16279 ( .A1(n13101), .A2(n13131), .A3(n13100), .A4(n13099), .ZN(
        n13102) );
  AOI21_X2 U16280 ( .B1(n15289), .B2(n9975), .A(n15283), .ZN(n15278) );
  AOI22_X1 U16281 ( .A1(n13129), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13133), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13110) );
  NAND2_X1 U16282 ( .A1(n9587), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n13107) );
  NAND2_X1 U16283 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n13106) );
  NAND2_X1 U16284 ( .A1(n10376), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n13105) );
  NAND2_X1 U16285 ( .A1(n10375), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n13104) );
  AND4_X1 U16286 ( .A1(n13107), .A2(n13106), .A3(n13105), .A4(n13104), .ZN(
        n13109) );
  AOI22_X1 U16287 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n9590), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13108) );
  NAND4_X1 U16288 ( .A1(n13110), .A2(n13109), .A3(n13108), .A4(n13134), .ZN(
        n13119) );
  NAND2_X1 U16289 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n13114) );
  NAND2_X1 U16290 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n13113) );
  NAND2_X1 U16291 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n13112) );
  NAND2_X1 U16292 ( .A1(n10375), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n13111) );
  AND4_X1 U16293 ( .A1(n13114), .A2(n13113), .A3(n13112), .A4(n13111), .ZN(
        n13117) );
  AOI22_X1 U16294 ( .A1(n13133), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13116) );
  AOI22_X1 U16295 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9586), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13115) );
  NAND4_X1 U16296 ( .A1(n13117), .A2(n13131), .A3(n13116), .A4(n13115), .ZN(
        n13118) );
  NAND2_X1 U16297 ( .A1(n13119), .A2(n13118), .ZN(n13124) );
  INV_X1 U16298 ( .A(n15283), .ZN(n13120) );
  NAND2_X1 U16299 ( .A1(n13297), .A2(n13120), .ZN(n13122) );
  OR2_X1 U16300 ( .A1(n15282), .A2(n13122), .ZN(n13123) );
  NOR2_X1 U16301 ( .A1(n13123), .A2(n13124), .ZN(n13125) );
  AOI21_X1 U16302 ( .B1(n13124), .B2(n13123), .A(n13125), .ZN(n15277) );
  INV_X1 U16303 ( .A(n13125), .ZN(n13126) );
  AOI22_X1 U16304 ( .A1(n13133), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13128) );
  AOI22_X1 U16305 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9587), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13127) );
  NAND2_X1 U16306 ( .A1(n13128), .A2(n13127), .ZN(n13143) );
  AOI22_X1 U16307 ( .A1(n13129), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9596), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13132) );
  AOI22_X1 U16308 ( .A1(n9590), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13130) );
  NAND3_X1 U16309 ( .A1(n13132), .A2(n13131), .A3(n13130), .ZN(n13142) );
  AOI22_X1 U16310 ( .A1(n13133), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9590), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13136) );
  AOI22_X1 U16311 ( .A1(n10374), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10375), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13135) );
  NAND3_X1 U16312 ( .A1(n13136), .A2(n13135), .A3(n13134), .ZN(n13141) );
  AOI22_X1 U16313 ( .A1(n13137), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10235), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13139) );
  AOI22_X1 U16314 ( .A1(n9596), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10376), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13138) );
  NAND2_X1 U16315 ( .A1(n13139), .A2(n13138), .ZN(n13140) );
  OAI22_X1 U16316 ( .A1(n13143), .A2(n13142), .B1(n13141), .B2(n13140), .ZN(
        n13144) );
  AND2_X1 U16317 ( .A1(n13145), .A2(n19721), .ZN(n16348) );
  AOI22_X1 U16318 ( .A1(n16340), .A2(n16334), .B1(n16350), .B2(n16348), .ZN(
        n13975) );
  NAND2_X1 U16319 ( .A1(n13975), .A2(n13146), .ZN(n13147) );
  NOR2_X1 U16320 ( .A1(n19167), .A2(n13298), .ZN(n13150) );
  NOR4_X1 U16321 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13154) );
  NOR4_X1 U16322 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n13153) );
  NOR4_X1 U16323 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13152) );
  NOR4_X1 U16324 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13151) );
  NAND4_X1 U16325 ( .A1(n13154), .A2(n13153), .A3(n13152), .A4(n13151), .ZN(
        n13159) );
  NOR4_X1 U16326 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n13157) );
  NOR4_X1 U16327 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13156) );
  NOR4_X1 U16328 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13155) );
  INV_X1 U16329 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19743) );
  NAND4_X1 U16330 ( .A1(n13157), .A2(n13156), .A3(n13155), .A4(n19743), .ZN(
        n13158) );
  INV_X1 U16331 ( .A(n13161), .ZN(n13162) );
  NAND2_X1 U16332 ( .A1(n14276), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13165) );
  INV_X1 U16333 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n13163) );
  OR2_X1 U16334 ( .A1(n14276), .A2(n13163), .ZN(n13164) );
  NAND2_X1 U16335 ( .A1(n13165), .A2(n13164), .ZN(n19106) );
  INV_X1 U16336 ( .A(n19106), .ZN(n13167) );
  INV_X1 U16337 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13166) );
  OAI22_X1 U16338 ( .A1(n15410), .A2(n13167), .B1(n19041), .B2(n13166), .ZN(
        n13173) );
  NAND2_X1 U16339 ( .A1(n19041), .A2(n19167), .ZN(n15385) );
  INV_X1 U16340 ( .A(n19010), .ZN(n15412) );
  INV_X1 U16341 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n14529) );
  OAI22_X1 U16342 ( .A1(n14548), .A2(n15385), .B1(n15412), .B2(n14529), .ZN(
        n13172) );
  AOI211_X1 U16343 ( .C1(n19011), .C2(BUF2_REG_30__SCAN_IN), .A(n13173), .B(
        n13172), .ZN(n13174) );
  NAND2_X1 U16344 ( .A1(n13175), .A2(n13174), .ZN(P2_U2889) );
  INV_X1 U16345 ( .A(n16340), .ZN(n16335) );
  NAND2_X1 U16346 ( .A1(n16335), .A2(n16339), .ZN(n13973) );
  NAND2_X1 U16347 ( .A1(n13973), .A2(n13177), .ZN(n13178) );
  NAND2_X1 U16348 ( .A1(n13179), .A2(n15342), .ZN(n13185) );
  NAND2_X1 U16349 ( .A1(n15419), .A2(n15316), .ZN(n13183) );
  INV_X1 U16350 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n13182) );
  NAND2_X1 U16351 ( .A1(n13185), .A2(n13184), .ZN(P2_U2857) );
  AOI21_X1 U16352 ( .B1(n15439), .B2(n13187), .A(n12849), .ZN(n15443) );
  AOI21_X1 U16353 ( .B1(n15484), .B2(n13188), .A(n13189), .ZN(n15487) );
  NOR2_X1 U16354 ( .A1(n13191), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13192) );
  NOR2_X1 U16355 ( .A1(n13190), .A2(n13192), .ZN(n15522) );
  AOI21_X1 U16356 ( .B1(n14244), .B2(n13193), .A(n13194), .ZN(n15566) );
  AOI21_X1 U16357 ( .B1(n16189), .B2(n13195), .A(n13196), .ZN(n16178) );
  NOR2_X1 U16358 ( .A1(n16206), .A2(n13197), .ZN(n13205) );
  AOI21_X1 U16359 ( .B1(n16206), .B2(n13197), .A(n13205), .ZN(n16199) );
  AOI21_X1 U16360 ( .B1(n16227), .B2(n13198), .A(n13199), .ZN(n18960) );
  AOI21_X1 U16361 ( .B1(n18973), .B2(n13200), .A(n13201), .ZN(n18971) );
  AOI21_X1 U16362 ( .B1(n16264), .B2(n13202), .A(n9623), .ZN(n16254) );
  AOI21_X1 U16363 ( .B1(n13984), .B2(n13203), .A(n13204), .ZN(n13982) );
  OAI22_X1 U16364 ( .A1(n13325), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n19003) );
  INV_X1 U16365 ( .A(n19003), .ZN(n13962) );
  AOI22_X1 U16366 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14051), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n13325), .ZN(n14048) );
  NOR2_X1 U16367 ( .A1(n13962), .A2(n14048), .ZN(n14011) );
  OAI21_X1 U16368 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n13203), .ZN(n14012) );
  NAND2_X1 U16369 ( .A1(n14011), .A2(n14012), .ZN(n13980) );
  NOR2_X1 U16370 ( .A1(n13982), .A2(n13980), .ZN(n13900) );
  OAI21_X1 U16371 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13204), .A(
        n13202), .ZN(n19124) );
  NAND2_X1 U16372 ( .A1(n13900), .A2(n19124), .ZN(n13993) );
  NOR2_X1 U16373 ( .A1(n16254), .A2(n13993), .ZN(n13889) );
  OAI21_X1 U16374 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n9623), .A(
        n13200), .ZN(n16253) );
  NAND2_X1 U16375 ( .A1(n13889), .A2(n16253), .ZN(n18969) );
  NOR2_X1 U16376 ( .A1(n18971), .A2(n18969), .ZN(n13863) );
  OAI21_X1 U16377 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13201), .A(
        n13198), .ZN(n16245) );
  NAND2_X1 U16378 ( .A1(n13863), .A2(n16245), .ZN(n18959) );
  NOR2_X1 U16379 ( .A1(n18960), .A2(n18959), .ZN(n13877) );
  OAI21_X1 U16380 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n13199), .A(
        n13197), .ZN(n16220) );
  NAND2_X1 U16381 ( .A1(n13877), .A2(n16220), .ZN(n13847) );
  NOR2_X1 U16382 ( .A1(n16199), .A2(n13847), .ZN(n13914) );
  OAI21_X1 U16383 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n13205), .A(
        n13195), .ZN(n16198) );
  NAND2_X1 U16384 ( .A1(n13914), .A2(n16198), .ZN(n14034) );
  NOR2_X1 U16385 ( .A1(n16178), .A2(n14034), .ZN(n18943) );
  OAI21_X1 U16386 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n13196), .A(
        n13193), .ZN(n18945) );
  NAND2_X1 U16387 ( .A1(n18943), .A2(n18945), .ZN(n14237) );
  NOR2_X1 U16388 ( .A1(n15566), .A2(n14237), .ZN(n18933) );
  OAI21_X1 U16389 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n13194), .A(
        n9696), .ZN(n18934) );
  AND2_X1 U16390 ( .A1(n18933), .A2(n18934), .ZN(n13206) );
  AOI21_X1 U16391 ( .B1(n9696), .B2(n15542), .A(n13208), .ZN(n18923) );
  NOR2_X1 U16392 ( .A1(n18922), .A2(n10114), .ZN(n18912) );
  NOR2_X1 U16393 ( .A1(n13208), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13209) );
  OR2_X1 U16394 ( .A1(n13191), .A2(n13209), .ZN(n18911) );
  OAI21_X1 U16395 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n13190), .A(
        n10777), .ZN(n15510) );
  INV_X1 U16396 ( .A(n15510), .ZN(n18903) );
  NOR2_X1 U16397 ( .A1(n9951), .A2(n18902), .ZN(n18886) );
  NOR2_X1 U16398 ( .A1(n18886), .A2(n18887), .ZN(n15888) );
  OAI21_X1 U16399 ( .B1(n9694), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n13188), .ZN(n15890) );
  AOI21_X1 U16400 ( .B1(n15888), .B2(n15890), .A(n9951), .ZN(n15254) );
  NOR2_X1 U16401 ( .A1(n15487), .A2(n15254), .ZN(n15255) );
  NOR2_X1 U16402 ( .A1(n9951), .A2(n15255), .ZN(n16151) );
  OR2_X1 U16403 ( .A1(n13189), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13211) );
  NAND2_X1 U16404 ( .A1(n13210), .A2(n13211), .ZN(n15473) );
  INV_X1 U16405 ( .A(n15473), .ZN(n16153) );
  NOR2_X1 U16406 ( .A1(n16151), .A2(n16153), .ZN(n16152) );
  NOR2_X1 U16407 ( .A1(n9951), .A2(n16152), .ZN(n15228) );
  AOI21_X1 U16408 ( .B1(n15467), .B2(n13210), .A(n13212), .ZN(n15465) );
  NOR2_X1 U16409 ( .A1(n15228), .A2(n15465), .ZN(n15229) );
  NOR2_X1 U16410 ( .A1(n9951), .A2(n15229), .ZN(n15217) );
  INV_X1 U16411 ( .A(n13187), .ZN(n13213) );
  AOI21_X1 U16412 ( .B1(n15449), .B2(n13214), .A(n13213), .ZN(n15452) );
  OR2_X1 U16413 ( .A1(n15217), .A2(n15452), .ZN(n15218) );
  INV_X1 U16414 ( .A(n13216), .ZN(n13217) );
  NOR2_X1 U16415 ( .A1(n15177), .A2(n15435), .ZN(n15165) );
  NOR2_X1 U16416 ( .A1(n9951), .A2(n15165), .ZN(n13218) );
  XNOR2_X1 U16417 ( .A(n13216), .B(n13234), .ZN(n15423) );
  XNOR2_X1 U16418 ( .A(n13218), .B(n15423), .ZN(n13219) );
  NAND4_X1 U16419 ( .A1(n13325), .A2(n19848), .A3(n19791), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19717) );
  NAND2_X1 U16420 ( .A1(n13219), .A2(n18984), .ZN(n13243) );
  NAND2_X1 U16421 ( .A1(n19791), .A2(n16347), .ZN(n16360) );
  NOR2_X1 U16422 ( .A1(n14548), .A2(n18989), .ZN(n13241) );
  OR2_X1 U16423 ( .A1(n19841), .A2(n13221), .ZN(n13224) );
  NAND2_X1 U16424 ( .A1(n19791), .A2(n19721), .ZN(n13222) );
  NAND2_X1 U16425 ( .A1(n15419), .A2(n18999), .ZN(n13239) );
  INV_X1 U16426 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n13223) );
  INV_X1 U16427 ( .A(n13222), .ZN(n13229) );
  INV_X2 U16428 ( .A(n19113), .ZN(n15534) );
  AND3_X1 U16429 ( .A1(n19848), .A2(n19714), .A3(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n16365) );
  NOR2_X1 U16430 ( .A1(n18984), .A2(n16365), .ZN(n13225) );
  AND2_X1 U16431 ( .A1(n15534), .A2(n13225), .ZN(n13226) );
  NAND2_X1 U16432 ( .A1(n19109), .A2(n16360), .ZN(n13232) );
  INV_X1 U16433 ( .A(n13275), .ZN(n13268) );
  NOR2_X1 U16434 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13229), .ZN(n13230) );
  NAND2_X1 U16435 ( .A1(n13268), .A2(n13230), .ZN(n13231) );
  NAND2_X2 U16436 ( .A1(n13232), .A2(n13231), .ZN(n18992) );
  AOI22_X1 U16437 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n18992), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n18951), .ZN(n13233) );
  OAI21_X1 U16438 ( .B1(n13234), .B2(n18974), .A(n13233), .ZN(n13235) );
  AOI21_X1 U16439 ( .B1(n13237), .B2(n13236), .A(n13235), .ZN(n13238) );
  NAND2_X1 U16440 ( .A1(n13243), .A2(n13242), .ZN(P2_U2825) );
  NOR2_X1 U16441 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13245) );
  NOR4_X1 U16442 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13244) );
  NAND4_X1 U16443 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13245), .A4(n13244), .ZN(n13248) );
  INV_X1 U16444 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20737) );
  NOR3_X1 U16445 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20737), .ZN(n13247) );
  NOR4_X1 U16446 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13246) );
  NAND4_X1 U16447 ( .A1(n20053), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13247), .A4(
        n13246), .ZN(U214) );
  NOR2_X1 U16448 ( .A1(n14276), .A2(n13248), .ZN(n16443) );
  NAND2_X1 U16449 ( .A1(n16443), .A2(U214), .ZN(U212) );
  INV_X1 U16450 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17552) );
  OR2_X1 U16451 ( .A1(n16912), .A2(n17575), .ZN(n17549) );
  NOR2_X1 U16452 ( .A1(n17574), .A2(n17549), .ZN(n13250) );
  NAND2_X1 U16453 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n13250), .ZN(
        n13249) );
  NOR2_X1 U16454 ( .A1(n16912), .A2(n17543), .ZN(n17513) );
  AOI21_X1 U16455 ( .B1(n17552), .B2(n13249), .A(n17513), .ZN(n17555) );
  XOR2_X1 U16456 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n13250), .Z(
        n17566) );
  AOI21_X1 U16457 ( .B1(n17574), .B2(n17549), .A(n13250), .ZN(n17576) );
  INV_X1 U16458 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17602) );
  INV_X1 U16459 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17590) );
  NOR2_X1 U16460 ( .A1(n17602), .A2(n17590), .ZN(n17586) );
  INV_X1 U16461 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16578) );
  NAND2_X1 U16462 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16398), .ZN(
        n13251) );
  XOR2_X2 U16463 ( .A(n16578), .B(n13251), .Z(n16876) );
  NAND2_X1 U16464 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17635) );
  NAND2_X1 U16465 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17634), .ZN(
        n17629) );
  NOR2_X1 U16466 ( .A1(n17635), .A2(n17629), .ZN(n16712) );
  NAND2_X1 U16467 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16712), .ZN(
        n17588) );
  OAI21_X1 U16468 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17588), .A(
        n16876), .ZN(n16693) );
  OAI21_X1 U16469 ( .B1(n17586), .B2(n9919), .A(n16693), .ZN(n16673) );
  NOR2_X1 U16470 ( .A1(n17555), .A2(n13252), .ZN(n16567) );
  NAND4_X1 U16471 ( .A1(n18688), .A2(n15851), .A3(n18841), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n18694) );
  AOI211_X1 U16472 ( .C1(n17555), .C2(n13252), .A(n16567), .B(n18694), .ZN(
        n13266) );
  NOR3_X1 U16473 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16893) );
  INV_X1 U16474 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17183) );
  NAND2_X1 U16475 ( .A1(n16893), .A2(n17183), .ZN(n16880) );
  NOR2_X1 U16476 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16880), .ZN(n16859) );
  INV_X1 U16477 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16854) );
  NAND2_X1 U16478 ( .A1(n16859), .A2(n16854), .ZN(n16853) );
  INV_X1 U16479 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17167) );
  NAND2_X1 U16480 ( .A1(n16834), .A2(n17167), .ZN(n16823) );
  NAND2_X1 U16481 ( .A1(n16805), .A2(n17123), .ZN(n16801) );
  INV_X1 U16482 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17094) );
  NAND2_X1 U16483 ( .A1(n16789), .A2(n17094), .ZN(n16779) );
  INV_X1 U16484 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16761) );
  NAND2_X1 U16485 ( .A1(n16762), .A2(n16761), .ZN(n16758) );
  INV_X1 U16486 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17064) );
  NAND2_X1 U16487 ( .A1(n16739), .A2(n17064), .ZN(n16734) );
  INV_X1 U16488 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16704) );
  NAND2_X1 U16489 ( .A1(n16716), .A2(n16704), .ZN(n16702) );
  INV_X1 U16490 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16686) );
  NAND2_X1 U16491 ( .A1(n16694), .A2(n16686), .ZN(n16684) );
  INV_X1 U16492 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16667) );
  NAND2_X1 U16493 ( .A1(n16674), .A2(n16667), .ZN(n16665) );
  NAND2_X1 U16494 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18843) );
  NOR2_X4 U16495 ( .A1(n13254), .A2(n13253), .ZN(n15853) );
  NAND2_X1 U16496 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18193), .ZN(n13258) );
  AOI211_X4 U16497 ( .C1(n18841), .C2(n18843), .A(n13260), .B(n13258), .ZN(
        n16881) );
  AOI211_X1 U16498 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16665), .A(n16660), .B(
        n16916), .ZN(n13265) );
  NAND2_X1 U16499 ( .A1(n18688), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18562) );
  OR2_X1 U16500 ( .A1(n18690), .A2(n18562), .ZN(n18685) );
  INV_X1 U16501 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n16925) );
  NOR2_X1 U16502 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18703) );
  NOR3_X1 U16503 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18725), .A3(n18703), 
        .ZN(n15863) );
  OAI211_X1 U16504 ( .C1(n18193), .C2(n15863), .A(n18843), .B(n18841), .ZN(
        n18680) );
  OAI211_X2 U16505 ( .C1(n16925), .C2(n18842), .A(n18680), .B(n13259), .ZN(
        n16917) );
  INV_X1 U16506 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16949) );
  OAI22_X1 U16507 ( .A1(n17552), .A2(n16907), .B1(n16917), .B2(n16949), .ZN(
        n13264) );
  INV_X1 U16508 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18759) );
  INV_X1 U16509 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18756) );
  INV_X1 U16510 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18754) );
  NOR3_X1 U16511 ( .A1(n18759), .A2(n18756), .A3(n18754), .ZN(n13261) );
  NAND3_X1 U16512 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16556) );
  INV_X1 U16513 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18742) );
  INV_X1 U16514 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18738) );
  INV_X1 U16515 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18734) );
  INV_X1 U16516 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18726) );
  NAND3_X1 U16517 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16863) );
  NOR2_X1 U16518 ( .A1(n18726), .A2(n16863), .ZN(n16847) );
  NAND2_X1 U16519 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16847), .ZN(n16825) );
  NAND2_X1 U16520 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n16809) );
  NOR3_X1 U16521 ( .A1(n18734), .A2(n16825), .A3(n16809), .ZN(n16808) );
  NAND2_X1 U16522 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16808), .ZN(n16788) );
  NOR2_X1 U16523 ( .A1(n18738), .A2(n16788), .ZN(n16771) );
  NAND2_X1 U16524 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16771), .ZN(n16770) );
  NOR2_X1 U16525 ( .A1(n18742), .A2(n16770), .ZN(n16740) );
  NAND4_X1 U16526 ( .A1(n16869), .A2(P3_REIP_REG_14__SCAN_IN), .A3(
        P3_REIP_REG_13__SCAN_IN), .A4(n16740), .ZN(n16726) );
  NOR2_X1 U16527 ( .A1(n16556), .A2(n16726), .ZN(n16691) );
  NAND2_X1 U16528 ( .A1(n13261), .A2(n16691), .ZN(n16671) );
  XNOR2_X1 U16529 ( .A(P3_REIP_REG_22__SCAN_IN), .B(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n13262) );
  INV_X1 U16530 ( .A(n13261), .ZN(n16555) );
  NAND3_X1 U16531 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n16740), .ZN(n16720) );
  OR3_X1 U16532 ( .A1(n16919), .A2(n16720), .A3(n16556), .ZN(n16701) );
  NOR2_X1 U16533 ( .A1(n16919), .A2(n16869), .ZN(n16722) );
  INV_X1 U16534 ( .A(n16722), .ZN(n16922) );
  OAI21_X1 U16535 ( .B1(n16555), .B2(n16701), .A(n16922), .ZN(n16679) );
  INV_X1 U16536 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18762) );
  OAI22_X1 U16537 ( .A1(n16671), .A2(n13262), .B1(n16679), .B2(n18762), .ZN(
        n13263) );
  OR4_X1 U16538 ( .A1(n13266), .A2(n13265), .A3(n13264), .A4(n13263), .ZN(
        P3_U2649) );
  OR2_X1 U16539 ( .A1(n10966), .A2(n18863), .ZN(n13321) );
  OR2_X1 U16540 ( .A1(n16337), .A2(n13321), .ZN(n18985) );
  INV_X1 U16541 ( .A(n18985), .ZN(n13270) );
  INV_X1 U16542 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13269) );
  NOR2_X1 U16543 ( .A1(n13268), .A2(n13267), .ZN(n13272) );
  OAI21_X1 U16544 ( .B1(n13270), .B2(n13269), .A(n13272), .ZN(P2_U2814) );
  INV_X1 U16545 ( .A(n19841), .ZN(n13273) );
  NOR2_X1 U16546 ( .A1(n13270), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n13271)
         );
  AOI22_X1 U16547 ( .A1(n13274), .A2(n13273), .B1(n13272), .B2(n13271), .ZN(
        P2_U3612) );
  INV_X1 U16548 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13279) );
  NOR2_X1 U16549 ( .A1(n13275), .A2(n19849), .ZN(n13276) );
  OR2_X1 U16550 ( .A1(n19109), .A2(n13276), .ZN(n13311) );
  INV_X1 U16551 ( .A(n19107), .ZN(n13278) );
  AOI22_X1 U16552 ( .A1(n14278), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14276), .ZN(n19017) );
  INV_X1 U16553 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13277) );
  OAI222_X1 U16554 ( .A1(n13279), .A2(n13311), .B1(n13278), .B2(n19017), .C1(
        n13532), .C2(n13277), .ZN(P2_U2982) );
  NOR2_X1 U16555 ( .A1(n11789), .A2(n13285), .ZN(n13284) );
  NAND2_X1 U16556 ( .A1(n13284), .A2(n13280), .ZN(n14562) );
  NOR2_X1 U16557 ( .A1(n11470), .A2(n13281), .ZN(n13283) );
  NOR2_X1 U16558 ( .A1(n20573), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14228) );
  OAI21_X1 U16559 ( .B1(n14228), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n20738), 
        .ZN(n13282) );
  OAI21_X1 U16560 ( .B1(n20738), .B2(n13283), .A(n13282), .ZN(P1_U3487) );
  OAI22_X1 U16561 ( .A1(n15927), .A2(n13284), .B1(n11470), .B2(n13444), .ZN(
        n19863) );
  AOI21_X1 U16562 ( .B1(n13477), .B2(n15956), .A(n20741), .ZN(n20746) );
  NOR2_X1 U16563 ( .A1(n19863), .A2(n20746), .ZN(n15916) );
  NOR2_X1 U16564 ( .A1(n15916), .A2(n19862), .ZN(n19871) );
  INV_X1 U16565 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13296) );
  INV_X1 U16566 ( .A(n13285), .ZN(n13294) );
  INV_X1 U16567 ( .A(n15920), .ZN(n13287) );
  NAND2_X1 U16568 ( .A1(n13287), .A2(n13286), .ZN(n13288) );
  OR2_X1 U16569 ( .A1(n13288), .A2(n15927), .ZN(n13289) );
  NAND2_X1 U16570 ( .A1(n13289), .A2(n15936), .ZN(n13293) );
  INV_X1 U16571 ( .A(n13290), .ZN(n13291) );
  NAND2_X1 U16572 ( .A1(n13444), .A2(n13291), .ZN(n13292) );
  OAI211_X1 U16573 ( .C1(n13294), .C2(n11789), .A(n13293), .B(n13292), .ZN(
        n15918) );
  NAND2_X1 U16574 ( .A1(n19871), .A2(n15918), .ZN(n13295) );
  OAI21_X1 U16575 ( .B1(n19871), .B2(n13296), .A(n13295), .ZN(P1_U3484) );
  INV_X1 U16576 ( .A(n13968), .ZN(n13301) );
  NAND2_X1 U16577 ( .A1(n13297), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13299) );
  NAND4_X1 U16578 ( .A1(n13299), .A2(n13298), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19839), .ZN(n13300) );
  MUX2_X1 U16579 ( .A(n10554), .B(n13963), .S(n15316), .Z(n13302) );
  OAI21_X1 U16580 ( .B1(n18986), .B2(n15350), .A(n13302), .ZN(P2_U2887) );
  XOR2_X1 U16581 ( .A(n18994), .B(n13304), .Z(n13414) );
  NOR2_X1 U16582 ( .A1(n15534), .A2(n18988), .ZN(n13412) );
  AOI21_X1 U16583 ( .B1(n13305), .B2(n13304), .A(n13303), .ZN(n13306) );
  INV_X1 U16584 ( .A(n13306), .ZN(n13410) );
  NOR2_X1 U16585 ( .A1(n16256), .A2(n13410), .ZN(n13307) );
  AOI211_X1 U16586 ( .C1(n19121), .C2(n13414), .A(n13412), .B(n13307), .ZN(
        n13310) );
  OAI21_X1 U16587 ( .B1(n19114), .B2(n13308), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13309) );
  OAI211_X1 U16588 ( .C1(n16247), .C2(n13963), .A(n13310), .B(n13309), .ZN(
        P2_U3014) );
  INV_X1 U16589 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13332) );
  INV_X2 U16590 ( .A(n13311), .ZN(n19110) );
  NAND2_X1 U16591 ( .A1(n19110), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13314) );
  NAND2_X1 U16592 ( .A1(n14276), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13313) );
  INV_X1 U16593 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16474) );
  OR2_X1 U16594 ( .A1(n14276), .A2(n16474), .ZN(n13312) );
  NAND2_X1 U16595 ( .A1(n13313), .A2(n13312), .ZN(n19023) );
  NAND2_X1 U16596 ( .A1(n19107), .A2(n19023), .ZN(n13526) );
  OAI211_X1 U16597 ( .C1(n13332), .C2(n13532), .A(n13314), .B(n13526), .ZN(
        P2_U2964) );
  NAND2_X1 U16598 ( .A1(n19110), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13317) );
  NAND2_X1 U16599 ( .A1(n14276), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13316) );
  INV_X1 U16600 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16478) );
  OR2_X1 U16601 ( .A1(n14276), .A2(n16478), .ZN(n13315) );
  NAND2_X1 U16602 ( .A1(n13316), .A2(n13315), .ZN(n19028) );
  NAND2_X1 U16603 ( .A1(n19107), .A2(n19028), .ZN(n13530) );
  OAI211_X1 U16604 ( .C1(n15370), .C2(n13532), .A(n13317), .B(n13530), .ZN(
        P2_U2962) );
  INV_X1 U16605 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13334) );
  NAND2_X1 U16606 ( .A1(n19110), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13320) );
  NAND2_X1 U16607 ( .A1(n14276), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13319) );
  INV_X1 U16608 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16481) );
  OR2_X1 U16609 ( .A1(n14276), .A2(n16481), .ZN(n13318) );
  NAND2_X1 U16610 ( .A1(n13319), .A2(n13318), .ZN(n19034) );
  NAND2_X1 U16611 ( .A1(n19107), .A2(n19034), .ZN(n13528) );
  OAI211_X1 U16612 ( .C1(n13334), .C2(n13532), .A(n13320), .B(n13528), .ZN(
        P2_U2960) );
  INV_X1 U16613 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n15409) );
  OAI21_X1 U16614 ( .B1(n13322), .B2(n13321), .A(n13532), .ZN(n13323) );
  NAND2_X1 U16615 ( .A1(n14270), .A2(n13325), .ZN(n19843) );
  INV_X2 U16616 ( .A(n19843), .ZN(n19099) );
  AOI22_X1 U16617 ( .A1(n19099), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13326) );
  OAI21_X1 U16618 ( .B1(n15409), .B2(n19067), .A(n13326), .ZN(P2_U2932) );
  AOI22_X1 U16619 ( .A1(n19099), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13327) );
  OAI21_X1 U16620 ( .B1(n20882), .B2(n19067), .A(n13327), .ZN(P2_U2924) );
  AOI22_X1 U16621 ( .A1(n19099), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13328) );
  OAI21_X1 U16622 ( .B1(n15376), .B2(n19067), .A(n13328), .ZN(P2_U2926) );
  AOI22_X1 U16623 ( .A1(n19099), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13329) );
  OAI21_X1 U16624 ( .B1(n15370), .B2(n19067), .A(n13329), .ZN(P2_U2925) );
  AOI22_X1 U16625 ( .A1(n19099), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13330) );
  OAI21_X1 U16626 ( .B1(n11238), .B2(n19067), .A(n13330), .ZN(P2_U2929) );
  AOI22_X1 U16627 ( .A1(n19099), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13331) );
  OAI21_X1 U16628 ( .B1(n13332), .B2(n19067), .A(n13331), .ZN(P2_U2923) );
  AOI22_X1 U16629 ( .A1(n19099), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13333) );
  OAI21_X1 U16630 ( .B1(n13334), .B2(n19067), .A(n13333), .ZN(P2_U2927) );
  INV_X1 U16631 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15389) );
  AOI22_X1 U16632 ( .A1(n19099), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13335) );
  OAI21_X1 U16633 ( .B1(n15389), .B2(n19067), .A(n13335), .ZN(P2_U2928) );
  AOI22_X1 U16634 ( .A1(n19099), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13336) );
  OAI21_X1 U16635 ( .B1(n11232), .B2(n19067), .A(n13336), .ZN(P2_U2933) );
  AOI22_X1 U16636 ( .A1(n19099), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13337) );
  OAI21_X1 U16637 ( .B1(n15352), .B2(n19067), .A(n13337), .ZN(P2_U2922) );
  INV_X1 U16638 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13339) );
  AOI22_X1 U16639 ( .A1(n19099), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13338) );
  OAI21_X1 U16640 ( .B1(n13339), .B2(n19067), .A(n13338), .ZN(P2_U2935) );
  INV_X1 U16641 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13341) );
  AOI22_X1 U16642 ( .A1(n19099), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13340) );
  OAI21_X1 U16643 ( .B1(n13341), .B2(n19067), .A(n13340), .ZN(P2_U2931) );
  AOI22_X1 U16644 ( .A1(n19099), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13342) );
  OAI21_X1 U16645 ( .B1(n14254), .B2(n19067), .A(n13342), .ZN(P2_U2934) );
  AOI22_X1 U16646 ( .A1(n19099), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13343) );
  OAI21_X1 U16647 ( .B1(n15403), .B2(n19067), .A(n13343), .ZN(P2_U2930) );
  AOI21_X1 U16648 ( .B1(n13345), .B2(n14181), .A(n13344), .ZN(n13346) );
  XOR2_X1 U16649 ( .A(n13346), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n15795) );
  NOR2_X1 U16650 ( .A1(n15534), .A2(n10272), .ZN(n15794) );
  OAI21_X1 U16651 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13348), .A(
        n13347), .ZN(n15791) );
  NOR2_X1 U16652 ( .A1(n16256), .A2(n15791), .ZN(n13349) );
  AOI211_X1 U16653 ( .C1(n19121), .C2(n15795), .A(n15794), .B(n13349), .ZN(
        n13351) );
  MUX2_X1 U16654 ( .A(n19125), .B(n16265), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n13350) );
  OAI211_X1 U16655 ( .C1(n15792), .C2(n16247), .A(n13351), .B(n13350), .ZN(
        P2_U3013) );
  AOI22_X1 U16656 ( .A1(n19110), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(
        P2_EAX_REG_16__SCAN_IN), .B2(n19109), .ZN(n13352) );
  OAI22_X1 U16657 ( .A1(n14276), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n14278), .ZN(n14283) );
  INV_X1 U16658 ( .A(n14283), .ZN(n19008) );
  NAND2_X1 U16659 ( .A1(n19107), .A2(n19008), .ZN(n13501) );
  NAND2_X1 U16660 ( .A1(n13352), .A2(n13501), .ZN(P2_U2952) );
  AOI22_X1 U16661 ( .A1(n19110), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n19109), .ZN(n13353) );
  OAI22_X1 U16662 ( .A1(n14276), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14278), .ZN(n19150) );
  INV_X1 U16663 ( .A(n19150), .ZN(n16168) );
  NAND2_X1 U16664 ( .A1(n19107), .A2(n16168), .ZN(n13503) );
  NAND2_X1 U16665 ( .A1(n13353), .A2(n13503), .ZN(P2_U2954) );
  AOI22_X1 U16666 ( .A1(n19110), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19109), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n13357) );
  INV_X1 U16667 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14795) );
  OR2_X1 U16668 ( .A1(n14276), .A2(n14795), .ZN(n13355) );
  NAND2_X1 U16669 ( .A1(n14276), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13354) );
  AND2_X1 U16670 ( .A1(n13355), .A2(n13354), .ZN(n19021) );
  INV_X1 U16671 ( .A(n19021), .ZN(n13356) );
  NAND2_X1 U16672 ( .A1(n19107), .A2(n13356), .ZN(n13511) );
  NAND2_X1 U16673 ( .A1(n13357), .A2(n13511), .ZN(P2_U2980) );
  AOI22_X1 U16674 ( .A1(n19110), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n19109), .ZN(n13362) );
  INV_X1 U16675 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13358) );
  OR2_X1 U16676 ( .A1(n14276), .A2(n13358), .ZN(n13360) );
  NAND2_X1 U16677 ( .A1(n14276), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13359) );
  AND2_X1 U16678 ( .A1(n13360), .A2(n13359), .ZN(n19026) );
  INV_X1 U16679 ( .A(n19026), .ZN(n13361) );
  NAND2_X1 U16680 ( .A1(n19107), .A2(n13361), .ZN(n13509) );
  NAND2_X1 U16681 ( .A1(n13362), .A2(n13509), .ZN(P2_U2963) );
  AOI22_X1 U16682 ( .A1(n19110), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19109), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13364) );
  AOI22_X1 U16683 ( .A1(n14278), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14276), .ZN(n19155) );
  INV_X1 U16684 ( .A(n19155), .ZN(n13363) );
  NAND2_X1 U16685 ( .A1(n19107), .A2(n13363), .ZN(n13515) );
  NAND2_X1 U16686 ( .A1(n13364), .A2(n13515), .ZN(P2_U2955) );
  AOI22_X1 U16687 ( .A1(n19110), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n19109), .ZN(n13368) );
  INV_X1 U16688 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n14330) );
  OR2_X1 U16689 ( .A1(n14276), .A2(n14330), .ZN(n13366) );
  NAND2_X1 U16690 ( .A1(n14276), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13365) );
  AND2_X1 U16691 ( .A1(n13366), .A2(n13365), .ZN(n19031) );
  INV_X1 U16692 ( .A(n19031), .ZN(n13367) );
  NAND2_X1 U16693 ( .A1(n19107), .A2(n13367), .ZN(n13499) );
  NAND2_X1 U16694 ( .A1(n13368), .A2(n13499), .ZN(P2_U2961) );
  AOI22_X1 U16695 ( .A1(n19110), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19109), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13370) );
  AOI22_X1 U16696 ( .A1(n14278), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14276), .ZN(n19169) );
  INV_X1 U16697 ( .A(n19169), .ZN(n13369) );
  NAND2_X1 U16698 ( .A1(n19107), .A2(n13369), .ZN(n13495) );
  NAND2_X1 U16699 ( .A1(n13370), .A2(n13495), .ZN(P2_U2959) );
  AOI22_X1 U16700 ( .A1(n19110), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n19109), .ZN(n13372) );
  AOI22_X1 U16701 ( .A1(n14278), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n14276), .ZN(n19038) );
  INV_X1 U16702 ( .A(n19038), .ZN(n13371) );
  NAND2_X1 U16703 ( .A1(n19107), .A2(n13371), .ZN(n13497) );
  NAND2_X1 U16704 ( .A1(n13372), .A2(n13497), .ZN(P2_U2958) );
  AOI22_X1 U16705 ( .A1(n19110), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19109), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13374) );
  AOI22_X1 U16706 ( .A1(n14278), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n14276), .ZN(n19065) );
  INV_X1 U16707 ( .A(n19065), .ZN(n13373) );
  NAND2_X1 U16708 ( .A1(n19107), .A2(n13373), .ZN(n13505) );
  NAND2_X1 U16709 ( .A1(n13374), .A2(n13505), .ZN(P2_U2953) );
  AOI22_X1 U16710 ( .A1(n19110), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19109), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13376) );
  AOI22_X1 U16711 ( .A1(n14278), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14276), .ZN(n19040) );
  INV_X1 U16712 ( .A(n19040), .ZN(n13375) );
  NAND2_X1 U16713 ( .A1(n19107), .A2(n13375), .ZN(n13507) );
  NAND2_X1 U16714 ( .A1(n13376), .A2(n13507), .ZN(P2_U2957) );
  AOI22_X1 U16715 ( .A1(n19110), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n19109), .ZN(n13377) );
  OAI22_X1 U16716 ( .A1(n14276), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n14278), .ZN(n19159) );
  INV_X1 U16717 ( .A(n19159), .ZN(n16163) );
  NAND2_X1 U16718 ( .A1(n19107), .A2(n16163), .ZN(n13513) );
  NAND2_X1 U16719 ( .A1(n13377), .A2(n13513), .ZN(P2_U2956) );
  AOI21_X1 U16720 ( .B1(n9607), .B2(n13379), .A(n11064), .ZN(n13413) );
  INV_X1 U16721 ( .A(n13413), .ZN(n18990) );
  NOR2_X1 U16722 ( .A1(n18986), .A2(n18990), .ZN(n19059) );
  INV_X1 U16723 ( .A(n19059), .ZN(n13380) );
  OAI211_X1 U16724 ( .C1(n19825), .C2(n13413), .A(n13380), .B(n13149), .ZN(
        n13382) );
  AOI22_X1 U16725 ( .A1(n19056), .A2(n13413), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19055), .ZN(n13381) );
  OAI211_X1 U16726 ( .C1(n19064), .C2(n14283), .A(n13382), .B(n13381), .ZN(
        P2_U2919) );
  NOR2_X1 U16727 ( .A1(n15792), .A2(n13618), .ZN(n13386) );
  AOI21_X1 U16728 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n13618), .A(n13386), .ZN(
        n13387) );
  OAI21_X1 U16729 ( .B1(n19816), .B2(n15350), .A(n13387), .ZN(P2_U2886) );
  AND2_X1 U16730 ( .A1(n11496), .A2(n20741), .ZN(n13388) );
  OR2_X1 U16731 ( .A1(n20026), .A2(n20076), .ZN(n13587) );
  INV_X1 U16732 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13392) );
  OR2_X1 U16733 ( .A1(n20026), .A2(n15926), .ZN(n13588) );
  INV_X1 U16734 ( .A(n20053), .ZN(n20054) );
  INV_X1 U16735 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13389) );
  NOR2_X1 U16736 ( .A1(n20054), .A2(n13389), .ZN(n13390) );
  AOI21_X1 U16737 ( .B1(DATAI_15_), .B2(n20054), .A(n13390), .ZN(n14860) );
  INV_X1 U16738 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13391) );
  OAI222_X1 U16739 ( .A1(n13587), .A2(n13392), .B1(n13588), .B2(n14860), .C1(
        n13391), .C2(n13596), .ZN(P1_U2967) );
  XNOR2_X1 U16740 ( .A(n13394), .B(n13393), .ZN(n19134) );
  INV_X1 U16741 ( .A(n14012), .ZN(n13401) );
  XNOR2_X1 U16742 ( .A(n13396), .B(n13395), .ZN(n19136) );
  NAND2_X1 U16743 ( .A1(n19114), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13398) );
  OR2_X1 U16744 ( .A1(n15534), .A2(n13397), .ZN(n19145) );
  OAI211_X1 U16745 ( .C1(n16256), .C2(n19136), .A(n13398), .B(n19145), .ZN(
        n13400) );
  NOR2_X1 U16746 ( .A1(n19139), .A2(n16247), .ZN(n13399) );
  AOI211_X1 U16747 ( .C1(n16255), .C2(n13401), .A(n13400), .B(n13399), .ZN(
        n13402) );
  OAI21_X1 U16748 ( .B1(n16258), .B2(n19134), .A(n13402), .ZN(P2_U3012) );
  INV_X1 U16749 ( .A(n13403), .ZN(n13406) );
  OR2_X1 U16750 ( .A1(n13404), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13405) );
  AND2_X1 U16751 ( .A1(n13406), .A2(n13405), .ZN(n14107) );
  INV_X1 U16752 ( .A(n14107), .ZN(n13409) );
  XNOR2_X1 U16753 ( .A(n13408), .B(n13407), .ZN(n14114) );
  OAI222_X1 U16754 ( .A1(n19985), .A2(n13409), .B1(n11872), .B2(n19997), .C1(
        n19992), .C2(n14114), .ZN(P1_U2872) );
  OAI22_X1 U16755 ( .A1(n13963), .A2(n19138), .B1(n19137), .B2(n13410), .ZN(
        n13411) );
  AOI211_X1 U16756 ( .C1(n19130), .C2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13412), .B(n13411), .ZN(n13416) );
  AOI22_X1 U16757 ( .A1(n16300), .A2(n13414), .B1(n16298), .B2(n13413), .ZN(
        n13415) );
  OAI211_X1 U16758 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n15766), .A(
        n13416), .B(n13415), .ZN(P2_U3046) );
  INV_X1 U16759 ( .A(n13463), .ZN(n13417) );
  OAI22_X1 U16760 ( .A1(n14564), .A2(n20076), .B1(n13417), .B2(n13643), .ZN(
        n13419) );
  NAND2_X1 U16761 ( .A1(n19998), .A2(n20061), .ZN(n13633) );
  NAND2_X1 U16762 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16145) );
  NAND2_X1 U16763 ( .A1(n20744), .A2(n13672), .ZN(n20740) );
  NOR2_X4 U16764 ( .A1(n19998), .A2(n20017), .ZN(n20016) );
  AOI22_X1 U16765 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13420) );
  OAI21_X1 U16766 ( .B1(n14802), .B2(n13633), .A(n13420), .ZN(P1_U2908) );
  AOI22_X1 U16767 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13421) );
  OAI21_X1 U16768 ( .B1(n14810), .B2(n13633), .A(n13421), .ZN(P1_U2910) );
  AOI22_X1 U16769 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13422) );
  OAI21_X1 U16770 ( .B1(n14797), .B2(n13633), .A(n13422), .ZN(P1_U2907) );
  INV_X1 U16771 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13424) );
  AOI22_X1 U16772 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13423) );
  OAI21_X1 U16773 ( .B1(n13424), .B2(n13633), .A(n13423), .ZN(P1_U2912) );
  AOI22_X1 U16774 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13425) );
  OAI21_X1 U16775 ( .B1(n12411), .B2(n13633), .A(n13425), .ZN(P1_U2909) );
  INV_X1 U16776 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13427) );
  AOI22_X1 U16777 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13426) );
  OAI21_X1 U16778 ( .B1(n13427), .B2(n13633), .A(n13426), .ZN(P1_U2906) );
  AOI22_X1 U16779 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13428) );
  OAI21_X1 U16780 ( .B1(n14814), .B2(n13633), .A(n13428), .ZN(P1_U2911) );
  NAND3_X1 U16781 ( .A1(n11855), .A2(n13431), .A3(n13430), .ZN(n13432) );
  NOR2_X1 U16782 ( .A1(n13433), .A2(n13432), .ZN(n13434) );
  NAND2_X1 U16783 ( .A1(n13434), .A2(n12512), .ZN(n14555) );
  INV_X1 U16784 ( .A(n14555), .ZN(n13484) );
  OR2_X1 U16785 ( .A1(n20537), .A2(n13484), .ZN(n13441) );
  INV_X1 U16786 ( .A(n13435), .ZN(n13443) );
  INV_X1 U16787 ( .A(n13663), .ZN(n13437) );
  NAND3_X1 U16788 ( .A1(n13478), .A2(n13443), .A3(n13437), .ZN(n13438) );
  OAI21_X1 U16789 ( .B1(n13643), .B2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13438), .ZN(n13439) );
  INV_X1 U16790 ( .A(n13439), .ZN(n13440) );
  NAND2_X1 U16791 ( .A1(n13441), .A2(n13440), .ZN(n15902) );
  INV_X1 U16792 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13442) );
  OAI22_X1 U16793 ( .A1(n9866), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n13442), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13489) );
  NAND2_X1 U16794 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13490) );
  NOR2_X1 U16795 ( .A1(n13489), .A2(n13490), .ZN(n13446) );
  INV_X1 U16796 ( .A(n13443), .ZN(n13639) );
  NOR3_X1 U16797 ( .A1(n13663), .A2(n13639), .A3(n20705), .ZN(n13445) );
  AOI211_X1 U16798 ( .C1(n15902), .C2(n14558), .A(n13446), .B(n13445), .ZN(
        n13459) );
  INV_X1 U16799 ( .A(n13447), .ZN(n13457) );
  NAND2_X1 U16800 ( .A1(n13643), .A2(n11855), .ZN(n13451) );
  INV_X1 U16801 ( .A(n13448), .ZN(n13450) );
  NAND2_X1 U16802 ( .A1(n12514), .A2(n15956), .ZN(n13449) );
  NAND3_X1 U16803 ( .A1(n13451), .A2(n13450), .A3(n13449), .ZN(n13455) );
  OR2_X1 U16804 ( .A1(n14091), .A2(n11477), .ZN(n13452) );
  AND4_X1 U16805 ( .A1(n13455), .A2(n13454), .A3(n13453), .A4(n13452), .ZN(
        n13456) );
  INV_X1 U16806 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19870) );
  NAND2_X1 U16807 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13672), .ZN(n16150) );
  OAI22_X1 U16808 ( .A1(n13665), .A2(n19862), .B1(n19870), .B2(n16150), .ZN(
        n13472) );
  AOI21_X1 U16809 ( .B1(n20744), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n13472), 
        .ZN(n14560) );
  NAND2_X1 U16810 ( .A1(n13648), .A2(n14560), .ZN(n13458) );
  OAI21_X1 U16811 ( .B1(n13459), .B2(n14560), .A(n13458), .ZN(P1_U3473) );
  AND3_X1 U16812 ( .A1(n20744), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n13460) );
  OAI21_X1 U16813 ( .B1(n13462), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13461), .ZN(n13522) );
  INV_X1 U16814 ( .A(n13522), .ZN(n13468) );
  AND2_X1 U16815 ( .A1(n16118), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13519) );
  AND2_X1 U16816 ( .A1(n13464), .A2(n20573), .ZN(n20739) );
  OR2_X1 U16817 ( .A1(n20739), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13465) );
  AND2_X2 U16818 ( .A1(n19869), .A2(n13465), .ZN(n16060) );
  INV_X1 U16819 ( .A(n16060), .ZN(n14973) );
  NAND2_X1 U16820 ( .A1(n20744), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15928) );
  NAND2_X1 U16821 ( .A1(n20742), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13466) );
  AND2_X1 U16822 ( .A1(n15928), .A2(n13466), .ZN(n13785) );
  AOI21_X1 U16823 ( .B1(n14973), .B2(n13785), .A(n14101), .ZN(n13467) );
  AOI211_X1 U16824 ( .C1(n13468), .C2(n16065), .A(n13519), .B(n13467), .ZN(
        n13469) );
  OAI21_X1 U16825 ( .B1(n14114), .B2(n20055), .A(n13469), .ZN(P1_U2999) );
  INV_X1 U16826 ( .A(n14560), .ZN(n20707) );
  INV_X1 U16827 ( .A(n20212), .ZN(n20458) );
  OR2_X1 U16828 ( .A1(n13470), .A2(n20458), .ZN(n13471) );
  XNOR2_X1 U16829 ( .A(n13471), .B(n13664), .ZN(n19933) );
  NAND2_X1 U16830 ( .A1(n14558), .A2(n13472), .ZN(n20710) );
  OR3_X1 U16831 ( .A1(n19933), .A2(n12512), .A3(n20710), .ZN(n13473) );
  OAI21_X1 U16832 ( .B1(n13664), .B2(n20707), .A(n13473), .ZN(P1_U3468) );
  OR2_X1 U16833 ( .A1(n13476), .A2(n13484), .ZN(n13486) );
  XNOR2_X1 U16834 ( .A(n13639), .B(n13474), .ZN(n13488) );
  XNOR2_X1 U16836 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13648), .ZN(
        n13481) );
  NOR2_X1 U16837 ( .A1(n13477), .A2(n11480), .ZN(n13479) );
  AND2_X1 U16838 ( .A1(n13479), .A2(n13478), .ZN(n13641) );
  INV_X1 U16839 ( .A(n13641), .ZN(n13480) );
  OAI22_X1 U16840 ( .A1(n13643), .A2(n13481), .B1(n13488), .B2(n13480), .ZN(
        n13482) );
  AOI21_X1 U16841 ( .B1(n13484), .B2(n13483), .A(n13482), .ZN(n13485) );
  NAND2_X1 U16842 ( .A1(n13486), .A2(n13485), .ZN(n13658) );
  INV_X1 U16843 ( .A(n20710), .ZN(n13487) );
  NAND2_X1 U16844 ( .A1(n13658), .A2(n13487), .ZN(n13494) );
  INV_X1 U16845 ( .A(n13489), .ZN(n13491) );
  OAI22_X1 U16846 ( .A1(n9844), .A2(n20705), .B1(n13491), .B2(n13490), .ZN(
        n13492) );
  NAND2_X1 U16847 ( .A1(n13492), .A2(n20707), .ZN(n13493) );
  OAI211_X1 U16848 ( .C1(n20707), .C2(n13474), .A(n13494), .B(n13493), .ZN(
        P1_U3472) );
  AOI22_X1 U16849 ( .A1(n19110), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19109), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13496) );
  NAND2_X1 U16850 ( .A1(n13496), .A2(n13495), .ZN(P2_U2974) );
  AOI22_X1 U16851 ( .A1(n19110), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19109), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13498) );
  NAND2_X1 U16852 ( .A1(n13498), .A2(n13497), .ZN(P2_U2973) );
  AOI22_X1 U16853 ( .A1(n19110), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19109), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n13500) );
  NAND2_X1 U16854 ( .A1(n13500), .A2(n13499), .ZN(P2_U2976) );
  AOI22_X1 U16855 ( .A1(n19110), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19109), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n13502) );
  NAND2_X1 U16856 ( .A1(n13502), .A2(n13501), .ZN(P2_U2967) );
  AOI22_X1 U16857 ( .A1(n19110), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19109), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13504) );
  NAND2_X1 U16858 ( .A1(n13504), .A2(n13503), .ZN(P2_U2969) );
  AOI22_X1 U16859 ( .A1(n19110), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19109), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13506) );
  NAND2_X1 U16860 ( .A1(n13506), .A2(n13505), .ZN(P2_U2968) );
  AOI22_X1 U16861 ( .A1(n19110), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19109), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13508) );
  NAND2_X1 U16862 ( .A1(n13508), .A2(n13507), .ZN(P2_U2972) );
  AOI22_X1 U16863 ( .A1(n19110), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19109), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13510) );
  NAND2_X1 U16864 ( .A1(n13510), .A2(n13509), .ZN(P2_U2978) );
  AOI22_X1 U16865 ( .A1(n19110), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n19109), .ZN(n13512) );
  NAND2_X1 U16866 ( .A1(n13512), .A2(n13511), .ZN(P2_U2965) );
  AOI22_X1 U16867 ( .A1(n19110), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19109), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n13514) );
  NAND2_X1 U16868 ( .A1(n13514), .A2(n13513), .ZN(P2_U2971) );
  AOI22_X1 U16869 ( .A1(n19110), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19109), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n13516) );
  NAND2_X1 U16870 ( .A1(n13516), .A2(n13515), .ZN(P2_U2970) );
  AOI21_X1 U16871 ( .B1(n15121), .B2(n13552), .A(n15119), .ZN(n13691) );
  INV_X1 U16872 ( .A(n15097), .ZN(n13551) );
  NOR3_X1 U16873 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15121), .A3(
        n13550), .ZN(n13517) );
  AOI21_X1 U16874 ( .B1(n13691), .B2(n13551), .A(n13517), .ZN(n13518) );
  INV_X1 U16875 ( .A(n13518), .ZN(n13521) );
  AOI21_X1 U16876 ( .B1(n16119), .B2(n14107), .A(n13519), .ZN(n13520) );
  OAI211_X1 U16877 ( .C1(n16137), .C2(n13522), .A(n13521), .B(n13520), .ZN(
        P1_U3031) );
  MUX2_X1 U16878 ( .A(n19139), .B(n14014), .S(n15347), .Z(n13525) );
  OAI21_X1 U16879 ( .B1(n19804), .B2(n15350), .A(n13525), .ZN(P2_U2885) );
  INV_X1 U16880 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19078) );
  NAND2_X1 U16881 ( .A1(n19110), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13527) );
  OAI211_X1 U16882 ( .C1(n19078), .C2(n13532), .A(n13527), .B(n13526), .ZN(
        P2_U2979) );
  INV_X1 U16883 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19086) );
  NAND2_X1 U16884 ( .A1(n19110), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13529) );
  OAI211_X1 U16885 ( .C1(n19086), .C2(n13532), .A(n13529), .B(n13528), .ZN(
        P2_U2975) );
  INV_X1 U16886 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19082) );
  NAND2_X1 U16887 ( .A1(n19110), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13531) );
  OAI211_X1 U16888 ( .C1(n19082), .C2(n13532), .A(n13531), .B(n13530), .ZN(
        P2_U2977) );
  NOR2_X1 U16889 ( .A1(n13534), .A2(n13533), .ZN(n13535) );
  XNOR2_X1 U16890 ( .A(n13536), .B(n11914), .ZN(n19969) );
  OAI222_X1 U16891 ( .A1(n19977), .A2(n19992), .B1(n9864), .B2(n19997), .C1(
        n19969), .C2(n19985), .ZN(P1_U2871) );
  NOR2_X1 U16892 ( .A1(n12870), .A2(n13618), .ZN(n13542) );
  AOI21_X1 U16893 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n13618), .A(n13542), .ZN(
        n13543) );
  OAI21_X1 U16894 ( .B1(n19795), .B2(n15350), .A(n13543), .ZN(P2_U2884) );
  XNOR2_X1 U16895 ( .A(n13545), .B(n13544), .ZN(n13791) );
  NAND3_X1 U16896 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n15121), .ZN(n13546) );
  OAI211_X1 U16897 ( .C1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n16092), .A(
        n13547), .B(n13546), .ZN(n13559) );
  XNOR2_X1 U16898 ( .A(n13549), .B(n13548), .ZN(n19967) );
  INV_X1 U16899 ( .A(n13550), .ZN(n13553) );
  OAI21_X1 U16900 ( .B1(n13553), .B2(n13552), .A(n13551), .ZN(n16099) );
  NAND3_X1 U16901 ( .A1(n16099), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n13554), .ZN(n13557) );
  NAND2_X1 U16902 ( .A1(n15121), .A2(n13706), .ZN(n13705) );
  INV_X1 U16903 ( .A(n13705), .ZN(n13555) );
  AND2_X1 U16904 ( .A1(n16118), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n13786) );
  NOR2_X1 U16905 ( .A1(n13555), .A2(n13786), .ZN(n13556) );
  OAI211_X1 U16906 ( .C1(n19967), .C2(n16136), .A(n13557), .B(n13556), .ZN(
        n13558) );
  AOI21_X1 U16907 ( .B1(n13559), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n13558), .ZN(n13560) );
  OAI21_X1 U16908 ( .B1(n13791), .B2(n16137), .A(n13560), .ZN(P1_U3029) );
  AND2_X1 U16909 ( .A1(n13562), .A2(n13563), .ZN(n13725) );
  NAND2_X1 U16910 ( .A1(n13562), .A2(n13564), .ZN(n13731) );
  OAI211_X1 U16911 ( .C1(n13725), .C2(n13565), .A(n13731), .B(n15342), .ZN(
        n13570) );
  NAND2_X1 U16912 ( .A1(n13726), .A2(n13566), .ZN(n13567) );
  NAND2_X1 U16913 ( .A1(n9682), .A2(n13567), .ZN(n16291) );
  INV_X1 U16914 ( .A(n16291), .ZN(n13568) );
  NAND2_X1 U16915 ( .A1(n13568), .A2(n15316), .ZN(n13569) );
  OAI211_X1 U16916 ( .C1(n15316), .C2(n9890), .A(n13570), .B(n13569), .ZN(
        P2_U2877) );
  AND2_X1 U16917 ( .A1(n13562), .A2(n13571), .ZN(n13723) );
  XNOR2_X1 U16918 ( .A(n13723), .B(n13722), .ZN(n13576) );
  AND2_X1 U16919 ( .A1(n13697), .A2(n13572), .ZN(n13573) );
  OR2_X1 U16920 ( .A1(n13573), .A2(n13728), .ZN(n16239) );
  INV_X1 U16921 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n13574) );
  MUX2_X1 U16922 ( .A(n16239), .B(n13574), .S(n15347), .Z(n13575) );
  OAI21_X1 U16923 ( .B1(n13576), .B2(n15350), .A(n13575), .ZN(P2_U2879) );
  INV_X1 U16924 ( .A(n13580), .ZN(n13578) );
  NAND2_X1 U16925 ( .A1(n13579), .A2(n13578), .ZN(n13581) );
  NAND2_X1 U16926 ( .A1(n13562), .A2(n13580), .ZN(n13614) );
  OAI21_X1 U16927 ( .B1(n13577), .B2(n13581), .A(n13614), .ZN(n19043) );
  NOR2_X1 U16928 ( .A1(n13583), .A2(n13582), .ZN(n13584) );
  OR2_X1 U16929 ( .A1(n9693), .A2(n13584), .ZN(n19115) );
  MUX2_X1 U16930 ( .A(n19115), .B(n13585), .S(n15347), .Z(n13586) );
  OAI21_X1 U16931 ( .B1(n19043), .B2(n15350), .A(n13586), .ZN(P2_U2883) );
  INV_X2 U16932 ( .A(n13587), .ZN(n20050) );
  AOI22_X1 U16933 ( .A1(n20050), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20049), .ZN(n13592) );
  NAND2_X1 U16934 ( .A1(n20054), .A2(DATAI_6_), .ZN(n13590) );
  NAND2_X1 U16935 ( .A1(n20053), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13589) );
  AND2_X1 U16936 ( .A1(n13590), .A2(n13589), .ZN(n20099) );
  INV_X1 U16937 ( .A(n20099), .ZN(n13591) );
  NAND2_X1 U16938 ( .A1(n20037), .A2(n13591), .ZN(n13939) );
  NAND2_X1 U16939 ( .A1(n13592), .A2(n13939), .ZN(P1_U2958) );
  AOI22_X1 U16940 ( .A1(n20050), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20049), .ZN(n13595) );
  NAND2_X1 U16941 ( .A1(n20054), .A2(DATAI_5_), .ZN(n13594) );
  NAND2_X1 U16942 ( .A1(n20053), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13593) );
  AND2_X1 U16943 ( .A1(n13594), .A2(n13593), .ZN(n20095) );
  INV_X1 U16944 ( .A(n20095), .ZN(n14833) );
  NAND2_X1 U16945 ( .A1(n20037), .A2(n14833), .ZN(n13929) );
  NAND2_X1 U16946 ( .A1(n13595), .A2(n13929), .ZN(P1_U2957) );
  INV_X1 U16947 ( .A(n13596), .ZN(n20049) );
  AOI22_X1 U16948 ( .A1(n20050), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20049), .ZN(n13599) );
  INV_X1 U16949 ( .A(DATAI_11_), .ZN(n13598) );
  NAND2_X1 U16950 ( .A1(n20053), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13597) );
  OAI21_X1 U16951 ( .B1(n20053), .B2(n13598), .A(n13597), .ZN(n14806) );
  NAND2_X1 U16952 ( .A1(n20037), .A2(n14806), .ZN(n13935) );
  NAND2_X1 U16953 ( .A1(n13599), .A2(n13935), .ZN(P1_U2963) );
  AOI22_X1 U16954 ( .A1(n20050), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20049), .ZN(n13603) );
  NAND2_X1 U16955 ( .A1(n20054), .A2(DATAI_7_), .ZN(n13601) );
  NAND2_X1 U16956 ( .A1(n20053), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13600) );
  AND2_X1 U16957 ( .A1(n13601), .A2(n13600), .ZN(n20107) );
  INV_X1 U16958 ( .A(n20107), .ZN(n13602) );
  NAND2_X1 U16959 ( .A1(n20037), .A2(n13602), .ZN(n13931) );
  NAND2_X1 U16960 ( .A1(n13603), .A2(n13931), .ZN(P1_U2959) );
  OR2_X1 U16961 ( .A1(n13735), .A2(n13604), .ZN(n13606) );
  NAND2_X1 U16962 ( .A1(n13606), .A2(n13605), .ZN(n16191) );
  INV_X1 U16963 ( .A(n13732), .ZN(n13607) );
  NOR2_X1 U16964 ( .A1(n13731), .A2(n13607), .ZN(n13610) );
  OAI211_X1 U16965 ( .C1(n13610), .C2(n13609), .A(n13608), .B(n15342), .ZN(
        n13612) );
  NAND2_X1 U16966 ( .A1(n15347), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13611) );
  OAI211_X1 U16967 ( .C1(n16191), .C2(n13618), .A(n13612), .B(n13611), .ZN(
        P2_U2875) );
  OAI21_X1 U16968 ( .B1(n9693), .B2(n13613), .A(n13715), .ZN(n14204) );
  INV_X1 U16969 ( .A(n13614), .ZN(n13615) );
  OR2_X1 U16970 ( .A1(n13614), .A2(n14295), .ZN(n13713) );
  OAI211_X1 U16971 ( .C1(n13615), .C2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n15342), .B(n13713), .ZN(n13617) );
  NAND2_X1 U16972 ( .A1(n15347), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n13616) );
  OAI211_X1 U16973 ( .C1(n14204), .C2(n13618), .A(n13617), .B(n13616), .ZN(
        P2_U2882) );
  NAND2_X1 U16974 ( .A1(n11482), .A2(n12000), .ZN(n13619) );
  NAND2_X1 U16975 ( .A1(n20054), .A2(DATAI_1_), .ZN(n13621) );
  NAND2_X1 U16976 ( .A1(n20053), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13620) );
  AND2_X1 U16977 ( .A1(n13621), .A2(n13620), .ZN(n20078) );
  OAI222_X1 U16978 ( .A1(n14869), .A2(n19977), .B1(n14867), .B2(n12009), .C1(
        n14866), .C2(n20078), .ZN(P1_U2903) );
  AOI22_X1 U16979 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13622) );
  OAI21_X1 U16980 ( .B1(n14822), .B2(n13633), .A(n13622), .ZN(P1_U2913) );
  INV_X1 U16981 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13624) );
  AOI22_X1 U16982 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13623) );
  OAI21_X1 U16983 ( .B1(n13624), .B2(n13633), .A(n13623), .ZN(P1_U2915) );
  INV_X1 U16984 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13626) );
  AOI22_X1 U16985 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13625) );
  OAI21_X1 U16986 ( .B1(n13626), .B2(n13633), .A(n13625), .ZN(P1_U2916) );
  AOI22_X1 U16987 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13627) );
  OAI21_X1 U16988 ( .B1(n14826), .B2(n13633), .A(n13627), .ZN(P1_U2914) );
  AOI22_X1 U16989 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13628) );
  OAI21_X1 U16990 ( .B1(n14847), .B2(n13633), .A(n13628), .ZN(P1_U2918) );
  INV_X1 U16991 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13630) );
  AOI22_X1 U16992 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13629) );
  OAI21_X1 U16993 ( .B1(n13630), .B2(n13633), .A(n13629), .ZN(P1_U2919) );
  AOI22_X1 U16994 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13631) );
  OAI21_X1 U16995 ( .B1(n14843), .B2(n13633), .A(n13631), .ZN(P1_U2917) );
  INV_X1 U16996 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13634) );
  AOI22_X1 U16997 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13632) );
  OAI21_X1 U16998 ( .B1(n13634), .B2(n13633), .A(n13632), .ZN(P1_U2920) );
  NAND2_X1 U16999 ( .A1(n13639), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13635) );
  NAND2_X1 U17000 ( .A1(n13635), .A2(n20708), .ZN(n13636) );
  INV_X1 U17001 ( .A(n13638), .ZN(n13646) );
  MUX2_X1 U17002 ( .A(n13640), .B(n11321), .S(n13639), .Z(n13642) );
  OAI21_X1 U17003 ( .B1(n13638), .B2(n13642), .A(n13641), .ZN(n13650) );
  INV_X1 U17004 ( .A(n13643), .ZN(n15903) );
  NAND2_X1 U17005 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13644) );
  NAND2_X1 U17006 ( .A1(n13644), .A2(n20708), .ZN(n13645) );
  NAND2_X1 U17007 ( .A1(n13646), .A2(n13645), .ZN(n13647) );
  OAI211_X1 U17008 ( .C1(n20708), .C2(n13648), .A(n15903), .B(n13647), .ZN(
        n13649) );
  OAI211_X1 U17009 ( .C1(n14555), .C2(n13651), .A(n13650), .B(n13649), .ZN(
        n13652) );
  AOI21_X1 U17010 ( .B1(n20717), .B2(n14555), .A(n13652), .ZN(n20711) );
  OR2_X1 U17011 ( .A1(n20711), .A2(n13665), .ZN(n13654) );
  NAND2_X1 U17012 ( .A1(n13665), .A2(n20708), .ZN(n13653) );
  NAND2_X1 U17013 ( .A1(n13654), .A2(n13653), .ZN(n15913) );
  NAND2_X1 U17014 ( .A1(n15913), .A2(n16149), .ZN(n13656) );
  AND2_X1 U17015 ( .A1(n19870), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13668) );
  NAND2_X1 U17016 ( .A1(n20708), .A2(n13668), .ZN(n13655) );
  NAND2_X1 U17017 ( .A1(n13656), .A2(n13655), .ZN(n13662) );
  NAND2_X1 U17018 ( .A1(n13665), .A2(n13474), .ZN(n13657) );
  OAI21_X1 U17019 ( .B1(n13658), .B2(n13665), .A(n13657), .ZN(n15912) );
  NAND2_X1 U17020 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n13668), .ZN(
        n13660) );
  OAI21_X1 U17021 ( .B1(n15912), .B2(P1_STATE2_REG_1__SCAN_IN), .A(n13660), 
        .ZN(n13661) );
  NAND2_X1 U17022 ( .A1(n13662), .A2(n13661), .ZN(n15922) );
  OR2_X1 U17023 ( .A1(n15922), .A2(n13663), .ZN(n13675) );
  INV_X1 U17024 ( .A(n13665), .ZN(n15901) );
  OAI21_X1 U17025 ( .B1(n19933), .B2(n12512), .A(n15901), .ZN(n13667) );
  AOI21_X1 U17026 ( .B1(n13665), .B2(n13664), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n13666) );
  NAND2_X1 U17027 ( .A1(n13667), .A2(n13666), .ZN(n13670) );
  NAND2_X1 U17028 ( .A1(n13668), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13669) );
  NAND2_X1 U17029 ( .A1(n13670), .A2(n13669), .ZN(n15921) );
  NOR2_X1 U17030 ( .A1(n15921), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n13671) );
  AOI21_X1 U17031 ( .B1(n13675), .B2(n13671), .A(n16150), .ZN(n13673) );
  NOR2_X1 U17032 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20748) );
  NOR2_X1 U17033 ( .A1(n15921), .A2(n16145), .ZN(n13674) );
  NAND2_X1 U17034 ( .A1(n13675), .A2(n13674), .ZN(n15938) );
  INV_X1 U17035 ( .A(n15938), .ZN(n13678) );
  NOR2_X1 U17036 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n16149), .ZN(n20715) );
  INV_X1 U17037 ( .A(n9594), .ZN(n13676) );
  OAI22_X1 U17038 ( .A1(n12013), .A2(n20573), .B1(n20715), .B2(n13676), .ZN(
        n13677) );
  OAI21_X1 U17039 ( .B1(n13678), .B2(n13677), .A(n20725), .ZN(n13679) );
  OAI21_X1 U17040 ( .B1(n20725), .B2(n20499), .A(n13679), .ZN(P1_U3478) );
  INV_X1 U17041 ( .A(n9595), .ZN(n13682) );
  NAND2_X1 U17042 ( .A1(n20718), .A2(n20742), .ZN(n13681) );
  OAI22_X1 U17043 ( .A1(n13682), .A2(n13681), .B1(n20715), .B2(n20537), .ZN(
        n13683) );
  OAI21_X1 U17044 ( .B1(n10125), .B2(n13683), .A(n20725), .ZN(n13684) );
  OAI21_X1 U17045 ( .B1(n20386), .B2(n20725), .A(n13684), .ZN(P1_U3477) );
  NAND2_X1 U17046 ( .A1(n9595), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20428) );
  NAND2_X1 U17047 ( .A1(n20428), .A2(n20718), .ZN(n13685) );
  OR2_X1 U17048 ( .A1(n20428), .A2(n20573), .ZN(n20712) );
  MUX2_X1 U17049 ( .A(n13685), .B(n20712), .S(n11999), .Z(n13686) );
  OAI21_X1 U17050 ( .B1(n20715), .B2(n13476), .A(n13686), .ZN(n13687) );
  NAND2_X1 U17051 ( .A1(n20725), .A2(n13687), .ZN(n13688) );
  OAI21_X1 U17052 ( .B1(n20725), .B2(n11803), .A(n13688), .ZN(P1_U3476) );
  XOR2_X1 U17053 ( .A(n13689), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n14031) );
  INV_X1 U17054 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20729) );
  OAI22_X1 U17055 ( .A1(n16136), .A2(n19969), .B1(n20729), .B2(n16134), .ZN(
        n13695) );
  NOR2_X1 U17056 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15097), .ZN(
        n13690) );
  NOR2_X1 U17057 ( .A1(n16071), .A2(n13690), .ZN(n13693) );
  INV_X1 U17058 ( .A(n13691), .ZN(n13692) );
  MUX2_X1 U17059 ( .A(n13693), .B(n13692), .S(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n13694) );
  AOI211_X1 U17060 ( .C1(n16122), .C2(n14031), .A(n13695), .B(n13694), .ZN(
        n13696) );
  INV_X1 U17061 ( .A(n13696), .ZN(P1_U3030) );
  OAI21_X1 U17062 ( .B1(n10801), .B2(n10136), .A(n13697), .ZN(n18979) );
  INV_X1 U17063 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14291) );
  NOR2_X1 U17064 ( .A1(n13713), .A2(n14291), .ZN(n13699) );
  INV_X1 U17065 ( .A(n13723), .ZN(n13698) );
  OAI211_X1 U17066 ( .C1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .C2(n13699), .A(
        n13698), .B(n15342), .ZN(n13701) );
  NAND2_X1 U17067 ( .A1(n15347), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n13700) );
  OAI211_X1 U17068 ( .C1(n18979), .C2(n15347), .A(n13701), .B(n13700), .ZN(
        P2_U2880) );
  XNOR2_X1 U17069 ( .A(n13703), .B(n13702), .ZN(n13862) );
  NOR2_X1 U17070 ( .A1(n16092), .A2(n13796), .ZN(n13704) );
  NOR2_X1 U17071 ( .A1(n13704), .A2(n15119), .ZN(n14220) );
  NAND2_X1 U17072 ( .A1(n14220), .A2(n13705), .ZN(n13770) );
  AOI21_X1 U17073 ( .B1(n13796), .B2(n16099), .A(n15121), .ZN(n15145) );
  NOR2_X1 U17074 ( .A1(n13706), .A2(n15145), .ZN(n14152) );
  AOI22_X1 U17075 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13770), .B1(
        n14152), .B2(n11880), .ZN(n13712) );
  OR2_X1 U17076 ( .A1(n13708), .A2(n13707), .ZN(n13709) );
  NAND2_X1 U17077 ( .A1(n13772), .A2(n13709), .ZN(n19954) );
  INV_X1 U17078 ( .A(n19954), .ZN(n13710) );
  INV_X1 U17079 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20657) );
  NOR2_X1 U17080 ( .A1(n16134), .A2(n20657), .ZN(n13857) );
  AOI21_X1 U17081 ( .B1(n13710), .B2(n16119), .A(n13857), .ZN(n13711) );
  OAI211_X1 U17082 ( .C1(n13862), .C2(n16137), .A(n13712), .B(n13711), .ZN(
        P1_U3028) );
  XOR2_X1 U17083 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B(n13713), .Z(n13720)
         );
  NAND2_X1 U17084 ( .A1(n13715), .A2(n13714), .ZN(n13716) );
  NAND2_X1 U17085 ( .A1(n13717), .A2(n13716), .ZN(n16246) );
  NOR2_X1 U17086 ( .A1(n16246), .A2(n13618), .ZN(n13718) );
  AOI21_X1 U17087 ( .B1(P2_EBX_REG_6__SCAN_IN), .B2(n13618), .A(n13718), .ZN(
        n13719) );
  OAI21_X1 U17088 ( .B1(n13720), .B2(n15350), .A(n13719), .ZN(P2_U2881) );
  AOI21_X1 U17089 ( .B1(n13723), .B2(n13722), .A(n13721), .ZN(n13724) );
  OR3_X1 U17090 ( .A1(n13725), .A2(n13724), .A3(n15350), .ZN(n13730) );
  OAI21_X1 U17091 ( .B1(n13728), .B2(n13727), .A(n13726), .ZN(n18964) );
  INV_X1 U17092 ( .A(n18964), .ZN(n16224) );
  NAND2_X1 U17093 ( .A1(n16224), .A2(n15316), .ZN(n13729) );
  OAI211_X1 U17094 ( .C1(n15316), .C2(n10629), .A(n13730), .B(n13729), .ZN(
        P2_U2878) );
  XOR2_X1 U17095 ( .A(n13732), .B(n13731), .Z(n13738) );
  AND2_X1 U17096 ( .A1(n9682), .A2(n13733), .ZN(n13734) );
  OR2_X1 U17097 ( .A1(n13735), .A2(n13734), .ZN(n15771) );
  MUX2_X1 U17098 ( .A(n15771), .B(n13736), .S(n15347), .Z(n13737) );
  OAI21_X1 U17099 ( .B1(n13738), .B2(n15350), .A(n13737), .ZN(P2_U2876) );
  XNOR2_X1 U17100 ( .A(n13739), .B(n13740), .ZN(n19962) );
  NAND2_X1 U17101 ( .A1(n20054), .A2(DATAI_2_), .ZN(n13742) );
  NAND2_X1 U17102 ( .A1(n20053), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13741) );
  AND2_X1 U17103 ( .A1(n13742), .A2(n13741), .ZN(n20082) );
  OAI222_X1 U17104 ( .A1(n14869), .A2(n19962), .B1(n14867), .B2(n12002), .C1(
        n14866), .C2(n20082), .ZN(P1_U2902) );
  OAI222_X1 U17105 ( .A1(n19967), .A2(n19985), .B1(n19997), .B2(n11876), .C1(
        n19962), .C2(n19992), .ZN(P1_U2870) );
  NAND2_X1 U17106 ( .A1(n13743), .A2(n13605), .ZN(n13745) );
  INV_X1 U17107 ( .A(n13837), .ZN(n13744) );
  AND2_X1 U17108 ( .A1(n13745), .A2(n13744), .ZN(n16186) );
  INV_X1 U17109 ( .A(n16186), .ZN(n16280) );
  INV_X1 U17110 ( .A(n13608), .ZN(n13748) );
  INV_X1 U17111 ( .A(n13746), .ZN(n13747) );
  OAI211_X1 U17112 ( .C1(n13748), .C2(n9679), .A(n13747), .B(n15342), .ZN(
        n13750) );
  NAND2_X1 U17113 ( .A1(n15347), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13749) );
  OAI211_X1 U17114 ( .C1(n16280), .C2(n15347), .A(n13750), .B(n13749), .ZN(
        P2_U2874) );
  NAND2_X1 U17115 ( .A1(n13752), .A2(n13751), .ZN(n13755) );
  INV_X1 U17116 ( .A(n13753), .ZN(n13754) );
  AND2_X1 U17117 ( .A1(n13755), .A2(n13754), .ZN(n19806) );
  XNOR2_X1 U17118 ( .A(n19804), .B(n19806), .ZN(n13762) );
  XNOR2_X1 U17119 ( .A(n13757), .B(n13756), .ZN(n19820) );
  INV_X1 U17120 ( .A(n19820), .ZN(n13758) );
  NAND2_X1 U17121 ( .A1(n19816), .A2(n13758), .ZN(n13759) );
  OAI21_X1 U17122 ( .B1(n19816), .B2(n13758), .A(n13759), .ZN(n19058) );
  NOR2_X1 U17123 ( .A1(n19058), .A2(n19059), .ZN(n19057) );
  INV_X1 U17124 ( .A(n13759), .ZN(n13760) );
  NOR2_X1 U17125 ( .A1(n19057), .A2(n13760), .ZN(n13761) );
  NOR2_X1 U17126 ( .A1(n13761), .A2(n13762), .ZN(n14118) );
  AOI21_X1 U17127 ( .B1(n13762), .B2(n13761), .A(n14118), .ZN(n13766) );
  AOI22_X1 U17128 ( .A1(n19033), .A2(n16168), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19055), .ZN(n13765) );
  INV_X1 U17129 ( .A(n19806), .ZN(n13763) );
  NAND2_X1 U17130 ( .A1(n13763), .A2(n19056), .ZN(n13764) );
  OAI211_X1 U17131 ( .C1(n13766), .C2(n19060), .A(n13765), .B(n13764), .ZN(
        P2_U2917) );
  XNOR2_X1 U17132 ( .A(n13768), .B(n13767), .ZN(n14010) );
  AOI21_X1 U17133 ( .B1(n11680), .B2(n11880), .A(n13797), .ZN(n13769) );
  AOI22_X1 U17134 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13770), .B1(
        n14152), .B2(n13769), .ZN(n13776) );
  NAND2_X1 U17135 ( .A1(n13772), .A2(n13771), .ZN(n13773) );
  AND2_X1 U17136 ( .A1(n16128), .A2(n13773), .ZN(n19990) );
  INV_X1 U17137 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n13774) );
  NOR2_X1 U17138 ( .A1(n16134), .A2(n13774), .ZN(n14005) );
  AOI21_X1 U17139 ( .B1(n19990), .B2(n16119), .A(n14005), .ZN(n13775) );
  OAI211_X1 U17140 ( .C1(n14010), .C2(n16137), .A(n13776), .B(n13775), .ZN(
        P1_U3027) );
  OAI21_X1 U17141 ( .B1(n13777), .B2(n13780), .A(n13779), .ZN(n19950) );
  NAND2_X1 U17142 ( .A1(n20054), .A2(DATAI_3_), .ZN(n13782) );
  NAND2_X1 U17143 ( .A1(n20053), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13781) );
  AND2_X1 U17144 ( .A1(n13782), .A2(n13781), .ZN(n20086) );
  OAI222_X1 U17145 ( .A1(n14869), .A2(n19950), .B1(n14867), .B2(n12029), .C1(
        n14866), .C2(n20086), .ZN(P1_U2901) );
  NAND2_X1 U17146 ( .A1(n20054), .A2(DATAI_0_), .ZN(n13784) );
  NAND2_X1 U17147 ( .A1(n20053), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13783) );
  AND2_X1 U17148 ( .A1(n13784), .A2(n13783), .ZN(n20069) );
  OAI222_X1 U17149 ( .A1(n14866), .A2(n20069), .B1(n14869), .B2(n14114), .C1(
        n12015), .C2(n14867), .ZN(P1_U2904) );
  INV_X1 U17150 ( .A(n19962), .ZN(n13789) );
  INV_X1 U17151 ( .A(n20055), .ZN(n16066) );
  AOI21_X1 U17152 ( .B1(n16060), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n13786), .ZN(n13787) );
  OAI21_X1 U17153 ( .B1(n16069), .B2(n19956), .A(n13787), .ZN(n13788) );
  AOI21_X1 U17154 ( .B1(n13789), .B2(n16066), .A(n13788), .ZN(n13790) );
  OAI21_X1 U17155 ( .B1(n19869), .B2(n13791), .A(n13790), .ZN(P1_U2997) );
  XNOR2_X1 U17156 ( .A(n13794), .B(n13793), .ZN(n14027) );
  AOI21_X1 U17157 ( .B1(n15121), .B2(n13795), .A(n15119), .ZN(n16097) );
  OAI221_X1 U17158 ( .B1(n16092), .B2(n13796), .C1(n16092), .C2(n13797), .A(
        n16097), .ZN(n14150) );
  AND2_X1 U17159 ( .A1(n20852), .A2(n13797), .ZN(n14151) );
  AOI22_X1 U17160 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14150), .B1(
        n14152), .B2(n14151), .ZN(n13799) );
  XNOR2_X1 U17161 ( .A(n16128), .B(n16130), .ZN(n19922) );
  INV_X1 U17162 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n19926) );
  NOR2_X1 U17163 ( .A1(n16134), .A2(n19926), .ZN(n14022) );
  AOI21_X1 U17164 ( .B1(n19922), .B2(n16119), .A(n14022), .ZN(n13798) );
  OAI211_X1 U17165 ( .C1(n14027), .C2(n16137), .A(n13799), .B(n13798), .ZN(
        P1_U3026) );
  INV_X1 U17166 ( .A(n19950), .ZN(n13860) );
  INV_X1 U17167 ( .A(n19992), .ZN(n16014) );
  INV_X1 U17168 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13800) );
  OAI22_X1 U17169 ( .A1(n19954), .A2(n19985), .B1(n13800), .B2(n19997), .ZN(
        n13801) );
  AOI21_X1 U17170 ( .B1(n13860), .B2(n16014), .A(n13801), .ZN(n13802) );
  INV_X1 U17171 ( .A(n13802), .ZN(P1_U2869) );
  AND2_X1 U17172 ( .A1(n13779), .A2(n13805), .ZN(n13806) );
  OR2_X1 U17173 ( .A1(n13804), .A2(n13806), .ZN(n19993) );
  INV_X1 U17174 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n13809) );
  NAND2_X1 U17175 ( .A1(n20054), .A2(DATAI_4_), .ZN(n13808) );
  NAND2_X1 U17176 ( .A1(n20053), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13807) );
  AND2_X1 U17177 ( .A1(n13808), .A2(n13807), .ZN(n20090) );
  OAI222_X1 U17178 ( .A1(n19993), .A2(n14869), .B1(n13809), .B2(n14867), .C1(
        n14866), .C2(n20090), .ZN(P1_U2900) );
  INV_X1 U17179 ( .A(n13988), .ZN(n13810) );
  NAND2_X1 U17180 ( .A1(n13811), .A2(n13810), .ZN(n13814) );
  XOR2_X1 U17181 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n13812), .Z(
        n13813) );
  XNOR2_X1 U17182 ( .A(n13814), .B(n13813), .ZN(n13835) );
  XOR2_X1 U17183 ( .A(n13816), .B(n13815), .Z(n13833) );
  NOR2_X1 U17184 ( .A1(n15534), .A2(n13817), .ZN(n13829) );
  NOR2_X1 U17185 ( .A1(n16265), .A2(n13984), .ZN(n13818) );
  AOI211_X1 U17186 ( .C1(n16255), .C2(n13982), .A(n13829), .B(n13818), .ZN(
        n13819) );
  OAI21_X1 U17187 ( .B1(n13541), .B2(n16247), .A(n13819), .ZN(n13820) );
  AOI21_X1 U17188 ( .B1(n13833), .B2(n19118), .A(n13820), .ZN(n13821) );
  OAI21_X1 U17189 ( .B1(n16258), .B2(n13835), .A(n13821), .ZN(P2_U3011) );
  OR2_X1 U17190 ( .A1(n13823), .A2(n13822), .ZN(n13825) );
  NAND2_X1 U17191 ( .A1(n13825), .A2(n13824), .ZN(n14119) );
  INV_X1 U17192 ( .A(n13826), .ZN(n13828) );
  MUX2_X1 U17193 ( .A(n13828), .B(n13827), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n13831) );
  AOI21_X1 U17194 ( .B1(n16302), .B2(n10350), .A(n13829), .ZN(n13830) );
  OAI211_X1 U17195 ( .C1(n14119), .C2(n19143), .A(n13831), .B(n13830), .ZN(
        n13832) );
  AOI21_X1 U17196 ( .B1(n13833), .B2(n16271), .A(n13832), .ZN(n13834) );
  OAI21_X1 U17197 ( .B1(n19133), .B2(n13835), .A(n13834), .ZN(P2_U3043) );
  XNOR2_X1 U17198 ( .A(n13746), .B(n13836), .ZN(n13840) );
  OAI21_X1 U17199 ( .B1(n13838), .B2(n13837), .A(n13958), .ZN(n18952) );
  MUX2_X1 U17200 ( .A(n10659), .B(n18952), .S(n15316), .Z(n13839) );
  OAI21_X1 U17201 ( .B1(n13840), .B2(n15350), .A(n13839), .ZN(P2_U2873) );
  OAI21_X1 U17202 ( .B1(n13804), .B2(n13842), .A(n13841), .ZN(n19924) );
  AOI22_X1 U17203 ( .A1(n19922), .A2(n12508), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n12469), .ZN(n13843) );
  OAI21_X1 U17204 ( .B1(n19924), .B2(n19992), .A(n13843), .ZN(P1_U2867) );
  OAI21_X1 U17205 ( .B1(n13844), .B2(n13846), .A(n13845), .ZN(n19027) );
  AOI21_X1 U17206 ( .B1(n16199), .B2(n13847), .A(n13914), .ZN(n13848) );
  OAI221_X1 U17207 ( .B1(n9951), .B2(n13848), .C1(n9949), .C2(n16199), .A(
        n18984), .ZN(n13856) );
  INV_X1 U17208 ( .A(n15771), .ZN(n16203) );
  OAI22_X1 U17209 ( .A1(n16206), .A2(n18974), .B1(n10812), .B2(n18987), .ZN(
        n13854) );
  INV_X1 U17210 ( .A(n18992), .ZN(n15201) );
  INV_X1 U17211 ( .A(n13849), .ZN(n13851) );
  NAND3_X1 U17212 ( .A1(n13851), .A2(n13236), .A3(n13850), .ZN(n13852) );
  OAI211_X1 U17213 ( .C1(n15201), .C2(n13736), .A(n13852), .B(n15534), .ZN(
        n13853) );
  AOI211_X1 U17214 ( .C1(n16203), .C2(n18999), .A(n13854), .B(n13853), .ZN(
        n13855) );
  OAI211_X1 U17215 ( .C1(n19027), .C2(n18989), .A(n13856), .B(n13855), .ZN(
        P2_U2844) );
  AOI21_X1 U17216 ( .B1(n16060), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n13857), .ZN(n13858) );
  OAI21_X1 U17217 ( .B1(n16069), .B2(n19949), .A(n13858), .ZN(n13859) );
  AOI21_X1 U17218 ( .B1(n13860), .B2(n16066), .A(n13859), .ZN(n13861) );
  OAI21_X1 U17219 ( .B1(n19869), .B2(n13862), .A(n13861), .ZN(P1_U2996) );
  NOR2_X1 U17220 ( .A1(n9951), .A2(n13863), .ZN(n13864) );
  XNOR2_X1 U17221 ( .A(n13864), .B(n16245), .ZN(n13865) );
  NAND2_X1 U17222 ( .A1(n13865), .A2(n18984), .ZN(n13876) );
  INV_X1 U17223 ( .A(n14352), .ZN(n13866) );
  OR2_X1 U17224 ( .A1(n13867), .A2(n13866), .ZN(n13870) );
  INV_X1 U17225 ( .A(n13868), .ZN(n13869) );
  NAND2_X1 U17226 ( .A1(n13870), .A2(n13869), .ZN(n19036) );
  AOI22_X1 U17227 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19000), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n18951), .ZN(n13871) );
  OAI211_X1 U17228 ( .C1(n18989), .C2(n19036), .A(n13871), .B(n15534), .ZN(
        n13873) );
  NOR2_X1 U17229 ( .A1(n15201), .A2(n13574), .ZN(n13872) );
  AOI211_X1 U17230 ( .C1(n13236), .C2(n13874), .A(n13873), .B(n13872), .ZN(
        n13875) );
  OAI211_X1 U17231 ( .C1(n16239), .C2(n18978), .A(n13876), .B(n13875), .ZN(
        P2_U2847) );
  NOR2_X1 U17232 ( .A1(n9951), .A2(n13877), .ZN(n13878) );
  XNOR2_X1 U17233 ( .A(n13878), .B(n16220), .ZN(n13879) );
  NAND2_X1 U17234 ( .A1(n13879), .A2(n18984), .ZN(n13888) );
  INV_X1 U17235 ( .A(n13880), .ZN(n13881) );
  XNOR2_X1 U17236 ( .A(n13882), .B(n13881), .ZN(n19030) );
  AOI22_X1 U17237 ( .A1(P2_EBX_REG_10__SCAN_IN), .A2(n18992), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19000), .ZN(n13883) );
  OAI211_X1 U17238 ( .C1(n18989), .C2(n19030), .A(n13883), .B(n15534), .ZN(
        n13886) );
  NOR2_X1 U17239 ( .A1(n13884), .A2(n18995), .ZN(n13885) );
  AOI211_X1 U17240 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n18951), .A(n13886), 
        .B(n13885), .ZN(n13887) );
  OAI211_X1 U17241 ( .C1(n16291), .C2(n18978), .A(n13888), .B(n13887), .ZN(
        P2_U2845) );
  NOR2_X1 U17242 ( .A1(n9951), .A2(n13889), .ZN(n13890) );
  XNOR2_X1 U17243 ( .A(n13890), .B(n16253), .ZN(n13891) );
  NAND2_X1 U17244 ( .A1(n13891), .A2(n18984), .ZN(n13899) );
  XNOR2_X1 U17245 ( .A(n13892), .B(n13893), .ZN(n19039) );
  AOI22_X1 U17246 ( .A1(P2_EBX_REG_6__SCAN_IN), .A2(n18992), .B1(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19000), .ZN(n13894) );
  OAI211_X1 U17247 ( .C1(n18989), .C2(n19039), .A(n13894), .B(n15534), .ZN(
        n13897) );
  NOR2_X1 U17248 ( .A1(n13895), .A2(n18995), .ZN(n13896) );
  AOI211_X1 U17249 ( .C1(P2_REIP_REG_6__SCAN_IN), .C2(n18951), .A(n13897), .B(
        n13896), .ZN(n13898) );
  OAI211_X1 U17250 ( .C1(n16246), .C2(n18978), .A(n13899), .B(n13898), .ZN(
        P2_U2849) );
  INV_X1 U17251 ( .A(n19124), .ZN(n13903) );
  NOR2_X1 U17252 ( .A1(n9951), .A2(n13900), .ZN(n13902) );
  AOI21_X1 U17253 ( .B1(n13903), .B2(n13902), .A(n19717), .ZN(n13901) );
  OAI21_X1 U17254 ( .B1(n13903), .B2(n13902), .A(n13901), .ZN(n13912) );
  XNOR2_X1 U17255 ( .A(n13824), .B(n13904), .ZN(n14121) );
  OAI21_X1 U17256 ( .B1(n18974), .B2(n10785), .A(n15534), .ZN(n13905) );
  AOI21_X1 U17257 ( .B1(n18954), .B2(n14121), .A(n13905), .ZN(n13907) );
  NAND2_X1 U17258 ( .A1(n18992), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n13906) );
  OAI211_X1 U17259 ( .C1(n18987), .C2(n11084), .A(n13907), .B(n13906), .ZN(
        n13909) );
  NOR2_X1 U17260 ( .A1(n19115), .A2(n18978), .ZN(n13908) );
  AOI211_X1 U17261 ( .C1(n13236), .C2(n13910), .A(n13909), .B(n13908), .ZN(
        n13911) );
  OAI211_X1 U17262 ( .C1(n18985), .C2(n19043), .A(n13912), .B(n13911), .ZN(
        P2_U2851) );
  XNOR2_X1 U17263 ( .A(n13845), .B(n13913), .ZN(n19025) );
  NOR2_X1 U17264 ( .A1(n9951), .A2(n13914), .ZN(n13915) );
  XNOR2_X1 U17265 ( .A(n16198), .B(n13915), .ZN(n13916) );
  NAND2_X1 U17266 ( .A1(n13916), .A2(n18984), .ZN(n13924) );
  INV_X1 U17267 ( .A(n16191), .ZN(n13922) );
  INV_X1 U17268 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n13917) );
  OAI22_X1 U17269 ( .A1(n13917), .A2(n18974), .B1(n11176), .B2(n18987), .ZN(
        n13921) );
  AOI21_X1 U17270 ( .B1(n18992), .B2(P2_EBX_REG_12__SCAN_IN), .A(n16279), .ZN(
        n13918) );
  OAI21_X1 U17271 ( .B1(n13919), .B2(n18995), .A(n13918), .ZN(n13920) );
  AOI211_X1 U17272 ( .C1(n13922), .C2(n18999), .A(n13921), .B(n13920), .ZN(
        n13923) );
  OAI211_X1 U17273 ( .C1(n19025), .C2(n18989), .A(n13924), .B(n13923), .ZN(
        P2_U2843) );
  AOI22_X1 U17274 ( .A1(n20050), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20049), .ZN(n13926) );
  INV_X1 U17275 ( .A(n20078), .ZN(n13925) );
  NAND2_X1 U17276 ( .A1(n20037), .A2(n13925), .ZN(n13941) );
  NAND2_X1 U17277 ( .A1(n13926), .A2(n13941), .ZN(P1_U2953) );
  AOI22_X1 U17278 ( .A1(n20050), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20049), .ZN(n13928) );
  INV_X1 U17279 ( .A(n20069), .ZN(n13927) );
  NAND2_X1 U17280 ( .A1(n20037), .A2(n13927), .ZN(n13937) );
  NAND2_X1 U17281 ( .A1(n13928), .A2(n13937), .ZN(P1_U2937) );
  AOI22_X1 U17282 ( .A1(n20050), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20049), .ZN(n13930) );
  NAND2_X1 U17283 ( .A1(n13930), .A2(n13929), .ZN(P1_U2942) );
  AOI22_X1 U17284 ( .A1(n20050), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20049), .ZN(n13932) );
  NAND2_X1 U17285 ( .A1(n13932), .A2(n13931), .ZN(P1_U2944) );
  AOI22_X1 U17286 ( .A1(n20050), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20049), .ZN(n13934) );
  INV_X1 U17287 ( .A(n20090), .ZN(n13933) );
  NAND2_X1 U17288 ( .A1(n20037), .A2(n13933), .ZN(n13951) );
  NAND2_X1 U17289 ( .A1(n13934), .A2(n13951), .ZN(P1_U2941) );
  AOI22_X1 U17290 ( .A1(n20050), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20049), .ZN(n13936) );
  NAND2_X1 U17291 ( .A1(n13936), .A2(n13935), .ZN(P1_U2948) );
  AOI22_X1 U17292 ( .A1(n20050), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20049), .ZN(n13938) );
  NAND2_X1 U17293 ( .A1(n13938), .A2(n13937), .ZN(P1_U2952) );
  AOI22_X1 U17294 ( .A1(n20050), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20049), .ZN(n13940) );
  NAND2_X1 U17295 ( .A1(n13940), .A2(n13939), .ZN(P1_U2943) );
  AOI22_X1 U17296 ( .A1(n20050), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20049), .ZN(n13942) );
  NAND2_X1 U17297 ( .A1(n13942), .A2(n13941), .ZN(P1_U2938) );
  AOI22_X1 U17298 ( .A1(n20050), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20049), .ZN(n13944) );
  INV_X1 U17299 ( .A(n20082), .ZN(n13943) );
  NAND2_X1 U17300 ( .A1(n20037), .A2(n13943), .ZN(n13945) );
  NAND2_X1 U17301 ( .A1(n13944), .A2(n13945), .ZN(P1_U2939) );
  AOI22_X1 U17302 ( .A1(n20050), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20049), .ZN(n13946) );
  NAND2_X1 U17303 ( .A1(n13946), .A2(n13945), .ZN(P1_U2954) );
  AOI22_X1 U17304 ( .A1(n20050), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20049), .ZN(n13948) );
  INV_X1 U17305 ( .A(n20086), .ZN(n13947) );
  NAND2_X1 U17306 ( .A1(n20037), .A2(n13947), .ZN(n13949) );
  NAND2_X1 U17307 ( .A1(n13948), .A2(n13949), .ZN(P1_U2940) );
  AOI22_X1 U17308 ( .A1(n20050), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20049), .ZN(n13950) );
  NAND2_X1 U17309 ( .A1(n13950), .A2(n13949), .ZN(P1_U2955) );
  AOI22_X1 U17310 ( .A1(n20050), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20049), .ZN(n13952) );
  NAND2_X1 U17311 ( .A1(n13952), .A2(n13951), .ZN(P1_U2956) );
  OAI211_X1 U17312 ( .C1(n9686), .C2(n13955), .A(n15342), .B(n13954), .ZN(
        n13961) );
  INV_X1 U17313 ( .A(n13956), .ZN(n13957) );
  AOI21_X1 U17314 ( .B1(n13959), .B2(n13958), .A(n13957), .ZN(n16270) );
  NAND2_X1 U17315 ( .A1(n16270), .A2(n15316), .ZN(n13960) );
  OAI211_X1 U17316 ( .C1(n15316), .C2(n14249), .A(n13961), .B(n13960), .ZN(
        P2_U2872) );
  AOI22_X1 U17317 ( .A1(n9951), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n13962), .B2(n9949), .ZN(n14052) );
  INV_X1 U17318 ( .A(n13963), .ZN(n18998) );
  INV_X1 U17319 ( .A(n15801), .ZN(n13967) );
  NAND2_X1 U17320 ( .A1(n13964), .A2(n11249), .ZN(n14129) );
  MUX2_X1 U17321 ( .A(n11048), .B(n14129), .S(n13965), .Z(n13966) );
  AOI21_X1 U17322 ( .B1(n18998), .B2(n13967), .A(n13966), .ZN(n16315) );
  OAI22_X1 U17323 ( .A1(n16315), .A2(n15857), .B1(n13968), .B2(n16359), .ZN(
        n13969) );
  AOI21_X1 U17324 ( .B1(n14052), .B2(P2_STATE2_REG_1__SCAN_IN), .A(n13969), 
        .ZN(n13979) );
  NAND2_X1 U17325 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14270), .ZN(n16375) );
  INV_X1 U17326 ( .A(n16375), .ZN(n15958) );
  NOR2_X1 U17327 ( .A1(n10966), .A2(n13970), .ZN(n13971) );
  NAND2_X1 U17328 ( .A1(n13972), .A2(n13971), .ZN(n13976) );
  AND4_X1 U17329 ( .A1(n13976), .A2(n13975), .A3(n13974), .A4(n13973), .ZN(
        n16333) );
  OAI22_X1 U17330 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19839), .B1(n16333), 
        .B2(n18863), .ZN(n13977) );
  AOI21_X1 U17331 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n15958), .A(n13977), .ZN(
        n15818) );
  NAND2_X1 U17332 ( .A1(n15818), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13978) );
  OAI21_X1 U17333 ( .B1(n13979), .B2(n15818), .A(n13978), .ZN(P2_U3601) );
  NAND2_X1 U17334 ( .A1(n9949), .A2(n13980), .ZN(n13981) );
  XNOR2_X1 U17335 ( .A(n13982), .B(n13981), .ZN(n13983) );
  NAND2_X1 U17336 ( .A1(n13983), .A2(n18984), .ZN(n13992) );
  INV_X1 U17337 ( .A(n14119), .ZN(n19801) );
  NOR2_X1 U17338 ( .A1(n18974), .A2(n13984), .ZN(n13987) );
  INV_X1 U17339 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13985) );
  OAI22_X1 U17340 ( .A1(n15201), .A2(n13985), .B1(n13817), .B2(n18987), .ZN(
        n13986) );
  AOI211_X1 U17341 ( .C1(n13236), .C2(n13988), .A(n13987), .B(n13986), .ZN(
        n13989) );
  OAI21_X1 U17342 ( .B1(n13541), .B2(n18978), .A(n13989), .ZN(n13990) );
  AOI21_X1 U17343 ( .B1(n18954), .B2(n19801), .A(n13990), .ZN(n13991) );
  OAI211_X1 U17344 ( .C1(n19795), .C2(n18985), .A(n13992), .B(n13991), .ZN(
        P2_U2852) );
  NAND2_X1 U17345 ( .A1(n9949), .A2(n13993), .ZN(n13994) );
  XNOR2_X1 U17346 ( .A(n16254), .B(n13994), .ZN(n13995) );
  NAND2_X1 U17347 ( .A1(n13995), .A2(n18984), .ZN(n14003) );
  XNOR2_X1 U17348 ( .A(n13997), .B(n13996), .ZN(n19047) );
  AOI22_X1 U17349 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19000), .B1(
        P2_REIP_REG_5__SCAN_IN), .B2(n18951), .ZN(n13998) );
  OAI211_X1 U17350 ( .C1(n18989), .C2(n19047), .A(n13998), .B(n15534), .ZN(
        n14001) );
  NOR2_X1 U17351 ( .A1(n18995), .A2(n13999), .ZN(n14000) );
  AOI211_X1 U17352 ( .C1(P2_EBX_REG_5__SCAN_IN), .C2(n18992), .A(n14001), .B(
        n14000), .ZN(n14002) );
  OAI211_X1 U17353 ( .C1(n14204), .C2(n18978), .A(n14003), .B(n14002), .ZN(
        P2_U2850) );
  OAI222_X1 U17354 ( .A1(n14869), .A2(n19924), .B1(n14867), .B2(n12050), .C1(
        n14866), .C2(n20095), .ZN(P1_U2899) );
  INV_X1 U17355 ( .A(n19993), .ZN(n14008) );
  INV_X1 U17356 ( .A(n14004), .ZN(n19936) );
  AOI21_X1 U17357 ( .B1(n16060), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n14005), .ZN(n14006) );
  OAI21_X1 U17358 ( .B1(n16069), .B2(n19936), .A(n14006), .ZN(n14007) );
  AOI21_X1 U17359 ( .B1(n14008), .B2(n16066), .A(n14007), .ZN(n14009) );
  OAI21_X1 U17360 ( .B1(n19869), .B2(n14010), .A(n14009), .ZN(P1_U2995) );
  NOR2_X1 U17361 ( .A1(n9951), .A2(n14011), .ZN(n14049) );
  XNOR2_X1 U17362 ( .A(n14049), .B(n14012), .ZN(n14013) );
  NAND2_X1 U17363 ( .A1(n14013), .A2(n18984), .ZN(n14021) );
  OAI22_X1 U17364 ( .A1(n15201), .A2(n14014), .B1(n13397), .B2(n18987), .ZN(
        n14015) );
  AOI21_X1 U17365 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19000), .A(
        n14015), .ZN(n14016) );
  OAI21_X1 U17366 ( .B1(n18995), .B2(n14017), .A(n14016), .ZN(n14019) );
  NOR2_X1 U17367 ( .A1(n19806), .A2(n18989), .ZN(n14018) );
  AOI211_X1 U17368 ( .C1(n18999), .C2(n12860), .A(n14019), .B(n14018), .ZN(
        n14020) );
  OAI211_X1 U17369 ( .C1(n19804), .C2(n18985), .A(n14021), .B(n14020), .ZN(
        P2_U2853) );
  INV_X1 U17370 ( .A(n19924), .ZN(n14025) );
  AOI21_X1 U17371 ( .B1(n16060), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n14022), .ZN(n14023) );
  OAI21_X1 U17372 ( .B1(n16069), .B2(n19929), .A(n14023), .ZN(n14024) );
  AOI21_X1 U17373 ( .B1(n14025), .B2(n16066), .A(n14024), .ZN(n14026) );
  OAI21_X1 U17374 ( .B1(n19869), .B2(n14027), .A(n14026), .ZN(P1_U2994) );
  AOI22_X1 U17375 ( .A1(n16060), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n16118), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n14029) );
  NAND2_X1 U17376 ( .A1(n16055), .A2(n12008), .ZN(n14028) );
  OAI211_X1 U17377 ( .C1(n19977), .C2(n20055), .A(n14029), .B(n14028), .ZN(
        n14030) );
  AOI21_X1 U17378 ( .B1(n16065), .B2(n14031), .A(n14030), .ZN(n14032) );
  INV_X1 U17379 ( .A(n14032), .ZN(P1_U2998) );
  INV_X1 U17380 ( .A(n14033), .ZN(n14047) );
  NAND2_X1 U17381 ( .A1(n9949), .A2(n14034), .ZN(n14035) );
  XNOR2_X1 U17382 ( .A(n16178), .B(n14035), .ZN(n14036) );
  NAND2_X1 U17383 ( .A1(n14036), .A2(n18984), .ZN(n14046) );
  OR2_X1 U17384 ( .A1(n14038), .A2(n14037), .ZN(n14040) );
  NAND2_X1 U17385 ( .A1(n14040), .A2(n14039), .ZN(n19022) );
  AOI22_X1 U17386 ( .A1(P2_EBX_REG_13__SCAN_IN), .A2(n18992), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19000), .ZN(n14041) );
  OAI211_X1 U17387 ( .C1(n18989), .C2(n19022), .A(n14041), .B(n15534), .ZN(
        n14044) );
  NOR2_X1 U17388 ( .A1(n18987), .A2(n14042), .ZN(n14043) );
  AOI211_X1 U17389 ( .C1(n16186), .C2(n18999), .A(n14044), .B(n14043), .ZN(
        n14045) );
  OAI211_X1 U17390 ( .C1(n18995), .C2(n14047), .A(n14046), .B(n14045), .ZN(
        P2_U2842) );
  INV_X1 U17391 ( .A(n14048), .ZN(n14050) );
  OAI21_X1 U17392 ( .B1(n19003), .B2(n14050), .A(n14049), .ZN(n14179) );
  OAI21_X1 U17393 ( .B1(n9949), .B2(n14051), .A(n14179), .ZN(n14127) );
  NOR2_X1 U17394 ( .A1(n14052), .A2(n10302), .ZN(n14125) );
  NOR2_X1 U17395 ( .A1(n16334), .A2(n16339), .ZN(n15810) );
  INV_X1 U17396 ( .A(n15810), .ZN(n14059) );
  NOR2_X1 U17397 ( .A1(n14053), .A2(n16322), .ZN(n15809) );
  INV_X1 U17398 ( .A(n15809), .ZN(n15804) );
  NAND2_X1 U17399 ( .A1(n15804), .A2(n15802), .ZN(n14058) );
  OR2_X1 U17400 ( .A1(n11049), .A2(n11032), .ZN(n15803) );
  INV_X1 U17401 ( .A(n15803), .ZN(n14056) );
  INV_X1 U17402 ( .A(n14054), .ZN(n15807) );
  NAND2_X1 U17403 ( .A1(n11048), .A2(n15807), .ZN(n15805) );
  NOR2_X1 U17404 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n16322), .ZN(
        n14055) );
  OAI22_X1 U17405 ( .A1(n14056), .A2(n14058), .B1(n15805), .B2(n14055), .ZN(
        n14057) );
  AOI21_X1 U17406 ( .B1(n14059), .B2(n14058), .A(n14057), .ZN(n14060) );
  OAI21_X1 U17407 ( .B1(n19139), .B2(n15801), .A(n14060), .ZN(n16321) );
  INV_X1 U17408 ( .A(n16321), .ZN(n14061) );
  OAI22_X1 U17409 ( .A1(n19804), .A2(n16359), .B1(n15857), .B2(n14061), .ZN(
        n14062) );
  AOI21_X1 U17410 ( .B1(n14127), .B2(n14125), .A(n14062), .ZN(n14064) );
  NAND2_X1 U17411 ( .A1(n15818), .A2(n16322), .ZN(n14063) );
  OAI21_X1 U17412 ( .B1(n14064), .B2(n15818), .A(n14063), .ZN(P2_U3599) );
  NAND2_X1 U17413 ( .A1(n13841), .A2(n14066), .ZN(n14067) );
  NAND2_X1 U17414 ( .A1(n14166), .A2(n14067), .ZN(n19986) );
  OAI222_X1 U17415 ( .A1(n19986), .A2(n14869), .B1(n14068), .B2(n14867), .C1(
        n14866), .C2(n20099), .ZN(P1_U2898) );
  AOI21_X1 U17416 ( .B1(n14069), .B2(n13954), .A(n9677), .ZN(n19013) );
  NAND2_X1 U17417 ( .A1(n19013), .A2(n15342), .ZN(n14073) );
  NAND2_X1 U17418 ( .A1(n13956), .A2(n14070), .ZN(n14071) );
  AND2_X1 U17419 ( .A1(n14136), .A2(n14071), .ZN(n18939) );
  NAND2_X1 U17420 ( .A1(n15316), .A2(n18939), .ZN(n14072) );
  OAI211_X1 U17421 ( .C1(n15316), .C2(n14074), .A(n14073), .B(n14072), .ZN(
        P2_U2871) );
  NAND2_X1 U17422 ( .A1(n14076), .A2(n14075), .ZN(n14077) );
  XNOR2_X1 U17423 ( .A(n14077), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19119) );
  INV_X1 U17424 ( .A(n19119), .ZN(n14086) );
  XOR2_X1 U17425 ( .A(n14079), .B(n14078), .Z(n19120) );
  NOR2_X1 U17426 ( .A1(n14197), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14084) );
  NOR2_X1 U17427 ( .A1(n11084), .A2(n15534), .ZN(n14080) );
  AOI21_X1 U17428 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n14203), .A(
        n14080), .ZN(n14082) );
  NAND2_X1 U17429 ( .A1(n16298), .A2(n14121), .ZN(n14081) );
  OAI211_X1 U17430 ( .C1(n19115), .C2(n19138), .A(n14082), .B(n14081), .ZN(
        n14083) );
  AOI211_X1 U17431 ( .C1(n19120), .C2(n16300), .A(n14084), .B(n14083), .ZN(
        n14085) );
  OAI21_X1 U17432 ( .B1(n19137), .B2(n14086), .A(n14085), .ZN(P2_U3042) );
  NAND2_X1 U17433 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20748), .ZN(n15935) );
  AND2_X1 U17434 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20744), .ZN(n14087) );
  NAND2_X1 U17435 ( .A1(n12499), .A2(n14087), .ZN(n14088) );
  OAI211_X1 U17436 ( .C1(n15935), .C2(n20744), .A(n16134), .B(n14088), .ZN(
        n14089) );
  INV_X1 U17437 ( .A(n14089), .ZN(n14090) );
  NOR2_X1 U17438 ( .A1(n14112), .A2(n14091), .ZN(n19980) );
  NAND2_X1 U17439 ( .A1(n20647), .A2(n20742), .ZN(n14103) );
  INV_X1 U17440 ( .A(n14103), .ZN(n14093) );
  INV_X1 U17441 ( .A(n19972), .ZN(n19948) );
  NAND2_X1 U17442 ( .A1(n19888), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n14110) );
  AND2_X1 U17443 ( .A1(n20076), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n14104) );
  OR2_X1 U17444 ( .A1(n15925), .A2(n14104), .ZN(n14096) );
  INV_X1 U17445 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14098) );
  INV_X1 U17446 ( .A(n14492), .ZN(n14100) );
  AOI21_X1 U17447 ( .B1(n19975), .B2(n19983), .A(n14101), .ZN(n14102) );
  AOI21_X1 U17448 ( .B1(n9585), .B2(P1_EBX_REG_0__SCAN_IN), .A(n14102), .ZN(
        n14109) );
  NAND2_X1 U17449 ( .A1(n14104), .A2(n14103), .ZN(n14105) );
  NAND2_X1 U17450 ( .A1(n19971), .A2(n14107), .ZN(n14108) );
  NAND3_X1 U17451 ( .A1(n14110), .A2(n14109), .A3(n14108), .ZN(n14116) );
  OR2_X1 U17452 ( .A1(n14112), .A2(n14111), .ZN(n14113) );
  NOR2_X1 U17453 ( .A1(n14114), .A2(n19976), .ZN(n14115) );
  AOI211_X1 U17454 ( .C1(n19980), .C2(n9594), .A(n14116), .B(n14115), .ZN(
        n14117) );
  INV_X1 U17455 ( .A(n14117), .ZN(P1_U2840) );
  AOI21_X1 U17456 ( .B1(n19806), .B2(n19804), .A(n14118), .ZN(n19051) );
  XNOR2_X1 U17457 ( .A(n19795), .B(n14119), .ZN(n19050) );
  NOR2_X1 U17458 ( .A1(n19051), .A2(n19050), .ZN(n19049) );
  AOI21_X1 U17459 ( .B1(n19795), .B2(n14119), .A(n19049), .ZN(n14120) );
  NOR2_X1 U17460 ( .A1(n14120), .A2(n14121), .ZN(n19044) );
  XNOR2_X1 U17461 ( .A(n19044), .B(n19043), .ZN(n14124) );
  AOI22_X1 U17462 ( .A1(n19056), .A2(n14121), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19055), .ZN(n14123) );
  NAND2_X1 U17463 ( .A1(n19033), .A2(n16163), .ZN(n14122) );
  OAI211_X1 U17464 ( .C1(n14124), .C2(n19060), .A(n14123), .B(n14122), .ZN(
        P2_U2915) );
  INV_X1 U17465 ( .A(n15818), .ZN(n15861) );
  INV_X1 U17466 ( .A(n14125), .ZN(n14126) );
  NOR2_X1 U17467 ( .A1(n14127), .A2(n14126), .ZN(n14133) );
  NOR2_X1 U17468 ( .A1(n14128), .A2(n14053), .ZN(n14130) );
  AOI22_X1 U17469 ( .A1(n11048), .A2(n14135), .B1(n14130), .B2(n14129), .ZN(
        n14131) );
  OAI21_X1 U17470 ( .B1(n15792), .B2(n15801), .A(n14131), .ZN(n16316) );
  INV_X1 U17471 ( .A(n16316), .ZN(n16317) );
  OAI22_X1 U17472 ( .A1(n19816), .A2(n16359), .B1(n15857), .B2(n16317), .ZN(
        n14132) );
  OAI21_X1 U17473 ( .B1(n14133), .B2(n14132), .A(n15861), .ZN(n14134) );
  OAI21_X1 U17474 ( .B1(n15861), .B2(n14135), .A(n14134), .ZN(P2_U3600) );
  OAI21_X1 U17475 ( .B1(n9677), .B2(n9699), .A(n9626), .ZN(n14262) );
  NAND2_X1 U17476 ( .A1(n15347), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n14139) );
  AOI21_X1 U17477 ( .B1(n14137), .B2(n14136), .A(n14174), .ZN(n18929) );
  NAND2_X1 U17478 ( .A1(n18929), .A2(n15316), .ZN(n14138) );
  OAI211_X1 U17479 ( .C1(n14262), .C2(n15350), .A(n14139), .B(n14138), .ZN(
        P2_U2870) );
  XNOR2_X1 U17480 ( .A(n14141), .B(n14140), .ZN(n16138) );
  INV_X1 U17481 ( .A(n19986), .ZN(n14144) );
  AOI22_X1 U17482 ( .A1(n16060), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n16118), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n14142) );
  OAI21_X1 U17483 ( .B1(n16069), .B2(n19916), .A(n14142), .ZN(n14143) );
  AOI21_X1 U17484 ( .B1(n14144), .B2(n16066), .A(n14143), .ZN(n14145) );
  OAI21_X1 U17485 ( .B1(n19869), .B2(n16138), .A(n14145), .ZN(P1_U2993) );
  XOR2_X1 U17486 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n14147), .Z(
        n14148) );
  XNOR2_X1 U17487 ( .A(n14149), .B(n14148), .ZN(n14311) );
  AOI21_X1 U17488 ( .B1(n16099), .B2(n14151), .A(n14150), .ZN(n16144) );
  OAI21_X1 U17489 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16071), .A(
        n16144), .ZN(n16121) );
  NAND2_X1 U17490 ( .A1(n14153), .A2(n14152), .ZN(n16127) );
  AOI211_X1 U17491 ( .C1(n14155), .C2(n14154), .A(n16142), .B(n16127), .ZN(
        n14157) );
  NAND2_X1 U17492 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n14156) );
  AOI22_X1 U17493 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n16121), .B1(
        n14157), .B2(n14156), .ZN(n14162) );
  AOI21_X1 U17494 ( .B1(n16132), .B2(n14167), .A(n14158), .ZN(n14159) );
  OR2_X1 U17495 ( .A1(n14215), .A2(n14159), .ZN(n14263) );
  INV_X1 U17496 ( .A(n14263), .ZN(n14229) );
  INV_X1 U17497 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n14160) );
  NOR2_X1 U17498 ( .A1(n16134), .A2(n14160), .ZN(n14307) );
  AOI21_X1 U17499 ( .B1(n14229), .B2(n16119), .A(n14307), .ZN(n14161) );
  OAI211_X1 U17500 ( .C1(n14311), .C2(n16137), .A(n14162), .B(n14161), .ZN(
        P1_U3023) );
  INV_X1 U17501 ( .A(n14164), .ZN(n14165) );
  AOI21_X1 U17502 ( .B1(n14163), .B2(n14166), .A(n14165), .ZN(n19900) );
  INV_X1 U17503 ( .A(n19900), .ZN(n14169) );
  INV_X1 U17504 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n14168) );
  XNOR2_X1 U17505 ( .A(n16132), .B(n14167), .ZN(n19896) );
  OAI222_X1 U17506 ( .A1(n19992), .A2(n14169), .B1(n14168), .B2(n19997), .C1(
        n19985), .C2(n19896), .ZN(P1_U2865) );
  OAI222_X1 U17507 ( .A1(n14869), .A2(n14169), .B1(n14867), .B2(n12062), .C1(
        n14866), .C2(n20107), .ZN(P1_U2897) );
  INV_X1 U17508 ( .A(n14170), .ZN(n14171) );
  AOI21_X1 U17509 ( .B1(n14171), .B2(n9626), .A(n9676), .ZN(n16169) );
  NAND2_X1 U17510 ( .A1(n16169), .A2(n15342), .ZN(n14177) );
  OR2_X1 U17511 ( .A1(n14174), .A2(n14173), .ZN(n14175) );
  AND2_X1 U17512 ( .A1(n14172), .A2(n14175), .ZN(n18917) );
  NAND2_X1 U17513 ( .A1(n18917), .A2(n15316), .ZN(n14176) );
  OAI211_X1 U17514 ( .C1(n15316), .C2(n14178), .A(n14177), .B(n14176), .ZN(
        P2_U2869) );
  AOI221_X1 U17515 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n14179), .C1(
        n9949), .C2(n14179), .A(n19717), .ZN(n14180) );
  INV_X1 U17516 ( .A(n14180), .ZN(n14188) );
  INV_X1 U17517 ( .A(n14181), .ZN(n14184) );
  AOI22_X1 U17518 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19000), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n18951), .ZN(n14183) );
  NAND2_X1 U17519 ( .A1(n18992), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n14182) );
  OAI211_X1 U17520 ( .C1(n18995), .C2(n14184), .A(n14183), .B(n14182), .ZN(
        n14186) );
  NOR2_X1 U17521 ( .A1(n15792), .A2(n18978), .ZN(n14185) );
  AOI211_X1 U17522 ( .C1(n18954), .C2(n19820), .A(n14186), .B(n14185), .ZN(
        n14187) );
  OAI211_X1 U17523 ( .C1(n19816), .C2(n18985), .A(n14188), .B(n14187), .ZN(
        P2_U2854) );
  XNOR2_X1 U17524 ( .A(n14190), .B(n14189), .ZN(n16259) );
  AND2_X1 U17525 ( .A1(n14192), .A2(n14191), .ZN(n14193) );
  OAI22_X1 U17526 ( .A1(n14196), .A2(n14195), .B1(n14194), .B2(n14193), .ZN(
        n16257) );
  NOR2_X1 U17527 ( .A1(n11089), .A2(n15534), .ZN(n14202) );
  AOI211_X1 U17528 ( .C1(n14200), .C2(n14199), .A(n14198), .B(n14197), .ZN(
        n14201) );
  AOI211_X1 U17529 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n14203), .A(
        n14202), .B(n14201), .ZN(n14207) );
  INV_X1 U17530 ( .A(n14204), .ZN(n16261) );
  INV_X1 U17531 ( .A(n19047), .ZN(n14205) );
  AOI22_X1 U17532 ( .A1(n16261), .A2(n16302), .B1(n16298), .B2(n14205), .ZN(
        n14206) );
  OAI211_X1 U17533 ( .C1(n16257), .C2(n19137), .A(n14207), .B(n14206), .ZN(
        n14208) );
  INV_X1 U17534 ( .A(n14208), .ZN(n14209) );
  OAI21_X1 U17535 ( .B1(n19133), .B2(n16259), .A(n14209), .ZN(P2_U3041) );
  MUX2_X1 U17536 ( .A(n11751), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .S(
        n15131), .Z(n14210) );
  XNOR2_X1 U17537 ( .A(n14211), .B(n14210), .ZN(n14377) );
  NAND2_X1 U17538 ( .A1(n14213), .A2(n14212), .ZN(n14218) );
  NOR2_X1 U17539 ( .A1(n15145), .A2(n14218), .ZN(n15161) );
  OR2_X1 U17540 ( .A1(n14215), .A2(n14214), .ZN(n14216) );
  NAND2_X1 U17541 ( .A1(n14335), .A2(n14216), .ZN(n14368) );
  INV_X1 U17542 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n16001) );
  OAI22_X1 U17543 ( .A1(n14368), .A2(n16136), .B1(n16001), .B2(n16134), .ZN(
        n14217) );
  AOI21_X1 U17544 ( .B1(n15161), .B2(n11751), .A(n14217), .ZN(n14223) );
  INV_X1 U17545 ( .A(n14218), .ZN(n14221) );
  AOI21_X1 U17546 ( .B1(n14221), .B2(n14220), .A(n14219), .ZN(n15162) );
  NAND2_X1 U17547 ( .A1(n15162), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14222) );
  OAI211_X1 U17548 ( .C1(n14377), .C2(n16137), .A(n14223), .B(n14222), .ZN(
        P1_U3022) );
  AND2_X1 U17549 ( .A1(n14164), .A2(n14224), .ZN(n14226) );
  OR2_X1 U17550 ( .A1(n14226), .A2(n14225), .ZN(n14303) );
  INV_X1 U17551 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n14305) );
  OAI22_X1 U17552 ( .A1(n14305), .A2(n19975), .B1(n19983), .B2(n14227), .ZN(
        n14232) );
  INV_X1 U17553 ( .A(n14228), .ZN(n14563) );
  INV_X1 U17554 ( .A(n19918), .ZN(n19931) );
  NAND4_X1 U17555 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n14497)
         );
  INV_X1 U17556 ( .A(n19888), .ZN(n14676) );
  NAND4_X1 U17557 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n14498)
         );
  NOR2_X1 U17558 ( .A1(n19972), .A2(n14498), .ZN(n19887) );
  NOR2_X1 U17559 ( .A1(n14676), .A2(n19887), .ZN(n19935) );
  AOI21_X1 U17560 ( .B1(n14497), .B2(n19888), .A(n19935), .ZN(n14748) );
  AOI22_X1 U17561 ( .A1(n19971), .A2(n14229), .B1(n9585), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n14230) );
  OAI21_X1 U17562 ( .B1(n14748), .B2(n14160), .A(n14230), .ZN(n14231) );
  NOR3_X1 U17563 ( .A1(n14232), .A2(n19931), .A3(n14231), .ZN(n14236) );
  NAND3_X1 U17564 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n14234) );
  NAND3_X1 U17565 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n14233) );
  NOR2_X1 U17566 ( .A1(n19942), .A2(n14233), .ZN(n19930) );
  NAND2_X1 U17567 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n19930), .ZN(n19917) );
  NOR2_X1 U17568 ( .A1(n14234), .A2(n19917), .ZN(n14363) );
  NAND2_X1 U17569 ( .A1(n14363), .A2(n14160), .ZN(n14235) );
  OAI211_X1 U17570 ( .C1(n14303), .C2(n19903), .A(n14236), .B(n14235), .ZN(
        P1_U2832) );
  NAND2_X1 U17571 ( .A1(n9949), .A2(n14237), .ZN(n14238) );
  XNOR2_X1 U17572 ( .A(n15566), .B(n14238), .ZN(n14239) );
  NAND2_X1 U17573 ( .A1(n14239), .A2(n18984), .ZN(n14252) );
  OR2_X1 U17574 ( .A1(n14241), .A2(n14240), .ZN(n14243) );
  NAND2_X1 U17575 ( .A1(n14243), .A2(n14242), .ZN(n19018) );
  INV_X1 U17576 ( .A(n19018), .ZN(n14247) );
  OAI21_X1 U17577 ( .B1(n11227), .B2(n18987), .A(n15534), .ZN(n14246) );
  NOR2_X1 U17578 ( .A1(n18974), .A2(n14244), .ZN(n14245) );
  AOI211_X1 U17579 ( .C1(n18954), .C2(n14247), .A(n14246), .B(n14245), .ZN(
        n14248) );
  OAI21_X1 U17580 ( .B1(n15201), .B2(n14249), .A(n14248), .ZN(n14250) );
  AOI21_X1 U17581 ( .B1(n18999), .B2(n16270), .A(n14250), .ZN(n14251) );
  OAI211_X1 U17582 ( .C1(n18995), .C2(n14253), .A(n14252), .B(n14251), .ZN(
        P2_U2840) );
  OAI22_X1 U17583 ( .A1(n15410), .A2(n19065), .B1(n19041), .B2(n14254), .ZN(
        n14259) );
  NAND2_X1 U17584 ( .A1(n15718), .A2(n14256), .ZN(n14257) );
  NAND2_X1 U17585 ( .A1(n15685), .A2(n14257), .ZN(n18927) );
  NOR2_X1 U17586 ( .A1(n15385), .A2(n18927), .ZN(n14258) );
  NOR2_X1 U17587 ( .A1(n14259), .A2(n14258), .ZN(n14261) );
  AOI22_X1 U17588 ( .A1(n19011), .A2(BUF2_REG_17__SCAN_IN), .B1(n19010), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n14260) );
  OAI211_X1 U17589 ( .C1(n14262), .C2(n19060), .A(n14261), .B(n14260), .ZN(
        P2_U2902) );
  INV_X1 U17590 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14264) );
  OAI222_X1 U17591 ( .A1(n14303), .A2(n19992), .B1(n14264), .B2(n19997), .C1(
        n14263), .C2(n19985), .ZN(P1_U2864) );
  INV_X1 U17592 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n14266) );
  INV_X1 U17593 ( .A(DATAI_8_), .ZN(n14265) );
  MUX2_X1 U17594 ( .A(n14265), .B(n16481), .S(n20053), .Z(n20020) );
  OAI222_X1 U17595 ( .A1(n14303), .A2(n14869), .B1(n14266), .B2(n14867), .C1(
        n14866), .C2(n20020), .ZN(P1_U2896) );
  NOR2_X2 U17596 ( .A1(n19420), .A2(n19327), .ZN(n19200) );
  OAI21_X1 U17597 ( .B1(n19708), .B2(n19200), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n14267) );
  NAND2_X1 U17598 ( .A1(n14267), .A2(n19793), .ZN(n14282) );
  INV_X1 U17599 ( .A(n14282), .ZN(n14275) );
  INV_X1 U17600 ( .A(n14268), .ZN(n14269) );
  AND2_X1 U17601 ( .A1(n14269), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19703) );
  NAND2_X1 U17602 ( .A1(n19803), .A2(n19813), .ZN(n19233) );
  INV_X1 U17603 ( .A(n19233), .ZN(n19234) );
  NAND2_X1 U17604 ( .A1(n19234), .A2(n19822), .ZN(n19178) );
  NOR2_X1 U17605 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19178), .ZN(
        n19168) );
  NOR2_X1 U17606 ( .A1(n19703), .A2(n19168), .ZN(n14281) );
  AOI211_X1 U17607 ( .C1(n10482), .C2(n19839), .A(n19168), .B(n19793), .ZN(
        n14274) );
  NOR2_X1 U17608 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19850) );
  INV_X1 U17609 ( .A(n19850), .ZN(n14272) );
  INV_X1 U17610 ( .A(n14270), .ZN(n14271) );
  NAND2_X1 U17611 ( .A1(n14272), .A2(n14271), .ZN(n14273) );
  INV_X1 U17612 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14287) );
  AOI22_X1 U17613 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19171), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19170), .ZN(n19668) );
  INV_X1 U17614 ( .A(n19668), .ZN(n19613) );
  AOI22_X1 U17615 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19171), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19170), .ZN(n19625) );
  INV_X1 U17616 ( .A(n19200), .ZN(n14297) );
  INV_X1 U17617 ( .A(n19168), .ZN(n14296) );
  NAND2_X1 U17618 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19662), .ZN(n19166) );
  NAND2_X1 U17619 ( .A1(n10274), .A2(n19149), .ZN(n19489) );
  OAI22_X1 U17620 ( .A1(n19625), .A2(n14297), .B1(n14296), .B2(n19489), .ZN(
        n14279) );
  AOI21_X1 U17621 ( .B1(n19708), .B2(n19613), .A(n14279), .ZN(n14286) );
  OAI21_X1 U17622 ( .B1(n10482), .B2(n19168), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14280) );
  NAND2_X1 U17623 ( .A1(n19172), .A2(n14284), .ZN(n14285) );
  OAI211_X1 U17624 ( .C1(n19176), .C2(n14287), .A(n14286), .B(n14285), .ZN(
        P2_U3048) );
  AOI22_X1 U17625 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19170), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19171), .ZN(n19702) );
  INV_X1 U17626 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16459) );
  INV_X1 U17627 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n20902) );
  NAND2_X1 U17628 ( .A1(n10214), .A2(n19149), .ZN(n19526) );
  OAI22_X1 U17629 ( .A1(n19604), .A2(n14297), .B1(n14296), .B2(n19526), .ZN(
        n14288) );
  AOI21_X1 U17630 ( .B1(n19708), .B2(n19600), .A(n14288), .ZN(n14290) );
  NOR2_X2 U17631 ( .A1(n19038), .A2(n19363), .ZN(n19698) );
  NAND2_X1 U17632 ( .A1(n19172), .A2(n19698), .ZN(n14289) );
  OAI211_X1 U17633 ( .C1(n19176), .C2(n14291), .A(n14290), .B(n14289), .ZN(
        P2_U3054) );
  AOI22_X1 U17634 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19170), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19171), .ZN(n19696) );
  INV_X1 U17635 ( .A(n19696), .ZN(n19640) );
  INV_X1 U17636 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20843) );
  INV_X1 U17637 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n18212) );
  NAND2_X1 U17638 ( .A1(n10038), .A2(n19149), .ZN(n19521) );
  OAI22_X1 U17639 ( .A1(n19643), .A2(n14297), .B1(n14296), .B2(n19521), .ZN(
        n14292) );
  AOI21_X1 U17640 ( .B1(n19708), .B2(n19640), .A(n14292), .ZN(n14294) );
  NOR2_X2 U17641 ( .A1(n19040), .A2(n19363), .ZN(n19692) );
  NAND2_X1 U17642 ( .A1(n19172), .A2(n19692), .ZN(n14293) );
  OAI211_X1 U17643 ( .C1(n19176), .C2(n14295), .A(n14294), .B(n14293), .ZN(
        P2_U3053) );
  AOI22_X1 U17644 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19171), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19170), .ZN(n19673) );
  INV_X1 U17645 ( .A(n19673), .ZN(n19626) );
  AOI22_X1 U17646 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19171), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19170), .ZN(n19629) );
  NAND2_X1 U17647 ( .A1(n9600), .A2(n19149), .ZN(n19499) );
  OAI22_X1 U17648 ( .A1(n19629), .A2(n14297), .B1(n14296), .B2(n19499), .ZN(
        n14298) );
  AOI21_X1 U17649 ( .B1(n19708), .B2(n19626), .A(n14298), .ZN(n14301) );
  NAND2_X1 U17650 ( .A1(n19172), .A2(n14299), .ZN(n14300) );
  OAI211_X1 U17651 ( .C1(n19176), .C2(n14302), .A(n14301), .B(n14300), .ZN(
        P2_U3049) );
  INV_X1 U17652 ( .A(n14303), .ZN(n14304) );
  NAND2_X1 U17653 ( .A1(n14304), .A2(n16066), .ZN(n14310) );
  NOR2_X1 U17654 ( .A1(n14973), .A2(n14305), .ZN(n14306) );
  AOI211_X1 U17655 ( .C1(n16055), .C2(n14308), .A(n14307), .B(n14306), .ZN(
        n14309) );
  OAI211_X1 U17656 ( .C1(n14311), .C2(n19869), .A(n14310), .B(n14309), .ZN(
        P1_U2991) );
  OAI21_X1 U17657 ( .B1(n14313), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n14312), .ZN(n16248) );
  XOR2_X1 U17658 ( .A(n14315), .B(n14314), .Z(n16250) );
  NAND2_X1 U17659 ( .A1(n16250), .A2(n16300), .ZN(n14325) );
  INV_X1 U17660 ( .A(n14316), .ZN(n14323) );
  INV_X1 U17661 ( .A(n19039), .ZN(n14319) );
  NOR2_X1 U17662 ( .A1(n15534), .A2(n14317), .ZN(n14318) );
  AOI21_X1 U17663 ( .B1(n16298), .B2(n14319), .A(n14318), .ZN(n14320) );
  OAI21_X1 U17664 ( .B1(n16246), .B2(n19138), .A(n14320), .ZN(n14322) );
  AOI211_X1 U17665 ( .C1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n14323), .A(
        n14322), .B(n14321), .ZN(n14324) );
  OAI211_X1 U17666 ( .C1(n16248), .C2(n19137), .A(n14325), .B(n14324), .ZN(
        P2_U3040) );
  NOR2_X1 U17667 ( .A1(n14225), .A2(n14327), .ZN(n14328) );
  OR2_X1 U17668 ( .A1(n14326), .A2(n14328), .ZN(n14362) );
  INV_X1 U17669 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n14329) );
  OAI222_X1 U17670 ( .A1(n14362), .A2(n19992), .B1(n19997), .B2(n14329), .C1(
        n14368), .C2(n19985), .ZN(P1_U2863) );
  INV_X1 U17671 ( .A(DATAI_9_), .ZN(n14331) );
  MUX2_X1 U17672 ( .A(n14331), .B(n14330), .S(n20053), .Z(n20023) );
  OAI222_X1 U17673 ( .A1(n14362), .A2(n14869), .B1(n14332), .B2(n14867), .C1(
        n14866), .C2(n20023), .ZN(P1_U2895) );
  OAI21_X1 U17674 ( .B1(n14326), .B2(n14334), .A(n14333), .ZN(n15999) );
  INV_X1 U17675 ( .A(n14382), .ZN(n14741) );
  AOI21_X1 U17676 ( .B1(n14336), .B2(n14335), .A(n14741), .ZN(n16003) );
  AOI22_X1 U17677 ( .A1(n16003), .A2(n12508), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n12469), .ZN(n14337) );
  OAI21_X1 U17678 ( .B1(n15999), .B2(n19992), .A(n14337), .ZN(P1_U2862) );
  INV_X1 U17679 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14339) );
  INV_X1 U17680 ( .A(DATAI_10_), .ZN(n14338) );
  MUX2_X1 U17681 ( .A(n14338), .B(n16478), .S(n20053), .Z(n20027) );
  OAI222_X1 U17682 ( .A1(n15999), .A2(n14869), .B1(n14339), .B2(n14867), .C1(
        n14866), .C2(n20027), .ZN(P1_U2894) );
  NAND2_X1 U17683 ( .A1(n16233), .A2(n16232), .ZN(n14341) );
  XOR2_X1 U17684 ( .A(n14341), .B(n14340), .Z(n14361) );
  XNOR2_X1 U17685 ( .A(n14343), .B(n14342), .ZN(n14344) );
  XNOR2_X1 U17686 ( .A(n14345), .B(n14344), .ZN(n14359) );
  OAI22_X1 U17687 ( .A1(n16265), .A2(n18973), .B1(n10797), .B2(n15534), .ZN(
        n14346) );
  AOI21_X1 U17688 ( .B1(n16255), .B2(n18971), .A(n14346), .ZN(n14347) );
  OAI21_X1 U17689 ( .B1(n18979), .B2(n16247), .A(n14347), .ZN(n14348) );
  AOI21_X1 U17690 ( .B1(n14359), .B2(n19118), .A(n14348), .ZN(n14349) );
  OAI21_X1 U17691 ( .B1(n14361), .B2(n16258), .A(n14349), .ZN(P2_U3007) );
  INV_X1 U17692 ( .A(n16310), .ZN(n14357) );
  NOR2_X1 U17693 ( .A1(n18979), .A2(n19138), .ZN(n14355) );
  OR2_X1 U17694 ( .A1(n14351), .A2(n14350), .ZN(n14353) );
  NAND2_X1 U17695 ( .A1(n14353), .A2(n14352), .ZN(n19037) );
  OAI22_X1 U17696 ( .A1(n19143), .A2(n19037), .B1(n10797), .B2(n15534), .ZN(
        n14354) );
  AOI211_X1 U17697 ( .C1(n16299), .C2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n14355), .B(n14354), .ZN(n14356) );
  OAI21_X1 U17698 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n14357), .A(
        n14356), .ZN(n14358) );
  AOI21_X1 U17699 ( .B1(n14359), .B2(n16271), .A(n14358), .ZN(n14360) );
  OAI21_X1 U17700 ( .B1(n14361), .B2(n19133), .A(n14360), .ZN(P2_U3039) );
  INV_X1 U17701 ( .A(n14362), .ZN(n14375) );
  NAND2_X1 U17702 ( .A1(n14375), .A2(n19899), .ZN(n14371) );
  NAND2_X1 U17703 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14363), .ZN(n16000) );
  INV_X1 U17704 ( .A(n16000), .ZN(n14747) );
  OR2_X1 U17705 ( .A1(n19975), .A2(n14364), .ZN(n14365) );
  OAI211_X1 U17706 ( .C1(n14373), .C2(n19983), .A(n14365), .B(n19918), .ZN(
        n14366) );
  AOI21_X1 U17707 ( .B1(n9585), .B2(P1_EBX_REG_9__SCAN_IN), .A(n14366), .ZN(
        n14367) );
  OAI21_X1 U17708 ( .B1(n14368), .B2(n19968), .A(n14367), .ZN(n14369) );
  AOI21_X1 U17709 ( .B1(n14747), .B2(n16001), .A(n14369), .ZN(n14370) );
  OAI211_X1 U17710 ( .C1(n16001), .C2(n14748), .A(n14371), .B(n14370), .ZN(
        P1_U2831) );
  AOI22_X1 U17711 ( .A1(n16060), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n16118), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n14372) );
  OAI21_X1 U17712 ( .B1(n16069), .B2(n14373), .A(n14372), .ZN(n14374) );
  AOI21_X1 U17713 ( .B1(n14375), .B2(n16066), .A(n14374), .ZN(n14376) );
  OAI21_X1 U17714 ( .B1(n14377), .B2(n19869), .A(n14376), .ZN(P1_U2990) );
  OR2_X1 U17715 ( .A1(n14380), .A2(n14379), .ZN(n14381) );
  AND2_X1 U17716 ( .A1(n14378), .A2(n14381), .ZN(n15995) );
  INV_X1 U17717 ( .A(n15995), .ZN(n14385) );
  XNOR2_X1 U17718 ( .A(n14382), .B(n14740), .ZN(n16112) );
  AOI22_X1 U17719 ( .A1(n16112), .A2(n12508), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n12469), .ZN(n14383) );
  OAI21_X1 U17720 ( .B1(n14385), .B2(n19992), .A(n14383), .ZN(P1_U2861) );
  INV_X1 U17721 ( .A(n14806), .ZN(n14384) );
  OAI222_X1 U17722 ( .A1(n14385), .A2(n14869), .B1(n20005), .B2(n14867), .C1(
        n14866), .C2(n14384), .ZN(P1_U2893) );
  AOI22_X1 U17723 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n17143), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17127), .ZN(n14395) );
  AOI22_X1 U17724 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n15823), .ZN(n14394) );
  AOI22_X1 U17725 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n17109), .ZN(n14386) );
  OAI21_X1 U17726 ( .B1(n20813), .B2(n14457), .A(n14386), .ZN(n14392) );
  AOI22_X1 U17727 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17108), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n17125), .ZN(n14390) );
  AOI22_X1 U17728 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n12692), .B1(
        n12703), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14389) );
  AOI22_X1 U17729 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14388) );
  AOI22_X1 U17730 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n14458), .ZN(n14387) );
  NAND4_X1 U17731 ( .A1(n14390), .A2(n14389), .A3(n14388), .A4(n14387), .ZN(
        n14391) );
  AOI211_X1 U17732 ( .C1(n17116), .C2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n14392), .B(n14391), .ZN(n14393) );
  NAND3_X1 U17733 ( .A1(n14395), .A2(n14394), .A3(n14393), .ZN(n14480) );
  AOI22_X1 U17734 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14399) );
  AOI22_X1 U17735 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14398) );
  AOI22_X1 U17736 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14397) );
  AOI22_X1 U17737 ( .A1(n17108), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14396) );
  NAND4_X1 U17738 ( .A1(n14399), .A2(n14398), .A3(n14397), .A4(n14396), .ZN(
        n14405) );
  AOI22_X1 U17739 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14403) );
  AOI22_X1 U17740 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14402) );
  AOI22_X1 U17741 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14401) );
  AOI22_X1 U17742 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14400) );
  NAND4_X1 U17743 ( .A1(n14403), .A2(n14402), .A3(n14401), .A4(n14400), .ZN(
        n14404) );
  NOR2_X1 U17744 ( .A1(n14405), .A2(n14404), .ZN(n16930) );
  AOI22_X1 U17745 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14409) );
  AOI22_X1 U17746 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14408) );
  AOI22_X1 U17747 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14407) );
  AOI22_X1 U17748 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14406) );
  NAND4_X1 U17749 ( .A1(n14409), .A2(n14408), .A3(n14407), .A4(n14406), .ZN(
        n14415) );
  AOI22_X1 U17750 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14413) );
  AOI22_X1 U17751 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14412) );
  AOI22_X1 U17752 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12703), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14411) );
  AOI22_X1 U17753 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14410) );
  NAND4_X1 U17754 ( .A1(n14413), .A2(n14412), .A3(n14411), .A4(n14410), .ZN(
        n14414) );
  NOR2_X1 U17755 ( .A1(n14415), .A2(n14414), .ZN(n16929) );
  AOI22_X1 U17756 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12703), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14419) );
  AOI22_X1 U17757 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14418) );
  AOI22_X1 U17758 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17132), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14417) );
  AOI22_X1 U17759 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14416) );
  NAND4_X1 U17760 ( .A1(n14419), .A2(n14418), .A3(n14417), .A4(n14416), .ZN(
        n14425) );
  AOI22_X1 U17761 ( .A1(n12689), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14423) );
  AOI22_X1 U17762 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14422) );
  AOI22_X1 U17763 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15823), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14421) );
  AOI22_X1 U17764 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14420) );
  NAND4_X1 U17765 ( .A1(n14423), .A2(n14422), .A3(n14421), .A4(n14420), .ZN(
        n14424) );
  NOR2_X1 U17766 ( .A1(n14425), .A2(n14424), .ZN(n16940) );
  AOI22_X1 U17767 ( .A1(n12689), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17132), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14429) );
  AOI22_X1 U17768 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14428) );
  AOI22_X1 U17769 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14427) );
  AOI22_X1 U17770 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14426) );
  NAND4_X1 U17771 ( .A1(n14429), .A2(n14428), .A3(n14427), .A4(n14426), .ZN(
        n14435) );
  AOI22_X1 U17772 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14433) );
  AOI22_X1 U17773 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14432) );
  AOI22_X1 U17774 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14431) );
  AOI22_X1 U17775 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14430) );
  NAND4_X1 U17776 ( .A1(n14433), .A2(n14432), .A3(n14431), .A4(n14430), .ZN(
        n14434) );
  NOR2_X1 U17777 ( .A1(n14435), .A2(n14434), .ZN(n16946) );
  AOI22_X1 U17778 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12703), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14445) );
  AOI22_X1 U17779 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14444) );
  AOI22_X1 U17780 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14436) );
  OAI21_X1 U17781 ( .B1(n14457), .B2(n17146), .A(n14436), .ZN(n14442) );
  AOI22_X1 U17782 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14440) );
  AOI22_X1 U17783 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14439) );
  AOI22_X1 U17784 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14438) );
  AOI22_X1 U17785 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14437) );
  NAND4_X1 U17786 ( .A1(n14440), .A2(n14439), .A3(n14438), .A4(n14437), .ZN(
        n14441) );
  AOI211_X1 U17787 ( .C1(n17045), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n14442), .B(n14441), .ZN(n14443) );
  NAND3_X1 U17788 ( .A1(n14445), .A2(n14444), .A3(n14443), .ZN(n16953) );
  AOI22_X1 U17789 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17125), .ZN(n14455) );
  AOI22_X1 U17790 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17132), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14454) );
  AOI22_X1 U17791 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n17127), .ZN(n14446) );
  OAI21_X1 U17792 ( .B1(n20813), .B2(n9635), .A(n14446), .ZN(n14452) );
  AOI22_X1 U17793 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n17108), .ZN(n14450) );
  AOI22_X1 U17794 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17159), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17109), .ZN(n14449) );
  AOI22_X1 U17795 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n17149), .ZN(n14448) );
  AOI22_X1 U17796 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n14458), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14447) );
  NAND4_X1 U17797 ( .A1(n14450), .A2(n14449), .A3(n14448), .A4(n14447), .ZN(
        n14451) );
  AOI211_X1 U17798 ( .C1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .C2(n12689), .A(
        n14452), .B(n14451), .ZN(n14453) );
  NAND3_X1 U17799 ( .A1(n14455), .A2(n14454), .A3(n14453), .ZN(n16954) );
  NAND2_X1 U17800 ( .A1(n16953), .A2(n16954), .ZN(n16952) );
  NOR2_X1 U17801 ( .A1(n16946), .A2(n16952), .ZN(n16944) );
  AOI22_X1 U17802 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12692), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14467) );
  AOI22_X1 U17803 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14466) );
  AOI22_X1 U17804 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14456) );
  OAI21_X1 U17805 ( .B1(n14457), .B2(n17191), .A(n14456), .ZN(n14464) );
  AOI22_X1 U17806 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14462) );
  AOI22_X1 U17807 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14461) );
  AOI22_X1 U17808 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14460) );
  AOI22_X1 U17809 ( .A1(n12689), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14459) );
  NAND4_X1 U17810 ( .A1(n14462), .A2(n14461), .A3(n14460), .A4(n14459), .ZN(
        n14463) );
  AOI211_X1 U17811 ( .C1(n17159), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n14464), .B(n14463), .ZN(n14465) );
  NAND3_X1 U17812 ( .A1(n14467), .A2(n14466), .A3(n14465), .ZN(n16943) );
  NAND2_X1 U17813 ( .A1(n16944), .A2(n16943), .ZN(n16942) );
  NOR2_X1 U17814 ( .A1(n16940), .A2(n16942), .ZN(n16937) );
  AOI22_X1 U17815 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14478) );
  AOI22_X1 U17816 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14477) );
  AOI22_X1 U17817 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14468) );
  OAI21_X1 U17818 ( .B1(n14469), .B2(n20795), .A(n14468), .ZN(n14475) );
  AOI22_X1 U17819 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n15823), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14473) );
  AOI22_X1 U17820 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14472) );
  AOI22_X1 U17821 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12703), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14471) );
  AOI22_X1 U17822 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14470) );
  NAND4_X1 U17823 ( .A1(n14473), .A2(n14472), .A3(n14471), .A4(n14470), .ZN(
        n14474) );
  AOI211_X1 U17824 ( .C1(n17159), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n14475), .B(n14474), .ZN(n14476) );
  NAND3_X1 U17825 ( .A1(n14478), .A2(n14477), .A3(n14476), .ZN(n16936) );
  NAND2_X1 U17826 ( .A1(n16937), .A2(n16936), .ZN(n16935) );
  NOR3_X1 U17827 ( .A1(n16930), .A2(n16929), .A3(n16935), .ZN(n14479) );
  XNOR2_X1 U17828 ( .A(n14480), .B(n14479), .ZN(n17214) );
  INV_X1 U17829 ( .A(n17214), .ZN(n14488) );
  INV_X1 U17830 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16643) );
  INV_X1 U17831 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n14485) );
  INV_X1 U17832 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16982) );
  INV_X1 U17833 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17020) );
  INV_X1 U17834 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17050) );
  NOR2_X1 U17835 ( .A1(n18207), .A2(n18225), .ZN(n14481) );
  INV_X1 U17836 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n16903) );
  INV_X1 U17837 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17200) );
  INV_X1 U17838 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17194) );
  NOR2_X1 U17839 ( .A1(n17200), .A2(n17194), .ZN(n17189) );
  INV_X1 U17840 ( .A(n17189), .ZN(n16904) );
  NOR2_X1 U17841 ( .A1(n16903), .A2(n16904), .ZN(n17179) );
  NAND3_X1 U17842 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17179), .ZN(n17172) );
  NAND3_X1 U17843 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .A3(n17176), .ZN(n17166) );
  NAND3_X1 U17844 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(n17080), .ZN(n17036) );
  NAND2_X1 U17845 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n15820), .ZN(n16979) );
  AND2_X1 U17846 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n15821) );
  NAND4_X1 U17847 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(n15821), .ZN(n14484) );
  NAND3_X1 U17848 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(P3_EBX_REG_29__SCAN_IN), 
        .A3(n16927), .ZN(n16926) );
  INV_X1 U17849 ( .A(n16926), .ZN(n16924) );
  AOI21_X1 U17850 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16927), .A(
        P3_EBX_REG_30__SCAN_IN), .ZN(n14486) );
  NOR2_X1 U17851 ( .A1(n16924), .A2(n14486), .ZN(n14487) );
  MUX2_X1 U17852 ( .A(n14488), .B(n14487), .S(n17192), .Z(P3_U2673) );
  INV_X1 U17853 ( .A(n14489), .ZN(n14516) );
  AOI21_X1 U17854 ( .B1(n16060), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14490), .ZN(n14491) );
  OAI21_X1 U17855 ( .B1(n16069), .B2(n14492), .A(n14491), .ZN(n14493) );
  AOI21_X1 U17856 ( .B1(n14494), .B2(n16065), .A(n14493), .ZN(n14495) );
  OAI21_X1 U17857 ( .B1(n14516), .B2(n20055), .A(n14495), .ZN(P1_U2968) );
  INV_X1 U17858 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20672) );
  INV_X1 U17859 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n14496) );
  NAND2_X1 U17860 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n14746) );
  NAND2_X1 U17861 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n15982) );
  NOR3_X1 U17862 ( .A1(n14496), .A2(n14746), .A3(n15982), .ZN(n14725) );
  NAND2_X1 U17863 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n14725), .ZN(n14710) );
  NOR3_X1 U17864 ( .A1(n14498), .A2(n14497), .A3(n14710), .ZN(n14499) );
  NAND3_X1 U17865 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .A3(n14499), .ZN(n14501) );
  AND3_X1 U17866 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(P1_REIP_REG_20__SCAN_IN), .ZN(n14502) );
  NAND2_X1 U17867 ( .A1(n14692), .A2(n14502), .ZN(n14657) );
  NAND2_X1 U17868 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14500) );
  NOR2_X1 U17869 ( .A1(n14657), .A2(n14500), .ZN(n14641) );
  NAND2_X1 U17870 ( .A1(n14641), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14621) );
  NAND3_X1 U17871 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .A3(P1_REIP_REG_26__SCAN_IN), .ZN(n14506) );
  NAND2_X1 U17872 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14508) );
  NAND2_X1 U17873 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14510) );
  NOR3_X1 U17874 ( .A1(n14532), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14510), 
        .ZN(n14513) );
  NOR3_X1 U17875 ( .A1(n19972), .A2(n14501), .A3(n20672), .ZN(n14675) );
  NAND2_X1 U17876 ( .A1(n14675), .A2(n14502), .ZN(n14503) );
  NAND3_X1 U17877 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .A3(P1_REIP_REG_22__SCAN_IN), .ZN(n14504) );
  AND2_X1 U17878 ( .A1(n19888), .A2(n14504), .ZN(n14505) );
  AND2_X1 U17879 ( .A1(n19888), .A2(n14506), .ZN(n14507) );
  NOR2_X1 U17880 ( .A1(n14640), .A2(n14507), .ZN(n14607) );
  NAND2_X1 U17881 ( .A1(n19888), .A2(n14508), .ZN(n14509) );
  NAND2_X1 U17882 ( .A1(n14607), .A2(n14509), .ZN(n14577) );
  AOI21_X1 U17883 ( .B1(n14510), .B2(n19888), .A(n14577), .ZN(n14536) );
  AOI22_X1 U17884 ( .A1(n9585), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19959), .ZN(n14511) );
  OAI21_X1 U17885 ( .B1(n14536), .B2(n20696), .A(n14511), .ZN(n14512) );
  AOI211_X1 U17886 ( .C1(n14514), .C2(n19971), .A(n14513), .B(n14512), .ZN(
        n14515) );
  OAI21_X1 U17887 ( .B1(n14516), .B2(n19903), .A(n14515), .ZN(P1_U2809) );
  NOR2_X1 U17888 ( .A1(n14517), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14520) );
  NOR2_X1 U17889 ( .A1(n14518), .A2(n15020), .ZN(n14519) );
  MUX2_X1 U17890 ( .A(n14520), .B(n14519), .S(n15131), .Z(n14521) );
  XNOR2_X1 U17891 ( .A(n14521), .B(n15010), .ZN(n15008) );
  NAND2_X1 U17892 ( .A1(n16055), .A2(n14533), .ZN(n14522) );
  NAND2_X1 U17893 ( .A1(n16118), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n15011) );
  OAI211_X1 U17894 ( .C1(n14973), .C2(n20877), .A(n14522), .B(n15011), .ZN(
        n14523) );
  AOI21_X1 U17895 ( .B1(n15008), .B2(n16065), .A(n14523), .ZN(n14524) );
  OAI21_X1 U17896 ( .B1(n14540), .B2(n20055), .A(n14524), .ZN(P1_U2969) );
  NOR3_X1 U17897 ( .A1(n14861), .A2(n14525), .A3(n20093), .ZN(n14834) );
  INV_X1 U17898 ( .A(DATAI_14_), .ZN(n14527) );
  NAND2_X1 U17899 ( .A1(n20053), .A2(BUF1_REG_14__SCAN_IN), .ZN(n14526) );
  OAI21_X1 U17900 ( .B1(n20053), .B2(n14527), .A(n14526), .ZN(n20036) );
  AOI22_X1 U17901 ( .A1(n14834), .A2(n20036), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n14861), .ZN(n14528) );
  OAI21_X1 U17902 ( .B1(n14529), .B2(n14836), .A(n14528), .ZN(n14530) );
  AOI21_X1 U17903 ( .B1(n12532), .B2(DATAI_30_), .A(n14530), .ZN(n14531) );
  OAI21_X1 U17904 ( .B1(n14540), .B2(n14869), .A(n14531), .ZN(P1_U2874) );
  INV_X1 U17905 ( .A(n14532), .ZN(n14570) );
  AOI21_X1 U17906 ( .B1(n14570), .B2(P1_REIP_REG_29__SCAN_IN), .A(
        P1_REIP_REG_30__SCAN_IN), .ZN(n14537) );
  AOI22_X1 U17907 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19959), .B1(
        n19958), .B2(n14533), .ZN(n14535) );
  NAND2_X1 U17908 ( .A1(n9585), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n14534) );
  OAI211_X1 U17909 ( .C1(n14537), .C2(n14536), .A(n14535), .B(n14534), .ZN(
        n14538) );
  AOI21_X1 U17910 ( .B1(n12509), .B2(n19971), .A(n14538), .ZN(n14539) );
  OAI21_X1 U17911 ( .B1(n14540), .B2(n19903), .A(n14539), .ZN(P1_U2810) );
  XNOR2_X1 U17912 ( .A(n14541), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15427) );
  NAND2_X1 U17913 ( .A1(n14542), .A2(n15429), .ZN(n14547) );
  INV_X1 U17914 ( .A(n14543), .ZN(n14545) );
  NAND2_X1 U17915 ( .A1(n14545), .A2(n14544), .ZN(n14546) );
  XNOR2_X1 U17916 ( .A(n14547), .B(n14546), .ZN(n15425) );
  AOI21_X1 U17917 ( .B1(n15579), .B2(n15581), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14549) );
  NOR2_X1 U17918 ( .A1(n15534), .A2(n14551), .ZN(n15420) );
  AOI21_X1 U17919 ( .B1(n15425), .B2(n16300), .A(n14552), .ZN(n14553) );
  OAI21_X1 U17920 ( .B1(n15427), .B2(n19137), .A(n14553), .ZN(P2_U3016) );
  NOR2_X1 U17921 ( .A1(n11787), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14554) );
  AOI21_X1 U17922 ( .B1(n9594), .B2(n14555), .A(n14554), .ZN(n15905) );
  INV_X1 U17923 ( .A(n15905), .ZN(n14557) );
  OAI22_X1 U17924 ( .A1(n16149), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20705), .ZN(n14556) );
  AOI21_X1 U17925 ( .B1(n14557), .B2(n14558), .A(n14556), .ZN(n14561) );
  AOI21_X1 U17926 ( .B1(n15903), .B2(n14558), .A(n14560), .ZN(n14559) );
  OAI22_X1 U17927 ( .A1(n14561), .A2(n14560), .B1(n14559), .B2(n9840), .ZN(
        P1_U3474) );
  NAND2_X1 U17928 ( .A1(n14562), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n14565)
         );
  NAND3_X1 U17929 ( .A1(n14565), .A2(n14564), .A3(n14563), .ZN(P1_U2801) );
  INV_X1 U17930 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20692) );
  OAI22_X1 U17931 ( .A1(n12456), .A2(n19975), .B1(n19983), .B2(n14874), .ZN(
        n14566) );
  AOI21_X1 U17932 ( .B1(n9585), .B2(P1_EBX_REG_29__SCAN_IN), .A(n14566), .ZN(
        n14568) );
  NAND2_X1 U17933 ( .A1(n14577), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14567) );
  OAI211_X1 U17934 ( .C1(n15019), .C2(n19968), .A(n14568), .B(n14567), .ZN(
        n14569) );
  AOI21_X1 U17935 ( .B1(n14570), .B2(n20692), .A(n14569), .ZN(n14571) );
  OAI21_X1 U17936 ( .B1(n14877), .B2(n19903), .A(n14571), .ZN(P1_U2811) );
  NOR2_X1 U17937 ( .A1(n14591), .A2(n14574), .ZN(n14575) );
  INV_X1 U17938 ( .A(n15036), .ZN(n14585) );
  NAND2_X1 U17939 ( .A1(n14577), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14582) );
  INV_X1 U17940 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14579) );
  INV_X1 U17941 ( .A(n14578), .ZN(n14886) );
  OAI22_X1 U17942 ( .A1(n14579), .A2(n19975), .B1(n19983), .B2(n14886), .ZN(
        n14580) );
  AOI21_X1 U17943 ( .B1(n9585), .B2(P1_EBX_REG_28__SCAN_IN), .A(n14580), .ZN(
        n14581) );
  NAND2_X1 U17944 ( .A1(n14582), .A2(n14581), .ZN(n14584) );
  INV_X1 U17945 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n14894) );
  NOR3_X1 U17946 ( .A1(n14599), .A2(P1_REIP_REG_28__SCAN_IN), .A3(n14894), 
        .ZN(n14583) );
  AOI211_X1 U17947 ( .C1(n14585), .C2(n19971), .A(n14584), .B(n14583), .ZN(
        n14586) );
  OAI21_X1 U17948 ( .B1(n14889), .B2(n19903), .A(n14586), .ZN(P1_U2812) );
  AOI21_X1 U17949 ( .B1(n14588), .B2(n14587), .A(n14572), .ZN(n14758) );
  NAND2_X1 U17950 ( .A1(n14758), .A2(n19899), .ZN(n14598) );
  NOR2_X1 U17951 ( .A1(n14604), .A2(n14589), .ZN(n14590) );
  INV_X1 U17952 ( .A(n15041), .ZN(n14596) );
  OAI22_X1 U17953 ( .A1(n14592), .A2(n19975), .B1(n19983), .B2(n14896), .ZN(
        n14593) );
  AOI21_X1 U17954 ( .B1(n9585), .B2(P1_EBX_REG_27__SCAN_IN), .A(n14593), .ZN(
        n14594) );
  OAI21_X1 U17955 ( .B1(n14607), .B2(n14894), .A(n14594), .ZN(n14595) );
  AOI21_X1 U17956 ( .B1(n14596), .B2(n19971), .A(n14595), .ZN(n14597) );
  OAI211_X1 U17957 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14599), .A(n14598), 
        .B(n14597), .ZN(P1_U2813) );
  OAI21_X1 U17958 ( .B1(n14600), .B2(n14601), .A(n14587), .ZN(n14910) );
  AND2_X1 U17959 ( .A1(n14616), .A2(n14602), .ZN(n14603) );
  NOR2_X1 U17960 ( .A1(n14604), .A2(n14603), .ZN(n15050) );
  INV_X1 U17961 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n20866) );
  AOI22_X1 U17962 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19959), .B1(
        n19958), .B2(n14902), .ZN(n14606) );
  NAND2_X1 U17963 ( .A1(n9585), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n14605) );
  OAI211_X1 U17964 ( .C1(n14607), .C2(n20866), .A(n14606), .B(n14605), .ZN(
        n14609) );
  INV_X1 U17965 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14925) );
  INV_X1 U17966 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20684) );
  NOR4_X1 U17967 ( .A1(n14621), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n14925), 
        .A4(n20684), .ZN(n14608) );
  AOI211_X1 U17968 ( .C1(n15050), .C2(n19971), .A(n14609), .B(n14608), .ZN(
        n14610) );
  OAI21_X1 U17969 ( .B1(n14910), .B2(n19903), .A(n14610), .ZN(P1_U2814) );
  AOI21_X1 U17970 ( .B1(n14613), .B2(n14612), .A(n14600), .ZN(n14918) );
  INV_X1 U17971 ( .A(n14918), .ZN(n14818) );
  NAND2_X1 U17972 ( .A1(n14626), .A2(n14614), .ZN(n14615) );
  NAND2_X1 U17973 ( .A1(n14616), .A2(n14615), .ZN(n14761) );
  INV_X1 U17974 ( .A(n14761), .ZN(n15059) );
  INV_X1 U17975 ( .A(n14916), .ZN(n14617) );
  AOI22_X1 U17976 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19959), .B1(
        n19958), .B2(n14617), .ZN(n14618) );
  OAI21_X1 U17977 ( .B1(n19944), .B2(n14762), .A(n14618), .ZN(n14620) );
  NOR3_X1 U17978 ( .A1(n14621), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n14925), 
        .ZN(n14619) );
  AOI211_X1 U17979 ( .C1(n15059), .C2(n19971), .A(n14620), .B(n14619), .ZN(
        n14623) );
  NOR2_X1 U17980 ( .A1(n14621), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14631) );
  OAI21_X1 U17981 ( .B1(n14631), .B2(n14640), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14622) );
  OAI211_X1 U17982 ( .C1(n14818), .C2(n19903), .A(n14623), .B(n14622), .ZN(
        P1_U2815) );
  OAI21_X1 U17983 ( .B1(n14624), .B2(n14625), .A(n14612), .ZN(n14923) );
  AOI21_X1 U17984 ( .B1(n14627), .B2(n9627), .A(n9881), .ZN(n15069) );
  INV_X1 U17985 ( .A(n14640), .ZN(n14630) );
  AOI22_X1 U17986 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19959), .B1(
        n19958), .B2(n14924), .ZN(n14629) );
  NAND2_X1 U17987 ( .A1(n9585), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n14628) );
  OAI211_X1 U17988 ( .C1(n14630), .C2(n14925), .A(n14629), .B(n14628), .ZN(
        n14632) );
  AOI211_X1 U17989 ( .C1(n15069), .C2(n19971), .A(n14632), .B(n14631), .ZN(
        n14633) );
  OAI21_X1 U17990 ( .B1(n14923), .B2(n19903), .A(n14633), .ZN(P1_U2816) );
  XNOR2_X1 U17991 ( .A(n14634), .B(n14635), .ZN(n14937) );
  OAI22_X1 U17992 ( .A1(n14636), .A2(n19975), .B1(n19983), .B2(n14934), .ZN(
        n14639) );
  OAI21_X1 U17993 ( .B1(n14651), .B2(n14637), .A(n9627), .ZN(n14764) );
  NOR2_X1 U17994 ( .A1(n14764), .A2(n19968), .ZN(n14638) );
  AOI211_X1 U17995 ( .C1(n9585), .C2(P1_EBX_REG_23__SCAN_IN), .A(n14639), .B(
        n14638), .ZN(n14643) );
  OAI21_X1 U17996 ( .B1(n14641), .B2(P1_REIP_REG_23__SCAN_IN), .A(n14640), 
        .ZN(n14642) );
  OAI211_X1 U17997 ( .C1(n14937), .C2(n19903), .A(n14643), .B(n14642), .ZN(
        P1_U2817) );
  NAND2_X1 U17998 ( .A1(n14645), .A2(n14660), .ZN(n14831) );
  NOR2_X1 U17999 ( .A1(n14831), .A2(n14832), .ZN(n14830) );
  OAI21_X1 U18000 ( .B1(n14830), .B2(n14646), .A(n14634), .ZN(n14947) );
  INV_X1 U18001 ( .A(n15945), .ZN(n14649) );
  INV_X1 U18002 ( .A(n14647), .ZN(n14648) );
  AOI21_X1 U18003 ( .B1(n15946), .B2(n14649), .A(n14648), .ZN(n14650) );
  OR2_X1 U18004 ( .A1(n14651), .A2(n14650), .ZN(n15085) );
  INV_X1 U18005 ( .A(n15085), .ZN(n14656) );
  INV_X1 U18006 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14766) );
  AOI22_X1 U18007 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19959), .B1(
        n19958), .B2(n14941), .ZN(n14652) );
  OAI21_X1 U18008 ( .B1(n19944), .B2(n14766), .A(n14652), .ZN(n14655) );
  INV_X1 U18009 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n14653) );
  NOR3_X1 U18010 ( .A1(n14657), .A2(P1_REIP_REG_22__SCAN_IN), .A3(n14653), 
        .ZN(n14654) );
  AOI211_X1 U18011 ( .C1(n14656), .C2(n19971), .A(n14655), .B(n14654), .ZN(
        n14659) );
  NOR2_X1 U18012 ( .A1(n14657), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15967) );
  OAI21_X1 U18013 ( .B1(n15967), .B2(n15968), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14658) );
  OAI211_X1 U18014 ( .C1(n14947), .C2(n19903), .A(n14659), .B(n14658), .ZN(
        P1_U2818) );
  OAI21_X1 U18015 ( .B1(n14645), .B2(n14660), .A(n14831), .ZN(n14959) );
  INV_X1 U18016 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n15110) );
  NAND2_X1 U18017 ( .A1(n14692), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14677) );
  INV_X1 U18018 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20678) );
  OAI21_X1 U18019 ( .B1(n15110), .B2(n14677), .A(n20678), .ZN(n14666) );
  AND2_X1 U18020 ( .A1(n14672), .A2(n14661), .ZN(n14662) );
  OR2_X1 U18021 ( .A1(n14662), .A2(n15946), .ZN(n15102) );
  NOR2_X1 U18022 ( .A1(n15102), .A2(n19968), .ZN(n14665) );
  INV_X1 U18023 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14767) );
  AOI22_X1 U18024 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19959), .B1(
        n19958), .B2(n14954), .ZN(n14663) );
  OAI21_X1 U18025 ( .B1(n19944), .B2(n14767), .A(n14663), .ZN(n14664) );
  AOI211_X1 U18026 ( .C1(n14666), .C2(n15968), .A(n14665), .B(n14664), .ZN(
        n14667) );
  OAI21_X1 U18027 ( .B1(n14959), .B2(n19903), .A(n14667), .ZN(P1_U2820) );
  OR2_X1 U18028 ( .A1(n10145), .A2(n14645), .ZN(n16023) );
  NAND2_X1 U18029 ( .A1(n9659), .A2(n14670), .ZN(n14671) );
  AND2_X1 U18030 ( .A1(n14672), .A2(n14671), .ZN(n15116) );
  OAI21_X1 U18031 ( .B1(n19983), .B2(n16027), .A(n19918), .ZN(n14673) );
  AOI21_X1 U18032 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19959), .A(
        n14673), .ZN(n14674) );
  OAI21_X1 U18033 ( .B1(n19944), .B2(n14770), .A(n14674), .ZN(n14680) );
  INV_X1 U18034 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n14691) );
  NOR2_X1 U18035 ( .A1(n14676), .A2(n14675), .ZN(n14705) );
  AOI21_X1 U18036 ( .B1(n14692), .B2(n14691), .A(n14705), .ZN(n14678) );
  AOI22_X1 U18037 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n14678), .B1(n14677), 
        .B2(n15110), .ZN(n14679) );
  AOI211_X1 U18038 ( .C1(n15116), .C2(n19971), .A(n14680), .B(n14679), .ZN(
        n14681) );
  OAI21_X1 U18039 ( .B1(n16023), .B2(n19903), .A(n14681), .ZN(P1_U2821) );
  OAI21_X1 U18040 ( .B1(n9606), .B2(n12235), .A(n14668), .ZN(n14966) );
  OAI21_X1 U18041 ( .B1(n14699), .B2(n14683), .A(n9659), .ZN(n15127) );
  INV_X1 U18042 ( .A(n14684), .ZN(n14964) );
  INV_X1 U18043 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14687) );
  NOR2_X1 U18044 ( .A1(n19975), .A2(n14960), .ZN(n14685) );
  AOI211_X1 U18045 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n14705), .A(n19931), 
        .B(n14685), .ZN(n14686) );
  OAI21_X1 U18046 ( .B1(n14687), .B2(n19944), .A(n14686), .ZN(n14688) );
  AOI21_X1 U18047 ( .B1(n14964), .B2(n19958), .A(n14688), .ZN(n14689) );
  OAI21_X1 U18048 ( .B1(n15127), .B2(n19968), .A(n14689), .ZN(n14690) );
  AOI21_X1 U18049 ( .B1(n14692), .B2(n14691), .A(n14690), .ZN(n14693) );
  OAI21_X1 U18050 ( .B1(n14966), .B2(n19903), .A(n14693), .ZN(P1_U2822) );
  AOI21_X1 U18051 ( .B1(n14695), .B2(n14694), .A(n9606), .ZN(n16029) );
  INV_X1 U18052 ( .A(n16029), .ZN(n14854) );
  NAND2_X1 U18053 ( .A1(n20672), .A2(n14696), .ZN(n14706) );
  NOR2_X1 U18054 ( .A1(n14712), .A2(n14697), .ZN(n14698) );
  OR2_X1 U18055 ( .A1(n14699), .A2(n14698), .ZN(n15139) );
  OAI21_X1 U18056 ( .B1(n19975), .B2(n14700), .A(n19918), .ZN(n14702) );
  INV_X1 U18057 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14773) );
  NOR2_X1 U18058 ( .A1(n19944), .A2(n14773), .ZN(n14701) );
  AOI211_X1 U18059 ( .C1(n16028), .C2(n19958), .A(n14702), .B(n14701), .ZN(
        n14703) );
  OAI21_X1 U18060 ( .B1(n15139), .B2(n19968), .A(n14703), .ZN(n14704) );
  AOI21_X1 U18061 ( .B1(n14706), .B2(n14705), .A(n14704), .ZN(n14707) );
  OAI21_X1 U18062 ( .B1(n14854), .B2(n19903), .A(n14707), .ZN(P1_U2823) );
  OAI21_X1 U18063 ( .B1(n14708), .B2(n14709), .A(n14694), .ZN(n14974) );
  INV_X1 U18064 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20670) );
  NOR4_X1 U18065 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n14710), .A3(n20670), 
        .A4(n16000), .ZN(n14719) );
  NOR3_X1 U18066 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n14710), .A3(n16000), 
        .ZN(n15976) );
  INV_X1 U18067 ( .A(n14710), .ZN(n14711) );
  OAI21_X1 U18068 ( .B1(n14711), .B2(n19942), .A(n14748), .ZN(n15971) );
  OAI21_X1 U18069 ( .B1(n15976), .B2(n15971), .A(P1_REIP_REG_16__SCAN_IN), 
        .ZN(n14717) );
  AOI21_X1 U18070 ( .B1(n9678), .B2(n14713), .A(n14712), .ZN(n16073) );
  AOI22_X1 U18071 ( .A1(P1_EBX_REG_16__SCAN_IN), .A2(n9585), .B1(n19958), .B2(
        n14977), .ZN(n14714) );
  OAI211_X1 U18072 ( .C1(n19975), .C2(n14972), .A(n14714), .B(n19918), .ZN(
        n14715) );
  AOI21_X1 U18073 ( .B1(n16073), .B2(n19971), .A(n14715), .ZN(n14716) );
  NAND2_X1 U18074 ( .A1(n14717), .A2(n14716), .ZN(n14718) );
  NOR2_X1 U18075 ( .A1(n14719), .A2(n14718), .ZN(n14720) );
  OAI21_X1 U18076 ( .B1(n14974), .B2(n19903), .A(n14720), .ZN(P1_U2824) );
  INV_X1 U18077 ( .A(n14721), .ZN(n14786) );
  OAI21_X1 U18078 ( .B1(n14786), .B2(n12172), .A(n14724), .ZN(n14985) );
  OAI221_X1 U18079 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n14725), .C1(
        P1_REIP_REG_14__SCAN_IN), .C2(n14747), .A(n15971), .ZN(n14732) );
  INV_X1 U18080 ( .A(n14987), .ZN(n14730) );
  NAND2_X1 U18081 ( .A1(n14791), .A2(n14726), .ZN(n14727) );
  NAND2_X1 U18082 ( .A1(n14780), .A2(n14727), .ZN(n15147) );
  AOI22_X1 U18083 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19959), .B1(
        P1_EBX_REG_14__SCAN_IN), .B2(n9585), .ZN(n14728) );
  OAI211_X1 U18084 ( .C1(n19968), .C2(n15147), .A(n14728), .B(n19918), .ZN(
        n14729) );
  AOI21_X1 U18085 ( .B1(n19958), .B2(n14730), .A(n14729), .ZN(n14731) );
  OAI211_X1 U18086 ( .C1(n14985), .C2(n19903), .A(n14732), .B(n14731), .ZN(
        P1_U2826) );
  INV_X1 U18087 ( .A(n14733), .ZN(n14735) );
  NOR2_X1 U18088 ( .A1(n14735), .A2(n14734), .ZN(n14738) );
  INV_X1 U18089 ( .A(n14736), .ZN(n14737) );
  AOI21_X1 U18090 ( .B1(n14738), .B2(n14378), .A(n14737), .ZN(n14999) );
  INV_X1 U18091 ( .A(n14999), .ZN(n14870) );
  INV_X1 U18092 ( .A(n14997), .ZN(n14754) );
  INV_X1 U18093 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n14745) );
  AOI21_X1 U18094 ( .B1(n14741), .B2(n14740), .A(n14739), .ZN(n14742) );
  OR2_X1 U18095 ( .A1(n14742), .A2(n14789), .ZN(n16100) );
  INV_X1 U18096 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14794) );
  OAI22_X1 U18097 ( .A1(n16100), .A2(n19968), .B1(n19944), .B2(n14794), .ZN(
        n14743) );
  INV_X1 U18098 ( .A(n14743), .ZN(n14744) );
  OAI211_X1 U18099 ( .C1(n19975), .C2(n14745), .A(n14744), .B(n19918), .ZN(
        n14753) );
  INV_X1 U18100 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n14751) );
  INV_X1 U18101 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n14750) );
  INV_X1 U18102 ( .A(n14746), .ZN(n14749) );
  NAND2_X1 U18103 ( .A1(n14749), .A2(n14747), .ZN(n15998) );
  INV_X1 U18104 ( .A(n19942), .ZN(n19973) );
  OAI21_X1 U18105 ( .B1(n14749), .B2(n19942), .A(n14748), .ZN(n16002) );
  AOI21_X1 U18106 ( .B1(n19973), .B2(n15982), .A(n16002), .ZN(n15983) );
  AOI221_X1 U18107 ( .B1(n14751), .B2(n14750), .C1(n15998), .C2(n14750), .A(
        n15983), .ZN(n14752) );
  AOI211_X1 U18108 ( .C1(n19958), .C2(n14754), .A(n14753), .B(n14752), .ZN(
        n14755) );
  OAI21_X1 U18109 ( .B1(n14870), .B2(n19903), .A(n14755), .ZN(P1_U2828) );
  INV_X1 U18110 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14756) );
  INV_X1 U18111 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14757) );
  OAI222_X1 U18112 ( .A1(n15036), .A2(n19985), .B1(n14757), .B2(n19997), .C1(
        n14889), .C2(n19992), .ZN(P1_U2844) );
  INV_X1 U18113 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14759) );
  OAI222_X1 U18114 ( .A1(n15041), .A2(n19985), .B1(n14759), .B2(n19997), .C1(
        n14899), .C2(n19992), .ZN(P1_U2845) );
  AOI22_X1 U18115 ( .A1(n15050), .A2(n12508), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n12469), .ZN(n14760) );
  OAI21_X1 U18116 ( .B1(n14910), .B2(n19992), .A(n14760), .ZN(P1_U2846) );
  OAI222_X1 U18117 ( .A1(n14818), .A2(n19992), .B1(n14762), .B2(n19997), .C1(
        n14761), .C2(n19985), .ZN(P1_U2847) );
  AOI22_X1 U18118 ( .A1(n15069), .A2(n12508), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n12469), .ZN(n14763) );
  OAI21_X1 U18119 ( .B1(n14923), .B2(n19992), .A(n14763), .ZN(P1_U2848) );
  INV_X1 U18120 ( .A(n14764), .ZN(n15080) );
  AOI22_X1 U18121 ( .A1(n15080), .A2(n12508), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n12469), .ZN(n14765) );
  OAI21_X1 U18122 ( .B1(n14937), .B2(n19992), .A(n14765), .ZN(P1_U2849) );
  OAI222_X1 U18123 ( .A1(n15085), .A2(n19985), .B1(n14766), .B2(n19997), .C1(
        n14947), .C2(n19992), .ZN(P1_U2850) );
  OAI22_X1 U18124 ( .A1(n15102), .A2(n19985), .B1(n14767), .B2(n19997), .ZN(
        n14768) );
  INV_X1 U18125 ( .A(n14768), .ZN(n14769) );
  OAI21_X1 U18126 ( .B1(n14959), .B2(n19992), .A(n14769), .ZN(P1_U2852) );
  NOR2_X1 U18127 ( .A1(n19997), .A2(n14770), .ZN(n14771) );
  AOI21_X1 U18128 ( .B1(n15116), .B2(n12508), .A(n14771), .ZN(n14772) );
  OAI21_X1 U18129 ( .B1(n16023), .B2(n19992), .A(n14772), .ZN(P1_U2853) );
  OAI222_X1 U18130 ( .A1(n15127), .A2(n19985), .B1(n14687), .B2(n19997), .C1(
        n14966), .C2(n19992), .ZN(P1_U2854) );
  OAI22_X1 U18131 ( .A1(n15139), .A2(n19985), .B1(n14773), .B2(n19997), .ZN(
        n14774) );
  AOI21_X1 U18132 ( .B1(n16029), .B2(n16014), .A(n14774), .ZN(n14775) );
  INV_X1 U18133 ( .A(n14775), .ZN(P1_U2855) );
  AOI22_X1 U18134 ( .A1(n16073), .A2(n12508), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n12469), .ZN(n14776) );
  OAI21_X1 U18135 ( .B1(n14974), .B2(n19992), .A(n14776), .ZN(P1_U2856) );
  AND2_X1 U18136 ( .A1(n14724), .A2(n14777), .ZN(n14778) );
  OR2_X1 U18137 ( .A1(n14778), .A2(n14708), .ZN(n16041) );
  INV_X1 U18138 ( .A(n16041), .ZN(n15977) );
  NAND2_X1 U18139 ( .A1(n14780), .A2(n14779), .ZN(n14781) );
  NAND2_X1 U18140 ( .A1(n9678), .A2(n14781), .ZN(n16078) );
  OAI22_X1 U18141 ( .A1(n16078), .A2(n19985), .B1(n14782), .B2(n19997), .ZN(
        n14783) );
  AOI21_X1 U18142 ( .B1(n15977), .B2(n16014), .A(n14783), .ZN(n14784) );
  INV_X1 U18143 ( .A(n14784), .ZN(P1_U2857) );
  INV_X1 U18144 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14785) );
  OAI222_X1 U18145 ( .A1(n14985), .A2(n19992), .B1(n19997), .B2(n14785), .C1(
        n15147), .C2(n19985), .ZN(P1_U2858) );
  AOI21_X1 U18146 ( .B1(n14787), .B2(n14736), .A(n14786), .ZN(n16051) );
  OR2_X1 U18147 ( .A1(n14789), .A2(n14788), .ZN(n14790) );
  NAND2_X1 U18148 ( .A1(n14791), .A2(n14790), .ZN(n16085) );
  INV_X1 U18149 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15980) );
  OAI22_X1 U18150 ( .A1(n16085), .A2(n19985), .B1(n15980), .B2(n19997), .ZN(
        n14792) );
  AOI21_X1 U18151 ( .B1(n16051), .B2(n16014), .A(n14792), .ZN(n14793) );
  INV_X1 U18152 ( .A(n14793), .ZN(P1_U2859) );
  OAI222_X1 U18153 ( .A1(n16100), .A2(n19985), .B1(n14794), .B2(n19997), .C1(
        n14870), .C2(n19992), .ZN(P1_U2860) );
  INV_X1 U18154 ( .A(DATAI_13_), .ZN(n14796) );
  MUX2_X1 U18155 ( .A(n14796), .B(n14795), .S(n20053), .Z(n20033) );
  OAI22_X1 U18156 ( .A1(n14855), .A2(n20033), .B1(n14867), .B2(n14797), .ZN(
        n14798) );
  AOI21_X1 U18157 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n14857), .A(n14798), .ZN(
        n14800) );
  NAND2_X1 U18158 ( .A1(n12532), .A2(DATAI_29_), .ZN(n14799) );
  OAI211_X1 U18159 ( .C1(n14877), .C2(n14869), .A(n14800), .B(n14799), .ZN(
        P1_U2875) );
  INV_X1 U18160 ( .A(DATAI_12_), .ZN(n14801) );
  MUX2_X1 U18161 ( .A(n14801), .B(n16474), .S(n20053), .Z(n20030) );
  OAI22_X1 U18162 ( .A1(n14855), .A2(n20030), .B1(n14867), .B2(n14802), .ZN(
        n14803) );
  AOI21_X1 U18163 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n14857), .A(n14803), .ZN(
        n14805) );
  NAND2_X1 U18164 ( .A1(n12532), .A2(DATAI_28_), .ZN(n14804) );
  OAI211_X1 U18165 ( .C1(n14889), .C2(n14869), .A(n14805), .B(n14804), .ZN(
        P1_U2876) );
  INV_X1 U18166 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16450) );
  AOI22_X1 U18167 ( .A1(n14834), .A2(n14806), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n14861), .ZN(n14807) );
  OAI21_X1 U18168 ( .B1(n14836), .B2(n16450), .A(n14807), .ZN(n14808) );
  AOI21_X1 U18169 ( .B1(n12532), .B2(DATAI_27_), .A(n14808), .ZN(n14809) );
  OAI21_X1 U18170 ( .B1(n14899), .B2(n14869), .A(n14809), .ZN(P1_U2877) );
  OAI22_X1 U18171 ( .A1(n14855), .A2(n20027), .B1(n14867), .B2(n14810), .ZN(
        n14811) );
  AOI21_X1 U18172 ( .B1(n14857), .B2(BUF1_REG_26__SCAN_IN), .A(n14811), .ZN(
        n14813) );
  NAND2_X1 U18173 ( .A1(n12532), .A2(DATAI_26_), .ZN(n14812) );
  OAI211_X1 U18174 ( .C1(n14910), .C2(n14869), .A(n14813), .B(n14812), .ZN(
        P1_U2878) );
  OAI22_X1 U18175 ( .A1(n14855), .A2(n20023), .B1(n14867), .B2(n14814), .ZN(
        n14815) );
  AOI21_X1 U18176 ( .B1(n14857), .B2(BUF1_REG_25__SCAN_IN), .A(n14815), .ZN(
        n14817) );
  NAND2_X1 U18177 ( .A1(n12532), .A2(DATAI_25_), .ZN(n14816) );
  OAI211_X1 U18178 ( .C1(n14818), .C2(n14869), .A(n14817), .B(n14816), .ZN(
        P1_U2879) );
  OAI22_X1 U18179 ( .A1(n14855), .A2(n20020), .B1(n14867), .B2(n13424), .ZN(
        n14819) );
  AOI21_X1 U18180 ( .B1(n14857), .B2(BUF1_REG_24__SCAN_IN), .A(n14819), .ZN(
        n14821) );
  NAND2_X1 U18181 ( .A1(n12532), .A2(DATAI_24_), .ZN(n14820) );
  OAI211_X1 U18182 ( .C1(n14923), .C2(n14869), .A(n14821), .B(n14820), .ZN(
        P1_U2880) );
  OAI22_X1 U18183 ( .A1(n14855), .A2(n20107), .B1(n14867), .B2(n14822), .ZN(
        n14823) );
  AOI21_X1 U18184 ( .B1(n14857), .B2(BUF1_REG_23__SCAN_IN), .A(n14823), .ZN(
        n14825) );
  NAND2_X1 U18185 ( .A1(n12532), .A2(DATAI_23_), .ZN(n14824) );
  OAI211_X1 U18186 ( .C1(n14937), .C2(n14869), .A(n14825), .B(n14824), .ZN(
        P1_U2881) );
  OAI22_X1 U18187 ( .A1(n14855), .A2(n20099), .B1(n14867), .B2(n14826), .ZN(
        n14827) );
  AOI21_X1 U18188 ( .B1(n14857), .B2(BUF1_REG_22__SCAN_IN), .A(n14827), .ZN(
        n14829) );
  NAND2_X1 U18189 ( .A1(n12532), .A2(DATAI_22_), .ZN(n14828) );
  OAI211_X1 U18190 ( .C1(n14947), .C2(n14869), .A(n14829), .B(n14828), .ZN(
        P1_U2882) );
  AOI21_X1 U18191 ( .B1(n14832), .B2(n14831), .A(n14830), .ZN(n16018) );
  INV_X1 U18192 ( .A(n16018), .ZN(n14839) );
  AOI22_X1 U18193 ( .A1(n14834), .A2(n14833), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n14861), .ZN(n14835) );
  OAI21_X1 U18194 ( .B1(n20843), .B2(n14836), .A(n14835), .ZN(n14837) );
  AOI21_X1 U18195 ( .B1(n12532), .B2(DATAI_21_), .A(n14837), .ZN(n14838) );
  OAI21_X1 U18196 ( .B1(n14839), .B2(n14869), .A(n14838), .ZN(P1_U2883) );
  OAI22_X1 U18197 ( .A1(n14855), .A2(n20090), .B1(n14867), .B2(n13626), .ZN(
        n14840) );
  AOI21_X1 U18198 ( .B1(n14857), .B2(BUF1_REG_20__SCAN_IN), .A(n14840), .ZN(
        n14842) );
  NAND2_X1 U18199 ( .A1(n12532), .A2(DATAI_20_), .ZN(n14841) );
  OAI211_X1 U18200 ( .C1(n14959), .C2(n14869), .A(n14842), .B(n14841), .ZN(
        P1_U2884) );
  OAI22_X1 U18201 ( .A1(n14855), .A2(n20086), .B1(n14867), .B2(n14843), .ZN(
        n14844) );
  AOI21_X1 U18202 ( .B1(n14857), .B2(BUF1_REG_19__SCAN_IN), .A(n14844), .ZN(
        n14846) );
  NAND2_X1 U18203 ( .A1(n12532), .A2(DATAI_19_), .ZN(n14845) );
  OAI211_X1 U18204 ( .C1(n16023), .C2(n14869), .A(n14846), .B(n14845), .ZN(
        P1_U2885) );
  OAI22_X1 U18205 ( .A1(n14855), .A2(n20082), .B1(n14867), .B2(n14847), .ZN(
        n14848) );
  AOI21_X1 U18206 ( .B1(n14857), .B2(BUF1_REG_18__SCAN_IN), .A(n14848), .ZN(
        n14850) );
  NAND2_X1 U18207 ( .A1(n12532), .A2(DATAI_18_), .ZN(n14849) );
  OAI211_X1 U18208 ( .C1(n14966), .C2(n14869), .A(n14850), .B(n14849), .ZN(
        P1_U2886) );
  OAI22_X1 U18209 ( .A1(n14855), .A2(n20078), .B1(n14867), .B2(n13630), .ZN(
        n14851) );
  AOI21_X1 U18210 ( .B1(n14857), .B2(BUF1_REG_17__SCAN_IN), .A(n14851), .ZN(
        n14853) );
  NAND2_X1 U18211 ( .A1(n12532), .A2(DATAI_17_), .ZN(n14852) );
  OAI211_X1 U18212 ( .C1(n14854), .C2(n14869), .A(n14853), .B(n14852), .ZN(
        P1_U2887) );
  OAI22_X1 U18213 ( .A1(n14855), .A2(n20069), .B1(n14867), .B2(n13634), .ZN(
        n14856) );
  AOI21_X1 U18214 ( .B1(n14857), .B2(BUF1_REG_16__SCAN_IN), .A(n14856), .ZN(
        n14859) );
  NAND2_X1 U18215 ( .A1(n12532), .A2(DATAI_16_), .ZN(n14858) );
  OAI211_X1 U18216 ( .C1(n14974), .C2(n14869), .A(n14859), .B(n14858), .ZN(
        P1_U2888) );
  OAI222_X1 U18217 ( .A1(n14869), .A2(n16041), .B1(n14867), .B2(n13392), .C1(
        n14866), .C2(n14860), .ZN(P1_U2889) );
  INV_X1 U18218 ( .A(n14866), .ZN(n14862) );
  AOI22_X1 U18219 ( .A1(n14862), .A2(n20036), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14861), .ZN(n14863) );
  OAI21_X1 U18220 ( .B1(n14985), .B2(n14869), .A(n14863), .ZN(P1_U2890) );
  INV_X1 U18221 ( .A(n16051), .ZN(n14865) );
  INV_X1 U18222 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14864) );
  OAI222_X1 U18223 ( .A1(n14865), .A2(n14869), .B1(n14864), .B2(n14867), .C1(
        n14866), .C2(n20033), .ZN(P1_U2891) );
  OAI222_X1 U18224 ( .A1(n14870), .A2(n14869), .B1(n14868), .B2(n14867), .C1(
        n14866), .C2(n20030), .ZN(P1_U2892) );
  XNOR2_X1 U18225 ( .A(n15136), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14871) );
  XNOR2_X1 U18226 ( .A(n14872), .B(n14871), .ZN(n15018) );
  NOR2_X1 U18227 ( .A1(n16134), .A2(n20692), .ZN(n15023) );
  AOI21_X1 U18228 ( .B1(n16060), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15023), .ZN(n14873) );
  OAI21_X1 U18229 ( .B1(n16069), .B2(n14874), .A(n14873), .ZN(n14875) );
  AOI21_X1 U18230 ( .B1(n15018), .B2(n16065), .A(n14875), .ZN(n14876) );
  OAI21_X1 U18231 ( .B1(n14877), .B2(n20055), .A(n14876), .ZN(P1_U2970) );
  AOI21_X2 U18232 ( .B1(n14878), .B2(n15131), .A(n14932), .ZN(n14881) );
  INV_X1 U18233 ( .A(n14881), .ZN(n14880) );
  INV_X1 U18234 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14892) );
  INV_X1 U18235 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15052) );
  NAND4_X1 U18236 ( .A1(n14880), .A2(n14879), .A3(n14892), .A4(n15052), .ZN(
        n14883) );
  NAND3_X1 U18237 ( .A1(n14881), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14882) );
  MUX2_X1 U18238 ( .A(n14883), .B(n14882), .S(n15131), .Z(n14884) );
  XNOR2_X1 U18239 ( .A(n14884), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15038) );
  NAND2_X1 U18240 ( .A1(n16118), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15028) );
  NAND2_X1 U18241 ( .A1(n16060), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14885) );
  OAI211_X1 U18242 ( .C1(n16069), .C2(n14886), .A(n15028), .B(n14885), .ZN(
        n14887) );
  AOI21_X1 U18243 ( .B1(n15038), .B2(n16065), .A(n14887), .ZN(n14888) );
  OAI21_X1 U18244 ( .B1(n14889), .B2(n20055), .A(n14888), .ZN(P1_U2971) );
  MUX2_X1 U18245 ( .A(n14890), .B(n14891), .S(n15941), .Z(n14893) );
  XNOR2_X1 U18246 ( .A(n14893), .B(n14892), .ZN(n15040) );
  NOR2_X1 U18247 ( .A1(n16134), .A2(n14894), .ZN(n15043) );
  AOI21_X1 U18248 ( .B1(n16060), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15043), .ZN(n14895) );
  OAI21_X1 U18249 ( .B1(n16069), .B2(n14896), .A(n14895), .ZN(n14897) );
  AOI21_X1 U18250 ( .B1(n15040), .B2(n16065), .A(n14897), .ZN(n14898) );
  OAI21_X1 U18251 ( .B1(n14899), .B2(n20055), .A(n14898), .ZN(P1_U2972) );
  NOR2_X1 U18252 ( .A1(n16134), .A2(n20866), .ZN(n15049) );
  INV_X1 U18253 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14900) );
  NOR2_X1 U18254 ( .A1(n14973), .A2(n14900), .ZN(n14901) );
  AOI211_X1 U18255 ( .C1(n16055), .C2(n14902), .A(n15049), .B(n14901), .ZN(
        n14909) );
  INV_X1 U18256 ( .A(n14932), .ZN(n14904) );
  NAND2_X1 U18257 ( .A1(n14904), .A2(n14903), .ZN(n14905) );
  MUX2_X1 U18258 ( .A(n14906), .B(n14905), .S(n15131), .Z(n14907) );
  XNOR2_X1 U18259 ( .A(n14907), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15047) );
  NAND2_X1 U18260 ( .A1(n15047), .A2(n16065), .ZN(n14908) );
  OAI211_X1 U18261 ( .C1(n14910), .C2(n20055), .A(n14909), .B(n14908), .ZN(
        P1_U2973) );
  NAND2_X1 U18262 ( .A1(n14911), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14920) );
  INV_X1 U18263 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15070) );
  NAND2_X1 U18264 ( .A1(n14932), .A2(n15077), .ZN(n14912) );
  MUX2_X1 U18265 ( .A(n15070), .B(n14912), .S(n15941), .Z(n14913) );
  AOI21_X1 U18266 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14920), .A(
        n14913), .ZN(n14914) );
  XNOR2_X1 U18267 ( .A(n14914), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15064) );
  NOR2_X1 U18268 ( .A1(n16134), .A2(n20684), .ZN(n15058) );
  AOI21_X1 U18269 ( .B1(n16060), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15058), .ZN(n14915) );
  OAI21_X1 U18270 ( .B1(n16069), .B2(n14916), .A(n14915), .ZN(n14917) );
  AOI21_X1 U18271 ( .B1(n14918), .B2(n16066), .A(n14917), .ZN(n14919) );
  OAI21_X1 U18272 ( .B1(n19869), .B2(n15064), .A(n14919), .ZN(P1_U2974) );
  NAND2_X1 U18273 ( .A1(n14920), .A2(n14932), .ZN(n14921) );
  MUX2_X1 U18274 ( .A(n14921), .B(n14920), .S(n15136), .Z(n14922) );
  XOR2_X1 U18275 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n14922), .Z(
        n15073) );
  INV_X1 U18276 ( .A(n14923), .ZN(n14929) );
  INV_X1 U18277 ( .A(n14924), .ZN(n14927) );
  NOR2_X1 U18278 ( .A1(n16134), .A2(n14925), .ZN(n15068) );
  AOI21_X1 U18279 ( .B1(n16060), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15068), .ZN(n14926) );
  OAI21_X1 U18280 ( .B1(n16069), .B2(n14927), .A(n14926), .ZN(n14928) );
  AOI21_X1 U18281 ( .B1(n14929), .B2(n16066), .A(n14928), .ZN(n14930) );
  OAI21_X1 U18282 ( .B1(n19869), .B2(n15073), .A(n14930), .ZN(P1_U2975) );
  XNOR2_X1 U18283 ( .A(n15136), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14931) );
  XNOR2_X1 U18284 ( .A(n14932), .B(n14931), .ZN(n15075) );
  INV_X1 U18285 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20682) );
  NOR2_X1 U18286 ( .A1(n16134), .A2(n20682), .ZN(n15079) );
  AOI21_X1 U18287 ( .B1(n16060), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15079), .ZN(n14933) );
  OAI21_X1 U18288 ( .B1(n16069), .B2(n14934), .A(n14933), .ZN(n14935) );
  AOI21_X1 U18289 ( .B1(n15075), .B2(n16065), .A(n14935), .ZN(n14936) );
  OAI21_X1 U18290 ( .B1(n14937), .B2(n20055), .A(n14936), .ZN(P1_U2976) );
  INV_X1 U18291 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n14938) );
  NOR2_X1 U18292 ( .A1(n16134), .A2(n14938), .ZN(n15087) );
  INV_X1 U18293 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14939) );
  NOR2_X1 U18294 ( .A1(n14973), .A2(n14939), .ZN(n14940) );
  AOI211_X1 U18295 ( .C1(n16055), .C2(n14941), .A(n15087), .B(n14940), .ZN(
        n14946) );
  NAND2_X1 U18296 ( .A1(n14943), .A2(n14942), .ZN(n14944) );
  XNOR2_X1 U18297 ( .A(n14944), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15084) );
  NAND2_X1 U18298 ( .A1(n15084), .A2(n16065), .ZN(n14945) );
  OAI211_X1 U18299 ( .C1(n14947), .C2(n20055), .A(n14946), .B(n14945), .ZN(
        P1_U2977) );
  NAND2_X1 U18300 ( .A1(n15131), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14952) );
  INV_X1 U18301 ( .A(n14949), .ZN(n14951) );
  NAND3_X1 U18302 ( .A1(n14951), .A2(n15941), .A3(n14950), .ZN(n15943) );
  OAI21_X1 U18303 ( .B1(n14948), .B2(n14952), .A(n15943), .ZN(n14953) );
  XNOR2_X1 U18304 ( .A(n14953), .B(n15104), .ZN(n15094) );
  NAND2_X1 U18305 ( .A1(n16055), .A2(n14954), .ZN(n14955) );
  NAND2_X1 U18306 ( .A1(n16118), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15100) );
  OAI211_X1 U18307 ( .C1(n14956), .C2(n14973), .A(n14955), .B(n15100), .ZN(
        n14957) );
  AOI21_X1 U18308 ( .B1(n15094), .B2(n16065), .A(n14957), .ZN(n14958) );
  OAI21_X1 U18309 ( .B1(n14959), .B2(n20055), .A(n14958), .ZN(P1_U2979) );
  NAND2_X1 U18310 ( .A1(n16118), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15125) );
  OAI21_X1 U18311 ( .B1(n14973), .B2(n14960), .A(n15125), .ZN(n14963) );
  OAI21_X1 U18312 ( .B1(n14949), .B2(n14961), .A(n14948), .ZN(n15130) );
  NOR2_X1 U18313 ( .A1(n15130), .A2(n19869), .ZN(n14962) );
  AOI211_X1 U18314 ( .C1(n16055), .C2(n14964), .A(n14963), .B(n14962), .ZN(
        n14965) );
  OAI21_X1 U18315 ( .B1(n14966), .B2(n20055), .A(n14965), .ZN(P1_U2981) );
  INV_X1 U18316 ( .A(n14980), .ZN(n16046) );
  OAI21_X1 U18317 ( .B1(n15001), .B2(n14967), .A(n16046), .ZN(n16035) );
  OAI21_X1 U18318 ( .B1(n16035), .B2(n14968), .A(n16036), .ZN(n14969) );
  XOR2_X1 U18319 ( .A(n14970), .B(n14969), .Z(n16072) );
  INV_X1 U18320 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14971) );
  OAI22_X1 U18321 ( .A1(n14973), .A2(n14972), .B1(n16134), .B2(n14971), .ZN(
        n14976) );
  NOR2_X1 U18322 ( .A1(n14974), .A2(n20055), .ZN(n14975) );
  AOI211_X1 U18323 ( .C1(n16055), .C2(n14977), .A(n14976), .B(n14975), .ZN(
        n14978) );
  OAI21_X1 U18324 ( .B1(n19869), .B2(n16072), .A(n14978), .ZN(P1_U2983) );
  INV_X1 U18325 ( .A(n15001), .ZN(n15154) );
  OAI21_X1 U18326 ( .B1(n15154), .B2(n14980), .A(n14979), .ZN(n14982) );
  NAND2_X1 U18327 ( .A1(n14982), .A2(n14981), .ZN(n14984) );
  XNOR2_X1 U18328 ( .A(n15136), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14983) );
  XNOR2_X1 U18329 ( .A(n14984), .B(n14983), .ZN(n15152) );
  INV_X1 U18330 ( .A(n14985), .ZN(n14989) );
  AOI22_X1 U18331 ( .A1(n16060), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16118), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n14986) );
  OAI21_X1 U18332 ( .B1(n16069), .B2(n14987), .A(n14986), .ZN(n14988) );
  AOI21_X1 U18333 ( .B1(n14989), .B2(n16066), .A(n14988), .ZN(n14990) );
  OAI21_X1 U18334 ( .B1(n15152), .B2(n19869), .A(n14990), .ZN(P1_U2985) );
  NAND2_X1 U18335 ( .A1(n9846), .A2(n14991), .ZN(n14995) );
  OR2_X1 U18336 ( .A1(n15001), .A2(n14992), .ZN(n16047) );
  NAND2_X1 U18337 ( .A1(n16047), .A2(n14993), .ZN(n14994) );
  XOR2_X1 U18338 ( .A(n14995), .B(n14994), .Z(n16103) );
  NOR2_X1 U18339 ( .A1(n16134), .A2(n14750), .ZN(n16101) );
  AOI21_X1 U18340 ( .B1(n16060), .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16101), .ZN(n14996) );
  OAI21_X1 U18341 ( .B1(n16069), .B2(n14997), .A(n14996), .ZN(n14998) );
  AOI21_X1 U18342 ( .B1(n14999), .B2(n16066), .A(n14998), .ZN(n15000) );
  OAI21_X1 U18343 ( .B1(n16103), .B2(n19869), .A(n15000), .ZN(P1_U2987) );
  INV_X1 U18344 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15159) );
  NOR3_X1 U18345 ( .A1(n15001), .A2(n15941), .A3(n15159), .ZN(n15157) );
  NOR3_X1 U18346 ( .A1(n15153), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15136), .ZN(n15002) );
  NOR2_X1 U18347 ( .A1(n15157), .A2(n15002), .ZN(n15003) );
  XNOR2_X1 U18348 ( .A(n15003), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16114) );
  INV_X1 U18349 ( .A(n16114), .ZN(n15007) );
  NOR2_X1 U18350 ( .A1(n16134), .A2(n14751), .ZN(n16111) );
  AOI21_X1 U18351 ( .B1(n16060), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16111), .ZN(n15004) );
  OAI21_X1 U18352 ( .B1(n16069), .B2(n15993), .A(n15004), .ZN(n15005) );
  AOI21_X1 U18353 ( .B1(n15995), .B2(n16066), .A(n15005), .ZN(n15006) );
  OAI21_X1 U18354 ( .B1(n15007), .B2(n19869), .A(n15006), .ZN(P1_U2988) );
  INV_X1 U18355 ( .A(n15008), .ZN(n15017) );
  INV_X1 U18356 ( .A(n15009), .ZN(n15027) );
  OAI21_X1 U18357 ( .B1(n15027), .B2(n15020), .A(n15010), .ZN(n15014) );
  OAI21_X1 U18358 ( .B1(n15012), .B2(n16136), .A(n15011), .ZN(n15013) );
  AOI21_X1 U18359 ( .B1(n15015), .B2(n15014), .A(n15013), .ZN(n15016) );
  OAI21_X1 U18360 ( .B1(n15017), .B2(n16137), .A(n15016), .ZN(P1_U3001) );
  NAND2_X1 U18361 ( .A1(n15018), .A2(n16122), .ZN(n15026) );
  INV_X1 U18362 ( .A(n15019), .ZN(n15024) );
  NOR2_X1 U18363 ( .A1(n15021), .A2(n15020), .ZN(n15022) );
  AOI211_X1 U18364 ( .C1(n15024), .C2(n16119), .A(n15023), .B(n15022), .ZN(
        n15025) );
  OAI211_X1 U18365 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15027), .A(
        n15026), .B(n15025), .ZN(P1_U3002) );
  INV_X1 U18366 ( .A(n15028), .ZN(n15029) );
  AOI21_X1 U18367 ( .B1(n9605), .B2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15029), .ZN(n15035) );
  INV_X1 U18368 ( .A(n15046), .ZN(n15033) );
  INV_X1 U18369 ( .A(n15030), .ZN(n15031) );
  NAND3_X1 U18370 ( .A1(n15033), .A2(n15032), .A3(n15031), .ZN(n15034) );
  OAI211_X1 U18371 ( .C1(n15036), .C2(n16136), .A(n15035), .B(n15034), .ZN(
        n15037) );
  AOI21_X1 U18372 ( .B1(n15038), .B2(n16122), .A(n15037), .ZN(n15039) );
  INV_X1 U18373 ( .A(n15039), .ZN(P1_U3003) );
  NAND2_X1 U18374 ( .A1(n15040), .A2(n16122), .ZN(n15045) );
  NOR2_X1 U18375 ( .A1(n15041), .A2(n16136), .ZN(n15042) );
  AOI211_X1 U18376 ( .C1(n9605), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15043), .B(n15042), .ZN(n15044) );
  OAI211_X1 U18377 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15046), .A(
        n15045), .B(n15044), .ZN(P1_U3004) );
  INV_X1 U18378 ( .A(n15047), .ZN(n15055) );
  NOR2_X1 U18379 ( .A1(n15056), .A2(n15052), .ZN(n15048) );
  AOI211_X1 U18380 ( .C1(n15050), .C2(n16119), .A(n15049), .B(n15048), .ZN(
        n15054) );
  INV_X1 U18381 ( .A(n15051), .ZN(n15061) );
  NAND3_X1 U18382 ( .A1(n15061), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n15052), .ZN(n15053) );
  OAI211_X1 U18383 ( .C1(n15055), .C2(n16137), .A(n15054), .B(n15053), .ZN(
        P1_U3005) );
  NOR2_X1 U18384 ( .A1(n15056), .A2(n15060), .ZN(n15057) );
  AOI211_X1 U18385 ( .C1(n15059), .C2(n16119), .A(n15058), .B(n15057), .ZN(
        n15063) );
  NAND2_X1 U18386 ( .A1(n15061), .A2(n15060), .ZN(n15062) );
  OAI211_X1 U18387 ( .C1(n15064), .C2(n16137), .A(n15063), .B(n15062), .ZN(
        P1_U3006) );
  NAND2_X1 U18388 ( .A1(n16099), .A2(n15077), .ZN(n15066) );
  AOI21_X1 U18389 ( .B1(n15066), .B2(n15065), .A(n15070), .ZN(n15067) );
  AOI211_X1 U18390 ( .C1(n15069), .C2(n16119), .A(n15068), .B(n15067), .ZN(
        n15072) );
  NAND3_X1 U18391 ( .A1(n15074), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n15070), .ZN(n15071) );
  OAI211_X1 U18392 ( .C1(n15073), .C2(n16137), .A(n15072), .B(n15071), .ZN(
        P1_U3007) );
  INV_X1 U18393 ( .A(n15074), .ZN(n15083) );
  NAND2_X1 U18394 ( .A1(n15075), .A2(n16122), .ZN(n15082) );
  NOR2_X1 U18395 ( .A1(n15077), .A2(n15076), .ZN(n15078) );
  AOI211_X1 U18396 ( .C1(n15080), .C2(n16119), .A(n15079), .B(n15078), .ZN(
        n15081) );
  OAI211_X1 U18397 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n15083), .A(
        n15082), .B(n15081), .ZN(P1_U3008) );
  INV_X1 U18398 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15093) );
  INV_X1 U18399 ( .A(n15940), .ZN(n15092) );
  NAND2_X1 U18400 ( .A1(n15084), .A2(n16122), .ZN(n15091) );
  AOI21_X1 U18401 ( .B1(n11937), .B2(n15093), .A(n15949), .ZN(n15089) );
  NOR2_X1 U18402 ( .A1(n15085), .A2(n16136), .ZN(n15086) );
  AOI211_X1 U18403 ( .C1(n15089), .C2(n15088), .A(n15087), .B(n15086), .ZN(
        n15090) );
  OAI211_X1 U18404 ( .C1(n15093), .C2(n15092), .A(n15091), .B(n15090), .ZN(
        P1_U3009) );
  INV_X1 U18405 ( .A(n15094), .ZN(n15107) );
  NOR3_X1 U18406 ( .A1(n15097), .A2(n15096), .A3(n15095), .ZN(n15098) );
  NOR2_X1 U18407 ( .A1(n15098), .A2(n15111), .ZN(n15099) );
  NAND2_X1 U18408 ( .A1(n15099), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15101) );
  OAI211_X1 U18409 ( .C1(n15102), .C2(n16136), .A(n15101), .B(n15100), .ZN(
        n15103) );
  AOI21_X1 U18410 ( .B1(n15105), .B2(n15104), .A(n15103), .ZN(n15106) );
  OAI21_X1 U18411 ( .B1(n15107), .B2(n16137), .A(n15106), .ZN(P1_U3011) );
  NOR2_X1 U18412 ( .A1(n15131), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15108) );
  MUX2_X1 U18413 ( .A(n15136), .B(n15108), .S(n14948), .Z(n15109) );
  XNOR2_X1 U18414 ( .A(n15109), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16022) );
  NOR2_X1 U18415 ( .A1(n16134), .A2(n15110), .ZN(n15115) );
  AOI21_X1 U18416 ( .B1(n15113), .B2(n15112), .A(n15111), .ZN(n15114) );
  AOI211_X1 U18417 ( .C1(n16119), .C2(n15116), .A(n15115), .B(n15114), .ZN(
        n15117) );
  OAI21_X1 U18418 ( .B1(n16022), .B2(n16137), .A(n15117), .ZN(P1_U3012) );
  NOR2_X1 U18419 ( .A1(n16092), .A2(n15118), .ZN(n15120) );
  AOI211_X1 U18420 ( .C1(n15121), .C2(n15144), .A(n15120), .B(n15119), .ZN(
        n16091) );
  OAI21_X1 U18421 ( .B1(n16071), .B2(n15122), .A(n16091), .ZN(n15141) );
  NOR2_X1 U18422 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15123), .ZN(
        n15124) );
  NAND2_X1 U18423 ( .A1(n15138), .A2(n15124), .ZN(n15126) );
  OAI211_X1 U18424 ( .C1(n15127), .C2(n16136), .A(n15126), .B(n15125), .ZN(
        n15128) );
  AOI21_X1 U18425 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15141), .A(
        n15128), .ZN(n15129) );
  OAI21_X1 U18426 ( .B1(n15130), .B2(n16137), .A(n15129), .ZN(P1_U3013) );
  NOR2_X1 U18427 ( .A1(n15131), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15135) );
  OAI21_X1 U18428 ( .B1(n15154), .B2(n15133), .A(n15132), .ZN(n15134) );
  MUX2_X1 U18429 ( .A(n15136), .B(n15135), .S(n15134), .Z(n15137) );
  XOR2_X1 U18430 ( .A(n11923), .B(n15137), .Z(n16032) );
  NAND2_X1 U18431 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16070) );
  NAND2_X1 U18432 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15138), .ZN(
        n16084) );
  OAI21_X1 U18433 ( .B1(n16070), .B2(n16084), .A(n11923), .ZN(n15142) );
  OAI22_X1 U18434 ( .A1(n15139), .A2(n16136), .B1(n16134), .B2(n20672), .ZN(
        n15140) );
  AOI21_X1 U18435 ( .B1(n15142), .B2(n15141), .A(n15140), .ZN(n15143) );
  OAI21_X1 U18436 ( .B1(n16032), .B2(n16137), .A(n15143), .ZN(P1_U3014) );
  INV_X1 U18437 ( .A(n16091), .ZN(n15150) );
  NOR3_X1 U18438 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15145), .A3(
        n15144), .ZN(n15149) );
  INV_X1 U18439 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n15146) );
  OAI22_X1 U18440 ( .A1(n15147), .A2(n16136), .B1(n15146), .B2(n16134), .ZN(
        n15148) );
  AOI211_X1 U18441 ( .C1(n15150), .C2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15149), .B(n15148), .ZN(n15151) );
  OAI21_X1 U18442 ( .B1(n15152), .B2(n16137), .A(n15151), .ZN(P1_U3017) );
  XOR2_X1 U18443 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n15153), .Z(
        n15156) );
  NOR2_X1 U18444 ( .A1(n15154), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15155) );
  MUX2_X1 U18445 ( .A(n15156), .B(n15155), .S(n15131), .Z(n15158) );
  OR2_X1 U18446 ( .A1(n15158), .A2(n15157), .ZN(n16059) );
  AOI22_X1 U18447 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(n11751), .B2(n15159), .ZN(
        n15160) );
  AOI22_X1 U18448 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15162), .B1(
        n15161), .B2(n15160), .ZN(n15164) );
  AOI22_X1 U18449 ( .A1(n16003), .A2(n16119), .B1(n16118), .B2(
        P1_REIP_REG_10__SCAN_IN), .ZN(n15163) );
  OAI211_X1 U18450 ( .C1(n16059), .C2(n16137), .A(n15164), .B(n15163), .ZN(
        P1_U3021) );
  NAND4_X1 U18451 ( .A1(n15165), .A2(n18984), .A3(n9949), .A4(n15423), .ZN(
        n15173) );
  INV_X1 U18452 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19782) );
  NAND3_X1 U18453 ( .A1(n19109), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n16360), 
        .ZN(n15168) );
  INV_X1 U18454 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n15166) );
  OR2_X1 U18455 ( .A1(n18974), .A2(n15166), .ZN(n15167) );
  OAI211_X1 U18456 ( .C1(n18987), .C2(n19782), .A(n15168), .B(n15167), .ZN(
        n15170) );
  NOR2_X1 U18457 ( .A1(n19004), .A2(n18989), .ZN(n15169) );
  AOI211_X1 U18458 ( .C1(n13236), .C2(n15171), .A(n15170), .B(n15169), .ZN(
        n15172) );
  OAI211_X1 U18459 ( .C1(n15276), .C2(n18978), .A(n15173), .B(n15172), .ZN(
        P2_U2824) );
  NAND2_X1 U18460 ( .A1(n11044), .A2(n15174), .ZN(n15175) );
  INV_X1 U18461 ( .A(n13169), .ZN(n15182) );
  NAND2_X1 U18462 ( .A1(n11305), .A2(n15180), .ZN(n15181) );
  NAND2_X1 U18463 ( .A1(n15182), .A2(n15181), .ZN(n15577) );
  AOI22_X1 U18464 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19000), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n18951), .ZN(n15184) );
  NAND2_X1 U18465 ( .A1(n18992), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15183) );
  OAI211_X1 U18466 ( .C1(n15577), .C2(n18989), .A(n15184), .B(n15183), .ZN(
        n15185) );
  AOI21_X1 U18467 ( .B1(n15186), .B2(n13236), .A(n15185), .ZN(n15187) );
  OAI211_X1 U18468 ( .C1(n15573), .C2(n18978), .A(n15188), .B(n15187), .ZN(
        P2_U2826) );
  OAI211_X1 U18469 ( .C1(n9952), .C2(n15189), .A(n18984), .B(n9618), .ZN(
        n15195) );
  NOR2_X1 U18470 ( .A1(n15360), .A2(n18989), .ZN(n15192) );
  AOI22_X1 U18471 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n18992), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n18951), .ZN(n15190) );
  OAI21_X1 U18472 ( .B1(n9928), .B2(n18974), .A(n15190), .ZN(n15191) );
  AOI211_X1 U18473 ( .C1(n15193), .C2(n13236), .A(n15192), .B(n15191), .ZN(
        n15194) );
  OAI211_X1 U18474 ( .C1(n18978), .C2(n15287), .A(n15195), .B(n15194), .ZN(
        P2_U2827) );
  AOI21_X1 U18475 ( .B1(n15197), .B2(n15443), .A(n15196), .ZN(n15198) );
  NAND2_X1 U18476 ( .A1(n15198), .A2(n18984), .ZN(n15211) );
  INV_X1 U18477 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n15200) );
  AOI22_X1 U18478 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19000), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n18951), .ZN(n15199) );
  OAI21_X1 U18479 ( .B1(n15201), .B2(n15200), .A(n15199), .ZN(n15209) );
  INV_X1 U18480 ( .A(n15202), .ZN(n15207) );
  INV_X1 U18481 ( .A(n15203), .ZN(n15206) );
  INV_X1 U18482 ( .A(n15204), .ZN(n15205) );
  AOI211_X1 U18483 ( .C1(n15207), .C2(n15206), .A(n18995), .B(n15205), .ZN(
        n15208) );
  AOI211_X1 U18484 ( .C1(n18954), .C2(n15365), .A(n15209), .B(n15208), .ZN(
        n15210) );
  OAI211_X1 U18485 ( .C1(n18978), .C2(n15440), .A(n15211), .B(n15210), .ZN(
        P2_U2828) );
  INV_X1 U18486 ( .A(n11286), .ZN(n15212) );
  OAI21_X1 U18487 ( .B1(n15233), .B2(n15213), .A(n15212), .ZN(n15595) );
  NAND2_X1 U18488 ( .A1(n15237), .A2(n15214), .ZN(n15215) );
  AND2_X1 U18489 ( .A1(n15216), .A2(n15215), .ZN(n15592) );
  AOI22_X1 U18490 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n18992), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19000), .ZN(n15222) );
  INV_X1 U18491 ( .A(n15218), .ZN(n15219) );
  AOI211_X1 U18492 ( .C1(n15452), .C2(n15217), .A(n19717), .B(n15219), .ZN(
        n15220) );
  INV_X1 U18493 ( .A(n15220), .ZN(n15221) );
  OAI211_X1 U18494 ( .C1(n18987), .C2(n15223), .A(n15222), .B(n15221), .ZN(
        n15226) );
  AOI211_X1 U18495 ( .C1(P2_EBX_REG_26__SCAN_IN), .C2(n9646), .A(n18995), .B(
        n15224), .ZN(n15225) );
  AOI211_X1 U18496 ( .C1(n15592), .C2(n18954), .A(n15226), .B(n15225), .ZN(
        n15227) );
  OAI21_X1 U18497 ( .B1(n15595), .B2(n18978), .A(n15227), .ZN(P2_U2829) );
  AOI211_X1 U18498 ( .C1(n15228), .C2(n15465), .A(n19717), .B(n15229), .ZN(
        n15230) );
  INV_X1 U18499 ( .A(n15230), .ZN(n15242) );
  AND2_X1 U18500 ( .A1(n15312), .A2(n15231), .ZN(n15232) );
  NOR2_X1 U18501 ( .A1(n15233), .A2(n15232), .ZN(n15608) );
  NAND2_X1 U18502 ( .A1(n15234), .A2(n15235), .ZN(n15236) );
  NAND2_X1 U18503 ( .A1(n15237), .A2(n15236), .ZN(n15606) );
  AOI22_X1 U18504 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19000), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n18951), .ZN(n15239) );
  NAND2_X1 U18505 ( .A1(n18992), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n15238) );
  OAI211_X1 U18506 ( .C1(n15606), .C2(n18989), .A(n15239), .B(n15238), .ZN(
        n15240) );
  AOI21_X1 U18507 ( .B1(n15608), .B2(n18999), .A(n15240), .ZN(n15241) );
  OAI211_X1 U18508 ( .C1(n18995), .C2(n15243), .A(n15242), .B(n15241), .ZN(
        P2_U2830) );
  NAND2_X1 U18509 ( .A1(n15244), .A2(n15245), .ZN(n15246) );
  NAND2_X1 U18510 ( .A1(n15310), .A2(n15246), .ZN(n15631) );
  NOR2_X1 U18511 ( .A1(n15248), .A2(n15249), .ZN(n15250) );
  AOI22_X1 U18512 ( .A1(P2_EBX_REG_23__SCAN_IN), .A2(n18992), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n18951), .ZN(n15251) );
  OAI21_X1 U18513 ( .B1(n15484), .B2(n18974), .A(n15251), .ZN(n15252) );
  AOI21_X1 U18514 ( .B1(n9658), .B2(n18954), .A(n15252), .ZN(n15253) );
  OAI21_X1 U18515 ( .B1(n15631), .B2(n18978), .A(n15253), .ZN(n15257) );
  AOI211_X1 U18516 ( .C1(n15254), .C2(n15487), .A(n19717), .B(n15255), .ZN(
        n15256) );
  AOI211_X1 U18517 ( .C1(n13236), .C2(n15258), .A(n15257), .B(n15256), .ZN(
        n15259) );
  INV_X1 U18518 ( .A(n15259), .ZN(P2_U2832) );
  AOI211_X1 U18519 ( .C1(n15260), .C2(n15522), .A(n19717), .B(n15261), .ZN(
        n15274) );
  INV_X1 U18520 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15262) );
  OAI22_X1 U18521 ( .A1(n15263), .A2(n18995), .B1(n18974), .B2(n15262), .ZN(
        n15264) );
  AOI211_X1 U18522 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n18992), .A(n19113), .B(
        n15264), .ZN(n15265) );
  OAI21_X1 U18523 ( .B1(n19760), .B2(n18987), .A(n15265), .ZN(n15273) );
  NAND2_X1 U18524 ( .A1(n14172), .A2(n15266), .ZN(n15267) );
  NAND2_X1 U18525 ( .A1(n15336), .A2(n15267), .ZN(n15674) );
  NOR2_X1 U18526 ( .A1(n15269), .A2(n15270), .ZN(n15271) );
  OR2_X1 U18527 ( .A1(n15268), .A2(n15271), .ZN(n15408) );
  OAI22_X1 U18528 ( .A1(n15674), .A2(n18978), .B1(n18989), .B2(n15408), .ZN(
        n15272) );
  OR3_X1 U18529 ( .A1(n15274), .A2(n15273), .A3(n15272), .ZN(P2_U2836) );
  NAND2_X1 U18530 ( .A1(n15347), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n15275) );
  OAI21_X1 U18531 ( .B1(n15276), .B2(n13618), .A(n15275), .ZN(P2_U2856) );
  OR2_X1 U18532 ( .A1(n15278), .A2(n15277), .ZN(n15351) );
  NAND3_X1 U18533 ( .A1(n15351), .A2(n15279), .A3(n15342), .ZN(n15281) );
  NAND2_X1 U18534 ( .A1(n15347), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15280) );
  OAI211_X1 U18535 ( .C1(n15347), .C2(n15573), .A(n15281), .B(n15280), .ZN(
        P2_U2858) );
  NAND2_X1 U18536 ( .A1(n9975), .A2(n15282), .ZN(n15284) );
  XNOR2_X1 U18537 ( .A(n15284), .B(n15283), .ZN(n15362) );
  NAND2_X1 U18538 ( .A1(n15362), .A2(n15342), .ZN(n15286) );
  NAND2_X1 U18539 ( .A1(n15347), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n15285) );
  OAI211_X1 U18540 ( .C1(n15287), .C2(n13618), .A(n15286), .B(n15285), .ZN(
        P2_U2859) );
  OAI21_X1 U18541 ( .B1(n15288), .B2(n15290), .A(n15289), .ZN(n15368) );
  NOR2_X1 U18542 ( .A1(n15440), .A2(n13618), .ZN(n15291) );
  AOI21_X1 U18543 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n13618), .A(n15291), .ZN(
        n15292) );
  OAI21_X1 U18544 ( .B1(n15368), .B2(n15350), .A(n15292), .ZN(P2_U2860) );
  AOI21_X1 U18545 ( .B1(n15293), .B2(n15295), .A(n15294), .ZN(n15369) );
  NAND2_X1 U18546 ( .A1(n15369), .A2(n15342), .ZN(n15297) );
  NAND2_X1 U18547 ( .A1(n15347), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15296) );
  OAI211_X1 U18548 ( .C1(n15595), .C2(n15347), .A(n15297), .B(n15296), .ZN(
        P2_U2861) );
  OAI21_X1 U18549 ( .B1(n15298), .B2(n15300), .A(n15299), .ZN(n15381) );
  NOR2_X1 U18550 ( .A1(n15316), .A2(n15301), .ZN(n15302) );
  AOI21_X1 U18551 ( .B1(n15608), .B2(n15316), .A(n15302), .ZN(n15303) );
  OAI21_X1 U18552 ( .B1(n15381), .B2(n15350), .A(n15303), .ZN(P2_U2862) );
  AOI21_X1 U18553 ( .B1(n15304), .B2(n15306), .A(n15305), .ZN(n15308) );
  XNOR2_X1 U18554 ( .A(n15308), .B(n15307), .ZN(n15387) );
  NAND2_X1 U18555 ( .A1(n15387), .A2(n15342), .ZN(n15314) );
  NAND2_X1 U18556 ( .A1(n15310), .A2(n15309), .ZN(n15311) );
  AND2_X1 U18557 ( .A1(n15312), .A2(n15311), .ZN(n16160) );
  NAND2_X1 U18558 ( .A1(n16160), .A2(n15316), .ZN(n15313) );
  OAI211_X1 U18559 ( .C1(n15316), .C2(n15315), .A(n15314), .B(n15313), .ZN(
        P2_U2863) );
  INV_X1 U18560 ( .A(n15318), .ZN(n15319) );
  AOI21_X1 U18561 ( .B1(n15317), .B2(n15320), .A(n15319), .ZN(n15321) );
  INV_X1 U18562 ( .A(n15321), .ZN(n15393) );
  MUX2_X1 U18563 ( .A(n15631), .B(n10916), .S(n15347), .Z(n15322) );
  OAI21_X1 U18564 ( .B1(n15393), .B2(n15350), .A(n15322), .ZN(P2_U2864) );
  AOI21_X1 U18565 ( .B1(n15325), .B2(n15324), .A(n13016), .ZN(n15326) );
  INV_X1 U18566 ( .A(n15326), .ZN(n15400) );
  OAI21_X1 U18567 ( .B1(n15328), .B2(n15327), .A(n15244), .ZN(n15896) );
  NOR2_X1 U18568 ( .A1(n15896), .A2(n13618), .ZN(n15329) );
  AOI21_X1 U18569 ( .B1(P2_EBX_REG_22__SCAN_IN), .B2(n13618), .A(n15329), .ZN(
        n15330) );
  OAI21_X1 U18570 ( .B1(n15400), .B2(n15350), .A(n15330), .ZN(P2_U2865) );
  INV_X1 U18571 ( .A(n15331), .ZN(n15332) );
  OAI21_X1 U18572 ( .B1(n15332), .B2(n10137), .A(n15324), .ZN(n15407) );
  MUX2_X1 U18573 ( .A(n18892), .B(n15333), .S(n15347), .Z(n15334) );
  OAI21_X1 U18574 ( .B1(n15407), .B2(n15350), .A(n15334), .ZN(P2_U2866) );
  AND2_X1 U18575 ( .A1(n15336), .A2(n15335), .ZN(n15338) );
  OR2_X1 U18576 ( .A1(n15338), .A2(n15337), .ZN(n18899) );
  OR2_X1 U18577 ( .A1(n15339), .A2(n15340), .ZN(n15341) );
  AND2_X1 U18578 ( .A1(n15341), .A2(n15331), .ZN(n16164) );
  NAND2_X1 U18579 ( .A1(n16164), .A2(n15342), .ZN(n15344) );
  NAND2_X1 U18580 ( .A1(n15347), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n15343) );
  OAI211_X1 U18581 ( .C1(n18899), .C2(n15347), .A(n15344), .B(n15343), .ZN(
        P2_U2867) );
  INV_X1 U18582 ( .A(n15339), .ZN(n15345) );
  OAI21_X1 U18583 ( .B1(n9676), .B2(n15346), .A(n15345), .ZN(n15418) );
  MUX2_X1 U18584 ( .A(n15674), .B(n15348), .S(n15347), .Z(n15349) );
  OAI21_X1 U18585 ( .B1(n15418), .B2(n15350), .A(n15349), .ZN(P2_U2868) );
  NAND3_X1 U18586 ( .A1(n15351), .A2(n15279), .A3(n13149), .ZN(n15357) );
  INV_X1 U18587 ( .A(n15577), .ZN(n15354) );
  OAI22_X1 U18588 ( .A1(n15410), .A2(n19021), .B1(n19041), .B2(n15352), .ZN(
        n15353) );
  AOI21_X1 U18589 ( .B1(n15354), .B2(n19056), .A(n15353), .ZN(n15356) );
  AOI22_X1 U18590 ( .A1(n19011), .A2(BUF2_REG_29__SCAN_IN), .B1(n19010), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n15355) );
  NAND3_X1 U18591 ( .A1(n15357), .A2(n15356), .A3(n15355), .ZN(P2_U2890) );
  AOI22_X1 U18592 ( .A1(n19009), .A2(n19023), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n19055), .ZN(n15359) );
  AOI22_X1 U18593 ( .A1(n19011), .A2(BUF2_REG_28__SCAN_IN), .B1(n19010), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15358) );
  OAI211_X1 U18594 ( .C1(n15360), .C2(n15385), .A(n15359), .B(n15358), .ZN(
        n15361) );
  AOI21_X1 U18595 ( .B1(n15362), .B2(n13149), .A(n15361), .ZN(n15363) );
  INV_X1 U18596 ( .A(n15363), .ZN(P2_U2891) );
  OAI22_X1 U18597 ( .A1(n15410), .A2(n19026), .B1(n19041), .B2(n20882), .ZN(
        n15364) );
  AOI21_X1 U18598 ( .B1(n15365), .B2(n19056), .A(n15364), .ZN(n15367) );
  AOI22_X1 U18599 ( .A1(n19011), .A2(BUF2_REG_27__SCAN_IN), .B1(n19010), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15366) );
  OAI211_X1 U18600 ( .C1(n15368), .C2(n19060), .A(n15367), .B(n15366), .ZN(
        P2_U2892) );
  INV_X1 U18601 ( .A(n15369), .ZN(n15375) );
  INV_X1 U18602 ( .A(n19028), .ZN(n15371) );
  OAI22_X1 U18603 ( .A1(n15410), .A2(n15371), .B1(n19041), .B2(n15370), .ZN(
        n15372) );
  AOI21_X1 U18604 ( .B1(n15592), .B2(n19056), .A(n15372), .ZN(n15374) );
  AOI22_X1 U18605 ( .A1(n19011), .A2(BUF2_REG_26__SCAN_IN), .B1(n19010), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15373) );
  OAI211_X1 U18606 ( .C1(n15375), .C2(n19060), .A(n15374), .B(n15373), .ZN(
        P2_U2893) );
  INV_X1 U18607 ( .A(n15606), .ZN(n15378) );
  OAI22_X1 U18608 ( .A1(n15410), .A2(n19031), .B1(n19041), .B2(n15376), .ZN(
        n15377) );
  AOI21_X1 U18609 ( .B1(n15378), .B2(n19056), .A(n15377), .ZN(n15380) );
  AOI22_X1 U18610 ( .A1(n19011), .A2(BUF2_REG_25__SCAN_IN), .B1(n19010), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15379) );
  OAI211_X1 U18611 ( .C1(n15381), .C2(n19060), .A(n15380), .B(n15379), .ZN(
        P2_U2894) );
  OAI21_X1 U18612 ( .B1(n15247), .B2(n15382), .A(n15234), .ZN(n16158) );
  AOI22_X1 U18613 ( .A1(n19011), .A2(BUF2_REG_24__SCAN_IN), .B1(n19010), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n15384) );
  AOI22_X1 U18614 ( .A1(n19009), .A2(n19034), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n19055), .ZN(n15383) );
  OAI211_X1 U18615 ( .C1(n15385), .C2(n16158), .A(n15384), .B(n15383), .ZN(
        n15386) );
  AOI21_X1 U18616 ( .B1(n15387), .B2(n13149), .A(n15386), .ZN(n15388) );
  INV_X1 U18617 ( .A(n15388), .ZN(P2_U2895) );
  OAI22_X1 U18618 ( .A1(n15410), .A2(n19169), .B1(n19041), .B2(n15389), .ZN(
        n15390) );
  AOI21_X1 U18619 ( .B1(n19056), .B2(n9658), .A(n15390), .ZN(n15392) );
  AOI22_X1 U18620 ( .A1(n19011), .A2(BUF2_REG_23__SCAN_IN), .B1(n19010), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n15391) );
  OAI211_X1 U18621 ( .C1(n15393), .C2(n19060), .A(n15392), .B(n15391), .ZN(
        P2_U2896) );
  AND2_X1 U18622 ( .A1(n15395), .A2(n15394), .ZN(n15396) );
  NOR2_X1 U18623 ( .A1(n15248), .A2(n15396), .ZN(n15894) );
  OAI22_X1 U18624 ( .A1(n15410), .A2(n19038), .B1(n19041), .B2(n11238), .ZN(
        n15398) );
  INV_X1 U18625 ( .A(n19011), .ZN(n15414) );
  OAI22_X1 U18626 ( .A1(n15414), .A2(n20902), .B1(n15412), .B2(n16459), .ZN(
        n15397) );
  AOI211_X1 U18627 ( .C1(n19056), .C2(n15894), .A(n15398), .B(n15397), .ZN(
        n15399) );
  OAI21_X1 U18628 ( .B1(n15400), .B2(n19060), .A(n15399), .ZN(P2_U2897) );
  XNOR2_X1 U18629 ( .A(n15401), .B(n10032), .ZN(n18893) );
  OAI22_X1 U18630 ( .A1(n15410), .A2(n19040), .B1(n19041), .B2(n15403), .ZN(
        n15405) );
  OAI22_X1 U18631 ( .A1(n15414), .A2(n18212), .B1(n15412), .B2(n20843), .ZN(
        n15404) );
  AOI211_X1 U18632 ( .C1(n19056), .C2(n18893), .A(n15405), .B(n15404), .ZN(
        n15406) );
  OAI21_X1 U18633 ( .B1(n15407), .B2(n19060), .A(n15406), .ZN(P2_U2898) );
  INV_X1 U18634 ( .A(n15408), .ZN(n15673) );
  OAI22_X1 U18635 ( .A1(n15410), .A2(n19155), .B1(n19041), .B2(n15409), .ZN(
        n15416) );
  INV_X1 U18636 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n15413) );
  INV_X1 U18637 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n15411) );
  OAI22_X1 U18638 ( .A1(n15414), .A2(n15413), .B1(n15412), .B2(n15411), .ZN(
        n15415) );
  AOI211_X1 U18639 ( .C1(n19056), .C2(n15673), .A(n15416), .B(n15415), .ZN(
        n15417) );
  OAI21_X1 U18640 ( .B1(n15418), .B2(n19060), .A(n15417), .ZN(P2_U2900) );
  NAND2_X1 U18641 ( .A1(n15419), .A2(n19117), .ZN(n15422) );
  AOI21_X1 U18642 ( .B1(n19114), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15420), .ZN(n15421) );
  OAI211_X1 U18643 ( .C1(n19125), .C2(n15423), .A(n15422), .B(n15421), .ZN(
        n15424) );
  AOI21_X1 U18644 ( .B1(n15425), .B2(n19121), .A(n15424), .ZN(n15426) );
  OAI21_X1 U18645 ( .B1(n15427), .B2(n16256), .A(n15426), .ZN(P2_U2984) );
  NAND2_X1 U18646 ( .A1(n15430), .A2(n15429), .ZN(n15431) );
  XOR2_X1 U18647 ( .A(n15428), .B(n15431), .Z(n15590) );
  NAND2_X1 U18648 ( .A1(n15571), .A2(n19118), .ZN(n15437) );
  NAND2_X1 U18649 ( .A1(n19113), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15575) );
  OAI21_X1 U18650 ( .B1(n16265), .B2(n15432), .A(n15575), .ZN(n15434) );
  NOR2_X1 U18651 ( .A1(n15573), .A2(n16247), .ZN(n15433) );
  AOI211_X1 U18652 ( .C1(n16255), .C2(n15435), .A(n15434), .B(n15433), .ZN(
        n15436) );
  OAI211_X1 U18653 ( .C1(n15590), .C2(n16258), .A(n15437), .B(n15436), .ZN(
        P2_U2985) );
  OAI21_X1 U18654 ( .B1(n16265), .B2(n15439), .A(n15438), .ZN(n15442) );
  NOR2_X1 U18655 ( .A1(n15440), .A2(n16247), .ZN(n15441) );
  AOI211_X1 U18656 ( .C1(n16255), .C2(n15443), .A(n15442), .B(n15441), .ZN(
        n15446) );
  NAND3_X1 U18657 ( .A1(n15444), .A2(n11285), .A3(n19121), .ZN(n15445) );
  OAI211_X1 U18658 ( .C1(n15447), .C2(n16256), .A(n15446), .B(n15445), .ZN(
        P2_U2987) );
  OAI21_X1 U18659 ( .B1(n15448), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11281), .ZN(n15602) );
  NAND2_X1 U18660 ( .A1(n19113), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15594) );
  OAI21_X1 U18661 ( .B1(n16265), .B2(n15449), .A(n15594), .ZN(n15451) );
  NOR2_X1 U18662 ( .A1(n15595), .A2(n16247), .ZN(n15450) );
  AOI211_X1 U18663 ( .C1(n16255), .C2(n15452), .A(n15451), .B(n15450), .ZN(
        n15458) );
  INV_X1 U18664 ( .A(n15459), .ZN(n15454) );
  OAI21_X1 U18665 ( .B1(n15461), .B2(n15454), .A(n15460), .ZN(n15456) );
  XNOR2_X1 U18666 ( .A(n15456), .B(n15455), .ZN(n15599) );
  NAND2_X1 U18667 ( .A1(n15599), .A2(n19121), .ZN(n15457) );
  OAI211_X1 U18668 ( .C1(n15602), .C2(n16256), .A(n15458), .B(n15457), .ZN(
        P2_U2988) );
  NAND2_X1 U18669 ( .A1(n15460), .A2(n15459), .ZN(n15462) );
  XOR2_X1 U18670 ( .A(n15462), .B(n15461), .Z(n15615) );
  INV_X1 U18671 ( .A(n15448), .ZN(n15604) );
  NAND2_X1 U18672 ( .A1(n15463), .A2(n15464), .ZN(n15603) );
  NAND3_X1 U18673 ( .A1(n15604), .A2(n19118), .A3(n15603), .ZN(n15470) );
  NAND2_X1 U18674 ( .A1(n16255), .A2(n15465), .ZN(n15466) );
  NAND2_X1 U18675 ( .A1(n19113), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15605) );
  OAI211_X1 U18676 ( .C1(n16265), .C2(n15467), .A(n15466), .B(n15605), .ZN(
        n15468) );
  AOI21_X1 U18677 ( .B1(n15608), .B2(n19117), .A(n15468), .ZN(n15469) );
  OAI211_X1 U18678 ( .C1(n16258), .C2(n15615), .A(n15470), .B(n15469), .ZN(
        P2_U2989) );
  OAI21_X1 U18679 ( .B1(n15471), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15463), .ZN(n15626) );
  NAND2_X1 U18680 ( .A1(n19113), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15620) );
  NAND2_X1 U18681 ( .A1(n19114), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15472) );
  OAI211_X1 U18682 ( .C1(n19125), .C2(n15473), .A(n15620), .B(n15472), .ZN(
        n15474) );
  AOI21_X1 U18683 ( .B1(n16160), .B2(n19117), .A(n15474), .ZN(n15480) );
  NAND2_X1 U18684 ( .A1(n10883), .A2(n15476), .ZN(n15477) );
  XNOR2_X1 U18685 ( .A(n15478), .B(n15477), .ZN(n15624) );
  NAND2_X1 U18686 ( .A1(n15624), .A2(n19121), .ZN(n15479) );
  OAI211_X1 U18687 ( .C1(n15626), .C2(n16256), .A(n15480), .B(n15479), .ZN(
        P2_U2990) );
  INV_X1 U18688 ( .A(n15481), .ZN(n15483) );
  INV_X1 U18689 ( .A(n15471), .ZN(n15482) );
  OAI21_X1 U18690 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15483), .A(
        n15482), .ZN(n15627) );
  OR2_X1 U18691 ( .A1(n15534), .A2(n19767), .ZN(n15628) );
  OAI21_X1 U18692 ( .B1(n16265), .B2(n15484), .A(n15628), .ZN(n15486) );
  NOR2_X1 U18693 ( .A1(n15631), .A2(n16247), .ZN(n15485) );
  AOI211_X1 U18694 ( .C1(n16255), .C2(n15487), .A(n15486), .B(n15485), .ZN(
        n15492) );
  OR2_X1 U18695 ( .A1(n15489), .A2(n15488), .ZN(n15634) );
  NAND3_X1 U18696 ( .A1(n15634), .A2(n15490), .A3(n19121), .ZN(n15491) );
  OAI211_X1 U18697 ( .C1(n15627), .C2(n16256), .A(n15492), .B(n15491), .ZN(
        P2_U2991) );
  NAND2_X1 U18698 ( .A1(n15494), .A2(n15493), .ZN(n15496) );
  XOR2_X1 U18699 ( .A(n15496), .B(n15495), .Z(n15649) );
  NAND2_X1 U18700 ( .A1(n10853), .A2(n15640), .ZN(n15639) );
  NAND3_X1 U18701 ( .A1(n15481), .A2(n19118), .A3(n15639), .ZN(n15501) );
  INV_X1 U18702 ( .A(n15896), .ZN(n15499) );
  NOR2_X1 U18703 ( .A1(n15534), .A2(n19765), .ZN(n15642) );
  AOI21_X1 U18704 ( .B1(n19114), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15642), .ZN(n15497) );
  OAI21_X1 U18705 ( .B1(n19125), .B2(n15890), .A(n15497), .ZN(n15498) );
  AOI21_X1 U18706 ( .B1(n15499), .B2(n19117), .A(n15498), .ZN(n15500) );
  OAI211_X1 U18707 ( .C1(n15649), .C2(n16258), .A(n15501), .B(n15500), .ZN(
        P2_U2992) );
  NAND2_X1 U18708 ( .A1(n15503), .A2(n15502), .ZN(n15504) );
  XNOR2_X1 U18709 ( .A(n15505), .B(n15504), .ZN(n15671) );
  OR2_X2 U18710 ( .A1(n15506), .A2(n15702), .ZN(n15544) );
  NOR2_X2 U18711 ( .A1(n15544), .A2(n15688), .ZN(n15532) );
  AND2_X1 U18712 ( .A1(n15532), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15521) );
  INV_X1 U18713 ( .A(n15521), .ZN(n15507) );
  AOI21_X1 U18714 ( .B1(n15508), .B2(n15507), .A(n10773), .ZN(n15669) );
  NOR2_X1 U18715 ( .A1(n15534), .A2(n15509), .ZN(n15664) );
  NOR2_X1 U18716 ( .A1(n19125), .A2(n15510), .ZN(n15511) );
  AOI211_X1 U18717 ( .C1(n19114), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15664), .B(n15511), .ZN(n15512) );
  OAI21_X1 U18718 ( .B1(n16247), .B2(n18899), .A(n15512), .ZN(n15513) );
  AOI21_X1 U18719 ( .B1(n15669), .B2(n19118), .A(n15513), .ZN(n15514) );
  OAI21_X1 U18720 ( .B1(n15671), .B2(n16258), .A(n15514), .ZN(P2_U2994) );
  NAND2_X1 U18721 ( .A1(n15515), .A2(n15528), .ZN(n15519) );
  NAND2_X1 U18722 ( .A1(n15517), .A2(n15516), .ZN(n15518) );
  XNOR2_X1 U18723 ( .A(n15519), .B(n15518), .ZN(n15682) );
  NOR2_X1 U18724 ( .A1(n15532), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15520) );
  NAND2_X1 U18725 ( .A1(n15522), .A2(n16255), .ZN(n15524) );
  NOR2_X1 U18726 ( .A1(n15534), .A2(n19760), .ZN(n15672) );
  AOI21_X1 U18727 ( .B1(n19114), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15672), .ZN(n15523) );
  OAI211_X1 U18728 ( .C1(n15674), .C2(n16247), .A(n15524), .B(n15523), .ZN(
        n15525) );
  AOI21_X1 U18729 ( .B1(n10140), .B2(n19118), .A(n15525), .ZN(n15526) );
  OAI21_X1 U18730 ( .B1(n15682), .B2(n16258), .A(n15526), .ZN(P2_U2995) );
  NAND2_X1 U18731 ( .A1(n15528), .A2(n15527), .ZN(n15529) );
  XNOR2_X1 U18732 ( .A(n15530), .B(n15529), .ZN(n15697) );
  AND2_X1 U18733 ( .A1(n15544), .A2(n15688), .ZN(n15531) );
  NOR2_X1 U18734 ( .A1(n15532), .A2(n15531), .ZN(n15695) );
  NOR2_X1 U18735 ( .A1(n15534), .A2(n15533), .ZN(n15687) );
  AOI21_X1 U18736 ( .B1(n19114), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15687), .ZN(n15536) );
  NAND2_X1 U18737 ( .A1(n18917), .A2(n19117), .ZN(n15535) );
  OAI211_X1 U18738 ( .C1(n19125), .C2(n18911), .A(n15536), .B(n15535), .ZN(
        n15537) );
  AOI21_X1 U18739 ( .B1(n15695), .B2(n19118), .A(n15537), .ZN(n15538) );
  OAI21_X1 U18740 ( .B1(n15697), .B2(n16258), .A(n15538), .ZN(P2_U2996) );
  XOR2_X1 U18741 ( .A(n15540), .B(n15539), .Z(n15710) );
  NAND2_X1 U18742 ( .A1(n18923), .A2(n16255), .ZN(n15541) );
  NAND2_X1 U18743 ( .A1(n19113), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15699) );
  OAI211_X1 U18744 ( .C1(n16265), .C2(n15542), .A(n15541), .B(n15699), .ZN(
        n15543) );
  AOI21_X1 U18745 ( .B1(n19117), .B2(n18929), .A(n15543), .ZN(n15547) );
  INV_X1 U18746 ( .A(n15506), .ZN(n15545) );
  OAI211_X1 U18747 ( .C1(n15545), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n19118), .B(n15544), .ZN(n15546) );
  OAI211_X1 U18748 ( .C1(n15710), .C2(n16258), .A(n15547), .B(n15546), .ZN(
        P2_U2997) );
  OAI21_X1 U18749 ( .B1(n15550), .B2(n15549), .A(n15548), .ZN(n15725) );
  OR2_X1 U18750 ( .A1(n15725), .A2(n16258), .ZN(n15559) );
  NOR2_X1 U18751 ( .A1(n11229), .A2(n15534), .ZN(n15551) );
  AOI21_X1 U18752 ( .B1(n19117), .B2(n18939), .A(n15551), .ZN(n15558) );
  OAI21_X1 U18753 ( .B1(n15552), .B2(n10667), .A(n15713), .ZN(n15553) );
  NAND3_X1 U18754 ( .A1(n15553), .A2(n19118), .A3(n15506), .ZN(n15557) );
  INV_X1 U18755 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15554) );
  OAI22_X1 U18756 ( .A1(n16265), .A2(n15554), .B1(n19125), .B2(n18934), .ZN(
        n15555) );
  INV_X1 U18757 ( .A(n15555), .ZN(n15556) );
  NAND4_X1 U18758 ( .A1(n15559), .A2(n15558), .A3(n15557), .A4(n15556), .ZN(
        P2_U2998) );
  NAND2_X1 U18759 ( .A1(n15561), .A2(n15560), .ZN(n15565) );
  INV_X1 U18760 ( .A(n15728), .ZN(n15562) );
  NOR2_X1 U18761 ( .A1(n15563), .A2(n15562), .ZN(n15564) );
  XOR2_X1 U18762 ( .A(n15565), .B(n15564), .Z(n16275) );
  XNOR2_X1 U18763 ( .A(n15552), .B(n10667), .ZN(n16269) );
  AOI22_X1 U18764 ( .A1(n19114), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n16255), .B2(n15566), .ZN(n15568) );
  AOI22_X1 U18765 ( .A1(n19117), .A2(n16270), .B1(P2_REIP_REG_15__SCAN_IN), 
        .B2(n19113), .ZN(n15567) );
  OAI211_X1 U18766 ( .C1(n16269), .C2(n16256), .A(n15568), .B(n15567), .ZN(
        n15569) );
  INV_X1 U18767 ( .A(n15569), .ZN(n15570) );
  OAI21_X1 U18768 ( .B1(n16275), .B2(n16258), .A(n15570), .ZN(P2_U2999) );
  NAND2_X1 U18769 ( .A1(n15571), .A2(n16271), .ZN(n15589) );
  INV_X1 U18770 ( .A(n15573), .ZN(n15574) );
  NAND2_X1 U18771 ( .A1(n15574), .A2(n16302), .ZN(n15576) );
  OAI211_X1 U18772 ( .C1(n15577), .C2(n19143), .A(n15576), .B(n15575), .ZN(
        n15578) );
  INV_X1 U18773 ( .A(n15578), .ZN(n15586) );
  INV_X1 U18774 ( .A(n15579), .ZN(n15580) );
  AOI211_X1 U18775 ( .C1(n15583), .C2(n15582), .A(n15581), .B(n15580), .ZN(
        n15584) );
  INV_X1 U18776 ( .A(n15584), .ZN(n15585) );
  INV_X1 U18777 ( .A(n15587), .ZN(n15588) );
  OAI211_X1 U18778 ( .C1(n15590), .C2(n19133), .A(n15589), .B(n15588), .ZN(
        P2_U3017) );
  INV_X1 U18779 ( .A(n15591), .ZN(n15612) );
  NAND2_X1 U18780 ( .A1(n15592), .A2(n16298), .ZN(n15593) );
  OAI211_X1 U18781 ( .C1(n15595), .C2(n19138), .A(n15594), .B(n15593), .ZN(
        n15598) );
  XNOR2_X1 U18782 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15596) );
  NOR2_X1 U18783 ( .A1(n15610), .A2(n15596), .ZN(n15597) );
  AOI211_X1 U18784 ( .C1(n15612), .C2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15598), .B(n15597), .ZN(n15601) );
  NAND2_X1 U18785 ( .A1(n15599), .A2(n16300), .ZN(n15600) );
  OAI211_X1 U18786 ( .C1(n15602), .C2(n19137), .A(n15601), .B(n15600), .ZN(
        P2_U3020) );
  NAND3_X1 U18787 ( .A1(n15604), .A2(n16271), .A3(n15603), .ZN(n15614) );
  OAI21_X1 U18788 ( .B1(n19143), .B2(n15606), .A(n15605), .ZN(n15607) );
  AOI21_X1 U18789 ( .B1(n15608), .B2(n16302), .A(n15607), .ZN(n15609) );
  OAI21_X1 U18790 ( .B1(n15610), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15609), .ZN(n15611) );
  AOI21_X1 U18791 ( .B1(n15612), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15611), .ZN(n15613) );
  OAI211_X1 U18792 ( .C1(n15615), .C2(n19133), .A(n15614), .B(n15613), .ZN(
        P2_U3021) );
  INV_X1 U18793 ( .A(n15616), .ZN(n15617) );
  AOI21_X1 U18794 ( .B1(n15619), .B2(n15618), .A(n15617), .ZN(n15623) );
  NAND2_X1 U18795 ( .A1(n16160), .A2(n16302), .ZN(n15621) );
  OAI211_X1 U18796 ( .C1(n19143), .C2(n16158), .A(n15621), .B(n15620), .ZN(
        n15622) );
  AOI211_X1 U18797 ( .C1(n15624), .C2(n16300), .A(n15623), .B(n15622), .ZN(
        n15625) );
  OAI21_X1 U18798 ( .B1(n15626), .B2(n19137), .A(n15625), .ZN(P2_U3022) );
  OR2_X1 U18799 ( .A1(n15627), .A2(n19137), .ZN(n15638) );
  XNOR2_X1 U18800 ( .A(n15640), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15633) );
  INV_X1 U18801 ( .A(n15628), .ZN(n15629) );
  AOI21_X1 U18802 ( .B1(n16298), .B2(n9658), .A(n15629), .ZN(n15630) );
  OAI21_X1 U18803 ( .B1(n15631), .B2(n19138), .A(n15630), .ZN(n15632) );
  AOI21_X1 U18804 ( .B1(n15641), .B2(n15633), .A(n15632), .ZN(n15637) );
  NAND3_X1 U18805 ( .A1(n15634), .A2(n15490), .A3(n16300), .ZN(n15636) );
  NAND2_X1 U18806 ( .A1(n15646), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15635) );
  NAND4_X1 U18807 ( .A1(n15638), .A2(n15637), .A3(n15636), .A4(n15635), .ZN(
        P2_U3023) );
  NAND3_X1 U18808 ( .A1(n15481), .A2(n16271), .A3(n15639), .ZN(n15648) );
  NAND2_X1 U18809 ( .A1(n15641), .A2(n15640), .ZN(n15644) );
  AOI21_X1 U18810 ( .B1(n16298), .B2(n15894), .A(n15642), .ZN(n15643) );
  OAI211_X1 U18811 ( .C1(n15896), .C2(n19138), .A(n15644), .B(n15643), .ZN(
        n15645) );
  AOI21_X1 U18812 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15646), .A(
        n15645), .ZN(n15647) );
  OAI211_X1 U18813 ( .C1(n15649), .C2(n19133), .A(n15648), .B(n15647), .ZN(
        P2_U3024) );
  NAND2_X1 U18814 ( .A1(n15650), .A2(n16300), .ZN(n15659) );
  INV_X1 U18815 ( .A(n15651), .ZN(n15657) );
  NAND2_X1 U18816 ( .A1(n16298), .A2(n18893), .ZN(n15652) );
  OAI211_X1 U18817 ( .C1(n18892), .C2(n19138), .A(n15653), .B(n15652), .ZN(
        n15656) );
  NOR2_X1 U18818 ( .A1(n15654), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15655) );
  AOI211_X1 U18819 ( .C1(n15657), .C2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15656), .B(n15655), .ZN(n15658) );
  OAI211_X1 U18820 ( .C1(n15660), .C2(n19137), .A(n15659), .B(n15658), .ZN(
        P2_U3025) );
  XNOR2_X1 U18821 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15667) );
  NAND2_X1 U18822 ( .A1(n15679), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15666) );
  OR2_X1 U18823 ( .A1(n15268), .A2(n15661), .ZN(n15662) );
  AND2_X1 U18824 ( .A1(n15401), .A2(n15662), .ZN(n18897) );
  NOR2_X1 U18825 ( .A1(n18899), .A2(n19138), .ZN(n15663) );
  AOI211_X1 U18826 ( .C1(n16298), .C2(n18897), .A(n15664), .B(n15663), .ZN(
        n15665) );
  OAI211_X1 U18827 ( .C1(n15677), .C2(n15667), .A(n15666), .B(n15665), .ZN(
        n15668) );
  AOI21_X1 U18828 ( .B1(n15669), .B2(n16271), .A(n15668), .ZN(n15670) );
  OAI21_X1 U18829 ( .B1(n15671), .B2(n19133), .A(n15670), .ZN(P2_U3026) );
  AOI21_X1 U18830 ( .B1(n16298), .B2(n15673), .A(n15672), .ZN(n15676) );
  OR2_X1 U18831 ( .A1(n15674), .A2(n19138), .ZN(n15675) );
  OAI211_X1 U18832 ( .C1(n15677), .C2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15676), .B(n15675), .ZN(n15678) );
  AOI21_X1 U18833 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15679), .A(
        n15678), .ZN(n15681) );
  NAND2_X1 U18834 ( .A1(n10140), .A2(n16271), .ZN(n15680) );
  OAI211_X1 U18835 ( .C1(n15682), .C2(n19133), .A(n15681), .B(n15680), .ZN(
        P2_U3027) );
  NAND2_X1 U18836 ( .A1(n15683), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15693) );
  AND2_X1 U18837 ( .A1(n15685), .A2(n15684), .ZN(n15686) );
  NOR2_X1 U18838 ( .A1(n15269), .A2(n15686), .ZN(n18916) );
  AOI21_X1 U18839 ( .B1(n16298), .B2(n18916), .A(n15687), .ZN(n15692) );
  NAND3_X1 U18840 ( .A1(n16268), .A2(n15689), .A3(n15688), .ZN(n15691) );
  NAND2_X1 U18841 ( .A1(n16302), .A2(n18917), .ZN(n15690) );
  NAND4_X1 U18842 ( .A1(n15693), .A2(n15692), .A3(n15691), .A4(n15690), .ZN(
        n15694) );
  AOI21_X1 U18843 ( .B1(n15695), .B2(n16271), .A(n15694), .ZN(n15696) );
  OAI21_X1 U18844 ( .B1(n15697), .B2(n19133), .A(n15696), .ZN(P2_U3028) );
  INV_X1 U18845 ( .A(n16268), .ZN(n15712) );
  OAI22_X1 U18846 ( .A1(n15506), .A2(n19137), .B1(n15698), .B2(n15712), .ZN(
        n15703) );
  NAND2_X1 U18847 ( .A1(n16302), .A2(n18929), .ZN(n15700) );
  OAI211_X1 U18848 ( .C1(n19143), .C2(n18927), .A(n15700), .B(n15699), .ZN(
        n15701) );
  AOI21_X1 U18849 ( .B1(n15703), .B2(n15702), .A(n15701), .ZN(n15709) );
  NAND2_X1 U18850 ( .A1(n19147), .A2(n19137), .ZN(n15706) );
  NOR2_X1 U18851 ( .A1(n19128), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15704) );
  OR2_X1 U18852 ( .A1(n16267), .A2(n15704), .ZN(n15705) );
  AOI21_X1 U18853 ( .B1(n15506), .B2(n15706), .A(n15705), .ZN(n15711) );
  OAI21_X1 U18854 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15766), .A(
        n15711), .ZN(n15707) );
  NAND2_X1 U18855 ( .A1(n15707), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15708) );
  OAI211_X1 U18856 ( .C1(n15710), .C2(n19133), .A(n15709), .B(n15708), .ZN(
        P2_U3029) );
  INV_X1 U18857 ( .A(n15711), .ZN(n15723) );
  OAI21_X1 U18858 ( .B1(n15552), .B2(n19137), .A(n15712), .ZN(n15714) );
  NAND3_X1 U18859 ( .A1(n15714), .A2(n15713), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15721) );
  OR2_X1 U18860 ( .A1(n15716), .A2(n15715), .ZN(n15717) );
  AND2_X1 U18861 ( .A1(n15718), .A2(n15717), .ZN(n19012) );
  AOI22_X1 U18862 ( .A1(n16298), .A2(n19012), .B1(P2_REIP_REG_16__SCAN_IN), 
        .B2(n19113), .ZN(n15720) );
  NAND2_X1 U18863 ( .A1(n16302), .A2(n18939), .ZN(n15719) );
  NAND3_X1 U18864 ( .A1(n15721), .A2(n15720), .A3(n15719), .ZN(n15722) );
  AOI21_X1 U18865 ( .B1(n15723), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15722), .ZN(n15724) );
  OAI21_X1 U18866 ( .B1(n15725), .B2(n19133), .A(n15724), .ZN(P2_U3030) );
  OAI21_X1 U18867 ( .B1(n15726), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15552), .ZN(n16173) );
  NAND2_X1 U18868 ( .A1(n15728), .A2(n15727), .ZN(n15729) );
  XNOR2_X1 U18869 ( .A(n15730), .B(n15729), .ZN(n16175) );
  NAND2_X1 U18870 ( .A1(n16175), .A2(n16300), .ZN(n15741) );
  INV_X1 U18871 ( .A(n15731), .ZN(n15732) );
  NOR3_X1 U18872 ( .A1(n15732), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n16276), .ZN(n15739) );
  AOI21_X1 U18873 ( .B1(n15733), .B2(n14039), .A(n14240), .ZN(n18953) );
  INV_X1 U18874 ( .A(n18953), .ZN(n19020) );
  OAI22_X1 U18875 ( .A1(n19143), .A2(n19020), .B1(n19138), .B2(n18952), .ZN(
        n15738) );
  AND3_X1 U18876 ( .A1(n10644), .A2(n15734), .A3(n15789), .ZN(n15751) );
  OAI21_X1 U18877 ( .B1(n15734), .B2(n15766), .A(n15783), .ZN(n15752) );
  NOR2_X1 U18878 ( .A1(n15751), .A2(n15752), .ZN(n16277) );
  NAND3_X1 U18879 ( .A1(n15734), .A2(n15789), .A3(n16276), .ZN(n16286) );
  NAND2_X1 U18880 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19113), .ZN(n15735) );
  OAI221_X1 U18881 ( .B1(n15736), .B2(n16277), .C1(n15736), .C2(n16286), .A(
        n15735), .ZN(n15737) );
  AOI211_X1 U18882 ( .C1(n15789), .C2(n15739), .A(n15738), .B(n15737), .ZN(
        n15740) );
  OAI211_X1 U18883 ( .C1(n16173), .C2(n19137), .A(n15741), .B(n15740), .ZN(
        P2_U3032) );
  OR2_X1 U18884 ( .A1(n10085), .A2(n15743), .ZN(n15744) );
  XNOR2_X1 U18885 ( .A(n15745), .B(n15744), .ZN(n16190) );
  AND2_X1 U18886 ( .A1(n15747), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16208) );
  NAND2_X1 U18887 ( .A1(n16208), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16207) );
  OAI21_X1 U18888 ( .B1(n16207), .B2(n15767), .A(n10644), .ZN(n15749) );
  NAND2_X1 U18889 ( .A1(n15749), .A2(n15748), .ZN(n16194) );
  NOR2_X1 U18890 ( .A1(n11176), .A2(n15534), .ZN(n15750) );
  AOI211_X1 U18891 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n15752), .A(
        n15751), .B(n15750), .ZN(n15755) );
  OAI22_X1 U18892 ( .A1(n19025), .A2(n19143), .B1(n19138), .B2(n16191), .ZN(
        n15753) );
  INV_X1 U18893 ( .A(n15753), .ZN(n15754) );
  OAI211_X1 U18894 ( .C1(n16194), .C2(n19137), .A(n15755), .B(n15754), .ZN(
        n15756) );
  AOI21_X1 U18895 ( .B1(n16300), .B2(n16190), .A(n15756), .ZN(n15757) );
  INV_X1 U18896 ( .A(n15757), .ZN(P2_U3034) );
  XNOR2_X1 U18897 ( .A(n16207), .B(n15767), .ZN(n16201) );
  INV_X1 U18898 ( .A(n15758), .ZN(n15759) );
  NAND2_X1 U18899 ( .A1(n15760), .A2(n15759), .ZN(n15765) );
  INV_X1 U18900 ( .A(n15761), .ZN(n15762) );
  NOR2_X1 U18901 ( .A1(n15763), .A2(n15762), .ZN(n15764) );
  XNOR2_X1 U18902 ( .A(n15765), .B(n15764), .ZN(n16200) );
  OAI21_X1 U18903 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15766), .A(
        n15783), .ZN(n16290) );
  NOR2_X1 U18904 ( .A1(n10812), .A2(n15534), .ZN(n15770) );
  NAND2_X1 U18905 ( .A1(n15789), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16287) );
  AOI221_X1 U18906 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C1(n15768), .C2(n15767), .A(
        n16287), .ZN(n15769) );
  AOI211_X1 U18907 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16290), .A(
        n15770), .B(n15769), .ZN(n15774) );
  OAI22_X1 U18908 ( .A1(n19027), .A2(n19143), .B1(n19138), .B2(n15771), .ZN(
        n15772) );
  INV_X1 U18909 ( .A(n15772), .ZN(n15773) );
  OAI211_X1 U18910 ( .C1(n16200), .C2(n19133), .A(n15774), .B(n15773), .ZN(
        n15775) );
  INV_X1 U18911 ( .A(n15775), .ZN(n15776) );
  OAI21_X1 U18912 ( .B1(n16201), .B2(n19137), .A(n15776), .ZN(P2_U3035) );
  INV_X1 U18913 ( .A(n16208), .ZN(n15777) );
  OAI21_X1 U18914 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15747), .A(
        n15777), .ZN(n16222) );
  NOR2_X1 U18915 ( .A1(n11130), .A2(n15534), .ZN(n15781) );
  OR2_X1 U18916 ( .A1(n15778), .A2(n13868), .ZN(n15779) );
  NAND2_X1 U18917 ( .A1(n15779), .A2(n13880), .ZN(n19032) );
  NOR2_X1 U18918 ( .A1(n19143), .A2(n19032), .ZN(n15780) );
  AOI211_X1 U18919 ( .C1(n16224), .C2(n16302), .A(n15781), .B(n15780), .ZN(
        n15782) );
  OAI21_X1 U18920 ( .B1(n15783), .B2(n15788), .A(n15782), .ZN(n15787) );
  NAND2_X1 U18921 ( .A1(n9692), .A2(n16209), .ZN(n15785) );
  XNOR2_X1 U18922 ( .A(n15784), .B(n15785), .ZN(n16221) );
  NOR2_X1 U18923 ( .A1(n16221), .A2(n19133), .ZN(n15786) );
  AOI211_X1 U18924 ( .C1(n15789), .C2(n15788), .A(n15787), .B(n15786), .ZN(
        n15790) );
  OAI21_X1 U18925 ( .B1(n16222), .B2(n19137), .A(n15790), .ZN(P2_U3037) );
  OAI22_X1 U18926 ( .A1(n15792), .A2(n19138), .B1(n19137), .B2(n15791), .ZN(
        n15793) );
  AOI211_X1 U18927 ( .C1(n19130), .C2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n15794), .B(n15793), .ZN(n15800) );
  AOI22_X1 U18928 ( .A1(n16300), .A2(n15795), .B1(n16298), .B2(n19820), .ZN(
        n15799) );
  OAI211_X1 U18929 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n15797), .B(n15796), .ZN(n15798) );
  NAND3_X1 U18930 ( .A1(n15800), .A2(n15799), .A3(n15798), .ZN(P2_U3045) );
  OR2_X1 U18931 ( .A1(n13541), .A2(n15801), .ZN(n15816) );
  NAND2_X1 U18932 ( .A1(n15803), .A2(n15802), .ZN(n15806) );
  NAND3_X1 U18933 ( .A1(n15806), .A2(n15805), .A3(n15804), .ZN(n15813) );
  INV_X1 U18934 ( .A(n11048), .ZN(n15808) );
  OAI22_X1 U18935 ( .A1(n15810), .A2(n15809), .B1(n15808), .B2(n15807), .ZN(
        n15812) );
  MUX2_X1 U18936 ( .A(n15813), .B(n15812), .S(n15811), .Z(n15814) );
  NOR2_X1 U18937 ( .A1(n15814), .A2(n10445), .ZN(n15815) );
  NAND2_X1 U18938 ( .A1(n15816), .A2(n15815), .ZN(n16323) );
  INV_X1 U18939 ( .A(n16323), .ZN(n15817) );
  OAI22_X1 U18940 ( .A1(n19795), .A2(n16359), .B1(n15857), .B2(n15817), .ZN(
        n15819) );
  MUX2_X1 U18941 ( .A(n15819), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15818), .Z(P2_U3596) );
  INV_X1 U18942 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16624) );
  INV_X1 U18943 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16950) );
  NOR2_X1 U18944 ( .A1(n18225), .A2(n16995), .ZN(n16980) );
  NAND2_X1 U18945 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16980), .ZN(n16968) );
  NAND2_X1 U18946 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n9636), .ZN(n16938) );
  XOR2_X1 U18947 ( .A(n16929), .B(n16935), .Z(n17219) );
  AOI22_X1 U18948 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16932), .B1(n17198), 
        .B2(n17219), .ZN(n15822) );
  OAI21_X1 U18949 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n16938), .A(n15822), .ZN(
        P3_U2675) );
  AOI22_X1 U18950 ( .A1(n12689), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15827) );
  AOI22_X1 U18951 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12692), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15826) );
  AOI22_X1 U18952 ( .A1(n15823), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15825) );
  AOI22_X1 U18953 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15824) );
  NAND4_X1 U18954 ( .A1(n15827), .A2(n15826), .A3(n15825), .A4(n15824), .ZN(
        n15834) );
  AOI22_X1 U18955 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12703), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15832) );
  AOI22_X1 U18956 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15831) );
  AOI22_X1 U18957 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n15828), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15830) );
  AOI22_X1 U18958 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15829) );
  NAND4_X1 U18959 ( .A1(n15832), .A2(n15831), .A3(n15830), .A4(n15829), .ZN(
        n15833) );
  NOR2_X1 U18960 ( .A1(n15834), .A2(n15833), .ZN(n17298) );
  AND2_X1 U18961 ( .A1(n16928), .A2(n17080), .ZN(n17077) );
  NAND2_X1 U18962 ( .A1(n17192), .A2(n15835), .ZN(n17091) );
  NOR2_X1 U18963 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17091), .ZN(n15836) );
  AOI211_X1 U18964 ( .C1(n17298), .C2(n17198), .A(n17077), .B(n15836), .ZN(
        P3_U2690) );
  NOR2_X1 U18965 ( .A1(n15851), .A2(n18801), .ZN(n18696) );
  NAND2_X1 U18966 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18696), .ZN(n18792) );
  INV_X1 U18967 ( .A(n18792), .ZN(n18699) );
  NAND3_X1 U18968 ( .A1(n9635), .A2(n15855), .A3(n18631), .ZN(n18174) );
  AOI221_X1 U18969 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n18699), .C1(n18174), .C2(
        n18699), .A(n18535), .ZN(n18178) );
  INV_X1 U18970 ( .A(n18178), .ZN(n18182) );
  NAND2_X1 U18971 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18637), .ZN(n18229) );
  NAND2_X1 U18972 ( .A1(n18182), .A2(n18229), .ZN(n15840) );
  NOR2_X1 U18973 ( .A1(n18638), .A2(n15840), .ZN(n15842) );
  INV_X1 U18974 ( .A(n15840), .ZN(n15838) );
  NAND2_X1 U18975 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17744) );
  AOI21_X1 U18976 ( .B1(n18173), .B2(n17744), .A(P3_STATE2_REG_3__SCAN_IN), 
        .ZN(n15837) );
  INV_X1 U18977 ( .A(n15837), .ZN(n15841) );
  AOI21_X1 U18978 ( .B1(n15838), .B2(n15841), .A(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15839) );
  AOI21_X1 U18979 ( .B1(n15842), .B2(n18532), .A(n15839), .ZN(P3_U2864) );
  NAND2_X1 U18980 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18352) );
  OAI22_X1 U18981 ( .A1(n18178), .A2(n15841), .B1(n15840), .B2(n18352), .ZN(
        n18179) );
  INV_X1 U18982 ( .A(n18532), .ZN(n18475) );
  AOI22_X1 U18983 ( .A1(n18475), .A2(n18182), .B1(n15842), .B2(n15841), .ZN(
        n18181) );
  AOI22_X1 U18984 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18179), .B1(
        n18181), .B2(n18670), .ZN(P3_U2865) );
  INV_X1 U18985 ( .A(n15843), .ZN(n15845) );
  AOI211_X1 U18986 ( .C1(n16537), .C2(n15846), .A(n15845), .B(n15844), .ZN(
        n15867) );
  INV_X1 U18987 ( .A(n18843), .ZN(n18836) );
  NOR2_X1 U18988 ( .A1(n18622), .A2(n18836), .ZN(n15849) );
  NAND2_X1 U18989 ( .A1(n18842), .A2(n17416), .ZN(n18681) );
  INV_X1 U18990 ( .A(n15863), .ZN(n18840) );
  AOI22_X1 U18991 ( .A1(n18627), .A2(n15848), .B1(n15849), .B2(n17352), .ZN(
        n15850) );
  NAND3_X1 U18992 ( .A1(n15867), .A2(n15850), .A3(n15963), .ZN(n18664) );
  INV_X1 U18993 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18175) );
  NAND2_X1 U18994 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n15851), .ZN(n18183) );
  OAI21_X1 U18995 ( .B1(n18175), .B2(n18792), .A(n18183), .ZN(n15852) );
  AOI21_X1 U18996 ( .B1(n18679), .B2(n18664), .A(n15852), .ZN(n18822) );
  INV_X1 U18997 ( .A(n18822), .ZN(n18819) );
  INV_X1 U18998 ( .A(n15853), .ZN(n15854) );
  AOI21_X1 U18999 ( .B1(n15855), .B2(n18631), .A(n15854), .ZN(n18677) );
  NAND3_X1 U19000 ( .A1(n18819), .A2(n18817), .A3(n18677), .ZN(n15856) );
  OAI21_X1 U19001 ( .B1(n18819), .B2(n18631), .A(n15856), .ZN(P3_U3284) );
  NOR4_X1 U19002 ( .A1(n10966), .A2(n16343), .A3(n15857), .A4(n13297), .ZN(
        n15858) );
  NAND2_X1 U19003 ( .A1(n15861), .A2(n15858), .ZN(n15859) );
  OAI21_X1 U19004 ( .B1(n15861), .B2(n15860), .A(n15859), .ZN(P2_U3595) );
  NAND2_X1 U19005 ( .A1(n15862), .A2(n18215), .ZN(n15868) );
  AOI21_X1 U19006 ( .B1(n18842), .B2(n18200), .A(n15863), .ZN(n15864) );
  AOI21_X1 U19007 ( .B1(n15864), .B2(n15872), .A(n18836), .ZN(n16536) );
  OAI211_X1 U19008 ( .C1(n17209), .C2(n18200), .A(n16536), .B(n15865), .ZN(
        n15866) );
  OAI211_X1 U19009 ( .C1(n15869), .C2(n15868), .A(n15867), .B(n15866), .ZN(
        n15871) );
  NOR2_X1 U19010 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17743), .ZN(
        n16426) );
  INV_X1 U19011 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17861) );
  NOR2_X1 U19012 ( .A1(n18658), .A2(n18654), .ZN(n18027) );
  INV_X1 U19013 ( .A(n18027), .ZN(n18059) );
  INV_X2 U19014 ( .A(n18122), .ZN(n18165) );
  NOR3_X1 U19015 ( .A1(n18118), .A2(n10066), .A3(n17786), .ZN(n17966) );
  AOI21_X1 U19016 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18115) );
  INV_X1 U19017 ( .A(n18115), .ZN(n15875) );
  NAND2_X1 U19018 ( .A1(n17966), .A2(n15875), .ZN(n18079) );
  NAND2_X1 U19019 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18076) );
  OR2_X1 U19020 ( .A1(n20851), .A2(n18076), .ZN(n17967) );
  NOR2_X1 U19021 ( .A1(n18079), .A2(n17967), .ZN(n18020) );
  NAND3_X1 U19022 ( .A1(n17963), .A2(n17850), .A3(n18020), .ZN(n17959) );
  NAND2_X1 U19023 ( .A1(n17878), .A2(n17849), .ZN(n15881) );
  OAI21_X1 U19024 ( .B1(n17959), .B2(n15881), .A(n18654), .ZN(n17855) );
  NAND2_X1 U19025 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17965) );
  INV_X1 U19026 ( .A(n17965), .ZN(n18116) );
  NAND2_X1 U19027 ( .A1(n17966), .A2(n18116), .ZN(n18077) );
  NOR2_X1 U19028 ( .A1(n17967), .A2(n18077), .ZN(n18021) );
  NAND2_X1 U19029 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18021), .ZN(
        n18065) );
  NOR2_X1 U19030 ( .A1(n17969), .A2(n18065), .ZN(n17980) );
  NAND2_X1 U19031 ( .A1(n15876), .A2(n17980), .ZN(n17852) );
  NAND2_X1 U19032 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17849), .ZN(
        n16425) );
  OAI21_X1 U19033 ( .B1(n17852), .B2(n16425), .A(n18633), .ZN(n15878) );
  NAND3_X1 U19034 ( .A1(n17963), .A2(n17850), .A3(n18021), .ZN(n15882) );
  OAI21_X1 U19035 ( .B1(n15881), .B2(n15882), .A(n18658), .ZN(n15877) );
  NAND4_X1 U19036 ( .A1(n18119), .A2(n17855), .A3(n15878), .A4(n15877), .ZN(
        n15951) );
  AOI21_X1 U19037 ( .B1(n17861), .B2(n18059), .A(n15951), .ZN(n16433) );
  NAND2_X1 U19038 ( .A1(n17918), .A2(n18162), .ZN(n18171) );
  INV_X1 U19039 ( .A(n18623), .ZN(n16428) );
  NOR2_X1 U19040 ( .A1(n18154), .A2(n18045), .ZN(n18087) );
  AOI22_X1 U19041 ( .A1(n18152), .A2(n16393), .B1(n18087), .B2(n16391), .ZN(
        n15955) );
  NOR2_X1 U19042 ( .A1(n18154), .A2(n18120), .ZN(n18157) );
  NAND2_X1 U19043 ( .A1(n18157), .A2(n17476), .ZN(n15880) );
  OAI211_X1 U19044 ( .C1(n18153), .C2(n16433), .A(n15955), .B(n15880), .ZN(
        n15886) );
  INV_X1 U19045 ( .A(n15881), .ZN(n15883) );
  AOI21_X1 U19046 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18633), .A(
        n18658), .ZN(n18138) );
  OAI22_X1 U19047 ( .A1(n18648), .A2(n17959), .B1(n15882), .B2(n18138), .ZN(
        n17877) );
  NAND2_X1 U19048 ( .A1(n15883), .A2(n17877), .ZN(n16413) );
  OAI21_X1 U19049 ( .B1(n16430), .B2(n18626), .A(n16413), .ZN(n15884) );
  AOI22_X1 U19050 ( .A1(n17475), .A2(n18087), .B1(n18162), .B2(n15884), .ZN(
        n15954) );
  OAI21_X1 U19051 ( .B1(n16431), .B2(n15954), .A(n12799), .ZN(n15885) );
  OAI21_X1 U19052 ( .B1(n12799), .B2(n15886), .A(n15885), .ZN(n15887) );
  NAND2_X1 U19053 ( .A1(n18153), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16402) );
  OAI211_X1 U19054 ( .C1(n18091), .C2(n16404), .A(n15887), .B(n16402), .ZN(
        P3_U2833) );
  NOR2_X1 U19055 ( .A1(n9951), .A2(n15888), .ZN(n15889) );
  XOR2_X1 U19056 ( .A(n15890), .B(n15889), .Z(n15900) );
  OAI22_X1 U19057 ( .A1(n15891), .A2(n18995), .B1(n18974), .B2(n9937), .ZN(
        n15892) );
  INV_X1 U19058 ( .A(n15892), .ZN(n15893) );
  OAI21_X1 U19059 ( .B1(n19765), .B2(n18987), .A(n15893), .ZN(n15898) );
  INV_X1 U19060 ( .A(n15894), .ZN(n15895) );
  OAI22_X1 U19061 ( .A1(n15896), .A2(n18978), .B1(n18989), .B2(n15895), .ZN(
        n15897) );
  AOI211_X1 U19062 ( .C1(P2_EBX_REG_22__SCAN_IN), .C2(n18992), .A(n15898), .B(
        n15897), .ZN(n15899) );
  OAI21_X1 U19063 ( .B1(n19717), .B2(n15900), .A(n15899), .ZN(P2_U2833) );
  NAND2_X1 U19064 ( .A1(n15902), .A2(n15901), .ZN(n15908) );
  AOI21_X1 U19065 ( .B1(n15903), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n20499), .ZN(n15904) );
  OAI211_X1 U19066 ( .C1(n15908), .C2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15905), .B(n15904), .ZN(n15906) );
  INV_X1 U19067 ( .A(n15906), .ZN(n15907) );
  AOI21_X1 U19068 ( .B1(n15908), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15907), .ZN(n15909) );
  NAND2_X1 U19069 ( .A1(n11803), .A2(n15909), .ZN(n15911) );
  INV_X1 U19070 ( .A(n15909), .ZN(n15910) );
  AOI22_X1 U19071 ( .A1(n15912), .A2(n15911), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15910), .ZN(n15914) );
  OR2_X1 U19072 ( .A1(n15914), .A2(n15913), .ZN(n15915) );
  AOI22_X1 U19073 ( .A1(n15915), .A2(n20727), .B1(n15914), .B2(n15913), .ZN(
        n15924) );
  OAI21_X1 U19074 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15916), .ZN(n15917) );
  INV_X1 U19075 ( .A(n15917), .ZN(n15919) );
  NOR4_X1 U19076 ( .A1(n15921), .A2(n15920), .A3(n15919), .A4(n15918), .ZN(
        n15923) );
  OAI211_X1 U19077 ( .C1(n15924), .C2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n15923), .B(n15922), .ZN(n15931) );
  NAND3_X1 U19078 ( .A1(n15927), .A2(n15926), .A3(n15925), .ZN(n15930) );
  OAI21_X1 U19079 ( .B1(n15928), .B2(n20647), .A(n20634), .ZN(n15929) );
  NAND2_X1 U19080 ( .A1(n15930), .A2(n15929), .ZN(n16147) );
  AOI221_X1 U19081 ( .B1(n20744), .B2(n16149), .C1(n15931), .C2(n16149), .A(
        n16147), .ZN(n15933) );
  NOR2_X1 U19082 ( .A1(n15933), .A2(n20744), .ZN(n20635) );
  OAI211_X1 U19083 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20647), .A(n20635), 
        .B(n15935), .ZN(n16148) );
  AOI21_X1 U19084 ( .B1(n15932), .B2(n15931), .A(n16148), .ZN(n15939) );
  INV_X1 U19085 ( .A(n15933), .ZN(n15934) );
  OAI21_X1 U19086 ( .B1(n15936), .B2(n15935), .A(n15934), .ZN(n15937) );
  AOI22_X1 U19087 ( .A1(n15939), .A2(n15938), .B1(n20744), .B2(n15937), .ZN(
        P1_U3161) );
  AOI22_X1 U19088 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15940), .B1(
        n16118), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15948) );
  OAI22_X1 U19089 ( .A1(n15943), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n15942), .B2(n15941), .ZN(n15944) );
  XNOR2_X1 U19090 ( .A(n15944), .B(n11937), .ZN(n16017) );
  XNOR2_X1 U19091 ( .A(n15946), .B(n15945), .ZN(n16013) );
  AOI22_X1 U19092 ( .A1(n16017), .A2(n16122), .B1(n16119), .B2(n16013), .ZN(
        n15947) );
  OAI211_X1 U19093 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15949), .A(
        n15948), .B(n15947), .ZN(P1_U3010) );
  INV_X1 U19094 ( .A(n15950), .ZN(n16415) );
  AOI22_X1 U19095 ( .A1(n18157), .A2(n16415), .B1(n18122), .B2(n15951), .ZN(
        n16412) );
  INV_X1 U19096 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20653) );
  INV_X1 U19097 ( .A(HOLD), .ZN(n20639) );
  NOR2_X1 U19098 ( .A1(n20653), .A2(n20639), .ZN(n20642) );
  AOI22_X1 U19099 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15957) );
  NAND2_X1 U19100 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20741), .ZN(n20638) );
  OAI211_X1 U19101 ( .C1(n20642), .C2(n15957), .A(n15956), .B(n20638), .ZN(
        P1_U3195) );
  AND2_X1 U19102 ( .A1(n20016), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR3_X1 U19103 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15959) );
  NOR2_X1 U19104 ( .A1(n13325), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19715) );
  AND2_X1 U19105 ( .A1(n19849), .A2(n19715), .ZN(n16366) );
  NOR4_X1 U19106 ( .A1(n15959), .A2(n19850), .A3(n16366), .A4(n15958), .ZN(
        P2_U3178) );
  INV_X1 U19107 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n20817) );
  INV_X1 U19108 ( .A(n19834), .ZN(n15960) );
  OAI221_X1 U19109 ( .B1(n20817), .B2(n16375), .C1(n15960), .C2(n16375), .A(
        n19363), .ZN(n19826) );
  NOR2_X1 U19110 ( .A1(n16330), .A2(n19826), .ZN(P2_U3047) );
  NAND2_X1 U19111 ( .A1(n16928), .A2(n17202), .ZN(n17292) );
  INV_X1 U19112 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17414) );
  AOI22_X1 U19113 ( .A1(n17348), .A2(BUF2_REG_0__SCAN_IN), .B1(n17317), .B2(
        n17842), .ZN(n15964) );
  OAI221_X1 U19114 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17292), .C1(n17414), 
        .C2(n17202), .A(n15964), .ZN(P3_U2735) );
  INV_X1 U19115 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15965) );
  OAI22_X1 U19116 ( .A1(n19944), .A2(n16016), .B1(n15965), .B2(n19975), .ZN(
        n15966) );
  AOI211_X1 U19117 ( .C1(n15968), .C2(P1_REIP_REG_21__SCAN_IN), .A(n15967), 
        .B(n15966), .ZN(n15970) );
  AOI22_X1 U19118 ( .A1(n16018), .A2(n19899), .B1(n19971), .B2(n16013), .ZN(
        n15969) );
  OAI211_X1 U19119 ( .C1(n16021), .C2(n19983), .A(n15970), .B(n15969), .ZN(
        P1_U2819) );
  AOI22_X1 U19120 ( .A1(n15972), .A2(n19958), .B1(P1_REIP_REG_15__SCAN_IN), 
        .B2(n15971), .ZN(n15979) );
  AOI21_X1 U19121 ( .B1(n19959), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n19931), .ZN(n15974) );
  NAND2_X1 U19122 ( .A1(n9585), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n15973) );
  OAI211_X1 U19123 ( .C1(n16078), .C2(n19968), .A(n15974), .B(n15973), .ZN(
        n15975) );
  AOI211_X1 U19124 ( .C1(n15977), .C2(n19899), .A(n15976), .B(n15975), .ZN(
        n15978) );
  NAND2_X1 U19125 ( .A1(n15979), .A2(n15978), .ZN(P1_U2825) );
  OAI22_X1 U19126 ( .A1(n16085), .A2(n19968), .B1(n15980), .B2(n19944), .ZN(
        n15981) );
  AOI211_X1 U19127 ( .C1(n19959), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n19931), .B(n15981), .ZN(n15988) );
  NOR2_X1 U19128 ( .A1(n15982), .A2(n15998), .ZN(n15985) );
  INV_X1 U19129 ( .A(n15983), .ZN(n15984) );
  MUX2_X1 U19130 ( .A(n15985), .B(n15984), .S(P1_REIP_REG_13__SCAN_IN), .Z(
        n15986) );
  AOI21_X1 U19131 ( .B1(n16051), .B2(n19899), .A(n15986), .ZN(n15987) );
  OAI211_X1 U19132 ( .C1(n15989), .C2(n19983), .A(n15988), .B(n15987), .ZN(
        P1_U2827) );
  AOI22_X1 U19133 ( .A1(n16002), .A2(P1_REIP_REG_11__SCAN_IN), .B1(n9585), 
        .B2(P1_EBX_REG_11__SCAN_IN), .ZN(n15990) );
  OAI211_X1 U19134 ( .C1(n19975), .C2(n15991), .A(n15990), .B(n19918), .ZN(
        n15992) );
  AOI21_X1 U19135 ( .B1(n19971), .B2(n16112), .A(n15992), .ZN(n15997) );
  NOR2_X1 U19136 ( .A1(n19983), .A2(n15993), .ZN(n15994) );
  AOI21_X1 U19137 ( .B1(n15995), .B2(n19899), .A(n15994), .ZN(n15996) );
  OAI211_X1 U19138 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n15998), .A(n15997), 
        .B(n15996), .ZN(P1_U2829) );
  INV_X1 U19139 ( .A(n15999), .ZN(n16056) );
  AOI22_X1 U19140 ( .A1(n16056), .A2(n19899), .B1(n19958), .B2(n16054), .ZN(
        n16012) );
  NOR3_X1 U19141 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n16001), .A3(n16000), 
        .ZN(n16010) );
  NAND2_X1 U19142 ( .A1(n9585), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n16008) );
  INV_X1 U19143 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16005) );
  AOI22_X1 U19144 ( .A1(n19971), .A2(n16003), .B1(P1_REIP_REG_10__SCAN_IN), 
        .B2(n16002), .ZN(n16004) );
  OAI211_X1 U19145 ( .C1(n19975), .C2(n16005), .A(n16004), .B(n19918), .ZN(
        n16006) );
  INV_X1 U19146 ( .A(n16006), .ZN(n16007) );
  NAND2_X1 U19147 ( .A1(n16008), .A2(n16007), .ZN(n16009) );
  NOR2_X1 U19148 ( .A1(n16010), .A2(n16009), .ZN(n16011) );
  NAND2_X1 U19149 ( .A1(n16012), .A2(n16011), .ZN(P1_U2830) );
  AOI22_X1 U19150 ( .A1(n16018), .A2(n16014), .B1(n12508), .B2(n16013), .ZN(
        n16015) );
  OAI21_X1 U19151 ( .B1(n19997), .B2(n16016), .A(n16015), .ZN(P1_U2851) );
  AOI22_X1 U19152 ( .A1(n16060), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n16118), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n16020) );
  AOI22_X1 U19153 ( .A1(n16018), .A2(n16066), .B1(n16065), .B2(n16017), .ZN(
        n16019) );
  OAI211_X1 U19154 ( .C1(n16069), .C2(n16021), .A(n16020), .B(n16019), .ZN(
        P1_U2978) );
  AOI22_X1 U19155 ( .A1(n16060), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n16118), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16026) );
  OAI22_X1 U19156 ( .A1(n16023), .A2(n20055), .B1(n19869), .B2(n16022), .ZN(
        n16024) );
  INV_X1 U19157 ( .A(n16024), .ZN(n16025) );
  OAI211_X1 U19158 ( .C1(n16069), .C2(n16027), .A(n16026), .B(n16025), .ZN(
        P1_U2980) );
  AOI22_X1 U19159 ( .A1(n16060), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n16118), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n16031) );
  AOI22_X1 U19160 ( .A1(n16029), .A2(n16066), .B1(n16055), .B2(n16028), .ZN(
        n16030) );
  OAI211_X1 U19161 ( .C1(n19869), .C2(n16032), .A(n16031), .B(n16030), .ZN(
        P1_U2982) );
  INV_X1 U19162 ( .A(n16033), .ZN(n16034) );
  NOR2_X1 U19163 ( .A1(n16035), .A2(n16034), .ZN(n16039) );
  NAND2_X1 U19164 ( .A1(n16037), .A2(n16036), .ZN(n16038) );
  XNOR2_X1 U19165 ( .A(n16039), .B(n16038), .ZN(n16079) );
  AOI22_X1 U19166 ( .A1(n16060), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n16118), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16044) );
  OAI22_X1 U19167 ( .A1(n16041), .A2(n20055), .B1(n16040), .B2(n16069), .ZN(
        n16042) );
  INV_X1 U19168 ( .A(n16042), .ZN(n16043) );
  OAI211_X1 U19169 ( .C1(n16079), .C2(n19869), .A(n16044), .B(n16043), .ZN(
        P1_U2984) );
  AOI21_X1 U19170 ( .B1(n16047), .B2(n16046), .A(n16045), .ZN(n16048) );
  XOR2_X1 U19171 ( .A(n16049), .B(n16048), .Z(n16086) );
  AOI22_X1 U19172 ( .A1(n16060), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n16118), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n16053) );
  AOI22_X1 U19173 ( .A1(n16051), .A2(n16066), .B1(n16050), .B2(n16055), .ZN(
        n16052) );
  OAI211_X1 U19174 ( .C1(n19869), .C2(n16086), .A(n16053), .B(n16052), .ZN(
        P1_U2986) );
  AOI22_X1 U19175 ( .A1(n16060), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n16118), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n16058) );
  AOI22_X1 U19176 ( .A1(n16056), .A2(n16066), .B1(n16055), .B2(n16054), .ZN(
        n16057) );
  OAI211_X1 U19177 ( .C1(n19869), .C2(n16059), .A(n16058), .B(n16057), .ZN(
        P1_U2989) );
  AOI22_X1 U19178 ( .A1(n16060), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16118), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16068) );
  NAND2_X1 U19179 ( .A1(n16063), .A2(n16062), .ZN(n16064) );
  XNOR2_X1 U19180 ( .A(n16061), .B(n16064), .ZN(n16123) );
  AOI22_X1 U19181 ( .A1(n19900), .A2(n16066), .B1(n16065), .B2(n16123), .ZN(
        n16067) );
  OAI211_X1 U19182 ( .C1(n16069), .C2(n19902), .A(n16068), .B(n16067), .ZN(
        P1_U2992) );
  OAI21_X1 U19183 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n16070), .ZN(n16077) );
  OAI21_X1 U19184 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16071), .A(
        n16091), .ZN(n16082) );
  AOI22_X1 U19185 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n16082), .B1(
        n16118), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16076) );
  INV_X1 U19186 ( .A(n16072), .ZN(n16074) );
  AOI22_X1 U19187 ( .A1(n16074), .A2(n16122), .B1(n16119), .B2(n16073), .ZN(
        n16075) );
  OAI211_X1 U19188 ( .C1(n16084), .C2(n16077), .A(n16076), .B(n16075), .ZN(
        P1_U3015) );
  NOR2_X1 U19189 ( .A1(n16134), .A2(n20670), .ZN(n16081) );
  OAI22_X1 U19190 ( .A1(n16079), .A2(n16137), .B1(n16136), .B2(n16078), .ZN(
        n16080) );
  AOI211_X1 U19191 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16082), .A(
        n16081), .B(n16080), .ZN(n16083) );
  OAI21_X1 U19192 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16084), .A(
        n16083), .ZN(P1_U3016) );
  OAI22_X1 U19193 ( .A1(n16086), .A2(n16137), .B1(n16136), .B2(n16085), .ZN(
        n16087) );
  AOI21_X1 U19194 ( .B1(n16118), .B2(P1_REIP_REG_13__SCAN_IN), .A(n16087), 
        .ZN(n16088) );
  OAI221_X1 U19195 ( .B1(n16091), .B2(n16090), .C1(n16091), .C2(n16089), .A(
        n16088), .ZN(P1_U3018) );
  NOR2_X1 U19196 ( .A1(n16094), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16110) );
  INV_X1 U19197 ( .A(n16092), .ZN(n16093) );
  OAI21_X1 U19198 ( .B1(n16095), .B2(n16094), .A(n16093), .ZN(n16096) );
  OAI211_X1 U19199 ( .C1(n16105), .C2(n16098), .A(n16097), .B(n16096), .ZN(
        n16113) );
  AOI21_X1 U19200 ( .B1(n16099), .B2(n16110), .A(n16113), .ZN(n16109) );
  INV_X1 U19201 ( .A(n16100), .ZN(n16102) );
  AOI21_X1 U19202 ( .B1(n16102), .B2(n16119), .A(n16101), .ZN(n16108) );
  INV_X1 U19203 ( .A(n16103), .ZN(n16106) );
  NOR2_X1 U19204 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16127), .ZN(
        n16104) );
  AOI22_X1 U19205 ( .A1(n16106), .A2(n16122), .B1(n16105), .B2(n16104), .ZN(
        n16107) );
  OAI211_X1 U19206 ( .C1(n16109), .C2(n11762), .A(n16108), .B(n16107), .ZN(
        P1_U3019) );
  INV_X1 U19207 ( .A(n16110), .ZN(n16117) );
  AOI21_X1 U19208 ( .B1(n16112), .B2(n16119), .A(n16111), .ZN(n16116) );
  AOI22_X1 U19209 ( .A1(n16114), .A2(n16122), .B1(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16113), .ZN(n16115) );
  OAI211_X1 U19210 ( .C1(n16127), .C2(n16117), .A(n16116), .B(n16115), .ZN(
        P1_U3020) );
  OR2_X1 U19211 ( .A1(n16142), .A2(n16127), .ZN(n16126) );
  INV_X1 U19212 ( .A(n19896), .ZN(n16120) );
  AOI22_X1 U19213 ( .A1(n16120), .A2(n16119), .B1(n16118), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16125) );
  AOI22_X1 U19214 ( .A1(n16123), .A2(n16122), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16121), .ZN(n16124) );
  OAI211_X1 U19215 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n16126), .A(
        n16125), .B(n16124), .ZN(P1_U3024) );
  INV_X1 U19216 ( .A(n16127), .ZN(n16141) );
  INV_X1 U19217 ( .A(n16128), .ZN(n16131) );
  AOI21_X1 U19218 ( .B1(n16131), .B2(n16130), .A(n16129), .ZN(n16133) );
  OR2_X1 U19219 ( .A1(n16133), .A2(n16132), .ZN(n19984) );
  INV_X1 U19220 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n16135) );
  OAI22_X1 U19221 ( .A1(n19984), .A2(n16136), .B1(n16135), .B2(n16134), .ZN(
        n16140) );
  NOR2_X1 U19222 ( .A1(n16138), .A2(n16137), .ZN(n16139) );
  AOI211_X1 U19223 ( .C1(n16142), .C2(n16141), .A(n16140), .B(n16139), .ZN(
        n16143) );
  OAI21_X1 U19224 ( .B1(n16144), .B2(n16142), .A(n16143), .ZN(P1_U3025) );
  OAI221_X1 U19225 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n20744), .C2(n20647), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n20636) );
  NAND2_X1 U19226 ( .A1(n16145), .A2(n20636), .ZN(n16146) );
  AOI22_X1 U19227 ( .A1(n16149), .A2(n16148), .B1(n16147), .B2(n16146), .ZN(
        P1_U3162) );
  OAI21_X1 U19228 ( .B1(n20635), .B2(n20338), .A(n16150), .ZN(P1_U3466) );
  AOI211_X1 U19229 ( .C1(n16153), .C2(n16151), .A(n16152), .B(n19717), .ZN(
        n16157) );
  AOI22_X1 U19230 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19000), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n18951), .ZN(n16154) );
  OAI21_X1 U19231 ( .B1(n16155), .B2(n18995), .A(n16154), .ZN(n16156) );
  AOI211_X1 U19232 ( .C1(P2_EBX_REG_24__SCAN_IN), .C2(n18992), .A(n16157), .B(
        n16156), .ZN(n16162) );
  INV_X1 U19233 ( .A(n16158), .ZN(n16159) );
  AOI22_X1 U19234 ( .A1(n16160), .A2(n18999), .B1(n18954), .B2(n16159), .ZN(
        n16161) );
  NAND2_X1 U19235 ( .A1(n16162), .A2(n16161), .ZN(P2_U2831) );
  AOI22_X1 U19236 ( .A1(n19009), .A2(n16163), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19055), .ZN(n16167) );
  AOI22_X1 U19237 ( .A1(n19011), .A2(BUF2_REG_20__SCAN_IN), .B1(n19010), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n16166) );
  AOI22_X1 U19238 ( .A1(n16164), .A2(n13149), .B1(n19056), .B2(n18897), .ZN(
        n16165) );
  NAND3_X1 U19239 ( .A1(n16167), .A2(n16166), .A3(n16165), .ZN(P2_U2899) );
  AOI22_X1 U19240 ( .A1(n19009), .A2(n16168), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19055), .ZN(n16172) );
  AOI22_X1 U19241 ( .A1(n19011), .A2(BUF2_REG_18__SCAN_IN), .B1(n19010), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n16171) );
  AOI22_X1 U19242 ( .A1(n16169), .A2(n13149), .B1(n19056), .B2(n18916), .ZN(
        n16170) );
  NAND3_X1 U19243 ( .A1(n16172), .A2(n16171), .A3(n16170), .ZN(P2_U2901) );
  AOI22_X1 U19244 ( .A1(n19114), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n16279), .ZN(n16177) );
  OAI22_X1 U19245 ( .A1(n16173), .A2(n16256), .B1(n16247), .B2(n18952), .ZN(
        n16174) );
  AOI21_X1 U19246 ( .B1(n16175), .B2(n19121), .A(n16174), .ZN(n16176) );
  OAI211_X1 U19247 ( .C1(n19125), .C2(n18945), .A(n16177), .B(n16176), .ZN(
        P2_U3000) );
  AOI22_X1 U19248 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n16279), .B1(n16255), 
        .B2(n16178), .ZN(n16188) );
  AND2_X1 U19249 ( .A1(n16180), .A2(n16179), .ZN(n16181) );
  XNOR2_X1 U19250 ( .A(n16182), .B(n16181), .ZN(n16283) );
  INV_X1 U19251 ( .A(n16283), .ZN(n16184) );
  AND2_X1 U19252 ( .A1(n15748), .A2(n16276), .ZN(n16183) );
  OR2_X1 U19253 ( .A1(n16183), .A2(n15726), .ZN(n16281) );
  OAI22_X1 U19254 ( .A1(n16184), .A2(n16258), .B1(n16256), .B2(n16281), .ZN(
        n16185) );
  AOI21_X1 U19255 ( .B1(n19117), .B2(n16186), .A(n16185), .ZN(n16187) );
  OAI211_X1 U19256 ( .C1(n16265), .C2(n16189), .A(n16188), .B(n16187), .ZN(
        P2_U3001) );
  AOI22_X1 U19257 ( .A1(n19114), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19113), .ZN(n16197) );
  NAND2_X1 U19258 ( .A1(n16190), .A2(n19121), .ZN(n16193) );
  OR2_X1 U19259 ( .A1(n16191), .A2(n16247), .ZN(n16192) );
  OAI211_X1 U19260 ( .C1(n16194), .C2(n16256), .A(n16193), .B(n16192), .ZN(
        n16195) );
  INV_X1 U19261 ( .A(n16195), .ZN(n16196) );
  OAI211_X1 U19262 ( .C1(n19125), .C2(n16198), .A(n16197), .B(n16196), .ZN(
        P2_U3002) );
  AOI22_X1 U19263 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19113), .B1(n16255), 
        .B2(n16199), .ZN(n16205) );
  OAI22_X1 U19264 ( .A1(n16201), .A2(n16256), .B1(n16200), .B2(n16258), .ZN(
        n16202) );
  AOI21_X1 U19265 ( .B1(n19117), .B2(n16203), .A(n16202), .ZN(n16204) );
  OAI211_X1 U19266 ( .C1(n16265), .C2(n16206), .A(n16205), .B(n16204), .ZN(
        P2_U3003) );
  AOI22_X1 U19267 ( .A1(n19114), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19113), .ZN(n16219) );
  OAI21_X1 U19268 ( .B1(n16208), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16207), .ZN(n16292) );
  OAI22_X1 U19269 ( .A1(n16292), .A2(n16256), .B1(n16247), .B2(n16291), .ZN(
        n16217) );
  INV_X1 U19270 ( .A(n16209), .ZN(n16210) );
  OR2_X1 U19271 ( .A1(n16211), .A2(n16210), .ZN(n16215) );
  AND2_X1 U19272 ( .A1(n16213), .A2(n16212), .ZN(n16214) );
  XNOR2_X1 U19273 ( .A(n16215), .B(n16214), .ZN(n16296) );
  NOR2_X1 U19274 ( .A1(n16296), .A2(n16258), .ZN(n16216) );
  NOR2_X1 U19275 ( .A1(n16217), .A2(n16216), .ZN(n16218) );
  OAI211_X1 U19276 ( .C1(n19125), .C2(n16220), .A(n16219), .B(n16218), .ZN(
        P2_U3004) );
  AOI22_X1 U19277 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n16279), .B1(n16255), 
        .B2(n18960), .ZN(n16226) );
  OAI22_X1 U19278 ( .A1(n16222), .A2(n16256), .B1(n16258), .B2(n16221), .ZN(
        n16223) );
  AOI21_X1 U19279 ( .B1(n19117), .B2(n16224), .A(n16223), .ZN(n16225) );
  OAI211_X1 U19280 ( .C1(n16265), .C2(n16227), .A(n16226), .B(n16225), .ZN(
        P2_U3005) );
  AOI22_X1 U19281 ( .A1(n19114), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19113), .ZN(n16244) );
  NAND2_X1 U19282 ( .A1(n16228), .A2(n16229), .ZN(n16230) );
  NAND2_X1 U19283 ( .A1(n16231), .A2(n16230), .ZN(n16306) );
  NAND2_X1 U19284 ( .A1(n14340), .A2(n16232), .ZN(n16234) );
  NAND2_X1 U19285 ( .A1(n16234), .A2(n16233), .ZN(n16238) );
  NAND2_X1 U19286 ( .A1(n16236), .A2(n16235), .ZN(n16237) );
  XNOR2_X1 U19287 ( .A(n16238), .B(n16237), .ZN(n16301) );
  NAND2_X1 U19288 ( .A1(n16301), .A2(n19121), .ZN(n16241) );
  INV_X1 U19289 ( .A(n16239), .ZN(n16303) );
  NAND2_X1 U19290 ( .A1(n16303), .A2(n19117), .ZN(n16240) );
  OAI211_X1 U19291 ( .C1(n16306), .C2(n16256), .A(n16241), .B(n16240), .ZN(
        n16242) );
  INV_X1 U19292 ( .A(n16242), .ZN(n16243) );
  OAI211_X1 U19293 ( .C1(n19125), .C2(n16245), .A(n16244), .B(n16243), .ZN(
        P2_U3006) );
  AOI22_X1 U19294 ( .A1(n19114), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n19113), .ZN(n16252) );
  OAI22_X1 U19295 ( .A1(n16248), .A2(n16256), .B1(n16247), .B2(n16246), .ZN(
        n16249) );
  AOI21_X1 U19296 ( .B1(n19121), .B2(n16250), .A(n16249), .ZN(n16251) );
  OAI211_X1 U19297 ( .C1(n19125), .C2(n16253), .A(n16252), .B(n16251), .ZN(
        P2_U3008) );
  AOI22_X1 U19298 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n16279), .B1(n16255), 
        .B2(n16254), .ZN(n16263) );
  OAI22_X1 U19299 ( .A1(n16259), .A2(n16258), .B1(n16257), .B2(n16256), .ZN(
        n16260) );
  AOI21_X1 U19300 ( .B1(n19117), .B2(n16261), .A(n16260), .ZN(n16262) );
  OAI211_X1 U19301 ( .C1(n16265), .C2(n16264), .A(n16263), .B(n16262), .ZN(
        P2_U3009) );
  OAI22_X1 U19302 ( .A1(n19143), .A2(n19018), .B1(n11227), .B2(n15534), .ZN(
        n16266) );
  AOI221_X1 U19303 ( .B1(n16268), .B2(n10667), .C1(n16267), .C2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(n16266), .ZN(n16274) );
  INV_X1 U19304 ( .A(n16269), .ZN(n16272) );
  AOI22_X1 U19305 ( .A1(n16272), .A2(n16271), .B1(n16302), .B2(n16270), .ZN(
        n16273) );
  OAI211_X1 U19306 ( .C1(n19133), .C2(n16275), .A(n16274), .B(n16273), .ZN(
        P2_U3031) );
  OAI22_X1 U19307 ( .A1(n16277), .A2(n16276), .B1(n19143), .B2(n19022), .ZN(
        n16278) );
  AOI21_X1 U19308 ( .B1(P2_REIP_REG_13__SCAN_IN), .B2(n16279), .A(n16278), 
        .ZN(n16285) );
  OAI22_X1 U19309 ( .A1(n16281), .A2(n19137), .B1(n19138), .B2(n16280), .ZN(
        n16282) );
  AOI21_X1 U19310 ( .B1(n16300), .B2(n16283), .A(n16282), .ZN(n16284) );
  OAI211_X1 U19311 ( .C1(n10644), .C2(n16286), .A(n16285), .B(n16284), .ZN(
        P2_U3033) );
  NOR2_X1 U19312 ( .A1(n11146), .A2(n15534), .ZN(n16289) );
  OAI22_X1 U19313 ( .A1(n16287), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n19030), .B2(n19143), .ZN(n16288) );
  AOI211_X1 U19314 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n16290), .A(
        n16289), .B(n16288), .ZN(n16295) );
  OAI22_X1 U19315 ( .A1(n16292), .A2(n19137), .B1(n19138), .B2(n16291), .ZN(
        n16293) );
  INV_X1 U19316 ( .A(n16293), .ZN(n16294) );
  OAI211_X1 U19317 ( .C1(n16296), .C2(n19133), .A(n16295), .B(n16294), .ZN(
        P2_U3036) );
  INV_X1 U19318 ( .A(n19036), .ZN(n16297) );
  AOI22_X1 U19319 ( .A1(n16299), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16298), .B2(n16297), .ZN(n16314) );
  NAND2_X1 U19320 ( .A1(n16301), .A2(n16300), .ZN(n16305) );
  NAND2_X1 U19321 ( .A1(n16303), .A2(n16302), .ZN(n16304) );
  OAI211_X1 U19322 ( .C1(n16306), .C2(n19137), .A(n16305), .B(n16304), .ZN(
        n16307) );
  INV_X1 U19323 ( .A(n16307), .ZN(n16313) );
  NAND2_X1 U19324 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19113), .ZN(n16312) );
  INV_X1 U19325 ( .A(n16308), .ZN(n16309) );
  OAI211_X1 U19326 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16310), .B(n16309), .ZN(n16311) );
  NAND4_X1 U19327 ( .A1(n16314), .A2(n16313), .A3(n16312), .A4(n16311), .ZN(
        P2_U3038) );
  AND2_X1 U19328 ( .A1(n16315), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n16319) );
  NAND2_X1 U19329 ( .A1(n19822), .A2(n16316), .ZN(n16318) );
  AOI221_X1 U19330 ( .B1(n16319), .B2(n16318), .C1(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n16317), .A(n16333), .ZN(
        n16327) );
  INV_X1 U19331 ( .A(n16333), .ZN(n16320) );
  AOI22_X1 U19332 ( .A1(n16333), .A2(n16322), .B1(n16321), .B2(n16320), .ZN(
        n16332) );
  NOR2_X1 U19333 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n16332), .ZN(
        n16326) );
  MUX2_X1 U19334 ( .A(n16323), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n16333), .Z(n16356) );
  INV_X1 U19335 ( .A(n16356), .ZN(n16324) );
  AOI21_X1 U19336 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16324), .A(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n16325) );
  AOI222_X1 U19337 ( .A1(n16327), .A2(n16326), .B1(n16327), .B2(n16325), .C1(
        n16326), .C2(n19813), .ZN(n16329) );
  NAND2_X1 U19338 ( .A1(n16356), .A2(n19803), .ZN(n16328) );
  NAND2_X1 U19339 ( .A1(n16329), .A2(n16328), .ZN(n16331) );
  NAND2_X1 U19340 ( .A1(n16331), .A2(n16330), .ZN(n16358) );
  INV_X1 U19341 ( .A(n16332), .ZN(n16355) );
  NAND2_X1 U19342 ( .A1(n16333), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n16353) );
  NAND2_X1 U19343 ( .A1(n16335), .A2(n16334), .ZN(n16342) );
  INV_X1 U19344 ( .A(n16336), .ZN(n16338) );
  AOI22_X1 U19345 ( .A1(n16340), .A2(n16339), .B1(n16338), .B2(n16337), .ZN(
        n16341) );
  AND2_X1 U19346 ( .A1(n16342), .A2(n16341), .ZN(n19835) );
  INV_X1 U19347 ( .A(n16343), .ZN(n16344) );
  NAND2_X1 U19348 ( .A1(n10364), .A2(n16344), .ZN(n16345) );
  OAI22_X1 U19349 ( .A1(n10966), .A2(n16345), .B1(n10727), .B2(n19846), .ZN(
        n16346) );
  INV_X1 U19350 ( .A(n16346), .ZN(n16352) );
  NOR2_X1 U19351 ( .A1(n16348), .A2(n16347), .ZN(n16349) );
  AND2_X1 U19352 ( .A1(n16350), .A2(n16349), .ZN(n18864) );
  OAI21_X1 U19353 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n18864), .ZN(n16351) );
  NAND4_X1 U19354 ( .A1(n16353), .A2(n19835), .A3(n16352), .A4(n16351), .ZN(
        n16354) );
  AOI21_X1 U19355 ( .B1(n16356), .B2(n16355), .A(n16354), .ZN(n16357) );
  AND2_X1 U19356 ( .A1(n16358), .A2(n16357), .ZN(n16374) );
  INV_X1 U19357 ( .A(n16359), .ZN(n16364) );
  INV_X1 U19358 ( .A(n16360), .ZN(n16362) );
  OR2_X1 U19359 ( .A1(n19840), .A2(n19848), .ZN(n16361) );
  AOI21_X1 U19360 ( .B1(n16363), .B2(n16362), .A(n16361), .ZN(n16370) );
  AOI22_X1 U19361 ( .A1(n16364), .A2(n19850), .B1(n19849), .B2(n16370), .ZN(
        n16367) );
  AOI211_X1 U19362 ( .C1(n16367), .C2(n13325), .A(n16366), .B(n16365), .ZN(
        n16373) );
  NAND2_X1 U19363 ( .A1(n16374), .A2(n10302), .ZN(n16369) );
  NAND2_X1 U19364 ( .A1(n16369), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16371) );
  OAI21_X1 U19365 ( .B1(n10121), .B2(n19719), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n16372) );
  OAI211_X1 U19366 ( .C1(n16374), .C2(n18863), .A(n16373), .B(n16372), .ZN(
        P2_U3176) );
  INV_X1 U19367 ( .A(n19719), .ZN(n16376) );
  OAI221_X1 U19368 ( .B1(n19839), .B2(P2_STATE2_REG_0__SCAN_IN), .C1(n19839), 
        .C2(n16376), .A(n16375), .ZN(P2_U3593) );
  INV_X1 U19369 ( .A(n16377), .ZN(n16378) );
  NOR2_X1 U19370 ( .A1(n17627), .A2(n16378), .ZN(n16386) );
  NAND2_X1 U19371 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17627), .ZN(
        n16381) );
  OAI211_X1 U19372 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n17627), .A(
        n16379), .B(n16381), .ZN(n16385) );
  OAI21_X1 U19373 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n20799), .A(
        n16380), .ZN(n16383) );
  OAI22_X1 U19374 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17627), .B1(
        n16381), .B2(n20799), .ZN(n16382) );
  OAI21_X1 U19375 ( .B1(n16386), .B2(n16383), .A(n16382), .ZN(n16384) );
  OAI21_X1 U19376 ( .B1(n16386), .B2(n16385), .A(n16384), .ZN(n16423) );
  INV_X1 U19377 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18779) );
  NOR2_X1 U19378 ( .A1(n18779), .A2(n18122), .ZN(n16417) );
  XNOR2_X1 U19379 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16388) );
  OAI22_X1 U19380 ( .A1(n16389), .A2(n16388), .B1(n16387), .B2(n16578), .ZN(
        n16390) );
  AOI211_X1 U19381 ( .C1(n17649), .C2(n16876), .A(n16417), .B(n16390), .ZN(
        n16396) );
  INV_X1 U19382 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18803) );
  OR2_X1 U19383 ( .A1(n20799), .A2(n16391), .ZN(n16392) );
  XOR2_X1 U19384 ( .A(n18803), .B(n16392), .Z(n16420) );
  OR2_X1 U19385 ( .A1(n20799), .A2(n16393), .ZN(n16394) );
  XOR2_X1 U19386 ( .A(n18803), .B(n16394), .Z(n16419) );
  AOI22_X1 U19387 ( .A1(n17753), .A2(n16420), .B1(n17837), .B2(n16419), .ZN(
        n16395) );
  OAI211_X1 U19388 ( .C1(n17756), .C2(n16423), .A(n16396), .B(n16395), .ZN(
        P3_U2799) );
  OR2_X1 U19389 ( .A1(n16431), .A2(n16430), .ZN(n16410) );
  AOI21_X1 U19390 ( .B1(n9925), .B2(n16399), .A(n16398), .ZN(n16591) );
  OAI21_X1 U19391 ( .B1(n16400), .B2(n17649), .A(n16591), .ZN(n16401) );
  OAI211_X1 U19392 ( .C1(n16403), .C2(n9926), .A(n16402), .B(n16401), .ZN(
        n16407) );
  NOR2_X1 U19393 ( .A1(n17858), .A2(n16431), .ZN(n16434) );
  NOR2_X1 U19394 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16434), .ZN(
        n16406) );
  OAI221_X1 U19395 ( .B1(n16411), .B2(n12799), .C1(n16411), .C2(n16410), .A(
        n16409), .ZN(P3_U2801) );
  INV_X1 U19396 ( .A(n18157), .ZN(n18082) );
  OAI21_X1 U19397 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18082), .A(
        n16412), .ZN(n16418) );
  NAND2_X1 U19398 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18803), .ZN(
        n16414) );
  NOR4_X1 U19399 ( .A1(n16415), .A2(n16414), .A3(n18154), .A4(n16413), .ZN(
        n16416) );
  AOI211_X1 U19400 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16418), .A(
        n16417), .B(n16416), .ZN(n16422) );
  AOI22_X1 U19401 ( .A1(n16420), .A2(n18087), .B1(n16419), .B2(n18152), .ZN(
        n16421) );
  OAI211_X1 U19402 ( .C1(n16423), .C2(n18091), .A(n16422), .B(n16421), .ZN(
        P3_U2831) );
  OAI22_X1 U19403 ( .A1(n18626), .A2(n17711), .B1(n17712), .B2(n18045), .ZN(
        n17968) );
  NOR2_X1 U19404 ( .A1(n17609), .A2(n17969), .ZN(n16424) );
  AOI21_X1 U19405 ( .B1(n17968), .B2(n16424), .A(n17877), .ZN(n17912) );
  OR2_X1 U19406 ( .A1(n18154), .A2(n17912), .ZN(n17930) );
  NOR2_X1 U19407 ( .A1(n17867), .A2(n17930), .ZN(n17892) );
  NOR2_X1 U19408 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16425), .ZN(
        n17482) );
  AOI22_X1 U19409 ( .A1(n18153), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n17892), 
        .B2(n17482), .ZN(n16440) );
  INV_X1 U19410 ( .A(n18169), .ZN(n18150) );
  NAND3_X1 U19411 ( .A1(n17488), .A2(n18150), .A3(n16426), .ZN(n16439) );
  AOI22_X1 U19412 ( .A1(n17627), .A2(n17476), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17743), .ZN(n17479) );
  NAND3_X1 U19413 ( .A1(n17487), .A2(n18072), .A3(n17479), .ZN(n16438) );
  INV_X1 U19414 ( .A(n17488), .ZN(n16427) );
  AOI21_X1 U19415 ( .B1(n17627), .B2(n16427), .A(n17487), .ZN(n17478) );
  NOR2_X1 U19416 ( .A1(n17479), .A2(n17478), .ZN(n17477) );
  NOR4_X1 U19417 ( .A1(n17321), .A2(n16429), .A3(n17477), .A4(n16428), .ZN(
        n16436) );
  OAI21_X1 U19418 ( .B1(n16431), .B2(n16430), .A(n17918), .ZN(n16432) );
  OAI211_X1 U19419 ( .C1(n16434), .C2(n18045), .A(n16433), .B(n16432), .ZN(
        n16435) );
  OAI211_X1 U19420 ( .C1(n16436), .C2(n16435), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18122), .ZN(n16437) );
  NAND4_X1 U19421 ( .A1(n16440), .A2(n16439), .A3(n16438), .A4(n16437), .ZN(
        P3_U2834) );
  NOR3_X1 U19422 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16442) );
  NOR4_X1 U19423 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16441) );
  NAND4_X1 U19424 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16442), .A3(n16441), .A4(
        U215), .ZN(U213) );
  INV_X1 U19425 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16526) );
  INV_X2 U19426 ( .A(U214), .ZN(n16490) );
  NOR2_X2 U19427 ( .A1(n16490), .A2(n16443), .ZN(n16491) );
  INV_X1 U19428 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19066) );
  OAI222_X1 U19429 ( .A1(U214), .A2(n16526), .B1(n16494), .B2(n19165), .C1(
        U212), .C2(n19066), .ZN(U216) );
  INV_X1 U19430 ( .A(U212), .ZN(n16487) );
  AOI222_X1 U19431 ( .A1(n16490), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16491), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n16487), .C2(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n16444) );
  INV_X1 U19432 ( .A(n16444), .ZN(U217) );
  INV_X1 U19433 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16446) );
  AOI22_X1 U19434 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n16487), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n16490), .ZN(n16445) );
  OAI21_X1 U19435 ( .B1(n16446), .B2(n16494), .A(n16445), .ZN(U218) );
  INV_X1 U19436 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16448) );
  AOI22_X1 U19437 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16487), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16490), .ZN(n16447) );
  OAI21_X1 U19438 ( .B1(n16448), .B2(n16494), .A(n16447), .ZN(U219) );
  AOI22_X1 U19439 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16487), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16490), .ZN(n16449) );
  OAI21_X1 U19440 ( .B1(n16450), .B2(n16494), .A(n16449), .ZN(U220) );
  INV_X1 U19441 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16452) );
  AOI22_X1 U19442 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16487), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16490), .ZN(n16451) );
  OAI21_X1 U19443 ( .B1(n16452), .B2(n16494), .A(n16451), .ZN(U221) );
  INV_X1 U19444 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n20901) );
  AOI22_X1 U19445 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n16491), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n16490), .ZN(n16453) );
  OAI21_X1 U19446 ( .B1(n20901), .B2(U212), .A(n16453), .ZN(U222) );
  INV_X1 U19447 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16455) );
  AOI22_X1 U19448 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16487), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16490), .ZN(n16454) );
  OAI21_X1 U19449 ( .B1(n16455), .B2(n16494), .A(n16454), .ZN(U223) );
  INV_X1 U19450 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16457) );
  AOI22_X1 U19451 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16487), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16490), .ZN(n16456) );
  OAI21_X1 U19452 ( .B1(n16457), .B2(n16494), .A(n16456), .ZN(U224) );
  AOI22_X1 U19453 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16487), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16490), .ZN(n16458) );
  OAI21_X1 U19454 ( .B1(n16459), .B2(n16494), .A(n16458), .ZN(U225) );
  AOI222_X1 U19455 ( .A1(n16490), .A2(P1_DATAO_REG_21__SCAN_IN), .B1(n16491), 
        .B2(BUF1_REG_21__SCAN_IN), .C1(n16487), .C2(P2_DATAO_REG_21__SCAN_IN), 
        .ZN(n16460) );
  INV_X1 U19456 ( .A(n16460), .ZN(U226) );
  INV_X1 U19457 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16462) );
  AOI22_X1 U19458 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16487), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16490), .ZN(n16461) );
  OAI21_X1 U19459 ( .B1(n16462), .B2(n16494), .A(n16461), .ZN(U227) );
  AOI22_X1 U19460 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n16487), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16490), .ZN(n16463) );
  OAI21_X1 U19461 ( .B1(n15411), .B2(n16494), .A(n16463), .ZN(U228) );
  INV_X1 U19462 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16465) );
  AOI22_X1 U19463 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16487), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16490), .ZN(n16464) );
  OAI21_X1 U19464 ( .B1(n16465), .B2(n16494), .A(n16464), .ZN(U229) );
  INV_X1 U19465 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20826) );
  AOI22_X1 U19466 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16487), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16490), .ZN(n16466) );
  OAI21_X1 U19467 ( .B1(n20826), .B2(n16494), .A(n16466), .ZN(U230) );
  INV_X1 U19468 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16468) );
  AOI22_X1 U19469 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16487), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16490), .ZN(n16467) );
  OAI21_X1 U19470 ( .B1(n16468), .B2(n16494), .A(n16467), .ZN(U231) );
  INV_X1 U19471 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n16510) );
  AOI22_X1 U19472 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n16491), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16490), .ZN(n16469) );
  OAI21_X1 U19473 ( .B1(n16510), .B2(U212), .A(n16469), .ZN(U232) );
  INV_X1 U19474 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n16471) );
  AOI22_X1 U19475 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n16491), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16490), .ZN(n16470) );
  OAI21_X1 U19476 ( .B1(n16471), .B2(U212), .A(n16470), .ZN(U233) );
  INV_X1 U19477 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n20802) );
  AOI22_X1 U19478 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n16491), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16487), .ZN(n16472) );
  OAI21_X1 U19479 ( .B1(n20802), .B2(U214), .A(n16472), .ZN(U234) );
  AOI22_X1 U19480 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n16487), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16490), .ZN(n16473) );
  OAI21_X1 U19481 ( .B1(n16474), .B2(n16494), .A(n16473), .ZN(U235) );
  INV_X1 U19482 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16476) );
  AOI22_X1 U19483 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n16491), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16490), .ZN(n16475) );
  OAI21_X1 U19484 ( .B1(n16476), .B2(U212), .A(n16475), .ZN(U236) );
  AOI22_X1 U19485 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n16487), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16490), .ZN(n16477) );
  OAI21_X1 U19486 ( .B1(n16478), .B2(n16494), .A(n16477), .ZN(U237) );
  INV_X1 U19487 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16504) );
  AOI22_X1 U19488 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16491), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16490), .ZN(n16479) );
  OAI21_X1 U19489 ( .B1(n16504), .B2(U212), .A(n16479), .ZN(U238) );
  AOI22_X1 U19490 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n16487), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16490), .ZN(n16480) );
  OAI21_X1 U19491 ( .B1(n16481), .B2(n16494), .A(n16480), .ZN(U239) );
  INV_X1 U19492 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16502) );
  AOI22_X1 U19493 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16491), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16490), .ZN(n16482) );
  OAI21_X1 U19494 ( .B1(n16502), .B2(U212), .A(n16482), .ZN(U240) );
  INV_X1 U19495 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16501) );
  AOI22_X1 U19496 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n16491), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16490), .ZN(n16483) );
  OAI21_X1 U19497 ( .B1(n16501), .B2(U212), .A(n16483), .ZN(U241) );
  INV_X1 U19498 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16500) );
  AOI22_X1 U19499 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16491), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16490), .ZN(n16484) );
  OAI21_X1 U19500 ( .B1(n16500), .B2(U212), .A(n16484), .ZN(U242) );
  INV_X1 U19501 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n20834) );
  AOI22_X1 U19502 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n16487), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16490), .ZN(n16485) );
  OAI21_X1 U19503 ( .B1(n20834), .B2(n16494), .A(n16485), .ZN(U243) );
  INV_X1 U19504 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16498) );
  AOI22_X1 U19505 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16491), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16490), .ZN(n16486) );
  OAI21_X1 U19506 ( .B1(n16498), .B2(U212), .A(n16486), .ZN(U244) );
  INV_X1 U19507 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16489) );
  AOI22_X1 U19508 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n16487), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16490), .ZN(n16488) );
  OAI21_X1 U19509 ( .B1(n16489), .B2(n16494), .A(n16488), .ZN(U245) );
  INV_X1 U19510 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16496) );
  AOI22_X1 U19511 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16491), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16490), .ZN(n16492) );
  OAI21_X1 U19512 ( .B1(n16496), .B2(U212), .A(n16492), .ZN(U246) );
  INV_X1 U19513 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n20816) );
  INV_X1 U19514 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16493) );
  INV_X1 U19515 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16495) );
  OAI222_X1 U19516 ( .A1(U214), .A2(n20816), .B1(n16494), .B2(n16493), .C1(
        U212), .C2(n16495), .ZN(U247) );
  INV_X1 U19517 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18186) );
  AOI22_X1 U19518 ( .A1(n16523), .A2(n16495), .B1(n18186), .B2(U215), .ZN(U251) );
  INV_X1 U19519 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18195) );
  AOI22_X1 U19520 ( .A1(n16523), .A2(n16496), .B1(n18195), .B2(U215), .ZN(U252) );
  OAI22_X1 U19521 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16523), .ZN(n16497) );
  INV_X1 U19522 ( .A(n16497), .ZN(U253) );
  INV_X1 U19523 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n20912) );
  AOI22_X1 U19524 ( .A1(n16523), .A2(n16498), .B1(n20912), .B2(U215), .ZN(U254) );
  OAI22_X1 U19525 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16523), .ZN(n16499) );
  INV_X1 U19526 ( .A(n16499), .ZN(U255) );
  INV_X1 U19527 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18213) );
  AOI22_X1 U19528 ( .A1(n16523), .A2(n16500), .B1(n18213), .B2(U215), .ZN(U256) );
  INV_X1 U19529 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18218) );
  AOI22_X1 U19530 ( .A1(n16523), .A2(n16501), .B1(n18218), .B2(U215), .ZN(U257) );
  INV_X1 U19531 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18222) );
  AOI22_X1 U19532 ( .A1(n16523), .A2(n16502), .B1(n18222), .B2(U215), .ZN(U258) );
  OAI22_X1 U19533 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16523), .ZN(n16503) );
  INV_X1 U19534 ( .A(n16503), .ZN(U259) );
  INV_X1 U19535 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17450) );
  AOI22_X1 U19536 ( .A1(n16525), .A2(n16504), .B1(n17450), .B2(U215), .ZN(U260) );
  OAI22_X1 U19537 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16523), .ZN(n16505) );
  INV_X1 U19538 ( .A(n16505), .ZN(U261) );
  OAI22_X1 U19539 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16523), .ZN(n16506) );
  INV_X1 U19540 ( .A(n16506), .ZN(U262) );
  OAI22_X1 U19541 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16523), .ZN(n16507) );
  INV_X1 U19542 ( .A(n16507), .ZN(U263) );
  OAI22_X1 U19543 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16523), .ZN(n16508) );
  INV_X1 U19544 ( .A(n16508), .ZN(U264) );
  OAI22_X1 U19545 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16523), .ZN(n16509) );
  INV_X1 U19546 ( .A(n16509), .ZN(U265) );
  INV_X1 U19547 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n17291) );
  AOI22_X1 U19548 ( .A1(n16523), .A2(n16510), .B1(n17291), .B2(U215), .ZN(U266) );
  OAI22_X1 U19549 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16523), .ZN(n16511) );
  INV_X1 U19550 ( .A(n16511), .ZN(U267) );
  OAI22_X1 U19551 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16525), .ZN(n16512) );
  INV_X1 U19552 ( .A(n16512), .ZN(U268) );
  OAI22_X1 U19553 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16525), .ZN(n16513) );
  INV_X1 U19554 ( .A(n16513), .ZN(U269) );
  OAI22_X1 U19555 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16525), .ZN(n16514) );
  INV_X1 U19556 ( .A(n16514), .ZN(U270) );
  OAI22_X1 U19557 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16525), .ZN(n16515) );
  INV_X1 U19558 ( .A(n16515), .ZN(U271) );
  INV_X1 U19559 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n20911) );
  AOI22_X1 U19560 ( .A1(n16523), .A2(n20911), .B1(n18212), .B2(U215), .ZN(U272) );
  OAI22_X1 U19561 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16525), .ZN(n16516) );
  INV_X1 U19562 ( .A(n16516), .ZN(U273) );
  OAI22_X1 U19563 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16525), .ZN(n16517) );
  INV_X1 U19564 ( .A(n16517), .ZN(U274) );
  OAI22_X1 U19565 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16525), .ZN(n16518) );
  INV_X1 U19566 ( .A(n16518), .ZN(U275) );
  INV_X1 U19567 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18194) );
  AOI22_X1 U19568 ( .A1(n16525), .A2(n20901), .B1(n18194), .B2(U215), .ZN(U276) );
  OAI22_X1 U19569 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16523), .ZN(n16519) );
  INV_X1 U19570 ( .A(n16519), .ZN(U277) );
  OAI22_X1 U19571 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16523), .ZN(n16520) );
  INV_X1 U19572 ( .A(n16520), .ZN(U278) );
  OAI22_X1 U19573 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16523), .ZN(n16521) );
  INV_X1 U19574 ( .A(n16521), .ZN(U279) );
  OAI22_X1 U19575 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16523), .ZN(n16522) );
  INV_X1 U19576 ( .A(n16522), .ZN(U280) );
  OAI22_X1 U19577 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16523), .ZN(n16524) );
  INV_X1 U19578 ( .A(n16524), .ZN(U281) );
  INV_X1 U19579 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19163) );
  AOI22_X1 U19580 ( .A1(n16525), .A2(n19066), .B1(n19163), .B2(U215), .ZN(U282) );
  INV_X1 U19581 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n20915) );
  AOI222_X1 U19582 ( .A1(n19066), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16526), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n20915), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16527) );
  INV_X2 U19583 ( .A(n16529), .ZN(n16528) );
  INV_X1 U19584 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18739) );
  INV_X1 U19585 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19750) );
  AOI22_X1 U19586 ( .A1(n16528), .A2(n18739), .B1(n19750), .B2(n16529), .ZN(
        U347) );
  INV_X1 U19587 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18737) );
  INV_X1 U19588 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19749) );
  AOI22_X1 U19589 ( .A1(n16528), .A2(n18737), .B1(n19749), .B2(n16529), .ZN(
        U348) );
  INV_X1 U19590 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18735) );
  INV_X1 U19591 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19748) );
  AOI22_X1 U19592 ( .A1(n16528), .A2(n18735), .B1(n19748), .B2(n16529), .ZN(
        U349) );
  INV_X1 U19593 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18733) );
  INV_X1 U19594 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19747) );
  AOI22_X1 U19595 ( .A1(n16528), .A2(n18733), .B1(n19747), .B2(n16529), .ZN(
        U350) );
  INV_X1 U19596 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18731) );
  INV_X1 U19597 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19746) );
  AOI22_X1 U19598 ( .A1(n16528), .A2(n18731), .B1(n19746), .B2(n16529), .ZN(
        U351) );
  INV_X1 U19599 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18728) );
  INV_X1 U19600 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19745) );
  AOI22_X1 U19601 ( .A1(n16528), .A2(n18728), .B1(n19745), .B2(n16529), .ZN(
        U352) );
  INV_X1 U19602 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18727) );
  INV_X1 U19603 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19744) );
  AOI22_X1 U19604 ( .A1(n16528), .A2(n18727), .B1(n19744), .B2(n16529), .ZN(
        U353) );
  INV_X1 U19605 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18724) );
  AOI22_X1 U19606 ( .A1(n16528), .A2(n18724), .B1(n19743), .B2(n16529), .ZN(
        U354) );
  INV_X1 U19607 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18781) );
  INV_X1 U19608 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19781) );
  AOI22_X1 U19609 ( .A1(n16528), .A2(n18781), .B1(n19781), .B2(n16529), .ZN(
        U355) );
  INV_X1 U19610 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18778) );
  INV_X1 U19611 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20829) );
  AOI22_X1 U19612 ( .A1(n16528), .A2(n18778), .B1(n20829), .B2(n16529), .ZN(
        U356) );
  INV_X1 U19613 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18775) );
  INV_X1 U19614 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19777) );
  AOI22_X1 U19615 ( .A1(n16528), .A2(n18775), .B1(n19777), .B2(n16529), .ZN(
        U357) );
  INV_X1 U19616 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18774) );
  INV_X1 U19617 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19774) );
  AOI22_X1 U19618 ( .A1(n16528), .A2(n18774), .B1(n19774), .B2(n16529), .ZN(
        U358) );
  INV_X1 U19619 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18772) );
  INV_X1 U19620 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19773) );
  AOI22_X1 U19621 ( .A1(n16528), .A2(n18772), .B1(n19773), .B2(n16529), .ZN(
        U359) );
  INV_X1 U19622 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18770) );
  INV_X1 U19623 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19772) );
  AOI22_X1 U19624 ( .A1(n16528), .A2(n18770), .B1(n19772), .B2(n16529), .ZN(
        U360) );
  INV_X1 U19625 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18767) );
  INV_X1 U19626 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19770) );
  AOI22_X1 U19627 ( .A1(n16528), .A2(n18767), .B1(n19770), .B2(n16529), .ZN(
        U361) );
  INV_X1 U19628 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18765) );
  INV_X1 U19629 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19768) );
  AOI22_X1 U19630 ( .A1(n16528), .A2(n18765), .B1(n19768), .B2(n16529), .ZN(
        U362) );
  INV_X1 U19631 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18763) );
  INV_X1 U19632 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19766) );
  AOI22_X1 U19633 ( .A1(n16528), .A2(n18763), .B1(n19766), .B2(n16529), .ZN(
        U363) );
  INV_X1 U19634 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18761) );
  INV_X1 U19635 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19764) );
  AOI22_X1 U19636 ( .A1(n16528), .A2(n18761), .B1(n19764), .B2(n16529), .ZN(
        U364) );
  INV_X1 U19637 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18722) );
  INV_X1 U19638 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19742) );
  AOI22_X1 U19639 ( .A1(n16528), .A2(n18722), .B1(n19742), .B2(n16529), .ZN(
        U365) );
  INV_X1 U19640 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18758) );
  INV_X1 U19641 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19762) );
  AOI22_X1 U19642 ( .A1(n16528), .A2(n18758), .B1(n19762), .B2(n16529), .ZN(
        U366) );
  INV_X1 U19643 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18757) );
  INV_X1 U19644 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19761) );
  AOI22_X1 U19645 ( .A1(n16528), .A2(n18757), .B1(n19761), .B2(n16529), .ZN(
        U367) );
  INV_X1 U19646 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18755) );
  INV_X1 U19647 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19759) );
  AOI22_X1 U19648 ( .A1(n16528), .A2(n18755), .B1(n19759), .B2(n16529), .ZN(
        U368) );
  INV_X1 U19649 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18752) );
  INV_X1 U19650 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19758) );
  AOI22_X1 U19651 ( .A1(n16528), .A2(n18752), .B1(n19758), .B2(n16529), .ZN(
        U369) );
  INV_X1 U19652 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18751) );
  INV_X1 U19653 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19756) );
  AOI22_X1 U19654 ( .A1(n16528), .A2(n18751), .B1(n19756), .B2(n16529), .ZN(
        U370) );
  INV_X1 U19655 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18749) );
  INV_X1 U19656 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19755) );
  AOI22_X1 U19657 ( .A1(n16528), .A2(n18749), .B1(n19755), .B2(n16529), .ZN(
        U371) );
  INV_X1 U19658 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18746) );
  INV_X1 U19659 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19754) );
  AOI22_X1 U19660 ( .A1(n16528), .A2(n18746), .B1(n19754), .B2(n16529), .ZN(
        U372) );
  INV_X1 U19661 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18745) );
  INV_X1 U19662 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19753) );
  AOI22_X1 U19663 ( .A1(n16528), .A2(n18745), .B1(n19753), .B2(n16529), .ZN(
        U373) );
  INV_X1 U19664 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18743) );
  INV_X1 U19665 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19752) );
  AOI22_X1 U19666 ( .A1(n16528), .A2(n18743), .B1(n19752), .B2(n16529), .ZN(
        U374) );
  INV_X1 U19667 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18741) );
  INV_X1 U19668 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19751) );
  AOI22_X1 U19669 ( .A1(n16528), .A2(n18741), .B1(n19751), .B2(n16529), .ZN(
        U375) );
  INV_X1 U19670 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18719) );
  INV_X1 U19671 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19741) );
  AOI22_X1 U19672 ( .A1(n16528), .A2(n18719), .B1(n19741), .B2(n16529), .ZN(
        U376) );
  INV_X1 U19673 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18716) );
  NOR2_X1 U19674 ( .A1(n18705), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18707) );
  OAI22_X1 U19675 ( .A1(n18716), .A2(n18707), .B1(n18705), .B2(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18701) );
  INV_X1 U19676 ( .A(n18701), .ZN(n18702) );
  AOI21_X1 U19677 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18702), .ZN(n16530) );
  INV_X1 U19678 ( .A(n16530), .ZN(P3_U2633) );
  NAND2_X1 U19679 ( .A1(n18688), .A2(n18794), .ZN(n16534) );
  NOR2_X1 U19680 ( .A1(n17416), .A2(n16531), .ZN(n16532) );
  OAI21_X1 U19681 ( .B1(n16532), .B2(n17417), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16533) );
  OAI21_X1 U19682 ( .B1(n16534), .B2(n18690), .A(n16533), .ZN(P3_U2634) );
  INV_X1 U19683 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18718) );
  AOI21_X1 U19684 ( .B1(n18716), .B2(n18718), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16535) );
  AOI22_X1 U19685 ( .A1(n18786), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16535), 
        .B2(n18851), .ZN(P3_U2635) );
  OAI21_X1 U19686 ( .B1(n18703), .B2(BS16), .A(n18702), .ZN(n18788) );
  OAI21_X1 U19687 ( .B1(n18702), .B2(n18841), .A(n18788), .ZN(P3_U2636) );
  AOI211_X1 U19688 ( .C1(n17418), .C2(n16537), .A(n16536), .B(n18622), .ZN(
        n18628) );
  NOR2_X1 U19689 ( .A1(n18628), .A2(n18839), .ZN(n18833) );
  INV_X1 U19690 ( .A(n16538), .ZN(n16539) );
  OAI21_X1 U19691 ( .B1(n18833), .B2(n18175), .A(n16539), .ZN(P3_U2637) );
  NOR4_X1 U19692 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16543) );
  NOR4_X1 U19693 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16542) );
  NOR4_X1 U19694 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16541) );
  NOR4_X1 U19695 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16540) );
  NAND4_X1 U19696 ( .A1(n16543), .A2(n16542), .A3(n16541), .A4(n16540), .ZN(
        n16549) );
  NOR4_X1 U19697 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_3__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n16547) );
  AOI211_X1 U19698 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_13__SCAN_IN), .B(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16546) );
  NOR4_X1 U19699 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A3(P3_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16545) );
  NOR4_X1 U19700 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n16544) );
  NAND4_X1 U19701 ( .A1(n16547), .A2(n16546), .A3(n16545), .A4(n16544), .ZN(
        n16548) );
  NOR2_X1 U19702 ( .A1(n16549), .A2(n16548), .ZN(n18831) );
  INV_X1 U19703 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16551) );
  NOR3_X1 U19704 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16552) );
  OAI21_X1 U19705 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16552), .A(n18831), .ZN(
        n16550) );
  OAI21_X1 U19706 ( .B1(n18831), .B2(n16551), .A(n16550), .ZN(P3_U2638) );
  INV_X1 U19707 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16554) );
  NOR2_X1 U19708 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18825) );
  OAI21_X1 U19709 ( .B1(n16552), .B2(n18825), .A(n18831), .ZN(n16553) );
  OAI21_X1 U19710 ( .B1(n18831), .B2(n16554), .A(n16553), .ZN(P3_U2639) );
  INV_X1 U19711 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18782) );
  INV_X1 U19712 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18769) );
  INV_X1 U19713 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18764) );
  NOR3_X1 U19714 ( .A1(n16720), .A2(n16556), .A3(n16555), .ZN(n16557) );
  NAND3_X1 U19715 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .A3(n16557), .ZN(n16656) );
  NOR2_X1 U19716 ( .A1(n18764), .A2(n16656), .ZN(n16654) );
  NAND2_X1 U19717 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16654), .ZN(n16635) );
  NOR2_X1 U19718 ( .A1(n18769), .A2(n16635), .ZN(n16619) );
  NAND2_X1 U19719 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16619), .ZN(n16568) );
  NAND4_X1 U19720 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16614), .ZN(n16571) );
  NOR3_X1 U19721 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18782), .A3(n16571), 
        .ZN(n16558) );
  AOI21_X1 U19722 ( .B1(n16878), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16558), .ZN(
        n16577) );
  NAND2_X1 U19723 ( .A1(n16660), .A2(n16950), .ZN(n16659) );
  NAND2_X1 U19724 ( .A1(n16631), .A2(n16643), .ZN(n16621) );
  INV_X1 U19725 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16616) );
  NAND2_X1 U19726 ( .A1(n16620), .A2(n16616), .ZN(n16615) );
  NOR2_X1 U19727 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16615), .ZN(n16600) );
  INV_X1 U19728 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n20863) );
  NAND2_X1 U19729 ( .A1(n16600), .A2(n20863), .ZN(n16579) );
  NOR2_X1 U19730 ( .A1(n16916), .A2(n16579), .ZN(n16586) );
  INV_X1 U19731 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16575) );
  INV_X1 U19732 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17503) );
  NAND2_X1 U19733 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17512), .ZN(
        n16565) );
  NOR3_X1 U19734 ( .A1(n16561), .A2(n17503), .A3(n16565), .ZN(n16562) );
  NAND2_X1 U19735 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16562), .ZN(
        n16560) );
  AOI21_X1 U19736 ( .B1(n17471), .B2(n16560), .A(n16559), .ZN(n17474) );
  OAI21_X1 U19737 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16562), .A(
        n16560), .ZN(n17497) );
  INV_X1 U19738 ( .A(n17497), .ZN(n16611) );
  NOR2_X1 U19739 ( .A1(n16561), .A2(n16565), .ZN(n17468) );
  INV_X1 U19740 ( .A(n17468), .ZN(n16563) );
  AOI21_X1 U19741 ( .B1(n17503), .B2(n16563), .A(n16562), .ZN(n17505) );
  INV_X1 U19742 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17527) );
  NOR2_X1 U19743 ( .A1(n17527), .A2(n16565), .ZN(n16564) );
  OAI21_X1 U19744 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16564), .A(
        n16563), .ZN(n17515) );
  INV_X1 U19745 ( .A(n17515), .ZN(n16634) );
  AOI21_X1 U19746 ( .B1(n17527), .B2(n16565), .A(n16564), .ZN(n17533) );
  OAI21_X1 U19747 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17513), .A(
        n16565), .ZN(n16566) );
  INV_X1 U19748 ( .A(n16566), .ZN(n17540) );
  NOR2_X1 U19749 ( .A1(n16567), .A2(n9919), .ZN(n16653) );
  NOR2_X1 U19750 ( .A1(n16634), .A2(n16633), .ZN(n16632) );
  NOR2_X1 U19751 ( .A1(n16632), .A2(n9919), .ZN(n16623) );
  NOR2_X1 U19752 ( .A1(n17505), .A2(n16623), .ZN(n16622) );
  NOR2_X1 U19753 ( .A1(n16622), .A2(n9919), .ZN(n16610) );
  NOR2_X1 U19754 ( .A1(n16591), .A2(n16590), .ZN(n16589) );
  NOR2_X1 U19755 ( .A1(n16589), .A2(n9919), .ZN(n16580) );
  NOR2_X1 U19756 ( .A1(n9919), .A2(n18694), .ZN(n16877) );
  INV_X1 U19757 ( .A(n16877), .ZN(n16908) );
  NOR3_X1 U19758 ( .A1(n16581), .A2(n16580), .A3(n16908), .ZN(n16574) );
  NAND3_X1 U19759 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16570) );
  NAND2_X1 U19760 ( .A1(n16869), .A2(n16568), .ZN(n16569) );
  NAND2_X1 U19761 ( .A1(n16807), .A2(n16569), .ZN(n16608) );
  AOI21_X1 U19762 ( .B1(n16869), .B2(n16570), .A(n16608), .ZN(n16599) );
  NOR2_X1 U19763 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16571), .ZN(n16584) );
  INV_X1 U19764 ( .A(n16584), .ZN(n16572) );
  AOI21_X1 U19765 ( .B1(n16599), .B2(n16572), .A(n18779), .ZN(n16573) );
  AOI211_X1 U19766 ( .C1(n16586), .C2(n16575), .A(n16574), .B(n16573), .ZN(
        n16576) );
  OAI211_X1 U19767 ( .C1(n16578), .C2(n16907), .A(n16577), .B(n16576), .ZN(
        P3_U2640) );
  NAND2_X1 U19768 ( .A1(n16881), .A2(n16579), .ZN(n16595) );
  XOR2_X1 U19769 ( .A(n16581), .B(n16580), .Z(n16585) );
  INV_X1 U19770 ( .A(n18694), .ZN(n16851) );
  OAI22_X1 U19771 ( .A1(n16599), .A2(n18782), .B1(n16582), .B2(n16907), .ZN(
        n16583) );
  AOI211_X1 U19772 ( .C1(n16585), .C2(n16851), .A(n16584), .B(n16583), .ZN(
        n16588) );
  OAI21_X1 U19773 ( .B1(n16878), .B2(n16586), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16587) );
  INV_X1 U19774 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18777) );
  AOI211_X1 U19775 ( .C1(n16591), .C2(n16590), .A(n16589), .B(n18694), .ZN(
        n16594) );
  NAND3_X1 U19776 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16614), .ZN(n16592) );
  OAI22_X1 U19777 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16592), .B1(n9925), 
        .B2(n16907), .ZN(n16593) );
  AOI211_X1 U19778 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16878), .A(n16594), .B(
        n16593), .ZN(n16598) );
  INV_X1 U19779 ( .A(n16595), .ZN(n16596) );
  OAI21_X1 U19780 ( .B1(n16600), .B2(n20863), .A(n16596), .ZN(n16597) );
  OAI211_X1 U19781 ( .C1(n16599), .C2(n18777), .A(n16598), .B(n16597), .ZN(
        P3_U2642) );
  AOI22_X1 U19782 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16879), .B1(
        n16878), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16607) );
  AOI211_X1 U19783 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16615), .A(n16600), .B(
        n16916), .ZN(n16603) );
  AOI211_X1 U19784 ( .C1(n17474), .C2(n16601), .A(n9656), .B(n18694), .ZN(
        n16602) );
  AOI211_X1 U19785 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16608), .A(n16603), 
        .B(n16602), .ZN(n16606) );
  NAND2_X1 U19786 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n16604) );
  OAI211_X1 U19787 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16614), .B(n16604), .ZN(n16605) );
  NAND3_X1 U19788 ( .A1(n16607), .A2(n16606), .A3(n16605), .ZN(P3_U2643) );
  INV_X1 U19789 ( .A(n16608), .ZN(n16630) );
  INV_X1 U19790 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18773) );
  AOI211_X1 U19791 ( .C1(n16611), .C2(n16610), .A(n16609), .B(n18694), .ZN(
        n16613) );
  OAI22_X1 U19792 ( .A1(n17470), .A2(n16907), .B1(n16917), .B2(n16616), .ZN(
        n16612) );
  AOI211_X1 U19793 ( .C1(n16614), .C2(n18773), .A(n16613), .B(n16612), .ZN(
        n16618) );
  OAI211_X1 U19794 ( .C1(n16620), .C2(n16616), .A(n16881), .B(n16615), .ZN(
        n16617) );
  OAI211_X1 U19795 ( .C1(n16630), .C2(n18773), .A(n16618), .B(n16617), .ZN(
        P3_U2644) );
  AOI21_X1 U19796 ( .B1(n16869), .B2(n16619), .A(P3_REIP_REG_26__SCAN_IN), 
        .ZN(n16629) );
  AOI211_X1 U19797 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16621), .A(n16620), .B(
        n16916), .ZN(n16627) );
  AOI211_X1 U19798 ( .C1(n17505), .C2(n16623), .A(n16622), .B(n18694), .ZN(
        n16626) );
  OAI22_X1 U19799 ( .A1(n17503), .A2(n16907), .B1(n16917), .B2(n16624), .ZN(
        n16625) );
  NOR3_X1 U19800 ( .A1(n16627), .A2(n16626), .A3(n16625), .ZN(n16628) );
  OAI21_X1 U19801 ( .B1(n16630), .B2(n16629), .A(n16628), .ZN(P3_U2645) );
  OR2_X1 U19802 ( .A1(n16916), .A2(n16631), .ZN(n16645) );
  AOI21_X1 U19803 ( .B1(n16881), .B2(n16631), .A(n16878), .ZN(n16642) );
  AOI211_X1 U19804 ( .C1(n16634), .C2(n16633), .A(n16632), .B(n18694), .ZN(
        n16640) );
  NOR2_X1 U19805 ( .A1(n16909), .A2(n16635), .ZN(n16638) );
  INV_X1 U19806 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18766) );
  OAI21_X1 U19807 ( .B1(n16654), .B2(n16909), .A(n16807), .ZN(n16651) );
  AOI21_X1 U19808 ( .B1(n16869), .B2(n18766), .A(n16651), .ZN(n16636) );
  INV_X1 U19809 ( .A(n16636), .ZN(n16637) );
  MUX2_X1 U19810 ( .A(n16638), .B(n16637), .S(P3_REIP_REG_25__SCAN_IN), .Z(
        n16639) );
  AOI211_X1 U19811 ( .C1(n16879), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16640), .B(n16639), .ZN(n16641) );
  OAI221_X1 U19812 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n16645), .C1(n16643), 
        .C2(n16642), .A(n16641), .ZN(P3_U2646) );
  NOR2_X1 U19813 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16909), .ZN(n16644) );
  AOI22_X1 U19814 ( .A1(n16878), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16654), 
        .B2(n16644), .ZN(n16650) );
  AOI21_X1 U19815 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16659), .A(n16645), .ZN(
        n16648) );
  AOI211_X1 U19816 ( .C1(n17533), .C2(n16646), .A(n9673), .B(n18694), .ZN(
        n16647) );
  AOI211_X1 U19817 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16651), .A(n16648), 
        .B(n16647), .ZN(n16649) );
  OAI211_X1 U19818 ( .C1(n17527), .C2(n16907), .A(n16650), .B(n16649), .ZN(
        P3_U2647) );
  INV_X1 U19819 ( .A(n16651), .ZN(n16663) );
  AOI211_X1 U19820 ( .C1(n17540), .C2(n16653), .A(n16652), .B(n18694), .ZN(
        n16658) );
  OR2_X1 U19821 ( .A1(n16909), .A2(n16654), .ZN(n16655) );
  OAI22_X1 U19822 ( .A1(n16917), .A2(n16950), .B1(n16656), .B2(n16655), .ZN(
        n16657) );
  AOI211_X1 U19823 ( .C1(n16879), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16658), .B(n16657), .ZN(n16662) );
  OAI211_X1 U19824 ( .C1(n16660), .C2(n16950), .A(n16881), .B(n16659), .ZN(
        n16661) );
  OAI211_X1 U19825 ( .C1(n16663), .C2(n18764), .A(n16662), .B(n16661), .ZN(
        P3_U2648) );
  INV_X1 U19826 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18760) );
  AOI211_X1 U19827 ( .C1(n17566), .C2(n9697), .A(n16664), .B(n18694), .ZN(
        n16669) );
  OAI211_X1 U19828 ( .C1(n16674), .C2(n16667), .A(n16881), .B(n16665), .ZN(
        n16666) );
  OAI21_X1 U19829 ( .B1(n16667), .B2(n16917), .A(n16666), .ZN(n16668) );
  AOI211_X1 U19830 ( .C1(n16879), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16669), .B(n16668), .ZN(n16670) );
  OAI221_X1 U19831 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16671), .C1(n18760), 
        .C2(n16679), .A(n16670), .ZN(P3_U2650) );
  NAND3_X1 U19832 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .A3(n16691), .ZN(n16680) );
  AOI211_X1 U19833 ( .C1(n17576), .C2(n16673), .A(n16672), .B(n18694), .ZN(
        n16677) );
  AOI211_X1 U19834 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16684), .A(n16674), .B(
        n16916), .ZN(n16676) );
  OAI22_X1 U19835 ( .A1(n17574), .A2(n16907), .B1(n16917), .B2(n16982), .ZN(
        n16675) );
  NOR3_X1 U19836 ( .A1(n16677), .A2(n16676), .A3(n16675), .ZN(n16678) );
  OAI221_X1 U19837 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(n16680), .C1(n18759), 
        .C2(n16679), .A(n16678), .ZN(P3_U2651) );
  NAND2_X1 U19838 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16691), .ZN(n16690) );
  OAI21_X1 U19839 ( .B1(n18754), .B2(n16701), .A(n16922), .ZN(n16700) );
  NOR2_X1 U19840 ( .A1(n17602), .A2(n17588), .ZN(n16692) );
  OAI21_X1 U19841 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16692), .A(
        n17549), .ZN(n17589) );
  INV_X1 U19842 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17645) );
  NOR2_X1 U19843 ( .A1(n17645), .A2(n17629), .ZN(n16727) );
  INV_X1 U19844 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16918) );
  AND2_X1 U19845 ( .A1(n16727), .A2(n16918), .ZN(n16728) );
  AOI21_X1 U19846 ( .B1(n16692), .B2(n16728), .A(n9919), .ZN(n16681) );
  INV_X1 U19847 ( .A(n16681), .ZN(n16683) );
  OAI21_X1 U19848 ( .B1(n17589), .B2(n16683), .A(n16851), .ZN(n16682) );
  AOI21_X1 U19849 ( .B1(n17589), .B2(n16683), .A(n16682), .ZN(n16688) );
  OAI211_X1 U19850 ( .C1(n16694), .C2(n16686), .A(n16881), .B(n16684), .ZN(
        n16685) );
  OAI211_X1 U19851 ( .C1(n16917), .C2(n16686), .A(n18122), .B(n16685), .ZN(
        n16687) );
  AOI211_X1 U19852 ( .C1(n16879), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16688), .B(n16687), .ZN(n16689) );
  OAI221_X1 U19853 ( .B1(P3_REIP_REG_19__SCAN_IN), .B2(n16690), .C1(n18756), 
        .C2(n16700), .A(n16689), .ZN(P3_U2652) );
  NOR2_X1 U19854 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16691), .ZN(n16699) );
  AOI22_X1 U19855 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16879), .B1(
        n16878), .B2(P3_EBX_REG_18__SCAN_IN), .ZN(n16698) );
  AOI21_X1 U19856 ( .B1(n17602), .B2(n17588), .A(n16692), .ZN(n17605) );
  XNOR2_X1 U19857 ( .A(n17605), .B(n16693), .ZN(n16696) );
  AOI211_X1 U19858 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16702), .A(n16694), .B(
        n16916), .ZN(n16695) );
  AOI211_X1 U19859 ( .C1(n16851), .C2(n16696), .A(n18165), .B(n16695), .ZN(
        n16697) );
  OAI211_X1 U19860 ( .C1(n16700), .C2(n16699), .A(n16698), .B(n16697), .ZN(
        P3_U2653) );
  NAND2_X1 U19861 ( .A1(n16922), .A2(n16701), .ZN(n16711) );
  INV_X1 U19862 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18753) );
  INV_X1 U19863 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18750) );
  INV_X1 U19864 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18748) );
  NOR4_X1 U19865 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n18750), .A3(n18748), 
        .A4(n16726), .ZN(n16706) );
  OAI211_X1 U19866 ( .C1(n16716), .C2(n16704), .A(n16881), .B(n16702), .ZN(
        n16703) );
  OAI211_X1 U19867 ( .C1(n16917), .C2(n16704), .A(n18122), .B(n16703), .ZN(
        n16705) );
  AOI211_X1 U19868 ( .C1(n16879), .C2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16706), .B(n16705), .ZN(n16710) );
  OAI21_X1 U19869 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16712), .A(
        n17588), .ZN(n17614) );
  INV_X1 U19870 ( .A(n17614), .ZN(n16708) );
  AOI21_X1 U19871 ( .B1(n16918), .B2(n16712), .A(n9919), .ZN(n16707) );
  INV_X1 U19872 ( .A(n16707), .ZN(n16715) );
  OAI221_X1 U19873 ( .B1(n16708), .B2(n16707), .C1(n17614), .C2(n16715), .A(
        n16851), .ZN(n16709) );
  OAI211_X1 U19874 ( .C1(n16711), .C2(n18753), .A(n16710), .B(n16709), .ZN(
        P3_U2654) );
  NAND2_X1 U19875 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n18750), .ZN(n16725) );
  INV_X1 U19876 ( .A(n16712), .ZN(n16713) );
  OAI21_X1 U19877 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16727), .A(
        n16713), .ZN(n17631) );
  NAND2_X1 U19878 ( .A1(n16851), .A2(n9919), .ZN(n16896) );
  OAI21_X1 U19879 ( .B1(n16728), .B2(n17631), .A(n16851), .ZN(n16714) );
  AOI22_X1 U19880 ( .A1(n17631), .A2(n16715), .B1(n16896), .B2(n16714), .ZN(
        n16719) );
  AOI211_X1 U19881 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16734), .A(n16716), .B(
        n16916), .ZN(n16718) );
  INV_X1 U19882 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17632) );
  OAI22_X1 U19883 ( .A1(n17632), .A2(n16907), .B1(n16917), .B2(n17050), .ZN(
        n16717) );
  NOR4_X1 U19884 ( .A1(n18165), .A2(n16719), .A3(n16718), .A4(n16717), .ZN(
        n16724) );
  NOR2_X1 U19885 ( .A1(n16919), .A2(n16720), .ZN(n16721) );
  NOR2_X1 U19886 ( .A1(n16722), .A2(n16721), .ZN(n16741) );
  NOR2_X1 U19887 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16726), .ZN(n16732) );
  OAI21_X1 U19888 ( .B1(n16741), .B2(n16732), .A(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n16723) );
  OAI211_X1 U19889 ( .C1(n16726), .C2(n16725), .A(n16724), .B(n16723), .ZN(
        P3_U2655) );
  AOI21_X1 U19890 ( .B1(n17645), .B2(n17629), .A(n16727), .ZN(n17648) );
  NOR3_X1 U19891 ( .A1(n17648), .A2(n16728), .A3(n16908), .ZN(n16729) );
  AOI211_X1 U19892 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16879), .A(
        n18165), .B(n16729), .ZN(n16730) );
  OAI21_X1 U19893 ( .B1(n16917), .B2(n17064), .A(n16730), .ZN(n16731) );
  AOI211_X1 U19894 ( .C1(n16741), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16732), 
        .B(n16731), .ZN(n16737) );
  INV_X1 U19895 ( .A(n17629), .ZN(n16733) );
  AOI21_X1 U19896 ( .B1(n16876), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n18694), .ZN(n16911) );
  OAI211_X1 U19897 ( .C1(n16733), .C2(n9919), .A(n17648), .B(n16911), .ZN(
        n16736) );
  OAI211_X1 U19898 ( .C1(n16739), .C2(n17064), .A(n16881), .B(n16734), .ZN(
        n16735) );
  NAND3_X1 U19899 ( .A1(n16737), .A2(n16736), .A3(n16735), .ZN(P3_U2656) );
  NOR2_X1 U19900 ( .A1(n16912), .A2(n17678), .ZN(n17677) );
  INV_X1 U19901 ( .A(n17677), .ZN(n16773) );
  NOR2_X1 U19902 ( .A1(n17680), .A2(n16773), .ZN(n16748) );
  OAI21_X1 U19903 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16748), .A(
        n17629), .ZN(n17669) );
  AOI21_X1 U19904 ( .B1(n16748), .B2(n16918), .A(n9919), .ZN(n16738) );
  XOR2_X1 U19905 ( .A(n17669), .B(n16738), .Z(n16747) );
  AOI211_X1 U19906 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16758), .A(n16739), .B(
        n16916), .ZN(n16745) );
  INV_X1 U19907 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17076) );
  INV_X1 U19908 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18744) );
  NAND2_X1 U19909 ( .A1(n16869), .A2(n16740), .ZN(n16754) );
  NOR2_X1 U19910 ( .A1(n18744), .A2(n16754), .ZN(n16742) );
  OAI21_X1 U19911 ( .B1(P3_REIP_REG_14__SCAN_IN), .B2(n16742), .A(n16741), 
        .ZN(n16743) );
  OAI211_X1 U19912 ( .C1(n16917), .C2(n17076), .A(n18122), .B(n16743), .ZN(
        n16744) );
  AOI211_X1 U19913 ( .C1(n16879), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16745), .B(n16744), .ZN(n16746) );
  OAI21_X1 U19914 ( .B1(n18694), .B2(n16747), .A(n16746), .ZN(P3_U2657) );
  AOI21_X1 U19915 ( .B1(n16869), .B2(n16770), .A(n16919), .ZN(n16776) );
  OAI21_X1 U19916 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n16909), .A(n16776), 
        .ZN(n16757) );
  NOR2_X1 U19917 ( .A1(n17691), .A2(n16773), .ZN(n16749) );
  INV_X1 U19918 ( .A(n16748), .ZN(n16752) );
  OAI21_X1 U19919 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16749), .A(
        n16752), .ZN(n17683) );
  OAI21_X1 U19920 ( .B1(n9919), .B2(n16751), .A(n16911), .ZN(n16750) );
  OAI22_X1 U19921 ( .A1(n16751), .A2(n16907), .B1(n17683), .B2(n16750), .ZN(
        n16756) );
  OAI211_X1 U19922 ( .C1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n16752), .A(
        n16877), .B(n17683), .ZN(n16753) );
  OAI211_X1 U19923 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16754), .A(n18122), 
        .B(n16753), .ZN(n16755) );
  AOI211_X1 U19924 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16757), .A(n16756), 
        .B(n16755), .ZN(n16760) );
  OAI211_X1 U19925 ( .C1(n16762), .C2(n16761), .A(n16881), .B(n16758), .ZN(
        n16759) );
  OAI211_X1 U19926 ( .C1(n16761), .C2(n16917), .A(n16760), .B(n16759), .ZN(
        P3_U2658) );
  NAND2_X1 U19927 ( .A1(n16869), .A2(n18742), .ZN(n16769) );
  AOI21_X1 U19928 ( .B1(n16878), .B2(P3_EBX_REG_12__SCAN_IN), .A(n18165), .ZN(
        n16768) );
  AOI211_X1 U19929 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16779), .A(n16762), .B(
        n16916), .ZN(n16766) );
  AOI22_X1 U19930 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16773), .B1(
        n17677), .B2(n17691), .ZN(n17695) );
  OAI21_X1 U19931 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16773), .A(
        n16876), .ZN(n16763) );
  XNOR2_X1 U19932 ( .A(n17695), .B(n16763), .ZN(n16764) );
  OAI22_X1 U19933 ( .A1(n18694), .A2(n16764), .B1(n18742), .B2(n16776), .ZN(
        n16765) );
  AOI211_X1 U19934 ( .C1(n16879), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16766), .B(n16765), .ZN(n16767) );
  OAI211_X1 U19935 ( .C1(n16770), .C2(n16769), .A(n16768), .B(n16767), .ZN(
        P3_U2659) );
  INV_X1 U19936 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16782) );
  AOI21_X1 U19937 ( .B1(n16869), .B2(n16771), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16777) );
  INV_X1 U19938 ( .A(n17772), .ZN(n17771) );
  NAND2_X1 U19939 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17771), .ZN(
        n16833) );
  INV_X1 U19940 ( .A(n16833), .ZN(n16845) );
  NAND2_X1 U19941 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16845), .ZN(
        n16831) );
  NOR2_X1 U19942 ( .A1(n16772), .A2(n16831), .ZN(n16783) );
  AOI21_X1 U19943 ( .B1(n16783), .B2(n16918), .A(n9919), .ZN(n16774) );
  OAI21_X1 U19944 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16783), .A(
        n16773), .ZN(n17706) );
  XOR2_X1 U19945 ( .A(n16774), .B(n17706), .Z(n16775) );
  OAI22_X1 U19946 ( .A1(n16777), .A2(n16776), .B1(n18694), .B2(n16775), .ZN(
        n16778) );
  AOI211_X1 U19947 ( .C1(n16878), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18165), .B(
        n16778), .ZN(n16781) );
  OAI211_X1 U19948 ( .C1(n16789), .C2(n17094), .A(n16881), .B(n16779), .ZN(
        n16780) );
  OAI211_X1 U19949 ( .C1(n16907), .C2(n16782), .A(n16781), .B(n16780), .ZN(
        P3_U2660) );
  INV_X1 U19950 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18736) );
  INV_X1 U19951 ( .A(n16808), .ZN(n16798) );
  AOI221_X1 U19952 ( .B1(n18736), .B2(n16869), .C1(n16798), .C2(n16869), .A(
        n16919), .ZN(n16797) );
  AOI22_X1 U19953 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16879), .B1(
        n16878), .B2(P3_EBX_REG_10__SCAN_IN), .ZN(n16794) );
  INV_X1 U19954 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16784) );
  NOR2_X1 U19955 ( .A1(n17730), .A2(n16831), .ZN(n16785) );
  INV_X1 U19956 ( .A(n16785), .ZN(n16795) );
  AOI21_X1 U19957 ( .B1(n16784), .B2(n16795), .A(n16783), .ZN(n17721) );
  AOI21_X1 U19958 ( .B1(n16785), .B2(n16918), .A(n9919), .ZN(n16787) );
  OAI21_X1 U19959 ( .B1(n17721), .B2(n16787), .A(n16851), .ZN(n16786) );
  AOI21_X1 U19960 ( .B1(n17721), .B2(n16787), .A(n16786), .ZN(n16792) );
  NOR3_X1 U19961 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n16909), .A3(n16788), 
        .ZN(n16791) );
  AOI211_X1 U19962 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16801), .A(n16789), .B(
        n16916), .ZN(n16790) );
  NOR4_X1 U19963 ( .A1(n18165), .A2(n16792), .A3(n16791), .A4(n16790), .ZN(
        n16793) );
  OAI211_X1 U19964 ( .C1(n16797), .C2(n18738), .A(n16794), .B(n16793), .ZN(
        P3_U2661) );
  AOI22_X1 U19965 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16879), .B1(
        n16878), .B2(P3_EBX_REG_9__SCAN_IN), .ZN(n16804) );
  NOR2_X1 U19966 ( .A1(n17745), .A2(n16831), .ZN(n16810) );
  OAI21_X1 U19967 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16810), .A(
        n16795), .ZN(n17733) );
  AOI21_X1 U19968 ( .B1(n16810), .B2(n16918), .A(n9919), .ZN(n16796) );
  XNOR2_X1 U19969 ( .A(n17733), .B(n16796), .ZN(n16800) );
  AOI221_X1 U19970 ( .B1(n16909), .B2(n18736), .C1(n16798), .C2(n18736), .A(
        n16797), .ZN(n16799) );
  AOI21_X1 U19971 ( .B1(n16800), .B2(n16851), .A(n16799), .ZN(n16803) );
  OAI211_X1 U19972 ( .C1(n16805), .C2(n17123), .A(n16881), .B(n16801), .ZN(
        n16802) );
  NAND4_X1 U19973 ( .A1(n16804), .A2(n16803), .A3(n18122), .A4(n16802), .ZN(
        P3_U2662) );
  INV_X1 U19974 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16820) );
  AOI211_X1 U19975 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16823), .A(n16805), .B(
        n16916), .ZN(n16806) );
  AOI211_X1 U19976 ( .C1(n16878), .C2(P3_EBX_REG_8__SCAN_IN), .A(n18165), .B(
        n16806), .ZN(n16819) );
  OAI21_X1 U19977 ( .B1(n16808), .B2(n16909), .A(n16807), .ZN(n16817) );
  NAND3_X1 U19978 ( .A1(n16869), .A2(P3_REIP_REG_5__SCAN_IN), .A3(n16847), 
        .ZN(n16843) );
  NOR2_X1 U19979 ( .A1(n16809), .A2(n16843), .ZN(n16816) );
  INV_X1 U19980 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16822) );
  NOR2_X1 U19981 ( .A1(n16822), .A2(n16831), .ZN(n16821) );
  INV_X1 U19982 ( .A(n16810), .ZN(n16811) );
  OAI21_X1 U19983 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16821), .A(
        n16811), .ZN(n17748) );
  NAND2_X1 U19984 ( .A1(n16918), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16891) );
  INV_X1 U19985 ( .A(n16891), .ZN(n16871) );
  NAND2_X1 U19986 ( .A1(n17746), .A2(n16871), .ZN(n16812) );
  OAI21_X1 U19987 ( .B1(n16822), .B2(n16812), .A(n16876), .ZN(n16814) );
  OAI21_X1 U19988 ( .B1(n17748), .B2(n16814), .A(n16851), .ZN(n16813) );
  AOI21_X1 U19989 ( .B1(n17748), .B2(n16814), .A(n16813), .ZN(n16815) );
  AOI221_X1 U19990 ( .B1(n16817), .B2(P3_REIP_REG_8__SCAN_IN), .C1(n16816), 
        .C2(n18734), .A(n16815), .ZN(n16818) );
  OAI211_X1 U19991 ( .C1(n16820), .C2(n16907), .A(n16819), .B(n16818), .ZN(
        P3_U2663) );
  AOI21_X1 U19992 ( .B1(n17746), .B2(n16871), .A(n9919), .ZN(n16835) );
  AOI21_X1 U19993 ( .B1(n16822), .B2(n16831), .A(n16821), .ZN(n17762) );
  XNOR2_X1 U19994 ( .A(n16835), .B(n17762), .ZN(n16830) );
  OAI211_X1 U19995 ( .C1(n16834), .C2(n17167), .A(n16881), .B(n16823), .ZN(
        n16824) );
  OAI211_X1 U19996 ( .C1(n16917), .C2(n17167), .A(n18122), .B(n16824), .ZN(
        n16828) );
  XNOR2_X1 U19997 ( .A(P3_REIP_REG_7__SCAN_IN), .B(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n16826) );
  AOI21_X1 U19998 ( .B1(n16869), .B2(n16825), .A(n16919), .ZN(n16848) );
  INV_X1 U19999 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18732) );
  OAI22_X1 U20000 ( .A1(n16843), .A2(n16826), .B1(n16848), .B2(n18732), .ZN(
        n16827) );
  AOI211_X1 U20001 ( .C1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n16879), .A(
        n16828), .B(n16827), .ZN(n16829) );
  OAI21_X1 U20002 ( .B1(n18694), .B2(n16830), .A(n16829), .ZN(P3_U2664) );
  INV_X1 U20003 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18730) );
  OAI21_X1 U20004 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16845), .A(
        n16831), .ZN(n17781) );
  INV_X1 U20005 ( .A(n17781), .ZN(n16841) );
  NAND2_X1 U20006 ( .A1(n16851), .A2(n16918), .ZN(n16832) );
  OAI21_X1 U20007 ( .B1(n16833), .B2(n16832), .A(n16896), .ZN(n16840) );
  AOI211_X1 U20008 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16853), .A(n16834), .B(
        n16916), .ZN(n16839) );
  AOI22_X1 U20009 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16879), .B1(
        n16878), .B2(P3_EBX_REG_6__SCAN_IN), .ZN(n16837) );
  NAND3_X1 U20010 ( .A1(n16851), .A2(n16835), .A3(n17781), .ZN(n16836) );
  NAND3_X1 U20011 ( .A1(n16837), .A2(n18122), .A3(n16836), .ZN(n16838) );
  AOI211_X1 U20012 ( .C1(n16841), .C2(n16840), .A(n16839), .B(n16838), .ZN(
        n16842) );
  OAI221_X1 U20013 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n16843), .C1(n18730), 
        .C2(n16848), .A(n16842), .ZN(P3_U2665) );
  AOI22_X1 U20014 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n16879), .B1(
        n16878), .B2(P3_EBX_REG_5__SCAN_IN), .ZN(n16857) );
  AOI21_X1 U20015 ( .B1(n17782), .B2(n16871), .A(n9919), .ZN(n16862) );
  INV_X1 U20016 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16846) );
  NAND2_X1 U20017 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17782), .ZN(
        n16858) );
  AOI21_X1 U20018 ( .B1(n16846), .B2(n16858), .A(n16845), .ZN(n17791) );
  XOR2_X1 U20019 ( .A(n16862), .B(n17791), .Z(n16852) );
  INV_X1 U20020 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18729) );
  NAND2_X1 U20021 ( .A1(n16869), .A2(n16847), .ZN(n16849) );
  AOI21_X1 U20022 ( .B1(n18729), .B2(n16849), .A(n16848), .ZN(n16850) );
  AOI21_X1 U20023 ( .B1(n16852), .B2(n16851), .A(n16850), .ZN(n16856) );
  OAI211_X1 U20024 ( .C1(n16859), .C2(n16854), .A(n16881), .B(n16853), .ZN(
        n16855) );
  NAND4_X1 U20025 ( .A1(n16857), .A2(n16856), .A3(n18122), .A4(n16855), .ZN(
        P3_U2666) );
  NOR2_X1 U20026 ( .A1(n16912), .A2(n17804), .ZN(n16872) );
  OAI21_X1 U20027 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16872), .A(
        n16858), .ZN(n17806) );
  NOR3_X1 U20028 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16909), .A3(n16863), .ZN(
        n16861) );
  AOI211_X1 U20029 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16880), .A(n16859), .B(
        n16916), .ZN(n16860) );
  AOI211_X1 U20030 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16878), .A(n16861), .B(
        n16860), .ZN(n16868) );
  NOR2_X1 U20031 ( .A1(n18185), .A2(n18855), .ZN(n16906) );
  INV_X1 U20032 ( .A(n16906), .ZN(n18857) );
  OAI221_X1 U20033 ( .B1(n18857), .B2(n9604), .C1(n18857), .C2(n18631), .A(
        n18122), .ZN(n16866) );
  NOR2_X1 U20034 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17804), .ZN(
        n17809) );
  AOI22_X1 U20035 ( .A1(n16871), .A2(n17809), .B1(n16862), .B2(n17806), .ZN(
        n16864) );
  AOI21_X1 U20036 ( .B1(n16869), .B2(n16863), .A(n16919), .ZN(n16887) );
  OAI22_X1 U20037 ( .A1(n16864), .A2(n18694), .B1(n18726), .B2(n16887), .ZN(
        n16865) );
  AOI211_X1 U20038 ( .C1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n16879), .A(
        n16866), .B(n16865), .ZN(n16867) );
  OAI211_X1 U20039 ( .C1(n17806), .C2(n16896), .A(n16868), .B(n16867), .ZN(
        P3_U2667) );
  INV_X1 U20040 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18720) );
  INV_X1 U20041 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18721) );
  NOR2_X1 U20042 ( .A1(n18720), .A2(n18721), .ZN(n16895) );
  AOI21_X1 U20043 ( .B1(n16869), .B2(n16895), .A(P3_REIP_REG_3__SCAN_IN), .ZN(
        n16888) );
  NOR2_X1 U20044 ( .A1(n12565), .A2(n18808), .ZN(n18652) );
  INV_X1 U20045 ( .A(n18652), .ZN(n18657) );
  NOR2_X1 U20046 ( .A1(n18821), .A2(n18657), .ZN(n18660) );
  OAI21_X1 U20047 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18660), .A(
        n9604), .ZN(n16870) );
  INV_X1 U20048 ( .A(n16870), .ZN(n18795) );
  NAND2_X1 U20049 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n16871), .ZN(
        n16875) );
  INV_X1 U20050 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16873) );
  NAND2_X1 U20051 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16889) );
  AOI21_X1 U20052 ( .B1(n16873), .B2(n16889), .A(n16872), .ZN(n17818) );
  INV_X1 U20053 ( .A(n17818), .ZN(n16874) );
  AOI211_X1 U20054 ( .C1(n16876), .C2(n16875), .A(n18694), .B(n16874), .ZN(
        n16885) );
  INV_X1 U20055 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17831) );
  OAI21_X1 U20056 ( .B1(n17831), .B2(n16891), .A(n16877), .ZN(n16890) );
  AOI22_X1 U20057 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n16879), .B1(
        n16878), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n16883) );
  OAI211_X1 U20058 ( .C1(n16893), .C2(n17183), .A(n16881), .B(n16880), .ZN(
        n16882) );
  OAI211_X1 U20059 ( .C1(n17818), .C2(n16890), .A(n16883), .B(n16882), .ZN(
        n16884) );
  AOI211_X1 U20060 ( .C1(n16906), .C2(n18795), .A(n16885), .B(n16884), .ZN(
        n16886) );
  OAI21_X1 U20061 ( .B1(n16888), .B2(n16887), .A(n16886), .ZN(P3_U2668) );
  AOI21_X1 U20062 ( .B1(n18650), .B2(n18808), .A(n18660), .ZN(n18804) );
  AOI22_X1 U20063 ( .A1(n16919), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n18804), 
        .B2(n16906), .ZN(n16902) );
  OAI21_X1 U20064 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16889), .ZN(n17827) );
  INV_X1 U20065 ( .A(n17827), .ZN(n16892) );
  AOI21_X1 U20066 ( .B1(n16892), .B2(n16891), .A(n16890), .ZN(n16900) );
  NAND2_X1 U20067 ( .A1(n17200), .A2(n17194), .ZN(n16894) );
  AOI211_X1 U20068 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16894), .A(n16893), .B(
        n16916), .ZN(n16899) );
  AOI211_X1 U20069 ( .C1(n18720), .C2(n18721), .A(n16895), .B(n16909), .ZN(
        n16898) );
  OAI22_X1 U20070 ( .A1(n17831), .A2(n16907), .B1(n17827), .B2(n16896), .ZN(
        n16897) );
  NOR4_X1 U20071 ( .A1(n16900), .A2(n16899), .A3(n16898), .A4(n16897), .ZN(
        n16901) );
  OAI211_X1 U20072 ( .C1(n16917), .C2(n16903), .A(n16902), .B(n16901), .ZN(
        P3_U2669) );
  OAI21_X1 U20073 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n16904), .ZN(n17195) );
  AND2_X1 U20074 ( .A1(n18650), .A2(n16905), .ZN(n18812) );
  AOI22_X1 U20075 ( .A1(n16919), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18812), 
        .B2(n16906), .ZN(n16915) );
  OAI21_X1 U20076 ( .B1(n16918), .B2(n16908), .A(n16907), .ZN(n16913) );
  OAI22_X1 U20077 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16909), .B1(n16917), 
        .B2(n17194), .ZN(n16910) );
  AOI221_X1 U20078 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16913), .C1(
        n16912), .C2(n16911), .A(n16910), .ZN(n16914) );
  OAI211_X1 U20079 ( .C1(n16916), .C2(n17195), .A(n16915), .B(n16914), .ZN(
        P3_U2670) );
  AOI21_X1 U20080 ( .B1(n16917), .B2(n16916), .A(n17200), .ZN(n16921) );
  NOR3_X1 U20081 ( .A1(n18817), .A2(n16919), .A3(n16918), .ZN(n16920) );
  AOI211_X1 U20082 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(n16922), .A(n16921), .B(
        n16920), .ZN(n16923) );
  OAI21_X1 U20083 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18857), .A(
        n16923), .ZN(P3_U2671) );
  OAI33_X1 U20084 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18225), .A3(n16926), 
        .B1(n16925), .B2(n17198), .B3(n16924), .ZN(P3_U2672) );
  NAND2_X1 U20085 ( .A1(n16928), .A2(n16927), .ZN(n16934) );
  NOR2_X1 U20086 ( .A1(n16935), .A2(n16929), .ZN(n16931) );
  XNOR2_X1 U20087 ( .A(n16931), .B(n16930), .ZN(n17215) );
  AOI22_X1 U20088 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16932), .B1(n17198), 
        .B2(n17215), .ZN(n16933) );
  OAI21_X1 U20089 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16934), .A(n16933), .ZN(
        P3_U2674) );
  OAI21_X1 U20090 ( .B1(n16937), .B2(n16936), .A(n16935), .ZN(n17227) );
  OAI211_X1 U20091 ( .C1(n9636), .C2(P3_EBX_REG_27__SCAN_IN), .A(n17192), .B(
        n16938), .ZN(n16939) );
  OAI21_X1 U20092 ( .B1(n17227), .B2(n17192), .A(n16939), .ZN(P3_U2676) );
  AOI21_X1 U20093 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17192), .A(n9637), .ZN(
        n16941) );
  XNOR2_X1 U20094 ( .A(n16940), .B(n16942), .ZN(n17232) );
  OAI22_X1 U20095 ( .A1(n9636), .A2(n16941), .B1(n17192), .B2(n17232), .ZN(
        P3_U2677) );
  AOI21_X1 U20096 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17192), .A(n16948), .ZN(
        n16945) );
  OAI21_X1 U20097 ( .B1(n16944), .B2(n16943), .A(n16942), .ZN(n17237) );
  OAI22_X1 U20098 ( .A1(n9637), .A2(n16945), .B1(n17192), .B2(n17237), .ZN(
        P3_U2678) );
  AOI21_X1 U20099 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17192), .A(n16956), .ZN(
        n16947) );
  XNOR2_X1 U20100 ( .A(n16946), .B(n16952), .ZN(n17242) );
  OAI22_X1 U20101 ( .A1(n16948), .A2(n16947), .B1(n17192), .B2(n17242), .ZN(
        P3_U2679) );
  OAI22_X1 U20102 ( .A1(n16950), .A2(n17198), .B1(n16949), .B2(n16968), .ZN(
        n16951) );
  INV_X1 U20103 ( .A(n16951), .ZN(n16955) );
  OAI21_X1 U20104 ( .B1(n16954), .B2(n16953), .A(n16952), .ZN(n17247) );
  OAI22_X1 U20105 ( .A1(n16956), .A2(n16955), .B1(n17192), .B2(n17247), .ZN(
        P3_U2680) );
  AOI22_X1 U20106 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16960) );
  AOI22_X1 U20107 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16959) );
  AOI22_X1 U20108 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16958) );
  AOI22_X1 U20109 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16957) );
  NAND4_X1 U20110 ( .A1(n16960), .A2(n16959), .A3(n16958), .A4(n16957), .ZN(
        n16966) );
  AOI22_X1 U20111 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16964) );
  AOI22_X1 U20112 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16963) );
  AOI22_X1 U20113 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16962) );
  AOI22_X1 U20114 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17142), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16961) );
  NAND4_X1 U20115 ( .A1(n16964), .A2(n16963), .A3(n16962), .A4(n16961), .ZN(
        n16965) );
  NOR2_X1 U20116 ( .A1(n16966), .A2(n16965), .ZN(n17249) );
  NAND3_X1 U20117 ( .A1(n16968), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17192), 
        .ZN(n16967) );
  OAI221_X1 U20118 ( .B1(n16968), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17192), 
        .C2(n17249), .A(n16967), .ZN(P3_U2681) );
  AOI22_X1 U20119 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16972) );
  AOI22_X1 U20120 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16971) );
  AOI22_X1 U20121 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16970) );
  AOI22_X1 U20122 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16969) );
  NAND4_X1 U20123 ( .A1(n16972), .A2(n16971), .A3(n16970), .A4(n16969), .ZN(
        n16978) );
  AOI22_X1 U20124 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16976) );
  AOI22_X1 U20125 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16975) );
  AOI22_X1 U20126 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16974) );
  AOI22_X1 U20127 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16973) );
  NAND4_X1 U20128 ( .A1(n16976), .A2(n16975), .A3(n16974), .A4(n16973), .ZN(
        n16977) );
  NOR2_X1 U20129 ( .A1(n16978), .A2(n16977), .ZN(n17257) );
  OAI21_X1 U20130 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n16980), .A(n16979), .ZN(
        n16981) );
  AOI22_X1 U20131 ( .A1(n17198), .A2(n17257), .B1(n16981), .B2(n17192), .ZN(
        P3_U2682) );
  AOI21_X1 U20132 ( .B1(n16982), .B2(n17007), .A(n17198), .ZN(n16994) );
  AOI22_X1 U20133 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17132), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16993) );
  AOI22_X1 U20134 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16992) );
  AOI22_X1 U20135 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17142), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16983) );
  OAI21_X1 U20136 ( .B1(n16984), .B2(n20795), .A(n16983), .ZN(n16990) );
  AOI22_X1 U20137 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16988) );
  AOI22_X1 U20138 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16987) );
  AOI22_X1 U20139 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16986) );
  AOI22_X1 U20140 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16985) );
  NAND4_X1 U20141 ( .A1(n16988), .A2(n16987), .A3(n16986), .A4(n16985), .ZN(
        n16989) );
  AOI211_X1 U20142 ( .C1(n17045), .C2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        n16990), .B(n16989), .ZN(n16991) );
  NAND3_X1 U20143 ( .A1(n16993), .A2(n16992), .A3(n16991), .ZN(n17260) );
  AOI22_X1 U20144 ( .A1(n16995), .A2(n16994), .B1(n17260), .B2(n17198), .ZN(
        n16996) );
  INV_X1 U20145 ( .A(n16996), .ZN(P3_U2683) );
  AOI22_X1 U20146 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17000) );
  AOI22_X1 U20147 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16999) );
  AOI22_X1 U20148 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16998) );
  AOI22_X1 U20149 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16997) );
  NAND4_X1 U20150 ( .A1(n17000), .A2(n16999), .A3(n16998), .A4(n16997), .ZN(
        n17006) );
  AOI22_X1 U20151 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17004) );
  AOI22_X1 U20152 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17003) );
  AOI22_X1 U20153 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17002) );
  AOI22_X1 U20154 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n15823), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17001) );
  NAND4_X1 U20155 ( .A1(n17004), .A2(n17003), .A3(n17002), .A4(n17001), .ZN(
        n17005) );
  NOR2_X1 U20156 ( .A1(n17006), .A2(n17005), .ZN(n17269) );
  OAI21_X1 U20157 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17019), .A(n17007), .ZN(
        n17008) );
  AOI22_X1 U20158 ( .A1(n17198), .A2(n17269), .B1(n17008), .B2(n17192), .ZN(
        P3_U2684) );
  NAND3_X1 U20159 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(n17077), .ZN(n17051) );
  NOR2_X1 U20160 ( .A1(n17050), .A2(n17051), .ZN(n17034) );
  NAND2_X1 U20161 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17034), .ZN(n17033) );
  AOI22_X1 U20162 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17018) );
  AOI22_X1 U20163 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17017) );
  AOI22_X1 U20164 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17009) );
  OAI21_X1 U20165 ( .B1(n9635), .B2(n17191), .A(n17009), .ZN(n17015) );
  AOI22_X1 U20166 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17013) );
  AOI22_X1 U20167 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17012) );
  AOI22_X1 U20168 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17011) );
  AOI22_X1 U20169 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17010) );
  NAND4_X1 U20170 ( .A1(n17013), .A2(n17012), .A3(n17011), .A4(n17010), .ZN(
        n17014) );
  AOI211_X1 U20171 ( .C1(n17132), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n17015), .B(n17014), .ZN(n17016) );
  NAND3_X1 U20172 ( .A1(n17018), .A2(n17017), .A3(n17016), .ZN(n17270) );
  OAI21_X1 U20173 ( .B1(n17020), .B2(n17019), .A(n17192), .ZN(n17021) );
  OAI21_X1 U20174 ( .B1(n17192), .B2(n17270), .A(n17021), .ZN(n17022) );
  OAI21_X1 U20175 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17033), .A(n17022), .ZN(
        P3_U2685) );
  AOI22_X1 U20176 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17026) );
  AOI22_X1 U20177 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17025) );
  AOI22_X1 U20178 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17024) );
  AOI22_X1 U20179 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17023) );
  NAND4_X1 U20180 ( .A1(n17026), .A2(n17025), .A3(n17024), .A4(n17023), .ZN(
        n17032) );
  AOI22_X1 U20181 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17030) );
  AOI22_X1 U20182 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17029) );
  AOI22_X1 U20183 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U20184 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17027) );
  NAND4_X1 U20185 ( .A1(n17030), .A2(n17029), .A3(n17028), .A4(n17027), .ZN(
        n17031) );
  NOR2_X1 U20186 ( .A1(n17032), .A2(n17031), .ZN(n17280) );
  OAI211_X1 U20187 ( .C1(n17034), .C2(P3_EBX_REG_17__SCAN_IN), .A(n17192), .B(
        n17033), .ZN(n17035) );
  OAI21_X1 U20188 ( .B1(n17280), .B2(n17192), .A(n17035), .ZN(P3_U2686) );
  NAND2_X1 U20189 ( .A1(n17192), .A2(n17036), .ZN(n17063) );
  AOI22_X1 U20190 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17048) );
  AOI22_X1 U20191 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17127), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17047) );
  AOI22_X1 U20192 ( .A1(n17037), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17038) );
  OAI21_X1 U20193 ( .B1(n9635), .B2(n17146), .A(n17038), .ZN(n17044) );
  AOI22_X1 U20194 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17042) );
  AOI22_X1 U20195 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17132), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17041) );
  AOI22_X1 U20196 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17040) );
  AOI22_X1 U20197 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17039) );
  NAND4_X1 U20198 ( .A1(n17042), .A2(n17041), .A3(n17040), .A4(n17039), .ZN(
        n17043) );
  AOI211_X1 U20199 ( .C1(n17045), .C2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A(
        n17044), .B(n17043), .ZN(n17046) );
  NAND3_X1 U20200 ( .A1(n17048), .A2(n17047), .A3(n17046), .ZN(n17281) );
  NAND2_X1 U20201 ( .A1(n17198), .A2(n17281), .ZN(n17049) );
  OAI221_X1 U20202 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17051), .C1(n17050), 
        .C2(n17063), .A(n17049), .ZN(P3_U2687) );
  NAND2_X1 U20203 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17077), .ZN(n17065) );
  AOI22_X1 U20204 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17061) );
  AOI22_X1 U20205 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17125), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17060) );
  AOI22_X1 U20206 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n17127), .ZN(n17052) );
  OAI21_X1 U20207 ( .B1(n20813), .B2(n12600), .A(n17052), .ZN(n17058) );
  AOI22_X1 U20208 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__7__SCAN_IN), .B2(n17149), .ZN(n17056) );
  AOI22_X1 U20209 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17055) );
  AOI22_X1 U20210 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17054) );
  AOI22_X1 U20211 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17108), .ZN(n17053) );
  NAND4_X1 U20212 ( .A1(n17056), .A2(n17055), .A3(n17054), .A4(n17053), .ZN(
        n17057) );
  AOI211_X1 U20213 ( .C1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .C2(n17152), .A(
        n17058), .B(n17057), .ZN(n17059) );
  NAND3_X1 U20214 ( .A1(n17061), .A2(n17060), .A3(n17059), .ZN(n17289) );
  NAND2_X1 U20215 ( .A1(n17198), .A2(n17289), .ZN(n17062) );
  OAI221_X1 U20216 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17065), .C1(n17064), 
        .C2(n17063), .A(n17062), .ZN(P3_U2688) );
  NAND2_X1 U20217 ( .A1(n17192), .A2(P3_EBX_REG_14__SCAN_IN), .ZN(n17079) );
  AOI22_X1 U20218 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17142), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17075) );
  AOI22_X1 U20219 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17074) );
  AOI22_X1 U20220 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17066) );
  OAI21_X1 U20221 ( .B1(n12600), .B2(n17174), .A(n17066), .ZN(n17072) );
  AOI22_X1 U20222 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17070) );
  AOI22_X1 U20223 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17069) );
  AOI22_X1 U20224 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17127), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17068) );
  AOI22_X1 U20225 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17067) );
  NAND4_X1 U20226 ( .A1(n17070), .A2(n17069), .A3(n17068), .A4(n17067), .ZN(
        n17071) );
  AOI211_X1 U20227 ( .C1(n17159), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n17072), .B(n17071), .ZN(n17073) );
  NAND3_X1 U20228 ( .A1(n17075), .A2(n17074), .A3(n17073), .ZN(n17293) );
  AOI22_X1 U20229 ( .A1(n17198), .A2(n17293), .B1(n17077), .B2(n17076), .ZN(
        n17078) );
  OAI21_X1 U20230 ( .B1(n17080), .B2(n17079), .A(n17078), .ZN(P3_U2689) );
  AOI22_X1 U20231 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17084) );
  AOI22_X1 U20232 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17083) );
  AOI22_X1 U20233 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17082) );
  AOI22_X1 U20234 ( .A1(n17127), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17081) );
  NAND4_X1 U20235 ( .A1(n17084), .A2(n17083), .A3(n17082), .A4(n17081), .ZN(
        n17090) );
  AOI22_X1 U20236 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17142), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17088) );
  AOI22_X1 U20237 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17087) );
  AOI22_X1 U20238 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17086) );
  AOI22_X1 U20239 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17085) );
  NAND4_X1 U20240 ( .A1(n17088), .A2(n17087), .A3(n17086), .A4(n17085), .ZN(
        n17089) );
  NOR2_X1 U20241 ( .A1(n17090), .A2(n17089), .ZN(n17302) );
  NOR2_X1 U20242 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17093), .ZN(n17092) );
  OAI22_X1 U20243 ( .A1(n17302), .A2(n17192), .B1(n17092), .B2(n17091), .ZN(
        P3_U2691) );
  AOI21_X1 U20244 ( .B1(n17094), .B2(n17120), .A(n17198), .ZN(n17105) );
  AOI22_X1 U20245 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17142), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17104) );
  AOI22_X1 U20246 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17127), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17103) );
  INV_X1 U20247 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17185) );
  AOI22_X1 U20248 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17095) );
  OAI21_X1 U20249 ( .B1(n12600), .B2(n17185), .A(n17095), .ZN(n17101) );
  AOI22_X1 U20250 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17099) );
  AOI22_X1 U20251 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17098) );
  AOI22_X1 U20252 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17097) );
  AOI22_X1 U20253 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17096) );
  NAND4_X1 U20254 ( .A1(n17099), .A2(n17098), .A3(n17097), .A4(n17096), .ZN(
        n17100) );
  AOI211_X1 U20255 ( .C1(n17150), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n17101), .B(n17100), .ZN(n17102) );
  NAND3_X1 U20256 ( .A1(n17104), .A2(n17103), .A3(n17102), .ZN(n17305) );
  AOI22_X1 U20257 ( .A1(n9783), .A2(n17105), .B1(n17305), .B2(n17198), .ZN(
        n17106) );
  INV_X1 U20258 ( .A(n17106), .ZN(P3_U2692) );
  AOI22_X1 U20259 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17119) );
  AOI22_X1 U20260 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17118) );
  AOI22_X1 U20261 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17107) );
  OAI21_X1 U20262 ( .B1(n12600), .B2(n17191), .A(n17107), .ZN(n17115) );
  AOI22_X1 U20263 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17113) );
  AOI22_X1 U20264 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17142), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17112) );
  AOI22_X1 U20265 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17127), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17111) );
  AOI22_X1 U20266 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17108), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17110) );
  NAND4_X1 U20267 ( .A1(n17113), .A2(n17112), .A3(n17111), .A4(n17110), .ZN(
        n17114) );
  AOI211_X1 U20268 ( .C1(n17116), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n17115), .B(n17114), .ZN(n17117) );
  NAND3_X1 U20269 ( .A1(n17119), .A2(n17118), .A3(n17117), .ZN(n17308) );
  INV_X1 U20270 ( .A(n17308), .ZN(n17122) );
  OAI21_X1 U20271 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17141), .A(n17120), .ZN(
        n17121) );
  AOI22_X1 U20272 ( .A1(n17198), .A2(n17122), .B1(n17121), .B2(n17192), .ZN(
        P3_U2693) );
  AOI21_X1 U20273 ( .B1(n17123), .B2(n17163), .A(n17198), .ZN(n17124) );
  INV_X1 U20274 ( .A(n17124), .ZN(n17140) );
  AOI22_X1 U20275 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20276 ( .A1(n9588), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17130) );
  AOI22_X1 U20277 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17142), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17129) );
  AOI22_X1 U20278 ( .A1(n17127), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14458), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17128) );
  NAND4_X1 U20279 ( .A1(n17131), .A2(n17130), .A3(n17129), .A4(n17128), .ZN(
        n17139) );
  AOI22_X1 U20280 ( .A1(n17045), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17137) );
  AOI22_X1 U20281 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17136) );
  AOI22_X1 U20282 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17132), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17135) );
  AOI22_X1 U20283 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17134) );
  NAND4_X1 U20284 ( .A1(n17137), .A2(n17136), .A3(n17135), .A4(n17134), .ZN(
        n17138) );
  NOR2_X1 U20285 ( .A1(n17139), .A2(n17138), .ZN(n17313) );
  OAI22_X1 U20286 ( .A1(n17141), .A2(n17140), .B1(n17313), .B2(n17192), .ZN(
        P3_U2694) );
  AOI22_X1 U20287 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17037), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17162) );
  AOI22_X1 U20288 ( .A1(n17133), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17161) );
  AOI22_X1 U20289 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17145) );
  OAI21_X1 U20290 ( .B1(n12600), .B2(n17146), .A(n17145), .ZN(n17158) );
  AOI22_X1 U20291 ( .A1(n17148), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17147), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17156) );
  AOI22_X1 U20292 ( .A1(n17150), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17155) );
  AOI22_X1 U20293 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17154) );
  AOI22_X1 U20294 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9588), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17153) );
  NAND4_X1 U20295 ( .A1(n17156), .A2(n17155), .A3(n17154), .A4(n17153), .ZN(
        n17157) );
  AOI211_X1 U20296 ( .C1(n17159), .C2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n17158), .B(n17157), .ZN(n17160) );
  NAND3_X1 U20297 ( .A1(n17162), .A2(n17161), .A3(n17160), .ZN(n17316) );
  INV_X1 U20298 ( .A(n17316), .ZN(n17165) );
  OAI21_X1 U20299 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17170), .A(n17163), .ZN(
        n17164) );
  AOI22_X1 U20300 ( .A1(n17198), .A2(n17165), .B1(n17164), .B2(n17192), .ZN(
        P3_U2695) );
  AOI21_X1 U20301 ( .B1(n17167), .B2(n17166), .A(n17198), .ZN(n17168) );
  INV_X1 U20302 ( .A(n17168), .ZN(n17169) );
  OAI22_X1 U20303 ( .A1(n17170), .A2(n17169), .B1(n20813), .B2(n17192), .ZN(
        P3_U2696) );
  NOR2_X1 U20304 ( .A1(n18225), .A2(n17171), .ZN(n17197) );
  INV_X1 U20305 ( .A(n17197), .ZN(n17196) );
  NOR2_X1 U20306 ( .A1(n17172), .A2(n17196), .ZN(n17182) );
  NAND2_X1 U20307 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17182), .ZN(n17175) );
  NAND3_X1 U20308 ( .A1(n17175), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n17192), .ZN(
        n17173) );
  OAI221_X1 U20309 ( .B1(n17175), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n17192), 
        .C2(n17174), .A(n17173), .ZN(P3_U2697) );
  OAI211_X1 U20310 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n17176), .A(n17175), .B(
        n17192), .ZN(n17177) );
  OAI21_X1 U20311 ( .B1(n17192), .B2(n17178), .A(n17177), .ZN(P3_U2698) );
  NAND2_X1 U20312 ( .A1(n17179), .A2(n17197), .ZN(n17188) );
  NOR2_X1 U20313 ( .A1(n17183), .A2(n17188), .ZN(n17187) );
  AOI21_X1 U20314 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17192), .A(n17187), .ZN(
        n17181) );
  INV_X1 U20315 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17180) );
  OAI22_X1 U20316 ( .A1(n17182), .A2(n17181), .B1(n17180), .B2(n17192), .ZN(
        P3_U2699) );
  OAI21_X1 U20317 ( .B1(n17183), .B2(n17198), .A(n17188), .ZN(n17184) );
  INV_X1 U20318 ( .A(n17184), .ZN(n17186) );
  OAI22_X1 U20319 ( .A1(n17187), .A2(n17186), .B1(n17185), .B2(n17192), .ZN(
        P3_U2700) );
  OAI221_X1 U20320 ( .B1(P3_EBX_REG_2__SCAN_IN), .B2(n17201), .C1(
        P3_EBX_REG_2__SCAN_IN), .C2(n17189), .A(n17188), .ZN(n17190) );
  AOI22_X1 U20321 ( .A1(n17198), .A2(n17191), .B1(n17190), .B2(n17192), .ZN(
        P3_U2701) );
  INV_X1 U20322 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17193) );
  OAI222_X1 U20323 ( .A1(n17196), .A2(n17195), .B1(n17194), .B2(n17201), .C1(
        n17193), .C2(n17192), .ZN(P3_U2702) );
  AOI22_X1 U20324 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17198), .B1(
        n17197), .B2(n17200), .ZN(n17199) );
  OAI21_X1 U20325 ( .B1(n17201), .B2(n17200), .A(n17199), .ZN(P3_U2703) );
  INV_X1 U20326 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17359) );
  INV_X1 U20327 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17362) );
  INV_X1 U20328 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17384) );
  INV_X1 U20329 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17440) );
  NAND2_X1 U20330 ( .A1(n17202), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n17346) );
  INV_X1 U20331 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17403) );
  INV_X1 U20332 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17405) );
  INV_X1 U20333 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17407) );
  INV_X1 U20334 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17409) );
  NOR4_X1 U20335 ( .A1(n17403), .A2(n17405), .A3(n17407), .A4(n17409), .ZN(
        n17203) );
  NAND4_X1 U20336 ( .A1(n17344), .A2(P3_EAX_REG_7__SCAN_IN), .A3(
        P3_EAX_REG_6__SCAN_IN), .A4(n17203), .ZN(n17318) );
  NAND4_X1 U20337 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n17204)
         );
  NOR2_X1 U20338 ( .A1(n17318), .A2(n17204), .ZN(n17205) );
  NAND4_X1 U20339 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_8__SCAN_IN), .A4(n17205), .ZN(n17294) );
  NOR2_X2 U20340 ( .A1(n17384), .A2(n17294), .ZN(n17287) );
  NAND2_X1 U20341 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .ZN(n17248) );
  NAND4_X1 U20342 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_21__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17206)
         );
  NAND2_X1 U20343 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17244), .ZN(n17243) );
  NAND2_X1 U20344 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17239), .ZN(n17238) );
  NAND2_X1 U20345 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17228), .ZN(n17224) );
  NOR2_X2 U20346 ( .A1(n17359), .A2(n17224), .ZN(n17220) );
  NAND2_X1 U20347 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17220), .ZN(n17216) );
  NAND2_X1 U20348 ( .A1(n17211), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17210) );
  NAND2_X1 U20349 ( .A1(n18219), .A2(n17339), .ZN(n17256) );
  OAI22_X1 U20350 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17292), .B1(n17339), 
        .B2(n17211), .ZN(n17207) );
  AOI22_X1 U20351 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17282), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17207), .ZN(n17208) );
  OAI21_X1 U20352 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17210), .A(n17208), .ZN(
        P3_U2704) );
  NAND2_X1 U20353 ( .A1(n17209), .A2(n17339), .ZN(n17286) );
  AOI22_X1 U20354 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17274), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17282), .ZN(n17213) );
  OAI211_X1 U20355 ( .C1(n17211), .C2(P3_EAX_REG_30__SCAN_IN), .A(n20931), .B(
        n17210), .ZN(n17212) );
  OAI211_X1 U20356 ( .C1(n17214), .C2(n17350), .A(n17213), .B(n17212), .ZN(
        P3_U2705) );
  INV_X1 U20357 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18214) );
  AOI22_X1 U20358 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17274), .B1(n17215), .B2(
        n17317), .ZN(n17218) );
  OAI211_X1 U20359 ( .C1(n17220), .C2(P3_EAX_REG_29__SCAN_IN), .A(n20931), .B(
        n17216), .ZN(n17217) );
  OAI211_X1 U20360 ( .C1(n17256), .C2(n18214), .A(n17218), .B(n17217), .ZN(
        P3_U2706) );
  INV_X1 U20361 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18209) );
  AOI22_X1 U20362 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17274), .B1(n17219), .B2(
        n17317), .ZN(n17223) );
  AOI211_X1 U20363 ( .C1(n17359), .C2(n17224), .A(n17220), .B(n17339), .ZN(
        n17221) );
  INV_X1 U20364 ( .A(n17221), .ZN(n17222) );
  OAI211_X1 U20365 ( .C1(n17256), .C2(n18209), .A(n17223), .B(n17222), .ZN(
        P3_U2707) );
  AOI22_X1 U20366 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17274), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17282), .ZN(n17226) );
  OAI211_X1 U20367 ( .C1(n17228), .C2(P3_EAX_REG_27__SCAN_IN), .A(n20931), .B(
        n17224), .ZN(n17225) );
  OAI211_X1 U20368 ( .C1(n17350), .C2(n17227), .A(n17226), .B(n17225), .ZN(
        P3_U2708) );
  AOI22_X1 U20369 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17274), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17282), .ZN(n17231) );
  AOI211_X1 U20370 ( .C1(n17362), .C2(n17233), .A(n17228), .B(n17339), .ZN(
        n17229) );
  INV_X1 U20371 ( .A(n17229), .ZN(n17230) );
  OAI211_X1 U20372 ( .C1(n17232), .C2(n17350), .A(n17231), .B(n17230), .ZN(
        P3_U2709) );
  AOI22_X1 U20373 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17274), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17282), .ZN(n17236) );
  OAI211_X1 U20374 ( .C1(n17234), .C2(P3_EAX_REG_25__SCAN_IN), .A(n20931), .B(
        n17233), .ZN(n17235) );
  OAI211_X1 U20375 ( .C1(n17237), .C2(n17350), .A(n17236), .B(n17235), .ZN(
        P3_U2710) );
  AOI22_X1 U20376 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17274), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17282), .ZN(n17241) );
  OAI211_X1 U20377 ( .C1(n17239), .C2(P3_EAX_REG_24__SCAN_IN), .A(n20931), .B(
        n17238), .ZN(n17240) );
  OAI211_X1 U20378 ( .C1(n17242), .C2(n17350), .A(n17241), .B(n17240), .ZN(
        P3_U2711) );
  AOI22_X1 U20379 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17274), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17282), .ZN(n17246) );
  OAI211_X1 U20380 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17244), .A(n20931), .B(
        n17243), .ZN(n17245) );
  OAI211_X1 U20381 ( .C1(n17247), .C2(n17350), .A(n17246), .B(n17245), .ZN(
        P3_U2712) );
  INV_X1 U20382 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17421) );
  NAND2_X1 U20383 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17275), .ZN(n17271) );
  NOR2_X1 U20384 ( .A1(n17248), .A2(n17271), .ZN(n17251) );
  NAND2_X1 U20385 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17251), .ZN(n17255) );
  OAI22_X1 U20386 ( .A1(n20902), .A2(n17256), .B1(n17350), .B2(n17249), .ZN(
        n17250) );
  INV_X1 U20387 ( .A(n17250), .ZN(n17254) );
  INV_X1 U20388 ( .A(n17251), .ZN(n17261) );
  NAND2_X1 U20389 ( .A1(n20931), .A2(n17261), .ZN(n17264) );
  OAI21_X1 U20390 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17292), .A(n17264), .ZN(
        n17252) );
  AOI22_X1 U20391 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17274), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17252), .ZN(n17253) );
  OAI211_X1 U20392 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17255), .A(n17254), .B(
        n17253), .ZN(P3_U2713) );
  INV_X1 U20393 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17372) );
  OAI22_X1 U20394 ( .A1(n17257), .A2(n17350), .B1(n18212), .B2(n17256), .ZN(
        n17258) );
  AOI21_X1 U20395 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17274), .A(n17258), .ZN(
        n17259) );
  OAI221_X1 U20396 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17261), .C1(n17372), 
        .C2(n17264), .A(n17259), .ZN(P3_U2714) );
  INV_X1 U20397 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17374) );
  AOI22_X1 U20398 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17274), .B1(n17317), .B2(
        n17260), .ZN(n17263) );
  INV_X1 U20399 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17376) );
  NOR2_X1 U20400 ( .A1(n17376), .A2(n17271), .ZN(n17265) );
  AOI22_X1 U20401 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17282), .B1(n17265), .B2(
        n17261), .ZN(n17262) );
  OAI211_X1 U20402 ( .C1(n17374), .C2(n17264), .A(n17263), .B(n17262), .ZN(
        P3_U2715) );
  AOI22_X1 U20403 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17274), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17282), .ZN(n17268) );
  AOI211_X1 U20404 ( .C1(n17376), .C2(n17271), .A(n17265), .B(n17339), .ZN(
        n17266) );
  INV_X1 U20405 ( .A(n17266), .ZN(n17267) );
  OAI211_X1 U20406 ( .C1(n17269), .C2(n17350), .A(n17268), .B(n17267), .ZN(
        P3_U2716) );
  INV_X1 U20407 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18199) );
  AOI22_X1 U20408 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n17282), .B1(n17317), .B2(
        n17270), .ZN(n17273) );
  OAI211_X1 U20409 ( .C1(n17275), .C2(P3_EAX_REG_18__SCAN_IN), .A(n20931), .B(
        n17271), .ZN(n17272) );
  OAI211_X1 U20410 ( .C1(n17286), .C2(n18199), .A(n17273), .B(n17272), .ZN(
        P3_U2717) );
  AOI22_X1 U20411 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17274), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17282), .ZN(n17279) );
  INV_X1 U20412 ( .A(n17283), .ZN(n17277) );
  INV_X1 U20413 ( .A(n17275), .ZN(n17276) );
  OAI211_X1 U20414 ( .C1(n17277), .C2(P3_EAX_REG_17__SCAN_IN), .A(n20931), .B(
        n17276), .ZN(n17278) );
  OAI211_X1 U20415 ( .C1(n17280), .C2(n17350), .A(n17279), .B(n17278), .ZN(
        P3_U2718) );
  AOI22_X1 U20416 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n17282), .B1(n17317), .B2(
        n17281), .ZN(n17285) );
  OAI211_X1 U20417 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17287), .A(n20931), .B(
        n17283), .ZN(n17284) );
  OAI211_X1 U20418 ( .C1(n17286), .C2(n18186), .A(n17285), .B(n17284), .ZN(
        P3_U2719) );
  AOI211_X1 U20419 ( .C1(n17384), .C2(n17294), .A(n17339), .B(n17287), .ZN(
        n17288) );
  AOI21_X1 U20420 ( .B1(n17317), .B2(n17289), .A(n17288), .ZN(n17290) );
  OAI21_X1 U20421 ( .B1(n17291), .B2(n17343), .A(n17290), .ZN(P3_U2720) );
  INV_X1 U20422 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17454) );
  INV_X1 U20423 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17399) );
  INV_X1 U20424 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17401) );
  NAND2_X1 U20425 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17338), .ZN(n17334) );
  NAND2_X1 U20426 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17312), .ZN(n17310) );
  INV_X1 U20427 ( .A(n17310), .ZN(n17315) );
  NAND2_X1 U20428 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17315), .ZN(n17307) );
  NOR2_X1 U20429 ( .A1(n17454), .A2(n17307), .ZN(n17301) );
  NAND2_X1 U20430 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17304), .ZN(n17297) );
  AOI22_X1 U20431 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17348), .B1(n17317), .B2(
        n17293), .ZN(n17296) );
  NAND3_X1 U20432 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n20931), .A3(n17294), 
        .ZN(n17295) );
  OAI211_X1 U20433 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17297), .A(n17296), .B(
        n17295), .ZN(P3_U2721) );
  INV_X1 U20434 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17459) );
  INV_X1 U20435 ( .A(n17297), .ZN(n17300) );
  AOI21_X1 U20436 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n20931), .A(n17304), .ZN(
        n17299) );
  OAI222_X1 U20437 ( .A1(n17343), .A2(n17459), .B1(n17300), .B2(n17299), .C1(
        n17350), .C2(n17298), .ZN(P3_U2722) );
  INV_X1 U20438 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17456) );
  AOI21_X1 U20439 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n20931), .A(n17301), .ZN(
        n17303) );
  OAI222_X1 U20440 ( .A1(n17343), .A2(n17456), .B1(n17304), .B2(n17303), .C1(
        n17350), .C2(n17302), .ZN(P3_U2723) );
  NAND2_X1 U20441 ( .A1(n20931), .A2(n17307), .ZN(n17311) );
  AOI22_X1 U20442 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17348), .B1(n17317), .B2(
        n17305), .ZN(n17306) );
  OAI221_X1 U20443 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17307), .C1(n17454), 
        .C2(n17311), .A(n17306), .ZN(P3_U2724) );
  INV_X1 U20444 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17392) );
  AOI22_X1 U20445 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17348), .B1(n17317), .B2(
        n17308), .ZN(n17309) );
  OAI221_X1 U20446 ( .B1(n17311), .B2(n17392), .C1(n17311), .C2(n17310), .A(
        n17309), .ZN(P3_U2725) );
  AOI21_X1 U20447 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n20931), .A(n17312), .ZN(
        n17314) );
  OAI222_X1 U20448 ( .A1(n17343), .A2(n17450), .B1(n17315), .B2(n17314), .C1(
        n17350), .C2(n17313), .ZN(P3_U2726) );
  INV_X1 U20449 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17448) );
  INV_X1 U20450 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17396) );
  AOI22_X1 U20451 ( .A1(n17317), .A2(n17316), .B1(n17323), .B2(n17396), .ZN(
        n17320) );
  NAND3_X1 U20452 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n20931), .A3(n17318), .ZN(
        n17319) );
  OAI211_X1 U20453 ( .C1(n17343), .C2(n17448), .A(n17320), .B(n17319), .ZN(
        P3_U2727) );
  INV_X1 U20454 ( .A(n17324), .ZN(n17330) );
  AOI22_X1 U20455 ( .A1(n17330), .A2(P3_EAX_REG_6__SCAN_IN), .B1(
        P3_EAX_REG_7__SCAN_IN), .B2(n20931), .ZN(n17322) );
  OAI222_X1 U20456 ( .A1(n17343), .A2(n18222), .B1(n17323), .B2(n17322), .C1(
        n17350), .C2(n17321), .ZN(P3_U2728) );
  AOI21_X1 U20457 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n20931), .A(n17330), .ZN(
        n17327) );
  NOR2_X1 U20458 ( .A1(n17401), .A2(n17324), .ZN(n17326) );
  OAI222_X1 U20459 ( .A1(n17343), .A2(n18218), .B1(n17327), .B2(n17326), .C1(
        n17350), .C2(n17325), .ZN(P3_U2729) );
  AOI21_X1 U20460 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n20931), .A(n17333), .ZN(
        n17329) );
  OAI222_X1 U20461 ( .A1(n17343), .A2(n18213), .B1(n17330), .B2(n17329), .C1(
        n17350), .C2(n17328), .ZN(P3_U2730) );
  INV_X1 U20462 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18208) );
  AOI21_X1 U20463 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n20931), .A(n17337), .ZN(
        n17332) );
  OAI222_X1 U20464 ( .A1(n18208), .A2(n17343), .B1(n17333), .B2(n17332), .C1(
        n17350), .C2(n17331), .ZN(P3_U2731) );
  INV_X1 U20465 ( .A(n17334), .ZN(n17342) );
  AOI21_X1 U20466 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n20931), .A(n17342), .ZN(
        n17336) );
  OAI222_X1 U20467 ( .A1(n20912), .A2(n17343), .B1(n17337), .B2(n17336), .C1(
        n17350), .C2(n17335), .ZN(P3_U2732) );
  AOI21_X1 U20468 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n20931), .A(n17338), .ZN(
        n17341) );
  OAI222_X1 U20469 ( .A1(n18199), .A2(n17343), .B1(n17342), .B2(n17341), .C1(
        n17350), .C2(n17340), .ZN(P3_U2733) );
  AOI211_X1 U20470 ( .C1(n17440), .C2(n17346), .A(n17339), .B(n17344), .ZN(
        n17347) );
  AOI21_X1 U20471 ( .B1(n17348), .B2(BUF2_REG_1__SCAN_IN), .A(n17347), .ZN(
        n17349) );
  OAI21_X1 U20472 ( .B1(n17351), .B2(n17350), .A(n17349), .ZN(P3_U2734) );
  INV_X1 U20473 ( .A(n17844), .ZN(n17630) );
  NAND2_X1 U20474 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17630), .ZN(n18835) );
  NOR2_X1 U20475 ( .A1(n17354), .A2(n20915), .ZN(P3_U2736) );
  INV_X1 U20476 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17437) );
  INV_X2 U20477 ( .A(n18835), .ZN(n17411) );
  AOI22_X1 U20478 ( .A1(n17411), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17355) );
  OAI21_X1 U20479 ( .B1(n17437), .B2(n17381), .A(n17355), .ZN(P3_U2737) );
  INV_X1 U20480 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17357) );
  AOI22_X1 U20481 ( .A1(n17411), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17356) );
  OAI21_X1 U20482 ( .B1(n17357), .B2(n17381), .A(n17356), .ZN(P3_U2738) );
  AOI22_X1 U20483 ( .A1(n17411), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17358) );
  OAI21_X1 U20484 ( .B1(n17359), .B2(n17381), .A(n17358), .ZN(P3_U2739) );
  INV_X1 U20485 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17433) );
  AOI22_X1 U20486 ( .A1(n17411), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17360) );
  OAI21_X1 U20487 ( .B1(n17433), .B2(n17381), .A(n17360), .ZN(P3_U2740) );
  AOI22_X1 U20488 ( .A1(n17411), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17361) );
  OAI21_X1 U20489 ( .B1(n17362), .B2(n17381), .A(n17361), .ZN(P3_U2741) );
  INV_X1 U20490 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17364) );
  AOI22_X1 U20491 ( .A1(n17411), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17363) );
  OAI21_X1 U20492 ( .B1(n17364), .B2(n17381), .A(n17363), .ZN(P3_U2742) );
  INV_X1 U20493 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17366) );
  AOI22_X1 U20494 ( .A1(n17411), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17365) );
  OAI21_X1 U20495 ( .B1(n17366), .B2(n17381), .A(n17365), .ZN(P3_U2743) );
  INV_X1 U20496 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17368) );
  AOI22_X1 U20497 ( .A1(n17411), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17367) );
  OAI21_X1 U20498 ( .B1(n17368), .B2(n17381), .A(n17367), .ZN(P3_U2744) );
  INV_X1 U20499 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17370) );
  AOI22_X1 U20500 ( .A1(n17411), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17369) );
  OAI21_X1 U20501 ( .B1(n17370), .B2(n17381), .A(n17369), .ZN(P3_U2745) );
  AOI22_X1 U20502 ( .A1(n17411), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17371) );
  OAI21_X1 U20503 ( .B1(n17372), .B2(n17381), .A(n17371), .ZN(P3_U2746) );
  AOI22_X1 U20504 ( .A1(n17411), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17373) );
  OAI21_X1 U20505 ( .B1(n17374), .B2(n17381), .A(n17373), .ZN(P3_U2747) );
  AOI22_X1 U20506 ( .A1(n17411), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17375) );
  OAI21_X1 U20507 ( .B1(n17376), .B2(n17381), .A(n17375), .ZN(P3_U2748) );
  INV_X1 U20508 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17378) );
  AOI22_X1 U20509 ( .A1(n17411), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17377) );
  OAI21_X1 U20510 ( .B1(n17378), .B2(n17381), .A(n17377), .ZN(P3_U2749) );
  AOI22_X1 U20511 ( .A1(n17411), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17379) );
  OAI21_X1 U20512 ( .B1(n17421), .B2(n17381), .A(n17379), .ZN(P3_U2750) );
  INV_X1 U20513 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17382) );
  AOI22_X1 U20514 ( .A1(n17411), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17380) );
  OAI21_X1 U20515 ( .B1(n17382), .B2(n17381), .A(n17380), .ZN(P3_U2751) );
  AOI22_X1 U20516 ( .A1(n17411), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17383) );
  OAI21_X1 U20517 ( .B1(n17384), .B2(n17413), .A(n17383), .ZN(P3_U2752) );
  INV_X1 U20518 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17463) );
  AOI22_X1 U20519 ( .A1(n17411), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17385) );
  OAI21_X1 U20520 ( .B1(n17463), .B2(n17413), .A(n17385), .ZN(P3_U2753) );
  INV_X1 U20521 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17387) );
  AOI22_X1 U20522 ( .A1(n17411), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17386) );
  OAI21_X1 U20523 ( .B1(n17387), .B2(n17413), .A(n17386), .ZN(P3_U2754) );
  INV_X1 U20524 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17389) );
  AOI22_X1 U20525 ( .A1(n17411), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17388) );
  OAI21_X1 U20526 ( .B1(n17389), .B2(n17413), .A(n17388), .ZN(P3_U2755) );
  AOI22_X1 U20527 ( .A1(n17411), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17390) );
  OAI21_X1 U20528 ( .B1(n17454), .B2(n17413), .A(n17390), .ZN(P3_U2756) );
  AOI22_X1 U20529 ( .A1(n17411), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17391) );
  OAI21_X1 U20530 ( .B1(n17392), .B2(n17413), .A(n17391), .ZN(P3_U2757) );
  INV_X1 U20531 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17394) );
  AOI22_X1 U20532 ( .A1(n17411), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17393) );
  OAI21_X1 U20533 ( .B1(n17394), .B2(n17413), .A(n17393), .ZN(P3_U2758) );
  AOI22_X1 U20534 ( .A1(n17411), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17395) );
  OAI21_X1 U20535 ( .B1(n17396), .B2(n17413), .A(n17395), .ZN(P3_U2759) );
  AOI22_X1 U20536 ( .A1(n17411), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17398) );
  OAI21_X1 U20537 ( .B1(n17399), .B2(n17413), .A(n17398), .ZN(P3_U2760) );
  AOI22_X1 U20538 ( .A1(n17411), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17400) );
  OAI21_X1 U20539 ( .B1(n17401), .B2(n17413), .A(n17400), .ZN(P3_U2761) );
  AOI22_X1 U20540 ( .A1(n17411), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17402) );
  OAI21_X1 U20541 ( .B1(n17403), .B2(n17413), .A(n17402), .ZN(P3_U2762) );
  AOI22_X1 U20542 ( .A1(n17411), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17404) );
  OAI21_X1 U20543 ( .B1(n17405), .B2(n17413), .A(n17404), .ZN(P3_U2763) );
  AOI22_X1 U20544 ( .A1(n17411), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17406) );
  OAI21_X1 U20545 ( .B1(n17407), .B2(n17413), .A(n17406), .ZN(P3_U2764) );
  AOI22_X1 U20546 ( .A1(n17411), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17408) );
  OAI21_X1 U20547 ( .B1(n17409), .B2(n17413), .A(n17408), .ZN(P3_U2765) );
  AOI22_X1 U20548 ( .A1(n17411), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17410) );
  OAI21_X1 U20549 ( .B1(n17440), .B2(n17413), .A(n17410), .ZN(P3_U2766) );
  AOI22_X1 U20550 ( .A1(n17411), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17397), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17412) );
  OAI21_X1 U20551 ( .B1(n17414), .B2(n17413), .A(n17412), .ZN(P3_U2767) );
  NOR3_X1 U20552 ( .A1(n18193), .A2(n17418), .A3(n17417), .ZN(n17430) );
  AOI22_X1 U20553 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17464), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17465), .ZN(n17419) );
  OAI21_X1 U20554 ( .B1(n18186), .B2(n17458), .A(n17419), .ZN(P3_U2768) );
  AOI22_X1 U20555 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17466), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17465), .ZN(n17420) );
  OAI21_X1 U20556 ( .B1(n17421), .B2(n17462), .A(n17420), .ZN(P3_U2769) );
  AOI22_X1 U20557 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17464), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17465), .ZN(n17422) );
  OAI21_X1 U20558 ( .B1(n18199), .B2(n17458), .A(n17422), .ZN(P3_U2770) );
  AOI22_X1 U20559 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17464), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17465), .ZN(n17423) );
  OAI21_X1 U20560 ( .B1(n20912), .B2(n17458), .A(n17423), .ZN(P3_U2771) );
  AOI22_X1 U20561 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17464), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17465), .ZN(n17424) );
  OAI21_X1 U20562 ( .B1(n18208), .B2(n17458), .A(n17424), .ZN(P3_U2772) );
  AOI22_X1 U20563 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17464), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17465), .ZN(n17425) );
  OAI21_X1 U20564 ( .B1(n18213), .B2(n17458), .A(n17425), .ZN(P3_U2773) );
  AOI22_X1 U20565 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17430), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17465), .ZN(n17426) );
  OAI21_X1 U20566 ( .B1(n18218), .B2(n17458), .A(n17426), .ZN(P3_U2774) );
  AOI22_X1 U20567 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17430), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17465), .ZN(n17427) );
  OAI21_X1 U20568 ( .B1(n18222), .B2(n17458), .A(n17427), .ZN(P3_U2775) );
  AOI22_X1 U20569 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17430), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17465), .ZN(n17428) );
  OAI21_X1 U20570 ( .B1(n17448), .B2(n17458), .A(n17428), .ZN(P3_U2776) );
  AOI22_X1 U20571 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17430), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17465), .ZN(n17429) );
  OAI21_X1 U20572 ( .B1(n17450), .B2(n17458), .A(n17429), .ZN(P3_U2777) );
  INV_X1 U20573 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17452) );
  AOI22_X1 U20574 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17430), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17465), .ZN(n17431) );
  OAI21_X1 U20575 ( .B1(n17452), .B2(n17458), .A(n17431), .ZN(P3_U2778) );
  AOI22_X1 U20576 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17466), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17465), .ZN(n17432) );
  OAI21_X1 U20577 ( .B1(n17433), .B2(n17462), .A(n17432), .ZN(P3_U2779) );
  AOI22_X1 U20578 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17464), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17465), .ZN(n17434) );
  OAI21_X1 U20579 ( .B1(n17456), .B2(n17458), .A(n17434), .ZN(P3_U2780) );
  AOI22_X1 U20580 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17464), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17465), .ZN(n17435) );
  OAI21_X1 U20581 ( .B1(n17459), .B2(n17458), .A(n17435), .ZN(P3_U2781) );
  AOI22_X1 U20582 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17466), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17465), .ZN(n17436) );
  OAI21_X1 U20583 ( .B1(n17437), .B2(n17462), .A(n17436), .ZN(P3_U2782) );
  AOI22_X1 U20584 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17464), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17465), .ZN(n17438) );
  OAI21_X1 U20585 ( .B1(n18186), .B2(n17458), .A(n17438), .ZN(P3_U2783) );
  AOI22_X1 U20586 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17466), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17465), .ZN(n17439) );
  OAI21_X1 U20587 ( .B1(n17440), .B2(n17462), .A(n17439), .ZN(P3_U2784) );
  AOI22_X1 U20588 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17464), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17465), .ZN(n17441) );
  OAI21_X1 U20589 ( .B1(n18199), .B2(n17458), .A(n17441), .ZN(P3_U2785) );
  AOI22_X1 U20590 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17464), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17460), .ZN(n17442) );
  OAI21_X1 U20591 ( .B1(n20912), .B2(n17458), .A(n17442), .ZN(P3_U2786) );
  AOI22_X1 U20592 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17464), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17460), .ZN(n17443) );
  OAI21_X1 U20593 ( .B1(n18208), .B2(n17458), .A(n17443), .ZN(P3_U2787) );
  AOI22_X1 U20594 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17464), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17460), .ZN(n17444) );
  OAI21_X1 U20595 ( .B1(n18213), .B2(n17458), .A(n17444), .ZN(P3_U2788) );
  AOI22_X1 U20596 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17464), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17460), .ZN(n17445) );
  OAI21_X1 U20597 ( .B1(n18218), .B2(n17458), .A(n17445), .ZN(P3_U2789) );
  AOI22_X1 U20598 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17464), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17460), .ZN(n17446) );
  OAI21_X1 U20599 ( .B1(n18222), .B2(n17458), .A(n17446), .ZN(P3_U2790) );
  AOI22_X1 U20600 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17464), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17460), .ZN(n17447) );
  OAI21_X1 U20601 ( .B1(n17448), .B2(n17458), .A(n17447), .ZN(P3_U2791) );
  AOI22_X1 U20602 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17464), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17460), .ZN(n17449) );
  OAI21_X1 U20603 ( .B1(n17450), .B2(n17458), .A(n17449), .ZN(P3_U2792) );
  AOI22_X1 U20604 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17464), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17460), .ZN(n17451) );
  OAI21_X1 U20605 ( .B1(n17452), .B2(n17458), .A(n17451), .ZN(P3_U2793) );
  AOI22_X1 U20606 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17466), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17460), .ZN(n17453) );
  OAI21_X1 U20607 ( .B1(n17454), .B2(n17462), .A(n17453), .ZN(P3_U2794) );
  AOI22_X1 U20608 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17464), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17465), .ZN(n17455) );
  OAI21_X1 U20609 ( .B1(n17456), .B2(n17458), .A(n17455), .ZN(P3_U2795) );
  AOI22_X1 U20610 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17464), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17465), .ZN(n17457) );
  OAI21_X1 U20611 ( .B1(n17459), .B2(n17458), .A(n17457), .ZN(P3_U2796) );
  AOI22_X1 U20612 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17466), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17460), .ZN(n17461) );
  OAI21_X1 U20613 ( .B1(n17463), .B2(n17462), .A(n17461), .ZN(P3_U2797) );
  AOI222_X1 U20614 ( .A1(n17466), .A2(BUF2_REG_15__SCAN_IN), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17465), .C1(P3_EAX_REG_15__SCAN_IN), 
        .C2(n17464), .ZN(n17467) );
  INV_X1 U20615 ( .A(n17467), .ZN(P3_U2798) );
  INV_X1 U20616 ( .A(n17744), .ZN(n18697) );
  OAI21_X1 U20617 ( .B1(n17468), .B2(n17844), .A(n17843), .ZN(n17469) );
  AOI21_X1 U20618 ( .B1(n18697), .B2(n17492), .A(n17469), .ZN(n17501) );
  OAI21_X1 U20619 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17500), .A(
        n17501), .ZN(n17486) );
  NOR2_X1 U20620 ( .A1(n17679), .A2(n17492), .ZN(n17473) );
  XOR2_X1 U20621 ( .A(n17471), .B(n17470), .Z(n17472) );
  AOI22_X1 U20622 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17486), .B1(
        n17473), .B2(n17472), .ZN(n17485) );
  AOI22_X1 U20623 ( .A1(n18153), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n17649), 
        .B2(n17474), .ZN(n17484) );
  NOR2_X1 U20624 ( .A1(n17753), .A2(n17837), .ZN(n17582) );
  OAI22_X1 U20625 ( .A1(n17475), .A2(n17685), .B1(n17860), .B2(n17848), .ZN(
        n17507) );
  NOR2_X1 U20626 ( .A1(n17861), .A2(n17507), .ZN(n17490) );
  NOR3_X1 U20627 ( .A1(n17582), .A2(n17490), .A3(n17476), .ZN(n17481) );
  AOI211_X1 U20628 ( .C1(n17479), .C2(n17478), .A(n17477), .B(n17756), .ZN(
        n17480) );
  AOI211_X1 U20629 ( .C1(n17482), .C2(n17506), .A(n17481), .B(n17480), .ZN(
        n17483) );
  NAND3_X1 U20630 ( .A1(n17485), .A2(n17484), .A3(n17483), .ZN(P3_U2802) );
  AOI22_X1 U20631 ( .A1(n18165), .A2(P3_REIP_REG_27__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n17486), .ZN(n17496) );
  NOR2_X1 U20632 ( .A1(n17488), .A2(n17487), .ZN(n17489) );
  XOR2_X1 U20633 ( .A(n17489), .B(n17743), .Z(n17862) );
  AOI21_X1 U20634 ( .B1(n17861), .B2(n17491), .A(n17490), .ZN(n17494) );
  NOR3_X1 U20635 ( .A1(n17679), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        n17492), .ZN(n17493) );
  AOI211_X1 U20636 ( .C1(n17738), .C2(n17862), .A(n17494), .B(n17493), .ZN(
        n17495) );
  OAI211_X1 U20637 ( .C1(n17696), .C2(n17497), .A(n17496), .B(n17495), .ZN(
        P3_U2803) );
  AOI21_X1 U20638 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17499), .A(
        n17498), .ZN(n17871) );
  NAND2_X1 U20639 ( .A1(n17696), .A2(n17500), .ZN(n17817) );
  INV_X1 U20640 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18771) );
  NOR2_X1 U20641 ( .A1(n18122), .A2(n18771), .ZN(n17872) );
  NAND3_X1 U20642 ( .A1(n18568), .A2(n17512), .A3(n17511), .ZN(n17502) );
  AOI21_X1 U20643 ( .B1(n17503), .B2(n17502), .A(n17501), .ZN(n17504) );
  AOI211_X1 U20644 ( .C1(n17505), .C2(n17817), .A(n17872), .B(n17504), .ZN(
        n17509) );
  NOR3_X1 U20645 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17880), .A3(
        n17876), .ZN(n17868) );
  AOI22_X1 U20646 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17507), .B1(
        n17506), .B2(n17868), .ZN(n17508) );
  OAI211_X1 U20647 ( .C1(n17871), .C2(n17756), .A(n17509), .B(n17508), .ZN(
        P3_U2804) );
  XOR2_X1 U20648 ( .A(n17880), .B(n17510), .Z(n17889) );
  INV_X1 U20649 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17516) );
  INV_X1 U20650 ( .A(n17679), .ZN(n17633) );
  NAND2_X1 U20651 ( .A1(n17512), .A2(n17633), .ZN(n17528) );
  AOI211_X1 U20652 ( .C1(n17527), .C2(n17516), .A(n17511), .B(n17528), .ZN(
        n17518) );
  OR2_X1 U20653 ( .A1(n18285), .A2(n17512), .ZN(n17544) );
  OAI211_X1 U20654 ( .C1(n17513), .C2(n17844), .A(n17544), .B(n17843), .ZN(
        n17541) );
  AOI21_X1 U20655 ( .B1(n17577), .B2(n17514), .A(n17541), .ZN(n17526) );
  OAI22_X1 U20656 ( .A1(n17526), .A2(n17516), .B1(n17696), .B2(n17515), .ZN(
        n17517) );
  AOI211_X1 U20657 ( .C1(P3_REIP_REG_25__SCAN_IN), .C2(n18165), .A(n17518), 
        .B(n17517), .ZN(n17524) );
  XOR2_X1 U20658 ( .A(n17519), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17886) );
  AOI21_X1 U20659 ( .B1(n17521), .B2(n17743), .A(n17520), .ZN(n17522) );
  XOR2_X1 U20660 ( .A(n17522), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17885) );
  AOI22_X1 U20661 ( .A1(n17753), .A2(n17886), .B1(n17738), .B2(n17885), .ZN(
        n17523) );
  OAI211_X1 U20662 ( .C1(n17848), .C2(n17889), .A(n17524), .B(n17523), .ZN(
        P3_U2805) );
  AOI22_X1 U20663 ( .A1(n17753), .A2(n17893), .B1(n17837), .B2(n17894), .ZN(
        n17547) );
  NAND2_X1 U20664 ( .A1(n18153), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17525) );
  OAI221_X1 U20665 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17528), .C1(
        n17527), .C2(n17526), .A(n17525), .ZN(n17532) );
  AOI21_X1 U20666 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17530), .A(
        n17529), .ZN(n17904) );
  NAND2_X1 U20667 ( .A1(n17535), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17890) );
  OAI22_X1 U20668 ( .A1(n17904), .A2(n17756), .B1(n17548), .B2(n17890), .ZN(
        n17531) );
  AOI211_X1 U20669 ( .C1(n17649), .C2(n17533), .A(n17532), .B(n17531), .ZN(
        n17534) );
  OAI21_X1 U20670 ( .B1(n17547), .B2(n17535), .A(n17534), .ZN(P3_U2806) );
  AOI22_X1 U20671 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17743), .B1(
        n17537), .B2(n17556), .ZN(n17538) );
  NAND2_X1 U20672 ( .A1(n17536), .A2(n17538), .ZN(n17539) );
  XOR2_X1 U20673 ( .A(n17539), .B(n17898), .Z(n17905) );
  AOI22_X1 U20674 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17541), .B1(
        n17540), .B2(n17817), .ZN(n17542) );
  NAND2_X1 U20675 ( .A1(n18165), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17909) );
  OAI211_X1 U20676 ( .C1(n17544), .C2(n17543), .A(n17542), .B(n17909), .ZN(
        n17545) );
  AOI21_X1 U20677 ( .B1(n17738), .B2(n17905), .A(n17545), .ZN(n17546) );
  OAI221_X1 U20678 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17548), 
        .C1(n17898), .C2(n17547), .A(n17546), .ZN(P3_U2807) );
  INV_X1 U20679 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17563) );
  NAND2_X1 U20680 ( .A1(n17551), .A2(n17633), .ZN(n17564) );
  AOI221_X1 U20681 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C1(n17563), .C2(n17552), .A(
        n17564), .ZN(n17554) );
  AOI21_X1 U20682 ( .B1(n17630), .B2(n17549), .A(n17803), .ZN(n17550) );
  OAI21_X1 U20683 ( .B1(n17551), .B2(n17744), .A(n17550), .ZN(n17581) );
  AOI21_X1 U20684 ( .B1(n17577), .B2(n17574), .A(n17581), .ZN(n17562) );
  NAND2_X1 U20685 ( .A1(n18153), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17927) );
  OAI21_X1 U20686 ( .B1(n17562), .B2(n17552), .A(n17927), .ZN(n17553) );
  AOI211_X1 U20687 ( .C1(n17555), .C2(n17649), .A(n17554), .B(n17553), .ZN(
        n17561) );
  NOR2_X1 U20688 ( .A1(n17609), .A2(n17911), .ZN(n17919) );
  NOR2_X1 U20689 ( .A1(n17913), .A2(n17685), .ZN(n17652) );
  NOR2_X1 U20690 ( .A1(n17993), .A2(n17848), .ZN(n17651) );
  NOR2_X1 U20691 ( .A1(n17652), .A2(n17651), .ZN(n17640) );
  OAI21_X1 U20692 ( .B1(n17582), .B2(n17919), .A(n17640), .ZN(n17571) );
  INV_X1 U20693 ( .A(n17556), .ZN(n17557) );
  OAI221_X1 U20694 ( .B1(n17557), .B2(n17919), .C1(n17557), .C2(n17626), .A(
        n17536), .ZN(n17558) );
  XOR2_X1 U20695 ( .A(n17929), .B(n17558), .Z(n17926) );
  AOI22_X1 U20696 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17571), .B1(
        n17738), .B2(n17926), .ZN(n17560) );
  NAND3_X1 U20697 ( .A1(n17620), .A2(n17919), .A3(n17929), .ZN(n17559) );
  NAND3_X1 U20698 ( .A1(n17561), .A2(n17560), .A3(n17559), .ZN(P3_U2808) );
  NAND2_X1 U20699 ( .A1(n17937), .A2(n17932), .ZN(n17943) );
  NAND3_X1 U20700 ( .A1(n17963), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17620), .ZN(n17598) );
  NAND2_X1 U20701 ( .A1(n18165), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n17941) );
  OAI221_X1 U20702 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17564), .C1(
        n17563), .C2(n17562), .A(n17941), .ZN(n17565) );
  AOI21_X1 U20703 ( .B1(n17649), .B2(n17566), .A(n17565), .ZN(n17573) );
  INV_X1 U20704 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17931) );
  NOR3_X1 U20705 ( .A1(n17743), .A2(n17931), .A3(n17567), .ZN(n17593) );
  INV_X1 U20706 ( .A(n17568), .ZN(n17607) );
  AOI22_X1 U20707 ( .A1(n17937), .A2(n17593), .B1(n17607), .B2(n17569), .ZN(
        n17570) );
  XOR2_X1 U20708 ( .A(n17932), .B(n17570), .Z(n17940) );
  AOI22_X1 U20709 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17571), .B1(
        n17738), .B2(n17940), .ZN(n17572) );
  OAI211_X1 U20710 ( .C1(n17943), .C2(n17598), .A(n17573), .B(n17572), .ZN(
        P3_U2809) );
  OR2_X1 U20711 ( .A1(n20876), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17953) );
  OAI21_X1 U20712 ( .B1(n17575), .B2(n18285), .A(n17574), .ZN(n17580) );
  INV_X1 U20713 ( .A(n17576), .ZN(n17578) );
  NAND2_X1 U20714 ( .A1(n18165), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17951) );
  OAI221_X1 U20715 ( .B1(n17578), .B2(n17696), .C1(n17578), .C2(n17500), .A(
        n17951), .ZN(n17579) );
  AOI21_X1 U20716 ( .B1(n17581), .B2(n17580), .A(n17579), .ZN(n17585) );
  NOR2_X1 U20717 ( .A1(n17609), .A2(n17931), .ZN(n17933) );
  NAND2_X1 U20718 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17933), .ZN(
        n17915) );
  INV_X1 U20719 ( .A(n17915), .ZN(n17945) );
  OAI21_X1 U20720 ( .B1(n17582), .B2(n17945), .A(n17640), .ZN(n17595) );
  OAI221_X1 U20721 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17606), 
        .C1(n20876), .C2(n17593), .A(n17536), .ZN(n17583) );
  XNOR2_X1 U20722 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17583), .ZN(
        n17949) );
  AOI22_X1 U20723 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17595), .B1(
        n17738), .B2(n17949), .ZN(n17584) );
  OAI211_X1 U20724 ( .C1(n17598), .C2(n17953), .A(n17585), .B(n17584), .ZN(
        P3_U2810) );
  NAND2_X1 U20725 ( .A1(n17587), .A2(n17633), .ZN(n17603) );
  AOI211_X1 U20726 ( .C1(n17602), .C2(n17590), .A(n17586), .B(n17603), .ZN(
        n17592) );
  OAI21_X1 U20727 ( .B1(n17587), .B2(n17744), .A(n17843), .ZN(n17617) );
  AOI21_X1 U20728 ( .B1(n17630), .B2(n17588), .A(n17617), .ZN(n17601) );
  OAI22_X1 U20729 ( .A1(n17601), .A2(n17590), .B1(n17696), .B2(n17589), .ZN(
        n17591) );
  AOI211_X1 U20730 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n18165), .A(n17592), 
        .B(n17591), .ZN(n17597) );
  AOI21_X1 U20731 ( .B1(n17606), .B2(n17607), .A(n17593), .ZN(n17594) );
  XOR2_X1 U20732 ( .A(n20876), .B(n17594), .Z(n17954) );
  AOI22_X1 U20733 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17595), .B1(
        n17738), .B2(n17954), .ZN(n17596) );
  OAI211_X1 U20734 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17598), .A(
        n17597), .B(n17596), .ZN(P3_U2811) );
  INV_X1 U20735 ( .A(n17620), .ZN(n17641) );
  OAI21_X1 U20736 ( .B1(n17641), .B2(n17963), .A(n17640), .ZN(n17599) );
  INV_X1 U20737 ( .A(n17599), .ZN(n17623) );
  NAND2_X1 U20738 ( .A1(n18165), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17600) );
  OAI221_X1 U20739 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17603), .C1(
        n17602), .C2(n17601), .A(n17600), .ZN(n17604) );
  AOI21_X1 U20740 ( .B1(n17649), .B2(n17605), .A(n17604), .ZN(n17611) );
  AOI21_X1 U20741 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17627), .A(
        n17606), .ZN(n17608) );
  XOR2_X1 U20742 ( .A(n17608), .B(n17607), .Z(n17971) );
  NOR2_X1 U20743 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17609), .ZN(
        n17970) );
  AOI22_X1 U20744 ( .A1(n17738), .A2(n17971), .B1(n17620), .B2(n17970), .ZN(
        n17610) );
  OAI211_X1 U20745 ( .C1(n17623), .C2(n17931), .A(n17611), .B(n17610), .ZN(
        P3_U2812) );
  OAI21_X1 U20746 ( .B1(n18285), .B2(n17613), .A(n17612), .ZN(n17616) );
  INV_X2 U20747 ( .A(n17817), .ZN(n17840) );
  OAI22_X1 U20748 ( .A1(n17840), .A2(n17614), .B1(n18122), .B2(n18753), .ZN(
        n17615) );
  AOI21_X1 U20749 ( .B1(n17617), .B2(n17616), .A(n17615), .ZN(n17622) );
  OAI21_X1 U20750 ( .B1(n17619), .B2(n17964), .A(n17618), .ZN(n17976) );
  NOR2_X1 U20751 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17982), .ZN(
        n17975) );
  AOI22_X1 U20752 ( .A1(n17738), .A2(n17976), .B1(n17620), .B2(n17975), .ZN(
        n17621) );
  OAI211_X1 U20753 ( .C1(n17623), .C2(n17964), .A(n17622), .B(n17621), .ZN(
        P3_U2813) );
  NOR2_X1 U20754 ( .A1(n17743), .A2(n17624), .ZN(n17727) );
  INV_X1 U20755 ( .A(n17727), .ZN(n17625) );
  OAI22_X1 U20756 ( .A1(n17627), .A2(n17626), .B1(n17625), .B2(n17969), .ZN(
        n17628) );
  XOR2_X1 U20757 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17628), .Z(
        n17984) );
  OAI21_X1 U20758 ( .B1(n17634), .B2(n17744), .A(n17843), .ZN(n17659) );
  AOI21_X1 U20759 ( .B1(n17630), .B2(n17629), .A(n17659), .ZN(n17644) );
  OAI22_X1 U20760 ( .A1(n17644), .A2(n17632), .B1(n17696), .B2(n17631), .ZN(
        n17638) );
  NAND2_X1 U20761 ( .A1(n17634), .A2(n17633), .ZN(n17646) );
  OAI21_X1 U20762 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17635), .ZN(n17636) );
  OAI22_X1 U20763 ( .A1(n18122), .A2(n18750), .B1(n17646), .B2(n17636), .ZN(
        n17637) );
  AOI211_X1 U20764 ( .C1(n17738), .C2(n17984), .A(n17638), .B(n17637), .ZN(
        n17639) );
  OAI221_X1 U20765 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17641), 
        .C1(n17982), .C2(n17640), .A(n17639), .ZN(P3_U2814) );
  NAND2_X1 U20766 ( .A1(n17670), .A2(n17727), .ZN(n17660) );
  NAND3_X1 U20767 ( .A1(n17689), .A2(n17743), .A3(n18000), .ZN(n17661) );
  NOR2_X1 U20768 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18042), .ZN(
        n18017) );
  AOI221_X1 U20769 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17660), 
        .C1(n18005), .C2(n17661), .A(n18017), .ZN(n17642) );
  XOR2_X1 U20770 ( .A(n17642), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Z(
        n17996) );
  INV_X1 U20771 ( .A(n17996), .ZN(n17655) );
  NAND2_X1 U20772 ( .A1(n18165), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n17643) );
  OAI221_X1 U20773 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17646), .C1(
        n17645), .C2(n17644), .A(n17643), .ZN(n17647) );
  AOI21_X1 U20774 ( .B1(n17649), .B2(n17648), .A(n17647), .ZN(n17654) );
  NAND2_X1 U20775 ( .A1(n17663), .A2(n17650), .ZN(n17991) );
  INV_X1 U20776 ( .A(n17987), .ZN(n18004) );
  OAI21_X1 U20777 ( .B1(n17711), .B2(n18004), .A(n17650), .ZN(n17994) );
  AOI22_X1 U20778 ( .A1(n17652), .A2(n17991), .B1(n17651), .B2(n17994), .ZN(
        n17653) );
  OAI211_X1 U20779 ( .C1(n17756), .C2(n17655), .A(n17654), .B(n17653), .ZN(
        P3_U2815) );
  NOR2_X1 U20780 ( .A1(n18285), .A2(n17678), .ZN(n17707) );
  AOI21_X1 U20781 ( .B1(n17656), .B2(n17707), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17657) );
  INV_X1 U20782 ( .A(n17657), .ZN(n17658) );
  AOI22_X1 U20783 ( .A1(n18153), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n17659), 
        .B2(n17658), .ZN(n17668) );
  AOI21_X1 U20784 ( .B1(n17661), .B2(n17660), .A(n18017), .ZN(n17662) );
  XOR2_X1 U20785 ( .A(n17662), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n18012) );
  OAI21_X1 U20786 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17664), .A(
        n17663), .ZN(n18009) );
  NOR2_X1 U20787 ( .A1(n17711), .A2(n18003), .ZN(n18023) );
  NAND2_X1 U20788 ( .A1(n17987), .A2(n18044), .ZN(n17665) );
  OAI221_X1 U20789 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18023), .A(n17665), .ZN(
        n18016) );
  OAI22_X1 U20790 ( .A1(n17685), .A2(n18009), .B1(n17848), .B2(n18016), .ZN(
        n17666) );
  AOI21_X1 U20791 ( .B1(n17738), .B2(n18012), .A(n17666), .ZN(n17667) );
  OAI211_X1 U20792 ( .C1(n17840), .C2(n17669), .A(n17668), .B(n17667), .ZN(
        P3_U2816) );
  AOI22_X1 U20793 ( .A1(n17671), .A2(n17670), .B1(n17743), .B2(n18042), .ZN(
        n17674) );
  INV_X1 U20794 ( .A(n17672), .ZN(n17673) );
  NOR2_X1 U20795 ( .A1(n17674), .A2(n17673), .ZN(n17675) );
  XOR2_X1 U20796 ( .A(n17675), .B(n18000), .Z(n18032) );
  AOI21_X1 U20797 ( .B1(n18697), .B2(n17678), .A(n17803), .ZN(n17676) );
  OAI21_X1 U20798 ( .B1(n17677), .B2(n17844), .A(n17676), .ZN(n17693) );
  NOR2_X1 U20799 ( .A1(n17679), .A2(n17678), .ZN(n17692) );
  OAI211_X1 U20800 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17692), .B(n17680), .ZN(n17682) );
  NAND2_X1 U20801 ( .A1(n18153), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17681) );
  OAI211_X1 U20802 ( .C1(n17696), .C2(n17683), .A(n17682), .B(n17681), .ZN(
        n17684) );
  AOI21_X1 U20803 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17693), .A(
        n17684), .ZN(n17688) );
  OAI22_X1 U20804 ( .A1(n17686), .A2(n17685), .B1(n18023), .B2(n17848), .ZN(
        n17698) );
  NOR2_X1 U20805 ( .A1(n17741), .A2(n18036), .ZN(n17699) );
  AOI22_X1 U20806 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17698), .B1(
        n18017), .B2(n17699), .ZN(n17687) );
  OAI211_X1 U20807 ( .C1(n17756), .C2(n18032), .A(n17688), .B(n17687), .ZN(
        P3_U2817) );
  AND2_X1 U20808 ( .A1(n18051), .A2(n17727), .ZN(n17703) );
  AOI22_X1 U20809 ( .A1(n17703), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n17689), .B2(n17743), .ZN(n17690) );
  XOR2_X1 U20810 ( .A(n18042), .B(n17690), .Z(n18039) );
  INV_X1 U20811 ( .A(n18039), .ZN(n17701) );
  AOI22_X1 U20812 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17693), .B1(
        n17692), .B2(n17691), .ZN(n17694) );
  NAND2_X1 U20813 ( .A1(n18153), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18040) );
  OAI211_X1 U20814 ( .C1(n17696), .C2(n17695), .A(n17694), .B(n18040), .ZN(
        n17697) );
  AOI221_X1 U20815 ( .B1(n17699), .B2(n18042), .C1(n17698), .C2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17697), .ZN(n17700) );
  OAI21_X1 U20816 ( .B1(n17701), .B2(n17756), .A(n17700), .ZN(P3_U2818) );
  INV_X1 U20817 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18019) );
  NAND2_X1 U20818 ( .A1(n18051), .A2(n18019), .ZN(n18056) );
  NAND2_X1 U20819 ( .A1(n12781), .A2(n12780), .ZN(n17722) );
  INV_X1 U20820 ( .A(n17722), .ZN(n17704) );
  AND2_X1 U20821 ( .A1(n17702), .A2(n20851), .ZN(n17728) );
  AOI21_X1 U20822 ( .B1(n17704), .B2(n17728), .A(n17703), .ZN(n17705) );
  XOR2_X1 U20823 ( .A(n18019), .B(n17705), .Z(n18043) );
  INV_X1 U20824 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18740) );
  NOR2_X1 U20825 ( .A1(n18122), .A2(n18740), .ZN(n17710) );
  NAND3_X1 U20826 ( .A1(n18568), .A2(n17771), .A3(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17760) );
  INV_X1 U20827 ( .A(n17760), .ZN(n17731) );
  NAND2_X1 U20828 ( .A1(n17843), .A2(n17744), .ZN(n17836) );
  AOI22_X1 U20829 ( .A1(n17718), .A2(n17731), .B1(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17836), .ZN(n17708) );
  OAI22_X1 U20830 ( .A1(n17708), .A2(n17707), .B1(n17840), .B2(n17706), .ZN(
        n17709) );
  AOI211_X1 U20831 ( .C1(n17738), .C2(n18043), .A(n17710), .B(n17709), .ZN(
        n17714) );
  NOR2_X1 U20832 ( .A1(n18051), .A2(n17741), .ZN(n17723) );
  AOI22_X1 U20833 ( .A1(n17712), .A2(n17753), .B1(n17837), .B2(n17711), .ZN(
        n17740) );
  INV_X1 U20834 ( .A(n17740), .ZN(n17724) );
  OAI21_X1 U20835 ( .B1(n17723), .B2(n17724), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17713) );
  OAI211_X1 U20836 ( .C1(n17741), .C2(n18056), .A(n17714), .B(n17713), .ZN(
        P3_U2819) );
  AOI22_X1 U20837 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17727), .B1(
        n17728), .B2(n12781), .ZN(n17715) );
  XOR2_X1 U20838 ( .A(n17715), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .Z(
        n18064) );
  AOI22_X1 U20839 ( .A1(n17716), .A2(n17731), .B1(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17836), .ZN(n17717) );
  AOI21_X1 U20840 ( .B1(n17731), .B2(n17718), .A(n17717), .ZN(n17720) );
  NOR2_X1 U20841 ( .A1(n18122), .A2(n18738), .ZN(n17719) );
  AOI211_X1 U20842 ( .C1(n17721), .C2(n17817), .A(n17720), .B(n17719), .ZN(
        n17726) );
  AOI22_X1 U20843 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17724), .B1(
        n17723), .B2(n17722), .ZN(n17725) );
  OAI211_X1 U20844 ( .C1(n18064), .C2(n17756), .A(n17726), .B(n17725), .ZN(
        P3_U2820) );
  NOR2_X1 U20845 ( .A1(n17728), .A2(n17727), .ZN(n17729) );
  XOR2_X1 U20846 ( .A(n17729), .B(n12781), .Z(n18071) );
  NOR2_X1 U20847 ( .A1(n18122), .A2(n18736), .ZN(n17737) );
  NOR2_X1 U20848 ( .A1(n17730), .A2(n17760), .ZN(n17735) );
  AOI22_X1 U20849 ( .A1(n17732), .A2(n17731), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17836), .ZN(n17734) );
  OAI22_X1 U20850 ( .A1(n17735), .A2(n17734), .B1(n17840), .B2(n17733), .ZN(
        n17736) );
  AOI211_X1 U20851 ( .C1(n17738), .C2(n18071), .A(n17737), .B(n17736), .ZN(
        n17739) );
  OAI221_X1 U20852 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17741), .C1(
        n12781), .C2(n17740), .A(n17739), .ZN(P3_U2821) );
  AOI21_X1 U20853 ( .B1(n17743), .B2(n17750), .A(n17742), .ZN(n18092) );
  OAI21_X1 U20854 ( .B1(n17746), .B2(n17744), .A(n17843), .ZN(n17766) );
  NOR2_X1 U20855 ( .A1(n18122), .A2(n18734), .ZN(n18083) );
  OAI211_X1 U20856 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n17746), .B(n17745), .ZN(n17747)
         );
  OAI22_X1 U20857 ( .A1(n17840), .A2(n17748), .B1(n18285), .B2(n17747), .ZN(
        n17749) );
  AOI211_X1 U20858 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17766), .A(
        n18083), .B(n17749), .ZN(n17755) );
  INV_X1 U20859 ( .A(n17750), .ZN(n18088) );
  AOI21_X1 U20860 ( .B1(n17752), .B2(n20851), .A(n17751), .ZN(n18086) );
  AOI22_X1 U20861 ( .A1(n17753), .A2(n18088), .B1(n17837), .B2(n18086), .ZN(
        n17754) );
  OAI211_X1 U20862 ( .C1(n18092), .C2(n17756), .A(n17755), .B(n17754), .ZN(
        P3_U2822) );
  NAND2_X1 U20863 ( .A1(n17758), .A2(n17757), .ZN(n17759) );
  XOR2_X1 U20864 ( .A(n17759), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18100) );
  OAI22_X1 U20865 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17760), .B1(
        n18122), .B2(n18732), .ZN(n17761) );
  AOI21_X1 U20866 ( .B1(n17762), .B2(n17817), .A(n17761), .ZN(n17768) );
  INV_X1 U20867 ( .A(n17763), .ZN(n17764) );
  AOI21_X1 U20868 ( .B1(n18094), .B2(n17765), .A(n17764), .ZN(n18096) );
  AOI22_X1 U20869 ( .A1(n17833), .A2(n18096), .B1(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17766), .ZN(n17767) );
  OAI211_X1 U20870 ( .C1(n17848), .C2(n18100), .A(n17768), .B(n17767), .ZN(
        P3_U2823) );
  AOI21_X1 U20871 ( .B1(n18095), .B2(n17770), .A(n17769), .ZN(n18105) );
  NAND2_X1 U20872 ( .A1(n18568), .A2(n17771), .ZN(n17778) );
  OAI21_X1 U20873 ( .B1(n17772), .B2(n18285), .A(n17836), .ZN(n17794) );
  AOI21_X1 U20874 ( .B1(n17775), .B2(n17774), .A(n17773), .ZN(n18104) );
  AOI22_X1 U20875 ( .A1(n17833), .A2(n18104), .B1(n18153), .B2(
        P3_REIP_REG_6__SCAN_IN), .ZN(n17776) );
  OAI221_X1 U20876 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17778), .C1(
        n17777), .C2(n17794), .A(n17776), .ZN(n17779) );
  AOI21_X1 U20877 ( .B1(n17837), .B2(n18105), .A(n17779), .ZN(n17780) );
  OAI21_X1 U20878 ( .B1(n17840), .B2(n17781), .A(n17780), .ZN(P3_U2824) );
  AOI21_X1 U20879 ( .B1(n17782), .B2(n17843), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17795) );
  OAI21_X1 U20880 ( .B1(n17785), .B2(n17783), .A(n17784), .ZN(n17787) );
  XOR2_X1 U20881 ( .A(n17787), .B(n17786), .Z(n18110) );
  AOI22_X1 U20882 ( .A1(n17833), .A2(n18110), .B1(n18153), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17793) );
  AOI21_X1 U20883 ( .B1(n17790), .B2(n17789), .A(n17788), .ZN(n18109) );
  AOI22_X1 U20884 ( .A1(n17837), .A2(n18109), .B1(n17791), .B2(n17817), .ZN(
        n17792) );
  OAI211_X1 U20885 ( .C1(n17795), .C2(n17794), .A(n17793), .B(n17792), .ZN(
        P3_U2825) );
  OAI21_X1 U20886 ( .B1(n17798), .B2(n17797), .A(n17796), .ZN(n17799) );
  XOR2_X1 U20887 ( .A(n17799), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n18121) );
  OAI21_X1 U20888 ( .B1(n17801), .B2(n9630), .A(n17800), .ZN(n17802) );
  XOR2_X1 U20889 ( .A(n17802), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n18127) );
  OAI22_X1 U20890 ( .A1(n17847), .A2(n18127), .B1(n18122), .B2(n18726), .ZN(
        n17808) );
  AOI21_X1 U20891 ( .B1(n18697), .B2(n17804), .A(n17803), .ZN(n17821) );
  OAI22_X1 U20892 ( .A1(n17840), .A2(n17806), .B1(n17821), .B2(n17805), .ZN(
        n17807) );
  AOI211_X1 U20893 ( .C1(n18568), .C2(n17809), .A(n17808), .B(n17807), .ZN(
        n17810) );
  OAI21_X1 U20894 ( .B1(n17848), .B2(n18121), .A(n17810), .ZN(P3_U2826) );
  AOI21_X1 U20895 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17843), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17822) );
  AOI21_X1 U20896 ( .B1(n17813), .B2(n17812), .A(n17811), .ZN(n18129) );
  AOI22_X1 U20897 ( .A1(n17833), .A2(n18129), .B1(n18153), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17820) );
  AOI21_X1 U20898 ( .B1(n17816), .B2(n17815), .A(n17814), .ZN(n18130) );
  AOI22_X1 U20899 ( .A1(n17837), .A2(n18130), .B1(n17818), .B2(n17817), .ZN(
        n17819) );
  OAI211_X1 U20900 ( .C1(n17822), .C2(n17821), .A(n17820), .B(n17819), .ZN(
        P3_U2827) );
  NAND2_X1 U20901 ( .A1(n18153), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18146) );
  INV_X1 U20902 ( .A(n18146), .ZN(n17829) );
  XNOR2_X1 U20903 ( .A(n17826), .B(n17825), .ZN(n18148) );
  OAI22_X1 U20904 ( .A1(n17840), .A2(n17827), .B1(n17848), .B2(n18148), .ZN(
        n17828) );
  AOI211_X1 U20905 ( .C1(n17833), .C2(n18141), .A(n17829), .B(n17828), .ZN(
        n17830) );
  OAI221_X1 U20906 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18285), .C1(
        n17831), .C2(n17843), .A(n17830), .ZN(P3_U2828) );
  AOI21_X1 U20907 ( .B1(n17841), .B2(n17834), .A(n17832), .ZN(n18149) );
  AOI22_X1 U20908 ( .A1(n17833), .A2(n18149), .B1(n18153), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17839) );
  NOR2_X1 U20909 ( .A1(n17842), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17835) );
  XNOR2_X1 U20910 ( .A(n17835), .B(n17834), .ZN(n18151) );
  AOI22_X1 U20911 ( .A1(n17837), .A2(n18151), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17836), .ZN(n17838) );
  OAI211_X1 U20912 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n17840), .A(
        n17839), .B(n17838), .ZN(P3_U2829) );
  OAI21_X1 U20913 ( .B1(n17842), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17841), .ZN(n18170) );
  INV_X1 U20914 ( .A(n18170), .ZN(n18172) );
  NAND3_X1 U20915 ( .A1(n18801), .A2(n17844), .A3(n17843), .ZN(n17845) );
  AOI22_X1 U20916 ( .A1(n18165), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17845), .ZN(n17846) );
  OAI221_X1 U20917 ( .B1(n18172), .B2(n17848), .C1(n18170), .C2(n17847), .A(
        n17846), .ZN(P3_U2830) );
  AOI22_X1 U20918 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18162), .B1(
        n17849), .B2(n17892), .ZN(n17866) );
  NAND2_X1 U20919 ( .A1(n17850), .A2(n18021), .ZN(n17960) );
  INV_X1 U20920 ( .A(n17919), .ZN(n17851) );
  NOR2_X1 U20921 ( .A1(n17960), .A2(n17851), .ZN(n17853) );
  OAI21_X1 U20922 ( .B1(n17929), .B2(n18633), .A(n17852), .ZN(n17922) );
  INV_X1 U20923 ( .A(n18078), .ZN(n18136) );
  AOI21_X1 U20924 ( .B1(n17853), .B2(n17922), .A(n18136), .ZN(n17895) );
  AOI22_X1 U20925 ( .A1(n18633), .A2(n17854), .B1(n18078), .B2(n17876), .ZN(
        n17856) );
  OAI211_X1 U20926 ( .C1(n18634), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17856), .B(n17855), .ZN(n17857) );
  AOI211_X1 U20927 ( .C1(n18026), .C2(n17858), .A(n17895), .B(n17857), .ZN(
        n17859) );
  OAI21_X1 U20928 ( .B1(n17860), .B2(n18626), .A(n17859), .ZN(n17869) );
  AOI211_X1 U20929 ( .C1(n18658), .C2(n17875), .A(n17861), .B(n17869), .ZN(
        n17865) );
  AOI22_X1 U20930 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18156), .B1(
        n18072), .B2(n17862), .ZN(n17864) );
  NAND2_X1 U20931 ( .A1(n18153), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17863) );
  OAI211_X1 U20932 ( .C1(n17866), .C2(n17865), .A(n17864), .B(n17863), .ZN(
        P3_U2835) );
  NOR2_X1 U20933 ( .A1(n17912), .A2(n17867), .ZN(n17907) );
  AOI22_X1 U20934 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17869), .B1(
        n17868), .B2(n17907), .ZN(n17870) );
  OAI22_X1 U20935 ( .A1(n17871), .A2(n18091), .B1(n17870), .B2(n18154), .ZN(
        n17873) );
  NOR2_X1 U20936 ( .A1(n17873), .A2(n17872), .ZN(n17874) );
  OAI21_X1 U20937 ( .B1(n17875), .B2(n18119), .A(n17874), .ZN(P3_U2836) );
  NOR2_X1 U20938 ( .A1(n18122), .A2(n18769), .ZN(n17884) );
  INV_X1 U20939 ( .A(n17959), .ZN(n17917) );
  AOI21_X1 U20940 ( .B1(n17878), .B2(n17917), .A(n18648), .ZN(n17899) );
  AOI211_X1 U20941 ( .C1(n18081), .C2(n17876), .A(n17899), .B(n17895), .ZN(
        n17882) );
  NAND3_X1 U20942 ( .A1(n17879), .A2(n17878), .A3(n17877), .ZN(n17881) );
  AOI221_X1 U20943 ( .B1(n17882), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), 
        .C1(n17881), .C2(n17880), .A(n18154), .ZN(n17883) );
  AOI211_X1 U20944 ( .C1(n18156), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17884), .B(n17883), .ZN(n17888) );
  AOI22_X1 U20945 ( .A1(n18087), .A2(n17886), .B1(n18072), .B2(n17885), .ZN(
        n17887) );
  OAI211_X1 U20946 ( .C1(n18171), .C2(n17889), .A(n17888), .B(n17887), .ZN(
        P3_U2837) );
  INV_X1 U20947 ( .A(n17890), .ZN(n17891) );
  AOI22_X1 U20948 ( .A1(n18165), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n17892), 
        .B2(n17891), .ZN(n17903) );
  AOI22_X1 U20949 ( .A1(n17918), .A2(n17894), .B1(n18026), .B2(n17893), .ZN(
        n17897) );
  INV_X1 U20950 ( .A(n17895), .ZN(n17896) );
  NAND3_X1 U20951 ( .A1(n17897), .A2(n18119), .A3(n17896), .ZN(n17901) );
  NOR3_X1 U20952 ( .A1(n17899), .A2(n17898), .A3(n17901), .ZN(n17900) );
  NOR2_X1 U20953 ( .A1(n18165), .A2(n17900), .ZN(n17906) );
  OAI211_X1 U20954 ( .C1(n18081), .C2(n17901), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17906), .ZN(n17902) );
  OAI211_X1 U20955 ( .C1(n17904), .C2(n18091), .A(n17903), .B(n17902), .ZN(
        P3_U2838) );
  INV_X1 U20956 ( .A(n17905), .ZN(n17910) );
  OAI221_X1 U20957 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17907), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n18119), .A(n17906), .ZN(
        n17908) );
  OAI211_X1 U20958 ( .C1(n17910), .C2(n18091), .A(n17909), .B(n17908), .ZN(
        P3_U2839) );
  AOI221_X1 U20959 ( .B1(n17912), .B2(n17929), .C1(n17911), .C2(n17929), .A(
        n18154), .ZN(n17925) );
  NOR2_X1 U20960 ( .A1(n17913), .A2(n18045), .ZN(n17992) );
  AOI21_X1 U20961 ( .B1(n17918), .B2(n17914), .A(n17992), .ZN(n17934) );
  OAI21_X1 U20962 ( .B1(n17960), .B2(n17915), .A(n18658), .ZN(n17916) );
  OAI221_X1 U20963 ( .B1(n18648), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), 
        .C1(n18648), .C2(n17917), .A(n17916), .ZN(n17947) );
  NOR2_X1 U20964 ( .A1(n17918), .A2(n18026), .ZN(n18050) );
  OAI22_X1 U20965 ( .A1(n18634), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n17919), .B2(n18050), .ZN(n17920) );
  NOR2_X1 U20966 ( .A1(n17947), .A2(n17920), .ZN(n17936) );
  AOI22_X1 U20967 ( .A1(n18654), .A2(n17921), .B1(n17932), .B2(n18059), .ZN(
        n17923) );
  NAND4_X1 U20968 ( .A1(n17934), .A2(n17936), .A3(n17923), .A4(n17922), .ZN(
        n17924) );
  AOI22_X1 U20969 ( .A1(n18072), .A2(n17926), .B1(n17925), .B2(n17924), .ZN(
        n17928) );
  OAI211_X1 U20970 ( .C1(n18119), .C2(n17929), .A(n17928), .B(n17927), .ZN(
        P3_U2840) );
  NOR2_X1 U20971 ( .A1(n18165), .A2(n17932), .ZN(n17939) );
  NOR2_X1 U20972 ( .A1(n18654), .A2(n18633), .ZN(n18155) );
  AOI21_X1 U20973 ( .B1(n17980), .B2(n17933), .A(n18635), .ZN(n17935) );
  NAND2_X1 U20974 ( .A1(n18162), .A2(n17934), .ZN(n17981) );
  NOR2_X1 U20975 ( .A1(n17935), .A2(n17981), .ZN(n17944) );
  OAI211_X1 U20976 ( .C1(n17937), .C2(n18155), .A(n17936), .B(n17944), .ZN(
        n17938) );
  AOI22_X1 U20977 ( .A1(n18072), .A2(n17940), .B1(n17939), .B2(n17938), .ZN(
        n17942) );
  OAI211_X1 U20978 ( .C1(n17943), .C2(n17957), .A(n17942), .B(n17941), .ZN(
        P3_U2841) );
  NAND2_X1 U20979 ( .A1(n20876), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17948) );
  OAI21_X1 U20980 ( .B1(n17945), .B2(n18050), .A(n17944), .ZN(n17946) );
  OAI21_X1 U20981 ( .B1(n17947), .B2(n17946), .A(n18122), .ZN(n17956) );
  OAI21_X1 U20982 ( .B1(n18155), .B2(n17948), .A(n17956), .ZN(n17950) );
  AOI22_X1 U20983 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17950), .B1(
        n18072), .B2(n17949), .ZN(n17952) );
  OAI211_X1 U20984 ( .C1(n17957), .C2(n17953), .A(n17952), .B(n17951), .ZN(
        P3_U2842) );
  AOI22_X1 U20985 ( .A1(n18153), .A2(P3_REIP_REG_19__SCAN_IN), .B1(n18072), 
        .B2(n17954), .ZN(n17955) );
  OAI221_X1 U20986 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17957), 
        .C1(n20876), .C2(n17956), .A(n17955), .ZN(P3_U2843) );
  NAND2_X1 U20987 ( .A1(n18633), .A2(n18818), .ZN(n18137) );
  INV_X1 U20988 ( .A(n18137), .ZN(n17958) );
  AOI211_X1 U20989 ( .C1(n18654), .C2(n17959), .A(n17958), .B(n17981), .ZN(
        n17962) );
  OAI21_X1 U20990 ( .B1(n17982), .B2(n17960), .A(n18078), .ZN(n17961) );
  OAI211_X1 U20991 ( .C1(n17963), .C2(n18050), .A(n17962), .B(n17961), .ZN(
        n17974) );
  OAI221_X1 U20992 ( .B1(n17974), .B2(n18078), .C1(n17974), .C2(n17964), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17973) );
  OAI22_X1 U20993 ( .A1(n18115), .A2(n18648), .B1(n17965), .B2(n18138), .ZN(
        n18128) );
  NAND2_X1 U20994 ( .A1(n17966), .A2(n18128), .ZN(n18101) );
  NOR2_X1 U20995 ( .A1(n17967), .A2(n18101), .ZN(n18001) );
  OAI21_X1 U20996 ( .B1(n18001), .B2(n17968), .A(n18162), .ZN(n18075) );
  NOR2_X1 U20997 ( .A1(n17969), .A2(n18075), .ZN(n17983) );
  AOI22_X1 U20998 ( .A1(n18072), .A2(n17971), .B1(n17983), .B2(n17970), .ZN(
        n17972) );
  OAI221_X1 U20999 ( .B1(n18165), .B2(n17973), .C1(n18122), .C2(n18754), .A(
        n17972), .ZN(P3_U2844) );
  NAND2_X1 U21000 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17974), .ZN(
        n17978) );
  AOI22_X1 U21001 ( .A1(n18072), .A2(n17976), .B1(n17983), .B2(n17975), .ZN(
        n17977) );
  OAI221_X1 U21002 ( .B1(n18153), .B2(n17978), .C1(n18122), .C2(n18753), .A(
        n17977), .ZN(P3_U2845) );
  NAND2_X1 U21003 ( .A1(n18658), .A2(n20851), .ZN(n18067) );
  OAI21_X1 U21004 ( .B1(n18076), .B2(n18077), .A(n18658), .ZN(n18057) );
  OAI211_X1 U21005 ( .C1(n18020), .C2(n18648), .A(n18067), .B(n18057), .ZN(
        n18008) );
  AOI21_X1 U21006 ( .B1(n18004), .B2(n18059), .A(n18008), .ZN(n17979) );
  OAI211_X1 U21007 ( .C1(n17980), .C2(n18635), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17979), .ZN(n17990) );
  OAI221_X1 U21008 ( .B1(n17981), .B2(n18081), .C1(n17981), .C2(n17990), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17986) );
  AOI22_X1 U21009 ( .A1(n18072), .A2(n17984), .B1(n17983), .B2(n17982), .ZN(
        n17985) );
  OAI221_X1 U21010 ( .B1(n18165), .B2(n17986), .C1(n18122), .C2(n18750), .A(
        n17985), .ZN(P3_U2846) );
  AOI21_X1 U21011 ( .B1(n17987), .B2(n18001), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17988) );
  INV_X1 U21012 ( .A(n17988), .ZN(n17989) );
  AOI22_X1 U21013 ( .A1(n17992), .A2(n17991), .B1(n17990), .B2(n17989), .ZN(
        n17999) );
  AOI22_X1 U21014 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18156), .B1(
        n18165), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n17998) );
  NOR2_X1 U21015 ( .A1(n17993), .A2(n18171), .ZN(n17995) );
  AOI22_X1 U21016 ( .A1(n18072), .A2(n17996), .B1(n17995), .B2(n17994), .ZN(
        n17997) );
  OAI211_X1 U21017 ( .C1(n17999), .C2(n18154), .A(n17998), .B(n17997), .ZN(
        P3_U2847) );
  AOI22_X1 U21018 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18156), .B1(
        n18153), .B2(P3_REIP_REG_14__SCAN_IN), .ZN(n18015) );
  NOR2_X1 U21019 ( .A1(n18003), .A2(n18000), .ZN(n18002) );
  AOI21_X1 U21020 ( .B1(n18002), .B2(n18001), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18011) );
  NOR2_X1 U21021 ( .A1(n18003), .A2(n18065), .ZN(n18035) );
  NOR2_X1 U21022 ( .A1(n18635), .A2(n18035), .ZN(n18029) );
  OAI21_X1 U21023 ( .B1(n18005), .B2(n18059), .A(n18004), .ZN(n18006) );
  OAI21_X1 U21024 ( .B1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n18155), .A(
        n18006), .ZN(n18007) );
  NOR3_X1 U21025 ( .A1(n18029), .A2(n18008), .A3(n18007), .ZN(n18010) );
  OAI22_X1 U21026 ( .A1(n18011), .A2(n18010), .B1(n18045), .B2(n18009), .ZN(
        n18013) );
  AOI22_X1 U21027 ( .A1(n18162), .A2(n18013), .B1(n18072), .B2(n18012), .ZN(
        n18014) );
  OAI211_X1 U21028 ( .C1(n18171), .C2(n18016), .A(n18015), .B(n18014), .ZN(
        P3_U2848) );
  NOR2_X1 U21029 ( .A1(n18036), .A2(n18075), .ZN(n18018) );
  AOI22_X1 U21030 ( .A1(n18165), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18018), 
        .B2(n18017), .ZN(n18031) );
  AOI21_X1 U21031 ( .B1(n18658), .B2(n18019), .A(n18042), .ZN(n18034) );
  NOR2_X1 U21032 ( .A1(n18020), .A2(n18648), .ZN(n18048) );
  AOI21_X1 U21033 ( .B1(n18051), .B2(n18021), .A(n18634), .ZN(n18022) );
  AOI21_X1 U21034 ( .B1(n18654), .B2(n18036), .A(n18022), .ZN(n18052) );
  OAI21_X1 U21035 ( .B1(n18023), .B2(n18626), .A(n18052), .ZN(n18024) );
  AOI211_X1 U21036 ( .C1(n18026), .C2(n18025), .A(n18048), .B(n18024), .ZN(
        n18033) );
  OAI211_X1 U21037 ( .C1(n18027), .C2(n18034), .A(n18162), .B(n18033), .ZN(
        n18028) );
  OAI211_X1 U21038 ( .C1(n18029), .C2(n18028), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18122), .ZN(n18030) );
  OAI211_X1 U21039 ( .C1(n18091), .C2(n18032), .A(n18031), .B(n18030), .ZN(
        P3_U2849) );
  OAI211_X1 U21040 ( .C1(n18035), .C2(n18635), .A(n18034), .B(n18033), .ZN(
        n18038) );
  OAI22_X1 U21041 ( .A1(n18036), .A2(n18075), .B1(n18042), .B2(n18154), .ZN(
        n18037) );
  AOI22_X1 U21042 ( .A1(n18072), .A2(n18039), .B1(n18038), .B2(n18037), .ZN(
        n18041) );
  OAI211_X1 U21043 ( .C1(n18119), .C2(n18042), .A(n18041), .B(n18040), .ZN(
        P3_U2850) );
  AOI22_X1 U21044 ( .A1(n18165), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18072), 
        .B2(n18043), .ZN(n18055) );
  OAI22_X1 U21045 ( .A1(n18046), .A2(n18045), .B1(n18626), .B2(n18044), .ZN(
        n18047) );
  NOR2_X1 U21046 ( .A1(n18048), .A2(n18047), .ZN(n18066) );
  OAI21_X1 U21047 ( .B1(n12781), .B2(n18065), .A(n18633), .ZN(n18049) );
  OAI211_X1 U21048 ( .C1(n18051), .C2(n18050), .A(n18066), .B(n18049), .ZN(
        n18058) );
  OAI211_X1 U21049 ( .C1(n18635), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18052), .B(n18119), .ZN(n18053) );
  OAI211_X1 U21050 ( .C1(n18058), .C2(n18053), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18122), .ZN(n18054) );
  OAI211_X1 U21051 ( .C1(n18056), .C2(n18075), .A(n18055), .B(n18054), .ZN(
        P3_U2851) );
  NAND2_X1 U21052 ( .A1(n18162), .A2(n18057), .ZN(n18070) );
  AOI211_X1 U21053 ( .C1(n12781), .C2(n18059), .A(n18058), .B(n18070), .ZN(
        n18060) );
  AOI21_X1 U21054 ( .B1(n18060), .B2(n18067), .A(n12780), .ZN(n18062) );
  NOR3_X1 U21055 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n12781), .A3(
        n18075), .ZN(n18061) );
  AOI221_X1 U21056 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n18165), .C1(n18062), 
        .C2(n18122), .A(n18061), .ZN(n18063) );
  OAI21_X1 U21057 ( .B1(n18064), .B2(n18091), .A(n18063), .ZN(P3_U2852) );
  INV_X1 U21058 ( .A(n18065), .ZN(n18068) );
  OAI211_X1 U21059 ( .C1(n18068), .C2(n18635), .A(n18067), .B(n18066), .ZN(
        n18069) );
  OAI21_X1 U21060 ( .B1(n18070), .B2(n18069), .A(n18122), .ZN(n18074) );
  AOI22_X1 U21061 ( .A1(n18153), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18072), 
        .B2(n18071), .ZN(n18073) );
  OAI221_X1 U21062 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18075), .C1(
        n12781), .C2(n18074), .A(n18073), .ZN(P3_U2853) );
  NOR3_X1 U21063 ( .A1(n18154), .A2(n18076), .A3(n18101), .ZN(n18085) );
  AOI22_X1 U21064 ( .A1(n18654), .A2(n18079), .B1(n18078), .B2(n18077), .ZN(
        n18080) );
  NAND2_X1 U21065 ( .A1(n18080), .A2(n18137), .ZN(n18102) );
  AOI211_X1 U21066 ( .C1(n18081), .C2(n18095), .A(n18094), .B(n18102), .ZN(
        n18093) );
  OAI21_X1 U21067 ( .B1(n18093), .B2(n18082), .A(n18119), .ZN(n18084) );
  AOI221_X1 U21068 ( .B1(n18085), .B2(n20851), .C1(n18084), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18083), .ZN(n18090) );
  AOI22_X1 U21069 ( .A1(n18088), .A2(n18087), .B1(n18152), .B2(n18086), .ZN(
        n18089) );
  OAI211_X1 U21070 ( .C1(n18092), .C2(n18091), .A(n18090), .B(n18089), .ZN(
        P3_U2854) );
  AOI22_X1 U21071 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18156), .B1(
        n18165), .B2(P3_REIP_REG_7__SCAN_IN), .ZN(n18099) );
  AOI221_X1 U21072 ( .B1(n18095), .B2(n18094), .C1(n18101), .C2(n18094), .A(
        n18093), .ZN(n18097) );
  AOI22_X1 U21073 ( .A1(n18162), .A2(n18097), .B1(n18150), .B2(n18096), .ZN(
        n18098) );
  OAI211_X1 U21074 ( .C1(n18171), .C2(n18100), .A(n18099), .B(n18098), .ZN(
        P3_U2855) );
  OR2_X1 U21075 ( .A1(n18154), .A2(n18101), .ZN(n18108) );
  AOI21_X1 U21076 ( .B1(n18102), .B2(n18162), .A(n18156), .ZN(n18103) );
  INV_X1 U21077 ( .A(n18103), .ZN(n18111) );
  AOI22_X1 U21078 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18111), .B1(
        n18153), .B2(P3_REIP_REG_6__SCAN_IN), .ZN(n18107) );
  AOI22_X1 U21079 ( .A1(n18152), .A2(n18105), .B1(n18150), .B2(n18104), .ZN(
        n18106) );
  OAI211_X1 U21080 ( .C1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n18108), .A(
        n18107), .B(n18106), .ZN(P3_U2856) );
  NAND4_X1 U21081 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n18162), .A4(n18128), .ZN(
        n18114) );
  AOI22_X1 U21082 ( .A1(n18153), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18152), 
        .B2(n18109), .ZN(n18113) );
  AOI22_X1 U21083 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18111), .B1(
        n18150), .B2(n18110), .ZN(n18112) );
  OAI211_X1 U21084 ( .C1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n18114), .A(
        n18113), .B(n18112), .ZN(P3_U2857) );
  NAND2_X1 U21085 ( .A1(n18654), .A2(n18115), .ZN(n18143) );
  OAI211_X1 U21086 ( .C1(n18136), .C2(n18116), .A(n18137), .B(n18143), .ZN(
        n18117) );
  OAI21_X1 U21087 ( .B1(n18118), .B2(n18117), .A(n18162), .ZN(n18133) );
  OAI21_X1 U21088 ( .B1(n18120), .B2(n18133), .A(n18119), .ZN(n18124) );
  OAI22_X1 U21089 ( .A1(n18122), .A2(n18726), .B1(n18171), .B2(n18121), .ZN(
        n18123) );
  AOI21_X1 U21090 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18124), .A(
        n18123), .ZN(n18126) );
  NAND4_X1 U21091 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18162), .A3(
        n10066), .A4(n18128), .ZN(n18125) );
  OAI211_X1 U21092 ( .C1(n18127), .C2(n18169), .A(n18126), .B(n18125), .ZN(
        P3_U2858) );
  NOR2_X1 U21093 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18128), .ZN(
        n18134) );
  AOI22_X1 U21094 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18156), .B1(
        n18153), .B2(P3_REIP_REG_3__SCAN_IN), .ZN(n18132) );
  AOI22_X1 U21095 ( .A1(n18152), .A2(n18130), .B1(n18150), .B2(n18129), .ZN(
        n18131) );
  OAI211_X1 U21096 ( .C1(n18134), .C2(n18133), .A(n18132), .B(n18131), .ZN(
        P3_U2859) );
  AOI211_X1 U21097 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n18137), .A(
        n18136), .B(n18135), .ZN(n18140) );
  NOR3_X1 U21098 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18802), .A3(
        n18138), .ZN(n18139) );
  AOI211_X1 U21099 ( .C1(n18141), .C2(n18623), .A(n18140), .B(n18139), .ZN(
        n18144) );
  NAND4_X1 U21100 ( .A1(n18654), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18142) );
  NAND3_X1 U21101 ( .A1(n18144), .A2(n18143), .A3(n18142), .ZN(n18145) );
  AOI22_X1 U21102 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18156), .B1(
        n18162), .B2(n18145), .ZN(n18147) );
  OAI211_X1 U21103 ( .C1(n18148), .C2(n18171), .A(n18147), .B(n18146), .ZN(
        P3_U2860) );
  AOI22_X1 U21104 ( .A1(n18152), .A2(n18151), .B1(n18150), .B2(n18149), .ZN(
        n18161) );
  NAND2_X1 U21105 ( .A1(n18153), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18160) );
  NOR3_X1 U21106 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18155), .A3(
        n18154), .ZN(n18164) );
  OAI21_X1 U21107 ( .B1(n18156), .B2(n18164), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18159) );
  OAI211_X1 U21108 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18658), .A(
        n18157), .B(n18802), .ZN(n18158) );
  NAND4_X1 U21109 ( .A1(n18161), .A2(n18160), .A3(n18159), .A4(n18158), .ZN(
        P3_U2861) );
  AOI21_X1 U21110 ( .B1(n18634), .B2(n18162), .A(n18818), .ZN(n18163) );
  NOR2_X1 U21111 ( .A1(n18164), .A2(n18163), .ZN(n18167) );
  INV_X1 U21112 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18166) );
  MUX2_X1 U21113 ( .A(n18167), .B(n18166), .S(n18165), .Z(n18168) );
  OAI221_X1 U21114 ( .B1(n18172), .B2(n18171), .C1(n18170), .C2(n18169), .A(
        n18168), .ZN(P3_U2862) );
  AOI21_X1 U21115 ( .B1(n18175), .B2(n18174), .A(n18173), .ZN(n18682) );
  INV_X1 U21116 ( .A(n18682), .ZN(n18177) );
  OAI21_X1 U21117 ( .B1(n18178), .B2(n18838), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18176) );
  OAI221_X1 U21118 ( .B1(n18178), .B2(n18177), .C1(n18178), .C2(n18229), .A(
        n18176), .ZN(P3_U2863) );
  NAND2_X1 U21119 ( .A1(n18670), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18451) );
  INV_X1 U21120 ( .A(n18451), .ZN(n18474) );
  NAND2_X1 U21121 ( .A1(n18665), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18330) );
  INV_X1 U21122 ( .A(n18330), .ZN(n18354) );
  NOR2_X1 U21123 ( .A1(n18474), .A2(n18354), .ZN(n18180) );
  OAI22_X1 U21124 ( .A1(n18181), .A2(n18180), .B1(n18665), .B2(n18179), .ZN(
        P3_U2866) );
  INV_X1 U21125 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18666) );
  NOR2_X1 U21126 ( .A1(n18666), .A2(n18182), .ZN(P3_U2867) );
  NOR2_X1 U21127 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18641) );
  NAND2_X1 U21128 ( .A1(n18670), .A2(n18665), .ZN(n18268) );
  INV_X1 U21129 ( .A(n18268), .ZN(n18269) );
  NAND2_X1 U21130 ( .A1(n18641), .A2(n18269), .ZN(n18282) );
  NOR2_X1 U21131 ( .A1(n18184), .A2(n18183), .ZN(n18224) );
  NAND2_X1 U21132 ( .A1(n18185), .A2(n18224), .ZN(n18481) );
  NAND2_X1 U21133 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18568), .ZN(n18572) );
  INV_X1 U21134 ( .A(n18572), .ZN(n18473) );
  NAND2_X1 U21135 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18529) );
  NOR2_X1 U21136 ( .A1(n18529), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18567) );
  NAND2_X1 U21137 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18567), .ZN(
        n18510) );
  INV_X1 U21138 ( .A(n18510), .ZN(n18610) );
  NOR2_X2 U21139 ( .A1(n18376), .A2(n18186), .ZN(n18564) );
  INV_X1 U21140 ( .A(n18562), .ZN(n18691) );
  NOR2_X1 U21141 ( .A1(n18665), .A2(n18352), .ZN(n18566) );
  NAND2_X1 U21142 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18566), .ZN(
        n18579) );
  NOR2_X1 U21143 ( .A1(n20755), .A2(n18614), .ZN(n18248) );
  NOR2_X1 U21144 ( .A1(n18691), .A2(n18248), .ZN(n18223) );
  AOI22_X1 U21145 ( .A1(n18473), .A2(n18610), .B1(n18564), .B2(n18223), .ZN(
        n18192) );
  INV_X1 U21146 ( .A(n18529), .ZN(n18190) );
  NAND2_X1 U21147 ( .A1(n18638), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18399) );
  INV_X1 U21148 ( .A(n18399), .ZN(n18187) );
  NOR2_X1 U21149 ( .A1(n18638), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18331) );
  NOR2_X1 U21150 ( .A1(n18187), .A2(n18331), .ZN(n18477) );
  INV_X1 U21151 ( .A(n18477), .ZN(n18329) );
  NAND2_X1 U21152 ( .A1(n18190), .A2(n18329), .ZN(n18531) );
  OAI21_X1 U21153 ( .B1(n18532), .B2(n18531), .A(n18248), .ZN(n18188) );
  OAI211_X1 U21154 ( .C1(n20755), .C2(n18794), .A(n18535), .B(n18188), .ZN(
        n18226) );
  INV_X1 U21155 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18189) );
  NOR2_X2 U21156 ( .A1(n18285), .A2(n18189), .ZN(n18563) );
  NAND2_X1 U21157 ( .A1(n18331), .A2(n18190), .ZN(n18540) );
  AOI22_X1 U21158 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18226), .B1(
        n18563), .B2(n18557), .ZN(n18191) );
  OAI211_X1 U21159 ( .C1(n18282), .C2(n18481), .A(n18192), .B(n18191), .ZN(
        P3_U2868) );
  NAND2_X1 U21160 ( .A1(n18193), .A2(n18224), .ZN(n18580) );
  NOR2_X2 U21161 ( .A1(n18376), .A2(n18195), .ZN(n18573) );
  AOI22_X1 U21162 ( .A1(n18575), .A2(n18610), .B1(n18573), .B2(n18223), .ZN(
        n18198) );
  INV_X1 U21163 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n18196) );
  NOR2_X2 U21164 ( .A1(n18285), .A2(n18196), .ZN(n18576) );
  AOI22_X1 U21165 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18226), .B1(
        n18576), .B2(n18557), .ZN(n18197) );
  OAI211_X1 U21166 ( .C1(n18282), .C2(n18580), .A(n18198), .B(n18197), .ZN(
        P3_U2869) );
  NAND2_X1 U21167 ( .A1(n18568), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18514) );
  NOR2_X2 U21168 ( .A1(n18376), .A2(n18199), .ZN(n18582) );
  AOI22_X1 U21169 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18226), .B1(
        n18582), .B2(n18223), .ZN(n18203) );
  NAND2_X1 U21170 ( .A1(n18200), .A2(n18224), .ZN(n18409) );
  INV_X1 U21171 ( .A(n18409), .ZN(n18583) );
  INV_X1 U21172 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18201) );
  NOR2_X1 U21173 ( .A1(n18201), .A2(n18285), .ZN(n18511) );
  AOI22_X1 U21174 ( .A1(n20755), .A2(n18583), .B1(n18511), .B2(n18610), .ZN(
        n18202) );
  OAI211_X1 U21175 ( .C1(n18514), .C2(n18540), .A(n18203), .B(n18202), .ZN(
        P3_U2870) );
  NAND2_X1 U21176 ( .A1(n18568), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18546) );
  NOR2_X2 U21177 ( .A1(n18376), .A2(n20912), .ZN(n18587) );
  AOI22_X1 U21178 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18226), .B1(
        n18587), .B2(n18223), .ZN(n18206) );
  NAND2_X1 U21179 ( .A1(n18204), .A2(n18224), .ZN(n18412) );
  INV_X1 U21180 ( .A(n18412), .ZN(n18589) );
  NAND2_X1 U21181 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18568), .ZN(n18592) );
  INV_X1 U21182 ( .A(n18592), .ZN(n18543) );
  AOI22_X1 U21183 ( .A1(n20755), .A2(n18589), .B1(n18543), .B2(n18610), .ZN(
        n18205) );
  OAI211_X1 U21184 ( .C1(n18546), .C2(n18540), .A(n18206), .B(n18205), .ZN(
        P3_U2871) );
  NAND2_X1 U21185 ( .A1(n18207), .A2(n18224), .ZN(n18492) );
  NOR2_X2 U21186 ( .A1(n18376), .A2(n18208), .ZN(n18594) );
  AOI22_X1 U21187 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18226), .B1(
        n18594), .B2(n18223), .ZN(n18211) );
  NOR2_X1 U21188 ( .A1(n18209), .A2(n18285), .ZN(n18489) );
  AND2_X1 U21189 ( .A1(n18568), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18593) );
  AOI22_X1 U21190 ( .A1(n18489), .A2(n18610), .B1(n18593), .B2(n18557), .ZN(
        n18210) );
  OAI211_X1 U21191 ( .C1(n18282), .C2(n18492), .A(n18211), .B(n18210), .ZN(
        P3_U2872) );
  NOR2_X1 U21192 ( .A1(n18212), .A2(n18285), .ZN(n18599) );
  NOR2_X2 U21193 ( .A1(n18213), .A2(n18376), .ZN(n20757) );
  NOR2_X2 U21194 ( .A1(n18214), .A2(n18285), .ZN(n20756) );
  AOI22_X1 U21195 ( .A1(n20757), .A2(n18223), .B1(n20756), .B2(n18610), .ZN(
        n18217) );
  NAND2_X1 U21196 ( .A1(n18224), .A2(n18215), .ZN(n20760) );
  INV_X1 U21197 ( .A(n20760), .ZN(n18600) );
  AOI22_X1 U21198 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18226), .B1(
        n18600), .B2(n20755), .ZN(n18216) );
  OAI211_X1 U21199 ( .C1(n20762), .C2(n18540), .A(n18217), .B(n18216), .ZN(
        P3_U2873) );
  NOR2_X2 U21200 ( .A1(n20902), .A2(n18285), .ZN(n18605) );
  INV_X1 U21201 ( .A(n18605), .ZN(n18498) );
  NOR2_X2 U21202 ( .A1(n18218), .A2(n18376), .ZN(n18604) );
  AOI22_X1 U21203 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18226), .B1(
        n18604), .B2(n18223), .ZN(n18221) );
  NAND2_X1 U21204 ( .A1(n18219), .A2(n18224), .ZN(n18420) );
  INV_X1 U21205 ( .A(n18420), .ZN(n18606) );
  NAND2_X1 U21206 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18568), .ZN(n18609) );
  INV_X1 U21207 ( .A(n18609), .ZN(n18495) );
  AOI22_X1 U21208 ( .A1(n20755), .A2(n18606), .B1(n18495), .B2(n18610), .ZN(
        n18220) );
  OAI211_X1 U21209 ( .C1(n18498), .C2(n18540), .A(n18221), .B(n18220), .ZN(
        P3_U2874) );
  NOR2_X1 U21210 ( .A1(n18285), .A2(n19163), .ZN(n18556) );
  INV_X1 U21211 ( .A(n18556), .ZN(n18620) );
  NOR2_X2 U21212 ( .A1(n18222), .A2(n18376), .ZN(n18613) );
  NAND2_X1 U21213 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18568), .ZN(n18561) );
  INV_X1 U21214 ( .A(n18561), .ZN(n18611) );
  AOI22_X1 U21215 ( .A1(n18613), .A2(n18223), .B1(n18611), .B2(n18557), .ZN(
        n18228) );
  AND2_X1 U21216 ( .A1(n18225), .A2(n18224), .ZN(n18615) );
  AOI22_X1 U21217 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18226), .B1(
        n20755), .B2(n18615), .ZN(n18227) );
  OAI211_X1 U21218 ( .C1(n18620), .C2(n18510), .A(n18228), .B(n18227), .ZN(
        P3_U2875) );
  NOR2_X1 U21219 ( .A1(n18268), .A2(n18399), .ZN(n18300) );
  INV_X1 U21220 ( .A(n18300), .ZN(n20763) );
  NAND2_X1 U21221 ( .A1(n18638), .A2(n18562), .ZN(n18400) );
  NOR2_X1 U21222 ( .A1(n18268), .A2(n18400), .ZN(n18244) );
  AOI22_X1 U21223 ( .A1(n18473), .A2(n18557), .B1(n18564), .B2(n18244), .ZN(
        n18231) );
  NAND2_X1 U21224 ( .A1(n18535), .A2(n18229), .ZN(n18401) );
  NOR2_X1 U21225 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18401), .ZN(
        n18307) );
  AOI22_X1 U21226 ( .A1(n18568), .A2(n18566), .B1(n18269), .B2(n18307), .ZN(
        n18245) );
  AOI22_X1 U21227 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18245), .B1(
        n18563), .B2(n18614), .ZN(n18230) );
  OAI211_X1 U21228 ( .C1(n20763), .C2(n18481), .A(n18231), .B(n18230), .ZN(
        P3_U2876) );
  AOI22_X1 U21229 ( .A1(n18576), .A2(n18614), .B1(n18573), .B2(n18244), .ZN(
        n18233) );
  AOI22_X1 U21230 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18245), .B1(
        n18575), .B2(n18557), .ZN(n18232) );
  OAI211_X1 U21231 ( .C1(n20763), .C2(n18580), .A(n18233), .B(n18232), .ZN(
        P3_U2877) );
  AOI22_X1 U21232 ( .A1(n18511), .A2(n18557), .B1(n18582), .B2(n18244), .ZN(
        n18235) );
  INV_X1 U21233 ( .A(n18514), .ZN(n18581) );
  AOI22_X1 U21234 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18245), .B1(
        n18581), .B2(n18614), .ZN(n18234) );
  OAI211_X1 U21235 ( .C1(n20763), .C2(n18409), .A(n18235), .B(n18234), .ZN(
        P3_U2878) );
  AOI22_X1 U21236 ( .A1(n18587), .A2(n18244), .B1(n18543), .B2(n18557), .ZN(
        n18237) );
  INV_X1 U21237 ( .A(n18546), .ZN(n18588) );
  AOI22_X1 U21238 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18245), .B1(
        n18588), .B2(n18614), .ZN(n18236) );
  OAI211_X1 U21239 ( .C1(n20763), .C2(n18412), .A(n18237), .B(n18236), .ZN(
        P3_U2879) );
  AOI22_X1 U21240 ( .A1(n18594), .A2(n18244), .B1(n18593), .B2(n18614), .ZN(
        n18239) );
  AOI22_X1 U21241 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18245), .B1(
        n18489), .B2(n18557), .ZN(n18238) );
  OAI211_X1 U21242 ( .C1(n20763), .C2(n18492), .A(n18239), .B(n18238), .ZN(
        P3_U2880) );
  AOI22_X1 U21243 ( .A1(n18599), .A2(n18614), .B1(n20757), .B2(n18244), .ZN(
        n18241) );
  AOI22_X1 U21244 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18245), .B1(
        n20756), .B2(n18557), .ZN(n18240) );
  OAI211_X1 U21245 ( .C1(n20763), .C2(n20760), .A(n18241), .B(n18240), .ZN(
        P3_U2881) );
  AOI22_X1 U21246 ( .A1(n18604), .A2(n18244), .B1(n18495), .B2(n18557), .ZN(
        n18243) );
  AOI22_X1 U21247 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18245), .B1(
        n18605), .B2(n18614), .ZN(n18242) );
  OAI211_X1 U21248 ( .C1(n20763), .C2(n18420), .A(n18243), .B(n18242), .ZN(
        P3_U2882) );
  AOI22_X1 U21249 ( .A1(n18613), .A2(n18244), .B1(n18611), .B2(n18614), .ZN(
        n18247) );
  AOI22_X1 U21250 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18245), .B1(
        n18300), .B2(n18615), .ZN(n18246) );
  OAI211_X1 U21251 ( .C1(n18620), .C2(n18540), .A(n18247), .B(n18246), .ZN(
        P3_U2883) );
  INV_X1 U21252 ( .A(n18331), .ZN(n18426) );
  NOR2_X2 U21253 ( .A1(n18268), .A2(n18426), .ZN(n18319) );
  INV_X1 U21254 ( .A(n18319), .ZN(n18328) );
  NOR2_X1 U21255 ( .A1(n18300), .A2(n18319), .ZN(n18286) );
  NOR2_X1 U21256 ( .A1(n18691), .A2(n18286), .ZN(n18264) );
  AOI22_X1 U21257 ( .A1(n20755), .A2(n18563), .B1(n18564), .B2(n18264), .ZN(
        n18251) );
  OAI21_X1 U21258 ( .B1(n18248), .B2(n18532), .A(n18286), .ZN(n18249) );
  OAI211_X1 U21259 ( .C1(n18319), .C2(n18794), .A(n18535), .B(n18249), .ZN(
        n18265) );
  AOI22_X1 U21260 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18265), .B1(
        n18473), .B2(n18614), .ZN(n18250) );
  OAI211_X1 U21261 ( .C1(n18481), .C2(n18328), .A(n18251), .B(n18250), .ZN(
        P3_U2884) );
  AOI22_X1 U21262 ( .A1(n18575), .A2(n18614), .B1(n18573), .B2(n18264), .ZN(
        n18253) );
  AOI22_X1 U21263 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18265), .B1(
        n20755), .B2(n18576), .ZN(n18252) );
  OAI211_X1 U21264 ( .C1(n18580), .C2(n18328), .A(n18253), .B(n18252), .ZN(
        P3_U2885) );
  AOI22_X1 U21265 ( .A1(n18511), .A2(n18614), .B1(n18582), .B2(n18264), .ZN(
        n18255) );
  AOI22_X1 U21266 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18265), .B1(
        n18583), .B2(n18319), .ZN(n18254) );
  OAI211_X1 U21267 ( .C1(n18282), .C2(n18514), .A(n18255), .B(n18254), .ZN(
        P3_U2886) );
  AOI22_X1 U21268 ( .A1(n18587), .A2(n18264), .B1(n18543), .B2(n18614), .ZN(
        n18257) );
  AOI22_X1 U21269 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18265), .B1(
        n18589), .B2(n18319), .ZN(n18256) );
  OAI211_X1 U21270 ( .C1(n18282), .C2(n18546), .A(n18257), .B(n18256), .ZN(
        P3_U2887) );
  AOI22_X1 U21271 ( .A1(n20755), .A2(n18593), .B1(n18594), .B2(n18264), .ZN(
        n18259) );
  AOI22_X1 U21272 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18265), .B1(
        n18489), .B2(n18614), .ZN(n18258) );
  OAI211_X1 U21273 ( .C1(n18492), .C2(n18328), .A(n18259), .B(n18258), .ZN(
        P3_U2888) );
  AOI22_X1 U21274 ( .A1(n18599), .A2(n20755), .B1(n20757), .B2(n18264), .ZN(
        n18261) );
  AOI22_X1 U21275 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18265), .B1(
        n20756), .B2(n18614), .ZN(n18260) );
  OAI211_X1 U21276 ( .C1(n20760), .C2(n18328), .A(n18261), .B(n18260), .ZN(
        P3_U2889) );
  AOI22_X1 U21277 ( .A1(n20755), .A2(n18605), .B1(n18604), .B2(n18264), .ZN(
        n18263) );
  AOI22_X1 U21278 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18265), .B1(
        n18495), .B2(n18614), .ZN(n18262) );
  OAI211_X1 U21279 ( .C1(n18420), .C2(n18328), .A(n18263), .B(n18262), .ZN(
        P3_U2890) );
  AOI22_X1 U21280 ( .A1(n18556), .A2(n18614), .B1(n18613), .B2(n18264), .ZN(
        n18267) );
  AOI22_X1 U21281 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18265), .B1(
        n18615), .B2(n18319), .ZN(n18266) );
  OAI211_X1 U21282 ( .C1(n18282), .C2(n18561), .A(n18267), .B(n18266), .ZN(
        P3_U2891) );
  NOR2_X1 U21283 ( .A1(n18638), .A2(n18268), .ZN(n18308) );
  AND2_X1 U21284 ( .A1(n18308), .A2(n18562), .ZN(n20758) );
  AOI22_X1 U21285 ( .A1(n18300), .A2(n18563), .B1(n20758), .B2(n18564), .ZN(
        n18271) );
  NAND2_X1 U21286 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18308), .ZN(
        n20761) );
  OAI21_X1 U21287 ( .B1(n18376), .B2(n18638), .A(n18285), .ZN(n18353) );
  OAI211_X1 U21288 ( .C1(n18346), .C2(n18794), .A(n18269), .B(n18353), .ZN(
        n20766) );
  INV_X1 U21289 ( .A(n18481), .ZN(n18569) );
  AOI22_X1 U21290 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20766), .B1(
        n18346), .B2(n18569), .ZN(n18270) );
  OAI211_X1 U21291 ( .C1(n18282), .C2(n18572), .A(n18271), .B(n18270), .ZN(
        P3_U2892) );
  INV_X1 U21292 ( .A(n18575), .ZN(n18434) );
  AOI22_X1 U21293 ( .A1(n18300), .A2(n18576), .B1(n20758), .B2(n18573), .ZN(
        n18273) );
  INV_X1 U21294 ( .A(n18580), .ZN(n18431) );
  AOI22_X1 U21295 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20766), .B1(
        n18346), .B2(n18431), .ZN(n18272) );
  OAI211_X1 U21296 ( .C1(n18282), .C2(n18434), .A(n18273), .B(n18272), .ZN(
        P3_U2893) );
  AOI22_X1 U21297 ( .A1(n20758), .A2(n18582), .B1(n20755), .B2(n18511), .ZN(
        n18275) );
  AOI22_X1 U21298 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20766), .B1(
        n18346), .B2(n18583), .ZN(n18274) );
  OAI211_X1 U21299 ( .C1(n20763), .C2(n18514), .A(n18275), .B(n18274), .ZN(
        P3_U2894) );
  AOI22_X1 U21300 ( .A1(n18300), .A2(n18588), .B1(n20758), .B2(n18587), .ZN(
        n18277) );
  AOI22_X1 U21301 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20766), .B1(
        n18346), .B2(n18589), .ZN(n18276) );
  OAI211_X1 U21302 ( .C1(n18282), .C2(n18592), .A(n18277), .B(n18276), .ZN(
        P3_U2895) );
  INV_X1 U21303 ( .A(n18489), .ZN(n18598) );
  AOI22_X1 U21304 ( .A1(n18300), .A2(n18593), .B1(n20758), .B2(n18594), .ZN(
        n18279) );
  INV_X1 U21305 ( .A(n18492), .ZN(n18595) );
  AOI22_X1 U21306 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20766), .B1(
        n18346), .B2(n18595), .ZN(n18278) );
  OAI211_X1 U21307 ( .C1(n18282), .C2(n18598), .A(n18279), .B(n18278), .ZN(
        P3_U2896) );
  AOI22_X1 U21308 ( .A1(n18300), .A2(n18605), .B1(n20758), .B2(n18604), .ZN(
        n18281) );
  AOI22_X1 U21309 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20766), .B1(
        n18346), .B2(n18606), .ZN(n18280) );
  OAI211_X1 U21310 ( .C1(n18282), .C2(n18609), .A(n18281), .B(n18280), .ZN(
        P3_U2898) );
  AOI22_X1 U21311 ( .A1(n20758), .A2(n18613), .B1(n20755), .B2(n18556), .ZN(
        n18284) );
  AOI22_X1 U21312 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20766), .B1(
        n18346), .B2(n18615), .ZN(n18283) );
  OAI211_X1 U21313 ( .C1(n20763), .C2(n18561), .A(n18284), .B(n18283), .ZN(
        P3_U2899) );
  NAND2_X1 U21314 ( .A1(n18641), .A2(n18354), .ZN(n18369) );
  NOR2_X1 U21315 ( .A1(n18346), .A2(n18371), .ZN(n18332) );
  NOR2_X1 U21316 ( .A1(n18691), .A2(n18332), .ZN(n18303) );
  AOI22_X1 U21317 ( .A1(n18564), .A2(n18303), .B1(n18563), .B2(n18319), .ZN(
        n18289) );
  OAI22_X1 U21318 ( .A1(n18332), .A2(n18376), .B1(n18286), .B2(n18285), .ZN(
        n18287) );
  OAI21_X1 U21319 ( .B1(n18371), .B2(n18794), .A(n18287), .ZN(n18304) );
  AOI22_X1 U21320 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18304), .B1(
        n18371), .B2(n18569), .ZN(n18288) );
  OAI211_X1 U21321 ( .C1(n20763), .C2(n18572), .A(n18289), .B(n18288), .ZN(
        P3_U2900) );
  AOI22_X1 U21322 ( .A1(n18576), .A2(n18319), .B1(n18573), .B2(n18303), .ZN(
        n18291) );
  AOI22_X1 U21323 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18304), .B1(
        n18371), .B2(n18431), .ZN(n18290) );
  OAI211_X1 U21324 ( .C1(n20763), .C2(n18434), .A(n18291), .B(n18290), .ZN(
        P3_U2901) );
  INV_X1 U21325 ( .A(n18511), .ZN(n18586) );
  AOI22_X1 U21326 ( .A1(n18582), .A2(n18303), .B1(n18581), .B2(n18319), .ZN(
        n18293) );
  AOI22_X1 U21327 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18304), .B1(
        n18371), .B2(n18583), .ZN(n18292) );
  OAI211_X1 U21328 ( .C1(n20763), .C2(n18586), .A(n18293), .B(n18292), .ZN(
        P3_U2902) );
  AOI22_X1 U21329 ( .A1(n18300), .A2(n18543), .B1(n18587), .B2(n18303), .ZN(
        n18295) );
  AOI22_X1 U21330 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18304), .B1(
        n18371), .B2(n18589), .ZN(n18294) );
  OAI211_X1 U21331 ( .C1(n18546), .C2(n18328), .A(n18295), .B(n18294), .ZN(
        P3_U2903) );
  AOI22_X1 U21332 ( .A1(n18300), .A2(n18489), .B1(n18594), .B2(n18303), .ZN(
        n18297) );
  AOI22_X1 U21333 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18304), .B1(
        n18593), .B2(n18319), .ZN(n18296) );
  OAI211_X1 U21334 ( .C1(n18369), .C2(n18492), .A(n18297), .B(n18296), .ZN(
        P3_U2904) );
  INV_X1 U21335 ( .A(n20756), .ZN(n18603) );
  AOI22_X1 U21336 ( .A1(n18599), .A2(n18319), .B1(n20757), .B2(n18303), .ZN(
        n18299) );
  AOI22_X1 U21337 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18304), .B1(
        n18600), .B2(n18371), .ZN(n18298) );
  OAI211_X1 U21338 ( .C1(n20763), .C2(n18603), .A(n18299), .B(n18298), .ZN(
        P3_U2905) );
  AOI22_X1 U21339 ( .A1(n18300), .A2(n18495), .B1(n18604), .B2(n18303), .ZN(
        n18302) );
  AOI22_X1 U21340 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18304), .B1(
        n18371), .B2(n18606), .ZN(n18301) );
  OAI211_X1 U21341 ( .C1(n18498), .C2(n18328), .A(n18302), .B(n18301), .ZN(
        P3_U2906) );
  AOI22_X1 U21342 ( .A1(n18613), .A2(n18303), .B1(n18611), .B2(n18319), .ZN(
        n18306) );
  AOI22_X1 U21343 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18304), .B1(
        n18371), .B2(n18615), .ZN(n18305) );
  OAI211_X1 U21344 ( .C1(n20763), .C2(n18620), .A(n18306), .B(n18305), .ZN(
        P3_U2907) );
  NOR2_X1 U21345 ( .A1(n18330), .A2(n18400), .ZN(n18324) );
  AOI22_X1 U21346 ( .A1(n18346), .A2(n18563), .B1(n18564), .B2(n18324), .ZN(
        n18310) );
  AOI22_X1 U21347 ( .A1(n18568), .A2(n18308), .B1(n18354), .B2(n18307), .ZN(
        n18325) );
  NOR2_X2 U21348 ( .A1(n18330), .A2(n18399), .ZN(n18395) );
  AOI22_X1 U21349 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18325), .B1(
        n18395), .B2(n18569), .ZN(n18309) );
  OAI211_X1 U21350 ( .C1(n18572), .C2(n18328), .A(n18310), .B(n18309), .ZN(
        P3_U2908) );
  INV_X1 U21351 ( .A(n18395), .ZN(n18393) );
  AOI22_X1 U21352 ( .A1(n18575), .A2(n18319), .B1(n18573), .B2(n18324), .ZN(
        n18312) );
  AOI22_X1 U21353 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18325), .B1(
        n18346), .B2(n18576), .ZN(n18311) );
  OAI211_X1 U21354 ( .C1(n18393), .C2(n18580), .A(n18312), .B(n18311), .ZN(
        P3_U2909) );
  AOI22_X1 U21355 ( .A1(n18346), .A2(n18581), .B1(n18582), .B2(n18324), .ZN(
        n18314) );
  AOI22_X1 U21356 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18325), .B1(
        n18395), .B2(n18583), .ZN(n18313) );
  OAI211_X1 U21357 ( .C1(n18586), .C2(n18328), .A(n18314), .B(n18313), .ZN(
        P3_U2910) );
  AOI22_X1 U21358 ( .A1(n18346), .A2(n18588), .B1(n18587), .B2(n18324), .ZN(
        n18316) );
  AOI22_X1 U21359 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18325), .B1(
        n18395), .B2(n18589), .ZN(n18315) );
  OAI211_X1 U21360 ( .C1(n18592), .C2(n18328), .A(n18316), .B(n18315), .ZN(
        P3_U2911) );
  AOI22_X1 U21361 ( .A1(n18346), .A2(n18593), .B1(n18594), .B2(n18324), .ZN(
        n18318) );
  AOI22_X1 U21362 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18325), .B1(
        n18395), .B2(n18595), .ZN(n18317) );
  OAI211_X1 U21363 ( .C1(n18598), .C2(n18328), .A(n18318), .B(n18317), .ZN(
        P3_U2912) );
  AOI22_X1 U21364 ( .A1(n20757), .A2(n18324), .B1(n20756), .B2(n18319), .ZN(
        n18321) );
  AOI22_X1 U21365 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18325), .B1(
        n18600), .B2(n18395), .ZN(n18320) );
  OAI211_X1 U21366 ( .C1(n20762), .C2(n20761), .A(n18321), .B(n18320), .ZN(
        P3_U2913) );
  AOI22_X1 U21367 ( .A1(n18346), .A2(n18605), .B1(n18604), .B2(n18324), .ZN(
        n18323) );
  AOI22_X1 U21368 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18325), .B1(
        n18395), .B2(n18606), .ZN(n18322) );
  OAI211_X1 U21369 ( .C1(n18609), .C2(n18328), .A(n18323), .B(n18322), .ZN(
        P3_U2914) );
  AOI22_X1 U21370 ( .A1(n18346), .A2(n18611), .B1(n18613), .B2(n18324), .ZN(
        n18327) );
  AOI22_X1 U21371 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18325), .B1(
        n18395), .B2(n18615), .ZN(n18326) );
  OAI211_X1 U21372 ( .C1(n18620), .C2(n18328), .A(n18327), .B(n18326), .ZN(
        P3_U2915) );
  NAND2_X1 U21373 ( .A1(n18562), .A2(n18329), .ZN(n18530) );
  NOR2_X1 U21374 ( .A1(n18330), .A2(n18530), .ZN(n18375) );
  AOI22_X1 U21375 ( .A1(n18371), .A2(n18563), .B1(n18564), .B2(n18375), .ZN(
        n18335) );
  NAND2_X1 U21376 ( .A1(n18354), .A2(n18331), .ZN(n18425) );
  INV_X1 U21377 ( .A(n18425), .ZN(n18417) );
  AOI221_X1 U21378 ( .B1(n18332), .B2(n18393), .C1(n18532), .C2(n18393), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18333) );
  OAI21_X1 U21379 ( .B1(n18417), .B2(n18333), .A(n18535), .ZN(n18349) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18349), .B1(
        n18417), .B2(n18569), .ZN(n18334) );
  OAI211_X1 U21381 ( .C1(n20761), .C2(n18572), .A(n18335), .B(n18334), .ZN(
        P3_U2916) );
  AOI22_X1 U21382 ( .A1(n18371), .A2(n18576), .B1(n18375), .B2(n18573), .ZN(
        n18337) );
  AOI22_X1 U21383 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18349), .B1(
        n18417), .B2(n18431), .ZN(n18336) );
  OAI211_X1 U21384 ( .C1(n20761), .C2(n18434), .A(n18337), .B(n18336), .ZN(
        P3_U2917) );
  AOI22_X1 U21385 ( .A1(n18371), .A2(n18581), .B1(n18375), .B2(n18582), .ZN(
        n18339) );
  AOI22_X1 U21386 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18349), .B1(
        n18417), .B2(n18583), .ZN(n18338) );
  OAI211_X1 U21387 ( .C1(n20761), .C2(n18586), .A(n18339), .B(n18338), .ZN(
        P3_U2918) );
  AOI22_X1 U21388 ( .A1(n18346), .A2(n18543), .B1(n18375), .B2(n18587), .ZN(
        n18341) );
  AOI22_X1 U21389 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18349), .B1(
        n18417), .B2(n18589), .ZN(n18340) );
  OAI211_X1 U21390 ( .C1(n18369), .C2(n18546), .A(n18341), .B(n18340), .ZN(
        P3_U2919) );
  AOI22_X1 U21391 ( .A1(n18371), .A2(n18593), .B1(n18375), .B2(n18594), .ZN(
        n18343) );
  AOI22_X1 U21392 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18349), .B1(
        n18417), .B2(n18595), .ZN(n18342) );
  OAI211_X1 U21393 ( .C1(n20761), .C2(n18598), .A(n18343), .B(n18342), .ZN(
        P3_U2920) );
  AOI22_X1 U21394 ( .A1(n18346), .A2(n20756), .B1(n20757), .B2(n18375), .ZN(
        n18345) );
  AOI22_X1 U21395 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18349), .B1(
        n18600), .B2(n18417), .ZN(n18344) );
  OAI211_X1 U21396 ( .C1(n20762), .C2(n18369), .A(n18345), .B(n18344), .ZN(
        P3_U2921) );
  AOI22_X1 U21397 ( .A1(n18346), .A2(n18495), .B1(n18375), .B2(n18604), .ZN(
        n18348) );
  AOI22_X1 U21398 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18349), .B1(
        n18417), .B2(n18606), .ZN(n18347) );
  OAI211_X1 U21399 ( .C1(n18369), .C2(n18498), .A(n18348), .B(n18347), .ZN(
        P3_U2922) );
  AOI22_X1 U21400 ( .A1(n18371), .A2(n18611), .B1(n18375), .B2(n18613), .ZN(
        n18351) );
  AOI22_X1 U21401 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18349), .B1(
        n18417), .B2(n18615), .ZN(n18350) );
  OAI211_X1 U21402 ( .C1(n20761), .C2(n18620), .A(n18351), .B(n18350), .ZN(
        P3_U2923) );
  NOR2_X1 U21403 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18352), .ZN(
        n18402) );
  AND2_X1 U21404 ( .A1(n18562), .A2(n18402), .ZN(n18370) );
  AOI22_X1 U21405 ( .A1(n18395), .A2(n18563), .B1(n18564), .B2(n18370), .ZN(
        n18356) );
  NAND2_X1 U21406 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18402), .ZN(
        n18445) );
  OAI211_X1 U21407 ( .C1(n18447), .C2(n18794), .A(n18354), .B(n18353), .ZN(
        n18372) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18372), .B1(
        n18569), .B2(n18447), .ZN(n18355) );
  OAI211_X1 U21409 ( .C1(n18369), .C2(n18572), .A(n18356), .B(n18355), .ZN(
        P3_U2924) );
  AOI22_X1 U21410 ( .A1(n18371), .A2(n18575), .B1(n18573), .B2(n18370), .ZN(
        n18358) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18372), .B1(
        n18395), .B2(n18576), .ZN(n18357) );
  OAI211_X1 U21412 ( .C1(n18580), .C2(n18445), .A(n18358), .B(n18357), .ZN(
        P3_U2925) );
  AOI22_X1 U21413 ( .A1(n18371), .A2(n18511), .B1(n18582), .B2(n18370), .ZN(
        n18360) );
  AOI22_X1 U21414 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18372), .B1(
        n18583), .B2(n18447), .ZN(n18359) );
  OAI211_X1 U21415 ( .C1(n18393), .C2(n18514), .A(n18360), .B(n18359), .ZN(
        P3_U2926) );
  AOI22_X1 U21416 ( .A1(n18395), .A2(n18588), .B1(n18587), .B2(n18370), .ZN(
        n18362) );
  AOI22_X1 U21417 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18372), .B1(
        n18589), .B2(n18447), .ZN(n18361) );
  OAI211_X1 U21418 ( .C1(n18369), .C2(n18592), .A(n18362), .B(n18361), .ZN(
        P3_U2927) );
  AOI22_X1 U21419 ( .A1(n18371), .A2(n18489), .B1(n18594), .B2(n18370), .ZN(
        n18364) );
  AOI22_X1 U21420 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18372), .B1(
        n18395), .B2(n18593), .ZN(n18363) );
  OAI211_X1 U21421 ( .C1(n18492), .C2(n18445), .A(n18364), .B(n18363), .ZN(
        P3_U2928) );
  AOI22_X1 U21422 ( .A1(n18599), .A2(n18395), .B1(n20757), .B2(n18370), .ZN(
        n18366) );
  AOI22_X1 U21423 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18372), .B1(
        n18600), .B2(n18447), .ZN(n18365) );
  OAI211_X1 U21424 ( .C1(n18603), .C2(n18369), .A(n18366), .B(n18365), .ZN(
        P3_U2929) );
  AOI22_X1 U21425 ( .A1(n18395), .A2(n18605), .B1(n18604), .B2(n18370), .ZN(
        n18368) );
  AOI22_X1 U21426 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18372), .B1(
        n18606), .B2(n18447), .ZN(n18367) );
  OAI211_X1 U21427 ( .C1(n18369), .C2(n18609), .A(n18368), .B(n18367), .ZN(
        P3_U2930) );
  AOI22_X1 U21428 ( .A1(n18371), .A2(n18556), .B1(n18613), .B2(n18370), .ZN(
        n18374) );
  AOI22_X1 U21429 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18372), .B1(
        n18615), .B2(n18447), .ZN(n18373) );
  OAI211_X1 U21430 ( .C1(n18393), .C2(n18561), .A(n18374), .B(n18373), .ZN(
        P3_U2931) );
  NAND2_X1 U21431 ( .A1(n18641), .A2(n18474), .ZN(n18467) );
  AOI21_X1 U21432 ( .B1(n18467), .B2(n18445), .A(n18691), .ZN(n18394) );
  AOI22_X1 U21433 ( .A1(n18395), .A2(n18473), .B1(n18564), .B2(n18394), .ZN(
        n18380) );
  OAI221_X1 U21434 ( .B1(n18475), .B2(n18447), .C1(n18375), .C2(n18447), .A(
        n18794), .ZN(n18377) );
  AOI21_X1 U21435 ( .B1(n18467), .B2(n18377), .A(n18376), .ZN(n18378) );
  INV_X1 U21436 ( .A(n18378), .ZN(n18396) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18396), .B1(
        n18417), .B2(n18563), .ZN(n18379) );
  OAI211_X1 U21438 ( .C1(n18481), .C2(n18467), .A(n18380), .B(n18379), .ZN(
        P3_U2932) );
  AOI22_X1 U21439 ( .A1(n18417), .A2(n18576), .B1(n18573), .B2(n18394), .ZN(
        n18382) );
  INV_X1 U21440 ( .A(n18467), .ZN(n18469) );
  AOI22_X1 U21441 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18396), .B1(
        n18431), .B2(n18469), .ZN(n18381) );
  OAI211_X1 U21442 ( .C1(n18393), .C2(n18434), .A(n18382), .B(n18381), .ZN(
        P3_U2933) );
  AOI22_X1 U21443 ( .A1(n18417), .A2(n18581), .B1(n18582), .B2(n18394), .ZN(
        n18384) );
  AOI22_X1 U21444 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18396), .B1(
        n18583), .B2(n18469), .ZN(n18383) );
  OAI211_X1 U21445 ( .C1(n18393), .C2(n18586), .A(n18384), .B(n18383), .ZN(
        P3_U2934) );
  AOI22_X1 U21446 ( .A1(n18417), .A2(n18588), .B1(n18587), .B2(n18394), .ZN(
        n18386) );
  AOI22_X1 U21447 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18396), .B1(
        n18589), .B2(n18469), .ZN(n18385) );
  OAI211_X1 U21448 ( .C1(n18393), .C2(n18592), .A(n18386), .B(n18385), .ZN(
        P3_U2935) );
  AOI22_X1 U21449 ( .A1(n18395), .A2(n18489), .B1(n18594), .B2(n18394), .ZN(
        n18388) );
  AOI22_X1 U21450 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18396), .B1(
        n18417), .B2(n18593), .ZN(n18387) );
  OAI211_X1 U21451 ( .C1(n18492), .C2(n18467), .A(n18388), .B(n18387), .ZN(
        P3_U2936) );
  AOI22_X1 U21452 ( .A1(n20757), .A2(n18394), .B1(n20756), .B2(n18395), .ZN(
        n18390) );
  AOI22_X1 U21453 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18396), .B1(
        n18600), .B2(n18469), .ZN(n18389) );
  OAI211_X1 U21454 ( .C1(n20762), .C2(n18425), .A(n18390), .B(n18389), .ZN(
        P3_U2937) );
  AOI22_X1 U21455 ( .A1(n18417), .A2(n18605), .B1(n18604), .B2(n18394), .ZN(
        n18392) );
  AOI22_X1 U21456 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18396), .B1(
        n18606), .B2(n18469), .ZN(n18391) );
  OAI211_X1 U21457 ( .C1(n18393), .C2(n18609), .A(n18392), .B(n18391), .ZN(
        P3_U2938) );
  AOI22_X1 U21458 ( .A1(n18395), .A2(n18556), .B1(n18613), .B2(n18394), .ZN(
        n18398) );
  AOI22_X1 U21459 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18396), .B1(
        n18615), .B2(n18469), .ZN(n18397) );
  OAI211_X1 U21460 ( .C1(n18425), .C2(n18561), .A(n18398), .B(n18397), .ZN(
        P3_U2939) );
  NOR2_X2 U21461 ( .A1(n18451), .A2(n18399), .ZN(n18500) );
  INV_X1 U21462 ( .A(n18500), .ZN(n18488) );
  NOR2_X1 U21463 ( .A1(n18451), .A2(n18400), .ZN(n18421) );
  AOI22_X1 U21464 ( .A1(n18417), .A2(n18473), .B1(n18564), .B2(n18421), .ZN(
        n18404) );
  INV_X1 U21465 ( .A(n18401), .ZN(n18565) );
  NOR2_X1 U21466 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18451), .ZN(
        n18452) );
  AOI22_X1 U21467 ( .A1(n18568), .A2(n18402), .B1(n18565), .B2(n18452), .ZN(
        n18422) );
  AOI22_X1 U21468 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18422), .B1(
        n18563), .B2(n18447), .ZN(n18403) );
  OAI211_X1 U21469 ( .C1(n18481), .C2(n18488), .A(n18404), .B(n18403), .ZN(
        P3_U2940) );
  AOI22_X1 U21470 ( .A1(n18576), .A2(n18447), .B1(n18573), .B2(n18421), .ZN(
        n18406) );
  AOI22_X1 U21471 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18422), .B1(
        n18417), .B2(n18575), .ZN(n18405) );
  OAI211_X1 U21472 ( .C1(n18580), .C2(n18488), .A(n18406), .B(n18405), .ZN(
        P3_U2941) );
  AOI22_X1 U21473 ( .A1(n18417), .A2(n18511), .B1(n18582), .B2(n18421), .ZN(
        n18408) );
  AOI22_X1 U21474 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18422), .B1(
        n18581), .B2(n18447), .ZN(n18407) );
  OAI211_X1 U21475 ( .C1(n18409), .C2(n18488), .A(n18408), .B(n18407), .ZN(
        P3_U2942) );
  AOI22_X1 U21476 ( .A1(n18588), .A2(n18447), .B1(n18587), .B2(n18421), .ZN(
        n18411) );
  AOI22_X1 U21477 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18422), .B1(
        n18417), .B2(n18543), .ZN(n18410) );
  OAI211_X1 U21478 ( .C1(n18412), .C2(n18488), .A(n18411), .B(n18410), .ZN(
        P3_U2943) );
  AOI22_X1 U21479 ( .A1(n18417), .A2(n18489), .B1(n18594), .B2(n18421), .ZN(
        n18414) );
  AOI22_X1 U21480 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18422), .B1(
        n18593), .B2(n18447), .ZN(n18413) );
  OAI211_X1 U21481 ( .C1(n18492), .C2(n18488), .A(n18414), .B(n18413), .ZN(
        P3_U2944) );
  AOI22_X1 U21482 ( .A1(n20757), .A2(n18421), .B1(n20756), .B2(n18417), .ZN(
        n18416) );
  AOI22_X1 U21483 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18422), .B1(
        n18599), .B2(n18447), .ZN(n18415) );
  OAI211_X1 U21484 ( .C1(n20760), .C2(n18488), .A(n18416), .B(n18415), .ZN(
        P3_U2945) );
  AOI22_X1 U21485 ( .A1(n18417), .A2(n18495), .B1(n18604), .B2(n18421), .ZN(
        n18419) );
  AOI22_X1 U21486 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18422), .B1(
        n18605), .B2(n18447), .ZN(n18418) );
  OAI211_X1 U21487 ( .C1(n18420), .C2(n18488), .A(n18419), .B(n18418), .ZN(
        P3_U2946) );
  AOI22_X1 U21488 ( .A1(n18613), .A2(n18421), .B1(n18611), .B2(n18447), .ZN(
        n18424) );
  AOI22_X1 U21489 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18422), .B1(
        n18615), .B2(n18500), .ZN(n18423) );
  OAI211_X1 U21490 ( .C1(n18425), .C2(n18620), .A(n18424), .B(n18423), .ZN(
        P3_U2947) );
  NOR2_X2 U21491 ( .A1(n18451), .A2(n18426), .ZN(n18519) );
  INV_X1 U21492 ( .A(n18519), .ZN(n18528) );
  NOR2_X1 U21493 ( .A1(n18451), .A2(n18530), .ZN(n18446) );
  AOI22_X1 U21494 ( .A1(n18473), .A2(n18447), .B1(n18564), .B2(n18446), .ZN(
        n18430) );
  NOR2_X1 U21495 ( .A1(n18469), .A2(n18447), .ZN(n18427) );
  AOI221_X1 U21496 ( .B1(n18427), .B2(n18488), .C1(n18532), .C2(n18488), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18428) );
  OAI21_X1 U21497 ( .B1(n18519), .B2(n18428), .A(n18535), .ZN(n18448) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18448), .B1(
        n18563), .B2(n18469), .ZN(n18429) );
  OAI211_X1 U21499 ( .C1(n18481), .C2(n18528), .A(n18430), .B(n18429), .ZN(
        P3_U2948) );
  AOI22_X1 U21500 ( .A1(n18576), .A2(n18469), .B1(n18573), .B2(n18446), .ZN(
        n18433) );
  AOI22_X1 U21501 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18448), .B1(
        n18431), .B2(n18519), .ZN(n18432) );
  OAI211_X1 U21502 ( .C1(n18434), .C2(n18445), .A(n18433), .B(n18432), .ZN(
        P3_U2949) );
  AOI22_X1 U21503 ( .A1(n18511), .A2(n18447), .B1(n18582), .B2(n18446), .ZN(
        n18436) );
  AOI22_X1 U21504 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18448), .B1(
        n18583), .B2(n18519), .ZN(n18435) );
  OAI211_X1 U21505 ( .C1(n18514), .C2(n18467), .A(n18436), .B(n18435), .ZN(
        P3_U2950) );
  AOI22_X1 U21506 ( .A1(n18588), .A2(n18469), .B1(n18587), .B2(n18446), .ZN(
        n18438) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18448), .B1(
        n18589), .B2(n18519), .ZN(n18437) );
  OAI211_X1 U21508 ( .C1(n18592), .C2(n18445), .A(n18438), .B(n18437), .ZN(
        P3_U2951) );
  AOI22_X1 U21509 ( .A1(n18594), .A2(n18446), .B1(n18593), .B2(n18469), .ZN(
        n18440) );
  AOI22_X1 U21510 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18448), .B1(
        n18595), .B2(n18519), .ZN(n18439) );
  OAI211_X1 U21511 ( .C1(n18598), .C2(n18445), .A(n18440), .B(n18439), .ZN(
        P3_U2952) );
  AOI22_X1 U21512 ( .A1(n18599), .A2(n18469), .B1(n20757), .B2(n18446), .ZN(
        n18442) );
  AOI22_X1 U21513 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18448), .B1(
        n18600), .B2(n18519), .ZN(n18441) );
  OAI211_X1 U21514 ( .C1(n18603), .C2(n18445), .A(n18442), .B(n18441), .ZN(
        P3_U2953) );
  AOI22_X1 U21515 ( .A1(n18605), .A2(n18469), .B1(n18604), .B2(n18446), .ZN(
        n18444) );
  AOI22_X1 U21516 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18448), .B1(
        n18606), .B2(n18519), .ZN(n18443) );
  OAI211_X1 U21517 ( .C1(n18609), .C2(n18445), .A(n18444), .B(n18443), .ZN(
        P3_U2954) );
  AOI22_X1 U21518 ( .A1(n18556), .A2(n18447), .B1(n18613), .B2(n18446), .ZN(
        n18450) );
  AOI22_X1 U21519 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18448), .B1(
        n18615), .B2(n18519), .ZN(n18449) );
  OAI211_X1 U21520 ( .C1(n18561), .C2(n18467), .A(n18450), .B(n18449), .ZN(
        P3_U2955) );
  NOR2_X1 U21521 ( .A1(n18638), .A2(n18451), .ZN(n18505) );
  AND2_X1 U21522 ( .A1(n18562), .A2(n18505), .ZN(n18468) );
  AOI22_X1 U21523 ( .A1(n18564), .A2(n18468), .B1(n18563), .B2(n18500), .ZN(
        n18454) );
  AOI22_X1 U21524 ( .A1(n18568), .A2(n18452), .B1(n18565), .B2(n18505), .ZN(
        n18470) );
  NAND2_X1 U21525 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18505), .ZN(
        n18553) );
  INV_X1 U21526 ( .A(n18553), .ZN(n18555) );
  AOI22_X1 U21527 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18470), .B1(
        n18569), .B2(n18555), .ZN(n18453) );
  OAI211_X1 U21528 ( .C1(n18572), .C2(n18467), .A(n18454), .B(n18453), .ZN(
        P3_U2956) );
  AOI22_X1 U21529 ( .A1(n18575), .A2(n18469), .B1(n18573), .B2(n18468), .ZN(
        n18456) );
  AOI22_X1 U21530 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18470), .B1(
        n18576), .B2(n18500), .ZN(n18455) );
  OAI211_X1 U21531 ( .C1(n18580), .C2(n18553), .A(n18456), .B(n18455), .ZN(
        P3_U2957) );
  AOI22_X1 U21532 ( .A1(n18582), .A2(n18468), .B1(n18581), .B2(n18500), .ZN(
        n18458) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18470), .B1(
        n18583), .B2(n18555), .ZN(n18457) );
  OAI211_X1 U21534 ( .C1(n18586), .C2(n18467), .A(n18458), .B(n18457), .ZN(
        P3_U2958) );
  AOI22_X1 U21535 ( .A1(n18588), .A2(n18500), .B1(n18587), .B2(n18468), .ZN(
        n18460) );
  AOI22_X1 U21536 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18470), .B1(
        n18589), .B2(n18555), .ZN(n18459) );
  OAI211_X1 U21537 ( .C1(n18592), .C2(n18467), .A(n18460), .B(n18459), .ZN(
        P3_U2959) );
  AOI22_X1 U21538 ( .A1(n18594), .A2(n18468), .B1(n18593), .B2(n18500), .ZN(
        n18462) );
  AOI22_X1 U21539 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18470), .B1(
        n18595), .B2(n18555), .ZN(n18461) );
  OAI211_X1 U21540 ( .C1(n18598), .C2(n18467), .A(n18462), .B(n18461), .ZN(
        P3_U2960) );
  AOI22_X1 U21541 ( .A1(n20757), .A2(n18468), .B1(n20756), .B2(n18469), .ZN(
        n18464) );
  AOI22_X1 U21542 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18470), .B1(
        n18600), .B2(n18555), .ZN(n18463) );
  OAI211_X1 U21543 ( .C1(n20762), .C2(n18488), .A(n18464), .B(n18463), .ZN(
        P3_U2961) );
  AOI22_X1 U21544 ( .A1(n18605), .A2(n18500), .B1(n18604), .B2(n18468), .ZN(
        n18466) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18470), .B1(
        n18606), .B2(n18555), .ZN(n18465) );
  OAI211_X1 U21546 ( .C1(n18609), .C2(n18467), .A(n18466), .B(n18465), .ZN(
        P3_U2962) );
  AOI22_X1 U21547 ( .A1(n18556), .A2(n18469), .B1(n18613), .B2(n18468), .ZN(
        n18472) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18470), .B1(
        n18615), .B2(n18555), .ZN(n18471) );
  OAI211_X1 U21549 ( .C1(n18561), .C2(n18488), .A(n18472), .B(n18471), .ZN(
        P3_U2963) );
  INV_X1 U21550 ( .A(n18567), .ZN(n18504) );
  NOR2_X2 U21551 ( .A1(n18504), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18574) );
  INV_X1 U21552 ( .A(n18574), .ZN(n18619) );
  NOR2_X1 U21553 ( .A1(n18555), .A2(n18574), .ZN(n18533) );
  NOR2_X1 U21554 ( .A1(n18691), .A2(n18533), .ZN(n18499) );
  AOI22_X1 U21555 ( .A1(n18473), .A2(n18500), .B1(n18564), .B2(n18499), .ZN(
        n18480) );
  NAND2_X1 U21556 ( .A1(n18475), .A2(n18474), .ZN(n18476) );
  OAI21_X1 U21557 ( .B1(n18477), .B2(n18476), .A(n18533), .ZN(n18478) );
  OAI211_X1 U21558 ( .C1(n18574), .C2(n18794), .A(n18535), .B(n18478), .ZN(
        n18501) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18501), .B1(
        n18563), .B2(n18519), .ZN(n18479) );
  OAI211_X1 U21560 ( .C1(n18481), .C2(n18619), .A(n18480), .B(n18479), .ZN(
        P3_U2964) );
  AOI22_X1 U21561 ( .A1(n18575), .A2(n18500), .B1(n18573), .B2(n18499), .ZN(
        n18483) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18501), .B1(
        n18576), .B2(n18519), .ZN(n18482) );
  OAI211_X1 U21563 ( .C1(n18580), .C2(n18619), .A(n18483), .B(n18482), .ZN(
        P3_U2965) );
  AOI22_X1 U21564 ( .A1(n18511), .A2(n18500), .B1(n18582), .B2(n18499), .ZN(
        n18485) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18501), .B1(
        n18583), .B2(n18574), .ZN(n18484) );
  OAI211_X1 U21566 ( .C1(n18514), .C2(n18528), .A(n18485), .B(n18484), .ZN(
        P3_U2966) );
  AOI22_X1 U21567 ( .A1(n18588), .A2(n18519), .B1(n18587), .B2(n18499), .ZN(
        n18487) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18501), .B1(
        n18589), .B2(n18574), .ZN(n18486) );
  OAI211_X1 U21569 ( .C1(n18592), .C2(n18488), .A(n18487), .B(n18486), .ZN(
        P3_U2967) );
  AOI22_X1 U21570 ( .A1(n18489), .A2(n18500), .B1(n18594), .B2(n18499), .ZN(
        n18491) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18501), .B1(
        n18593), .B2(n18519), .ZN(n18490) );
  OAI211_X1 U21572 ( .C1(n18492), .C2(n18619), .A(n18491), .B(n18490), .ZN(
        P3_U2968) );
  AOI22_X1 U21573 ( .A1(n20757), .A2(n18499), .B1(n20756), .B2(n18500), .ZN(
        n18494) );
  AOI22_X1 U21574 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18501), .B1(
        n18600), .B2(n18574), .ZN(n18493) );
  OAI211_X1 U21575 ( .C1(n20762), .C2(n18528), .A(n18494), .B(n18493), .ZN(
        P3_U2969) );
  AOI22_X1 U21576 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18501), .B1(
        n18604), .B2(n18499), .ZN(n18497) );
  AOI22_X1 U21577 ( .A1(n18606), .A2(n18574), .B1(n18495), .B2(n18500), .ZN(
        n18496) );
  OAI211_X1 U21578 ( .C1(n18498), .C2(n18528), .A(n18497), .B(n18496), .ZN(
        P3_U2970) );
  AOI22_X1 U21579 ( .A1(n18556), .A2(n18500), .B1(n18613), .B2(n18499), .ZN(
        n18503) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18501), .B1(
        n18615), .B2(n18574), .ZN(n18502) );
  OAI211_X1 U21581 ( .C1(n18561), .C2(n18528), .A(n18503), .B(n18502), .ZN(
        P3_U2971) );
  NOR2_X1 U21582 ( .A1(n18691), .A2(n18504), .ZN(n18524) );
  AOI22_X1 U21583 ( .A1(n18564), .A2(n18524), .B1(n18563), .B2(n18555), .ZN(
        n18507) );
  AOI22_X1 U21584 ( .A1(n18568), .A2(n18505), .B1(n18567), .B2(n18565), .ZN(
        n18525) );
  AOI22_X1 U21585 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18525), .B1(
        n18569), .B2(n18610), .ZN(n18506) );
  OAI211_X1 U21586 ( .C1(n18572), .C2(n18528), .A(n18507), .B(n18506), .ZN(
        P3_U2972) );
  AOI22_X1 U21587 ( .A1(n18575), .A2(n18519), .B1(n18573), .B2(n18524), .ZN(
        n18509) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18525), .B1(
        n18576), .B2(n18555), .ZN(n18508) );
  OAI211_X1 U21589 ( .C1(n18580), .C2(n18510), .A(n18509), .B(n18508), .ZN(
        P3_U2973) );
  AOI22_X1 U21590 ( .A1(n18511), .A2(n18519), .B1(n18582), .B2(n18524), .ZN(
        n18513) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18525), .B1(
        n18583), .B2(n18610), .ZN(n18512) );
  OAI211_X1 U21592 ( .C1(n18514), .C2(n18553), .A(n18513), .B(n18512), .ZN(
        P3_U2974) );
  AOI22_X1 U21593 ( .A1(n18588), .A2(n18555), .B1(n18587), .B2(n18524), .ZN(
        n18516) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18525), .B1(
        n18589), .B2(n18610), .ZN(n18515) );
  OAI211_X1 U21595 ( .C1(n18592), .C2(n18528), .A(n18516), .B(n18515), .ZN(
        P3_U2975) );
  AOI22_X1 U21596 ( .A1(n18594), .A2(n18524), .B1(n18593), .B2(n18555), .ZN(
        n18518) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18525), .B1(
        n18595), .B2(n18610), .ZN(n18517) );
  OAI211_X1 U21598 ( .C1(n18598), .C2(n18528), .A(n18518), .B(n18517), .ZN(
        P3_U2976) );
  AOI22_X1 U21599 ( .A1(n20757), .A2(n18524), .B1(n20756), .B2(n18519), .ZN(
        n18521) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18525), .B1(
        n18600), .B2(n18610), .ZN(n18520) );
  OAI211_X1 U21601 ( .C1(n20762), .C2(n18553), .A(n18521), .B(n18520), .ZN(
        P3_U2977) );
  AOI22_X1 U21602 ( .A1(n18605), .A2(n18555), .B1(n18604), .B2(n18524), .ZN(
        n18523) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18525), .B1(
        n18606), .B2(n18610), .ZN(n18522) );
  OAI211_X1 U21604 ( .C1(n18609), .C2(n18528), .A(n18523), .B(n18522), .ZN(
        P3_U2978) );
  AOI22_X1 U21605 ( .A1(n18613), .A2(n18524), .B1(n18611), .B2(n18555), .ZN(
        n18527) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18525), .B1(
        n18615), .B2(n18610), .ZN(n18526) );
  OAI211_X1 U21607 ( .C1(n18620), .C2(n18528), .A(n18527), .B(n18526), .ZN(
        P3_U2979) );
  NOR2_X1 U21608 ( .A1(n18530), .A2(n18529), .ZN(n18554) );
  AOI22_X1 U21609 ( .A1(n18564), .A2(n18554), .B1(n18563), .B2(n18574), .ZN(
        n18537) );
  OAI21_X1 U21610 ( .B1(n18533), .B2(n18532), .A(n18531), .ZN(n18534) );
  OAI211_X1 U21611 ( .C1(n18557), .C2(n18794), .A(n18535), .B(n18534), .ZN(
        n18558) );
  AOI22_X1 U21612 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18558), .B1(
        n18569), .B2(n18557), .ZN(n18536) );
  OAI211_X1 U21613 ( .C1(n18572), .C2(n18553), .A(n18537), .B(n18536), .ZN(
        P3_U2980) );
  AOI22_X1 U21614 ( .A1(n18575), .A2(n18555), .B1(n18573), .B2(n18554), .ZN(
        n18539) );
  AOI22_X1 U21615 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18558), .B1(
        n18576), .B2(n18574), .ZN(n18538) );
  OAI211_X1 U21616 ( .C1(n18580), .C2(n18540), .A(n18539), .B(n18538), .ZN(
        P3_U2981) );
  AOI22_X1 U21617 ( .A1(n18582), .A2(n18554), .B1(n18581), .B2(n18574), .ZN(
        n18542) );
  AOI22_X1 U21618 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18558), .B1(
        n18583), .B2(n18557), .ZN(n18541) );
  OAI211_X1 U21619 ( .C1(n18586), .C2(n18553), .A(n18542), .B(n18541), .ZN(
        P3_U2982) );
  AOI22_X1 U21620 ( .A1(n18587), .A2(n18554), .B1(n18543), .B2(n18555), .ZN(
        n18545) );
  AOI22_X1 U21621 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18558), .B1(
        n18589), .B2(n18557), .ZN(n18544) );
  OAI211_X1 U21622 ( .C1(n18546), .C2(n18619), .A(n18545), .B(n18544), .ZN(
        P3_U2983) );
  AOI22_X1 U21623 ( .A1(n18594), .A2(n18554), .B1(n18593), .B2(n18574), .ZN(
        n18548) );
  AOI22_X1 U21624 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18558), .B1(
        n18595), .B2(n18557), .ZN(n18547) );
  OAI211_X1 U21625 ( .C1(n18598), .C2(n18553), .A(n18548), .B(n18547), .ZN(
        P3_U2984) );
  AOI22_X1 U21626 ( .A1(n20757), .A2(n18554), .B1(n20756), .B2(n18555), .ZN(
        n18550) );
  AOI22_X1 U21627 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18558), .B1(
        n18600), .B2(n18557), .ZN(n18549) );
  OAI211_X1 U21628 ( .C1(n20762), .C2(n18619), .A(n18550), .B(n18549), .ZN(
        P3_U2985) );
  AOI22_X1 U21629 ( .A1(n18605), .A2(n18574), .B1(n18604), .B2(n18554), .ZN(
        n18552) );
  AOI22_X1 U21630 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18558), .B1(
        n18606), .B2(n18557), .ZN(n18551) );
  OAI211_X1 U21631 ( .C1(n18609), .C2(n18553), .A(n18552), .B(n18551), .ZN(
        P3_U2986) );
  AOI22_X1 U21632 ( .A1(n18556), .A2(n18555), .B1(n18613), .B2(n18554), .ZN(
        n18560) );
  AOI22_X1 U21633 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18558), .B1(
        n18615), .B2(n18557), .ZN(n18559) );
  OAI211_X1 U21634 ( .C1(n18561), .C2(n18619), .A(n18560), .B(n18559), .ZN(
        P3_U2987) );
  AND2_X1 U21635 ( .A1(n18562), .A2(n18566), .ZN(n18612) );
  AOI22_X1 U21636 ( .A1(n18564), .A2(n18612), .B1(n18563), .B2(n18610), .ZN(
        n18571) );
  AOI22_X1 U21637 ( .A1(n18568), .A2(n18567), .B1(n18566), .B2(n18565), .ZN(
        n18616) );
  AOI22_X1 U21638 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18616), .B1(
        n18569), .B2(n18614), .ZN(n18570) );
  OAI211_X1 U21639 ( .C1(n18572), .C2(n18619), .A(n18571), .B(n18570), .ZN(
        P3_U2988) );
  AOI22_X1 U21640 ( .A1(n18575), .A2(n18574), .B1(n18573), .B2(n18612), .ZN(
        n18578) );
  AOI22_X1 U21641 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18616), .B1(
        n18576), .B2(n18610), .ZN(n18577) );
  OAI211_X1 U21642 ( .C1(n18580), .C2(n18579), .A(n18578), .B(n18577), .ZN(
        P3_U2989) );
  AOI22_X1 U21643 ( .A1(n18582), .A2(n18612), .B1(n18581), .B2(n18610), .ZN(
        n18585) );
  AOI22_X1 U21644 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18616), .B1(
        n18583), .B2(n18614), .ZN(n18584) );
  OAI211_X1 U21645 ( .C1(n18586), .C2(n18619), .A(n18585), .B(n18584), .ZN(
        P3_U2990) );
  AOI22_X1 U21646 ( .A1(n18588), .A2(n18610), .B1(n18587), .B2(n18612), .ZN(
        n18591) );
  AOI22_X1 U21647 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18616), .B1(
        n18589), .B2(n18614), .ZN(n18590) );
  OAI211_X1 U21648 ( .C1(n18592), .C2(n18619), .A(n18591), .B(n18590), .ZN(
        P3_U2991) );
  AOI22_X1 U21649 ( .A1(n18594), .A2(n18612), .B1(n18593), .B2(n18610), .ZN(
        n18597) );
  AOI22_X1 U21650 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18616), .B1(
        n18595), .B2(n18614), .ZN(n18596) );
  OAI211_X1 U21651 ( .C1(n18598), .C2(n18619), .A(n18597), .B(n18596), .ZN(
        P3_U2992) );
  AOI22_X1 U21652 ( .A1(n18599), .A2(n18610), .B1(n20757), .B2(n18612), .ZN(
        n18602) );
  AOI22_X1 U21653 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18616), .B1(
        n18600), .B2(n18614), .ZN(n18601) );
  OAI211_X1 U21654 ( .C1(n18603), .C2(n18619), .A(n18602), .B(n18601), .ZN(
        P3_U2993) );
  AOI22_X1 U21655 ( .A1(n18605), .A2(n18610), .B1(n18604), .B2(n18612), .ZN(
        n18608) );
  AOI22_X1 U21656 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18616), .B1(
        n18606), .B2(n18614), .ZN(n18607) );
  OAI211_X1 U21657 ( .C1(n18609), .C2(n18619), .A(n18608), .B(n18607), .ZN(
        P3_U2994) );
  AOI22_X1 U21658 ( .A1(n18613), .A2(n18612), .B1(n18611), .B2(n18610), .ZN(
        n18618) );
  AOI22_X1 U21659 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18616), .B1(
        n18615), .B2(n18614), .ZN(n18617) );
  OAI211_X1 U21660 ( .C1(n18620), .C2(n18619), .A(n18618), .B(n18617), .ZN(
        P3_U2995) );
  AOI22_X1 U21661 ( .A1(n18624), .A2(n18623), .B1(n18622), .B2(n18621), .ZN(
        n18625) );
  OAI221_X1 U21662 ( .B1(n18627), .B2(n18648), .C1(n18627), .C2(n18626), .A(
        n18625), .ZN(n18834) );
  OAI21_X1 U21663 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18628), .ZN(n18629) );
  OAI211_X1 U21664 ( .C1(n18631), .C2(n18664), .A(n18630), .B(n18629), .ZN(
        n18676) );
  OR2_X1 U21665 ( .A1(n18633), .A2(n18632), .ZN(n18636) );
  OAI21_X1 U21666 ( .B1(n18635), .B2(n18821), .A(n18634), .ZN(n18651) );
  AOI22_X1 U21667 ( .A1(n18812), .A2(n18636), .B1(n12565), .B2(n18651), .ZN(
        n18809) );
  AOI22_X1 U21668 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18658), .B1(
        n18636), .B2(n18821), .ZN(n18639) );
  INV_X1 U21669 ( .A(n18639), .ZN(n18816) );
  NOR3_X1 U21670 ( .A1(n18638), .A2(n18637), .A3(n18816), .ZN(n18640) );
  OAI22_X1 U21671 ( .A1(n18809), .A2(n18640), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18639), .ZN(n18642) );
  AOI21_X1 U21672 ( .B1(n18642), .B2(n18664), .A(n18641), .ZN(n18667) );
  NOR2_X1 U21673 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18667), .ZN(
        n18649) );
  OAI21_X1 U21674 ( .B1(n18645), .B2(n18644), .A(n18643), .ZN(n18656) );
  NAND3_X1 U21675 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18650), .A3(
        n18656), .ZN(n18647) );
  OAI211_X1 U21676 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n18651), .B(n18657), .ZN(
        n18646) );
  OAI211_X1 U21677 ( .C1(n18804), .C2(n18648), .A(n18647), .B(n18646), .ZN(
        n18806) );
  MUX2_X1 U21678 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n18806), .S(
        n18664), .Z(n18668) );
  AOI221_X1 U21679 ( .B1(n18649), .B2(n18666), .C1(n18665), .C2(n18666), .A(
        n18668), .ZN(n18674) );
  NAND2_X1 U21680 ( .A1(n18650), .A2(n18808), .ZN(n18653) );
  AOI22_X1 U21681 ( .A1(n18654), .A2(n18653), .B1(n18652), .B2(n18651), .ZN(
        n18655) );
  NOR2_X1 U21682 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18655), .ZN(
        n18796) );
  AOI21_X1 U21683 ( .B1(n18658), .B2(n18657), .A(n18656), .ZN(n18659) );
  OAI22_X1 U21684 ( .A1(n18661), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18660), .B2(n18659), .ZN(n18797) );
  INV_X1 U21685 ( .A(n18797), .ZN(n18662) );
  NAND2_X1 U21686 ( .A1(n18664), .A2(n18662), .ZN(n18663) );
  AOI22_X1 U21687 ( .A1(n18664), .A2(n18796), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18663), .ZN(n18673) );
  NAND2_X1 U21688 ( .A1(n18666), .A2(n18665), .ZN(n18672) );
  INV_X1 U21689 ( .A(n18667), .ZN(n18669) );
  AOI222_X1 U21690 ( .A1(n18670), .A2(n18669), .B1(n18670), .B2(n18668), .C1(
        n18669), .C2(n18668), .ZN(n18671) );
  OAI22_X1 U21691 ( .A1(n18674), .A2(n18673), .B1(n18672), .B2(n18671), .ZN(
        n18675) );
  NOR4_X1 U21692 ( .A1(n18677), .A2(n18834), .A3(n18676), .A4(n18675), .ZN(
        n18687) );
  AOI22_X1 U21693 ( .A1(n18815), .A2(n18845), .B1(n18836), .B2(n17411), .ZN(
        n18678) );
  INV_X1 U21694 ( .A(n18678), .ZN(n18684) );
  OAI211_X1 U21695 ( .C1(n18681), .C2(n18680), .A(n18679), .B(n18687), .ZN(
        n18793) );
  OAI21_X1 U21696 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18843), .A(n18793), 
        .ZN(n18689) );
  NOR2_X1 U21697 ( .A1(n18682), .A2(n18689), .ZN(n18683) );
  MUX2_X1 U21698 ( .A(n18684), .B(n18683), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18686) );
  OAI211_X1 U21699 ( .C1(n18687), .C2(n18839), .A(n18686), .B(n18685), .ZN(
        P3_U2996) );
  NAND2_X1 U21700 ( .A1(n18836), .A2(n17411), .ZN(n18693) );
  NAND3_X1 U21701 ( .A1(n18836), .A2(n18696), .A3(n18688), .ZN(n18695) );
  OR3_X1 U21702 ( .A1(n18691), .A2(n18690), .A3(n18689), .ZN(n18692) );
  NAND4_X1 U21703 ( .A1(n18694), .A2(n18693), .A3(n18695), .A4(n18692), .ZN(
        P3_U2997) );
  INV_X1 U21704 ( .A(n18695), .ZN(n18700) );
  NOR3_X1 U21705 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18697), .A3(n18696), 
        .ZN(n18698) );
  NOR3_X1 U21706 ( .A1(n18700), .A2(n18699), .A3(n18698), .ZN(P3_U2998) );
  AND2_X1 U21707 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18701), .ZN(
        P3_U2999) );
  AND2_X1 U21708 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18790), .ZN(
        P3_U3000) );
  AND2_X1 U21709 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18790), .ZN(
        P3_U3001) );
  AND2_X1 U21710 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18790), .ZN(
        P3_U3002) );
  AND2_X1 U21711 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18790), .ZN(
        P3_U3003) );
  AND2_X1 U21712 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18790), .ZN(
        P3_U3004) );
  AND2_X1 U21713 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18790), .ZN(
        P3_U3005) );
  AND2_X1 U21714 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18790), .ZN(
        P3_U3006) );
  AND2_X1 U21715 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18790), .ZN(
        P3_U3007) );
  AND2_X1 U21716 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18790), .ZN(
        P3_U3008) );
  AND2_X1 U21717 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18790), .ZN(
        P3_U3009) );
  AND2_X1 U21718 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18790), .ZN(
        P3_U3010) );
  AND2_X1 U21719 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18790), .ZN(
        P3_U3011) );
  AND2_X1 U21720 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18790), .ZN(
        P3_U3012) );
  AND2_X1 U21721 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18790), .ZN(
        P3_U3013) );
  AND2_X1 U21722 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18790), .ZN(
        P3_U3014) );
  AND2_X1 U21723 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18790), .ZN(
        P3_U3015) );
  AND2_X1 U21724 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18790), .ZN(
        P3_U3016) );
  AND2_X1 U21725 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18790), .ZN(
        P3_U3017) );
  AND2_X1 U21726 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18790), .ZN(
        P3_U3018) );
  AND2_X1 U21727 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18790), .ZN(
        P3_U3019) );
  AND2_X1 U21728 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18790), .ZN(
        P3_U3020) );
  AND2_X1 U21729 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18790), .ZN(P3_U3021) );
  AND2_X1 U21730 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18790), .ZN(P3_U3022) );
  AND2_X1 U21731 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18790), .ZN(P3_U3023) );
  AND2_X1 U21732 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18790), .ZN(P3_U3024) );
  AND2_X1 U21733 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18790), .ZN(P3_U3025) );
  AND2_X1 U21734 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18790), .ZN(P3_U3026) );
  AND2_X1 U21735 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18790), .ZN(P3_U3027) );
  AND2_X1 U21736 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18790), .ZN(P3_U3028) );
  NAND2_X1 U21737 ( .A1(n18836), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18712) );
  INV_X1 U21738 ( .A(n18712), .ZN(n18709) );
  OAI21_X1 U21739 ( .B1(n18703), .B2(n20639), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18704) );
  AOI22_X1 U21740 ( .A1(n18709), .A2(n18718), .B1(n18851), .B2(n18704), .ZN(
        n18706) );
  NAND3_X1 U21741 ( .A1(NA), .A2(n18716), .A3(n18705), .ZN(n18710) );
  OAI211_X1 U21742 ( .C1(P3_STATE_REG_0__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18706), .B(n18710), .ZN(P3_U3029) );
  NAND2_X1 U21743 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n18711) );
  AOI22_X1 U21744 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n18711), .B1(HOLD), 
        .B2(n18707), .ZN(n18708) );
  OAI211_X1 U21745 ( .C1(n18708), .C2(n18716), .A(n18712), .B(n18840), .ZN(
        P3_U3030) );
  AOI21_X1 U21746 ( .B1(n18716), .B2(n18710), .A(n18709), .ZN(n18717) );
  INV_X1 U21747 ( .A(n18711), .ZN(n18714) );
  OAI22_X1 U21748 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18712), .ZN(n18713) );
  OAI22_X1 U21749 ( .A1(n18714), .A2(n18713), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18715) );
  OAI22_X1 U21750 ( .A1(n18717), .A2(n18718), .B1(n18716), .B2(n18715), .ZN(
        P3_U3031) );
  OAI222_X1 U21751 ( .A1(n18720), .A2(n9591), .B1(n18719), .B2(n18850), .C1(
        n18721), .C2(n18768), .ZN(P3_U3032) );
  INV_X1 U21752 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18723) );
  OAI222_X1 U21753 ( .A1(n18768), .A2(n18723), .B1(n18722), .B2(n18780), .C1(
        n18721), .C2(n9591), .ZN(P3_U3033) );
  OAI222_X1 U21754 ( .A1(n18768), .A2(n18726), .B1(n18724), .B2(n18850), .C1(
        n18723), .C2(n9591), .ZN(P3_U3034) );
  OAI222_X1 U21755 ( .A1(n18768), .A2(n18729), .B1(n18727), .B2(n18780), .C1(
        n18726), .C2(n9591), .ZN(P3_U3035) );
  OAI222_X1 U21756 ( .A1(n18729), .A2(n9591), .B1(n18728), .B2(n18850), .C1(
        n18730), .C2(n18768), .ZN(P3_U3036) );
  OAI222_X1 U21757 ( .A1(n18768), .A2(n18732), .B1(n18731), .B2(n18850), .C1(
        n18730), .C2(n9591), .ZN(P3_U3037) );
  OAI222_X1 U21758 ( .A1(n18768), .A2(n18734), .B1(n18733), .B2(n18786), .C1(
        n18732), .C2(n9591), .ZN(P3_U3038) );
  OAI222_X1 U21759 ( .A1(n18768), .A2(n18736), .B1(n18735), .B2(n18850), .C1(
        n18734), .C2(n9591), .ZN(P3_U3039) );
  OAI222_X1 U21760 ( .A1(n18768), .A2(n18738), .B1(n18737), .B2(n18850), .C1(
        n18736), .C2(n9591), .ZN(P3_U3040) );
  OAI222_X1 U21761 ( .A1(n18768), .A2(n18740), .B1(n18739), .B2(n18850), .C1(
        n18738), .C2(n9591), .ZN(P3_U3041) );
  OAI222_X1 U21762 ( .A1(n18768), .A2(n18742), .B1(n18741), .B2(n18850), .C1(
        n18740), .C2(n9591), .ZN(P3_U3042) );
  OAI222_X1 U21763 ( .A1(n18768), .A2(n18744), .B1(n18743), .B2(n18850), .C1(
        n18742), .C2(n9591), .ZN(P3_U3043) );
  INV_X1 U21764 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18747) );
  OAI222_X1 U21765 ( .A1(n18768), .A2(n18747), .B1(n18745), .B2(n18850), .C1(
        n18744), .C2(n9591), .ZN(P3_U3044) );
  OAI222_X1 U21766 ( .A1(n18747), .A2(n9591), .B1(n18746), .B2(n18850), .C1(
        n18748), .C2(n18768), .ZN(P3_U3045) );
  OAI222_X1 U21767 ( .A1(n18768), .A2(n18750), .B1(n18749), .B2(n18850), .C1(
        n18748), .C2(n9591), .ZN(P3_U3046) );
  OAI222_X1 U21768 ( .A1(n18768), .A2(n18753), .B1(n18751), .B2(n18850), .C1(
        n18750), .C2(n9591), .ZN(P3_U3047) );
  OAI222_X1 U21769 ( .A1(n18753), .A2(n9591), .B1(n18752), .B2(n18850), .C1(
        n18754), .C2(n18768), .ZN(P3_U3048) );
  OAI222_X1 U21770 ( .A1(n18768), .A2(n18756), .B1(n18755), .B2(n18850), .C1(
        n18754), .C2(n9591), .ZN(P3_U3049) );
  OAI222_X1 U21771 ( .A1(n18768), .A2(n18759), .B1(n18757), .B2(n18850), .C1(
        n18756), .C2(n9591), .ZN(P3_U3050) );
  OAI222_X1 U21772 ( .A1(n18759), .A2(n9591), .B1(n18758), .B2(n18850), .C1(
        n18760), .C2(n18768), .ZN(P3_U3051) );
  OAI222_X1 U21773 ( .A1(n18768), .A2(n18762), .B1(n18761), .B2(n18850), .C1(
        n18760), .C2(n9591), .ZN(P3_U3052) );
  OAI222_X1 U21774 ( .A1(n18768), .A2(n18764), .B1(n18763), .B2(n18850), .C1(
        n18762), .C2(n9591), .ZN(P3_U3053) );
  OAI222_X1 U21775 ( .A1(n18768), .A2(n18766), .B1(n18765), .B2(n18780), .C1(
        n18764), .C2(n9591), .ZN(P3_U3054) );
  OAI222_X1 U21776 ( .A1(n18768), .A2(n18769), .B1(n18767), .B2(n18780), .C1(
        n18766), .C2(n9591), .ZN(P3_U3055) );
  OAI222_X1 U21777 ( .A1(n18768), .A2(n18771), .B1(n18770), .B2(n18780), .C1(
        n18769), .C2(n9591), .ZN(P3_U3056) );
  OAI222_X1 U21778 ( .A1(n18768), .A2(n18773), .B1(n18772), .B2(n18780), .C1(
        n18771), .C2(n9591), .ZN(P3_U3057) );
  INV_X1 U21779 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18776) );
  OAI222_X1 U21780 ( .A1(n18768), .A2(n18776), .B1(n18774), .B2(n18780), .C1(
        n18773), .C2(n9591), .ZN(P3_U3058) );
  OAI222_X1 U21781 ( .A1(n18776), .A2(n9591), .B1(n18775), .B2(n18780), .C1(
        n18777), .C2(n18768), .ZN(P3_U3059) );
  OAI222_X1 U21782 ( .A1(n18768), .A2(n18782), .B1(n18778), .B2(n18780), .C1(
        n18777), .C2(n9591), .ZN(P3_U3060) );
  OAI222_X1 U21783 ( .A1(n9591), .A2(n18782), .B1(n18781), .B2(n18780), .C1(
        n18779), .C2(n18768), .ZN(P3_U3061) );
  OAI22_X1 U21784 ( .A1(n18851), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18850), .ZN(n18783) );
  INV_X1 U21785 ( .A(n18783), .ZN(P3_U3274) );
  OAI22_X1 U21786 ( .A1(n18851), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18850), .ZN(n18784) );
  INV_X1 U21787 ( .A(n18784), .ZN(P3_U3275) );
  OAI22_X1 U21788 ( .A1(n18851), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18850), .ZN(n18785) );
  INV_X1 U21789 ( .A(n18785), .ZN(P3_U3276) );
  OAI22_X1 U21790 ( .A1(n18851), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18786), .ZN(n18787) );
  INV_X1 U21791 ( .A(n18787), .ZN(P3_U3277) );
  INV_X1 U21792 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18824) );
  INV_X1 U21793 ( .A(n18788), .ZN(n18789) );
  AOI21_X1 U21794 ( .B1(n18790), .B2(n18824), .A(n18789), .ZN(P3_U3280) );
  AOI21_X1 U21795 ( .B1(n18790), .B2(P3_DATAWIDTH_REG_1__SCAN_IN), .A(n18789), 
        .ZN(n18791) );
  INV_X1 U21796 ( .A(n18791), .ZN(P3_U3281) );
  OAI221_X1 U21797 ( .B1(n18794), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18794), 
        .C2(n18793), .A(n18792), .ZN(P3_U3282) );
  AOI22_X1 U21798 ( .A1(n18817), .A2(n18796), .B1(n18815), .B2(n18795), .ZN(
        n18800) );
  AOI21_X1 U21799 ( .B1(n18817), .B2(n18797), .A(n18822), .ZN(n18799) );
  OAI22_X1 U21800 ( .A1(n18822), .A2(n18800), .B1(n18799), .B2(n18798), .ZN(
        P3_U3285) );
  NOR2_X1 U21801 ( .A1(n18801), .A2(n18818), .ZN(n18810) );
  OAI22_X1 U21802 ( .A1(n18803), .A2(n18802), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18811) );
  INV_X1 U21803 ( .A(n18811), .ZN(n18805) );
  AOI222_X1 U21804 ( .A1(n18806), .A2(n18817), .B1(n18810), .B2(n18805), .C1(
        n18815), .C2(n18804), .ZN(n18807) );
  AOI22_X1 U21805 ( .A1(n18822), .A2(n18808), .B1(n18807), .B2(n18819), .ZN(
        P3_U3288) );
  INV_X1 U21806 ( .A(n18809), .ZN(n18813) );
  AOI222_X1 U21807 ( .A1(n18813), .A2(n18817), .B1(n18815), .B2(n18812), .C1(
        n18811), .C2(n18810), .ZN(n18814) );
  AOI22_X1 U21808 ( .A1(n18822), .A2(n12565), .B1(n18814), .B2(n18819), .ZN(
        P3_U3289) );
  AOI222_X1 U21809 ( .A1(n18818), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18817), 
        .B2(n18816), .C1(n18821), .C2(n18815), .ZN(n18820) );
  AOI22_X1 U21810 ( .A1(n18822), .A2(n18821), .B1(n18820), .B2(n18819), .ZN(
        P3_U3290) );
  NOR3_X1 U21811 ( .A1(n18824), .A2(P3_REIP_REG_0__SCAN_IN), .A3(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18823) );
  AOI221_X1 U21812 ( .B1(n18825), .B2(n18824), .C1(P3_REIP_REG_1__SCAN_IN), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n18823), .ZN(n18827) );
  INV_X1 U21813 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18826) );
  INV_X1 U21814 ( .A(n18831), .ZN(n18828) );
  AOI22_X1 U21815 ( .A1(n18831), .A2(n18827), .B1(n18826), .B2(n18828), .ZN(
        P3_U3292) );
  NOR2_X1 U21816 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n18830) );
  INV_X1 U21817 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18829) );
  AOI22_X1 U21818 ( .A1(n18831), .A2(n18830), .B1(n18829), .B2(n18828), .ZN(
        P3_U3293) );
  INV_X1 U21819 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18832) );
  AOI22_X1 U21820 ( .A1(n18850), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18832), 
        .B2(n18851), .ZN(P3_U3294) );
  MUX2_X1 U21821 ( .A(P3_MORE_REG_SCAN_IN), .B(n18834), .S(n18833), .Z(
        P3_U3295) );
  OAI21_X1 U21822 ( .B1(n18836), .B2(n18835), .A(n18855), .ZN(n18837) );
  AOI21_X1 U21823 ( .B1(n18839), .B2(n18838), .A(n18837), .ZN(n18849) );
  AOI21_X1 U21824 ( .B1(n18842), .B2(n18841), .A(n18840), .ZN(n18844) );
  OAI211_X1 U21825 ( .C1(n18854), .C2(n18844), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18843), .ZN(n18846) );
  AOI21_X1 U21826 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18846), .A(n18845), 
        .ZN(n18848) );
  NAND2_X1 U21827 ( .A1(n18849), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18847) );
  OAI21_X1 U21828 ( .B1(n18849), .B2(n18848), .A(n18847), .ZN(P3_U3296) );
  OAI22_X1 U21829 ( .A1(n18851), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18850), .ZN(n18852) );
  INV_X1 U21830 ( .A(n18852), .ZN(P3_U3297) );
  OAI21_X1 U21831 ( .B1(n18853), .B2(P3_STATE2_REG_2__SCAN_IN), .A(n18855), 
        .ZN(n18858) );
  OAI22_X1 U21832 ( .A1(n18858), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18855), 
        .B2(n18854), .ZN(n18856) );
  INV_X1 U21833 ( .A(n18856), .ZN(P3_U3298) );
  OAI21_X1 U21834 ( .B1(n18858), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n18857), 
        .ZN(n18859) );
  INV_X1 U21835 ( .A(n18859), .ZN(P3_U3299) );
  INV_X1 U21836 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19735) );
  NAND2_X1 U21837 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19740), .ZN(n19729) );
  NAND2_X1 U21838 ( .A1(n19735), .A2(n19722), .ZN(n19726) );
  OAI21_X1 U21839 ( .B1(n19735), .B2(n19729), .A(n19726), .ZN(n19789) );
  AOI21_X1 U21840 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19789), .ZN(n18860) );
  INV_X1 U21841 ( .A(n18860), .ZN(P2_U2815) );
  AOI22_X1 U21842 ( .A1(n19841), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19792), 
        .B2(n19715), .ZN(n18861) );
  INV_X1 U21843 ( .A(n18861), .ZN(P2_U2816) );
  INV_X2 U21844 ( .A(n19859), .ZN(n19858) );
  AOI21_X1 U21845 ( .B1(n19735), .B2(n19740), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18862) );
  AOI22_X1 U21846 ( .A1(n19858), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18862), 
        .B2(n19859), .ZN(P2_U2817) );
  OAI21_X1 U21847 ( .B1(n19733), .B2(BS16), .A(n19789), .ZN(n19787) );
  OAI21_X1 U21848 ( .B1(n19789), .B2(n19791), .A(n19787), .ZN(P2_U2818) );
  NOR2_X1 U21849 ( .A1(n18864), .A2(n18863), .ZN(n19837) );
  OAI21_X1 U21850 ( .B1(n19837), .B2(n20817), .A(n18865), .ZN(P2_U2819) );
  NOR4_X1 U21851 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18869) );
  NOR4_X1 U21852 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18868) );
  NOR4_X1 U21853 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18867) );
  NOR4_X1 U21854 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18866) );
  NAND4_X1 U21855 ( .A1(n18869), .A2(n18868), .A3(n18867), .A4(n18866), .ZN(
        n18875) );
  NOR4_X1 U21856 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18873) );
  AOI211_X1 U21857 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_24__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18872) );
  NOR4_X1 U21858 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18871) );
  NOR4_X1 U21859 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18870) );
  NAND4_X1 U21860 ( .A1(n18873), .A2(n18872), .A3(n18871), .A4(n18870), .ZN(
        n18874) );
  NOR2_X1 U21861 ( .A1(n18875), .A2(n18874), .ZN(n18885) );
  INV_X1 U21862 ( .A(n18885), .ZN(n18883) );
  NOR2_X1 U21863 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18883), .ZN(n18878) );
  INV_X1 U21864 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18876) );
  AOI22_X1 U21865 ( .A1(n18878), .A2(n18988), .B1(n18883), .B2(n18876), .ZN(
        P2_U2820) );
  OR3_X1 U21866 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18882) );
  INV_X1 U21867 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18877) );
  AOI22_X1 U21868 ( .A1(n18878), .A2(n18882), .B1(n18883), .B2(n18877), .ZN(
        P2_U2821) );
  INV_X1 U21869 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19788) );
  NAND2_X1 U21870 ( .A1(n18878), .A2(n19788), .ZN(n18881) );
  OAI21_X1 U21871 ( .B1(n10272), .B2(n18988), .A(n18885), .ZN(n18879) );
  OAI21_X1 U21872 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18885), .A(n18879), 
        .ZN(n18880) );
  OAI221_X1 U21873 ( .B1(n18881), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18881), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18880), .ZN(P2_U2822) );
  INV_X1 U21874 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18884) );
  OAI221_X1 U21875 ( .B1(n18885), .B2(n18884), .C1(n18883), .C2(n18882), .A(
        n18881), .ZN(P2_U2823) );
  AOI211_X1 U21876 ( .C1(n18887), .C2(n18886), .A(n15888), .B(n19717), .ZN(
        n18891) );
  AOI22_X1 U21877 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n19000), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n18951), .ZN(n18888) );
  OAI21_X1 U21878 ( .B1(n18889), .B2(n18995), .A(n18888), .ZN(n18890) );
  AOI211_X1 U21879 ( .C1(P2_EBX_REG_21__SCAN_IN), .C2(n18992), .A(n18891), .B(
        n18890), .ZN(n18896) );
  INV_X1 U21880 ( .A(n18892), .ZN(n18894) );
  AOI22_X1 U21881 ( .A1(n18894), .A2(n18999), .B1(n18954), .B2(n18893), .ZN(
        n18895) );
  NAND2_X1 U21882 ( .A1(n18896), .A2(n18895), .ZN(P2_U2834) );
  INV_X1 U21883 ( .A(n18897), .ZN(n18898) );
  OAI22_X1 U21884 ( .A1(n18899), .A2(n18978), .B1(n18989), .B2(n18898), .ZN(
        n18900) );
  INV_X1 U21885 ( .A(n18900), .ZN(n18910) );
  AOI211_X1 U21886 ( .C1(n18903), .C2(n18901), .A(n18902), .B(n19717), .ZN(
        n18908) );
  INV_X1 U21887 ( .A(n18904), .ZN(n18906) );
  AOI22_X1 U21888 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19000), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n18951), .ZN(n18905) );
  OAI21_X1 U21889 ( .B1(n18906), .B2(n18995), .A(n18905), .ZN(n18907) );
  AOI211_X1 U21890 ( .C1(P2_EBX_REG_20__SCAN_IN), .C2(n18992), .A(n18908), .B(
        n18907), .ZN(n18909) );
  NAND2_X1 U21891 ( .A1(n18910), .A2(n18909), .ZN(P2_U2835) );
  OAI21_X1 U21892 ( .B1(n18912), .B2(n18911), .A(n18984), .ZN(n18920) );
  AOI22_X1 U21893 ( .A1(P2_EBX_REG_18__SCAN_IN), .A2(n18992), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19000), .ZN(n18913) );
  OAI21_X1 U21894 ( .B1(n18914), .B2(n18995), .A(n18913), .ZN(n18915) );
  AOI211_X1 U21895 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n18951), .A(n19113), 
        .B(n18915), .ZN(n18919) );
  AOI22_X1 U21896 ( .A1(n18917), .A2(n18999), .B1(n18954), .B2(n18916), .ZN(
        n18918) );
  OAI211_X1 U21897 ( .C1(n18921), .C2(n18920), .A(n18919), .B(n18918), .ZN(
        P2_U2837) );
  XNOR2_X1 U21898 ( .A(n18923), .B(n18922), .ZN(n18932) );
  AOI22_X1 U21899 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19000), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n18951), .ZN(n18924) );
  OAI21_X1 U21900 ( .B1(n18925), .B2(n18995), .A(n18924), .ZN(n18926) );
  AOI211_X1 U21901 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n18992), .A(n19113), .B(
        n18926), .ZN(n18931) );
  INV_X1 U21902 ( .A(n18927), .ZN(n18928) );
  AOI22_X1 U21903 ( .A1(n18929), .A2(n18999), .B1(n18954), .B2(n18928), .ZN(
        n18930) );
  OAI211_X1 U21904 ( .C1(n19717), .C2(n18932), .A(n18931), .B(n18930), .ZN(
        P2_U2838) );
  NOR2_X1 U21905 ( .A1(n9951), .A2(n18933), .ZN(n18935) );
  XOR2_X1 U21906 ( .A(n18935), .B(n18934), .Z(n18942) );
  AOI22_X1 U21907 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n19000), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n18951), .ZN(n18936) );
  OAI21_X1 U21908 ( .B1(n18937), .B2(n18995), .A(n18936), .ZN(n18938) );
  AOI211_X1 U21909 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n18992), .A(n19113), .B(
        n18938), .ZN(n18941) );
  AOI22_X1 U21910 ( .A1(n18939), .A2(n18999), .B1(n18954), .B2(n19012), .ZN(
        n18940) );
  OAI211_X1 U21911 ( .C1(n19717), .C2(n18942), .A(n18941), .B(n18940), .ZN(
        P2_U2839) );
  NOR2_X1 U21912 ( .A1(n9951), .A2(n18943), .ZN(n18946) );
  XOR2_X1 U21913 ( .A(n18946), .B(n18945), .Z(n18958) );
  INV_X1 U21914 ( .A(n18947), .ZN(n18949) );
  AOI22_X1 U21915 ( .A1(P2_EBX_REG_14__SCAN_IN), .A2(n18992), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19000), .ZN(n18948) );
  OAI21_X1 U21916 ( .B1(n18949), .B2(n18995), .A(n18948), .ZN(n18950) );
  AOI211_X1 U21917 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n18951), .A(n19113), 
        .B(n18950), .ZN(n18957) );
  INV_X1 U21918 ( .A(n18952), .ZN(n18955) );
  AOI22_X1 U21919 ( .A1(n18999), .A2(n18955), .B1(n18954), .B2(n18953), .ZN(
        n18956) );
  OAI211_X1 U21920 ( .C1(n19717), .C2(n18958), .A(n18957), .B(n18956), .ZN(
        P2_U2841) );
  NAND2_X1 U21921 ( .A1(n9949), .A2(n18959), .ZN(n18961) );
  XOR2_X1 U21922 ( .A(n18961), .B(n18960), .Z(n18968) );
  AOI22_X1 U21923 ( .A1(n18962), .A2(n13236), .B1(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19000), .ZN(n18963) );
  OAI211_X1 U21924 ( .C1(n11130), .C2(n18987), .A(n18963), .B(n15534), .ZN(
        n18966) );
  OAI22_X1 U21925 ( .A1(n18964), .A2(n18978), .B1(n18989), .B2(n19032), .ZN(
        n18965) );
  AOI211_X1 U21926 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n18992), .A(n18966), .B(
        n18965), .ZN(n18967) );
  OAI21_X1 U21927 ( .B1(n18968), .B2(n19717), .A(n18967), .ZN(P2_U2846) );
  NAND2_X1 U21928 ( .A1(n9949), .A2(n18969), .ZN(n18972) );
  XOR2_X1 U21929 ( .A(n18972), .B(n18971), .Z(n18983) );
  NOR2_X1 U21930 ( .A1(n18974), .A2(n18973), .ZN(n18975) );
  AOI21_X1 U21931 ( .B1(n18976), .B2(n13236), .A(n18975), .ZN(n18977) );
  OAI211_X1 U21932 ( .C1(n10797), .C2(n18987), .A(n18977), .B(n15534), .ZN(
        n18981) );
  OAI22_X1 U21933 ( .A1(n18979), .A2(n18978), .B1(n18989), .B2(n19037), .ZN(
        n18980) );
  AOI211_X1 U21934 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n18992), .A(n18981), .B(
        n18980), .ZN(n18982) );
  OAI21_X1 U21935 ( .B1(n18983), .B2(n19717), .A(n18982), .ZN(P2_U2848) );
  NOR2_X1 U21936 ( .A1(n18986), .A2(n18985), .ZN(n18997) );
  OAI22_X1 U21937 ( .A1(n18990), .A2(n18989), .B1(n18988), .B2(n18987), .ZN(
        n18991) );
  AOI21_X1 U21938 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n18992), .A(n18991), .ZN(
        n18993) );
  OAI21_X1 U21939 ( .B1(n18995), .B2(n18994), .A(n18993), .ZN(n18996) );
  AOI211_X1 U21940 ( .C1(n18999), .C2(n18998), .A(n18997), .B(n18996), .ZN(
        n19002) );
  NAND2_X1 U21941 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19000), .ZN(
        n19001) );
  OAI211_X1 U21942 ( .C1(n19003), .C2(n19717), .A(n19002), .B(n19001), .ZN(
        P2_U2855) );
  INV_X1 U21943 ( .A(n19004), .ZN(n19005) );
  AOI22_X1 U21944 ( .A1(n19005), .A2(n19056), .B1(n19010), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n19007) );
  AOI22_X1 U21945 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19055), .B1(n19011), 
        .B2(BUF2_REG_31__SCAN_IN), .ZN(n19006) );
  NAND2_X1 U21946 ( .A1(n19007), .A2(n19006), .ZN(P2_U2888) );
  AOI22_X1 U21947 ( .A1(n19009), .A2(n19008), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n19055), .ZN(n19016) );
  AOI22_X1 U21948 ( .A1(n19011), .A2(BUF2_REG_16__SCAN_IN), .B1(n19010), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19015) );
  AOI22_X1 U21949 ( .A1(n19013), .A2(n13149), .B1(n19056), .B2(n19012), .ZN(
        n19014) );
  NAND3_X1 U21950 ( .A1(n19016), .A2(n19015), .A3(n19014), .ZN(P2_U2903) );
  OAI222_X1 U21951 ( .A1(n19018), .A2(n19048), .B1(n13277), .B2(n19041), .C1(
        n19017), .C2(n19064), .ZN(P2_U2904) );
  AOI22_X1 U21952 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19055), .B1(n19106), 
        .B2(n19033), .ZN(n19019) );
  OAI21_X1 U21953 ( .B1(n19048), .B2(n19020), .A(n19019), .ZN(P2_U2905) );
  INV_X1 U21954 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19076) );
  OAI222_X1 U21955 ( .A1(n19022), .A2(n19048), .B1(n19076), .B2(n19041), .C1(
        n19064), .C2(n19021), .ZN(P2_U2906) );
  AOI22_X1 U21956 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19055), .B1(n19023), 
        .B2(n19033), .ZN(n19024) );
  OAI21_X1 U21957 ( .B1(n19048), .B2(n19025), .A(n19024), .ZN(P2_U2907) );
  INV_X1 U21958 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19080) );
  OAI222_X1 U21959 ( .A1(n19027), .A2(n19048), .B1(n19080), .B2(n19041), .C1(
        n19064), .C2(n19026), .ZN(P2_U2908) );
  AOI22_X1 U21960 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19055), .B1(n19028), 
        .B2(n19033), .ZN(n19029) );
  OAI21_X1 U21961 ( .B1(n19048), .B2(n19030), .A(n19029), .ZN(P2_U2909) );
  INV_X1 U21962 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19084) );
  OAI222_X1 U21963 ( .A1(n19032), .A2(n19048), .B1(n19084), .B2(n19041), .C1(
        n19064), .C2(n19031), .ZN(P2_U2910) );
  AOI22_X1 U21964 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19055), .B1(n19034), .B2(
        n19033), .ZN(n19035) );
  OAI21_X1 U21965 ( .B1(n19048), .B2(n19036), .A(n19035), .ZN(P2_U2911) );
  INV_X1 U21966 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19088) );
  OAI222_X1 U21967 ( .A1(n19037), .A2(n19048), .B1(n19088), .B2(n19041), .C1(
        n19064), .C2(n19169), .ZN(P2_U2912) );
  INV_X1 U21968 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19090) );
  OAI222_X1 U21969 ( .A1(n19039), .A2(n19048), .B1(n19090), .B2(n19041), .C1(
        n19064), .C2(n19038), .ZN(P2_U2913) );
  INV_X1 U21970 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19092) );
  OAI22_X1 U21971 ( .A1(n19092), .A2(n19041), .B1(n19040), .B2(n19064), .ZN(
        n19042) );
  INV_X1 U21972 ( .A(n19042), .ZN(n19046) );
  OR3_X1 U21973 ( .A1(n19044), .A2(n19043), .A3(n19060), .ZN(n19045) );
  OAI211_X1 U21974 ( .C1(n19048), .C2(n19047), .A(n19046), .B(n19045), .ZN(
        P2_U2914) );
  AOI22_X1 U21975 ( .A1(n19801), .A2(n19056), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19055), .ZN(n19054) );
  AOI21_X1 U21976 ( .B1(n19051), .B2(n19050), .A(n19049), .ZN(n19052) );
  OR2_X1 U21977 ( .A1(n19052), .A2(n19060), .ZN(n19053) );
  OAI211_X1 U21978 ( .C1(n19155), .C2(n19064), .A(n19054), .B(n19053), .ZN(
        P2_U2916) );
  AOI22_X1 U21979 ( .A1(n19056), .A2(n19820), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19055), .ZN(n19063) );
  AOI21_X1 U21980 ( .B1(n19059), .B2(n19058), .A(n19057), .ZN(n19061) );
  OR2_X1 U21981 ( .A1(n19061), .A2(n19060), .ZN(n19062) );
  OAI211_X1 U21982 ( .C1(n19065), .C2(n19064), .A(n19063), .B(n19062), .ZN(
        P2_U2918) );
  NOR2_X1 U21983 ( .A1(n19071), .A2(n19066), .ZN(P2_U2920) );
  INV_X1 U21984 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19070) );
  INV_X1 U21985 ( .A(n19067), .ZN(n19068) );
  AOI22_X1 U21986 ( .A1(n19068), .A2(P2_EAX_REG_30__SCAN_IN), .B1(
        P2_UWORD_REG_14__SCAN_IN), .B2(n19099), .ZN(n19069) );
  OAI21_X1 U21987 ( .B1(n19071), .B2(n19070), .A(n19069), .ZN(P2_U2921) );
  AOI22_X1 U21988 ( .A1(n19099), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19072) );
  OAI21_X1 U21989 ( .B1(n13277), .B2(n19104), .A(n19072), .ZN(P2_U2936) );
  INV_X1 U21990 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19074) );
  AOI22_X1 U21991 ( .A1(n19099), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19073) );
  OAI21_X1 U21992 ( .B1(n19074), .B2(n19104), .A(n19073), .ZN(P2_U2937) );
  AOI22_X1 U21993 ( .A1(n19099), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19075) );
  OAI21_X1 U21994 ( .B1(n19076), .B2(n19104), .A(n19075), .ZN(P2_U2938) );
  AOI22_X1 U21995 ( .A1(n19099), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19077) );
  OAI21_X1 U21996 ( .B1(n19078), .B2(n19104), .A(n19077), .ZN(P2_U2939) );
  AOI22_X1 U21997 ( .A1(n19099), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19079) );
  OAI21_X1 U21998 ( .B1(n19080), .B2(n19104), .A(n19079), .ZN(P2_U2940) );
  AOI22_X1 U21999 ( .A1(n19099), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19081) );
  OAI21_X1 U22000 ( .B1(n19082), .B2(n19104), .A(n19081), .ZN(P2_U2941) );
  AOI22_X1 U22001 ( .A1(n19099), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19083) );
  OAI21_X1 U22002 ( .B1(n19084), .B2(n19104), .A(n19083), .ZN(P2_U2942) );
  AOI22_X1 U22003 ( .A1(n19099), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19085) );
  OAI21_X1 U22004 ( .B1(n19086), .B2(n19104), .A(n19085), .ZN(P2_U2943) );
  AOI22_X1 U22005 ( .A1(n19099), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19087) );
  OAI21_X1 U22006 ( .B1(n19088), .B2(n19104), .A(n19087), .ZN(P2_U2944) );
  AOI22_X1 U22007 ( .A1(n19099), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19089) );
  OAI21_X1 U22008 ( .B1(n19090), .B2(n19104), .A(n19089), .ZN(P2_U2945) );
  AOI22_X1 U22009 ( .A1(n19099), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19091) );
  OAI21_X1 U22010 ( .B1(n19092), .B2(n19104), .A(n19091), .ZN(P2_U2946) );
  INV_X1 U22011 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19094) );
  AOI22_X1 U22012 ( .A1(n19099), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19093) );
  OAI21_X1 U22013 ( .B1(n19094), .B2(n19104), .A(n19093), .ZN(P2_U2947) );
  INV_X1 U22014 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19096) );
  AOI22_X1 U22015 ( .A1(n19099), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19095) );
  OAI21_X1 U22016 ( .B1(n19096), .B2(n19104), .A(n19095), .ZN(P2_U2948) );
  INV_X1 U22017 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19098) );
  AOI22_X1 U22018 ( .A1(n19099), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19097) );
  OAI21_X1 U22019 ( .B1(n19098), .B2(n19104), .A(n19097), .ZN(P2_U2949) );
  INV_X1 U22020 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19101) );
  AOI22_X1 U22021 ( .A1(n19099), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19100) );
  OAI21_X1 U22022 ( .B1(n19101), .B2(n19104), .A(n19100), .ZN(P2_U2950) );
  INV_X1 U22023 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19105) );
  AOI22_X1 U22024 ( .A1(n19099), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19102), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19103) );
  OAI21_X1 U22025 ( .B1(n19105), .B2(n19104), .A(n19103), .ZN(P2_U2951) );
  AOI22_X1 U22026 ( .A1(n19110), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n19109), .ZN(n19108) );
  NAND2_X1 U22027 ( .A1(n19107), .A2(n19106), .ZN(n19111) );
  NAND2_X1 U22028 ( .A1(n19108), .A2(n19111), .ZN(P2_U2966) );
  AOI22_X1 U22029 ( .A1(n19110), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19109), 
        .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n19112) );
  NAND2_X1 U22030 ( .A1(n19112), .A2(n19111), .ZN(P2_U2981) );
  AOI22_X1 U22031 ( .A1(n19114), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19113), .ZN(n19123) );
  INV_X1 U22032 ( .A(n19115), .ZN(n19116) );
  AOI222_X1 U22033 ( .A1(n19121), .A2(n19120), .B1(n19119), .B2(n19118), .C1(
        n19117), .C2(n19116), .ZN(n19122) );
  OAI211_X1 U22034 ( .C1(n19125), .C2(n19124), .A(n19123), .B(n19122), .ZN(
        P2_U3010) );
  NOR2_X1 U22035 ( .A1(n19127), .A2(n19126), .ZN(n19148) );
  INV_X1 U22036 ( .A(n19128), .ZN(n19129) );
  NAND2_X1 U22037 ( .A1(n19129), .A2(n19148), .ZN(n19132) );
  NAND2_X1 U22038 ( .A1(n19130), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19131) );
  OAI211_X1 U22039 ( .C1(n19134), .C2(n19133), .A(n19132), .B(n19131), .ZN(
        n19135) );
  INV_X1 U22040 ( .A(n19135), .ZN(n19142) );
  OAI22_X1 U22041 ( .A1(n19139), .A2(n19138), .B1(n19137), .B2(n19136), .ZN(
        n19140) );
  INV_X1 U22042 ( .A(n19140), .ZN(n19141) );
  OAI211_X1 U22043 ( .C1(n19806), .C2(n19143), .A(n19142), .B(n19141), .ZN(
        n19144) );
  INV_X1 U22044 ( .A(n19144), .ZN(n19146) );
  OAI211_X1 U22045 ( .C1(n19148), .C2(n19147), .A(n19146), .B(n19145), .ZN(
        P2_U3044) );
  AOI22_X1 U22046 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19171), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19170), .ZN(n19678) );
  INV_X1 U22047 ( .A(n19678), .ZN(n19507) );
  AOI22_X1 U22048 ( .A1(n19507), .A2(n19708), .B1(n19168), .B2(n19674), .ZN(
        n19153) );
  AOI22_X1 U22049 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19171), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19170), .ZN(n19510) );
  INV_X1 U22050 ( .A(n19510), .ZN(n19675) );
  AOI22_X1 U22051 ( .A1(n19151), .A2(n19172), .B1(n19200), .B2(n19675), .ZN(
        n19152) );
  OAI211_X1 U22052 ( .C1(n19176), .C2(n12863), .A(n19153), .B(n19152), .ZN(
        P2_U3050) );
  INV_X1 U22053 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19158) );
  AOI22_X1 U22054 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19171), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19170), .ZN(n19684) );
  NOR2_X2 U22055 ( .A1(n19154), .A2(n19166), .ZN(n19679) );
  AOI22_X1 U22056 ( .A1(n19632), .A2(n19708), .B1(n19168), .B2(n19679), .ZN(
        n19157) );
  NOR2_X2 U22057 ( .A1(n19155), .A2(n19363), .ZN(n19680) );
  AOI22_X1 U22058 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19171), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19170), .ZN(n19635) );
  INV_X1 U22059 ( .A(n19635), .ZN(n19681) );
  AOI22_X1 U22060 ( .A1(n19680), .A2(n19172), .B1(n19200), .B2(n19681), .ZN(
        n19156) );
  OAI211_X1 U22061 ( .C1(n19176), .C2(n19158), .A(n19157), .B(n19156), .ZN(
        P2_U3051) );
  AOI22_X1 U22062 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19171), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19170), .ZN(n19690) );
  NOR2_X2 U22063 ( .A1(n10251), .A2(n19166), .ZN(n19685) );
  AOI22_X1 U22064 ( .A1(n19636), .A2(n19708), .B1(n19168), .B2(n19685), .ZN(
        n19161) );
  NOR2_X2 U22065 ( .A1(n19159), .A2(n19363), .ZN(n19686) );
  AOI22_X1 U22066 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19171), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19170), .ZN(n19639) );
  INV_X1 U22067 ( .A(n19639), .ZN(n19687) );
  AOI22_X1 U22068 ( .A1(n19686), .A2(n19172), .B1(n19200), .B2(n19687), .ZN(
        n19160) );
  OAI211_X1 U22069 ( .C1(n19176), .C2(n12883), .A(n19161), .B(n19160), .ZN(
        P2_U3052) );
  INV_X1 U22070 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19175) );
  NOR2_X2 U22071 ( .A1(n19167), .A2(n19166), .ZN(n19704) );
  AOI22_X1 U22072 ( .A1(n19650), .A2(n19708), .B1(n19168), .B2(n19704), .ZN(
        n19174) );
  NOR2_X2 U22073 ( .A1(n19169), .A2(n19363), .ZN(n19705) );
  AOI22_X1 U22074 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19171), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19170), .ZN(n19655) );
  AOI22_X1 U22075 ( .A1(n19705), .A2(n19172), .B1(n19200), .B2(n19707), .ZN(
        n19173) );
  OAI211_X1 U22076 ( .C1(n19176), .C2(n19175), .A(n19174), .B(n19173), .ZN(
        P2_U3055) );
  INV_X1 U22077 ( .A(n19793), .ZN(n19797) );
  NAND2_X1 U22078 ( .A1(n19822), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19421) );
  NOR2_X1 U22079 ( .A1(n19421), .A2(n19233), .ZN(n19198) );
  OAI21_X1 U22080 ( .B1(n19179), .B2(n19198), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19177) );
  OAI21_X1 U22081 ( .B1(n19178), .B2(n19797), .A(n19177), .ZN(n19199) );
  AOI22_X1 U22082 ( .A1(n19199), .A2(n14284), .B1(n19657), .B2(n19198), .ZN(
        n19185) );
  NAND2_X1 U22083 ( .A1(n19795), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19798) );
  OAI21_X1 U22084 ( .B1(n19798), .B2(n19420), .A(n19178), .ZN(n19183) );
  INV_X1 U22085 ( .A(n19179), .ZN(n19181) );
  INV_X1 U22086 ( .A(n19198), .ZN(n19180) );
  OAI211_X1 U22087 ( .C1(n19181), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19180), 
        .B(n19797), .ZN(n19182) );
  NAND3_X1 U22088 ( .A1(n19183), .A2(n19662), .A3(n19182), .ZN(n19201) );
  AOI22_X1 U22089 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19201), .B1(
        n19200), .B2(n19613), .ZN(n19184) );
  OAI211_X1 U22090 ( .C1(n19625), .C2(n19218), .A(n19185), .B(n19184), .ZN(
        P2_U3056) );
  AOI22_X1 U22091 ( .A1(n19199), .A2(n14299), .B1(n19669), .B2(n19198), .ZN(
        n19187) );
  AOI22_X1 U22092 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19201), .B1(
        n19200), .B2(n19626), .ZN(n19186) );
  OAI211_X1 U22093 ( .C1(n19629), .C2(n19218), .A(n19187), .B(n19186), .ZN(
        P2_U3057) );
  AOI22_X1 U22094 ( .A1(n19199), .A2(n19151), .B1(n19674), .B2(n19198), .ZN(
        n19189) );
  AOI22_X1 U22095 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19201), .B1(
        n19200), .B2(n19507), .ZN(n19188) );
  OAI211_X1 U22096 ( .C1(n19510), .C2(n19218), .A(n19189), .B(n19188), .ZN(
        P2_U3058) );
  AOI22_X1 U22097 ( .A1(n19199), .A2(n19680), .B1(n19679), .B2(n19198), .ZN(
        n19191) );
  AOI22_X1 U22098 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19201), .B1(
        n19200), .B2(n19632), .ZN(n19190) );
  OAI211_X1 U22099 ( .C1(n19635), .C2(n19218), .A(n19191), .B(n19190), .ZN(
        P2_U3059) );
  AOI22_X1 U22100 ( .A1(n19199), .A2(n19686), .B1(n19685), .B2(n19198), .ZN(
        n19193) );
  AOI22_X1 U22101 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19201), .B1(
        n19200), .B2(n19636), .ZN(n19192) );
  OAI211_X1 U22102 ( .C1(n19639), .C2(n19218), .A(n19193), .B(n19192), .ZN(
        P2_U3060) );
  AOI22_X1 U22103 ( .A1(n19199), .A2(n19692), .B1(n19691), .B2(n19198), .ZN(
        n19195) );
  AOI22_X1 U22104 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19201), .B1(
        n19200), .B2(n19640), .ZN(n19194) );
  OAI211_X1 U22105 ( .C1(n19643), .C2(n19218), .A(n19195), .B(n19194), .ZN(
        P2_U3061) );
  AOI22_X1 U22106 ( .A1(n19199), .A2(n19698), .B1(n19697), .B2(n19198), .ZN(
        n19197) );
  AOI22_X1 U22107 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19201), .B1(
        n19200), .B2(n19600), .ZN(n19196) );
  OAI211_X1 U22108 ( .C1(n19604), .C2(n19218), .A(n19197), .B(n19196), .ZN(
        P2_U3062) );
  AOI22_X1 U22109 ( .A1(n19199), .A2(n19705), .B1(n19704), .B2(n19198), .ZN(
        n19203) );
  AOI22_X1 U22110 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19201), .B1(
        n19200), .B2(n19650), .ZN(n19202) );
  OAI211_X1 U22111 ( .C1(n19655), .C2(n19218), .A(n19203), .B(n19202), .ZN(
        P2_U3063) );
  NOR2_X1 U22112 ( .A1(n19822), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19451) );
  AND2_X1 U22113 ( .A1(n19451), .A2(n19234), .ZN(n19227) );
  OAI21_X1 U22114 ( .B1(n10481), .B2(n19227), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19204) );
  NAND2_X1 U22115 ( .A1(n19450), .A2(n19234), .ZN(n19205) );
  NAND2_X1 U22116 ( .A1(n19204), .A2(n19205), .ZN(n19228) );
  AOI22_X1 U22117 ( .A1(n19228), .A2(n14284), .B1(n19657), .B2(n19227), .ZN(
        n19213) );
  OAI21_X1 U22118 ( .B1(n19249), .B2(n19229), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19206) );
  NAND2_X1 U22119 ( .A1(n19206), .A2(n19205), .ZN(n19210) );
  INV_X1 U22120 ( .A(n10481), .ZN(n19208) );
  INV_X1 U22121 ( .A(n19227), .ZN(n19207) );
  OAI21_X1 U22122 ( .B1(n19208), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19207), 
        .ZN(n19209) );
  MUX2_X1 U22123 ( .A(n19210), .B(n19209), .S(n19797), .Z(n19211) );
  NAND2_X1 U22124 ( .A1(n19211), .A2(n19662), .ZN(n19230) );
  AOI22_X1 U22125 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19230), .B1(
        n19249), .B2(n19665), .ZN(n19212) );
  OAI211_X1 U22126 ( .C1(n19668), .C2(n19218), .A(n19213), .B(n19212), .ZN(
        P2_U3064) );
  AOI22_X1 U22127 ( .A1(n19228), .A2(n14299), .B1(n19669), .B2(n19227), .ZN(
        n19215) );
  AOI22_X1 U22128 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19230), .B1(
        n19249), .B2(n19670), .ZN(n19214) );
  OAI211_X1 U22129 ( .C1(n19673), .C2(n19218), .A(n19215), .B(n19214), .ZN(
        P2_U3065) );
  AOI22_X1 U22130 ( .A1(n19228), .A2(n19151), .B1(n19674), .B2(n19227), .ZN(
        n19217) );
  AOI22_X1 U22131 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19230), .B1(
        n19249), .B2(n19675), .ZN(n19216) );
  OAI211_X1 U22132 ( .C1(n19678), .C2(n19218), .A(n19217), .B(n19216), .ZN(
        P2_U3066) );
  AOI22_X1 U22133 ( .A1(n19228), .A2(n19680), .B1(n19679), .B2(n19227), .ZN(
        n19220) );
  AOI22_X1 U22134 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19230), .B1(
        n19229), .B2(n19632), .ZN(n19219) );
  OAI211_X1 U22135 ( .C1(n19635), .C2(n19263), .A(n19220), .B(n19219), .ZN(
        P2_U3067) );
  AOI22_X1 U22136 ( .A1(n19228), .A2(n19686), .B1(n19685), .B2(n19227), .ZN(
        n19222) );
  AOI22_X1 U22137 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19230), .B1(
        n19229), .B2(n19636), .ZN(n19221) );
  OAI211_X1 U22138 ( .C1(n19639), .C2(n19263), .A(n19222), .B(n19221), .ZN(
        P2_U3068) );
  AOI22_X1 U22139 ( .A1(n19228), .A2(n19692), .B1(n19691), .B2(n19227), .ZN(
        n19224) );
  AOI22_X1 U22140 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19230), .B1(
        n19229), .B2(n19640), .ZN(n19223) );
  OAI211_X1 U22141 ( .C1(n19643), .C2(n19263), .A(n19224), .B(n19223), .ZN(
        P2_U3069) );
  AOI22_X1 U22142 ( .A1(n19228), .A2(n19698), .B1(n19697), .B2(n19227), .ZN(
        n19226) );
  AOI22_X1 U22143 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19230), .B1(
        n19229), .B2(n19600), .ZN(n19225) );
  OAI211_X1 U22144 ( .C1(n19604), .C2(n19263), .A(n19226), .B(n19225), .ZN(
        P2_U3070) );
  AOI22_X1 U22145 ( .A1(n19228), .A2(n19705), .B1(n19704), .B2(n19227), .ZN(
        n19232) );
  AOI22_X1 U22146 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19230), .B1(
        n19229), .B2(n19650), .ZN(n19231) );
  OAI211_X1 U22147 ( .C1(n19655), .C2(n19263), .A(n19232), .B(n19231), .ZN(
        P2_U3071) );
  NOR2_X1 U22148 ( .A1(n19482), .A2(n19233), .ZN(n19258) );
  AOI22_X1 U22149 ( .A1(n19613), .A2(n19249), .B1(n19657), .B2(n19258), .ZN(
        n19244) );
  OAI21_X1 U22150 ( .B1(n19798), .B2(n19481), .A(n19793), .ZN(n19242) );
  NAND2_X1 U22151 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19234), .ZN(
        n19241) );
  INV_X1 U22152 ( .A(n19241), .ZN(n19238) );
  INV_X1 U22153 ( .A(n19239), .ZN(n19236) );
  INV_X1 U22154 ( .A(n19258), .ZN(n19235) );
  OAI211_X1 U22155 ( .C1(n19236), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19235), 
        .B(n19797), .ZN(n19237) );
  OAI211_X1 U22156 ( .C1(n19242), .C2(n19238), .A(n19662), .B(n19237), .ZN(
        n19260) );
  OAI21_X1 U22157 ( .B1(n19239), .B2(n19258), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19240) );
  OAI21_X1 U22158 ( .B1(n19242), .B2(n19241), .A(n19240), .ZN(n19259) );
  AOI22_X1 U22159 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19260), .B1(
        n14284), .B2(n19259), .ZN(n19243) );
  OAI211_X1 U22160 ( .C1(n19625), .C2(n19294), .A(n19244), .B(n19243), .ZN(
        P2_U3072) );
  AOI22_X1 U22161 ( .A1(n19670), .A2(n19286), .B1(n19669), .B2(n19258), .ZN(
        n19246) );
  AOI22_X1 U22162 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19260), .B1(
        n14299), .B2(n19259), .ZN(n19245) );
  OAI211_X1 U22163 ( .C1(n19673), .C2(n19263), .A(n19246), .B(n19245), .ZN(
        P2_U3073) );
  AOI22_X1 U22164 ( .A1(n19675), .A2(n19286), .B1(n19258), .B2(n19674), .ZN(
        n19248) );
  AOI22_X1 U22165 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19260), .B1(
        n19151), .B2(n19259), .ZN(n19247) );
  OAI211_X1 U22166 ( .C1(n19678), .C2(n19263), .A(n19248), .B(n19247), .ZN(
        P2_U3074) );
  AOI22_X1 U22167 ( .A1(n19632), .A2(n19249), .B1(n19258), .B2(n19679), .ZN(
        n19251) );
  AOI22_X1 U22168 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19260), .B1(
        n19680), .B2(n19259), .ZN(n19250) );
  OAI211_X1 U22169 ( .C1(n19635), .C2(n19294), .A(n19251), .B(n19250), .ZN(
        P2_U3075) );
  AOI22_X1 U22170 ( .A1(n19687), .A2(n19286), .B1(n19258), .B2(n19685), .ZN(
        n19253) );
  AOI22_X1 U22171 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19260), .B1(
        n19686), .B2(n19259), .ZN(n19252) );
  OAI211_X1 U22172 ( .C1(n19690), .C2(n19263), .A(n19253), .B(n19252), .ZN(
        P2_U3076) );
  AOI22_X1 U22173 ( .A1(n19693), .A2(n19286), .B1(n19691), .B2(n19258), .ZN(
        n19255) );
  AOI22_X1 U22174 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19260), .B1(
        n19692), .B2(n19259), .ZN(n19254) );
  OAI211_X1 U22175 ( .C1(n19696), .C2(n19263), .A(n19255), .B(n19254), .ZN(
        P2_U3077) );
  AOI22_X1 U22176 ( .A1(n19699), .A2(n19286), .B1(n19697), .B2(n19258), .ZN(
        n19257) );
  AOI22_X1 U22177 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19260), .B1(
        n19698), .B2(n19259), .ZN(n19256) );
  OAI211_X1 U22178 ( .C1(n19702), .C2(n19263), .A(n19257), .B(n19256), .ZN(
        P2_U3078) );
  AOI22_X1 U22179 ( .A1(n19707), .A2(n19286), .B1(n19258), .B2(n19704), .ZN(
        n19262) );
  AOI22_X1 U22180 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19260), .B1(
        n19705), .B2(n19259), .ZN(n19261) );
  OAI211_X1 U22181 ( .C1(n19713), .C2(n19263), .A(n19262), .B(n19261), .ZN(
        P2_U3079) );
  INV_X1 U22182 ( .A(n19264), .ZN(n19266) );
  NOR2_X1 U22183 ( .A1(n19266), .A2(n19265), .ZN(n19550) );
  NAND2_X1 U22184 ( .A1(n19550), .A2(n19803), .ZN(n19272) );
  NAND3_X1 U22185 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19803), .A3(
        n19822), .ZN(n19302) );
  NOR2_X1 U22186 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19302), .ZN(
        n19289) );
  OAI21_X1 U22187 ( .B1(n19269), .B2(n19289), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19267) );
  OAI21_X1 U22188 ( .B1(n19272), .B2(n19797), .A(n19267), .ZN(n19290) );
  AOI22_X1 U22189 ( .A1(n19290), .A2(n14284), .B1(n19657), .B2(n19289), .ZN(
        n19275) );
  NOR2_X2 U22190 ( .A1(n19583), .A2(n19327), .ZN(n19321) );
  OAI21_X1 U22191 ( .B1(n19286), .B2(n19321), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19271) );
  AOI211_X1 U22192 ( .C1(n19269), .C2(n19839), .A(n19289), .B(n19793), .ZN(
        n19270) );
  AOI211_X1 U22193 ( .C1(n19272), .C2(n19271), .A(n19363), .B(n19270), .ZN(
        n19273) );
  AOI22_X1 U22194 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19291), .B1(
        n19321), .B2(n19665), .ZN(n19274) );
  OAI211_X1 U22195 ( .C1(n19668), .C2(n19294), .A(n19275), .B(n19274), .ZN(
        P2_U3080) );
  AOI22_X1 U22196 ( .A1(n19290), .A2(n14299), .B1(n19669), .B2(n19289), .ZN(
        n19277) );
  AOI22_X1 U22197 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19291), .B1(
        n19321), .B2(n19670), .ZN(n19276) );
  OAI211_X1 U22198 ( .C1(n19673), .C2(n19294), .A(n19277), .B(n19276), .ZN(
        P2_U3081) );
  INV_X1 U22199 ( .A(n19321), .ZN(n19318) );
  AOI22_X1 U22200 ( .A1(n19290), .A2(n19151), .B1(n19674), .B2(n19289), .ZN(
        n19279) );
  AOI22_X1 U22201 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19291), .B1(
        n19286), .B2(n19507), .ZN(n19278) );
  OAI211_X1 U22202 ( .C1(n19510), .C2(n19318), .A(n19279), .B(n19278), .ZN(
        P2_U3082) );
  AOI22_X1 U22203 ( .A1(n19290), .A2(n19680), .B1(n19679), .B2(n19289), .ZN(
        n19281) );
  AOI22_X1 U22204 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19291), .B1(
        n19286), .B2(n19632), .ZN(n19280) );
  OAI211_X1 U22205 ( .C1(n19635), .C2(n19318), .A(n19281), .B(n19280), .ZN(
        P2_U3083) );
  AOI22_X1 U22206 ( .A1(n19290), .A2(n19686), .B1(n19685), .B2(n19289), .ZN(
        n19283) );
  AOI22_X1 U22207 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19291), .B1(
        n19321), .B2(n19687), .ZN(n19282) );
  OAI211_X1 U22208 ( .C1(n19690), .C2(n19294), .A(n19283), .B(n19282), .ZN(
        P2_U3084) );
  AOI22_X1 U22209 ( .A1(n19290), .A2(n19692), .B1(n19691), .B2(n19289), .ZN(
        n19285) );
  AOI22_X1 U22210 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19291), .B1(
        n19321), .B2(n19693), .ZN(n19284) );
  OAI211_X1 U22211 ( .C1(n19696), .C2(n19294), .A(n19285), .B(n19284), .ZN(
        P2_U3085) );
  AOI22_X1 U22212 ( .A1(n19290), .A2(n19698), .B1(n19697), .B2(n19289), .ZN(
        n19288) );
  AOI22_X1 U22213 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19291), .B1(
        n19286), .B2(n19600), .ZN(n19287) );
  OAI211_X1 U22214 ( .C1(n19604), .C2(n19318), .A(n19288), .B(n19287), .ZN(
        P2_U3086) );
  AOI22_X1 U22215 ( .A1(n19290), .A2(n19705), .B1(n19704), .B2(n19289), .ZN(
        n19293) );
  AOI22_X1 U22216 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19291), .B1(
        n19321), .B2(n19707), .ZN(n19292) );
  OAI211_X1 U22217 ( .C1(n19713), .C2(n19294), .A(n19293), .B(n19292), .ZN(
        P2_U3087) );
  OAI21_X1 U22218 ( .B1(n19798), .B2(n19583), .A(n19793), .ZN(n19303) );
  INV_X1 U22219 ( .A(n19302), .ZN(n19295) );
  OR2_X1 U22220 ( .A1(n19303), .A2(n19295), .ZN(n19299) );
  NAND2_X1 U22221 ( .A1(n19300), .A2(n19839), .ZN(n19297) );
  NOR2_X1 U22222 ( .A1(n19828), .A2(n19302), .ZN(n19329) );
  NOR2_X1 U22223 ( .A1(n19793), .A2(n19329), .ZN(n19296) );
  AOI21_X1 U22224 ( .B1(n19297), .B2(n19296), .A(n19363), .ZN(n19298) );
  INV_X1 U22225 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n19306) );
  AOI22_X1 U22226 ( .A1(n19613), .A2(n19321), .B1(n19657), .B2(n19329), .ZN(
        n19305) );
  OAI21_X1 U22227 ( .B1(n19300), .B2(n19329), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19301) );
  OAI21_X1 U22228 ( .B1(n19303), .B2(n19302), .A(n19301), .ZN(n19322) );
  NOR2_X2 U22229 ( .A1(n19367), .A2(n19583), .ZN(n19354) );
  AOI22_X1 U22230 ( .A1(n14284), .A2(n19322), .B1(n19354), .B2(n19665), .ZN(
        n19304) );
  OAI211_X1 U22231 ( .C1(n19309), .C2(n19306), .A(n19305), .B(n19304), .ZN(
        P2_U3088) );
  AOI22_X1 U22232 ( .A1(n19670), .A2(n19354), .B1(n19669), .B2(n19329), .ZN(
        n19308) );
  AOI22_X1 U22233 ( .A1(n14299), .A2(n19322), .B1(n19321), .B2(n19626), .ZN(
        n19307) );
  OAI211_X1 U22234 ( .C1(n19309), .C2(n10386), .A(n19308), .B(n19307), .ZN(
        P2_U3089) );
  AOI22_X1 U22235 ( .A1(n19675), .A2(n19354), .B1(n19674), .B2(n19329), .ZN(
        n19311) );
  AOI22_X1 U22236 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19323), .B1(
        n19151), .B2(n19322), .ZN(n19310) );
  OAI211_X1 U22237 ( .C1(n19678), .C2(n19318), .A(n19311), .B(n19310), .ZN(
        P2_U3090) );
  INV_X1 U22238 ( .A(n19354), .ZN(n19326) );
  AOI22_X1 U22239 ( .A1(n19632), .A2(n19321), .B1(n19329), .B2(n19679), .ZN(
        n19313) );
  AOI22_X1 U22240 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19323), .B1(
        n19680), .B2(n19322), .ZN(n19312) );
  OAI211_X1 U22241 ( .C1(n19635), .C2(n19326), .A(n19313), .B(n19312), .ZN(
        P2_U3091) );
  AOI22_X1 U22242 ( .A1(n19636), .A2(n19321), .B1(n19685), .B2(n19329), .ZN(
        n19315) );
  AOI22_X1 U22243 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19323), .B1(
        n19686), .B2(n19322), .ZN(n19314) );
  OAI211_X1 U22244 ( .C1(n19639), .C2(n19326), .A(n19315), .B(n19314), .ZN(
        P2_U3092) );
  AOI22_X1 U22245 ( .A1(n19693), .A2(n19354), .B1(n19691), .B2(n19329), .ZN(
        n19317) );
  AOI22_X1 U22246 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19323), .B1(
        n19692), .B2(n19322), .ZN(n19316) );
  OAI211_X1 U22247 ( .C1(n19696), .C2(n19318), .A(n19317), .B(n19316), .ZN(
        P2_U3093) );
  AOI22_X1 U22248 ( .A1(n19600), .A2(n19321), .B1(n19697), .B2(n19329), .ZN(
        n19320) );
  AOI22_X1 U22249 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19323), .B1(
        n19698), .B2(n19322), .ZN(n19319) );
  OAI211_X1 U22250 ( .C1(n19604), .C2(n19326), .A(n19320), .B(n19319), .ZN(
        P2_U3094) );
  AOI22_X1 U22251 ( .A1(n19650), .A2(n19321), .B1(n19704), .B2(n19329), .ZN(
        n19325) );
  AOI22_X1 U22252 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19323), .B1(
        n19705), .B2(n19322), .ZN(n19324) );
  OAI211_X1 U22253 ( .C1(n19655), .C2(n19326), .A(n19325), .B(n19324), .ZN(
        P2_U3095) );
  NOR2_X1 U22254 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19328), .ZN(
        n19352) );
  NOR2_X1 U22255 ( .A1(n19329), .A2(n19352), .ZN(n19335) );
  INV_X1 U22256 ( .A(n19330), .ZN(n19333) );
  OAI21_X1 U22257 ( .B1(n19333), .B2(n19352), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19331) );
  OAI21_X1 U22258 ( .B1(n19335), .B2(n19797), .A(n19331), .ZN(n19353) );
  AOI22_X1 U22259 ( .A1(n19353), .A2(n14284), .B1(n19657), .B2(n19352), .ZN(
        n19339) );
  OAI21_X1 U22260 ( .B1(n19354), .B2(n19332), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19336) );
  AOI211_X1 U22261 ( .C1(n19333), .C2(n19839), .A(n19352), .B(n19793), .ZN(
        n19334) );
  AOI211_X1 U22262 ( .C1(n19336), .C2(n19335), .A(n19334), .B(n19363), .ZN(
        n19337) );
  AOI22_X1 U22263 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19355), .B1(
        n19354), .B2(n19613), .ZN(n19338) );
  OAI211_X1 U22264 ( .C1(n19625), .C2(n19389), .A(n19339), .B(n19338), .ZN(
        P2_U3096) );
  AOI22_X1 U22265 ( .A1(n19353), .A2(n14299), .B1(n19669), .B2(n19352), .ZN(
        n19341) );
  AOI22_X1 U22266 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19355), .B1(
        n19354), .B2(n19626), .ZN(n19340) );
  OAI211_X1 U22267 ( .C1(n19629), .C2(n19389), .A(n19341), .B(n19340), .ZN(
        P2_U3097) );
  AOI22_X1 U22268 ( .A1(n19353), .A2(n19151), .B1(n19674), .B2(n19352), .ZN(
        n19343) );
  AOI22_X1 U22269 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19355), .B1(
        n19354), .B2(n19507), .ZN(n19342) );
  OAI211_X1 U22270 ( .C1(n19510), .C2(n19389), .A(n19343), .B(n19342), .ZN(
        P2_U3098) );
  AOI22_X1 U22271 ( .A1(n19353), .A2(n19680), .B1(n19679), .B2(n19352), .ZN(
        n19345) );
  AOI22_X1 U22272 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19355), .B1(
        n19354), .B2(n19632), .ZN(n19344) );
  OAI211_X1 U22273 ( .C1(n19635), .C2(n19389), .A(n19345), .B(n19344), .ZN(
        P2_U3099) );
  AOI22_X1 U22274 ( .A1(n19353), .A2(n19686), .B1(n19685), .B2(n19352), .ZN(
        n19347) );
  AOI22_X1 U22275 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19355), .B1(
        n19354), .B2(n19636), .ZN(n19346) );
  OAI211_X1 U22276 ( .C1(n19639), .C2(n19389), .A(n19347), .B(n19346), .ZN(
        P2_U3100) );
  AOI22_X1 U22277 ( .A1(n19353), .A2(n19692), .B1(n19691), .B2(n19352), .ZN(
        n19349) );
  AOI22_X1 U22278 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19355), .B1(
        n19354), .B2(n19640), .ZN(n19348) );
  OAI211_X1 U22279 ( .C1(n19643), .C2(n19389), .A(n19349), .B(n19348), .ZN(
        P2_U3101) );
  AOI22_X1 U22280 ( .A1(n19353), .A2(n19698), .B1(n19697), .B2(n19352), .ZN(
        n19351) );
  AOI22_X1 U22281 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19355), .B1(
        n19354), .B2(n19600), .ZN(n19350) );
  OAI211_X1 U22282 ( .C1(n19604), .C2(n19389), .A(n19351), .B(n19350), .ZN(
        P2_U3102) );
  AOI22_X1 U22283 ( .A1(n19353), .A2(n19705), .B1(n19704), .B2(n19352), .ZN(
        n19357) );
  AOI22_X1 U22284 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19355), .B1(
        n19354), .B2(n19650), .ZN(n19356) );
  OAI211_X1 U22285 ( .C1(n19655), .C2(n19389), .A(n19357), .B(n19356), .ZN(
        P2_U3103) );
  NOR2_X1 U22286 ( .A1(n19395), .A2(n19848), .ZN(n19358) );
  AOI21_X1 U22287 ( .B1(n19839), .B2(n19361), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19360) );
  NOR2_X1 U22288 ( .A1(n19364), .A2(n19360), .ZN(n19385) );
  AOI22_X1 U22289 ( .A1(n19385), .A2(n14284), .B1(n19395), .B2(n19657), .ZN(
        n19369) );
  INV_X1 U22290 ( .A(n19798), .ZN(n19362) );
  AOI21_X1 U22291 ( .B1(n19362), .B2(n19610), .A(n19361), .ZN(n19365) );
  NOR3_X1 U22292 ( .A1(n19365), .A2(n19364), .A3(n19363), .ZN(n19366) );
  OAI21_X1 U22293 ( .B1(n19395), .B2(n19839), .A(n19366), .ZN(n19386) );
  AOI22_X1 U22294 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19386), .B1(
        n19411), .B2(n19665), .ZN(n19368) );
  OAI211_X1 U22295 ( .C1(n19668), .C2(n19389), .A(n19369), .B(n19368), .ZN(
        P2_U3104) );
  NOR2_X1 U22296 ( .A1(n19499), .A2(n19392), .ZN(n19370) );
  AOI21_X1 U22297 ( .B1(n19385), .B2(n14299), .A(n19370), .ZN(n19372) );
  AOI22_X1 U22298 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19386), .B1(
        n19411), .B2(n19670), .ZN(n19371) );
  OAI211_X1 U22299 ( .C1(n19673), .C2(n19389), .A(n19372), .B(n19371), .ZN(
        P2_U3105) );
  AOI22_X1 U22300 ( .A1(n19385), .A2(n19151), .B1(n19395), .B2(n19674), .ZN(
        n19374) );
  AOI22_X1 U22301 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19386), .B1(
        n19411), .B2(n19675), .ZN(n19373) );
  OAI211_X1 U22302 ( .C1(n19678), .C2(n19389), .A(n19374), .B(n19373), .ZN(
        P2_U3106) );
  AOI22_X1 U22303 ( .A1(n19385), .A2(n19680), .B1(n19395), .B2(n19679), .ZN(
        n19376) );
  AOI22_X1 U22304 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19386), .B1(
        n19411), .B2(n19681), .ZN(n19375) );
  OAI211_X1 U22305 ( .C1(n19684), .C2(n19389), .A(n19376), .B(n19375), .ZN(
        P2_U3107) );
  AOI22_X1 U22306 ( .A1(n19385), .A2(n19686), .B1(n19395), .B2(n19685), .ZN(
        n19378) );
  AOI22_X1 U22307 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19386), .B1(
        n19411), .B2(n19687), .ZN(n19377) );
  OAI211_X1 U22308 ( .C1(n19690), .C2(n19389), .A(n19378), .B(n19377), .ZN(
        P2_U3108) );
  NOR2_X1 U22309 ( .A1(n19521), .A2(n19392), .ZN(n19379) );
  AOI21_X1 U22310 ( .B1(n19385), .B2(n19692), .A(n19379), .ZN(n19381) );
  AOI22_X1 U22311 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19386), .B1(
        n19411), .B2(n19693), .ZN(n19380) );
  OAI211_X1 U22312 ( .C1(n19696), .C2(n19389), .A(n19381), .B(n19380), .ZN(
        P2_U3109) );
  NOR2_X1 U22313 ( .A1(n19526), .A2(n19392), .ZN(n19382) );
  AOI21_X1 U22314 ( .B1(n19385), .B2(n19698), .A(n19382), .ZN(n19384) );
  AOI22_X1 U22315 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19386), .B1(
        n19411), .B2(n19699), .ZN(n19383) );
  OAI211_X1 U22316 ( .C1(n19702), .C2(n19389), .A(n19384), .B(n19383), .ZN(
        P2_U3110) );
  AOI22_X1 U22317 ( .A1(n19385), .A2(n19705), .B1(n19395), .B2(n19704), .ZN(
        n19388) );
  AOI22_X1 U22318 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19386), .B1(
        n19411), .B2(n19707), .ZN(n19387) );
  OAI211_X1 U22319 ( .C1(n19713), .C2(n19389), .A(n19388), .B(n19387), .ZN(
        P2_U3111) );
  INV_X1 U22320 ( .A(n19420), .ZN(n19422) );
  INV_X1 U22321 ( .A(n19449), .ZN(n19437) );
  NAND2_X1 U22322 ( .A1(n19813), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19486) );
  INV_X1 U22323 ( .A(n19486), .ZN(n19483) );
  NAND2_X1 U22324 ( .A1(n19483), .A2(n19822), .ZN(n19427) );
  NOR2_X1 U22325 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19427), .ZN(
        n19414) );
  AOI22_X1 U22326 ( .A1(n19665), .A2(n19437), .B1(n19657), .B2(n19414), .ZN(
        n19400) );
  NAND2_X1 U22327 ( .A1(n19449), .A2(n19419), .ZN(n19390) );
  AOI21_X1 U22328 ( .B1(n19390), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19797), 
        .ZN(n19394) );
  AOI21_X1 U22329 ( .B1(n19396), .B2(n19839), .A(n19793), .ZN(n19391) );
  AOI21_X1 U22330 ( .B1(n19394), .B2(n19392), .A(n19391), .ZN(n19393) );
  OAI21_X1 U22331 ( .B1(n19414), .B2(n19393), .A(n19662), .ZN(n19416) );
  OAI21_X1 U22332 ( .B1(n19395), .B2(n19414), .A(n19394), .ZN(n19398) );
  OAI21_X1 U22333 ( .B1(n19396), .B2(n19414), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19397) );
  NAND2_X1 U22334 ( .A1(n19398), .A2(n19397), .ZN(n19415) );
  AOI22_X1 U22335 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19416), .B1(
        n14284), .B2(n19415), .ZN(n19399) );
  OAI211_X1 U22336 ( .C1(n19668), .C2(n19419), .A(n19400), .B(n19399), .ZN(
        P2_U3112) );
  AOI22_X1 U22337 ( .A1(n19670), .A2(n19437), .B1(n19669), .B2(n19414), .ZN(
        n19402) );
  AOI22_X1 U22338 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19416), .B1(
        n19415), .B2(n14299), .ZN(n19401) );
  OAI211_X1 U22339 ( .C1(n19673), .C2(n19419), .A(n19402), .B(n19401), .ZN(
        P2_U3113) );
  AOI22_X1 U22340 ( .A1(n19507), .A2(n19411), .B1(n19674), .B2(n19414), .ZN(
        n19404) );
  AOI22_X1 U22341 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19416), .B1(
        n19415), .B2(n19151), .ZN(n19403) );
  OAI211_X1 U22342 ( .C1(n19510), .C2(n19449), .A(n19404), .B(n19403), .ZN(
        P2_U3114) );
  AOI22_X1 U22343 ( .A1(n19632), .A2(n19411), .B1(n19679), .B2(n19414), .ZN(
        n19406) );
  AOI22_X1 U22344 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19416), .B1(
        n19415), .B2(n19680), .ZN(n19405) );
  OAI211_X1 U22345 ( .C1(n19635), .C2(n19449), .A(n19406), .B(n19405), .ZN(
        P2_U3115) );
  AOI22_X1 U22346 ( .A1(n19636), .A2(n19411), .B1(n19685), .B2(n19414), .ZN(
        n19408) );
  AOI22_X1 U22347 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19416), .B1(
        n19415), .B2(n19686), .ZN(n19407) );
  OAI211_X1 U22348 ( .C1(n19639), .C2(n19449), .A(n19408), .B(n19407), .ZN(
        P2_U3116) );
  AOI22_X1 U22349 ( .A1(n19640), .A2(n19411), .B1(n19691), .B2(n19414), .ZN(
        n19410) );
  AOI22_X1 U22350 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19416), .B1(
        n19415), .B2(n19692), .ZN(n19409) );
  OAI211_X1 U22351 ( .C1(n19643), .C2(n19449), .A(n19410), .B(n19409), .ZN(
        P2_U3117) );
  AOI22_X1 U22352 ( .A1(n19600), .A2(n19411), .B1(n19697), .B2(n19414), .ZN(
        n19413) );
  AOI22_X1 U22353 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19416), .B1(
        n19415), .B2(n19698), .ZN(n19412) );
  OAI211_X1 U22354 ( .C1(n19604), .C2(n19449), .A(n19413), .B(n19412), .ZN(
        P2_U3118) );
  AOI22_X1 U22355 ( .A1(n19707), .A2(n19437), .B1(n19704), .B2(n19414), .ZN(
        n19418) );
  AOI22_X1 U22356 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19416), .B1(
        n19415), .B2(n19705), .ZN(n19417) );
  OAI211_X1 U22357 ( .C1(n19713), .C2(n19419), .A(n19418), .B(n19417), .ZN(
        P2_U3119) );
  NOR2_X2 U22358 ( .A1(n19584), .A2(n19420), .ZN(n19471) );
  NOR2_X1 U22359 ( .A1(n19421), .A2(n19486), .ZN(n19444) );
  AOI22_X1 U22360 ( .A1(n19665), .A2(n19471), .B1(n19657), .B2(n19444), .ZN(
        n19430) );
  INV_X1 U22361 ( .A(n19444), .ZN(n19456) );
  NAND2_X1 U22362 ( .A1(n19456), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19424) );
  NOR2_X1 U22363 ( .A1(n19795), .A2(n19791), .ZN(n19659) );
  AOI21_X1 U22364 ( .B1(n19659), .B2(n19422), .A(n19797), .ZN(n19425) );
  AOI22_X1 U22365 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19456), .B1(n19425), 
        .B2(n19427), .ZN(n19423) );
  OAI211_X1 U22366 ( .C1(n10469), .C2(n19424), .A(n19662), .B(n19423), .ZN(
        n19446) );
  INV_X1 U22367 ( .A(n19425), .ZN(n19428) );
  OAI21_X1 U22368 ( .B1(n10469), .B2(n19444), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19426) );
  AOI22_X1 U22369 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19446), .B1(
        n14284), .B2(n19445), .ZN(n19429) );
  OAI211_X1 U22370 ( .C1(n19668), .C2(n19449), .A(n19430), .B(n19429), .ZN(
        P2_U3120) );
  AOI22_X1 U22371 ( .A1(n19670), .A2(n19471), .B1(n19669), .B2(n19444), .ZN(
        n19432) );
  AOI22_X1 U22372 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19446), .B1(
        n14299), .B2(n19445), .ZN(n19431) );
  OAI211_X1 U22373 ( .C1(n19673), .C2(n19449), .A(n19432), .B(n19431), .ZN(
        P2_U3121) );
  INV_X1 U22374 ( .A(n19471), .ZN(n19480) );
  AOI22_X1 U22375 ( .A1(n19507), .A2(n19437), .B1(n19674), .B2(n19444), .ZN(
        n19434) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19446), .B1(
        n19151), .B2(n19445), .ZN(n19433) );
  OAI211_X1 U22377 ( .C1(n19510), .C2(n19480), .A(n19434), .B(n19433), .ZN(
        P2_U3122) );
  AOI22_X1 U22378 ( .A1(n19681), .A2(n19471), .B1(n19679), .B2(n19444), .ZN(
        n19436) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19446), .B1(
        n19680), .B2(n19445), .ZN(n19435) );
  OAI211_X1 U22380 ( .C1(n19684), .C2(n19449), .A(n19436), .B(n19435), .ZN(
        P2_U3123) );
  AOI22_X1 U22381 ( .A1(n19636), .A2(n19437), .B1(n19685), .B2(n19444), .ZN(
        n19439) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19446), .B1(
        n19686), .B2(n19445), .ZN(n19438) );
  OAI211_X1 U22383 ( .C1(n19639), .C2(n19480), .A(n19439), .B(n19438), .ZN(
        P2_U3124) );
  AOI22_X1 U22384 ( .A1(n19693), .A2(n19471), .B1(n19691), .B2(n19444), .ZN(
        n19441) );
  AOI22_X1 U22385 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19446), .B1(
        n19692), .B2(n19445), .ZN(n19440) );
  OAI211_X1 U22386 ( .C1(n19696), .C2(n19449), .A(n19441), .B(n19440), .ZN(
        P2_U3125) );
  AOI22_X1 U22387 ( .A1(n19699), .A2(n19471), .B1(n19697), .B2(n19444), .ZN(
        n19443) );
  AOI22_X1 U22388 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19446), .B1(
        n19698), .B2(n19445), .ZN(n19442) );
  OAI211_X1 U22389 ( .C1(n19702), .C2(n19449), .A(n19443), .B(n19442), .ZN(
        P2_U3126) );
  AOI22_X1 U22390 ( .A1(n19707), .A2(n19471), .B1(n19704), .B2(n19444), .ZN(
        n19448) );
  AOI22_X1 U22391 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19446), .B1(
        n19705), .B2(n19445), .ZN(n19447) );
  OAI211_X1 U22392 ( .C1(n19713), .C2(n19449), .A(n19448), .B(n19447), .ZN(
        P2_U3127) );
  INV_X1 U22393 ( .A(n19450), .ZN(n19453) );
  AND2_X1 U22394 ( .A1(n19451), .A2(n19483), .ZN(n19475) );
  OAI21_X1 U22395 ( .B1(n19454), .B2(n19475), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19452) );
  OAI21_X1 U22396 ( .B1(n19486), .B2(n19453), .A(n19452), .ZN(n19476) );
  AOI22_X1 U22397 ( .A1(n19476), .A2(n14284), .B1(n19657), .B2(n19475), .ZN(
        n19460) );
  NAND2_X1 U22398 ( .A1(n19611), .A2(n19790), .ZN(n19474) );
  OAI21_X1 U22399 ( .B1(n19471), .B2(n19536), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19457) );
  NOR2_X1 U22400 ( .A1(n19454), .A2(n19848), .ZN(n19455) );
  AOI211_X1 U22401 ( .C1(n19457), .C2(n19456), .A(P2_STATE2_REG_3__SCAN_IN), 
        .B(n19455), .ZN(n19458) );
  OAI21_X1 U22402 ( .B1(n19458), .B2(n19475), .A(n19662), .ZN(n19477) );
  AOI22_X1 U22403 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19477), .B1(
        n19536), .B2(n19665), .ZN(n19459) );
  OAI211_X1 U22404 ( .C1(n19668), .C2(n19480), .A(n19460), .B(n19459), .ZN(
        P2_U3128) );
  AOI22_X1 U22405 ( .A1(n19476), .A2(n14299), .B1(n19669), .B2(n19475), .ZN(
        n19462) );
  AOI22_X1 U22406 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19477), .B1(
        n19536), .B2(n19670), .ZN(n19461) );
  OAI211_X1 U22407 ( .C1(n19673), .C2(n19480), .A(n19462), .B(n19461), .ZN(
        P2_U3129) );
  AOI22_X1 U22408 ( .A1(n19476), .A2(n19151), .B1(n19674), .B2(n19475), .ZN(
        n19464) );
  AOI22_X1 U22409 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19477), .B1(
        n19471), .B2(n19507), .ZN(n19463) );
  OAI211_X1 U22410 ( .C1(n19510), .C2(n19474), .A(n19464), .B(n19463), .ZN(
        P2_U3130) );
  AOI22_X1 U22411 ( .A1(n19476), .A2(n19680), .B1(n19679), .B2(n19475), .ZN(
        n19466) );
  AOI22_X1 U22412 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19477), .B1(
        n19471), .B2(n19632), .ZN(n19465) );
  OAI211_X1 U22413 ( .C1(n19635), .C2(n19474), .A(n19466), .B(n19465), .ZN(
        P2_U3131) );
  AOI22_X1 U22414 ( .A1(n19476), .A2(n19686), .B1(n19685), .B2(n19475), .ZN(
        n19468) );
  AOI22_X1 U22415 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19477), .B1(
        n19471), .B2(n19636), .ZN(n19467) );
  OAI211_X1 U22416 ( .C1(n19639), .C2(n19474), .A(n19468), .B(n19467), .ZN(
        P2_U3132) );
  AOI22_X1 U22417 ( .A1(n19476), .A2(n19692), .B1(n19691), .B2(n19475), .ZN(
        n19470) );
  AOI22_X1 U22418 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19477), .B1(
        n19471), .B2(n19640), .ZN(n19469) );
  OAI211_X1 U22419 ( .C1(n19643), .C2(n19474), .A(n19470), .B(n19469), .ZN(
        P2_U3133) );
  AOI22_X1 U22420 ( .A1(n19476), .A2(n19698), .B1(n19697), .B2(n19475), .ZN(
        n19473) );
  AOI22_X1 U22421 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19477), .B1(
        n19471), .B2(n19600), .ZN(n19472) );
  OAI211_X1 U22422 ( .C1(n19604), .C2(n19474), .A(n19473), .B(n19472), .ZN(
        P2_U3134) );
  AOI22_X1 U22423 ( .A1(n19476), .A2(n19705), .B1(n19704), .B2(n19475), .ZN(
        n19479) );
  AOI22_X1 U22424 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19477), .B1(
        n19536), .B2(n19707), .ZN(n19478) );
  OAI211_X1 U22425 ( .C1(n19713), .C2(n19480), .A(n19479), .B(n19478), .ZN(
        P2_U3135) );
  INV_X1 U22426 ( .A(n19482), .ZN(n19484) );
  NAND2_X1 U22427 ( .A1(n19484), .A2(n19483), .ZN(n19531) );
  NAND2_X1 U22428 ( .A1(n19531), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19485) );
  NOR2_X1 U22429 ( .A1(n19822), .A2(n19486), .ZN(n19496) );
  INV_X1 U22430 ( .A(n19496), .ZN(n19487) );
  OAI21_X1 U22431 ( .B1(n19487), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19848), 
        .ZN(n19488) );
  NAND2_X1 U22432 ( .A1(n19492), .A2(n19488), .ZN(n19534) );
  INV_X1 U22433 ( .A(n14284), .ZN(n19490) );
  OAI22_X1 U22434 ( .A1(n19534), .A2(n19490), .B1(n19489), .B2(n19531), .ZN(
        n19491) );
  INV_X1 U22435 ( .A(n19491), .ZN(n19498) );
  INV_X1 U22436 ( .A(n19531), .ZN(n19493) );
  OAI211_X1 U22437 ( .C1(n19493), .C2(n19839), .A(n19492), .B(n19662), .ZN(
        n19494) );
  INV_X1 U22438 ( .A(n19494), .ZN(n19495) );
  OAI221_X1 U22439 ( .B1(n19496), .B2(n19790), .C1(n19496), .C2(n19659), .A(
        n19495), .ZN(n19537) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19537), .B1(
        n19536), .B2(n19613), .ZN(n19497) );
  OAI211_X1 U22441 ( .C1(n19625), .C2(n19571), .A(n19498), .B(n19497), .ZN(
        P2_U3136) );
  INV_X1 U22442 ( .A(n14299), .ZN(n19500) );
  OAI22_X1 U22443 ( .A1(n19534), .A2(n19500), .B1(n19499), .B2(n19531), .ZN(
        n19501) );
  INV_X1 U22444 ( .A(n19501), .ZN(n19503) );
  AOI22_X1 U22445 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19537), .B1(
        n19536), .B2(n19626), .ZN(n19502) );
  OAI211_X1 U22446 ( .C1(n19629), .C2(n19571), .A(n19503), .B(n19502), .ZN(
        P2_U3137) );
  INV_X1 U22447 ( .A(n19151), .ZN(n19505) );
  INV_X1 U22448 ( .A(n19674), .ZN(n19504) );
  OAI22_X1 U22449 ( .A1(n19534), .A2(n19505), .B1(n19504), .B2(n19531), .ZN(
        n19506) );
  INV_X1 U22450 ( .A(n19506), .ZN(n19509) );
  AOI22_X1 U22451 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19537), .B1(
        n19536), .B2(n19507), .ZN(n19508) );
  OAI211_X1 U22452 ( .C1(n19510), .C2(n19571), .A(n19509), .B(n19508), .ZN(
        P2_U3138) );
  INV_X1 U22453 ( .A(n19680), .ZN(n19512) );
  INV_X1 U22454 ( .A(n19679), .ZN(n19511) );
  OAI22_X1 U22455 ( .A1(n19534), .A2(n19512), .B1(n19511), .B2(n19531), .ZN(
        n19513) );
  INV_X1 U22456 ( .A(n19513), .ZN(n19515) );
  AOI22_X1 U22457 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19537), .B1(
        n19536), .B2(n19632), .ZN(n19514) );
  OAI211_X1 U22458 ( .C1(n19635), .C2(n19571), .A(n19515), .B(n19514), .ZN(
        P2_U3139) );
  INV_X1 U22459 ( .A(n19686), .ZN(n19517) );
  INV_X1 U22460 ( .A(n19685), .ZN(n19516) );
  OAI22_X1 U22461 ( .A1(n19534), .A2(n19517), .B1(n19516), .B2(n19531), .ZN(
        n19518) );
  INV_X1 U22462 ( .A(n19518), .ZN(n19520) );
  AOI22_X1 U22463 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19537), .B1(
        n19536), .B2(n19636), .ZN(n19519) );
  OAI211_X1 U22464 ( .C1(n19639), .C2(n19571), .A(n19520), .B(n19519), .ZN(
        P2_U3140) );
  INV_X1 U22465 ( .A(n19692), .ZN(n19522) );
  OAI22_X1 U22466 ( .A1(n19534), .A2(n19522), .B1(n19521), .B2(n19531), .ZN(
        n19523) );
  INV_X1 U22467 ( .A(n19523), .ZN(n19525) );
  AOI22_X1 U22468 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19537), .B1(
        n19536), .B2(n19640), .ZN(n19524) );
  OAI211_X1 U22469 ( .C1(n19643), .C2(n19571), .A(n19525), .B(n19524), .ZN(
        P2_U3141) );
  INV_X1 U22470 ( .A(n19698), .ZN(n19527) );
  OAI22_X1 U22471 ( .A1(n19534), .A2(n19527), .B1(n19526), .B2(n19531), .ZN(
        n19528) );
  INV_X1 U22472 ( .A(n19528), .ZN(n19530) );
  AOI22_X1 U22473 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19537), .B1(
        n19536), .B2(n19600), .ZN(n19529) );
  OAI211_X1 U22474 ( .C1(n19604), .C2(n19571), .A(n19530), .B(n19529), .ZN(
        P2_U3142) );
  INV_X1 U22475 ( .A(n19705), .ZN(n19533) );
  INV_X1 U22476 ( .A(n19704), .ZN(n19532) );
  OAI22_X1 U22477 ( .A1(n19534), .A2(n19533), .B1(n19532), .B2(n19531), .ZN(
        n19535) );
  INV_X1 U22478 ( .A(n19535), .ZN(n19539) );
  AOI22_X1 U22479 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19537), .B1(
        n19536), .B2(n19650), .ZN(n19538) );
  OAI211_X1 U22480 ( .C1(n19655), .C2(n19571), .A(n19539), .B(n19538), .ZN(
        P2_U3143) );
  INV_X1 U22481 ( .A(n19540), .ZN(n19544) );
  INV_X1 U22482 ( .A(n19550), .ZN(n19543) );
  NAND3_X1 U22483 ( .A1(n19822), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19580) );
  NOR2_X1 U22484 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19580), .ZN(
        n19566) );
  OAI21_X1 U22485 ( .B1(n19541), .B2(n19566), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19542) );
  OAI21_X1 U22486 ( .B1(n19544), .B2(n19543), .A(n19542), .ZN(n19567) );
  AOI22_X1 U22487 ( .A1(n19567), .A2(n14284), .B1(n19657), .B2(n19566), .ZN(
        n19553) );
  INV_X1 U22488 ( .A(n19611), .ZN(n19545) );
  AOI21_X1 U22489 ( .B1(n19571), .B2(n19609), .A(n19791), .ZN(n19551) );
  INV_X1 U22490 ( .A(n19566), .ZN(n19546) );
  OAI211_X1 U22491 ( .C1(n19547), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19546), 
        .B(n19797), .ZN(n19548) );
  AND2_X1 U22492 ( .A1(n19548), .A2(n19662), .ZN(n19549) );
  OAI211_X1 U22493 ( .C1(n19551), .C2(n19550), .A(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n19549), .ZN(n19568) );
  AOI22_X1 U22494 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19568), .B1(
        n19601), .B2(n19665), .ZN(n19552) );
  OAI211_X1 U22495 ( .C1(n19668), .C2(n19571), .A(n19553), .B(n19552), .ZN(
        P2_U3144) );
  AOI22_X1 U22496 ( .A1(n19567), .A2(n14299), .B1(n19669), .B2(n19566), .ZN(
        n19555) );
  AOI22_X1 U22497 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19568), .B1(
        n19601), .B2(n19670), .ZN(n19554) );
  OAI211_X1 U22498 ( .C1(n19673), .C2(n19571), .A(n19555), .B(n19554), .ZN(
        P2_U3145) );
  AOI22_X1 U22499 ( .A1(n19567), .A2(n19151), .B1(n19674), .B2(n19566), .ZN(
        n19557) );
  AOI22_X1 U22500 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19568), .B1(
        n19601), .B2(n19675), .ZN(n19556) );
  OAI211_X1 U22501 ( .C1(n19678), .C2(n19571), .A(n19557), .B(n19556), .ZN(
        P2_U3146) );
  AOI22_X1 U22502 ( .A1(n19567), .A2(n19680), .B1(n19679), .B2(n19566), .ZN(
        n19559) );
  AOI22_X1 U22503 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19568), .B1(
        n19601), .B2(n19681), .ZN(n19558) );
  OAI211_X1 U22504 ( .C1(n19684), .C2(n19571), .A(n19559), .B(n19558), .ZN(
        P2_U3147) );
  AOI22_X1 U22505 ( .A1(n19567), .A2(n19686), .B1(n19685), .B2(n19566), .ZN(
        n19561) );
  AOI22_X1 U22506 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19568), .B1(
        n19601), .B2(n19687), .ZN(n19560) );
  OAI211_X1 U22507 ( .C1(n19690), .C2(n19571), .A(n19561), .B(n19560), .ZN(
        P2_U3148) );
  AOI22_X1 U22508 ( .A1(n19567), .A2(n19692), .B1(n19691), .B2(n19566), .ZN(
        n19563) );
  AOI22_X1 U22509 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19568), .B1(
        n19601), .B2(n19693), .ZN(n19562) );
  OAI211_X1 U22510 ( .C1(n19696), .C2(n19571), .A(n19563), .B(n19562), .ZN(
        P2_U3149) );
  AOI22_X1 U22511 ( .A1(n19567), .A2(n19698), .B1(n19697), .B2(n19566), .ZN(
        n19565) );
  AOI22_X1 U22512 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19568), .B1(
        n19601), .B2(n19699), .ZN(n19564) );
  OAI211_X1 U22513 ( .C1(n19702), .C2(n19571), .A(n19565), .B(n19564), .ZN(
        P2_U3150) );
  AOI22_X1 U22514 ( .A1(n19567), .A2(n19705), .B1(n19704), .B2(n19566), .ZN(
        n19570) );
  AOI22_X1 U22515 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19568), .B1(
        n19601), .B2(n19707), .ZN(n19569) );
  OAI211_X1 U22516 ( .C1(n19713), .C2(n19571), .A(n19570), .B(n19569), .ZN(
        P2_U3151) );
  INV_X1 U22517 ( .A(n19583), .ZN(n19572) );
  NAND2_X1 U22518 ( .A1(n19659), .A2(n19572), .ZN(n19573) );
  NAND2_X1 U22519 ( .A1(n19573), .A2(n19580), .ZN(n19579) );
  NOR2_X1 U22520 ( .A1(n19828), .A2(n19580), .ZN(n19615) );
  INV_X1 U22521 ( .A(n19615), .ZN(n19574) );
  AND2_X1 U22522 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19574), .ZN(n19575) );
  NAND2_X1 U22523 ( .A1(n19576), .A2(n19575), .ZN(n19582) );
  OAI211_X1 U22524 ( .C1(n19615), .C2(n19839), .A(n19582), .B(n19662), .ZN(
        n19577) );
  INV_X1 U22525 ( .A(n19577), .ZN(n19578) );
  INV_X1 U22526 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n19587) );
  OAI21_X1 U22527 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19580), .A(n19848), 
        .ZN(n19581) );
  AND2_X1 U22528 ( .A1(n19582), .A2(n19581), .ZN(n19605) );
  AOI22_X1 U22529 ( .A1(n19605), .A2(n14284), .B1(n19657), .B2(n19615), .ZN(
        n19586) );
  AOI22_X1 U22530 ( .A1(n19649), .A2(n19665), .B1(n19601), .B2(n19613), .ZN(
        n19585) );
  OAI211_X1 U22531 ( .C1(n19597), .C2(n19587), .A(n19586), .B(n19585), .ZN(
        P2_U3152) );
  AOI22_X1 U22532 ( .A1(n19605), .A2(n14299), .B1(n19669), .B2(n19615), .ZN(
        n19589) );
  AOI22_X1 U22533 ( .A1(n19649), .A2(n19670), .B1(n19601), .B2(n19626), .ZN(
        n19588) );
  OAI211_X1 U22534 ( .C1(n19597), .C2(n10421), .A(n19589), .B(n19588), .ZN(
        P2_U3153) );
  AOI22_X1 U22535 ( .A1(n19605), .A2(n19151), .B1(n19674), .B2(n19615), .ZN(
        n19591) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19606), .B1(
        n19649), .B2(n19675), .ZN(n19590) );
  OAI211_X1 U22537 ( .C1(n19678), .C2(n19609), .A(n19591), .B(n19590), .ZN(
        P2_U3154) );
  AOI22_X1 U22538 ( .A1(n19605), .A2(n19680), .B1(n19679), .B2(n19615), .ZN(
        n19593) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19606), .B1(
        n19649), .B2(n19681), .ZN(n19592) );
  OAI211_X1 U22540 ( .C1(n19684), .C2(n19609), .A(n19593), .B(n19592), .ZN(
        P2_U3155) );
  INV_X1 U22541 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n19596) );
  AOI22_X1 U22542 ( .A1(n19605), .A2(n19686), .B1(n19685), .B2(n19615), .ZN(
        n19595) );
  AOI22_X1 U22543 ( .A1(n19601), .A2(n19636), .B1(n19649), .B2(n19687), .ZN(
        n19594) );
  OAI211_X1 U22544 ( .C1(n19597), .C2(n19596), .A(n19595), .B(n19594), .ZN(
        P2_U3156) );
  AOI22_X1 U22545 ( .A1(n19605), .A2(n19692), .B1(n19691), .B2(n19615), .ZN(
        n19599) );
  AOI22_X1 U22546 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19606), .B1(
        n19649), .B2(n19693), .ZN(n19598) );
  OAI211_X1 U22547 ( .C1(n19696), .C2(n19609), .A(n19599), .B(n19598), .ZN(
        P2_U3157) );
  INV_X1 U22548 ( .A(n19649), .ZN(n19647) );
  AOI22_X1 U22549 ( .A1(n19605), .A2(n19698), .B1(n19697), .B2(n19615), .ZN(
        n19603) );
  AOI22_X1 U22550 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19606), .B1(
        n19601), .B2(n19600), .ZN(n19602) );
  OAI211_X1 U22551 ( .C1(n19604), .C2(n19647), .A(n19603), .B(n19602), .ZN(
        P2_U3158) );
  AOI22_X1 U22552 ( .A1(n19605), .A2(n19705), .B1(n19704), .B2(n19615), .ZN(
        n19608) );
  AOI22_X1 U22553 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19606), .B1(
        n19649), .B2(n19707), .ZN(n19607) );
  OAI211_X1 U22554 ( .C1(n19713), .C2(n19609), .A(n19608), .B(n19607), .ZN(
        P2_U3159) );
  NAND2_X1 U22555 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19612), .ZN(
        n19660) );
  NOR2_X1 U22556 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19660), .ZN(
        n19648) );
  AOI22_X1 U22557 ( .A1(n19613), .A2(n19649), .B1(n19657), .B2(n19648), .ZN(
        n19624) );
  INV_X1 U22558 ( .A(n19712), .ZN(n19644) );
  OAI21_X1 U22559 ( .B1(n19644), .B2(n19649), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19614) );
  NAND2_X1 U22560 ( .A1(n19614), .A2(n19793), .ZN(n19622) );
  NOR2_X1 U22561 ( .A1(n19648), .A2(n19615), .ZN(n19621) );
  INV_X1 U22562 ( .A(n19621), .ZN(n19618) );
  INV_X1 U22563 ( .A(n19648), .ZN(n19616) );
  OAI211_X1 U22564 ( .C1(n10474), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19616), 
        .B(n19797), .ZN(n19617) );
  OAI211_X1 U22565 ( .C1(n19622), .C2(n19618), .A(n19662), .B(n19617), .ZN(
        n19652) );
  INV_X1 U22566 ( .A(n10474), .ZN(n19619) );
  OAI21_X1 U22567 ( .B1(n19619), .B2(n19648), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19620) );
  AOI22_X1 U22568 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19652), .B1(
        n14284), .B2(n19651), .ZN(n19623) );
  OAI211_X1 U22569 ( .C1(n19625), .C2(n19712), .A(n19624), .B(n19623), .ZN(
        P2_U3160) );
  AOI22_X1 U22570 ( .A1(n19626), .A2(n19649), .B1(n19669), .B2(n19648), .ZN(
        n19628) );
  AOI22_X1 U22571 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19652), .B1(
        n14299), .B2(n19651), .ZN(n19627) );
  OAI211_X1 U22572 ( .C1(n19629), .C2(n19712), .A(n19628), .B(n19627), .ZN(
        P2_U3161) );
  AOI22_X1 U22573 ( .A1(n19675), .A2(n19644), .B1(n19674), .B2(n19648), .ZN(
        n19631) );
  AOI22_X1 U22574 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19652), .B1(
        n19151), .B2(n19651), .ZN(n19630) );
  OAI211_X1 U22575 ( .C1(n19678), .C2(n19647), .A(n19631), .B(n19630), .ZN(
        P2_U3162) );
  AOI22_X1 U22576 ( .A1(n19632), .A2(n19649), .B1(n19679), .B2(n19648), .ZN(
        n19634) );
  AOI22_X1 U22577 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19652), .B1(
        n19680), .B2(n19651), .ZN(n19633) );
  OAI211_X1 U22578 ( .C1(n19635), .C2(n19712), .A(n19634), .B(n19633), .ZN(
        P2_U3163) );
  AOI22_X1 U22579 ( .A1(n19636), .A2(n19649), .B1(n19685), .B2(n19648), .ZN(
        n19638) );
  AOI22_X1 U22580 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19652), .B1(
        n19686), .B2(n19651), .ZN(n19637) );
  OAI211_X1 U22581 ( .C1(n19639), .C2(n19712), .A(n19638), .B(n19637), .ZN(
        P2_U3164) );
  AOI22_X1 U22582 ( .A1(n19640), .A2(n19649), .B1(n19691), .B2(n19648), .ZN(
        n19642) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19652), .B1(
        n19692), .B2(n19651), .ZN(n19641) );
  OAI211_X1 U22584 ( .C1(n19643), .C2(n19712), .A(n19642), .B(n19641), .ZN(
        P2_U3165) );
  AOI22_X1 U22585 ( .A1(n19699), .A2(n19644), .B1(n19697), .B2(n19648), .ZN(
        n19646) );
  AOI22_X1 U22586 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19652), .B1(
        n19698), .B2(n19651), .ZN(n19645) );
  OAI211_X1 U22587 ( .C1(n19702), .C2(n19647), .A(n19646), .B(n19645), .ZN(
        P2_U3166) );
  AOI22_X1 U22588 ( .A1(n19650), .A2(n19649), .B1(n19704), .B2(n19648), .ZN(
        n19654) );
  AOI22_X1 U22589 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19652), .B1(
        n19705), .B2(n19651), .ZN(n19653) );
  OAI211_X1 U22590 ( .C1(n19655), .C2(n19712), .A(n19654), .B(n19653), .ZN(
        P2_U3167) );
  OAI21_X1 U22591 ( .B1(n10468), .B2(n19703), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19656) );
  OAI21_X1 U22592 ( .B1(n19660), .B2(n19797), .A(n19656), .ZN(n19706) );
  AOI22_X1 U22593 ( .A1(n19706), .A2(n14284), .B1(n19657), .B2(n19703), .ZN(
        n19667) );
  INV_X1 U22594 ( .A(n10468), .ZN(n19658) );
  AOI21_X1 U22595 ( .B1(n19658), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19664) );
  INV_X1 U22596 ( .A(n19659), .ZN(n19661) );
  OAI21_X1 U22597 ( .B1(n19661), .B2(n19796), .A(n19660), .ZN(n19663) );
  OAI211_X1 U22598 ( .C1(n19703), .C2(n19664), .A(n19663), .B(n19662), .ZN(
        n19709) );
  AOI22_X1 U22599 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19665), .ZN(n19666) );
  OAI211_X1 U22600 ( .C1(n19668), .C2(n19712), .A(n19667), .B(n19666), .ZN(
        P2_U3168) );
  AOI22_X1 U22601 ( .A1(n19706), .A2(n14299), .B1(n19669), .B2(n19703), .ZN(
        n19672) );
  AOI22_X1 U22602 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19670), .ZN(n19671) );
  OAI211_X1 U22603 ( .C1(n19673), .C2(n19712), .A(n19672), .B(n19671), .ZN(
        P2_U3169) );
  AOI22_X1 U22604 ( .A1(n19706), .A2(n19151), .B1(n19674), .B2(n19703), .ZN(
        n19677) );
  AOI22_X1 U22605 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19675), .ZN(n19676) );
  OAI211_X1 U22606 ( .C1(n19678), .C2(n19712), .A(n19677), .B(n19676), .ZN(
        P2_U3170) );
  AOI22_X1 U22607 ( .A1(n19706), .A2(n19680), .B1(n19679), .B2(n19703), .ZN(
        n19683) );
  AOI22_X1 U22608 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19681), .ZN(n19682) );
  OAI211_X1 U22609 ( .C1(n19684), .C2(n19712), .A(n19683), .B(n19682), .ZN(
        P2_U3171) );
  AOI22_X1 U22610 ( .A1(n19706), .A2(n19686), .B1(n19685), .B2(n19703), .ZN(
        n19689) );
  AOI22_X1 U22611 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19687), .ZN(n19688) );
  OAI211_X1 U22612 ( .C1(n19690), .C2(n19712), .A(n19689), .B(n19688), .ZN(
        P2_U3172) );
  AOI22_X1 U22613 ( .A1(n19706), .A2(n19692), .B1(n19691), .B2(n19703), .ZN(
        n19695) );
  AOI22_X1 U22614 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19693), .ZN(n19694) );
  OAI211_X1 U22615 ( .C1(n19696), .C2(n19712), .A(n19695), .B(n19694), .ZN(
        P2_U3173) );
  AOI22_X1 U22616 ( .A1(n19706), .A2(n19698), .B1(n19697), .B2(n19703), .ZN(
        n19701) );
  AOI22_X1 U22617 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19699), .ZN(n19700) );
  OAI211_X1 U22618 ( .C1(n19702), .C2(n19712), .A(n19701), .B(n19700), .ZN(
        P2_U3174) );
  AOI22_X1 U22619 ( .A1(n19706), .A2(n19705), .B1(n19704), .B2(n19703), .ZN(
        n19711) );
  AOI22_X1 U22620 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19709), .B1(
        n19708), .B2(n19707), .ZN(n19710) );
  OAI211_X1 U22621 ( .C1(n19713), .C2(n19712), .A(n19711), .B(n19710), .ZN(
        P2_U3175) );
  OAI221_X1 U22622 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19839), .C1(
        P2_STATE2_REG_2__SCAN_IN), .C2(n19721), .A(n19714), .ZN(n19718) );
  OAI211_X1 U22623 ( .C1(n19719), .C2(n19715), .A(n19849), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19716) );
  OAI211_X1 U22624 ( .C1(n19719), .C2(n19718), .A(n19717), .B(n19716), .ZN(
        P2_U3177) );
  AND2_X1 U22625 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19720), .ZN(
        P2_U3179) );
  AND2_X1 U22626 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19720), .ZN(
        P2_U3180) );
  AND2_X1 U22627 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19720), .ZN(
        P2_U3181) );
  AND2_X1 U22628 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19720), .ZN(
        P2_U3182) );
  AND2_X1 U22629 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19720), .ZN(
        P2_U3183) );
  AND2_X1 U22630 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19720), .ZN(
        P2_U3184) );
  AND2_X1 U22631 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19720), .ZN(
        P2_U3185) );
  AND2_X1 U22632 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19720), .ZN(
        P2_U3186) );
  AND2_X1 U22633 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19720), .ZN(
        P2_U3187) );
  AND2_X1 U22634 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19720), .ZN(
        P2_U3188) );
  AND2_X1 U22635 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19720), .ZN(
        P2_U3189) );
  AND2_X1 U22636 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19720), .ZN(
        P2_U3190) );
  AND2_X1 U22637 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19720), .ZN(
        P2_U3191) );
  AND2_X1 U22638 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19720), .ZN(
        P2_U3192) );
  AND2_X1 U22639 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19720), .ZN(
        P2_U3193) );
  AND2_X1 U22640 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19720), .ZN(
        P2_U3194) );
  AND2_X1 U22641 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19720), .ZN(
        P2_U3195) );
  AND2_X1 U22642 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19720), .ZN(
        P2_U3196) );
  AND2_X1 U22643 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19720), .ZN(
        P2_U3197) );
  AND2_X1 U22644 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19720), .ZN(
        P2_U3198) );
  AND2_X1 U22645 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19720), .ZN(
        P2_U3199) );
  AND2_X1 U22646 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19720), .ZN(
        P2_U3200) );
  AND2_X1 U22647 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19720), .ZN(P2_U3201) );
  AND2_X1 U22648 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19720), .ZN(P2_U3202) );
  AND2_X1 U22649 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19720), .ZN(P2_U3203) );
  AND2_X1 U22650 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19720), .ZN(P2_U3204) );
  AND2_X1 U22651 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19720), .ZN(P2_U3205) );
  AND2_X1 U22652 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19720), .ZN(P2_U3206) );
  AND2_X1 U22653 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19720), .ZN(P2_U3207) );
  AND2_X1 U22654 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19720), .ZN(P2_U3208) );
  NOR2_X1 U22655 ( .A1(n19722), .A2(n19721), .ZN(n19732) );
  INV_X1 U22656 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19856) );
  OR3_X1 U22657 ( .A1(n19732), .A2(n19856), .A3(n19735), .ZN(n19724) );
  AOI211_X1 U22658 ( .C1(n20639), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n19733), .B(n19858), .ZN(n19723) );
  INV_X1 U22659 ( .A(NA), .ZN(n20645) );
  NOR2_X1 U22660 ( .A1(n20645), .A2(n19726), .ZN(n19739) );
  AOI211_X1 U22661 ( .C1(n19740), .C2(n19724), .A(n19723), .B(n19739), .ZN(
        n19725) );
  INV_X1 U22662 ( .A(n19725), .ZN(P2_U3209) );
  AOI21_X1 U22663 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20639), .A(n19740), 
        .ZN(n19730) );
  NOR2_X1 U22664 ( .A1(n19856), .A2(n19730), .ZN(n19727) );
  AOI21_X1 U22665 ( .B1(n19727), .B2(n19726), .A(n19732), .ZN(n19728) );
  INV_X1 U22666 ( .A(n19845), .ZN(n19847) );
  OAI211_X1 U22667 ( .C1(n20639), .C2(n19729), .A(n19728), .B(n19847), .ZN(
        P2_U3210) );
  AOI21_X1 U22668 ( .B1(n19849), .B2(n19731), .A(n19730), .ZN(n19738) );
  AOI22_X1 U22669 ( .A1(n19856), .A2(n19733), .B1(n20645), .B2(n19732), .ZN(
        n19734) );
  AOI211_X1 U22670 ( .C1(n19856), .C2(n20639), .A(n19735), .B(n19734), .ZN(
        n19736) );
  INV_X1 U22671 ( .A(n19736), .ZN(n19737) );
  OAI21_X1 U22672 ( .B1(n19739), .B2(n19738), .A(n19737), .ZN(P2_U3211) );
  OAI222_X1 U22673 ( .A1(n19779), .A2(n13397), .B1(n19741), .B2(n19858), .C1(
        n10272), .C2(n19780), .ZN(P2_U3212) );
  OAI222_X1 U22674 ( .A1(n19779), .A2(n13817), .B1(n19742), .B2(n19858), .C1(
        n13397), .C2(n19780), .ZN(P2_U3213) );
  OAI222_X1 U22675 ( .A1(n19779), .A2(n11084), .B1(n19743), .B2(n19858), .C1(
        n13817), .C2(n19780), .ZN(P2_U3214) );
  OAI222_X1 U22676 ( .A1(n19779), .A2(n11089), .B1(n19744), .B2(n19858), .C1(
        n11084), .C2(n19780), .ZN(P2_U3215) );
  OAI222_X1 U22677 ( .A1(n19779), .A2(n14317), .B1(n19745), .B2(n19858), .C1(
        n11089), .C2(n19780), .ZN(P2_U3216) );
  OAI222_X1 U22678 ( .A1(n19779), .A2(n10797), .B1(n19746), .B2(n19858), .C1(
        n14317), .C2(n19780), .ZN(P2_U3217) );
  OAI222_X1 U22679 ( .A1(n19779), .A2(n11113), .B1(n19747), .B2(n19858), .C1(
        n10797), .C2(n19780), .ZN(P2_U3218) );
  OAI222_X1 U22680 ( .A1(n19779), .A2(n11130), .B1(n19748), .B2(n19858), .C1(
        n11113), .C2(n19780), .ZN(P2_U3219) );
  OAI222_X1 U22681 ( .A1(n19779), .A2(n11146), .B1(n19749), .B2(n19858), .C1(
        n11130), .C2(n19780), .ZN(P2_U3220) );
  OAI222_X1 U22682 ( .A1(n19779), .A2(n10812), .B1(n19750), .B2(n19858), .C1(
        n11146), .C2(n19780), .ZN(P2_U3221) );
  OAI222_X1 U22683 ( .A1(n19779), .A2(n11176), .B1(n19751), .B2(n19858), .C1(
        n10812), .C2(n19780), .ZN(P2_U3222) );
  OAI222_X1 U22684 ( .A1(n19779), .A2(n14042), .B1(n19752), .B2(n19858), .C1(
        n11176), .C2(n19780), .ZN(P2_U3223) );
  OAI222_X1 U22685 ( .A1(n19779), .A2(n11209), .B1(n19753), .B2(n19858), .C1(
        n14042), .C2(n19780), .ZN(P2_U3224) );
  OAI222_X1 U22686 ( .A1(n19779), .A2(n11227), .B1(n19754), .B2(n19858), .C1(
        n11209), .C2(n19780), .ZN(P2_U3225) );
  OAI222_X1 U22687 ( .A1(n19779), .A2(n11229), .B1(n19755), .B2(n19858), .C1(
        n11227), .C2(n19780), .ZN(P2_U3226) );
  INV_X1 U22688 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19757) );
  OAI222_X1 U22689 ( .A1(n19779), .A2(n19757), .B1(n19756), .B2(n19858), .C1(
        n11229), .C2(n19780), .ZN(P2_U3227) );
  OAI222_X1 U22690 ( .A1(n19779), .A2(n15533), .B1(n19758), .B2(n19858), .C1(
        n19757), .C2(n19780), .ZN(P2_U3228) );
  OAI222_X1 U22691 ( .A1(n19779), .A2(n19760), .B1(n19759), .B2(n19858), .C1(
        n15533), .C2(n19780), .ZN(P2_U3229) );
  OAI222_X1 U22692 ( .A1(n19779), .A2(n15509), .B1(n19761), .B2(n19858), .C1(
        n19760), .C2(n19780), .ZN(P2_U3230) );
  INV_X1 U22693 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19763) );
  OAI222_X1 U22694 ( .A1(n19779), .A2(n19763), .B1(n19762), .B2(n19858), .C1(
        n15509), .C2(n19780), .ZN(P2_U3231) );
  OAI222_X1 U22695 ( .A1(n19779), .A2(n19765), .B1(n19764), .B2(n19858), .C1(
        n19763), .C2(n19780), .ZN(P2_U3232) );
  OAI222_X1 U22696 ( .A1(n19779), .A2(n19767), .B1(n19766), .B2(n19858), .C1(
        n19765), .C2(n19780), .ZN(P2_U3233) );
  OAI222_X1 U22697 ( .A1(n19779), .A2(n19769), .B1(n19768), .B2(n19858), .C1(
        n19767), .C2(n19780), .ZN(P2_U3234) );
  INV_X1 U22698 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19771) );
  OAI222_X1 U22699 ( .A1(n19779), .A2(n19771), .B1(n19770), .B2(n19858), .C1(
        n19769), .C2(n19780), .ZN(P2_U3235) );
  OAI222_X1 U22700 ( .A1(n19779), .A2(n15223), .B1(n19772), .B2(n19858), .C1(
        n19771), .C2(n19780), .ZN(P2_U3236) );
  OAI222_X1 U22701 ( .A1(n19779), .A2(n19775), .B1(n19773), .B2(n19858), .C1(
        n15223), .C2(n19780), .ZN(P2_U3237) );
  OAI222_X1 U22702 ( .A1(n19780), .A2(n19775), .B1(n19774), .B2(n19858), .C1(
        n19776), .C2(n19779), .ZN(P2_U3238) );
  INV_X1 U22703 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19778) );
  OAI222_X1 U22704 ( .A1(n19779), .A2(n19778), .B1(n19777), .B2(n19858), .C1(
        n19776), .C2(n19780), .ZN(P2_U3239) );
  OAI222_X1 U22705 ( .A1(n19779), .A2(n14551), .B1(n20829), .B2(n19858), .C1(
        n19778), .C2(n19780), .ZN(P2_U3240) );
  OAI222_X1 U22706 ( .A1(n19779), .A2(n19782), .B1(n19781), .B2(n19858), .C1(
        n14551), .C2(n19780), .ZN(P2_U3241) );
  OAI22_X1 U22707 ( .A1(n19859), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19858), .ZN(n19783) );
  INV_X1 U22708 ( .A(n19783), .ZN(P2_U3585) );
  MUX2_X1 U22709 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19859), .Z(P2_U3586) );
  OAI22_X1 U22710 ( .A1(n19859), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19858), .ZN(n19784) );
  INV_X1 U22711 ( .A(n19784), .ZN(P2_U3587) );
  OAI22_X1 U22712 ( .A1(n19859), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19858), .ZN(n19785) );
  INV_X1 U22713 ( .A(n19785), .ZN(P2_U3588) );
  OAI21_X1 U22714 ( .B1(n19789), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19787), 
        .ZN(n19786) );
  INV_X1 U22715 ( .A(n19786), .ZN(P2_U3591) );
  OAI21_X1 U22716 ( .B1(n19789), .B2(n19788), .A(n19787), .ZN(P2_U3592) );
  INV_X1 U22717 ( .A(n19826), .ZN(n19829) );
  AND2_X1 U22718 ( .A1(n19793), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19817) );
  NAND2_X1 U22719 ( .A1(n19790), .A2(n19817), .ZN(n19807) );
  OR2_X1 U22720 ( .A1(n19816), .A2(n19791), .ZN(n19794) );
  AOI21_X1 U22721 ( .B1(n19794), .B2(n19793), .A(n19792), .ZN(n19805) );
  AOI21_X1 U22722 ( .B1(n19807), .B2(n19805), .A(n19795), .ZN(n19800) );
  NOR3_X1 U22723 ( .A1(n19798), .A2(n19797), .A3(n19796), .ZN(n19799) );
  AOI211_X1 U22724 ( .C1(n19801), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19800), 
        .B(n19799), .ZN(n19802) );
  AOI22_X1 U22725 ( .A1(n19829), .A2(n19803), .B1(n19802), .B2(n19826), .ZN(
        P2_U3602) );
  INV_X1 U22726 ( .A(n19804), .ZN(n19811) );
  INV_X1 U22727 ( .A(n19805), .ZN(n19810) );
  NOR2_X1 U22728 ( .A1(n19806), .A2(n19839), .ZN(n19809) );
  INV_X1 U22729 ( .A(n19807), .ZN(n19808) );
  AOI211_X1 U22730 ( .C1(n19811), .C2(n19810), .A(n19809), .B(n19808), .ZN(
        n19812) );
  AOI22_X1 U22731 ( .A1(n19829), .A2(n19813), .B1(n19812), .B2(n19826), .ZN(
        P2_U3603) );
  INV_X1 U22732 ( .A(n19824), .ZN(n19815) );
  NOR2_X1 U22733 ( .A1(n19815), .A2(n19814), .ZN(n19818) );
  MUX2_X1 U22734 ( .A(n19818), .B(n19817), .S(n19816), .Z(n19819) );
  AOI21_X1 U22735 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19820), .A(n19819), 
        .ZN(n19821) );
  AOI22_X1 U22736 ( .A1(n19829), .A2(n19822), .B1(n19821), .B2(n19826), .ZN(
        P2_U3604) );
  NOR2_X1 U22737 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19839), .ZN(
        n19823) );
  AOI211_X1 U22738 ( .C1(n19825), .C2(n19824), .A(n10121), .B(n19823), .ZN(
        n19827) );
  AOI22_X1 U22739 ( .A1(n19829), .A2(n19828), .B1(n19827), .B2(n19826), .ZN(
        P2_U3605) );
  INV_X1 U22740 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19830) );
  AOI22_X1 U22741 ( .A1(n19858), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19830), 
        .B2(n19859), .ZN(P2_U3608) );
  AOI22_X1 U22742 ( .A1(n19834), .A2(n19833), .B1(n19832), .B2(n19831), .ZN(
        n19836) );
  OAI21_X1 U22743 ( .B1(n19836), .B2(n10727), .A(n19835), .ZN(n19838) );
  MUX2_X1 U22744 ( .A(P2_MORE_REG_SCAN_IN), .B(n19838), .S(n19837), .Z(
        P2_U3609) );
  OAI21_X1 U22745 ( .B1(n19840), .B2(n19848), .A(n19839), .ZN(n19842) );
  OAI211_X1 U22746 ( .C1(n19849), .C2(n19843), .A(n19842), .B(n19841), .ZN(
        n19857) );
  AOI211_X1 U22747 ( .C1(P2_STATEBS16_REG_SCAN_IN), .C2(n19845), .A(n13325), 
        .B(n19844), .ZN(n19854) );
  NAND4_X1 U22748 ( .A1(n19847), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n19846), 
        .A4(n9600), .ZN(n19852) );
  OAI22_X1 U22749 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19850), .B1(n19849), 
        .B2(n19848), .ZN(n19851) );
  NAND2_X1 U22750 ( .A1(n19852), .A2(n19851), .ZN(n19853) );
  OAI21_X1 U22751 ( .B1(n19854), .B2(n19853), .A(n19857), .ZN(n19855) );
  OAI21_X1 U22752 ( .B1(n19857), .B2(n19856), .A(n19855), .ZN(P2_U3610) );
  OAI22_X1 U22753 ( .A1(n19859), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19858), .ZN(n19860) );
  INV_X1 U22754 ( .A(n19860), .ZN(P2_U3611) );
  AOI21_X1 U22755 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20653), .A(n20650), 
        .ZN(n19867) );
  INV_X1 U22756 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19861) );
  NAND2_X1 U22757 ( .A1(n20650), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20675) );
  AOI21_X1 U22758 ( .B1(n19867), .B2(n19861), .A(n20752), .ZN(P1_U2802) );
  OAI21_X1 U22759 ( .B1(n19863), .B2(n19862), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19864) );
  OAI21_X1 U22760 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n19865), .A(n19864), 
        .ZN(P1_U2803) );
  INV_X1 U22761 ( .A(n20752), .ZN(n20753) );
  NOR2_X1 U22762 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19868) );
  OAI21_X1 U22763 ( .B1(n19868), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20753), .ZN(
        n19866) );
  OAI21_X1 U22764 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20753), .A(n19866), 
        .ZN(P1_U2804) );
  NOR2_X1 U22765 ( .A1(n20752), .A2(n19867), .ZN(n20704) );
  OAI21_X1 U22766 ( .B1(BS16), .B2(n19868), .A(n20704), .ZN(n20702) );
  OAI21_X1 U22767 ( .B1(n20704), .B2(n20742), .A(n20702), .ZN(P1_U2805) );
  OAI21_X1 U22768 ( .B1(n19871), .B2(n19870), .A(n19869), .ZN(P1_U2806) );
  NOR4_X1 U22769 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19875) );
  NOR4_X1 U22770 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19874) );
  NOR4_X1 U22771 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19873) );
  NOR4_X1 U22772 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19872) );
  NAND4_X1 U22773 ( .A1(n19875), .A2(n19874), .A3(n19873), .A4(n19872), .ZN(
        n19881) );
  NOR4_X1 U22774 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19879) );
  AOI211_X1 U22775 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_30__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19878) );
  NOR4_X1 U22776 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19877) );
  NOR4_X1 U22777 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19876) );
  NAND4_X1 U22778 ( .A1(n19879), .A2(n19878), .A3(n19877), .A4(n19876), .ZN(
        n19880) );
  NOR2_X1 U22779 ( .A1(n19881), .A2(n19880), .ZN(n20736) );
  INV_X1 U22780 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19883) );
  NOR3_X1 U22781 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19884) );
  OAI21_X1 U22782 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19884), .A(n20736), .ZN(
        n19882) );
  OAI21_X1 U22783 ( .B1(n20736), .B2(n19883), .A(n19882), .ZN(P1_U2807) );
  INV_X1 U22784 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20703) );
  AOI21_X1 U22785 ( .B1(n20729), .B2(n20703), .A(n19884), .ZN(n19886) );
  INV_X1 U22786 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19885) );
  INV_X1 U22787 ( .A(n20736), .ZN(n20731) );
  AOI22_X1 U22788 ( .A1(n20736), .A2(n19886), .B1(n19885), .B2(n20731), .ZN(
        P1_U2808) );
  NAND2_X1 U22789 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19890) );
  NOR2_X1 U22790 ( .A1(n19890), .A2(n19917), .ZN(n19892) );
  INV_X1 U22791 ( .A(n19887), .ZN(n19889) );
  OAI21_X1 U22792 ( .B1(n19890), .B2(n19889), .A(n19888), .ZN(n19891) );
  INV_X1 U22793 ( .A(n19891), .ZN(n19904) );
  MUX2_X1 U22794 ( .A(n19892), .B(n19904), .S(P1_REIP_REG_7__SCAN_IN), .Z(
        n19898) );
  OAI21_X1 U22795 ( .B1(n19975), .B2(n19893), .A(n19918), .ZN(n19894) );
  AOI21_X1 U22796 ( .B1(n9585), .B2(P1_EBX_REG_7__SCAN_IN), .A(n19894), .ZN(
        n19895) );
  OAI21_X1 U22797 ( .B1(n19968), .B2(n19896), .A(n19895), .ZN(n19897) );
  AOI211_X1 U22798 ( .C1(n19900), .C2(n19899), .A(n19898), .B(n19897), .ZN(
        n19901) );
  OAI21_X1 U22799 ( .B1(n19902), .B2(n19983), .A(n19901), .ZN(P1_U2833) );
  NOR2_X1 U22800 ( .A1(n19986), .A2(n19903), .ZN(n19914) );
  NOR2_X1 U22801 ( .A1(n19926), .A2(n19917), .ZN(n19905) );
  MUX2_X1 U22802 ( .A(n19905), .B(n19904), .S(P1_REIP_REG_6__SCAN_IN), .Z(
        n19913) );
  INV_X1 U22803 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19906) );
  OAI21_X1 U22804 ( .B1(n19975), .B2(n19906), .A(n19918), .ZN(n19907) );
  AOI21_X1 U22805 ( .B1(n9585), .B2(P1_EBX_REG_6__SCAN_IN), .A(n19907), .ZN(
        n19911) );
  INV_X1 U22806 ( .A(n19984), .ZN(n19909) );
  NAND2_X1 U22807 ( .A1(n19909), .A2(n19971), .ZN(n19910) );
  NAND2_X1 U22808 ( .A1(n19911), .A2(n19910), .ZN(n19912) );
  NOR3_X1 U22809 ( .A1(n19914), .A2(n19913), .A3(n19912), .ZN(n19915) );
  OAI21_X1 U22810 ( .B1(n19916), .B2(n19983), .A(n19915), .ZN(P1_U2834) );
  INV_X1 U22811 ( .A(n19917), .ZN(n19927) );
  NAND2_X1 U22812 ( .A1(n9585), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n19919) );
  OAI211_X1 U22813 ( .C1(n19975), .C2(n19920), .A(n19919), .B(n19918), .ZN(
        n19921) );
  AOI21_X1 U22814 ( .B1(n19971), .B2(n19922), .A(n19921), .ZN(n19923) );
  OAI21_X1 U22815 ( .B1(n19924), .B2(n19976), .A(n19923), .ZN(n19925) );
  AOI221_X1 U22816 ( .B1(n19935), .B2(P1_REIP_REG_5__SCAN_IN), .C1(n19927), 
        .C2(n19926), .A(n19925), .ZN(n19928) );
  OAI21_X1 U22817 ( .B1(n19929), .B2(n19983), .A(n19928), .ZN(P1_U2835) );
  AOI22_X1 U22818 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19959), .B1(
        n19930), .B2(n13774), .ZN(n19941) );
  AOI21_X1 U22819 ( .B1(n19971), .B2(n19990), .A(n19931), .ZN(n19940) );
  INV_X1 U22820 ( .A(n19980), .ZN(n19932) );
  INV_X1 U22821 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n19996) );
  OAI22_X1 U22822 ( .A1(n19933), .A2(n19932), .B1(n19996), .B2(n19944), .ZN(
        n19934) );
  AOI21_X1 U22823 ( .B1(P1_REIP_REG_4__SCAN_IN), .B2(n19935), .A(n19934), .ZN(
        n19939) );
  OAI22_X1 U22824 ( .A1(n19993), .A2(n19976), .B1(n19936), .B2(n19983), .ZN(
        n19937) );
  INV_X1 U22825 ( .A(n19937), .ZN(n19938) );
  NAND4_X1 U22826 ( .A1(n19941), .A2(n19940), .A3(n19939), .A4(n19938), .ZN(
        P1_U2836) );
  NAND2_X1 U22827 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n19947) );
  NOR3_X1 U22828 ( .A1(n19942), .A2(n19947), .A3(P1_REIP_REG_3__SCAN_IN), .ZN(
        n19946) );
  OAI22_X1 U22829 ( .A1(n19944), .A2(n13800), .B1(n19943), .B2(n19975), .ZN(
        n19945) );
  NAND2_X1 U22830 ( .A1(n19973), .A2(n19947), .ZN(n19961) );
  NAND2_X1 U22831 ( .A1(n19961), .A2(n19948), .ZN(n19955) );
  OAI22_X1 U22832 ( .A1(n19950), .A2(n19976), .B1(n19949), .B2(n19983), .ZN(
        n19951) );
  AOI21_X1 U22833 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(n19955), .A(n19951), .ZN(
        n19952) );
  OAI211_X1 U22834 ( .C1(n19968), .C2(n19954), .A(n19953), .B(n19952), .ZN(
        P1_U2837) );
  AOI22_X1 U22835 ( .A1(n19955), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_EBX_REG_2__SCAN_IN), .B2(n9585), .ZN(n19966) );
  INV_X1 U22836 ( .A(n13476), .ZN(n20065) );
  INV_X1 U22837 ( .A(n19956), .ZN(n19957) );
  AOI22_X1 U22838 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19959), .B1(
        n19958), .B2(n19957), .ZN(n19960) );
  OAI21_X1 U22839 ( .B1(n19961), .B2(n20729), .A(n19960), .ZN(n19964) );
  NOR2_X1 U22840 ( .A1(n19962), .A2(n19976), .ZN(n19963) );
  AOI211_X1 U22841 ( .C1(n20065), .C2(n19980), .A(n19964), .B(n19963), .ZN(
        n19965) );
  OAI211_X1 U22842 ( .C1(n19968), .C2(n19967), .A(n19966), .B(n19965), .ZN(
        P1_U2838) );
  INV_X1 U22843 ( .A(n19969), .ZN(n19970) );
  AOI22_X1 U22844 ( .A1(n19971), .A2(n19970), .B1(n9585), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n19982) );
  INV_X1 U22845 ( .A(n20537), .ZN(n20538) );
  OAI22_X1 U22846 ( .A1(n19973), .A2(P1_REIP_REG_1__SCAN_IN), .B1(n19972), 
        .B2(n20729), .ZN(n19974) );
  OAI21_X1 U22847 ( .B1(n12008), .B2(n19975), .A(n19974), .ZN(n19979) );
  NOR2_X1 U22848 ( .A1(n19977), .A2(n19976), .ZN(n19978) );
  AOI211_X1 U22849 ( .C1(n19980), .C2(n20538), .A(n19979), .B(n19978), .ZN(
        n19981) );
  OAI211_X1 U22850 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19983), .A(
        n19982), .B(n19981), .ZN(P1_U2839) );
  INV_X1 U22851 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n19989) );
  OAI22_X1 U22852 ( .A1(n19986), .A2(n19992), .B1(n19985), .B2(n19984), .ZN(
        n19987) );
  INV_X1 U22853 ( .A(n19987), .ZN(n19988) );
  OAI21_X1 U22854 ( .B1(n19997), .B2(n19989), .A(n19988), .ZN(P1_U2866) );
  INV_X1 U22855 ( .A(n19990), .ZN(n19991) );
  OAI22_X1 U22856 ( .A1(n19993), .A2(n19992), .B1(n19985), .B2(n19991), .ZN(
        n19994) );
  INV_X1 U22857 ( .A(n19994), .ZN(n19995) );
  OAI21_X1 U22858 ( .B1(n19997), .B2(n19996), .A(n19995), .ZN(P1_U2868) );
  AOI22_X1 U22859 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19999) );
  OAI21_X1 U22860 ( .B1(n13392), .B2(n20019), .A(n19999), .ZN(P1_U2921) );
  INV_X1 U22861 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20001) );
  AOI22_X1 U22862 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20000) );
  OAI21_X1 U22863 ( .B1(n20001), .B2(n20019), .A(n20000), .ZN(P1_U2922) );
  AOI22_X1 U22864 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20002) );
  OAI21_X1 U22865 ( .B1(n14864), .B2(n20019), .A(n20002), .ZN(P1_U2923) );
  AOI22_X1 U22866 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20003) );
  OAI21_X1 U22867 ( .B1(n14868), .B2(n20019), .A(n20003), .ZN(P1_U2924) );
  AOI22_X1 U22868 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20004) );
  OAI21_X1 U22869 ( .B1(n20005), .B2(n20019), .A(n20004), .ZN(P1_U2925) );
  AOI22_X1 U22870 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20006) );
  OAI21_X1 U22871 ( .B1(n14339), .B2(n20019), .A(n20006), .ZN(P1_U2926) );
  AOI22_X1 U22872 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20007) );
  OAI21_X1 U22873 ( .B1(n14332), .B2(n20019), .A(n20007), .ZN(P1_U2927) );
  AOI22_X1 U22874 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20008) );
  OAI21_X1 U22875 ( .B1(n14266), .B2(n20019), .A(n20008), .ZN(P1_U2928) );
  AOI22_X1 U22876 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20009) );
  OAI21_X1 U22877 ( .B1(n12062), .B2(n20019), .A(n20009), .ZN(P1_U2929) );
  AOI22_X1 U22878 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20010) );
  OAI21_X1 U22879 ( .B1(n14068), .B2(n20019), .A(n20010), .ZN(P1_U2930) );
  AOI22_X1 U22880 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20011) );
  OAI21_X1 U22881 ( .B1(n12050), .B2(n20019), .A(n20011), .ZN(P1_U2931) );
  AOI22_X1 U22882 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20012) );
  OAI21_X1 U22883 ( .B1(n13809), .B2(n20019), .A(n20012), .ZN(P1_U2932) );
  AOI22_X1 U22884 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20013) );
  OAI21_X1 U22885 ( .B1(n12029), .B2(n20019), .A(n20013), .ZN(P1_U2933) );
  AOI22_X1 U22886 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20014) );
  OAI21_X1 U22887 ( .B1(n12002), .B2(n20019), .A(n20014), .ZN(P1_U2934) );
  AOI22_X1 U22888 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20015) );
  OAI21_X1 U22889 ( .B1(n12009), .B2(n20019), .A(n20015), .ZN(P1_U2935) );
  AOI22_X1 U22890 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20017), .B1(n20016), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20018) );
  OAI21_X1 U22891 ( .B1(n12015), .B2(n20019), .A(n20018), .ZN(P1_U2936) );
  AOI22_X1 U22892 ( .A1(n20050), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20026), .ZN(n20022) );
  INV_X1 U22893 ( .A(n20020), .ZN(n20021) );
  NAND2_X1 U22894 ( .A1(n20037), .A2(n20021), .ZN(n20039) );
  NAND2_X1 U22895 ( .A1(n20022), .A2(n20039), .ZN(P1_U2945) );
  AOI22_X1 U22896 ( .A1(n20050), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20026), .ZN(n20025) );
  INV_X1 U22897 ( .A(n20023), .ZN(n20024) );
  NAND2_X1 U22898 ( .A1(n20037), .A2(n20024), .ZN(n20041) );
  NAND2_X1 U22899 ( .A1(n20025), .A2(n20041), .ZN(P1_U2946) );
  AOI22_X1 U22900 ( .A1(n20050), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20026), .ZN(n20029) );
  INV_X1 U22901 ( .A(n20027), .ZN(n20028) );
  NAND2_X1 U22902 ( .A1(n20037), .A2(n20028), .ZN(n20043) );
  NAND2_X1 U22903 ( .A1(n20029), .A2(n20043), .ZN(P1_U2947) );
  AOI22_X1 U22904 ( .A1(n20050), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20049), .ZN(n20032) );
  INV_X1 U22905 ( .A(n20030), .ZN(n20031) );
  NAND2_X1 U22906 ( .A1(n20037), .A2(n20031), .ZN(n20045) );
  NAND2_X1 U22907 ( .A1(n20032), .A2(n20045), .ZN(P1_U2949) );
  AOI22_X1 U22908 ( .A1(n20050), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20049), .ZN(n20035) );
  INV_X1 U22909 ( .A(n20033), .ZN(n20034) );
  NAND2_X1 U22910 ( .A1(n20037), .A2(n20034), .ZN(n20047) );
  NAND2_X1 U22911 ( .A1(n20035), .A2(n20047), .ZN(P1_U2950) );
  AOI22_X1 U22912 ( .A1(n20050), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20049), .ZN(n20038) );
  NAND2_X1 U22913 ( .A1(n20037), .A2(n20036), .ZN(n20051) );
  NAND2_X1 U22914 ( .A1(n20038), .A2(n20051), .ZN(P1_U2951) );
  AOI22_X1 U22915 ( .A1(n20050), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20026), .ZN(n20040) );
  NAND2_X1 U22916 ( .A1(n20040), .A2(n20039), .ZN(P1_U2960) );
  AOI22_X1 U22917 ( .A1(n20050), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20049), .ZN(n20042) );
  NAND2_X1 U22918 ( .A1(n20042), .A2(n20041), .ZN(P1_U2961) );
  AOI22_X1 U22919 ( .A1(n20050), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20026), .ZN(n20044) );
  NAND2_X1 U22920 ( .A1(n20044), .A2(n20043), .ZN(P1_U2962) );
  AOI22_X1 U22921 ( .A1(n20050), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20049), .ZN(n20046) );
  NAND2_X1 U22922 ( .A1(n20046), .A2(n20045), .ZN(P1_U2964) );
  AOI22_X1 U22923 ( .A1(n20050), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20026), .ZN(n20048) );
  NAND2_X1 U22924 ( .A1(n20048), .A2(n20047), .ZN(P1_U2965) );
  AOI22_X1 U22925 ( .A1(n20050), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20049), .ZN(n20052) );
  NAND2_X1 U22926 ( .A1(n20052), .A2(n20051), .ZN(P1_U2966) );
  NOR2_X1 U22927 ( .A1(n11798), .A2(n20725), .ZN(P1_U3032) );
  AOI22_X1 U22928 ( .A1(DATAI_16_), .A2(n20103), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20102), .ZN(n20548) );
  INV_X1 U22929 ( .A(n20175), .ZN(n20057) );
  INV_X1 U22930 ( .A(n12013), .ZN(n20059) );
  NAND2_X1 U22931 ( .A1(n9595), .A2(n20059), .ZN(n20431) );
  INV_X1 U22932 ( .A(n20431), .ZN(n20308) );
  AOI22_X2 U22933 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20102), .B1(DATAI_24_), 
        .B2(n20103), .ZN(n20586) );
  NAND2_X1 U22934 ( .A1(n20104), .A2(n20061), .ZN(n20455) );
  NOR3_X1 U22935 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20116) );
  NAND2_X1 U22936 ( .A1(n20499), .A2(n20116), .ZN(n20105) );
  OAI22_X1 U22937 ( .A1(n20621), .A2(n20586), .B1(n20455), .B2(n20105), .ZN(
        n20062) );
  INV_X1 U22938 ( .A(n20062), .ZN(n20075) );
  INV_X1 U22939 ( .A(n20136), .ZN(n20063) );
  OAI21_X1 U22940 ( .B1(n20063), .B2(n20628), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20064) );
  NAND2_X1 U22941 ( .A1(n20064), .A2(n20718), .ZN(n20073) );
  OR2_X1 U22942 ( .A1(n20717), .A2(n20065), .ZN(n20141) );
  NOR2_X1 U22943 ( .A1(n20141), .A2(n20538), .ZN(n20070) );
  INV_X1 U22944 ( .A(n20071), .ZN(n20066) );
  NAND2_X1 U22945 ( .A1(n20066), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20536) );
  INV_X1 U22946 ( .A(n20393), .ZN(n20067) );
  OR2_X1 U22947 ( .A1(n20067), .A2(n20333), .ZN(n20213) );
  AOI22_X1 U22948 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20213), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20105), .ZN(n20068) );
  NOR2_X2 U22949 ( .A1(n20069), .A2(n20114), .ZN(n20577) );
  INV_X1 U22950 ( .A(n20070), .ZN(n20072) );
  NAND2_X1 U22951 ( .A1(n20071), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20394) );
  AOI22_X1 U22952 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20109), .B1(
        n20577), .B2(n20108), .ZN(n20074) );
  OAI211_X1 U22953 ( .C1(n20548), .C2(n20136), .A(n20075), .B(n20074), .ZN(
        P1_U3033) );
  AOI22_X1 U22954 ( .A1(DATAI_17_), .A2(n20103), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20102), .ZN(n20552) );
  AOI22_X2 U22955 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20102), .B1(DATAI_25_), 
        .B2(n20103), .ZN(n20592) );
  NAND2_X1 U22956 ( .A1(n20104), .A2(n20076), .ZN(n20467) );
  OAI22_X1 U22957 ( .A1(n20621), .A2(n20592), .B1(n20467), .B2(n20105), .ZN(
        n20077) );
  INV_X1 U22958 ( .A(n20077), .ZN(n20080) );
  NOR2_X2 U22959 ( .A1(n20078), .A2(n20114), .ZN(n20587) );
  AOI22_X1 U22960 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20109), .B1(
        n20587), .B2(n20108), .ZN(n20079) );
  OAI211_X1 U22961 ( .C1(n20552), .C2(n20136), .A(n20080), .B(n20079), .ZN(
        P1_U3034) );
  AOI22_X1 U22962 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20102), .B1(DATAI_26_), 
        .B2(n20103), .ZN(n20513) );
  NAND2_X1 U22963 ( .A1(n20104), .A2(n11477), .ZN(n20471) );
  OAI22_X1 U22964 ( .A1(n20621), .A2(n9703), .B1(n20471), .B2(n20105), .ZN(
        n20081) );
  INV_X1 U22965 ( .A(n20081), .ZN(n20084) );
  NOR2_X2 U22966 ( .A1(n20082), .A2(n20114), .ZN(n20593) );
  AOI22_X1 U22967 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20109), .B1(
        n20593), .B2(n20108), .ZN(n20083) );
  OAI211_X1 U22968 ( .C1(n20597), .C2(n20136), .A(n20084), .B(n20083), .ZN(
        P1_U3035) );
  AOI22_X1 U22969 ( .A1(DATAI_19_), .A2(n20103), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20102), .ZN(n20603) );
  OAI22_X1 U22970 ( .A1(n20621), .A2(n20517), .B1(n20475), .B2(n20105), .ZN(
        n20085) );
  INV_X1 U22971 ( .A(n20085), .ZN(n20088) );
  NOR2_X2 U22972 ( .A1(n20086), .A2(n20114), .ZN(n20598) );
  AOI22_X1 U22973 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20109), .B1(
        n20598), .B2(n20108), .ZN(n20087) );
  OAI211_X1 U22974 ( .C1(n20603), .C2(n20136), .A(n20088), .B(n20087), .ZN(
        P1_U3036) );
  AOI22_X1 U22975 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20102), .B1(DATAI_20_), 
        .B2(n20103), .ZN(n20560) );
  AOI22_X2 U22976 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20102), .B1(DATAI_28_), 
        .B2(n20103), .ZN(n20609) );
  NAND2_X1 U22977 ( .A1(n20104), .A2(n11483), .ZN(n20479) );
  OAI22_X1 U22978 ( .A1(n20621), .A2(n20609), .B1(n20479), .B2(n20105), .ZN(
        n20089) );
  INV_X1 U22979 ( .A(n20089), .ZN(n20092) );
  NOR2_X2 U22980 ( .A1(n20090), .A2(n20114), .ZN(n20604) );
  AOI22_X1 U22981 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20109), .B1(
        n20604), .B2(n20108), .ZN(n20091) );
  OAI211_X1 U22982 ( .C1(n20560), .C2(n20136), .A(n20092), .B(n20091), .ZN(
        P1_U3037) );
  AOI22_X1 U22983 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20102), .B1(DATAI_29_), 
        .B2(n20103), .ZN(n20523) );
  NAND2_X1 U22984 ( .A1(n20104), .A2(n20093), .ZN(n20483) );
  OAI22_X1 U22985 ( .A1(n20621), .A2(n20523), .B1(n20483), .B2(n20105), .ZN(
        n20094) );
  INV_X1 U22986 ( .A(n20094), .ZN(n20097) );
  NOR2_X2 U22987 ( .A1(n20095), .A2(n20114), .ZN(n20610) );
  AOI22_X1 U22988 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20109), .B1(
        n20610), .B2(n20108), .ZN(n20096) );
  OAI211_X1 U22989 ( .C1(n20615), .C2(n20136), .A(n20097), .B(n20096), .ZN(
        P1_U3038) );
  AOI22_X1 U22990 ( .A1(DATAI_22_), .A2(n20103), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20102), .ZN(n20622) );
  AOI22_X1 U22991 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20102), .B1(DATAI_30_), 
        .B2(n20103), .ZN(n20526) );
  NAND2_X1 U22992 ( .A1(n20104), .A2(n9843), .ZN(n20487) );
  OAI22_X1 U22993 ( .A1(n20621), .A2(n9707), .B1(n20487), .B2(n20105), .ZN(
        n20098) );
  INV_X1 U22994 ( .A(n20098), .ZN(n20101) );
  NOR2_X2 U22995 ( .A1(n20099), .A2(n20114), .ZN(n20616) );
  AOI22_X1 U22996 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20109), .B1(
        n20616), .B2(n20108), .ZN(n20100) );
  OAI211_X1 U22997 ( .C1(n9705), .C2(n20136), .A(n20101), .B(n20100), .ZN(
        P1_U3039) );
  AOI22_X1 U22998 ( .A1(DATAI_31_), .A2(n20103), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20102), .ZN(n20633) );
  NAND2_X1 U22999 ( .A1(n20104), .A2(n12000), .ZN(n20492) );
  OAI22_X1 U23000 ( .A1(n20621), .A2(n9709), .B1(n20492), .B2(n20105), .ZN(
        n20106) );
  INV_X1 U23001 ( .A(n20106), .ZN(n20111) );
  NOR2_X2 U23002 ( .A1(n20114), .A2(n20107), .ZN(n20624) );
  AOI22_X1 U23003 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20109), .B1(
        n20624), .B2(n20108), .ZN(n20110) );
  OAI211_X1 U23004 ( .C1(n20571), .C2(n20136), .A(n20111), .B(n20110), .ZN(
        P1_U3040) );
  INV_X1 U23005 ( .A(n20141), .ZN(n20178) );
  INV_X1 U23006 ( .A(n20502), .ZN(n20359) );
  INV_X1 U23007 ( .A(n20116), .ZN(n20112) );
  NOR2_X1 U23008 ( .A1(n20499), .A2(n20112), .ZN(n20131) );
  AOI21_X1 U23009 ( .B1(n20178), .B2(n20359), .A(n20131), .ZN(n20113) );
  OAI22_X1 U23010 ( .A1(n20113), .A2(n20573), .B1(n20112), .B2(n12409), .ZN(
        n20132) );
  AOI22_X1 U23011 ( .A1(n20132), .A2(n20577), .B1(n20578), .B2(n20131), .ZN(
        n20118) );
  OAI21_X1 U23012 ( .B1(n20175), .B2(n20742), .A(n20113), .ZN(n20115) );
  OAI221_X1 U23013 ( .B1(n20718), .B2(n20116), .C1(n20573), .C2(n20115), .A(
        n20581), .ZN(n20133) );
  INV_X1 U23014 ( .A(n20548), .ZN(n20583) );
  AOI22_X1 U23015 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20133), .B1(
        n20138), .B2(n20583), .ZN(n20117) );
  OAI211_X1 U23016 ( .C1(n20586), .C2(n20136), .A(n20118), .B(n20117), .ZN(
        P1_U3041) );
  AOI22_X1 U23017 ( .A1(n20132), .A2(n20587), .B1(n20588), .B2(n20131), .ZN(
        n20120) );
  INV_X1 U23018 ( .A(n20552), .ZN(n20589) );
  AOI22_X1 U23019 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20133), .B1(
        n20138), .B2(n20589), .ZN(n20119) );
  OAI211_X1 U23020 ( .C1(n20592), .C2(n20136), .A(n20120), .B(n20119), .ZN(
        P1_U3042) );
  AOI22_X1 U23021 ( .A1(n20132), .A2(n20593), .B1(n20594), .B2(n20131), .ZN(
        n20122) );
  INV_X1 U23022 ( .A(n20597), .ZN(n20510) );
  AOI22_X1 U23023 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20133), .B1(
        n20138), .B2(n20510), .ZN(n20121) );
  OAI211_X1 U23024 ( .C1(n9703), .C2(n20136), .A(n20122), .B(n20121), .ZN(
        P1_U3043) );
  AOI22_X1 U23025 ( .A1(n20132), .A2(n20598), .B1(n20599), .B2(n20131), .ZN(
        n20124) );
  INV_X1 U23026 ( .A(n20603), .ZN(n20514) );
  AOI22_X1 U23027 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20133), .B1(
        n20138), .B2(n20514), .ZN(n20123) );
  OAI211_X1 U23028 ( .C1(n20517), .C2(n20136), .A(n20124), .B(n20123), .ZN(
        P1_U3044) );
  AOI22_X1 U23029 ( .A1(n20132), .A2(n20604), .B1(n20605), .B2(n20131), .ZN(
        n20126) );
  INV_X1 U23030 ( .A(n20560), .ZN(n20606) );
  AOI22_X1 U23031 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20133), .B1(
        n20138), .B2(n20606), .ZN(n20125) );
  OAI211_X1 U23032 ( .C1(n20609), .C2(n20136), .A(n20126), .B(n20125), .ZN(
        P1_U3045) );
  AOI22_X1 U23033 ( .A1(n20132), .A2(n20610), .B1(n20611), .B2(n20131), .ZN(
        n20128) );
  INV_X1 U23034 ( .A(n20615), .ZN(n20520) );
  AOI22_X1 U23035 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20133), .B1(
        n20138), .B2(n20520), .ZN(n20127) );
  OAI211_X1 U23036 ( .C1(n20523), .C2(n20136), .A(n20128), .B(n20127), .ZN(
        P1_U3046) );
  AOI22_X1 U23037 ( .A1(n20132), .A2(n20616), .B1(n20617), .B2(n20131), .ZN(
        n20130) );
  AOI22_X1 U23038 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20133), .B1(
        n20138), .B2(n9704), .ZN(n20129) );
  OAI211_X1 U23039 ( .C1(n9707), .C2(n20136), .A(n20130), .B(n20129), .ZN(
        P1_U3047) );
  AOI22_X1 U23040 ( .A1(n20132), .A2(n20624), .B1(n20626), .B2(n20131), .ZN(
        n20135) );
  INV_X1 U23041 ( .A(n20571), .ZN(n20627) );
  AOI22_X1 U23042 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20133), .B1(
        n20138), .B2(n20627), .ZN(n20134) );
  OAI211_X1 U23043 ( .C1(n9709), .C2(n20136), .A(n20135), .B(n20134), .ZN(
        P1_U3048) );
  NAND2_X1 U23044 ( .A1(n9595), .A2(n12013), .ZN(n20385) );
  NAND3_X1 U23045 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20727), .A3(
        n11803), .ZN(n20181) );
  OR2_X1 U23046 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20181), .ZN(
        n20166) );
  OAI22_X1 U23047 ( .A1(n20167), .A2(n20586), .B1(n20166), .B2(n20455), .ZN(
        n20137) );
  INV_X1 U23048 ( .A(n20137), .ZN(n20147) );
  INV_X1 U23049 ( .A(n20205), .ZN(n20139) );
  OAI21_X1 U23050 ( .B1(n20139), .B2(n20138), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20140) );
  NAND2_X1 U23051 ( .A1(n20140), .A2(n20718), .ZN(n20145) );
  NOR2_X1 U23052 ( .A1(n20141), .A2(n20537), .ZN(n20143) );
  OR2_X1 U23053 ( .A1(n20393), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20272) );
  AND2_X1 U23054 ( .A1(n20272), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20268) );
  AOI21_X1 U23055 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20166), .A(n20268), 
        .ZN(n20142) );
  OAI211_X1 U23056 ( .C1(n20145), .C2(n20143), .A(n20391), .B(n20142), .ZN(
        n20170) );
  INV_X1 U23057 ( .A(n20143), .ZN(n20144) );
  AOI22_X1 U23058 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20170), .B1(
        n20577), .B2(n20169), .ZN(n20146) );
  OAI211_X1 U23059 ( .C1(n20548), .C2(n20205), .A(n20147), .B(n20146), .ZN(
        P1_U3049) );
  OAI22_X1 U23060 ( .A1(n20205), .A2(n20552), .B1(n20467), .B2(n20166), .ZN(
        n20148) );
  INV_X1 U23061 ( .A(n20148), .ZN(n20150) );
  AOI22_X1 U23062 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20170), .B1(
        n20587), .B2(n20169), .ZN(n20149) );
  OAI211_X1 U23063 ( .C1(n20592), .C2(n20167), .A(n20150), .B(n20149), .ZN(
        P1_U3050) );
  OAI22_X1 U23064 ( .A1(n20205), .A2(n20597), .B1(n20166), .B2(n20471), .ZN(
        n20151) );
  INV_X1 U23065 ( .A(n20151), .ZN(n20153) );
  AOI22_X1 U23066 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20170), .B1(
        n20593), .B2(n20169), .ZN(n20152) );
  OAI211_X1 U23067 ( .C1(n9703), .C2(n20167), .A(n20153), .B(n20152), .ZN(
        P1_U3051) );
  OAI22_X1 U23068 ( .A1(n20205), .A2(n20603), .B1(n20475), .B2(n20166), .ZN(
        n20154) );
  INV_X1 U23069 ( .A(n20154), .ZN(n20156) );
  AOI22_X1 U23070 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20170), .B1(
        n20598), .B2(n20169), .ZN(n20155) );
  OAI211_X1 U23071 ( .C1(n20517), .C2(n20167), .A(n20156), .B(n20155), .ZN(
        P1_U3052) );
  OAI22_X1 U23072 ( .A1(n20205), .A2(n20560), .B1(n20479), .B2(n20166), .ZN(
        n20157) );
  INV_X1 U23073 ( .A(n20157), .ZN(n20159) );
  AOI22_X1 U23074 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20170), .B1(
        n20604), .B2(n20169), .ZN(n20158) );
  OAI211_X1 U23075 ( .C1(n20609), .C2(n20167), .A(n20159), .B(n20158), .ZN(
        P1_U3053) );
  OAI22_X1 U23076 ( .A1(n20205), .A2(n20615), .B1(n20483), .B2(n20166), .ZN(
        n20160) );
  INV_X1 U23077 ( .A(n20160), .ZN(n20162) );
  AOI22_X1 U23078 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20170), .B1(
        n20610), .B2(n20169), .ZN(n20161) );
  OAI211_X1 U23079 ( .C1(n20523), .C2(n20167), .A(n20162), .B(n20161), .ZN(
        P1_U3054) );
  OAI22_X1 U23080 ( .A1(n20167), .A2(n9707), .B1(n20487), .B2(n20166), .ZN(
        n20163) );
  INV_X1 U23081 ( .A(n20163), .ZN(n20165) );
  AOI22_X1 U23082 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20170), .B1(
        n20616), .B2(n20169), .ZN(n20164) );
  OAI211_X1 U23083 ( .C1(n9705), .C2(n20205), .A(n20165), .B(n20164), .ZN(
        P1_U3055) );
  OAI22_X1 U23084 ( .A1(n20167), .A2(n9709), .B1(n20166), .B2(n20492), .ZN(
        n20168) );
  INV_X1 U23085 ( .A(n20168), .ZN(n20172) );
  AOI22_X1 U23086 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20170), .B1(
        n20624), .B2(n20169), .ZN(n20171) );
  OAI211_X1 U23087 ( .C1(n20571), .C2(n20205), .A(n20172), .B(n20171), .ZN(
        P1_U3056) );
  INV_X1 U23088 ( .A(n20424), .ZN(n20173) );
  NAND2_X1 U23089 ( .A1(n20173), .A2(n20727), .ZN(n20204) );
  OAI22_X1 U23090 ( .A1(n20205), .A2(n20586), .B1(n20204), .B2(n20455), .ZN(
        n20174) );
  INV_X1 U23091 ( .A(n20174), .ZN(n20185) );
  OAI21_X1 U23092 ( .B1(n20175), .B2(n20428), .A(n20718), .ZN(n20183) );
  AND2_X1 U23093 ( .A1(n20176), .A2(n9594), .ZN(n20572) );
  INV_X1 U23094 ( .A(n20204), .ZN(n20177) );
  AOI21_X1 U23095 ( .B1(n20178), .B2(n20572), .A(n20177), .ZN(n20182) );
  INV_X1 U23096 ( .A(n20182), .ZN(n20180) );
  NAND2_X1 U23097 ( .A1(n20573), .A2(n20181), .ZN(n20179) );
  OAI211_X1 U23098 ( .C1(n20183), .C2(n20180), .A(n20581), .B(n20179), .ZN(
        n20208) );
  OAI22_X1 U23099 ( .A1(n20183), .A2(n20182), .B1(n12409), .B2(n20181), .ZN(
        n20207) );
  AOI22_X1 U23100 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20208), .B1(
        n20577), .B2(n20207), .ZN(n20184) );
  OAI211_X1 U23101 ( .C1(n20548), .C2(n20230), .A(n20185), .B(n20184), .ZN(
        P1_U3057) );
  OAI22_X1 U23102 ( .A1(n20205), .A2(n20592), .B1(n20204), .B2(n20467), .ZN(
        n20186) );
  INV_X1 U23103 ( .A(n20186), .ZN(n20188) );
  AOI22_X1 U23104 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20208), .B1(
        n20587), .B2(n20207), .ZN(n20187) );
  OAI211_X1 U23105 ( .C1(n20552), .C2(n20230), .A(n20188), .B(n20187), .ZN(
        P1_U3058) );
  OAI22_X1 U23106 ( .A1(n20205), .A2(n9703), .B1(n20204), .B2(n20471), .ZN(
        n20189) );
  INV_X1 U23107 ( .A(n20189), .ZN(n20191) );
  AOI22_X1 U23108 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20208), .B1(
        n20593), .B2(n20207), .ZN(n20190) );
  OAI211_X1 U23109 ( .C1(n20597), .C2(n20230), .A(n20191), .B(n20190), .ZN(
        P1_U3059) );
  OAI22_X1 U23110 ( .A1(n20230), .A2(n20603), .B1(n20475), .B2(n20204), .ZN(
        n20192) );
  INV_X1 U23111 ( .A(n20192), .ZN(n20194) );
  AOI22_X1 U23112 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20208), .B1(
        n20598), .B2(n20207), .ZN(n20193) );
  OAI211_X1 U23113 ( .C1(n20517), .C2(n20205), .A(n20194), .B(n20193), .ZN(
        P1_U3060) );
  OAI22_X1 U23114 ( .A1(n20230), .A2(n20560), .B1(n20204), .B2(n20479), .ZN(
        n20195) );
  INV_X1 U23115 ( .A(n20195), .ZN(n20197) );
  AOI22_X1 U23116 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20208), .B1(
        n20604), .B2(n20207), .ZN(n20196) );
  OAI211_X1 U23117 ( .C1(n20609), .C2(n20205), .A(n20197), .B(n20196), .ZN(
        P1_U3061) );
  OAI22_X1 U23118 ( .A1(n20230), .A2(n20615), .B1(n20204), .B2(n20483), .ZN(
        n20198) );
  INV_X1 U23119 ( .A(n20198), .ZN(n20200) );
  AOI22_X1 U23120 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20208), .B1(
        n20610), .B2(n20207), .ZN(n20199) );
  OAI211_X1 U23121 ( .C1(n20523), .C2(n20205), .A(n20200), .B(n20199), .ZN(
        P1_U3062) );
  OAI22_X1 U23122 ( .A1(n20230), .A2(n9705), .B1(n20204), .B2(n20487), .ZN(
        n20201) );
  INV_X1 U23123 ( .A(n20201), .ZN(n20203) );
  AOI22_X1 U23124 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20208), .B1(
        n20616), .B2(n20207), .ZN(n20202) );
  OAI211_X1 U23125 ( .C1(n9707), .C2(n20205), .A(n20203), .B(n20202), .ZN(
        P1_U3063) );
  OAI22_X1 U23126 ( .A1(n20205), .A2(n9709), .B1(n20204), .B2(n20492), .ZN(
        n20206) );
  INV_X1 U23127 ( .A(n20206), .ZN(n20210) );
  AOI22_X1 U23128 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20208), .B1(
        n20624), .B2(n20207), .ZN(n20209) );
  OAI211_X1 U23129 ( .C1(n20571), .C2(n20230), .A(n20210), .B(n20209), .ZN(
        P1_U3064) );
  NOR3_X1 U23130 ( .A1(n11803), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20242) );
  INV_X1 U23131 ( .A(n20242), .ZN(n20239) );
  NOR2_X1 U23132 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20239), .ZN(
        n20234) );
  NOR2_X1 U23133 ( .A1(n13476), .A2(n20212), .ZN(n20302) );
  NAND2_X1 U23134 ( .A1(n20302), .A2(n20537), .ZN(n20214) );
  OAI22_X1 U23135 ( .A1(n20214), .A2(n20573), .B1(n20536), .B2(n20213), .ZN(
        n20233) );
  AOI22_X1 U23136 ( .A1(n20578), .A2(n20234), .B1(n20577), .B2(n20233), .ZN(
        n20219) );
  OAI21_X1 U23137 ( .B1(n20235), .B2(n20254), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20215) );
  NAND2_X1 U23138 ( .A1(n20215), .A2(n20214), .ZN(n20217) );
  INV_X1 U23139 ( .A(n20586), .ZN(n20545) );
  AOI22_X1 U23140 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20236), .B1(
        n20235), .B2(n20545), .ZN(n20218) );
  OAI211_X1 U23141 ( .C1(n20548), .C2(n20265), .A(n20219), .B(n20218), .ZN(
        P1_U3065) );
  AOI22_X1 U23142 ( .A1(n20588), .A2(n20234), .B1(n20587), .B2(n20233), .ZN(
        n20221) );
  AOI22_X1 U23143 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20236), .B1(
        n20254), .B2(n20589), .ZN(n20220) );
  OAI211_X1 U23144 ( .C1(n20592), .C2(n20230), .A(n20221), .B(n20220), .ZN(
        P1_U3066) );
  AOI22_X1 U23145 ( .A1(n20594), .A2(n20234), .B1(n20593), .B2(n20233), .ZN(
        n20223) );
  AOI22_X1 U23146 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20236), .B1(
        n20254), .B2(n20510), .ZN(n20222) );
  OAI211_X1 U23147 ( .C1(n9703), .C2(n20230), .A(n20223), .B(n20222), .ZN(
        P1_U3067) );
  AOI22_X1 U23148 ( .A1(n20599), .A2(n20234), .B1(n20598), .B2(n20233), .ZN(
        n20225) );
  AOI22_X1 U23149 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20236), .B1(
        n20254), .B2(n20514), .ZN(n20224) );
  OAI211_X1 U23150 ( .C1(n20517), .C2(n20230), .A(n20225), .B(n20224), .ZN(
        P1_U3068) );
  AOI22_X1 U23151 ( .A1(n20605), .A2(n20234), .B1(n20604), .B2(n20233), .ZN(
        n20227) );
  AOI22_X1 U23152 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20236), .B1(
        n20254), .B2(n20606), .ZN(n20226) );
  OAI211_X1 U23153 ( .C1(n20609), .C2(n20230), .A(n20227), .B(n20226), .ZN(
        P1_U3069) );
  AOI22_X1 U23154 ( .A1(n20611), .A2(n20234), .B1(n20610), .B2(n20233), .ZN(
        n20229) );
  AOI22_X1 U23155 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20236), .B1(
        n20254), .B2(n20520), .ZN(n20228) );
  OAI211_X1 U23156 ( .C1(n20523), .C2(n20230), .A(n20229), .B(n20228), .ZN(
        P1_U3070) );
  AOI22_X1 U23157 ( .A1(n20617), .A2(n20234), .B1(n20616), .B2(n20233), .ZN(
        n20232) );
  AOI22_X1 U23158 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20236), .B1(
        n20235), .B2(n9706), .ZN(n20231) );
  OAI211_X1 U23159 ( .C1(n9705), .C2(n20265), .A(n20232), .B(n20231), .ZN(
        P1_U3071) );
  AOI22_X1 U23160 ( .A1(n20626), .A2(n20234), .B1(n20624), .B2(n20233), .ZN(
        n20238) );
  AOI22_X1 U23161 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20236), .B1(
        n20235), .B2(n9708), .ZN(n20237) );
  OAI211_X1 U23162 ( .C1(n20571), .C2(n20265), .A(n20238), .B(n20237), .ZN(
        P1_U3072) );
  NOR2_X1 U23163 ( .A1(n20499), .A2(n20239), .ZN(n20259) );
  AOI21_X1 U23164 ( .B1(n20302), .B2(n20359), .A(n20259), .ZN(n20240) );
  OAI22_X1 U23165 ( .A1(n20240), .A2(n20573), .B1(n20239), .B2(n12409), .ZN(
        n20260) );
  AOI22_X1 U23166 ( .A1(n20577), .A2(n20260), .B1(n20578), .B2(n20259), .ZN(
        n20245) );
  OAI21_X1 U23167 ( .B1(n20305), .B2(n20742), .A(n20240), .ZN(n20241) );
  OAI221_X1 U23168 ( .B1(n20718), .B2(n20242), .C1(n20573), .C2(n20241), .A(
        n20581), .ZN(n20262) );
  INV_X1 U23169 ( .A(n20505), .ZN(n20243) );
  INV_X1 U23170 ( .A(n20301), .ZN(n20261) );
  AOI22_X1 U23171 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20262), .B1(
        n20261), .B2(n20583), .ZN(n20244) );
  OAI211_X1 U23172 ( .C1(n20586), .C2(n20265), .A(n20245), .B(n20244), .ZN(
        P1_U3073) );
  AOI22_X1 U23173 ( .A1(n20587), .A2(n20260), .B1(n20588), .B2(n20259), .ZN(
        n20247) );
  AOI22_X1 U23174 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20262), .B1(
        n20261), .B2(n20589), .ZN(n20246) );
  OAI211_X1 U23175 ( .C1(n20592), .C2(n20265), .A(n20247), .B(n20246), .ZN(
        P1_U3074) );
  AOI22_X1 U23176 ( .A1(n20593), .A2(n20260), .B1(n20594), .B2(n20259), .ZN(
        n20249) );
  AOI22_X1 U23177 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20262), .B1(
        n20261), .B2(n20510), .ZN(n20248) );
  OAI211_X1 U23178 ( .C1(n9703), .C2(n20265), .A(n20249), .B(n20248), .ZN(
        P1_U3075) );
  AOI22_X1 U23179 ( .A1(n20598), .A2(n20260), .B1(n20599), .B2(n20259), .ZN(
        n20251) );
  AOI22_X1 U23180 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20262), .B1(
        n20261), .B2(n20514), .ZN(n20250) );
  OAI211_X1 U23181 ( .C1(n20517), .C2(n20265), .A(n20251), .B(n20250), .ZN(
        P1_U3076) );
  AOI22_X1 U23182 ( .A1(n20604), .A2(n20260), .B1(n20605), .B2(n20259), .ZN(
        n20253) );
  INV_X1 U23183 ( .A(n20609), .ZN(n20557) );
  AOI22_X1 U23184 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20262), .B1(
        n20254), .B2(n20557), .ZN(n20252) );
  OAI211_X1 U23185 ( .C1(n20560), .C2(n20301), .A(n20253), .B(n20252), .ZN(
        P1_U3077) );
  AOI22_X1 U23186 ( .A1(n20610), .A2(n20260), .B1(n20611), .B2(n20259), .ZN(
        n20256) );
  INV_X1 U23187 ( .A(n20523), .ZN(n20612) );
  AOI22_X1 U23188 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20262), .B1(
        n20254), .B2(n20612), .ZN(n20255) );
  OAI211_X1 U23189 ( .C1(n20615), .C2(n20301), .A(n20256), .B(n20255), .ZN(
        P1_U3078) );
  AOI22_X1 U23190 ( .A1(n20616), .A2(n20260), .B1(n20617), .B2(n20259), .ZN(
        n20258) );
  AOI22_X1 U23191 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20262), .B1(
        n20261), .B2(n9704), .ZN(n20257) );
  OAI211_X1 U23192 ( .C1(n9707), .C2(n20265), .A(n20258), .B(n20257), .ZN(
        P1_U3079) );
  AOI22_X1 U23193 ( .A1(n20624), .A2(n20260), .B1(n20626), .B2(n20259), .ZN(
        n20264) );
  AOI22_X1 U23194 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20262), .B1(
        n20261), .B2(n20627), .ZN(n20263) );
  OAI211_X1 U23195 ( .C1(n9709), .C2(n20265), .A(n20264), .B(n20263), .ZN(
        P1_U3080) );
  INV_X1 U23196 ( .A(n20385), .ZN(n20533) );
  NOR2_X1 U23197 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20303), .ZN(
        n20270) );
  INV_X1 U23198 ( .A(n20270), .ZN(n20295) );
  OAI22_X1 U23199 ( .A1(n20319), .A2(n20548), .B1(n20455), .B2(n20295), .ZN(
        n20266) );
  INV_X1 U23200 ( .A(n20266), .ZN(n20276) );
  NAND2_X1 U23201 ( .A1(n20319), .A2(n20301), .ZN(n20267) );
  AOI21_X1 U23202 ( .B1(n20267), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20573), 
        .ZN(n20271) );
  NAND2_X1 U23203 ( .A1(n20302), .A2(n20538), .ZN(n20273) );
  AOI21_X1 U23204 ( .B1(n20271), .B2(n20273), .A(n20268), .ZN(n20269) );
  OAI211_X1 U23205 ( .C1(n20270), .C2(n20338), .A(n20543), .B(n20269), .ZN(
        n20298) );
  INV_X1 U23206 ( .A(n20271), .ZN(n20274) );
  AOI22_X1 U23207 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20298), .B1(
        n20577), .B2(n20297), .ZN(n20275) );
  OAI211_X1 U23208 ( .C1(n20586), .C2(n20301), .A(n20276), .B(n20275), .ZN(
        P1_U3081) );
  OAI22_X1 U23209 ( .A1(n20301), .A2(n20592), .B1(n20467), .B2(n20295), .ZN(
        n20277) );
  INV_X1 U23210 ( .A(n20277), .ZN(n20279) );
  AOI22_X1 U23211 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20298), .B1(
        n20587), .B2(n20297), .ZN(n20278) );
  OAI211_X1 U23212 ( .C1(n20552), .C2(n20319), .A(n20279), .B(n20278), .ZN(
        P1_U3082) );
  OAI22_X1 U23213 ( .A1(n20319), .A2(n20597), .B1(n20471), .B2(n20295), .ZN(
        n20280) );
  INV_X1 U23214 ( .A(n20280), .ZN(n20282) );
  AOI22_X1 U23215 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20298), .B1(
        n20593), .B2(n20297), .ZN(n20281) );
  OAI211_X1 U23216 ( .C1(n9703), .C2(n20301), .A(n20282), .B(n20281), .ZN(
        P1_U3083) );
  OAI22_X1 U23217 ( .A1(n20301), .A2(n20517), .B1(n20475), .B2(n20295), .ZN(
        n20283) );
  INV_X1 U23218 ( .A(n20283), .ZN(n20285) );
  AOI22_X1 U23219 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20298), .B1(
        n20598), .B2(n20297), .ZN(n20284) );
  OAI211_X1 U23220 ( .C1(n20603), .C2(n20319), .A(n20285), .B(n20284), .ZN(
        P1_U3084) );
  OAI22_X1 U23221 ( .A1(n20319), .A2(n20560), .B1(n20479), .B2(n20295), .ZN(
        n20286) );
  INV_X1 U23222 ( .A(n20286), .ZN(n20288) );
  AOI22_X1 U23223 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20298), .B1(
        n20604), .B2(n20297), .ZN(n20287) );
  OAI211_X1 U23224 ( .C1(n20609), .C2(n20301), .A(n20288), .B(n20287), .ZN(
        P1_U3085) );
  OAI22_X1 U23225 ( .A1(n20319), .A2(n20615), .B1(n20483), .B2(n20295), .ZN(
        n20289) );
  INV_X1 U23226 ( .A(n20289), .ZN(n20291) );
  AOI22_X1 U23227 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20298), .B1(
        n20610), .B2(n20297), .ZN(n20290) );
  OAI211_X1 U23228 ( .C1(n20523), .C2(n20301), .A(n20291), .B(n20290), .ZN(
        P1_U3086) );
  OAI22_X1 U23229 ( .A1(n20301), .A2(n9707), .B1(n20487), .B2(n20295), .ZN(
        n20292) );
  INV_X1 U23230 ( .A(n20292), .ZN(n20294) );
  AOI22_X1 U23231 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20298), .B1(
        n20616), .B2(n20297), .ZN(n20293) );
  OAI211_X1 U23232 ( .C1(n9705), .C2(n20319), .A(n20294), .B(n20293), .ZN(
        P1_U3087) );
  OAI22_X1 U23233 ( .A1(n20319), .A2(n20571), .B1(n20492), .B2(n20295), .ZN(
        n20296) );
  INV_X1 U23234 ( .A(n20296), .ZN(n20300) );
  AOI22_X1 U23235 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20298), .B1(
        n20624), .B2(n20297), .ZN(n20299) );
  OAI211_X1 U23236 ( .C1(n9709), .C2(n20301), .A(n20300), .B(n20299), .ZN(
        P1_U3088) );
  AOI21_X1 U23237 ( .B1(n20302), .B2(n20572), .A(n20324), .ZN(n20304) );
  OAI22_X1 U23238 ( .A1(n20304), .A2(n20573), .B1(n20303), .B2(n12409), .ZN(
        n20325) );
  AOI22_X1 U23239 ( .A1(n20577), .A2(n20325), .B1(n20578), .B2(n20324), .ZN(
        n20310) );
  INV_X1 U23240 ( .A(n20303), .ZN(n20307) );
  OAI21_X1 U23241 ( .B1(n20305), .B2(n20428), .A(n20304), .ZN(n20306) );
  OAI221_X1 U23242 ( .B1(n20718), .B2(n20307), .C1(n20573), .C2(n20306), .A(
        n20581), .ZN(n20327) );
  AOI22_X1 U23243 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20327), .B1(
        n20355), .B2(n20583), .ZN(n20309) );
  OAI211_X1 U23244 ( .C1(n20586), .C2(n20319), .A(n20310), .B(n20309), .ZN(
        P1_U3089) );
  AOI22_X1 U23245 ( .A1(n20587), .A2(n20325), .B1(n20588), .B2(n20324), .ZN(
        n20312) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20327), .B1(
        n20355), .B2(n20589), .ZN(n20311) );
  OAI211_X1 U23247 ( .C1(n20592), .C2(n20319), .A(n20312), .B(n20311), .ZN(
        P1_U3090) );
  AOI22_X1 U23248 ( .A1(n20593), .A2(n20325), .B1(n20594), .B2(n20324), .ZN(
        n20314) );
  INV_X1 U23249 ( .A(n20319), .ZN(n20326) );
  AOI22_X1 U23250 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20327), .B1(
        n20326), .B2(n9702), .ZN(n20313) );
  OAI211_X1 U23251 ( .C1(n20597), .C2(n20330), .A(n20314), .B(n20313), .ZN(
        P1_U3091) );
  AOI22_X1 U23252 ( .A1(n20598), .A2(n20325), .B1(n20599), .B2(n20324), .ZN(
        n20316) );
  INV_X1 U23253 ( .A(n20517), .ZN(n20600) );
  AOI22_X1 U23254 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20327), .B1(
        n20326), .B2(n20600), .ZN(n20315) );
  OAI211_X1 U23255 ( .C1(n20603), .C2(n20330), .A(n20316), .B(n20315), .ZN(
        P1_U3092) );
  AOI22_X1 U23256 ( .A1(n20604), .A2(n20325), .B1(n20605), .B2(n20324), .ZN(
        n20318) );
  AOI22_X1 U23257 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20327), .B1(
        n20355), .B2(n20606), .ZN(n20317) );
  OAI211_X1 U23258 ( .C1(n20609), .C2(n20319), .A(n20318), .B(n20317), .ZN(
        P1_U3093) );
  AOI22_X1 U23259 ( .A1(n20610), .A2(n20325), .B1(n20611), .B2(n20324), .ZN(
        n20321) );
  AOI22_X1 U23260 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20327), .B1(
        n20326), .B2(n20612), .ZN(n20320) );
  OAI211_X1 U23261 ( .C1(n20615), .C2(n20330), .A(n20321), .B(n20320), .ZN(
        P1_U3094) );
  AOI22_X1 U23262 ( .A1(n20616), .A2(n20325), .B1(n20617), .B2(n20324), .ZN(
        n20323) );
  AOI22_X1 U23263 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20327), .B1(
        n20326), .B2(n9706), .ZN(n20322) );
  OAI211_X1 U23264 ( .C1(n9705), .C2(n20330), .A(n20323), .B(n20322), .ZN(
        P1_U3095) );
  AOI22_X1 U23265 ( .A1(n20624), .A2(n20325), .B1(n20626), .B2(n20324), .ZN(
        n20329) );
  AOI22_X1 U23266 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20327), .B1(
        n20326), .B2(n9708), .ZN(n20328) );
  OAI211_X1 U23267 ( .C1(n20571), .C2(n20330), .A(n20329), .B(n20328), .ZN(
        P1_U3096) );
  INV_X1 U23268 ( .A(n11999), .ZN(n20331) );
  INV_X1 U23269 ( .A(n20432), .ZN(n20332) );
  NAND2_X1 U23270 ( .A1(n20717), .A2(n13476), .ZN(n20389) );
  INV_X1 U23271 ( .A(n20389), .ZN(n20425) );
  NOR3_X1 U23272 ( .A1(n20727), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20363) );
  INV_X1 U23273 ( .A(n20363), .ZN(n20360) );
  NOR2_X1 U23274 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20360), .ZN(
        n20353) );
  AOI21_X1 U23275 ( .B1(n20425), .B2(n20537), .A(n20353), .ZN(n20335) );
  NAND2_X1 U23276 ( .A1(n20333), .A2(n20393), .ZN(n20462) );
  OAI22_X1 U23277 ( .A1(n20335), .A2(n20573), .B1(n20462), .B2(n20394), .ZN(
        n20354) );
  AOI22_X1 U23278 ( .A1(n20354), .A2(n20577), .B1(n20578), .B2(n20353), .ZN(
        n20340) );
  INV_X1 U23279 ( .A(n20384), .ZN(n20334) );
  OAI21_X1 U23280 ( .B1(n20334), .B2(n20355), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20336) );
  NAND2_X1 U23281 ( .A1(n20336), .A2(n20335), .ZN(n20337) );
  AOI22_X1 U23282 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20356), .B1(
        n20355), .B2(n20545), .ZN(n20339) );
  OAI211_X1 U23283 ( .C1(n20548), .C2(n20384), .A(n20340), .B(n20339), .ZN(
        P1_U3097) );
  AOI22_X1 U23284 ( .A1(n20354), .A2(n20587), .B1(n20588), .B2(n20353), .ZN(
        n20342) );
  INV_X1 U23285 ( .A(n20592), .ZN(n20549) );
  AOI22_X1 U23286 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20356), .B1(
        n20355), .B2(n20549), .ZN(n20341) );
  OAI211_X1 U23287 ( .C1(n20552), .C2(n20384), .A(n20342), .B(n20341), .ZN(
        P1_U3098) );
  AOI22_X1 U23288 ( .A1(n20354), .A2(n20593), .B1(n20594), .B2(n20353), .ZN(
        n20344) );
  AOI22_X1 U23289 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20356), .B1(
        n20355), .B2(n9702), .ZN(n20343) );
  OAI211_X1 U23290 ( .C1(n20597), .C2(n20384), .A(n20344), .B(n20343), .ZN(
        P1_U3099) );
  AOI22_X1 U23291 ( .A1(n20354), .A2(n20598), .B1(n20599), .B2(n20353), .ZN(
        n20346) );
  AOI22_X1 U23292 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20356), .B1(
        n20355), .B2(n20600), .ZN(n20345) );
  OAI211_X1 U23293 ( .C1(n20603), .C2(n20384), .A(n20346), .B(n20345), .ZN(
        P1_U3100) );
  AOI22_X1 U23294 ( .A1(n20354), .A2(n20604), .B1(n20605), .B2(n20353), .ZN(
        n20348) );
  AOI22_X1 U23295 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20356), .B1(
        n20355), .B2(n20557), .ZN(n20347) );
  OAI211_X1 U23296 ( .C1(n20560), .C2(n20384), .A(n20348), .B(n20347), .ZN(
        P1_U3101) );
  AOI22_X1 U23297 ( .A1(n20354), .A2(n20610), .B1(n20611), .B2(n20353), .ZN(
        n20350) );
  AOI22_X1 U23298 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20356), .B1(
        n20355), .B2(n20612), .ZN(n20349) );
  OAI211_X1 U23299 ( .C1(n20615), .C2(n20384), .A(n20350), .B(n20349), .ZN(
        P1_U3102) );
  AOI22_X1 U23300 ( .A1(n20354), .A2(n20616), .B1(n20617), .B2(n20353), .ZN(
        n20352) );
  AOI22_X1 U23301 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20356), .B1(
        n20355), .B2(n9706), .ZN(n20351) );
  OAI211_X1 U23302 ( .C1(n9705), .C2(n20384), .A(n20352), .B(n20351), .ZN(
        P1_U3103) );
  AOI22_X1 U23303 ( .A1(n20354), .A2(n20624), .B1(n20626), .B2(n20353), .ZN(
        n20358) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20356), .B1(
        n20355), .B2(n9708), .ZN(n20357) );
  OAI211_X1 U23305 ( .C1(n20571), .C2(n20384), .A(n20358), .B(n20357), .ZN(
        P1_U3104) );
  NOR2_X1 U23306 ( .A1(n20499), .A2(n20360), .ZN(n20378) );
  AOI21_X1 U23307 ( .B1(n20425), .B2(n20359), .A(n20378), .ZN(n20361) );
  OAI22_X1 U23308 ( .A1(n20361), .A2(n20573), .B1(n20360), .B2(n12409), .ZN(
        n20379) );
  AOI22_X1 U23309 ( .A1(n20379), .A2(n20577), .B1(n20578), .B2(n20378), .ZN(
        n20365) );
  OAI21_X1 U23310 ( .B1(n20432), .B2(n20742), .A(n20361), .ZN(n20362) );
  OAI221_X1 U23311 ( .B1(n20718), .B2(n20363), .C1(n20573), .C2(n20362), .A(
        n20581), .ZN(n20381) );
  AOI22_X1 U23312 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20381), .B1(
        n20380), .B2(n20583), .ZN(n20364) );
  OAI211_X1 U23313 ( .C1(n20586), .C2(n20384), .A(n20365), .B(n20364), .ZN(
        P1_U3105) );
  AOI22_X1 U23314 ( .A1(n20379), .A2(n20587), .B1(n20588), .B2(n20378), .ZN(
        n20367) );
  AOI22_X1 U23315 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20381), .B1(
        n20380), .B2(n20589), .ZN(n20366) );
  OAI211_X1 U23316 ( .C1(n20592), .C2(n20384), .A(n20367), .B(n20366), .ZN(
        P1_U3106) );
  AOI22_X1 U23317 ( .A1(n20379), .A2(n20593), .B1(n20594), .B2(n20378), .ZN(
        n20369) );
  AOI22_X1 U23318 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20381), .B1(
        n20380), .B2(n20510), .ZN(n20368) );
  OAI211_X1 U23319 ( .C1(n9703), .C2(n20384), .A(n20369), .B(n20368), .ZN(
        P1_U3107) );
  AOI22_X1 U23320 ( .A1(n20379), .A2(n20598), .B1(n20599), .B2(n20378), .ZN(
        n20371) );
  AOI22_X1 U23321 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20381), .B1(
        n20380), .B2(n20514), .ZN(n20370) );
  OAI211_X1 U23322 ( .C1(n20517), .C2(n20384), .A(n20371), .B(n20370), .ZN(
        P1_U3108) );
  AOI22_X1 U23323 ( .A1(n20379), .A2(n20604), .B1(n20605), .B2(n20378), .ZN(
        n20373) );
  AOI22_X1 U23324 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20381), .B1(
        n20380), .B2(n20606), .ZN(n20372) );
  OAI211_X1 U23325 ( .C1(n20609), .C2(n20384), .A(n20373), .B(n20372), .ZN(
        P1_U3109) );
  AOI22_X1 U23326 ( .A1(n20379), .A2(n20610), .B1(n20611), .B2(n20378), .ZN(
        n20375) );
  AOI22_X1 U23327 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20381), .B1(
        n20380), .B2(n20520), .ZN(n20374) );
  OAI211_X1 U23328 ( .C1(n20523), .C2(n20384), .A(n20375), .B(n20374), .ZN(
        P1_U3110) );
  AOI22_X1 U23329 ( .A1(n20379), .A2(n20616), .B1(n20617), .B2(n20378), .ZN(
        n20377) );
  AOI22_X1 U23330 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20381), .B1(
        n20380), .B2(n9704), .ZN(n20376) );
  OAI211_X1 U23331 ( .C1(n9707), .C2(n20384), .A(n20377), .B(n20376), .ZN(
        P1_U3111) );
  AOI22_X1 U23332 ( .A1(n20379), .A2(n20624), .B1(n20626), .B2(n20378), .ZN(
        n20383) );
  AOI22_X1 U23333 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20381), .B1(
        n20380), .B2(n20627), .ZN(n20382) );
  OAI211_X1 U23334 ( .C1(n9709), .C2(n20384), .A(n20383), .B(n20382), .ZN(
        P1_U3112) );
  NOR3_X1 U23335 ( .A1(n20727), .A2(n20386), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20430) );
  NAND2_X1 U23336 ( .A1(n20499), .A2(n20430), .ZN(n20417) );
  OAI22_X1 U23337 ( .A1(n20423), .A2(n20586), .B1(n20455), .B2(n20417), .ZN(
        n20387) );
  INV_X1 U23338 ( .A(n20387), .ZN(n20398) );
  AOI21_X1 U23339 ( .B1(n20448), .B2(n20423), .A(n20742), .ZN(n20388) );
  NOR2_X1 U23340 ( .A1(n20388), .A2(n20573), .ZN(n20392) );
  OR2_X1 U23341 ( .A1(n20389), .A2(n20537), .ZN(n20395) );
  AOI22_X1 U23342 ( .A1(n20392), .A2(n20395), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20417), .ZN(n20390) );
  OAI21_X1 U23343 ( .B1(n20727), .B2(n20393), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n20542) );
  NAND3_X1 U23344 ( .A1(n20391), .A2(n20390), .A3(n20542), .ZN(n20420) );
  INV_X1 U23345 ( .A(n20392), .ZN(n20396) );
  OR2_X1 U23346 ( .A1(n20393), .A2(n20727), .ZN(n20535) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20420), .B1(
        n20577), .B2(n20419), .ZN(n20397) );
  OAI211_X1 U23348 ( .C1(n20548), .C2(n20448), .A(n20398), .B(n20397), .ZN(
        P1_U3113) );
  OAI22_X1 U23349 ( .A1(n20423), .A2(n20592), .B1(n20467), .B2(n20417), .ZN(
        n20399) );
  INV_X1 U23350 ( .A(n20399), .ZN(n20401) );
  AOI22_X1 U23351 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20420), .B1(
        n20587), .B2(n20419), .ZN(n20400) );
  OAI211_X1 U23352 ( .C1(n20552), .C2(n20448), .A(n20401), .B(n20400), .ZN(
        P1_U3114) );
  OAI22_X1 U23353 ( .A1(n20448), .A2(n20597), .B1(n20471), .B2(n20417), .ZN(
        n20402) );
  INV_X1 U23354 ( .A(n20402), .ZN(n20404) );
  AOI22_X1 U23355 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20420), .B1(
        n20593), .B2(n20419), .ZN(n20403) );
  OAI211_X1 U23356 ( .C1(n9703), .C2(n20423), .A(n20404), .B(n20403), .ZN(
        P1_U3115) );
  OAI22_X1 U23357 ( .A1(n20423), .A2(n20517), .B1(n20475), .B2(n20417), .ZN(
        n20405) );
  INV_X1 U23358 ( .A(n20405), .ZN(n20407) );
  AOI22_X1 U23359 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20420), .B1(
        n20598), .B2(n20419), .ZN(n20406) );
  OAI211_X1 U23360 ( .C1(n20603), .C2(n20448), .A(n20407), .B(n20406), .ZN(
        P1_U3116) );
  OAI22_X1 U23361 ( .A1(n20423), .A2(n20609), .B1(n20479), .B2(n20417), .ZN(
        n20408) );
  INV_X1 U23362 ( .A(n20408), .ZN(n20410) );
  AOI22_X1 U23363 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20420), .B1(
        n20604), .B2(n20419), .ZN(n20409) );
  OAI211_X1 U23364 ( .C1(n20560), .C2(n20448), .A(n20410), .B(n20409), .ZN(
        P1_U3117) );
  OAI22_X1 U23365 ( .A1(n20448), .A2(n20615), .B1(n20483), .B2(n20417), .ZN(
        n20411) );
  INV_X1 U23366 ( .A(n20411), .ZN(n20413) );
  AOI22_X1 U23367 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20420), .B1(
        n20610), .B2(n20419), .ZN(n20412) );
  OAI211_X1 U23368 ( .C1(n20523), .C2(n20423), .A(n20413), .B(n20412), .ZN(
        P1_U3118) );
  OAI22_X1 U23369 ( .A1(n20448), .A2(n9705), .B1(n20487), .B2(n20417), .ZN(
        n20414) );
  INV_X1 U23370 ( .A(n20414), .ZN(n20416) );
  AOI22_X1 U23371 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20420), .B1(
        n20616), .B2(n20419), .ZN(n20415) );
  OAI211_X1 U23372 ( .C1(n9707), .C2(n20423), .A(n20416), .B(n20415), .ZN(
        P1_U3119) );
  OAI22_X1 U23373 ( .A1(n20448), .A2(n20571), .B1(n20492), .B2(n20417), .ZN(
        n20418) );
  INV_X1 U23374 ( .A(n20418), .ZN(n20422) );
  AOI22_X1 U23375 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20420), .B1(
        n20624), .B2(n20419), .ZN(n20421) );
  OAI211_X1 U23376 ( .C1(n9709), .C2(n20423), .A(n20422), .B(n20421), .ZN(
        P1_U3120) );
  NOR2_X1 U23377 ( .A1(n20424), .A2(n20727), .ZN(n20449) );
  AOI21_X1 U23378 ( .B1(n20425), .B2(n20572), .A(n20449), .ZN(n20427) );
  INV_X1 U23379 ( .A(n20430), .ZN(n20426) );
  OAI22_X1 U23380 ( .A1(n20427), .A2(n20573), .B1(n20426), .B2(n12409), .ZN(
        n20450) );
  AOI22_X1 U23381 ( .A1(n20450), .A2(n20577), .B1(n20578), .B2(n20449), .ZN(
        n20434) );
  OAI21_X1 U23382 ( .B1(n20432), .B2(n20428), .A(n20427), .ZN(n20429) );
  OAI221_X1 U23383 ( .B1(n20718), .B2(n20430), .C1(n20573), .C2(n20429), .A(
        n20581), .ZN(n20452) );
  INV_X1 U23384 ( .A(n20498), .ZN(n20445) );
  AOI22_X1 U23385 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20452), .B1(
        n20445), .B2(n20583), .ZN(n20433) );
  OAI211_X1 U23386 ( .C1(n20586), .C2(n20448), .A(n20434), .B(n20433), .ZN(
        P1_U3121) );
  AOI22_X1 U23387 ( .A1(n20450), .A2(n20587), .B1(n20588), .B2(n20449), .ZN(
        n20436) );
  INV_X1 U23388 ( .A(n20448), .ZN(n20451) );
  AOI22_X1 U23389 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20452), .B1(
        n20451), .B2(n20549), .ZN(n20435) );
  OAI211_X1 U23390 ( .C1(n20552), .C2(n20498), .A(n20436), .B(n20435), .ZN(
        P1_U3122) );
  AOI22_X1 U23391 ( .A1(n20450), .A2(n20593), .B1(n20594), .B2(n20449), .ZN(
        n20438) );
  AOI22_X1 U23392 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20452), .B1(
        n20451), .B2(n9702), .ZN(n20437) );
  OAI211_X1 U23393 ( .C1(n20597), .C2(n20498), .A(n20438), .B(n20437), .ZN(
        P1_U3123) );
  AOI22_X1 U23394 ( .A1(n20450), .A2(n20598), .B1(n20599), .B2(n20449), .ZN(
        n20440) );
  AOI22_X1 U23395 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20452), .B1(
        n20445), .B2(n20514), .ZN(n20439) );
  OAI211_X1 U23396 ( .C1(n20517), .C2(n20448), .A(n20440), .B(n20439), .ZN(
        P1_U3124) );
  AOI22_X1 U23397 ( .A1(n20450), .A2(n20604), .B1(n20605), .B2(n20449), .ZN(
        n20442) );
  AOI22_X1 U23398 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20452), .B1(
        n20445), .B2(n20606), .ZN(n20441) );
  OAI211_X1 U23399 ( .C1(n20609), .C2(n20448), .A(n20442), .B(n20441), .ZN(
        P1_U3125) );
  AOI22_X1 U23400 ( .A1(n20450), .A2(n20610), .B1(n20611), .B2(n20449), .ZN(
        n20444) );
  AOI22_X1 U23401 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20452), .B1(
        n20451), .B2(n20612), .ZN(n20443) );
  OAI211_X1 U23402 ( .C1(n20615), .C2(n20498), .A(n20444), .B(n20443), .ZN(
        P1_U3126) );
  AOI22_X1 U23403 ( .A1(n20450), .A2(n20616), .B1(n20617), .B2(n20449), .ZN(
        n20447) );
  AOI22_X1 U23404 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20452), .B1(
        n20445), .B2(n9704), .ZN(n20446) );
  OAI211_X1 U23405 ( .C1(n9707), .C2(n20448), .A(n20447), .B(n20446), .ZN(
        P1_U3127) );
  AOI22_X1 U23406 ( .A1(n20450), .A2(n20624), .B1(n20626), .B2(n20449), .ZN(
        n20454) );
  AOI22_X1 U23407 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20452), .B1(
        n20451), .B2(n9708), .ZN(n20453) );
  OAI211_X1 U23408 ( .C1(n20571), .C2(n20498), .A(n20454), .B(n20453), .ZN(
        P1_U3128) );
  NOR3_X1 U23409 ( .A1(n11803), .A2(n20727), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20503) );
  NAND2_X1 U23410 ( .A1(n20499), .A2(n20503), .ZN(n20491) );
  OAI22_X1 U23411 ( .A1(n20532), .A2(n20548), .B1(n20455), .B2(n20491), .ZN(
        n20456) );
  INV_X1 U23412 ( .A(n20456), .ZN(n20466) );
  INV_X1 U23413 ( .A(n20462), .ZN(n20460) );
  AOI21_X1 U23414 ( .B1(n20498), .B2(n20532), .A(n20742), .ZN(n20457) );
  NOR2_X1 U23415 ( .A1(n20457), .A2(n20573), .ZN(n20461) );
  NOR2_X1 U23416 ( .A1(n13476), .A2(n20458), .ZN(n20539) );
  NAND2_X1 U23417 ( .A1(n20539), .A2(n20537), .ZN(n20463) );
  AOI22_X1 U23418 ( .A1(n20461), .A2(n20463), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20491), .ZN(n20459) );
  INV_X1 U23419 ( .A(n20461), .ZN(n20464) );
  AOI22_X1 U23420 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20495), .B1(
        n20577), .B2(n20494), .ZN(n20465) );
  OAI211_X1 U23421 ( .C1(n20586), .C2(n20498), .A(n20466), .B(n20465), .ZN(
        P1_U3129) );
  OAI22_X1 U23422 ( .A1(n20532), .A2(n20552), .B1(n20467), .B2(n20491), .ZN(
        n20468) );
  INV_X1 U23423 ( .A(n20468), .ZN(n20470) );
  AOI22_X1 U23424 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20495), .B1(
        n20587), .B2(n20494), .ZN(n20469) );
  OAI211_X1 U23425 ( .C1(n20592), .C2(n20498), .A(n20470), .B(n20469), .ZN(
        P1_U3130) );
  OAI22_X1 U23426 ( .A1(n20532), .A2(n20597), .B1(n20471), .B2(n20491), .ZN(
        n20472) );
  INV_X1 U23427 ( .A(n20472), .ZN(n20474) );
  AOI22_X1 U23428 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20495), .B1(
        n20593), .B2(n20494), .ZN(n20473) );
  OAI211_X1 U23429 ( .C1(n9703), .C2(n20498), .A(n20474), .B(n20473), .ZN(
        P1_U3131) );
  OAI22_X1 U23430 ( .A1(n20532), .A2(n20603), .B1(n20475), .B2(n20491), .ZN(
        n20476) );
  INV_X1 U23431 ( .A(n20476), .ZN(n20478) );
  AOI22_X1 U23432 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20495), .B1(
        n20598), .B2(n20494), .ZN(n20477) );
  OAI211_X1 U23433 ( .C1(n20517), .C2(n20498), .A(n20478), .B(n20477), .ZN(
        P1_U3132) );
  OAI22_X1 U23434 ( .A1(n20532), .A2(n20560), .B1(n20479), .B2(n20491), .ZN(
        n20480) );
  INV_X1 U23435 ( .A(n20480), .ZN(n20482) );
  AOI22_X1 U23436 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20495), .B1(
        n20604), .B2(n20494), .ZN(n20481) );
  OAI211_X1 U23437 ( .C1(n20609), .C2(n20498), .A(n20482), .B(n20481), .ZN(
        P1_U3133) );
  OAI22_X1 U23438 ( .A1(n20532), .A2(n20615), .B1(n20483), .B2(n20491), .ZN(
        n20484) );
  INV_X1 U23439 ( .A(n20484), .ZN(n20486) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20495), .B1(
        n20610), .B2(n20494), .ZN(n20485) );
  OAI211_X1 U23441 ( .C1(n20523), .C2(n20498), .A(n20486), .B(n20485), .ZN(
        P1_U3134) );
  OAI22_X1 U23442 ( .A1(n20532), .A2(n9705), .B1(n20487), .B2(n20491), .ZN(
        n20488) );
  INV_X1 U23443 ( .A(n20488), .ZN(n20490) );
  AOI22_X1 U23444 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20495), .B1(
        n20616), .B2(n20494), .ZN(n20489) );
  OAI211_X1 U23445 ( .C1(n9707), .C2(n20498), .A(n20490), .B(n20489), .ZN(
        P1_U3135) );
  OAI22_X1 U23446 ( .A1(n20532), .A2(n20571), .B1(n20492), .B2(n20491), .ZN(
        n20493) );
  INV_X1 U23447 ( .A(n20493), .ZN(n20497) );
  AOI22_X1 U23448 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20495), .B1(
        n20624), .B2(n20494), .ZN(n20496) );
  OAI211_X1 U23449 ( .C1(n9709), .C2(n20498), .A(n20497), .B(n20496), .ZN(
        P1_U3136) );
  INV_X1 U23450 ( .A(n20503), .ZN(n20500) );
  NOR2_X1 U23451 ( .A1(n20499), .A2(n20500), .ZN(n20528) );
  NAND2_X1 U23452 ( .A1(n20539), .A2(n20718), .ZN(n20576) );
  INV_X1 U23453 ( .A(n20528), .ZN(n20501) );
  OAI222_X1 U23454 ( .A1(n20576), .A2(n20502), .B1(n20501), .B2(n20573), .C1(
        n12409), .C2(n20500), .ZN(n20527) );
  AOI22_X1 U23455 ( .A1(n20578), .A2(n20528), .B1(n20527), .B2(n20577), .ZN(
        n20507) );
  NAND2_X1 U23456 ( .A1(n20534), .A2(n10125), .ZN(n20724) );
  INV_X1 U23457 ( .A(n20724), .ZN(n20504) );
  AOI22_X1 U23458 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20529), .B1(
        n20567), .B2(n20583), .ZN(n20506) );
  OAI211_X1 U23459 ( .C1(n20586), .C2(n20532), .A(n20507), .B(n20506), .ZN(
        P1_U3137) );
  AOI22_X1 U23460 ( .A1(n20588), .A2(n20528), .B1(n20527), .B2(n20587), .ZN(
        n20509) );
  AOI22_X1 U23461 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20529), .B1(
        n20567), .B2(n20589), .ZN(n20508) );
  OAI211_X1 U23462 ( .C1(n20592), .C2(n20532), .A(n20509), .B(n20508), .ZN(
        P1_U3138) );
  AOI22_X1 U23463 ( .A1(n20594), .A2(n20528), .B1(n20527), .B2(n20593), .ZN(
        n20512) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20529), .B1(
        n20567), .B2(n20510), .ZN(n20511) );
  OAI211_X1 U23465 ( .C1(n9703), .C2(n20532), .A(n20512), .B(n20511), .ZN(
        P1_U3139) );
  AOI22_X1 U23466 ( .A1(n20599), .A2(n20528), .B1(n20527), .B2(n20598), .ZN(
        n20516) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20529), .B1(
        n20567), .B2(n20514), .ZN(n20515) );
  OAI211_X1 U23468 ( .C1(n20517), .C2(n20532), .A(n20516), .B(n20515), .ZN(
        P1_U3140) );
  AOI22_X1 U23469 ( .A1(n20605), .A2(n20528), .B1(n20527), .B2(n20604), .ZN(
        n20519) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20529), .B1(
        n20567), .B2(n20606), .ZN(n20518) );
  OAI211_X1 U23471 ( .C1(n20609), .C2(n20532), .A(n20519), .B(n20518), .ZN(
        P1_U3141) );
  AOI22_X1 U23472 ( .A1(n20611), .A2(n20528), .B1(n20527), .B2(n20610), .ZN(
        n20522) );
  AOI22_X1 U23473 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20529), .B1(
        n20567), .B2(n20520), .ZN(n20521) );
  OAI211_X1 U23474 ( .C1(n20523), .C2(n20532), .A(n20522), .B(n20521), .ZN(
        P1_U3142) );
  AOI22_X1 U23475 ( .A1(n20617), .A2(n20528), .B1(n20527), .B2(n20616), .ZN(
        n20525) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20529), .B1(
        n20567), .B2(n9704), .ZN(n20524) );
  OAI211_X1 U23477 ( .C1(n9707), .C2(n20532), .A(n20525), .B(n20524), .ZN(
        P1_U3143) );
  AOI22_X1 U23478 ( .A1(n20626), .A2(n20528), .B1(n20624), .B2(n20527), .ZN(
        n20531) );
  AOI22_X1 U23479 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20529), .B1(
        n20567), .B2(n20627), .ZN(n20530) );
  OAI211_X1 U23480 ( .C1(n9709), .C2(n20532), .A(n20531), .B(n20530), .ZN(
        P1_U3144) );
  NOR2_X1 U23481 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20579), .ZN(
        n20566) );
  OAI22_X1 U23482 ( .A1(n20576), .A2(n20537), .B1(n20536), .B2(n20535), .ZN(
        n20565) );
  AOI22_X1 U23483 ( .A1(n20578), .A2(n20566), .B1(n20577), .B2(n20565), .ZN(
        n20547) );
  INV_X1 U23484 ( .A(n20632), .ZN(n20618) );
  OAI21_X1 U23485 ( .B1(n20618), .B2(n20567), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20541) );
  NAND2_X1 U23486 ( .A1(n20539), .A2(n20538), .ZN(n20540) );
  AOI21_X1 U23487 ( .B1(n20541), .B2(n20540), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20544) );
  AOI22_X1 U23488 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20568), .B1(
        n20567), .B2(n20545), .ZN(n20546) );
  OAI211_X1 U23489 ( .C1(n20548), .C2(n20632), .A(n20547), .B(n20546), .ZN(
        P1_U3145) );
  AOI22_X1 U23490 ( .A1(n20588), .A2(n20566), .B1(n20587), .B2(n20565), .ZN(
        n20551) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20568), .B1(
        n20567), .B2(n20549), .ZN(n20550) );
  OAI211_X1 U23492 ( .C1(n20552), .C2(n20632), .A(n20551), .B(n20550), .ZN(
        P1_U3146) );
  AOI22_X1 U23493 ( .A1(n20594), .A2(n20566), .B1(n20593), .B2(n20565), .ZN(
        n20554) );
  AOI22_X1 U23494 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20568), .B1(
        n20567), .B2(n9702), .ZN(n20553) );
  OAI211_X1 U23495 ( .C1(n20597), .C2(n20632), .A(n20554), .B(n20553), .ZN(
        P1_U3147) );
  AOI22_X1 U23496 ( .A1(n20599), .A2(n20566), .B1(n20598), .B2(n20565), .ZN(
        n20556) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20568), .B1(
        n20567), .B2(n20600), .ZN(n20555) );
  OAI211_X1 U23498 ( .C1(n20603), .C2(n20632), .A(n20556), .B(n20555), .ZN(
        P1_U3148) );
  AOI22_X1 U23499 ( .A1(n20605), .A2(n20566), .B1(n20604), .B2(n20565), .ZN(
        n20559) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20568), .B1(
        n20567), .B2(n20557), .ZN(n20558) );
  OAI211_X1 U23501 ( .C1(n20560), .C2(n20632), .A(n20559), .B(n20558), .ZN(
        P1_U3149) );
  AOI22_X1 U23502 ( .A1(n20611), .A2(n20566), .B1(n20610), .B2(n20565), .ZN(
        n20562) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20568), .B1(
        n20567), .B2(n20612), .ZN(n20561) );
  OAI211_X1 U23504 ( .C1(n20615), .C2(n20632), .A(n20562), .B(n20561), .ZN(
        P1_U3150) );
  AOI22_X1 U23505 ( .A1(n20617), .A2(n20566), .B1(n20616), .B2(n20565), .ZN(
        n20564) );
  AOI22_X1 U23506 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20568), .B1(
        n20567), .B2(n9706), .ZN(n20563) );
  OAI211_X1 U23507 ( .C1(n9705), .C2(n20632), .A(n20564), .B(n20563), .ZN(
        P1_U3151) );
  AOI22_X1 U23508 ( .A1(n20626), .A2(n20566), .B1(n20624), .B2(n20565), .ZN(
        n20570) );
  AOI22_X1 U23509 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20568), .B1(
        n20567), .B2(n9708), .ZN(n20569) );
  OAI211_X1 U23510 ( .C1(n20571), .C2(n20632), .A(n20570), .B(n20569), .ZN(
        P1_U3152) );
  INV_X1 U23511 ( .A(n20572), .ZN(n20575) );
  INV_X1 U23512 ( .A(n20625), .ZN(n20574) );
  OAI222_X1 U23513 ( .A1(n20576), .A2(n20575), .B1(n20574), .B2(n20573), .C1(
        n12409), .C2(n20579), .ZN(n20623) );
  AOI22_X1 U23514 ( .A1(n20578), .A2(n20625), .B1(n20623), .B2(n20577), .ZN(
        n20585) );
  OAI21_X1 U23515 ( .B1(n20580), .B2(n20712), .A(n20579), .ZN(n20582) );
  NAND2_X1 U23516 ( .A1(n20582), .A2(n20581), .ZN(n20629) );
  AOI22_X1 U23517 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20583), .ZN(n20584) );
  OAI211_X1 U23518 ( .C1(n20586), .C2(n20632), .A(n20585), .B(n20584), .ZN(
        P1_U3153) );
  AOI22_X1 U23519 ( .A1(n20588), .A2(n20625), .B1(n20623), .B2(n20587), .ZN(
        n20591) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20589), .ZN(n20590) );
  OAI211_X1 U23521 ( .C1(n20592), .C2(n20632), .A(n20591), .B(n20590), .ZN(
        P1_U3154) );
  AOI22_X1 U23522 ( .A1(n20594), .A2(n20625), .B1(n20623), .B2(n20593), .ZN(
        n20596) );
  AOI22_X1 U23523 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20629), .B1(
        n20618), .B2(n9702), .ZN(n20595) );
  OAI211_X1 U23524 ( .C1(n20597), .C2(n20621), .A(n20596), .B(n20595), .ZN(
        P1_U3155) );
  AOI22_X1 U23525 ( .A1(n20599), .A2(n20625), .B1(n20623), .B2(n20598), .ZN(
        n20602) );
  AOI22_X1 U23526 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20629), .B1(
        n20618), .B2(n20600), .ZN(n20601) );
  OAI211_X1 U23527 ( .C1(n20603), .C2(n20621), .A(n20602), .B(n20601), .ZN(
        P1_U3156) );
  AOI22_X1 U23528 ( .A1(n20605), .A2(n20625), .B1(n20623), .B2(n20604), .ZN(
        n20608) );
  AOI22_X1 U23529 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20606), .ZN(n20607) );
  OAI211_X1 U23530 ( .C1(n20609), .C2(n20632), .A(n20608), .B(n20607), .ZN(
        P1_U3157) );
  AOI22_X1 U23531 ( .A1(n20611), .A2(n20625), .B1(n20623), .B2(n20610), .ZN(
        n20614) );
  AOI22_X1 U23532 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20629), .B1(
        n20618), .B2(n20612), .ZN(n20613) );
  OAI211_X1 U23533 ( .C1(n20615), .C2(n20621), .A(n20614), .B(n20613), .ZN(
        P1_U3158) );
  AOI22_X1 U23534 ( .A1(n20617), .A2(n20625), .B1(n20623), .B2(n20616), .ZN(
        n20620) );
  AOI22_X1 U23535 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20629), .B1(
        n20618), .B2(n9706), .ZN(n20619) );
  OAI211_X1 U23536 ( .C1(n9705), .C2(n20621), .A(n20620), .B(n20619), .ZN(
        P1_U3159) );
  AOI22_X1 U23537 ( .A1(n20626), .A2(n20625), .B1(n20624), .B2(n20623), .ZN(
        n20631) );
  AOI22_X1 U23538 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20629), .B1(
        n20628), .B2(n20627), .ZN(n20630) );
  OAI211_X1 U23539 ( .C1(n9709), .C2(n20632), .A(n20631), .B(n20630), .ZN(
        P1_U3160) );
  OAI221_X1 U23540 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20636), .C1(n12409), 
        .C2(n20635), .A(n20634), .ZN(P1_U3163) );
  AND2_X1 U23541 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20637), .ZN(
        P1_U3164) );
  AND2_X1 U23542 ( .A1(n20637), .A2(P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(
        P1_U3165) );
  AND2_X1 U23543 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20637), .ZN(
        P1_U3166) );
  AND2_X1 U23544 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20637), .ZN(
        P1_U3167) );
  AND2_X1 U23545 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20637), .ZN(
        P1_U3168) );
  AND2_X1 U23546 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20637), .ZN(
        P1_U3169) );
  AND2_X1 U23547 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20637), .ZN(
        P1_U3170) );
  AND2_X1 U23548 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20637), .ZN(
        P1_U3171) );
  AND2_X1 U23549 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20637), .ZN(
        P1_U3172) );
  AND2_X1 U23550 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20637), .ZN(
        P1_U3173) );
  AND2_X1 U23551 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20637), .ZN(
        P1_U3174) );
  AND2_X1 U23552 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20637), .ZN(
        P1_U3175) );
  AND2_X1 U23553 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20637), .ZN(
        P1_U3176) );
  AND2_X1 U23554 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20637), .ZN(
        P1_U3177) );
  AND2_X1 U23555 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20637), .ZN(
        P1_U3178) );
  AND2_X1 U23556 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20637), .ZN(
        P1_U3179) );
  AND2_X1 U23557 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20637), .ZN(
        P1_U3180) );
  AND2_X1 U23558 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20637), .ZN(
        P1_U3181) );
  AND2_X1 U23559 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20637), .ZN(
        P1_U3182) );
  AND2_X1 U23560 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20637), .ZN(
        P1_U3183) );
  AND2_X1 U23561 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20637), .ZN(
        P1_U3184) );
  AND2_X1 U23562 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20637), .ZN(
        P1_U3185) );
  AND2_X1 U23563 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20637), .ZN(P1_U3186) );
  AND2_X1 U23564 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20637), .ZN(P1_U3187) );
  AND2_X1 U23565 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20637), .ZN(P1_U3188) );
  AND2_X1 U23566 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20637), .ZN(P1_U3189) );
  AND2_X1 U23567 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20637), .ZN(P1_U3190) );
  AND2_X1 U23568 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20637), .ZN(P1_U3191) );
  AND2_X1 U23569 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20637), .ZN(P1_U3192) );
  AND2_X1 U23570 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20637), .ZN(P1_U3193) );
  AND2_X1 U23571 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20638), .ZN(n20652) );
  INV_X1 U23572 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20750) );
  INV_X1 U23573 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20640) );
  OAI22_X1 U23574 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20645), .B1(n20640), 
        .B2(n20639), .ZN(n20641) );
  NOR3_X1 U23575 ( .A1(n20642), .A2(n20750), .A3(n20641), .ZN(n20643) );
  OAI22_X1 U23576 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20652), .B1(n20752), 
        .B2(n20643), .ZN(P1_U3194) );
  NOR2_X1 U23577 ( .A1(n20650), .A2(n20750), .ZN(n20644) );
  OAI22_X1 U23578 ( .A1(n20646), .A2(n20645), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20644), .ZN(n20651) );
  OAI211_X1 U23579 ( .C1(NA), .C2(n20647), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n20653), .ZN(n20648) );
  OAI211_X1 U23580 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20750), .A(HOLD), .B(
        n20648), .ZN(n20649) );
  OAI22_X1 U23581 ( .A1(n20652), .A2(n20651), .B1(n20650), .B2(n20649), .ZN(
        P1_U3196) );
  OR2_X1 U23582 ( .A1(n20753), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20695) );
  OR2_X1 U23583 ( .A1(n20653), .A2(n20675), .ZN(n20691) );
  INV_X1 U23584 ( .A(n20691), .ZN(n20693) );
  AOI222_X1 U23585 ( .A1(n20689), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20753), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20693), .ZN(n20654) );
  INV_X1 U23586 ( .A(n20654), .ZN(P1_U3197) );
  AOI222_X1 U23587 ( .A1(n20693), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20675), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20689), .ZN(n20655) );
  INV_X1 U23588 ( .A(n20655), .ZN(P1_U3198) );
  OAI222_X1 U23589 ( .A1(n20691), .A2(n20657), .B1(n20656), .B2(n20752), .C1(
        n13774), .C2(n20695), .ZN(P1_U3199) );
  AOI222_X1 U23590 ( .A1(n20689), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20675), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20693), .ZN(n20658) );
  INV_X1 U23591 ( .A(n20658), .ZN(P1_U3200) );
  AOI222_X1 U23592 ( .A1(n20693), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20753), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20689), .ZN(n20659) );
  INV_X1 U23593 ( .A(n20659), .ZN(P1_U3201) );
  AOI222_X1 U23594 ( .A1(n20693), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20675), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20689), .ZN(n20660) );
  INV_X1 U23595 ( .A(n20660), .ZN(P1_U3202) );
  INV_X1 U23596 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20661) );
  INV_X1 U23597 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20892) );
  OAI222_X1 U23598 ( .A1(n20691), .A2(n20661), .B1(n20892), .B2(n20752), .C1(
        n14160), .C2(n20695), .ZN(P1_U3203) );
  AOI222_X1 U23599 ( .A1(n20689), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20675), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20693), .ZN(n20662) );
  INV_X1 U23600 ( .A(n20662), .ZN(P1_U3204) );
  AOI222_X1 U23601 ( .A1(n20693), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20675), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20689), .ZN(n20663) );
  INV_X1 U23602 ( .A(n20663), .ZN(P1_U3205) );
  AOI222_X1 U23603 ( .A1(n20689), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20675), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20693), .ZN(n20664) );
  INV_X1 U23604 ( .A(n20664), .ZN(P1_U3206) );
  AOI222_X1 U23605 ( .A1(n20693), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20675), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20689), .ZN(n20665) );
  INV_X1 U23606 ( .A(n20665), .ZN(P1_U3207) );
  AOI222_X1 U23607 ( .A1(n20693), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20675), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20689), .ZN(n20666) );
  INV_X1 U23608 ( .A(n20666), .ZN(P1_U3208) );
  AOI222_X1 U23609 ( .A1(n20693), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20675), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20689), .ZN(n20667) );
  INV_X1 U23610 ( .A(n20667), .ZN(P1_U3209) );
  AOI222_X1 U23611 ( .A1(n20689), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20675), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20693), .ZN(n20668) );
  INV_X1 U23612 ( .A(n20668), .ZN(P1_U3210) );
  AOI22_X1 U23613 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n20675), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20689), .ZN(n20669) );
  OAI21_X1 U23614 ( .B1(n20670), .B2(n20691), .A(n20669), .ZN(P1_U3211) );
  AOI22_X1 U23615 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20675), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20693), .ZN(n20671) );
  OAI21_X1 U23616 ( .B1(n20672), .B2(n20695), .A(n20671), .ZN(P1_U3212) );
  AOI222_X1 U23617 ( .A1(n20689), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20675), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20693), .ZN(n20673) );
  INV_X1 U23618 ( .A(n20673), .ZN(P1_U3213) );
  AOI222_X1 U23619 ( .A1(n20693), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20675), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20689), .ZN(n20674) );
  INV_X1 U23620 ( .A(n20674), .ZN(P1_U3214) );
  AOI222_X1 U23621 ( .A1(n20693), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20675), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n20689), .ZN(n20676) );
  INV_X1 U23622 ( .A(n20676), .ZN(P1_U3215) );
  AOI22_X1 U23623 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20675), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(n20689), .ZN(n20677) );
  OAI21_X1 U23624 ( .B1(n20678), .B2(n20691), .A(n20677), .ZN(P1_U3216) );
  AOI22_X1 U23625 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(n20675), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n20689), .ZN(n20679) );
  OAI21_X1 U23626 ( .B1(n14653), .B2(n20691), .A(n20679), .ZN(P1_U3217) );
  AOI22_X1 U23627 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20675), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n20693), .ZN(n20680) );
  OAI21_X1 U23628 ( .B1(n20682), .B2(n20695), .A(n20680), .ZN(P1_U3218) );
  AOI22_X1 U23629 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20675), .B1(
        P1_REIP_REG_24__SCAN_IN), .B2(n20689), .ZN(n20681) );
  OAI21_X1 U23630 ( .B1(n20682), .B2(n20691), .A(n20681), .ZN(P1_U3219) );
  AOI22_X1 U23631 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(n20675), .B1(
        P1_REIP_REG_24__SCAN_IN), .B2(n20693), .ZN(n20683) );
  OAI21_X1 U23632 ( .B1(n20684), .B2(n20695), .A(n20683), .ZN(P1_U3220) );
  AOI222_X1 U23633 ( .A1(n20693), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20753), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20689), .ZN(n20685) );
  INV_X1 U23634 ( .A(n20685), .ZN(P1_U3221) );
  AOI222_X1 U23635 ( .A1(n20689), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20753), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20693), .ZN(n20686) );
  INV_X1 U23636 ( .A(n20686), .ZN(P1_U3222) );
  AOI222_X1 U23637 ( .A1(n20693), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20753), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20689), .ZN(n20687) );
  INV_X1 U23638 ( .A(n20687), .ZN(P1_U3223) );
  AOI222_X1 U23639 ( .A1(n20693), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20753), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20689), .ZN(n20688) );
  INV_X1 U23640 ( .A(n20688), .ZN(P1_U3224) );
  AOI22_X1 U23641 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(n20675), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(n20689), .ZN(n20690) );
  OAI21_X1 U23642 ( .B1(n20692), .B2(n20691), .A(n20690), .ZN(P1_U3225) );
  AOI22_X1 U23643 ( .A1(P1_ADDRESS_REG_29__SCAN_IN), .A2(n20675), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(n20693), .ZN(n20694) );
  OAI21_X1 U23644 ( .B1(n20696), .B2(n20695), .A(n20694), .ZN(P1_U3226) );
  OAI22_X1 U23645 ( .A1(n20753), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20752), .ZN(n20697) );
  INV_X1 U23646 ( .A(n20697), .ZN(P1_U3458) );
  OAI22_X1 U23647 ( .A1(n20753), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20752), .ZN(n20698) );
  INV_X1 U23648 ( .A(n20698), .ZN(P1_U3459) );
  OAI22_X1 U23649 ( .A1(n20753), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20752), .ZN(n20699) );
  INV_X1 U23650 ( .A(n20699), .ZN(P1_U3460) );
  OAI22_X1 U23651 ( .A1(n20753), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20752), .ZN(n20700) );
  INV_X1 U23652 ( .A(n20700), .ZN(P1_U3461) );
  OAI21_X1 U23653 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20704), .A(n20702), 
        .ZN(n20701) );
  INV_X1 U23654 ( .A(n20701), .ZN(P1_U3464) );
  OAI21_X1 U23655 ( .B1(n20704), .B2(n20703), .A(n20702), .ZN(P1_U3465) );
  OAI21_X1 U23656 ( .B1(n9701), .B2(n20705), .A(n20707), .ZN(n20706) );
  OAI21_X1 U23657 ( .B1(n20708), .B2(n20707), .A(n20706), .ZN(n20709) );
  OAI21_X1 U23658 ( .B1(n20711), .B2(n20710), .A(n20709), .ZN(P1_U3469) );
  INV_X1 U23659 ( .A(n20725), .ZN(n20728) );
  INV_X1 U23660 ( .A(n20712), .ZN(n20713) );
  NAND2_X1 U23661 ( .A1(n20714), .A2(n20713), .ZN(n20723) );
  INV_X1 U23662 ( .A(n20715), .ZN(n20716) );
  NAND2_X1 U23663 ( .A1(n20717), .A2(n20716), .ZN(n20722) );
  OAI21_X1 U23664 ( .B1(n11999), .B2(n20742), .A(n20718), .ZN(n20720) );
  OR2_X1 U23665 ( .A1(n20720), .A2(n20719), .ZN(n20721) );
  AND4_X1 U23666 ( .A1(n20724), .A2(n20723), .A3(n20722), .A4(n20721), .ZN(
        n20726) );
  AOI22_X1 U23667 ( .A1(n20728), .A2(n20727), .B1(n20726), .B2(n20725), .ZN(
        P1_U3475) );
  AOI21_X1 U23668 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20730) );
  AOI22_X1 U23669 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20730), .B2(n20729), .ZN(n20733) );
  INV_X1 U23670 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20732) );
  AOI22_X1 U23671 ( .A1(n20736), .A2(n20733), .B1(n20732), .B2(n20731), .ZN(
        P1_U3481) );
  INV_X1 U23672 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20735) );
  OAI21_X1 U23673 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20736), .ZN(n20734) );
  OAI21_X1 U23674 ( .B1(n20736), .B2(n20735), .A(n20734), .ZN(P1_U3482) );
  AOI22_X1 U23675 ( .A1(n20752), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20737), 
        .B2(n20753), .ZN(P1_U3483) );
  OAI211_X1 U23676 ( .C1(n20741), .C2(n20740), .A(n20739), .B(n20738), .ZN(
        n20751) );
  AOI21_X1 U23677 ( .B1(n20743), .B2(n20742), .A(n12409), .ZN(n20745) );
  AOI21_X1 U23678 ( .B1(n20746), .B2(n20745), .A(n20744), .ZN(n20747) );
  OAI21_X1 U23679 ( .B1(n20748), .B2(n20747), .A(n20751), .ZN(n20749) );
  OAI21_X1 U23680 ( .B1(n20751), .B2(n20750), .A(n20749), .ZN(P1_U3485) );
  OAI22_X1 U23681 ( .A1(n20753), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n20752), .ZN(n20754) );
  INV_X1 U23682 ( .A(n20754), .ZN(P1_U3486) );
  AOI22_X1 U23683 ( .A1(n20758), .A2(n20757), .B1(n20756), .B2(n20755), .ZN(
        n20759) );
  INV_X1 U23684 ( .A(n20759), .ZN(n20765) );
  OAI22_X1 U23685 ( .A1(n20763), .A2(n20762), .B1(n20761), .B2(n20760), .ZN(
        n20764) );
  AOI211_X1 U23686 ( .C1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .C2(n20766), .A(
        n20765), .B(n20764), .ZN(n20930) );
  NOR3_X1 U23687 ( .A1(keyinput8), .A2(keyinput36), .A3(keyinput34), .ZN(
        n20793) );
  NAND2_X1 U23688 ( .A1(keyinput1), .A2(keyinput7), .ZN(n20771) );
  NAND2_X1 U23689 ( .A1(keyinput25), .A2(keyinput47), .ZN(n20767) );
  NOR3_X1 U23690 ( .A1(keyinput10), .A2(keyinput29), .A3(n20767), .ZN(n20769)
         );
  INV_X1 U23691 ( .A(keyinput46), .ZN(n20768) );
  NAND4_X1 U23692 ( .A1(keyinput49), .A2(keyinput15), .A3(n20769), .A4(n20768), 
        .ZN(n20770) );
  NOR4_X1 U23693 ( .A1(keyinput60), .A2(keyinput20), .A3(n20771), .A4(n20770), 
        .ZN(n20792) );
  NAND3_X1 U23694 ( .A1(keyinput3), .A2(keyinput18), .A3(keyinput33), .ZN(
        n20790) );
  NOR2_X1 U23695 ( .A1(keyinput21), .A2(keyinput50), .ZN(n20775) );
  NAND3_X1 U23696 ( .A1(keyinput54), .A2(keyinput53), .A3(keyinput62), .ZN(
        n20773) );
  NAND3_X1 U23697 ( .A1(keyinput28), .A2(keyinput41), .A3(keyinput23), .ZN(
        n20772) );
  NOR4_X1 U23698 ( .A1(keyinput24), .A2(keyinput31), .A3(n20773), .A4(n20772), 
        .ZN(n20774) );
  NAND4_X1 U23699 ( .A1(keyinput39), .A2(keyinput22), .A3(n20775), .A4(n20774), 
        .ZN(n20789) );
  NOR3_X1 U23700 ( .A1(keyinput16), .A2(keyinput57), .A3(keyinput59), .ZN(
        n20787) );
  NAND2_X1 U23701 ( .A1(keyinput14), .A2(keyinput17), .ZN(n20779) );
  NOR2_X1 U23702 ( .A1(keyinput12), .A2(keyinput11), .ZN(n20777) );
  NOR4_X1 U23703 ( .A1(keyinput35), .A2(keyinput61), .A3(keyinput45), .A4(
        keyinput42), .ZN(n20776) );
  NAND4_X1 U23704 ( .A1(keyinput56), .A2(keyinput52), .A3(n20777), .A4(n20776), 
        .ZN(n20778) );
  NOR4_X1 U23705 ( .A1(keyinput30), .A2(keyinput55), .A3(n20779), .A4(n20778), 
        .ZN(n20786) );
  NAND4_X1 U23706 ( .A1(keyinput5), .A2(keyinput9), .A3(keyinput48), .A4(
        keyinput40), .ZN(n20784) );
  NAND3_X1 U23707 ( .A1(keyinput58), .A2(keyinput0), .A3(keyinput27), .ZN(
        n20783) );
  NOR3_X1 U23708 ( .A1(keyinput51), .A2(keyinput32), .A3(keyinput37), .ZN(
        n20781) );
  NOR3_X1 U23709 ( .A1(keyinput26), .A2(keyinput4), .A3(keyinput6), .ZN(n20780) );
  NAND4_X1 U23710 ( .A1(keyinput44), .A2(n20781), .A3(keyinput2), .A4(n20780), 
        .ZN(n20782) );
  NOR4_X1 U23711 ( .A1(keyinput13), .A2(n20784), .A3(n20783), .A4(n20782), 
        .ZN(n20785) );
  NAND4_X1 U23712 ( .A1(keyinput38), .A2(n20787), .A3(n20786), .A4(n20785), 
        .ZN(n20788) );
  NOR4_X1 U23713 ( .A1(keyinput63), .A2(n20790), .A3(n20789), .A4(n20788), 
        .ZN(n20791) );
  NAND4_X1 U23714 ( .A1(keyinput19), .A2(n20793), .A3(n20792), .A4(n20791), 
        .ZN(n20794) );
  AOI21_X1 U23715 ( .B1(keyinput43), .B2(n20794), .A(n20795), .ZN(n20928) );
  INV_X1 U23716 ( .A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n20797) );
  AOI22_X1 U23717 ( .A1(keyinput49), .A2(n20797), .B1(keyinput43), .B2(n20795), 
        .ZN(n20796) );
  OAI21_X1 U23718 ( .B1(n20797), .B2(keyinput49), .A(n20796), .ZN(n20810) );
  AOI22_X1 U23719 ( .A1(n20800), .A2(keyinput7), .B1(keyinput60), .B2(n20799), 
        .ZN(n20798) );
  OAI221_X1 U23720 ( .B1(n20800), .B2(keyinput7), .C1(n20799), .C2(keyinput60), 
        .A(n20798), .ZN(n20809) );
  AOI22_X1 U23721 ( .A1(n20803), .A2(keyinput46), .B1(keyinput1), .B2(n20802), 
        .ZN(n20801) );
  OAI221_X1 U23722 ( .B1(n20803), .B2(keyinput46), .C1(n20802), .C2(keyinput1), 
        .A(n20801), .ZN(n20808) );
  INV_X1 U23723 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20804) );
  XOR2_X1 U23724 ( .A(keyinput20), .B(n20804), .Z(n20806) );
  XNOR2_X1 U23725 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B(keyinput8), .ZN(
        n20805) );
  NAND2_X1 U23726 ( .A1(n20806), .A2(n20805), .ZN(n20807) );
  NOR4_X1 U23727 ( .A1(n20810), .A2(n20809), .A3(n20808), .A4(n20807), .ZN(
        n20860) );
  INV_X1 U23728 ( .A(keyinput19), .ZN(n20812) );
  AOI22_X1 U23729 ( .A1(n20813), .A2(keyinput36), .B1(P3_DATAO_REG_3__SCAN_IN), 
        .B2(n20812), .ZN(n20811) );
  OAI221_X1 U23730 ( .B1(n20813), .B2(keyinput36), .C1(n20812), .C2(
        P3_DATAO_REG_3__SCAN_IN), .A(n20811), .ZN(n20824) );
  INV_X1 U23731 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n20815) );
  AOI22_X1 U23732 ( .A1(n20816), .A2(keyinput10), .B1(n20815), .B2(keyinput25), 
        .ZN(n20814) );
  OAI221_X1 U23733 ( .B1(n20816), .B2(keyinput10), .C1(n20815), .C2(keyinput25), .A(n20814), .ZN(n20823) );
  XOR2_X1 U23734 ( .A(n12986), .B(keyinput47), .Z(n20821) );
  XOR2_X1 U23735 ( .A(n20817), .B(keyinput29), .Z(n20820) );
  XNOR2_X1 U23736 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B(keyinput34), .ZN(
        n20819) );
  XNOR2_X1 U23737 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B(keyinput14), .ZN(
        n20818) );
  NAND4_X1 U23738 ( .A1(n20821), .A2(n20820), .A3(n20819), .A4(n20818), .ZN(
        n20822) );
  NOR3_X1 U23739 ( .A1(n20824), .A2(n20823), .A3(n20822), .ZN(n20859) );
  INV_X1 U23740 ( .A(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n20827) );
  AOI22_X1 U23741 ( .A1(n20827), .A2(keyinput11), .B1(keyinput16), .B2(n20826), 
        .ZN(n20825) );
  OAI221_X1 U23742 ( .B1(n20827), .B2(keyinput11), .C1(n20826), .C2(keyinput16), .A(n20825), .ZN(n20840) );
  AOI22_X1 U23743 ( .A1(n20830), .A2(keyinput17), .B1(keyinput30), .B2(n20829), 
        .ZN(n20828) );
  OAI221_X1 U23744 ( .B1(n20830), .B2(keyinput17), .C1(n20829), .C2(keyinput30), .A(n20828), .ZN(n20839) );
  INV_X1 U23745 ( .A(DATAI_30_), .ZN(n20833) );
  INV_X1 U23746 ( .A(keyinput12), .ZN(n20832) );
  AOI22_X1 U23747 ( .A1(n20833), .A2(keyinput52), .B1(
        P3_DATAWIDTH_REG_14__SCAN_IN), .B2(n20832), .ZN(n20831) );
  OAI221_X1 U23748 ( .B1(n20833), .B2(keyinput52), .C1(n20832), .C2(
        P3_DATAWIDTH_REG_14__SCAN_IN), .A(n20831), .ZN(n20838) );
  XOR2_X1 U23749 ( .A(n20834), .B(keyinput56), .Z(n20836) );
  XNOR2_X1 U23750 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B(keyinput55), .ZN(
        n20835) );
  NAND2_X1 U23751 ( .A1(n20836), .A2(n20835), .ZN(n20837) );
  NOR4_X1 U23752 ( .A1(n20840), .A2(n20839), .A3(n20838), .A4(n20837), .ZN(
        n20858) );
  INV_X1 U23753 ( .A(keyinput57), .ZN(n20842) );
  AOI22_X1 U23754 ( .A1(n20843), .A2(keyinput38), .B1(P2_M_IO_N_REG_SCAN_IN), 
        .B2(n20842), .ZN(n20841) );
  OAI221_X1 U23755 ( .B1(n20843), .B2(keyinput38), .C1(n20842), .C2(
        P2_M_IO_N_REG_SCAN_IN), .A(n20841), .ZN(n20856) );
  INV_X1 U23756 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n20846) );
  AOI22_X1 U23757 ( .A1(n20846), .A2(keyinput59), .B1(n20845), .B2(keyinput35), 
        .ZN(n20844) );
  OAI221_X1 U23758 ( .B1(n20846), .B2(keyinput59), .C1(n20845), .C2(keyinput35), .A(n20844), .ZN(n20855) );
  INV_X1 U23759 ( .A(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n20848) );
  AOI22_X1 U23760 ( .A1(n20849), .A2(keyinput61), .B1(keyinput45), .B2(n20848), 
        .ZN(n20847) );
  OAI221_X1 U23761 ( .B1(n20849), .B2(keyinput61), .C1(n20848), .C2(keyinput45), .A(n20847), .ZN(n20854) );
  AOI22_X1 U23762 ( .A1(n20852), .A2(keyinput42), .B1(keyinput39), .B2(n20851), 
        .ZN(n20850) );
  OAI221_X1 U23763 ( .B1(n20852), .B2(keyinput42), .C1(n20851), .C2(keyinput39), .A(n20850), .ZN(n20853) );
  NOR4_X1 U23764 ( .A1(n20856), .A2(n20855), .A3(n20854), .A4(n20853), .ZN(
        n20857) );
  NAND4_X1 U23765 ( .A1(n20860), .A2(n20859), .A3(n20858), .A4(n20857), .ZN(
        n20927) );
  AOI22_X1 U23766 ( .A1(n20863), .A2(keyinput62), .B1(n20862), .B2(keyinput28), 
        .ZN(n20861) );
  OAI221_X1 U23767 ( .B1(n20863), .B2(keyinput62), .C1(n20862), .C2(keyinput28), .A(n20861), .ZN(n20874) );
  INV_X1 U23768 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n20865) );
  AOI22_X1 U23769 ( .A1(n20866), .A2(keyinput53), .B1(keyinput24), .B2(n20865), 
        .ZN(n20864) );
  OAI221_X1 U23770 ( .B1(n20866), .B2(keyinput53), .C1(n20865), .C2(keyinput24), .A(n20864), .ZN(n20873) );
  AOI22_X1 U23771 ( .A1(n18166), .A2(keyinput31), .B1(n10478), .B2(keyinput51), 
        .ZN(n20867) );
  OAI221_X1 U23772 ( .B1(n18166), .B2(keyinput31), .C1(n10478), .C2(keyinput51), .A(n20867), .ZN(n20872) );
  INV_X1 U23773 ( .A(keyinput23), .ZN(n20869) );
  AOI22_X1 U23774 ( .A1(n20870), .A2(keyinput41), .B1(
        P2_DATAWIDTH_REG_24__SCAN_IN), .B2(n20869), .ZN(n20868) );
  OAI221_X1 U23775 ( .B1(n20870), .B2(keyinput41), .C1(n20869), .C2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A(n20868), .ZN(n20871) );
  NOR4_X1 U23776 ( .A1(n20874), .A2(n20873), .A3(n20872), .A4(n20871), .ZN(
        n20925) );
  AOI22_X1 U23777 ( .A1(n20877), .A2(keyinput50), .B1(keyinput3), .B2(n20876), 
        .ZN(n20875) );
  OAI221_X1 U23778 ( .B1(n20877), .B2(keyinput50), .C1(n20876), .C2(keyinput3), 
        .A(n20875), .ZN(n20890) );
  INV_X1 U23779 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n20880) );
  INV_X1 U23780 ( .A(P3_LWORD_REG_5__SCAN_IN), .ZN(n20879) );
  AOI22_X1 U23781 ( .A1(n20880), .A2(keyinput22), .B1(keyinput21), .B2(n20879), 
        .ZN(n20878) );
  OAI221_X1 U23782 ( .B1(n20880), .B2(keyinput22), .C1(n20879), .C2(keyinput21), .A(n20878), .ZN(n20889) );
  AOI22_X1 U23783 ( .A1(n20883), .A2(keyinput63), .B1(n20882), .B2(keyinput54), 
        .ZN(n20881) );
  OAI221_X1 U23784 ( .B1(n20883), .B2(keyinput63), .C1(n20882), .C2(keyinput54), .A(n20881), .ZN(n20888) );
  INV_X1 U23785 ( .A(DATAI_29_), .ZN(n20886) );
  INV_X1 U23786 ( .A(keyinput33), .ZN(n20885) );
  AOI22_X1 U23787 ( .A1(n20886), .A2(keyinput18), .B1(
        P3_ADDRESS_REG_29__SCAN_IN), .B2(n20885), .ZN(n20884) );
  OAI221_X1 U23788 ( .B1(n20886), .B2(keyinput18), .C1(n20885), .C2(
        P3_ADDRESS_REG_29__SCAN_IN), .A(n20884), .ZN(n20887) );
  NOR4_X1 U23789 ( .A1(n20890), .A2(n20889), .A3(n20888), .A4(n20887), .ZN(
        n20924) );
  INV_X1 U23790 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n20893) );
  AOI22_X1 U23791 ( .A1(n20893), .A2(keyinput6), .B1(keyinput58), .B2(n20892), 
        .ZN(n20891) );
  OAI221_X1 U23792 ( .B1(n20893), .B2(keyinput6), .C1(n20892), .C2(keyinput58), 
        .A(n20891), .ZN(n20906) );
  INV_X1 U23793 ( .A(P2_UWORD_REG_13__SCAN_IN), .ZN(n20896) );
  INV_X1 U23794 ( .A(keyinput2), .ZN(n20895) );
  AOI22_X1 U23795 ( .A1(n20896), .A2(keyinput4), .B1(
        P1_DATAWIDTH_REG_30__SCAN_IN), .B2(n20895), .ZN(n20894) );
  OAI221_X1 U23796 ( .B1(n20896), .B2(keyinput4), .C1(n20895), .C2(
        P1_DATAWIDTH_REG_30__SCAN_IN), .A(n20894), .ZN(n20905) );
  INV_X1 U23797 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n20899) );
  INV_X1 U23798 ( .A(keyinput15), .ZN(n20898) );
  AOI22_X1 U23799 ( .A1(n20899), .A2(keyinput13), .B1(
        P3_DATAWIDTH_REG_13__SCAN_IN), .B2(n20898), .ZN(n20897) );
  OAI221_X1 U23800 ( .B1(n20899), .B2(keyinput13), .C1(n20898), .C2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A(n20897), .ZN(n20904) );
  AOI22_X1 U23801 ( .A1(n20902), .A2(keyinput0), .B1(keyinput27), .B2(n20901), 
        .ZN(n20900) );
  OAI221_X1 U23802 ( .B1(n20902), .B2(keyinput0), .C1(n20901), .C2(keyinput27), 
        .A(n20900), .ZN(n20903) );
  NOR4_X1 U23803 ( .A1(n20906), .A2(n20905), .A3(n20904), .A4(n20903), .ZN(
        n20923) );
  INV_X1 U23804 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n20909) );
  INV_X1 U23805 ( .A(keyinput48), .ZN(n20908) );
  AOI22_X1 U23806 ( .A1(n20909), .A2(keyinput9), .B1(
        P3_ADDRESS_REG_26__SCAN_IN), .B2(n20908), .ZN(n20907) );
  OAI221_X1 U23807 ( .B1(n20909), .B2(keyinput9), .C1(n20908), .C2(
        P3_ADDRESS_REG_26__SCAN_IN), .A(n20907), .ZN(n20921) );
  AOI22_X1 U23808 ( .A1(n20912), .A2(keyinput37), .B1(keyinput5), .B2(n20911), 
        .ZN(n20910) );
  OAI221_X1 U23809 ( .B1(n20912), .B2(keyinput37), .C1(n20911), .C2(keyinput5), 
        .A(n20910), .ZN(n20920) );
  INV_X1 U23810 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n20914) );
  AOI22_X1 U23811 ( .A1(n20915), .A2(keyinput40), .B1(n20914), .B2(keyinput26), 
        .ZN(n20913) );
  OAI221_X1 U23812 ( .B1(n20915), .B2(keyinput40), .C1(n20914), .C2(keyinput26), .A(n20913), .ZN(n20919) );
  XNOR2_X1 U23813 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(keyinput32), 
        .ZN(n20917) );
  XNOR2_X1 U23814 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B(keyinput44), 
        .ZN(n20916) );
  NAND2_X1 U23815 ( .A1(n20917), .A2(n20916), .ZN(n20918) );
  NOR4_X1 U23816 ( .A1(n20921), .A2(n20920), .A3(n20919), .A4(n20918), .ZN(
        n20922) );
  NAND4_X1 U23817 ( .A1(n20925), .A2(n20924), .A3(n20923), .A4(n20922), .ZN(
        n20926) );
  NOR3_X1 U23818 ( .A1(n20928), .A2(n20927), .A3(n20926), .ZN(n20929) );
  XNOR2_X1 U23819 ( .A(n20930), .B(n20929), .ZN(P3_U2897) );
  AND2_X1 U11336 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14053) );
  NAND4_X2 U11090 ( .A1(n11378), .A2(n11377), .A3(n11376), .A4(n11375), .ZN(
        n11483) );
  NAND2_X1 U11102 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18808), .ZN(
        n12561) );
  INV_X2 U15638 ( .A(n14457), .ZN(n17132) );
  BUF_X2 U12350 ( .A(n12692), .Z(n17037) );
  INV_X1 U11032 ( .A(n16876), .ZN(n9919) );
  INV_X2 U11154 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18808) );
  CLKBUF_X2 U11035 ( .A(n12677), .Z(n17152) );
  BUF_X2 U11039 ( .A(n12716), .Z(n9588) );
  BUF_X2 U11052 ( .A(n12599), .Z(n15828) );
  CLKBUF_X1 U11053 ( .A(n12290), .Z(n12478) );
  NAND3_X1 U11058 ( .A1(n10552), .A2(n9760), .A3(n11081), .ZN(n10577) );
  CLKBUF_X1 U11094 ( .A(n11415), .Z(n12314) );
  CLKBUF_X1 U11097 ( .A(n11407), .Z(n12487) );
  CLKBUF_X2 U11103 ( .A(n12342), .Z(n12479) );
  AND2_X1 U11132 ( .A1(n13436), .A2(n11328), .ZN(n11554) );
  CLKBUF_X1 U11139 ( .A(n11422), .Z(n11968) );
  AND2_X1 U11145 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13435) );
  CLKBUF_X1 U11147 ( .A(n11584), .Z(n11632) );
  NAND2_X2 U11351 ( .A1(n10264), .A2(n19154), .ZN(n10972) );
  INV_X1 U11413 ( .A(n12703), .ZN(n12742) );
  CLKBUF_X1 U11438 ( .A(n11879), .Z(n11499) );
  CLKBUF_X1 U11497 ( .A(n11938), .Z(n11960) );
  NAND2_X1 U11527 ( .A1(n13638), .A2(n13435), .ZN(n13637) );
  CLKBUF_X2 U11528 ( .A(n11631), .Z(n13470) );
  CLKBUF_X1 U11569 ( .A(n20056), .Z(n20719) );
  NOR2_X1 U11644 ( .A1(n13845), .A2(n13913), .ZN(n14037) );
  NOR2_X1 U11704 ( .A1(n13187), .A2(n15439), .ZN(n12849) );
  CLKBUF_X1 U11755 ( .A(n11894), .Z(n11914) );
  CLKBUF_X1 U11770 ( .A(n17460), .Z(n17465) );
  CLKBUF_X1 U11922 ( .A(n16525), .Z(n16523) );
  AND2_X1 U12281 ( .A1(n17202), .A2(n18225), .ZN(n17339) );
  INV_X1 U12289 ( .A(n17339), .ZN(n20931) );
endmodule

