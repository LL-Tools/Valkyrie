

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1,
         READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n11143, n11145, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
         n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
         n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
         n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220,
         n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
         n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
         n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
         n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
         n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
         n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
         n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
         n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
         n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
         n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
         n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
         n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
         n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
         n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
         n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404,
         n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412,
         n17413, n17414, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
         n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
         n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
         n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
         n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
         n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
         n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
         n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
         n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
         n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
         n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
         n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
         n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
         n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158,
         n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
         n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
         n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
         n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
         n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
         n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
         n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
         n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
         n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
         n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
         n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
         n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
         n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
         n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
         n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
         n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
         n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294,
         n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
         n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
         n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
         n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
         n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
         n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
         n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350,
         n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
         n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
         n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
         n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
         n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
         n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
         n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422,
         n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
         n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
         n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470,
         n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
         n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
         n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494,
         n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
         n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
         n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
         n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542,
         n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
         n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
         n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
         n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
         n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582,
         n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
         n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
         n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
         n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982,
         n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990,
         n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
         n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
         n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
         n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022,
         n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
         n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
         n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
         n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
         n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102,
         n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
         n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
         n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126,
         n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134,
         n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
         n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150,
         n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158,
         n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
         n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174,
         n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182,
         n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
         n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198,
         n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206,
         n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214,
         n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222,
         n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230,
         n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238,
         n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246,
         n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254,
         n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262,
         n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270,
         n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278,
         n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286,
         n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294,
         n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302,
         n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310,
         n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318,
         n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326,
         n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334,
         n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342,
         n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350,
         n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358,
         n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366,
         n21367, n21368, n21369, n21370, n21371, n21373, n21374, n21375,
         n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383,
         n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391,
         n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399,
         n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407,
         n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415,
         n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423,
         n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431,
         n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439,
         n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447,
         n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455,
         n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463,
         n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471,
         n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479,
         n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487,
         n21488, n21489, n21490, n21491, n21492, n21493, n21494, n21495,
         n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503,
         n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511,
         n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519,
         n21520, n21521, n21522, n21523, n21524, n21525, n21526, n21527,
         n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535,
         n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543,
         n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551,
         n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559,
         n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567,
         n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575,
         n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583,
         n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591,
         n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21599,
         n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607,
         n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615,
         n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623,
         n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631,
         n21632, n21633, n21634, n21635, n21636, n21637, n21638, n21639,
         n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647,
         n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655,
         n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663,
         n21664, n21665, n21666, n21667, n21668, n21669, n21670, n21671,
         n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679,
         n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687,
         n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695,
         n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703,
         n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711,
         n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719,
         n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727,
         n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735,
         n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743,
         n21744, n21745, n21746, n21747, n21748, n21749, n21750, n21751,
         n21752, n21753, n21754, n21755, n21756, n21757, n21758, n21759,
         n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767,
         n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775,
         n21776, n21777, n21778, n21779, n21780, n21781, n21782, n21783,
         n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791,
         n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799,
         n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807,
         n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815,
         n21816, n21817, n21818, n21819, n21820, n21821, n21822, n21823,
         n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831,
         n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839,
         n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847,
         n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855,
         n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863,
         n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871,
         n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879,
         n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887,
         n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895,
         n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903,
         n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911,
         n21912, n21913, n21914, n21915, n21916, n21917, n21918, n21919,
         n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927,
         n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
         n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943,
         n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951,
         n21952, n21953, n21954, n21955, n21956, n21957, n21958, n21959,
         n21960, n21961, n21962, n21963, n21964, n21965, n21966, n21967,
         n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975,
         n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983,
         n21984, n21985, n21986, n21987, n21988, n21989, n21990, n21991,
         n21992, n21993, n21994, n21995, n21996, n21997, n21998, n21999,
         n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007,
         n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015,
         n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023,
         n22024, n22025, n22026, n22027, n22028, n22029, n22030, n22031,
         n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039,
         n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047,
         n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055,
         n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22063,
         n22064, n22065, n22066, n22067, n22068, n22069, n22070, n22071,
         n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079,
         n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087,
         n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095,
         n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103,
         n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111,
         n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119,
         n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127,
         n22128, n22129, n22130, n22131, n22132, n22133, n22134, n22135,
         n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143,
         n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151,
         n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159,
         n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167,
         n22168, n22169, n22170, n22171, n22172, n22173, n22174, n22175,
         n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183,
         n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191,
         n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199,
         n22200, n22201, n22202, n22203, n22204, n22205, n22206, n22207,
         n22208, n22209, n22210, n22211, n22212, n22213, n22214, n22215,
         n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223,
         n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231,
         n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239,
         n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247,
         n22248, n22249, n22250, n22251, n22252, n22253, n22254, n22255,
         n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263,
         n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271,
         n22272, n22273, n22274, n22275, n22276, n22277, n22278, n22279,
         n22280, n22281, n22282, n22283, n22284, n22285, n22286, n22287,
         n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295,
         n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303,
         n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311,
         n22312, n22313, n22314, n22315, n22316, n22317, n22318, n22319,
         n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327,
         n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335,
         n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343,
         n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351,
         n22352, n22353, n22354, n22355, n22356, n22357, n22358, n22359,
         n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367,
         n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375,
         n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383,
         n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391,
         n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399,
         n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407,
         n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415,
         n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423,
         n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431,
         n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439,
         n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447,
         n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455,
         n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463,
         n22464, n22465, n22466, n22467, n22468, n22469, n22470, n22471,
         n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479,
         n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487,
         n22488, n22489, n22490, n22491, n22492, n22493, n22494, n22495,
         n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503,
         n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511,
         n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519,
         n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527,
         n22528, n22529, n22530, n22531, n22532, n22533, n22534, n22535,
         n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543,
         n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551,
         n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559,
         n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567,
         n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575,
         n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583,
         n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591,
         n22592, n22593, n22594, n22595, n22596, n22597, n22598, n22599,
         n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607,
         n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615,
         n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623,
         n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631,
         n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639,
         n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647,
         n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655,
         n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663,
         n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671,
         n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679,
         n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687,
         n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695,
         n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703,
         n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711,
         n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719,
         n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727,
         n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735,
         n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743,
         n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751,
         n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759,
         n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767,
         n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775,
         n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783,
         n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791,
         n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799,
         n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807,
         n22808, n22809, n22810, n22811, n22812;

  AOI211_X1 U11250 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n16260), .A(
        n21963), .B(n14170), .ZN(n14174) );
  INV_X2 U11251 ( .A(n11541), .ZN(n17250) );
  INV_X2 U11252 ( .A(n21524), .ZN(n21443) );
  NOR2_X1 U11253 ( .A1(n13915), .A2(n13914), .ZN(n21336) );
  NAND2_X1 U11254 ( .A1(n13039), .A2(n13038), .ZN(n14748) );
  NAND2_X1 U11255 ( .A1(n11192), .A2(n16320), .ZN(n16304) );
  CLKBUF_X1 U11258 ( .A(n12062), .Z(n11987) );
  INV_X1 U11259 ( .A(n16454), .ZN(n16472) );
  CLKBUF_X1 U11260 ( .A(n13771), .Z(n18539) );
  NAND2_X1 U11261 ( .A1(n13949), .A2(n21396), .ZN(n13793) );
  CLKBUF_X1 U11262 ( .A(n13441), .Z(n13592) );
  CLKBUF_X2 U11263 ( .A(n12969), .Z(n13591) );
  INV_X2 U11264 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19436) );
  AND2_X1 U11265 ( .A1(n11864), .A2(n16489), .ZN(n16482) );
  INV_X1 U11266 ( .A(n11206), .ZN(n18545) );
  CLKBUF_X1 U11267 ( .A(n13801), .Z(n13899) );
  INV_X1 U11268 ( .A(n11359), .ZN(n16724) );
  CLKBUF_X2 U11269 ( .A(n13806), .Z(n11157) );
  CLKBUF_X2 U11270 ( .A(n13771), .Z(n18522) );
  CLKBUF_X1 U11272 ( .A(n13845), .Z(n18523) );
  AND2_X1 U11273 ( .A1(n11537), .A2(n12603), .ZN(n11662) );
  NAND2_X1 U11274 ( .A1(n11677), .A2(n12603), .ZN(n11699) );
  INV_X2 U11275 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21550) );
  CLKBUF_X2 U11276 ( .A(n11658), .Z(n19921) );
  AND2_X1 U11277 ( .A1(n12816), .A2(n14508), .ZN(n12969) );
  INV_X2 U11278 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11571) );
  CLKBUF_X1 U11279 ( .A(n20425), .Z(n11143) );
  NOR3_X1 U11280 ( .A1(n22310), .A2(n16030), .A3(n19985), .ZN(n20425) );
  INV_X1 U11282 ( .A(n22812), .ZN(n11145) );
  INV_X1 U11284 ( .A(n22812), .ZN(n11147) );
  INV_X1 U11285 ( .A(n22812), .ZN(n11148) );
  INV_X4 U11286 ( .A(n14030), .ZN(n11153) );
  BUF_X2 U11287 ( .A(n11853), .Z(n11182) );
  CLKBUF_X2 U11288 ( .A(n12847), .Z(n13583) );
  OAI211_X1 U11289 ( .C1(n13689), .C2(n12950), .A(n14315), .B(n13678), .ZN(
        n12954) );
  AND2_X1 U11290 ( .A1(n12815), .A2(n12816), .ZN(n12847) );
  NAND2_X1 U11292 ( .A1(n13023), .A2(n13022), .ZN(n13168) );
  AND2_X1 U11293 ( .A1(n11865), .A2(n16489), .ZN(n16424) );
  INV_X1 U11294 ( .A(n20330), .ZN(n12603) );
  INV_X2 U11295 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11830) );
  CLKBUF_X3 U11296 ( .A(n16322), .Z(n11150) );
  AND2_X1 U11297 ( .A1(n11491), .A2(n11229), .ZN(n16900) );
  INV_X1 U11298 ( .A(n14882), .ZN(n14314) );
  XNOR2_X1 U11299 ( .A(n13168), .B(n13167), .ZN(n14760) );
  AND2_X1 U11300 ( .A1(n11862), .A2(n11571), .ZN(n16217) );
  CLKBUF_X2 U11301 ( .A(n11719), .Z(n12738) );
  AND2_X1 U11302 ( .A1(n11847), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12024) );
  BUF_X1 U11304 ( .A(n13808), .Z(n18381) );
  INV_X1 U11305 ( .A(n21936), .ZN(n21746) );
  CLKBUF_X3 U11306 ( .A(n14760), .Z(n11195) );
  NAND2_X1 U11307 ( .A1(n11666), .A2(n11872), .ZN(n12641) );
  BUF_X1 U11308 ( .A(n16057), .Z(n19263) );
  NOR2_X1 U11309 ( .A1(n17388), .A2(n17390), .ZN(n17389) );
  INV_X2 U11310 ( .A(n12211), .ZN(n20174) );
  NOR2_X2 U11311 ( .A1(n18807), .A2(n21299), .ZN(n18806) );
  NAND2_X1 U11312 ( .A1(n21405), .A2(n21404), .ZN(n21345) );
  AND2_X2 U11313 ( .A1(n20970), .A2(n14115), .ZN(n18624) );
  INV_X1 U11314 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18862) );
  NAND2_X1 U11315 ( .A1(n18934), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20943) );
  NAND2_X1 U11318 ( .A1(n15191), .A2(n15192), .ZN(n15368) );
  BUF_X1 U11319 ( .A(n11652), .Z(n11163) );
  INV_X1 U11320 ( .A(n21162), .ZN(n21179) );
  NAND2_X1 U11321 ( .A1(n18624), .A2(n18577), .ZN(n18600) );
  AOI211_X1 U11322 ( .C1(n20761), .C2(n16930), .A(n16929), .B(n16928), .ZN(
        n16931) );
  INV_X2 U11323 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n21535) );
  AND2_X1 U11324 ( .A1(n12601), .A2(n20429), .ZN(n11149) );
  INV_X1 U11325 ( .A(n19263), .ZN(n19314) );
  AOI21_X2 U11326 ( .B1(n14427), .B2(n22287), .A(n11357), .ZN(n14761) );
  INV_X2 U11327 ( .A(n11661), .ZN(n11649) );
  NAND2_X2 U11328 ( .A1(n13185), .A2(n13177), .ZN(n14939) );
  OAI21_X2 U11329 ( .B1(n12792), .B2(n12795), .A(n11535), .ZN(n12578) );
  AND4_X2 U11330 ( .A1(n12851), .A2(n12850), .A3(n12849), .A4(n12848), .ZN(
        n12857) );
  NAND2_X4 U11331 ( .A1(n11149), .A2(n11685), .ZN(n11733) );
  XNOR2_X2 U11332 ( .A(n13019), .B(n13020), .ZN(n13146) );
  NOR2_X1 U11333 ( .A1(n14310), .A2(n16710), .ZN(n14183) );
  XNOR2_X2 U11334 ( .A(n12448), .B(n11316), .ZN(n17914) );
  XNOR2_X2 U11335 ( .A(n12658), .B(n12659), .ZN(n15469) );
  AOI21_X2 U11336 ( .B1(n17582), .B2(n17579), .A(n12754), .ZN(n17567) );
  OAI21_X2 U11337 ( .B1(n16344), .B2(n15178), .A(n14375), .ZN(n14606) );
  BUF_X1 U11338 ( .A(n17497), .Z(n17518) );
  NOR2_X1 U11339 ( .A1(n17593), .A2(n12765), .ZN(n17575) );
  AOI211_X1 U11340 ( .C1(n12803), .C2(n12802), .A(n12801), .B(n16408), .ZN(
        n12807) );
  NAND2_X1 U11341 ( .A1(n16081), .A2(n16083), .ZN(n16082) );
  NOR2_X1 U11342 ( .A1(n16356), .A2(n11484), .ZN(n11483) );
  AND2_X2 U11343 ( .A1(n17740), .A2(n11239), .ZN(n17337) );
  CLKBUF_X3 U11344 ( .A(n19314), .Z(n11181) );
  OR2_X1 U11345 ( .A1(n12328), .A2(n12325), .ZN(n12371) );
  INV_X1 U11346 ( .A(n11176), .ZN(n12357) );
  OR2_X1 U11347 ( .A1(n12328), .A2(n12324), .ZN(n12368) );
  AND2_X1 U11348 ( .A1(n16005), .A2(n11362), .ZN(n16275) );
  OR2_X1 U11349 ( .A1(n14592), .A2(n12327), .ZN(n12314) );
  OR2_X1 U11350 ( .A1(n14592), .A2(n12325), .ZN(n12301) );
  OR2_X1 U11351 ( .A1(n17320), .A2(n17319), .ZN(n17322) );
  AND2_X1 U11352 ( .A1(n11716), .A2(n11697), .ZN(n12290) );
  NOR2_X1 U11353 ( .A1(n15200), .A2(n15375), .ZN(n16073) );
  NAND2_X1 U11354 ( .A1(n13676), .A2(n13675), .ZN(n16719) );
  AND2_X1 U11355 ( .A1(n15112), .A2(n11681), .ZN(n12744) );
  OR2_X1 U11356 ( .A1(n12703), .A2(n12597), .ZN(n11709) );
  AND2_X1 U11357 ( .A1(n11686), .A2(n12709), .ZN(n15127) );
  AND2_X1 U11358 ( .A1(n11681), .A2(n11668), .ZN(n12710) );
  NAND2_X1 U11359 ( .A1(n18594), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18675) );
  INV_X2 U11360 ( .A(n16322), .ZN(n11192) );
  INV_X2 U11362 ( .A(n11659), .ZN(n12192) );
  AND2_X1 U11364 ( .A1(n11626), .A2(n11625), .ZN(n11666) );
  INV_X4 U11365 ( .A(n14319), .ZN(n16710) );
  AND4_X1 U11366 ( .A1(n12829), .A2(n12828), .A3(n12827), .A4(n12826), .ZN(
        n12836) );
  INV_X1 U11367 ( .A(n13843), .ZN(n18279) );
  NAND2_X1 U11368 ( .A1(n18902), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18886) );
  CLKBUF_X3 U11369 ( .A(n13799), .Z(n11159) );
  CLKBUF_X1 U11370 ( .A(n11847), .Z(n11158) );
  BUF_X2 U11372 ( .A(n12860), .Z(n13585) );
  CLKBUF_X2 U11373 ( .A(n13115), .Z(n12920) );
  BUF_X2 U11374 ( .A(n12983), .Z(n13595) );
  CLKBUF_X1 U11375 ( .A(n11847), .Z(n11184) );
  NAND2_X1 U11376 ( .A1(n12819), .A2(n14508), .ZN(n12897) );
  CLKBUF_X1 U11377 ( .A(n12876), .Z(n11152) );
  NOR2_X1 U11378 ( .A1(n13715), .A2(n21549), .ZN(n13771) );
  NOR2_X4 U11379 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12816) );
  NAND2_X1 U11380 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12257) );
  AND2_X1 U11381 ( .A1(n17485), .A2(n17484), .ZN(n17486) );
  AND3_X1 U11382 ( .A1(n12807), .A2(n12806), .A3(n12805), .ZN(n12808) );
  AND2_X1 U11383 ( .A1(n12748), .A2(n12747), .ZN(n12749) );
  AND2_X1 U11384 ( .A1(n12736), .A2(n11531), .ZN(n12748) );
  NAND3_X1 U11385 ( .A1(n16376), .A2(n16375), .A3(n16374), .ZN(n17108) );
  OR2_X1 U11386 ( .A1(n14060), .A2(n18103), .ZN(n14047) );
  OR2_X1 U11387 ( .A1(n16396), .A2(n19375), .ZN(n12736) );
  AND2_X1 U11388 ( .A1(n18094), .A2(n18093), .ZN(n19384) );
  NAND2_X1 U11389 ( .A1(n11326), .A2(n11324), .ZN(n12788) );
  NAND2_X1 U11390 ( .A1(n11305), .A2(n12755), .ZN(n11309) );
  AND2_X1 U11391 ( .A1(n17537), .A2(n11325), .ZN(n11324) );
  AND2_X1 U11392 ( .A1(n17492), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17493) );
  OR2_X1 U11393 ( .A1(n16900), .A2(n11541), .ZN(n16363) );
  NAND2_X1 U11394 ( .A1(n17575), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17556) );
  XNOR2_X1 U11395 ( .A(n16382), .B(n13613), .ZN(n16380) );
  NOR2_X1 U11396 ( .A1(n17622), .A2(n17853), .ZN(n17623) );
  NAND2_X1 U11397 ( .A1(n17541), .A2(n12541), .ZN(n17527) );
  OR2_X1 U11398 ( .A1(n12764), .A2(n11322), .ZN(n17593) );
  OR2_X1 U11399 ( .A1(n17883), .A2(n17865), .ZN(n17622) );
  AOI21_X1 U11400 ( .B1(n17601), .B2(n12751), .A(n12750), .ZN(n17592) );
  AND2_X2 U11401 ( .A1(n11462), .A2(n11218), .ZN(n17540) );
  NOR2_X1 U11402 ( .A1(n17389), .A2(n16576), .ZN(n16621) );
  OAI21_X1 U11403 ( .B1(n12674), .B2(n11316), .A(n12684), .ZN(n11315) );
  NAND2_X1 U11404 ( .A1(n12279), .A2(n16406), .ZN(n19354) );
  XNOR2_X1 U11405 ( .A(n12743), .B(n12742), .ZN(n19350) );
  NAND2_X1 U11406 ( .A1(n18754), .A2(n18755), .ZN(n18753) );
  OAI21_X1 U11407 ( .B1(n17638), .B2(n11427), .A(n18060), .ZN(n11426) );
  AND2_X1 U11408 ( .A1(n16575), .A2(n11533), .ZN(n16576) );
  AND2_X1 U11409 ( .A1(n12673), .A2(n12672), .ZN(n12674) );
  AND2_X1 U11410 ( .A1(n11444), .A2(n14031), .ZN(n18754) );
  XNOR2_X1 U11411 ( .A(n16643), .B(n12737), .ZN(n16686) );
  NAND3_X1 U11412 ( .A1(n16067), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n16068), .ZN(n16069) );
  NAND2_X2 U11413 ( .A1(n17915), .A2(n17914), .ZN(n17913) );
  OR2_X1 U11414 ( .A1(n19330), .A2(n19329), .ZN(n19332) );
  XNOR2_X1 U11415 ( .A(n16644), .B(n11391), .ZN(n19331) );
  NOR2_X1 U11416 ( .A1(n16644), .A2(n16645), .ZN(n16643) );
  CLKBUF_X1 U11417 ( .A(n14078), .Z(n19318) );
  NAND2_X1 U11418 ( .A1(n11355), .A2(n11354), .ZN(n11482) );
  NAND2_X1 U11419 ( .A1(n14082), .A2(n14041), .ZN(n16644) );
  XNOR2_X1 U11420 ( .A(n16326), .B(n16325), .ZN(n17106) );
  OR2_X1 U11421 ( .A1(n16738), .A2(n16737), .ZN(n17126) );
  NOR2_X1 U11422 ( .A1(n17010), .A2(n17013), .ZN(n17251) );
  OR2_X1 U11423 ( .A1(n15471), .A2(n15470), .ZN(n15473) );
  AND2_X1 U11424 ( .A1(n11447), .A2(n11446), .ZN(n18761) );
  OR2_X1 U11425 ( .A1(n17028), .A2(n16349), .ZN(n17009) );
  NAND2_X1 U11426 ( .A1(n12657), .A2(n12656), .ZN(n12659) );
  NAND2_X1 U11427 ( .A1(n11312), .A2(n12652), .ZN(n15393) );
  NOR2_X1 U11428 ( .A1(n18719), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18718) );
  NOR3_X1 U11429 ( .A1(n16195), .A2(n11398), .A3(n17424), .ZN(n17350) );
  NAND2_X1 U11430 ( .A1(n15296), .A2(n15295), .ZN(n15575) );
  AND2_X1 U11431 ( .A1(n17043), .A2(n17040), .ZN(n17029) );
  XNOR2_X1 U11432 ( .A(n15592), .B(n22012), .ZN(n20747) );
  INV_X4 U11433 ( .A(n11541), .ZN(n17256) );
  AND2_X2 U11434 ( .A1(n15584), .A2(n15604), .ZN(n11541) );
  AND2_X1 U11435 ( .A1(n12444), .A2(n12443), .ZN(n12680) );
  NOR2_X1 U11436 ( .A1(n21449), .A2(n21450), .ZN(n21475) );
  NAND2_X1 U11437 ( .A1(n13108), .A2(n13107), .ZN(n15584) );
  XNOR2_X1 U11438 ( .A(n13195), .B(n13194), .ZN(n15576) );
  AND2_X1 U11439 ( .A1(n16172), .A2(n11418), .ZN(n17743) );
  OR2_X1 U11440 ( .A1(n15194), .A2(n11394), .ZN(n15539) );
  NOR2_X1 U11441 ( .A1(n12544), .A2(n12543), .ZN(n12542) );
  AND4_X1 U11442 ( .A1(n12339), .A2(n12338), .A3(n12337), .A4(n12336), .ZN(
        n12350) );
  NAND2_X1 U11443 ( .A1(n13175), .A2(n13174), .ZN(n13185) );
  OAI22_X1 U11444 ( .A1(n12343), .A2(n12373), .B1(n12371), .B2(n12342), .ZN(
        n12344) );
  INV_X1 U11445 ( .A(n13176), .ZN(n13175) );
  AND2_X1 U11446 ( .A1(n12308), .A2(n12303), .ZN(n19975) );
  CLKBUF_X1 U11447 ( .A(n12359), .Z(n20070) );
  INV_X1 U11448 ( .A(n12368), .ZN(n19936) );
  INV_X1 U11449 ( .A(n12373), .ZN(n19923) );
  OR2_X1 U11450 ( .A1(n12326), .A2(n12313), .ZN(n12346) );
  OR2_X1 U11451 ( .A1(n12328), .A2(n12327), .ZN(n12373) );
  AOI21_X1 U11452 ( .B1(n14612), .B2(n14611), .A(n14607), .ZN(n14715) );
  NOR2_X1 U11453 ( .A1(n14722), .A2(n14723), .ZN(n14724) );
  XNOR2_X1 U11454 ( .A(n14612), .B(n14611), .ZN(n19944) );
  CLKBUF_X1 U11455 ( .A(n14759), .Z(n11196) );
  AND2_X1 U11456 ( .A1(n12312), .A2(n12316), .ZN(n12356) );
  NOR2_X1 U11457 ( .A1(n21653), .A2(n11147), .ZN(n21939) );
  BUF_X2 U11458 ( .A(n14705), .Z(n12303) );
  CLKBUF_X1 U11459 ( .A(n16151), .Z(n16894) );
  XNOR2_X1 U11460 ( .A(n13148), .B(n13147), .ZN(n14759) );
  NAND2_X1 U11461 ( .A1(n12288), .A2(n12292), .ZN(n19105) );
  XNOR2_X1 U11462 ( .A(n14606), .B(n14604), .ZN(n14612) );
  NOR2_X1 U11463 ( .A1(n21405), .A2(n21519), .ZN(n21492) );
  OAI21_X1 U11464 ( .B1(n22418), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n13052), 
        .ZN(n13166) );
  NOR3_X1 U11465 ( .A1(n20897), .A2(n21954), .A3(n20896), .ZN(n21119) );
  NAND2_X1 U11466 ( .A1(n12300), .A2(n12299), .ZN(n12325) );
  NAND2_X1 U11467 ( .A1(n13037), .A2(n13036), .ZN(n11373) );
  AND2_X1 U11468 ( .A1(n11728), .A2(n11729), .ZN(n12284) );
  NOR2_X2 U11469 ( .A1(n11221), .A2(n17953), .ZN(n21936) );
  AOI21_X1 U11470 ( .B1(n22807), .B2(n14187), .A(n22811), .ZN(n21967) );
  OR2_X2 U11471 ( .A1(n12273), .A2(n12272), .ZN(n12275) );
  NAND2_X1 U11472 ( .A1(n15460), .A2(n15459), .ZN(n15458) );
  NAND2_X1 U11473 ( .A1(n11311), .A2(n11310), .ZN(n12297) );
  NAND2_X1 U11474 ( .A1(n11321), .A2(n11320), .ZN(n11729) );
  OAI21_X2 U11475 ( .B1(n21340), .B2(n21339), .A(n21338), .ZN(n21529) );
  NAND2_X1 U11476 ( .A1(n18014), .A2(n22807), .ZN(n22277) );
  AND2_X1 U11477 ( .A1(n20718), .A2(n15356), .ZN(n15460) );
  NOR2_X2 U11478 ( .A1(n20328), .A2(n20426), .ZN(n20329) );
  NOR2_X2 U11479 ( .A1(n16241), .A2(n20426), .ZN(n16029) );
  NOR2_X2 U11480 ( .A1(n19919), .A2(n20426), .ZN(n19920) );
  OR2_X1 U11481 ( .A1(n11740), .A2(n11741), .ZN(n11743) );
  NOR2_X1 U11482 ( .A1(n20699), .A2(n15338), .ZN(n20718) );
  NOR2_X2 U11483 ( .A1(n20114), .A2(n20426), .ZN(n20115) );
  NOR2_X2 U11484 ( .A1(n20230), .A2(n20426), .ZN(n20231) );
  NOR2_X2 U11485 ( .A1(n20172), .A2(n20426), .ZN(n20173) );
  NAND2_X1 U11486 ( .A1(n11718), .A2(n11717), .ZN(n11727) );
  AND2_X1 U11487 ( .A1(n11424), .A2(n11422), .ZN(n15199) );
  OAI211_X1 U11488 ( .C1(n11715), .C2(n19436), .A(n11714), .B(n11713), .ZN(
        n12293) );
  INV_X1 U11489 ( .A(n22416), .ZN(n11154) );
  NAND2_X1 U11490 ( .A1(n13035), .A2(n13034), .ZN(n13038) );
  NAND2_X1 U11491 ( .A1(n12955), .A2(n13013), .ZN(n13155) );
  NOR2_X1 U11492 ( .A1(n14686), .A2(n11367), .ZN(n11366) );
  AND2_X1 U11493 ( .A1(n13929), .A2(n11256), .ZN(n14145) );
  AND2_X1 U11494 ( .A1(n12715), .A2(n11708), .ZN(n11715) );
  AND2_X1 U11495 ( .A1(n12707), .A2(n11648), .ZN(n11708) );
  INV_X1 U11496 ( .A(n14685), .ZN(n14684) );
  OAI21_X1 U11497 ( .B1(n12962), .B2(n12946), .A(n14319), .ZN(n12938) );
  AND2_X1 U11498 ( .A1(n14683), .A2(n14682), .ZN(n14685) );
  NAND2_X1 U11499 ( .A1(n12245), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12266) );
  OAI21_X1 U11500 ( .B1(n16304), .B2(P1_EBX_REG_1__SCAN_IN), .A(n14648), .ZN(
        n14679) );
  NAND2_X1 U11501 ( .A1(n11471), .A2(n11647), .ZN(n11707) );
  NAND2_X1 U11502 ( .A1(n18648), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n18672) );
  INV_X1 U11503 ( .A(n16304), .ZN(n16293) );
  AND2_X2 U11504 ( .A1(n15127), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11720) );
  NOR2_X2 U11505 ( .A1(n18675), .A2(n20902), .ZN(n18648) );
  AND2_X1 U11506 ( .A1(n12940), .A2(n12939), .ZN(n16711) );
  NAND2_X1 U11507 ( .A1(n11192), .A2(n16385), .ZN(n16297) );
  INV_X1 U11508 ( .A(n12023), .ZN(n12086) );
  NAND2_X1 U11509 ( .A1(n14857), .A2(n16385), .ZN(n16323) );
  AND2_X1 U11510 ( .A1(n12882), .A2(n12881), .ZN(n12883) );
  AND2_X2 U11511 ( .A1(n12018), .A2(n12017), .ZN(n12685) );
  BUF_X2 U11512 ( .A(n12192), .Z(n12211) );
  AND3_X1 U11513 ( .A1(n16136), .A2(n20233), .A3(n12192), .ZN(n11663) );
  CLKBUF_X1 U11514 ( .A(n13617), .Z(n15602) );
  NAND2_X1 U11515 ( .A1(n13760), .A2(n13759), .ZN(n13949) );
  CLKBUF_X2 U11516 ( .A(n11601), .Z(n20233) );
  INV_X2 U11517 ( .A(n11666), .ZN(n19080) );
  NAND3_X1 U11518 ( .A1(n13854), .A2(n13853), .A3(n13852), .ZN(n20904) );
  NAND2_X1 U11519 ( .A1(n11579), .A2(n11578), .ZN(n11658) );
  OR2_X2 U11520 ( .A1(n20825), .A2(n20771), .ZN(n20811) );
  OR2_X1 U11521 ( .A1(n11243), .A2(n13811), .ZN(n21525) );
  NAND2_X1 U11523 ( .A1(n11599), .A2(n11598), .ZN(n16031) );
  NAND2_X1 U11524 ( .A1(n11566), .A2(n11565), .ZN(n11601) );
  OR2_X1 U11525 ( .A1(n13009), .A2(n13008), .ZN(n14636) );
  NAND2_X2 U11526 ( .A1(n12836), .A2(n12835), .ZN(n14882) );
  NAND2_X1 U11527 ( .A1(n11468), .A2(n11466), .ZN(n11661) );
  AND4_X1 U11528 ( .A1(n11618), .A2(n11617), .A3(n11616), .A4(n11615), .ZN(
        n11619) );
  AND4_X1 U11529 ( .A1(n12901), .A2(n12900), .A3(n12899), .A4(n12898), .ZN(
        n12907) );
  AND4_X1 U11530 ( .A1(n12919), .A2(n12918), .A3(n12917), .A4(n12916), .ZN(
        n12931) );
  AND4_X1 U11531 ( .A1(n12915), .A2(n12914), .A3(n12913), .A4(n12912), .ZN(
        n12932) );
  AND4_X1 U11532 ( .A1(n12880), .A2(n12879), .A3(n12878), .A4(n12877), .ZN(
        n11209) );
  AND4_X1 U11533 ( .A1(n12845), .A2(n12844), .A3(n12843), .A4(n12842), .ZN(
        n11540) );
  INV_X2 U11534 ( .A(U214), .ZN(n20825) );
  AND4_X1 U11535 ( .A1(n11623), .A2(n11622), .A3(n11621), .A4(n11620), .ZN(
        n11624) );
  AND4_X1 U11536 ( .A1(n12864), .A2(n12863), .A3(n12862), .A4(n12861), .ZN(
        n12869) );
  AND4_X1 U11537 ( .A1(n12834), .A2(n12833), .A3(n12832), .A4(n12831), .ZN(
        n12835) );
  CLKBUF_X1 U11538 ( .A(n19059), .Z(n22359) );
  AND4_X1 U11539 ( .A1(n12855), .A2(n12854), .A3(n12853), .A4(n12852), .ZN(
        n12856) );
  INV_X1 U11540 ( .A(n13746), .ZN(n13843) );
  AND4_X1 U11541 ( .A1(n12924), .A2(n12923), .A3(n12922), .A4(n12921), .ZN(
        n12930) );
  AND2_X2 U11542 ( .A1(n16676), .A2(n11571), .ZN(n16481) );
  AND4_X1 U11543 ( .A1(n12928), .A2(n12927), .A3(n12926), .A4(n12925), .ZN(
        n12929) );
  INV_X2 U11544 ( .A(n19811), .ZN(U215) );
  INV_X1 U11545 ( .A(n13710), .ZN(n18254) );
  BUF_X2 U11546 ( .A(n13845), .Z(n18497) );
  BUF_X2 U11547 ( .A(n13808), .Z(n18540) );
  INV_X2 U11548 ( .A(n22343), .ZN(n22352) );
  CLKBUF_X2 U11549 ( .A(n13807), .Z(n18548) );
  INV_X2 U11550 ( .A(n12897), .ZN(n12896) );
  BUF_X2 U11551 ( .A(n12830), .Z(n13561) );
  BUF_X2 U11552 ( .A(n12989), .Z(n13566) );
  OR2_X2 U11553 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18571), .ZN(n14030) );
  OR2_X1 U11554 ( .A1(n14159), .A2(n14172), .ZN(n18414) );
  AND2_X2 U11555 ( .A1(n11863), .A2(n11830), .ZN(n11853) );
  AND2_X2 U11556 ( .A1(n12818), .A2(n14746), .ZN(n11178) );
  INV_X2 U11557 ( .A(n20550), .ZN(n20600) );
  AND2_X2 U11558 ( .A1(n12818), .A2(n14746), .ZN(n13593) );
  BUF_X2 U11559 ( .A(n12984), .Z(n13594) );
  AND2_X2 U11560 ( .A1(n11477), .A2(n14508), .ZN(n12983) );
  BUF_X2 U11561 ( .A(n12990), .Z(n13596) );
  INV_X2 U11562 ( .A(n19068), .ZN(n22321) );
  NOR2_X1 U11563 ( .A1(n12257), .A2(n15402), .ZN(n12254) );
  AND2_X2 U11564 ( .A1(n11543), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11849) );
  AND2_X2 U11565 ( .A1(n11361), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12818) );
  AND2_X2 U11566 ( .A1(n11865), .A2(n11830), .ZN(n11639) );
  AND2_X2 U11567 ( .A1(n12809), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11477) );
  INV_X1 U11568 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21541) );
  INV_X1 U11569 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15402) );
  CLKBUF_X1 U11570 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n19360) );
  INV_X1 U11571 ( .A(n12945), .ZN(n11160) );
  NAND2_X2 U11572 ( .A1(n12846), .A2(n11540), .ZN(n13614) );
  AND2_X4 U11573 ( .A1(n11863), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11847) );
  NOR2_X1 U11574 ( .A1(n11664), .A2(n11161), .ZN(n11682) );
  NAND2_X1 U11575 ( .A1(n20429), .A2(n12188), .ZN(n11161) );
  AND2_X2 U11576 ( .A1(n11663), .A2(n11662), .ZN(n12601) );
  INV_X1 U11577 ( .A(n12933), .ZN(n11162) );
  NOR2_X1 U11578 ( .A1(n21167), .A2(n21168), .ZN(n21181) );
  NAND2_X1 U11579 ( .A1(n15575), .A2(n15574), .ZN(n20742) );
  AND2_X4 U11580 ( .A1(n12810), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12815) );
  INV_X2 U11581 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12810) );
  NOR2_X2 U11582 ( .A1(n21193), .A2(n21192), .ZN(n21208) );
  CLKBUF_X1 U11583 ( .A(n12744), .Z(n11164) );
  NAND2_X1 U11585 ( .A1(n11356), .A2(n11482), .ZN(n17004) );
  NAND2_X1 U11586 ( .A1(n11163), .A2(n16031), .ZN(n11166) );
  INV_X1 U11587 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11167) );
  NAND2_X1 U11588 ( .A1(n11661), .A2(n11659), .ZN(n11652) );
  INV_X2 U11589 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12809) );
  NAND2_X1 U11590 ( .A1(n20752), .A2(n15601), .ZN(n11168) );
  NAND2_X2 U11591 ( .A1(n20754), .A2(n20753), .ZN(n20752) );
  NOR2_X4 U11592 ( .A1(n21134), .A2(n18579), .ZN(n18594) );
  XNOR2_X2 U11593 ( .A(n18773), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n20908) );
  NAND2_X2 U11594 ( .A1(n11667), .A2(n11709), .ZN(n11698) );
  NOR2_X2 U11595 ( .A1(n21469), .A2(n21463), .ZN(n21462) );
  NOR4_X2 U11596 ( .A1(n21368), .A2(n21343), .A3(n21342), .A4(n21341), .ZN(
        n21403) );
  NOR2_X2 U11597 ( .A1(n13874), .A2(n13873), .ZN(n21524) );
  NAND2_X1 U11598 ( .A1(n12253), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11169) );
  OR2_X2 U11599 ( .A1(n11169), .A2(n11170), .ZN(n12250) );
  OR2_X1 U11600 ( .A1(n11171), .A2(n18077), .ZN(n11170) );
  INV_X1 U11601 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11171) );
  NAND2_X1 U11602 ( .A1(n12249), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11172) );
  OR2_X2 U11603 ( .A1(n11172), .A2(n11173), .ZN(n12244) );
  OR2_X1 U11604 ( .A1(n11174), .A2(n12246), .ZN(n11173) );
  INV_X1 U11605 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11174) );
  NOR2_X1 U11606 ( .A1(n12257), .A2(n15402), .ZN(n11175) );
  NOR2_X2 U11607 ( .A1(n17401), .A2(n17400), .ZN(n17402) );
  NOR2_X2 U11608 ( .A1(n17414), .A2(n17416), .ZN(n17410) );
  OR2_X1 U11609 ( .A1(n14705), .A2(n12301), .ZN(n11176) );
  NOR2_X1 U11610 ( .A1(n12326), .A2(n12325), .ZN(n20036) );
  NOR2_X4 U11611 ( .A1(n12244), .A2(n12231), .ZN(n12245) );
  INV_X2 U11612 ( .A(n12421), .ZN(n12317) );
  INV_X1 U11613 ( .A(n11149), .ZN(n12216) );
  NAND2_X1 U11614 ( .A1(n11847), .A2(n11571), .ZN(n16454) );
  NOR2_X4 U11615 ( .A1(n12250), .A2(n19177), .ZN(n12251) );
  NOR2_X2 U11616 ( .A1(n19289), .A2(n19288), .ZN(n19287) );
  NOR2_X2 U11617 ( .A1(n14099), .A2(n11181), .ZN(n19289) );
  NAND2_X2 U11618 ( .A1(n12251), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12262) );
  NOR2_X4 U11619 ( .A1(n12262), .A2(n17616), .ZN(n12249) );
  NAND2_X1 U11620 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n12249), .ZN(
        n12263) );
  NOR2_X1 U11621 ( .A1(n12263), .A2(n12246), .ZN(n12265) );
  INV_X2 U11622 ( .A(n14705), .ZN(n12312) );
  OR2_X1 U11623 ( .A1(n13687), .A2(n12948), .ZN(n14315) );
  NAND2_X1 U11624 ( .A1(n14314), .A2(n13614), .ZN(n14310) );
  AND2_X4 U11625 ( .A1(n12818), .A2(n12816), .ZN(n12968) );
  NOR2_X1 U11626 ( .A1(n12260), .A2(n18077), .ZN(n12252) );
  NAND2_X2 U11627 ( .A1(n12815), .A2(n14746), .ZN(n12875) );
  OAI21_X2 U11628 ( .B1(n17871), .B2(n12467), .A(n12466), .ZN(n17629) );
  NAND2_X2 U11629 ( .A1(n17913), .A2(n11201), .ZN(n17871) );
  AND2_X1 U11630 ( .A1(n12954), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13025) );
  AND2_X1 U11631 ( .A1(n12818), .A2(n14746), .ZN(n11177) );
  NAND2_X2 U11632 ( .A1(n11703), .A2(n11684), .ZN(n11719) );
  OAI21_X2 U11633 ( .B1(n11683), .B2(n11682), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n11684) );
  NOR2_X2 U11634 ( .A1(n14090), .A2(n19314), .ZN(n17359) );
  NOR2_X2 U11635 ( .A1(n14091), .A2(n19277), .ZN(n14090) );
  AND2_X1 U11636 ( .A1(n12815), .A2(n12816), .ZN(n11179) );
  NOR2_X4 U11637 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12817) );
  AND2_X1 U11640 ( .A1(n13082), .A2(n13175), .ZN(n13193) );
  NOR2_X2 U11641 ( .A1(n14815), .A2(n14816), .ZN(n14814) );
  OAI21_X1 U11642 ( .B1(n14939), .B2(n13289), .A(n13183), .ZN(n14868) );
  BUF_X1 U11643 ( .A(n14760), .Z(n11194) );
  AND2_X1 U11644 ( .A1(n16361), .A2(n11541), .ZN(n16362) );
  OAI21_X2 U11645 ( .B1(n17527), .B2(n17528), .A(n17529), .ZN(n17519) );
  NAND2_X2 U11646 ( .A1(n12982), .A2(n12981), .ZN(n13019) );
  XNOR2_X1 U11647 ( .A(n13185), .B(n13184), .ZN(n15288) );
  BUF_X8 U11648 ( .A(n11853), .Z(n11183) );
  NOR2_X2 U11649 ( .A1(n12266), .A2(n17558), .ZN(n12243) );
  XNOR2_X2 U11650 ( .A(n11349), .B(n11348), .ZN(n22416) );
  INV_X1 U11651 ( .A(n12947), .ZN(n11185) );
  INV_X4 U11652 ( .A(n12875), .ZN(n13453) );
  AND2_X1 U11653 ( .A1(n11849), .A2(n11830), .ZN(n11186) );
  AND2_X2 U11654 ( .A1(n11849), .A2(n11830), .ZN(n11187) );
  AND2_X1 U11655 ( .A1(n11849), .A2(n11830), .ZN(n11855) );
  AND2_X4 U11656 ( .A1(n11477), .A2(n12817), .ZN(n12860) );
  INV_X1 U11657 ( .A(n12897), .ZN(n11189) );
  INV_X1 U11658 ( .A(n12896), .ZN(n11190) );
  AND2_X1 U11659 ( .A1(n12819), .A2(n12815), .ZN(n11191) );
  NOR2_X2 U11660 ( .A1(n13211), .A2(n15311), .ZN(n15325) );
  OAI21_X2 U11661 ( .B1(n14939), .B2(n14938), .A(n14937), .ZN(n15285) );
  OAI21_X2 U11662 ( .B1(n12954), .B2(n12951), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n13029) );
  NOR2_X2 U11663 ( .A1(n16976), .A2(n17080), .ZN(n16358) );
  AOI22_X4 U11664 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12732), .B1(n16399), 
        .B2(n19436), .ZN(n16057) );
  XNOR2_X2 U11665 ( .A(n12234), .B(n12233), .ZN(n16399) );
  NOR2_X4 U11666 ( .A1(n16744), .A2(n16745), .ZN(n16263) );
  XNOR2_X2 U11667 ( .A(n14748), .B(n14823), .ZN(n14427) );
  AND2_X1 U11668 ( .A1(n14287), .A2(n16710), .ZN(n12935) );
  NAND2_X1 U11669 ( .A1(n13040), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13624) );
  NOR2_X1 U11670 ( .A1(n13715), .A2(n13716), .ZN(n13807) );
  INV_X1 U11671 ( .A(n13582), .ZN(n13557) );
  INV_X1 U11672 ( .A(n13204), .ZN(n13108) );
  INV_X1 U11673 ( .A(n13624), .ZN(n13674) );
  NAND2_X1 U11674 ( .A1(n12484), .A2(n12538), .ZN(n12544) );
  INV_X1 U11675 ( .A(n11726), .ZN(n11320) );
  INV_X1 U11676 ( .A(n11727), .ZN(n11321) );
  NOR2_X1 U11677 ( .A1(n11712), .A2(n11711), .ZN(n11713) );
  OAI22_X1 U11678 ( .A1(n11698), .A2(n11701), .B1(n19360), .B2(n11720), .ZN(
        n11705) );
  XNOR2_X1 U11679 ( .A(n12574), .B(n12213), .ZN(n12572) );
  NAND2_X1 U11680 ( .A1(n17629), .A2(n12482), .ZN(n11463) );
  NOR2_X1 U11681 ( .A1(n14644), .A2(n11415), .ZN(n11414) );
  INV_X1 U11682 ( .A(n14622), .ZN(n11415) );
  NAND2_X1 U11683 ( .A1(n11644), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11645) );
  NAND2_X1 U11684 ( .A1(n11638), .A2(n11571), .ZN(n11646) );
  NOR2_X1 U11685 ( .A1(n13719), .A2(n21549), .ZN(n13801) );
  NOR2_X1 U11686 ( .A1(n13715), .A2(n13718), .ZN(n13799) );
  NAND2_X1 U11687 ( .A1(n21559), .A2(n21550), .ZN(n13715) );
  NAND2_X1 U11688 ( .A1(n13791), .A2(n21376), .ZN(n13825) );
  NAND2_X1 U11689 ( .A1(n13553), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15064) );
  NAND2_X1 U11690 ( .A1(n16651), .A2(n12186), .ZN(n12701) );
  AND2_X1 U11691 ( .A1(n16649), .A2(n16648), .ZN(n16651) );
  OR2_X1 U11692 ( .A1(n20319), .A2(n14581), .ZN(n16141) );
  XNOR2_X1 U11693 ( .A(n12687), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18060) );
  NAND2_X1 U11694 ( .A1(n11456), .A2(n11454), .ZN(n12792) );
  INV_X1 U11695 ( .A(n11455), .ZN(n11454) );
  NAND2_X1 U11696 ( .A1(n12564), .A2(n11457), .ZN(n11456) );
  OAI21_X1 U11697 ( .B1(n12566), .B2(n11458), .A(n16696), .ZN(n11455) );
  NAND2_X1 U11698 ( .A1(n17567), .A2(n11306), .ZN(n11305) );
  NOR2_X1 U11699 ( .A1(n12756), .A2(n11307), .ZN(n11306) );
  INV_X1 U11700 ( .A(n17568), .ZN(n11307) );
  INV_X1 U11701 ( .A(n14145), .ZN(n14153) );
  NAND2_X1 U11702 ( .A1(n19331), .A2(n18091), .ZN(n11393) );
  AND2_X1 U11703 ( .A1(n11840), .A2(n11839), .ZN(n11842) );
  NOR2_X1 U11704 ( .A1(n14761), .A2(n13081), .ZN(n13082) );
  OR2_X1 U11705 ( .A1(n12979), .A2(n12978), .ZN(n14635) );
  OR2_X1 U11706 ( .A1(n12940), .A2(n14319), .ZN(n12936) );
  AOI22_X1 U11707 ( .A1(n12989), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12990), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11372) );
  NAND4_X1 U11708 ( .A1(n11955), .A2(n11521), .A3(n11954), .A4(n11953), .ZN(
        n12354) );
  NAND2_X1 U11709 ( .A1(n11328), .A2(n11327), .ZN(n12626) );
  NAND2_X1 U11710 ( .A1(n12194), .A2(n12641), .ZN(n11327) );
  NAND2_X1 U11711 ( .A1(n12351), .A2(n12581), .ZN(n11328) );
  AOI21_X1 U11712 ( .B1(n16217), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n11331), .ZN(n11330) );
  INV_X1 U11713 ( .A(n11930), .ZN(n11331) );
  INV_X1 U11714 ( .A(n12764), .ZN(n11430) );
  OAI22_X1 U11715 ( .A1(n12341), .A2(n12367), .B1(n12368), .B2(n12340), .ZN(
        n12345) );
  OR2_X1 U11716 ( .A1(n11895), .A2(n11894), .ZN(n12647) );
  AOI21_X1 U11717 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19952), .A(
        n11842), .ZN(n11843) );
  AOI22_X1 U11718 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11182), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11593) );
  NAND2_X1 U11719 ( .A1(n11559), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11560) );
  NAND2_X1 U11720 ( .A1(n11856), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11559) );
  NOR2_X1 U11721 ( .A1(n21391), .A2(n13793), .ZN(n13792) );
  AOI21_X1 U11722 ( .B1(n19524), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13987), .ZN(n13994) );
  AND2_X1 U11723 ( .A1(n13974), .A2(n11300), .ZN(n11299) );
  NAND2_X1 U11724 ( .A1(n11380), .A2(n11378), .ZN(n16744) );
  NOR2_X1 U11725 ( .A1(n11381), .A2(n11379), .ZN(n11378) );
  INV_X1 U11726 ( .A(n16790), .ZN(n11380) );
  INV_X1 U11727 ( .A(n16758), .ZN(n11379) );
  NAND2_X1 U11728 ( .A1(n16768), .A2(n11382), .ZN(n11381) );
  INV_X1 U11729 ( .A(n11383), .ZN(n11382) );
  NOR2_X1 U11730 ( .A1(n16801), .A2(n11377), .ZN(n11376) );
  INV_X1 U11731 ( .A(n16835), .ZN(n11377) );
  NAND2_X1 U11732 ( .A1(n14481), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13607) );
  NOR2_X1 U11733 ( .A1(n13286), .A2(n13285), .ZN(n13302) );
  NAND2_X1 U11734 ( .A1(n11237), .A2(n11204), .ZN(n11388) );
  NOR2_X1 U11735 ( .A1(n11490), .A2(n17097), .ZN(n11489) );
  INV_X1 U11736 ( .A(n16919), .ZN(n11490) );
  AND2_X1 U11737 ( .A1(n11483), .A2(n17256), .ZN(n11479) );
  INV_X1 U11738 ( .A(n16356), .ZN(n11354) );
  NAND2_X1 U11739 ( .A1(n17252), .A2(n16352), .ZN(n11355) );
  NOR2_X1 U11740 ( .A1(n11363), .A2(n16160), .ZN(n11362) );
  INV_X1 U11741 ( .A(n11364), .ZN(n11363) );
  NAND2_X1 U11742 ( .A1(n11352), .A2(n15591), .ZN(n15592) );
  NAND2_X1 U11743 ( .A1(n11353), .A2(n15584), .ZN(n11352) );
  OR2_X1 U11744 ( .A1(n13068), .A2(n13067), .ZN(n15289) );
  INV_X1 U11745 ( .A(n13025), .ZN(n11349) );
  OAI21_X1 U11746 ( .B1(n13029), .B2(n12810), .A(n12953), .ZN(n11348) );
  INV_X1 U11747 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18000) );
  INV_X1 U11748 ( .A(n12412), .ZN(n11336) );
  NOR2_X1 U11749 ( .A1(n12408), .A2(n12407), .ZN(n12413) );
  NOR2_X1 U11750 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16489) );
  INV_X1 U11751 ( .A(n17456), .ZN(n11408) );
  NAND2_X1 U11752 ( .A1(n11502), .A2(n17407), .ZN(n11501) );
  INV_X1 U11753 ( .A(n17411), .ZN(n11500) );
  NAND2_X1 U11754 ( .A1(n16129), .A2(n11236), .ZN(n17414) );
  AND2_X1 U11755 ( .A1(n12163), .A2(n12162), .ZN(n16238) );
  INV_X1 U11756 ( .A(n17767), .ZN(n11420) );
  AND2_X1 U11757 ( .A1(n14596), .A2(n19079), .ZN(n16597) );
  NAND2_X1 U11758 ( .A1(n11495), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11494) );
  NAND2_X1 U11759 ( .A1(n11493), .A2(n11571), .ZN(n11492) );
  INV_X1 U11760 ( .A(n16045), .ZN(n11402) );
  NOR2_X1 U11761 ( .A1(n11459), .A2(n11458), .ZN(n11457) );
  NAND2_X1 U11762 ( .A1(n11345), .A2(n11344), .ZN(n14035) );
  NOR2_X1 U11763 ( .A1(n17500), .A2(n17507), .ZN(n11344) );
  INV_X1 U11764 ( .A(n17499), .ZN(n11345) );
  NOR2_X1 U11765 ( .A1(n14080), .A2(n12685), .ZN(n14036) );
  OR2_X1 U11766 ( .A1(n19238), .A2(n12685), .ZN(n12525) );
  NOR2_X1 U11767 ( .A1(n14996), .A2(n11412), .ZN(n11411) );
  INV_X1 U11768 ( .A(n14819), .ZN(n11412) );
  OR2_X1 U11769 ( .A1(n12686), .A2(n12685), .ZN(n12687) );
  NAND2_X1 U11770 ( .A1(n15393), .A2(n12654), .ZN(n12658) );
  NAND2_X1 U11771 ( .A1(n11407), .A2(n11729), .ZN(n12287) );
  OR2_X1 U11772 ( .A1(n14380), .A2(n11898), .ZN(n11917) );
  OR2_X1 U11773 ( .A1(n19105), .A2(n12300), .ZN(n12313) );
  NAND2_X1 U11774 ( .A1(n11572), .A2(n11571), .ZN(n11579) );
  NOR2_X1 U11775 ( .A1(n11259), .A2(n11285), .ZN(n11284) );
  INV_X1 U11776 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11285) );
  OAI211_X1 U11777 ( .C1(n13755), .C2(n13754), .A(n13753), .B(n11517), .ZN(
        n13756) );
  NAND2_X1 U11778 ( .A1(n18480), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11246) );
  NOR2_X1 U11779 ( .A1(n13716), .A2(n13719), .ZN(n13806) );
  INV_X1 U11780 ( .A(n11437), .ZN(n11433) );
  OAI21_X1 U11781 ( .B1(n11441), .B2(n13819), .A(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11437) );
  INV_X1 U11782 ( .A(n11452), .ZN(n13836) );
  OAI21_X1 U11783 ( .B1(n18847), .B2(n11453), .A(n18845), .ZN(n11452) );
  NOR2_X1 U11784 ( .A1(n18755), .A2(n18877), .ZN(n14122) );
  OAI21_X1 U11785 ( .B1(n18892), .B2(n18891), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13961) );
  NAND2_X1 U11786 ( .A1(n18903), .A2(n13824), .ZN(n13826) );
  NOR2_X1 U11787 ( .A1(n13795), .A2(n13794), .ZN(n13797) );
  INV_X1 U11788 ( .A(n13793), .ZN(n13795) );
  NAND2_X1 U11789 ( .A1(n21345), .A2(n11301), .ZN(n13974) );
  NAND2_X1 U11790 ( .A1(n19727), .A2(n21336), .ZN(n11301) );
  AOI21_X1 U11791 ( .B1(n18393), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n11270), .ZN(n13862) );
  NOR2_X1 U11792 ( .A1(n18254), .A2(n11271), .ZN(n11270) );
  AOI21_X1 U11793 ( .B1(n18547), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n11260), .ZN(n13892) );
  NOR2_X1 U11794 ( .A1(n18254), .A2(n11261), .ZN(n11260) );
  NAND2_X1 U11795 ( .A1(n11297), .A2(n11296), .ZN(n13937) );
  AND2_X1 U11796 ( .A1(n22424), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13611) );
  NOR2_X2 U11797 ( .A1(n16729), .A2(n16383), .ZN(n16382) );
  AND2_X1 U11798 ( .A1(n13552), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13553) );
  OR2_X1 U11799 ( .A1(n16914), .A2(n13557), .ZN(n13581) );
  NAND2_X1 U11800 ( .A1(n13473), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13512) );
  NAND2_X1 U11801 ( .A1(n13326), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13340) );
  NAND2_X1 U11802 ( .A1(n16933), .A2(n17132), .ZN(n16899) );
  NAND2_X1 U11803 ( .A1(n15348), .A2(n15347), .ZN(n17320) );
  INV_X1 U11804 ( .A(n15349), .ZN(n15347) );
  INV_X1 U11805 ( .A(n15458), .ZN(n15348) );
  INV_X1 U11806 ( .A(n14686), .ZN(n11369) );
  NAND2_X1 U11807 ( .A1(n14684), .A2(n14860), .ZN(n11367) );
  NAND2_X1 U11808 ( .A1(n13058), .A2(n13057), .ZN(n14823) );
  NOR2_X1 U11809 ( .A1(n15033), .A2(n11195), .ZN(n22401) );
  INV_X1 U11810 ( .A(n11193), .ZN(n22471) );
  NAND2_X1 U11811 ( .A1(n22287), .A2(n14787), .ZN(n22678) );
  NAND2_X1 U11812 ( .A1(n13674), .A2(n13673), .ZN(n13675) );
  NAND2_X1 U11813 ( .A1(n13672), .A2(n13671), .ZN(n13676) );
  INV_X2 U11814 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n22424) );
  NAND2_X1 U11815 ( .A1(n12542), .A2(n11235), .ZN(n12550) );
  INV_X1 U11816 ( .A(n12547), .ZN(n11343) );
  OR2_X1 U11817 ( .A1(n15316), .A2(n15317), .ZN(n16171) );
  AND2_X1 U11818 ( .A1(n12157), .A2(n12156), .ZN(n16170) );
  NAND2_X1 U11819 ( .A1(n11508), .A2(n15370), .ZN(n11507) );
  OR2_X1 U11820 ( .A1(n11395), .A2(n15448), .ZN(n11394) );
  NAND2_X1 U11821 ( .A1(n11421), .A2(n11240), .ZN(n14085) );
  NAND2_X1 U11822 ( .A1(n16172), .A2(n11232), .ZN(n17770) );
  AND2_X1 U11823 ( .A1(n14381), .A2(n14382), .ZN(n14380) );
  INV_X1 U11824 ( .A(n11426), .ZN(n11425) );
  OAI21_X1 U11825 ( .B1(n12675), .B2(n11316), .A(n12678), .ZN(n11314) );
  OR2_X1 U11826 ( .A1(n16651), .A2(n12186), .ZN(n12187) );
  AND2_X1 U11827 ( .A1(n11414), .A2(n14667), .ZN(n11413) );
  NAND2_X1 U11828 ( .A1(n12678), .A2(n17911), .ZN(n17639) );
  NAND2_X1 U11829 ( .A1(n14471), .A2(n14470), .ZN(n14469) );
  INV_X1 U11830 ( .A(n11915), .ZN(n11424) );
  AOI21_X1 U11831 ( .B1(n14469), .B2(n11917), .A(n11916), .ZN(n11915) );
  NOR2_X1 U11832 ( .A1(n11872), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n14377) );
  NAND2_X1 U11833 ( .A1(n14718), .A2(n14717), .ZN(n14732) );
  NOR2_X1 U11834 ( .A1(n19944), .A2(n19929), .ZN(n20015) );
  OR2_X1 U11835 ( .A1(n19435), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16022) );
  NOR2_X1 U11836 ( .A1(n20058), .A2(n16017), .ZN(n19941) );
  NOR2_X1 U11837 ( .A1(n13766), .A2(n11449), .ZN(n11448) );
  AND2_X1 U11838 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11449) );
  INV_X1 U11839 ( .A(n11514), .ZN(n18538) );
  NOR2_X1 U11840 ( .A1(n18969), .A2(n18957), .ZN(n18682) );
  NAND2_X1 U11841 ( .A1(n18904), .A2(n18905), .ZN(n18903) );
  NAND2_X1 U11842 ( .A1(n18761), .A2(n18738), .ZN(n11445) );
  NAND2_X1 U11843 ( .A1(n18743), .A2(n14137), .ZN(n14017) );
  NAND2_X1 U11844 ( .A1(n14130), .A2(n13934), .ZN(n11257) );
  NOR2_X1 U11845 ( .A1(n11221), .A2(n20841), .ZN(n11255) );
  NOR2_X1 U11846 ( .A1(n13819), .A2(n11442), .ZN(n11441) );
  INV_X1 U11847 ( .A(n11435), .ZN(n11443) );
  NAND2_X1 U11848 ( .A1(n18938), .A2(n13815), .ZN(n18929) );
  INV_X1 U11849 ( .A(n21614), .ZN(n14137) );
  AND2_X1 U11850 ( .A1(n13983), .A2(n11219), .ZN(n11256) );
  OAI22_X1 U11851 ( .A1(n14114), .A2(n21847), .B1(n14136), .B2(n21614), .ZN(
        n14132) );
  NOR2_X1 U11852 ( .A1(n20904), .A2(n13937), .ZN(n20841) );
  AND2_X1 U11853 ( .A1(n16378), .A2(n15069), .ZN(n22266) );
  NAND2_X1 U11854 ( .A1(n13691), .A2(n14212), .ZN(n16054) );
  INV_X1 U11855 ( .A(n20728), .ZN(n20760) );
  INV_X1 U11856 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n22457) );
  NAND2_X1 U11857 ( .A1(n14761), .A2(n11195), .ZN(n14874) );
  OR2_X1 U11858 ( .A1(n14874), .A2(n15415), .ZN(n22742) );
  XNOR2_X1 U11859 ( .A(n12701), .B(n12700), .ZN(n19347) );
  INV_X1 U11860 ( .A(n20327), .ZN(n19914) );
  INV_X1 U11861 ( .A(n18127), .ZN(n16017) );
  AND2_X1 U11862 ( .A1(n14372), .A2(n14371), .ZN(n20319) );
  AND2_X1 U11863 ( .A1(n18076), .A2(n17961), .ZN(n18091) );
  INV_X1 U11864 ( .A(n12300), .ZN(n16344) );
  INV_X1 U11865 ( .A(n18091), .ZN(n18105) );
  INV_X1 U11866 ( .A(n18106), .ZN(n18079) );
  XNOR2_X1 U11867 ( .A(n12576), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12577) );
  INV_X1 U11868 ( .A(n16645), .ZN(n11391) );
  AOI21_X1 U11869 ( .B1(n11459), .B2(n12566), .A(n11458), .ZN(n11460) );
  NAND2_X1 U11870 ( .A1(n17556), .A2(n12780), .ZN(n11326) );
  NAND2_X1 U11871 ( .A1(n17550), .A2(n12780), .ZN(n11325) );
  OAI21_X1 U11872 ( .B1(n17548), .B2(n17550), .A(n11308), .ZN(n12761) );
  INV_X1 U11873 ( .A(n19375), .ZN(n19420) );
  OR2_X1 U11874 ( .A1(n12746), .A2(n12704), .ZN(n17928) );
  INV_X1 U11875 ( .A(n19929), .ZN(n20081) );
  INV_X1 U11876 ( .A(n20100), .ZN(n20096) );
  NAND2_X1 U11877 ( .A1(n14132), .A2(n21956), .ZN(n21964) );
  INV_X1 U11878 ( .A(n18793), .ZN(n18794) );
  OR2_X1 U11879 ( .A1(n18798), .A2(n11251), .ZN(n11250) );
  AND2_X1 U11880 ( .A1(n18808), .A2(n21314), .ZN(n11251) );
  INV_X1 U11881 ( .A(n18870), .ZN(n18881) );
  INV_X1 U11882 ( .A(n18974), .ZN(n18962) );
  NAND2_X1 U11883 ( .A1(n11720), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n11688) );
  AND4_X1 U11884 ( .A1(n12363), .A2(n12362), .A3(n12361), .A4(n12360), .ZN(
        n12380) );
  AOI21_X1 U11885 ( .B1(n12358), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n12188), .ZN(n12319) );
  INV_X1 U11886 ( .A(n12709), .ZN(n11471) );
  OR2_X1 U11887 ( .A1(n13993), .A2(n13994), .ZN(n13988) );
  NAND2_X1 U11888 ( .A1(n13193), .A2(n13194), .ZN(n13204) );
  AND2_X1 U11889 ( .A1(n13106), .A2(n13105), .ZN(n13203) );
  OR2_X1 U11890 ( .A1(n13092), .A2(n13091), .ZN(n15587) );
  NOR2_X1 U11891 ( .A1(n12499), .A2(n12485), .ZN(n12484) );
  NAND2_X1 U11892 ( .A1(n11698), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11718) );
  OR2_X1 U11893 ( .A1(n12582), .A2(n12395), .ZN(n11836) );
  AOI22_X1 U11894 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11583) );
  NAND2_X1 U11895 ( .A1(n12562), .A2(n12561), .ZN(n12570) );
  NAND2_X1 U11896 ( .A1(n12681), .A2(n12680), .ZN(n12686) );
  INV_X1 U11897 ( .A(n12679), .ZN(n12681) );
  BUF_X1 U11898 ( .A(n12385), .Z(n12657) );
  AOI22_X1 U11899 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n12365), .B1(
        n12366), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12347) );
  NOR2_X1 U11900 ( .A1(n12311), .A2(n12310), .ZN(n12332) );
  AOI22_X1 U11901 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12356), .B1(
        n19975), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U11902 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19942), .B1(
        n19936), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12330) );
  NOR2_X1 U11903 ( .A1(n12194), .A2(n11844), .ZN(n12592) );
  AOI21_X1 U11904 ( .B1(n11856), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11545) );
  AOI21_X1 U11905 ( .B1(n18540), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n11262), .ZN(n18406) );
  NOR2_X1 U11906 ( .A1(n11259), .A2(n11263), .ZN(n11262) );
  INV_X1 U11907 ( .A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11263) );
  AOI21_X1 U11908 ( .B1(n18393), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n11272), .ZN(n18397) );
  NOR2_X1 U11909 ( .A1(n11259), .A2(n11273), .ZN(n11272) );
  INV_X1 U11910 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11273) );
  AOI21_X1 U11911 ( .B1(n20948), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n11288), .ZN(n18370) );
  NOR2_X1 U11912 ( .A1(n11259), .A2(n11289), .ZN(n11288) );
  INV_X1 U11913 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11289) );
  NAND2_X1 U11914 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n21535), .ZN(
        n13716) );
  NAND2_X1 U11915 ( .A1(n21550), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13719) );
  NAND2_X1 U11916 ( .A1(n21541), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13718) );
  NAND2_X1 U11917 ( .A1(n11529), .A2(n11384), .ZN(n11383) );
  INV_X1 U11918 ( .A(n16791), .ZN(n11384) );
  INV_X1 U11919 ( .A(n13607), .ZN(n13573) );
  NOR2_X1 U11920 ( .A1(n17279), .A2(n11365), .ZN(n11364) );
  INV_X1 U11921 ( .A(n15555), .ZN(n11365) );
  OR2_X1 U11922 ( .A1(n17250), .A2(n16353), .ZN(n17040) );
  AND2_X1 U11923 ( .A1(n12933), .A2(n12941), .ZN(n12942) );
  NAND2_X1 U11924 ( .A1(n14289), .A2(n14314), .ZN(n12961) );
  OR2_X1 U11925 ( .A1(n12996), .A2(n12995), .ZN(n15606) );
  NAND2_X1 U11926 ( .A1(n12980), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12981) );
  OR2_X1 U11927 ( .A1(n14310), .A2(n16321), .ZN(n14428) );
  OR2_X1 U11928 ( .A1(n14458), .A2(n14457), .ZN(n17994) );
  AOI22_X1 U11929 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12830), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12834) );
  NOR2_X1 U11930 ( .A1(n12894), .A2(n12893), .ZN(n11360) );
  INV_X1 U11931 ( .A(n14757), .ZN(n14787) );
  OR2_X1 U11932 ( .A1(n13670), .A2(n13683), .ZN(n13671) );
  AND2_X2 U11933 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14746) );
  NAND2_X1 U11934 ( .A1(n19080), .A2(n12188), .ZN(n12589) );
  NAND2_X1 U11935 ( .A1(n12242), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12239) );
  INV_X1 U11936 ( .A(n12484), .ZN(n12539) );
  OR2_X1 U11937 ( .A1(n12490), .A2(n12491), .ZN(n12489) );
  NOR2_X1 U11938 ( .A1(n12511), .A2(n12504), .ZN(n12500) );
  NOR2_X1 U11939 ( .A1(n12517), .A2(n12516), .ZN(n11347) );
  OR2_X1 U11940 ( .A1(n12513), .A2(n12512), .ZN(n12517) );
  NOR2_X1 U11941 ( .A1(n11342), .A2(n11341), .ZN(n11340) );
  INV_X1 U11942 ( .A(n12456), .ZN(n11341) );
  INV_X1 U11943 ( .A(n12458), .ZN(n11342) );
  NOR2_X1 U11944 ( .A1(n12455), .A2(n12453), .ZN(n12459) );
  AND2_X1 U11945 ( .A1(n12459), .A2(n12458), .ZN(n12461) );
  NAND2_X1 U11946 ( .A1(n11319), .A2(n11716), .ZN(n11318) );
  INV_X1 U11947 ( .A(n16234), .ZN(n11512) );
  AND2_X1 U11948 ( .A1(n16131), .A2(n16211), .ZN(n11513) );
  AND2_X1 U11949 ( .A1(n11411), .A2(n15188), .ZN(n11410) );
  NOR2_X1 U11950 ( .A1(n11933), .A2(n11329), .ZN(n12351) );
  NAND2_X1 U11951 ( .A1(n12243), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12241) );
  OR2_X1 U11952 ( .A1(n11396), .A2(n15490), .ZN(n11395) );
  NAND2_X1 U11953 ( .A1(n11397), .A2(n15366), .ZN(n11396) );
  INV_X1 U11954 ( .A(n15195), .ZN(n11397) );
  OR2_X1 U11955 ( .A1(n11911), .A2(n11910), .ZN(n12645) );
  OR2_X1 U11956 ( .A1(n12570), .A2(n12569), .ZN(n12574) );
  INV_X1 U11957 ( .A(n12408), .ZN(n11335) );
  NOR2_X1 U11958 ( .A1(n11333), .A2(n12391), .ZN(n11332) );
  AND2_X1 U11959 ( .A1(n11406), .A2(n17335), .ZN(n11405) );
  INV_X1 U11960 ( .A(n17387), .ZN(n11406) );
  AND2_X1 U11961 ( .A1(n11429), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11428) );
  AND2_X1 U11962 ( .A1(n12693), .A2(n17707), .ZN(n11429) );
  AND2_X1 U11963 ( .A1(n11232), .A2(n11419), .ZN(n11418) );
  INV_X1 U11964 ( .A(n16238), .ZN(n11419) );
  NAND2_X1 U11965 ( .A1(n17611), .A2(n17612), .ZN(n17601) );
  AOI21_X1 U11966 ( .B1(n12482), .B2(n17628), .A(n11465), .ZN(n11464) );
  INV_X1 U11967 ( .A(n18087), .ZN(n11465) );
  AOI21_X1 U11968 ( .B1(n19180), .B2(n12019), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17628) );
  NOR2_X1 U11969 ( .A1(n12671), .A2(n12667), .ZN(n12664) );
  OAI21_X1 U11970 ( .B1(n11475), .B2(n12680), .A(n12665), .ZN(n12666) );
  NAND2_X1 U11971 ( .A1(n12662), .A2(n12661), .ZN(n12663) );
  AND3_X1 U11972 ( .A1(n11958), .A2(n11957), .A3(n11956), .ZN(n15375) );
  OR2_X1 U11973 ( .A1(n11871), .A2(n11870), .ZN(n12396) );
  INV_X1 U11974 ( .A(n12294), .ZN(n11311) );
  INV_X1 U11975 ( .A(n12293), .ZN(n11310) );
  AND2_X2 U11976 ( .A1(n11547), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11863) );
  INV_X1 U11977 ( .A(n11854), .ZN(n15126) );
  AND2_X1 U11978 ( .A1(n16597), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14597) );
  OR2_X1 U11979 ( .A1(n14600), .A2(n16516), .ZN(n14604) );
  AOI221_X1 U11980 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n11843), 
        .C1(n19364), .C2(n11843), .A(n11835), .ZN(n12631) );
  AND2_X1 U11981 ( .A1(n19436), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14704) );
  NAND2_X1 U11982 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n14155), .ZN(
        n14151) );
  AOI21_X1 U11983 ( .B1(n11156), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n11280), .ZN(n18413) );
  NOR2_X1 U11984 ( .A1(n11259), .A2(n11281), .ZN(n11280) );
  INV_X1 U11985 ( .A(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11281) );
  AOI21_X1 U11986 ( .B1(n11156), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n11278), .ZN(n18343) );
  NOR2_X1 U11987 ( .A1(n11259), .A2(n11279), .ZN(n11278) );
  INV_X1 U11988 ( .A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11279) );
  AOI21_X1 U11989 ( .B1(n20948), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n11290), .ZN(n18349) );
  NOR2_X1 U11990 ( .A1(n11259), .A2(n11291), .ZN(n11290) );
  INV_X1 U11991 ( .A(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11291) );
  AOI22_X1 U11992 ( .A1(n18480), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18546), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18268) );
  AOI21_X1 U11993 ( .B1(n11159), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n11264), .ZN(n18298) );
  NOR2_X1 U11994 ( .A1(n11259), .A2(n11265), .ZN(n11264) );
  INV_X1 U11995 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11265) );
  OR2_X1 U11996 ( .A1(n13716), .A2(n14172), .ZN(n11206) );
  NAND2_X1 U11997 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21559), .ZN(
        n13717) );
  NOR2_X1 U11998 ( .A1(n13717), .A2(n13718), .ZN(n13808) );
  AND2_X1 U11999 ( .A1(n18712), .A2(n18702), .ZN(n11522) );
  NOR2_X1 U12000 ( .A1(n21740), .A2(n21827), .ZN(n18737) );
  NAND2_X1 U12001 ( .A1(n21443), .A2(n13935), .ZN(n13976) );
  INV_X1 U12002 ( .A(n13961), .ZN(n13959) );
  NAND2_X1 U12003 ( .A1(n18942), .A2(n13951), .ZN(n13952) );
  NAND2_X1 U12004 ( .A1(n18952), .A2(n13813), .ZN(n13814) );
  NOR2_X1 U12005 ( .A1(n11253), .A2(n20841), .ZN(n14133) );
  INV_X1 U12006 ( .A(n11257), .ZN(n11253) );
  NAND2_X1 U12007 ( .A1(n21541), .A2(n21535), .ZN(n14159) );
  NAND2_X1 U12008 ( .A1(n11302), .A2(n11298), .ZN(n13933) );
  NAND2_X1 U12009 ( .A1(n13927), .A2(n11303), .ZN(n11302) );
  NAND2_X1 U12010 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14172) );
  AOI22_X1 U12011 ( .A1(n18480), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18546), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13913) );
  AOI21_X1 U12012 ( .B1(n18279), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n11286), .ZN(n13895) );
  NOR2_X1 U12013 ( .A1(n18254), .A2(n11287), .ZN(n11286) );
  AOI21_X1 U12014 ( .B1(n11156), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n11266), .ZN(n13879) );
  NOR2_X1 U12015 ( .A1(n18254), .A2(n11267), .ZN(n11266) );
  INV_X1 U12016 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15361) );
  NAND2_X1 U12017 ( .A1(n15067), .A2(n22066), .ZN(n22091) );
  NAND2_X1 U12018 ( .A1(n15079), .A2(n15078), .ZN(n22262) );
  AND2_X1 U12019 ( .A1(n16159), .A2(n16158), .ZN(n16160) );
  AOI21_X1 U12020 ( .B1(n14587), .B2(n14586), .A(n22331), .ZN(n20604) );
  INV_X1 U12021 ( .A(n14212), .ZN(n14357) );
  OR3_X1 U12022 ( .A1(n16719), .A2(n13689), .A3(n22302), .ZN(n14191) );
  NOR2_X1 U12023 ( .A1(n16731), .A2(n11390), .ZN(n11389) );
  INV_X1 U12024 ( .A(n16264), .ZN(n11390) );
  AND2_X1 U12025 ( .A1(n13513), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13514) );
  NOR2_X1 U12026 ( .A1(n13472), .A2(n16962), .ZN(n13473) );
  AND2_X1 U12027 ( .A1(n13495), .A2(n13494), .ZN(n16768) );
  OR2_X1 U12028 ( .A1(n13424), .A2(n16978), .ZN(n13425) );
  OR2_X1 U12029 ( .A1(n13425), .A2(n13448), .ZN(n13472) );
  AND2_X1 U12030 ( .A1(n11375), .A2(n11223), .ZN(n11374) );
  INV_X1 U12031 ( .A(n16872), .ZN(n11375) );
  AND2_X1 U12032 ( .A1(n13356), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13357) );
  NAND2_X1 U12033 ( .A1(n13357), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13389) );
  NOR2_X1 U12034 ( .A1(n13340), .A2(n22212), .ZN(n13356) );
  INV_X1 U12035 ( .A(n13321), .ZN(n13322) );
  NAND2_X1 U12036 ( .A1(n13302), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13321) );
  AND3_X1 U12037 ( .A1(n13306), .A2(n13305), .A3(n13304), .ZN(n16052) );
  NOR2_X1 U12038 ( .A1(n11388), .A2(n11386), .ZN(n11385) );
  INV_X1 U12039 ( .A(n15531), .ZN(n11386) );
  AND2_X1 U12040 ( .A1(n13226), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13227) );
  INV_X1 U12041 ( .A(n13205), .ZN(n13112) );
  NAND2_X1 U12042 ( .A1(n13112), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13140) );
  NAND2_X1 U12043 ( .A1(n13206), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13205) );
  NOR2_X1 U12044 ( .A1(n13196), .A2(n22119), .ZN(n13206) );
  CLKBUF_X1 U12045 ( .A(n14980), .Z(n14981) );
  NAND2_X1 U12046 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13178) );
  NOR2_X1 U12047 ( .A1(n13178), .A2(n14946), .ZN(n13188) );
  AOI21_X1 U12048 ( .B1(n14625), .B2(n13165), .A(n11518), .ZN(n13173) );
  NOR2_X1 U12049 ( .A1(n16910), .A2(n11516), .ZN(n16368) );
  INV_X1 U12050 ( .A(n11489), .ZN(n11351) );
  OR2_X1 U12051 ( .A1(n16771), .A2(n16759), .ZN(n11371) );
  NOR2_X1 U12052 ( .A1(n16825), .A2(n16793), .ZN(n16792) );
  NAND2_X1 U12053 ( .A1(n11370), .A2(n11241), .ZN(n16825) );
  NAND2_X1 U12054 ( .A1(n11481), .A2(n17256), .ZN(n11480) );
  NAND2_X1 U12055 ( .A1(n11482), .A2(n11242), .ZN(n11481) );
  NAND2_X1 U12056 ( .A1(n16830), .A2(n16829), .ZN(n17210) );
  NAND2_X1 U12057 ( .A1(n17061), .A2(n11483), .ZN(n11356) );
  NAND2_X1 U12058 ( .A1(n16005), .A2(n11364), .ZN(n17281) );
  AND2_X1 U12059 ( .A1(n15304), .A2(n15303), .ZN(n21992) );
  AND2_X1 U12060 ( .A1(n15346), .A2(n15345), .ZN(n15349) );
  AND2_X1 U12061 ( .A1(n15343), .A2(n15342), .ZN(n15459) );
  NAND2_X1 U12062 ( .A1(n11486), .A2(n11485), .ZN(n20754) );
  INV_X1 U12063 ( .A(n15583), .ZN(n11488) );
  OR2_X1 U12064 ( .A1(n15299), .A2(n15298), .ZN(n22030) );
  OR2_X1 U12065 ( .A1(n13029), .A2(n11361), .ZN(n12955) );
  OAI21_X1 U12066 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n13026), .A(
        n13025), .ZN(n13027) );
  OR2_X1 U12067 ( .A1(n13029), .A2(n12809), .ZN(n13035) );
  INV_X1 U12068 ( .A(n13069), .ZN(n11357) );
  BUF_X1 U12069 ( .A(n12911), .Z(n14462) );
  AND2_X1 U12070 ( .A1(n16722), .A2(n12947), .ZN(n14584) );
  INV_X1 U12071 ( .A(n15002), .ZN(n15034) );
  AND2_X1 U12072 ( .A1(n11196), .A2(n22280), .ZN(n15019) );
  AND2_X1 U12073 ( .A1(n15033), .A2(n14999), .ZN(n15020) );
  AND3_X1 U12074 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n22287), .A3(n14787), 
        .ZN(n22682) );
  INV_X1 U12075 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n15215) );
  INV_X1 U12076 ( .A(n15019), .ZN(n15415) );
  NAND2_X1 U12077 ( .A1(n11195), .A2(n13174), .ZN(n14841) );
  OR2_X1 U12078 ( .A1(n14775), .A2(n17060), .ZN(n22688) );
  AND2_X1 U12079 ( .A1(n14752), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17985) );
  NAND2_X1 U12080 ( .A1(n12589), .A2(n12641), .ZN(n14370) );
  OR2_X1 U12081 ( .A1(n15158), .A2(n12702), .ZN(n15166) );
  NAND2_X1 U12082 ( .A1(n12209), .A2(n12549), .ZN(n12558) );
  NOR2_X1 U12083 ( .A1(n12558), .A2(n12557), .ZN(n12562) );
  NAND2_X1 U12084 ( .A1(n12494), .A2(n12495), .ZN(n12499) );
  NOR2_X1 U12085 ( .A1(n12489), .A2(n12487), .ZN(n12494) );
  INV_X1 U12086 ( .A(n11347), .ZN(n12519) );
  NAND2_X1 U12087 ( .A1(n11347), .A2(n11346), .ZN(n12511) );
  INV_X1 U12088 ( .A(n12509), .ZN(n11346) );
  NAND2_X1 U12089 ( .A1(n12471), .A2(n12472), .ZN(n12513) );
  AND2_X1 U12090 ( .A1(n12459), .A2(n11338), .ZN(n12471) );
  NOR2_X1 U12091 ( .A1(n12468), .A2(n11339), .ZN(n11338) );
  INV_X1 U12092 ( .A(n11340), .ZN(n11339) );
  NOR2_X1 U12093 ( .A1(n20174), .A2(n12199), .ZN(n12468) );
  NAND2_X1 U12094 ( .A1(n12459), .A2(n11340), .ZN(n12470) );
  NOR2_X1 U12095 ( .A1(n11337), .A2(n11225), .ZN(n12446) );
  INV_X1 U12096 ( .A(n12413), .ZN(n11337) );
  INV_X1 U12097 ( .A(n14766), .ZN(n11511) );
  NOR3_X1 U12098 ( .A1(n17374), .A2(n12188), .A3(n16641), .ZN(n16659) );
  AND2_X1 U12099 ( .A1(n11238), .A2(n11499), .ZN(n11498) );
  NAND2_X1 U12100 ( .A1(n11502), .A2(n11500), .ZN(n11499) );
  INV_X1 U12101 ( .A(n17353), .ZN(n11409) );
  NAND2_X1 U12102 ( .A1(n17740), .A2(n12781), .ZN(n17352) );
  AND3_X1 U12104 ( .A1(n12155), .A2(n12154), .A3(n12153), .ZN(n15317) );
  AND3_X1 U12105 ( .A1(n12071), .A2(n12070), .A3(n12069), .ZN(n14737) );
  NAND2_X1 U12106 ( .A1(n12019), .A2(n11996), .ZN(n12020) );
  INV_X1 U12107 ( .A(n14619), .ZN(n11998) );
  AND2_X1 U12108 ( .A1(n14720), .A2(n14719), .ZN(n14721) );
  AND2_X1 U12109 ( .A1(n16597), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14740) );
  INV_X1 U12110 ( .A(n14566), .ZN(n11423) );
  AND2_X1 U12111 ( .A1(n14266), .A2(n19084), .ZN(n18147) );
  INV_X1 U12112 ( .A(n14536), .ZN(n14413) );
  INV_X1 U12113 ( .A(n16030), .ZN(n16139) );
  NAND2_X1 U12114 ( .A1(n17402), .A2(n11405), .ZN(n17385) );
  CLKBUF_X1 U12115 ( .A(n12235), .Z(n12271) );
  NAND2_X1 U12116 ( .A1(n11399), .A2(n12770), .ZN(n11398) );
  INV_X1 U12117 ( .A(n16216), .ZN(n11399) );
  NAND2_X1 U12118 ( .A1(n15569), .A2(n11224), .ZN(n16189) );
  INV_X1 U12119 ( .A(n16186), .ZN(n11401) );
  NOR2_X1 U12120 ( .A1(n16189), .A2(n16181), .ZN(n16194) );
  NAND2_X1 U12121 ( .A1(n15569), .A2(n11222), .ZN(n16187) );
  NOR2_X1 U12122 ( .A1(n15539), .A2(n15538), .ZN(n15569) );
  INV_X1 U12123 ( .A(n17635), .ZN(n11470) );
  AOI21_X1 U12124 ( .B1(n12572), .B2(n12019), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12795) );
  INV_X1 U12125 ( .A(n12563), .ZN(n11459) );
  INV_X1 U12126 ( .A(n11214), .ZN(n11458) );
  OR2_X1 U12127 ( .A1(n14036), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11536) );
  INV_X1 U12128 ( .A(n14035), .ZN(n14034) );
  INV_X1 U12129 ( .A(n12566), .ZN(n11461) );
  AND2_X1 U12130 ( .A1(n17402), .A2(n11403), .ZN(n14082) );
  AND2_X1 U12131 ( .A1(n11405), .A2(n11404), .ZN(n11403) );
  INV_X1 U12132 ( .A(n14083), .ZN(n11404) );
  NOR2_X1 U12133 ( .A1(n19306), .A2(n12685), .ZN(n14038) );
  NOR2_X1 U12134 ( .A1(n14037), .A2(n14036), .ZN(n17483) );
  NAND2_X1 U12135 ( .A1(n19295), .A2(n12019), .ZN(n12551) );
  OR2_X1 U12136 ( .A1(n12567), .A2(n17691), .ZN(n17508) );
  OR2_X1 U12137 ( .A1(n11474), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11472) );
  AND2_X1 U12138 ( .A1(n11474), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11473) );
  NAND2_X1 U12139 ( .A1(n19283), .A2(n12019), .ZN(n17520) );
  OR2_X1 U12140 ( .A1(n14104), .A2(n14106), .ZN(n17401) );
  NAND2_X1 U12141 ( .A1(n11430), .A2(n12693), .ZN(n17537) );
  OR2_X1 U12142 ( .A1(n19272), .A2(n12685), .ZN(n12757) );
  NAND2_X1 U12143 ( .A1(n17580), .A2(n12753), .ZN(n12754) );
  OR2_X1 U12144 ( .A1(n12764), .A2(n17815), .ZN(n11323) );
  AND2_X1 U12145 ( .A1(n12753), .A2(n12508), .ZN(n17591) );
  AND3_X1 U12146 ( .A1(n12106), .A2(n12105), .A3(n12104), .ZN(n14996) );
  AND3_X1 U12147 ( .A1(n12042), .A2(n12041), .A3(n12040), .ZN(n14644) );
  NAND2_X1 U12148 ( .A1(n12675), .A2(n12674), .ZN(n17912) );
  NAND2_X1 U12149 ( .A1(n17912), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17911) );
  NAND2_X1 U12150 ( .A1(n12663), .A2(n11475), .ZN(n16068) );
  NAND2_X1 U12151 ( .A1(n11313), .A2(n12662), .ZN(n16067) );
  AND2_X1 U12152 ( .A1(n12668), .A2(n12661), .ZN(n11313) );
  AOI21_X1 U12153 ( .B1(n12287), .B2(n12286), .A(n11744), .ZN(n14742) );
  INV_X1 U12154 ( .A(n15396), .ZN(n12652) );
  INV_X1 U12155 ( .A(n15395), .ZN(n11312) );
  OR2_X1 U12156 ( .A1(n12746), .A2(n15161), .ZN(n17923) );
  OR2_X1 U12157 ( .A1(n12746), .A2(n12716), .ZN(n17787) );
  XNOR2_X1 U12158 ( .A(n14380), .B(n11882), .ZN(n14471) );
  AND2_X1 U12159 ( .A1(n11897), .A2(n11896), .ZN(n14470) );
  CLKBUF_X1 U12160 ( .A(n11863), .Z(n11864) );
  INV_X1 U12161 ( .A(n12356), .ZN(n16023) );
  NOR2_X1 U12162 ( .A1(n20074), .A2(n19944), .ZN(n20097) );
  INV_X1 U12163 ( .A(n12364), .ZN(n20021) );
  INV_X1 U12164 ( .A(n12313), .ZN(n12295) );
  INV_X1 U12165 ( .A(n12367), .ZN(n19954) );
  NAND2_X1 U12166 ( .A1(n20086), .A2(n20100), .ZN(n19985) );
  NAND2_X1 U12167 ( .A1(n11592), .A2(n11571), .ZN(n11599) );
  NAND2_X1 U12168 ( .A1(n11597), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11598) );
  AND2_X1 U12169 ( .A1(n19944), .A2(n20081), .ZN(n20042) );
  INV_X1 U12170 ( .A(n20232), .ZN(n20428) );
  INV_X1 U12171 ( .A(n11143), .ZN(n20433) );
  AND2_X1 U12172 ( .A1(n21221), .A2(n21146), .ZN(n21222) );
  NOR2_X1 U12173 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n20958), .ZN(n20974) );
  AOI22_X1 U12174 ( .A1(n18480), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n18546), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18482) );
  AOI22_X1 U12175 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18546), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18327) );
  AOI21_X1 U12176 ( .B1(n18497), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n11284), .ZN(n18390) );
  AOI21_X1 U12177 ( .B1(n11159), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n11268), .ZN(n18434) );
  NOR2_X1 U12178 ( .A1(n11259), .A2(n11269), .ZN(n11268) );
  INV_X1 U12179 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11269) );
  AOI21_X1 U12180 ( .B1(n20948), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n11292), .ZN(n18493) );
  NOR2_X1 U12181 ( .A1(n11259), .A2(n11293), .ZN(n11292) );
  INV_X1 U12182 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11293) );
  AOI21_X1 U12183 ( .B1(n11156), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n11282), .ZN(n18516) );
  NOR2_X1 U12184 ( .A1(n11259), .A2(n11283), .ZN(n11282) );
  INV_X1 U12185 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11283) );
  AOI22_X1 U12186 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18546), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18244) );
  AOI22_X1 U12187 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18546), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16251) );
  AOI21_X1 U12188 ( .B1(n11156), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n11274), .ZN(n18282) );
  NOR2_X1 U12189 ( .A1(n11259), .A2(n11275), .ZN(n11274) );
  INV_X1 U12190 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11275) );
  AOI21_X1 U12191 ( .B1(n18279), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n11294), .ZN(n18219) );
  NOR2_X1 U12192 ( .A1(n11259), .A2(n11295), .ZN(n11294) );
  INV_X1 U12193 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11295) );
  AOI21_X1 U12194 ( .B1(n18523), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n11276), .ZN(n13713) );
  NOR2_X1 U12195 ( .A1(n18254), .A2(n11277), .ZN(n11276) );
  INV_X1 U12196 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11277) );
  AND2_X1 U12197 ( .A1(n13758), .A2(n13757), .ZN(n13759) );
  NOR2_X1 U12198 ( .A1(n14159), .A2(n13715), .ZN(n13710) );
  NAND2_X1 U12199 ( .A1(n18523), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11244) );
  NAND2_X1 U12200 ( .A1(n18522), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11247) );
  NAND2_X1 U12201 ( .A1(n18547), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11245) );
  NOR2_X1 U12202 ( .A1(n18568), .A2(n17952), .ZN(n19028) );
  NAND2_X1 U12203 ( .A1(n18753), .A2(n14031), .ZN(n18744) );
  INV_X1 U12204 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18633) );
  NAND2_X1 U12205 ( .A1(n13822), .A2(n11436), .ZN(n18904) );
  INV_X1 U12206 ( .A(n18682), .ZN(n18776) );
  NOR2_X1 U12207 ( .A1(n21337), .A2(n21964), .ZN(n14124) );
  INV_X1 U12208 ( .A(n14031), .ZN(n18800) );
  INV_X1 U12209 ( .A(n14016), .ZN(n11444) );
  NOR2_X1 U12210 ( .A1(n18645), .A2(n21739), .ZN(n11447) );
  INV_X1 U12211 ( .A(n18718), .ZN(n11446) );
  NOR2_X1 U12212 ( .A1(n21825), .A2(n21740), .ZN(n18736) );
  NAND2_X1 U12213 ( .A1(n21566), .A2(n18705), .ZN(n21825) );
  NAND2_X1 U12214 ( .A1(n18668), .A2(n13837), .ZN(n18719) );
  NOR2_X1 U12215 ( .A1(n21869), .A2(n14025), .ZN(n21566) );
  NAND2_X1 U12216 ( .A1(n21724), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n21869) );
  NAND2_X1 U12217 ( .A1(n13832), .A2(n13831), .ZN(n13833) );
  NAND2_X1 U12218 ( .A1(n13834), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13832) );
  NAND2_X1 U12219 ( .A1(n18825), .A2(n21882), .ZN(n18824) );
  NAND2_X1 U12220 ( .A1(n18876), .A2(n13829), .ZN(n18847) );
  INV_X1 U12221 ( .A(n13826), .ZN(n14121) );
  NAND2_X1 U12222 ( .A1(n18894), .A2(n13828), .ZN(n18877) );
  NAND2_X1 U12223 ( .A1(n18877), .A2(n18878), .ZN(n18876) );
  XNOR2_X1 U12224 ( .A(n13826), .B(n11451), .ZN(n18895) );
  INV_X1 U12225 ( .A(n13827), .ZN(n11451) );
  NAND2_X1 U12226 ( .A1(n18895), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18894) );
  NAND2_X1 U12227 ( .A1(n18900), .A2(n13958), .ZN(n18892) );
  XNOR2_X1 U12228 ( .A(n13952), .B(n21625), .ZN(n18927) );
  NAND2_X1 U12229 ( .A1(n18927), .A2(n18926), .ZN(n18925) );
  XNOR2_X1 U12230 ( .A(n13814), .B(n21626), .ZN(n18940) );
  NAND2_X1 U12231 ( .A1(n18940), .A2(n18939), .ZN(n18938) );
  AOI211_X1 U12232 ( .C1(n18279), .C2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A(
        n13851), .B(n13850), .ZN(n13852) );
  AOI21_X1 U12233 ( .B1(n14005), .B2(n14007), .A(n14004), .ZN(n14129) );
  INV_X1 U12234 ( .A(n21525), .ZN(n18968) );
  INV_X1 U12235 ( .A(n14146), .ZN(n14155) );
  NAND2_X1 U12236 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14146) );
  INV_X1 U12237 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19530) );
  NOR2_X1 U12238 ( .A1(n13864), .A2(n13863), .ZN(n19645) );
  NOR2_X1 U12239 ( .A1(n13894), .A2(n13893), .ZN(n21405) );
  INV_X1 U12240 ( .A(n22210), .ZN(n22200) );
  INV_X1 U12241 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n15457) );
  INV_X1 U12242 ( .A(n22269), .ZN(n22253) );
  INV_X1 U12243 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n22119) );
  INV_X1 U12244 ( .A(n22266), .ZN(n22257) );
  AND2_X1 U12245 ( .A1(n22091), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n22264) );
  AND2_X2 U12246 ( .A1(n14425), .A2(n14424), .ZN(n20727) );
  CLKBUF_X1 U12247 ( .A(n13703), .Z(n16892) );
  INV_X1 U12248 ( .A(n16149), .ZN(n16891) );
  INV_X1 U12249 ( .A(n16054), .ZN(n16890) );
  INV_X1 U12250 ( .A(n16056), .ZN(n16008) );
  BUF_X1 U12251 ( .A(n20620), .Z(n20632) );
  NOR2_X1 U12252 ( .A1(n20633), .A2(n20604), .ZN(n20620) );
  INV_X1 U12253 ( .A(n14587), .ZN(n22384) );
  OR2_X1 U12254 ( .A1(n15064), .A2(n16906), .ZN(n15065) );
  OR2_X1 U12255 ( .A1(n16263), .A2(n16264), .ZN(n16266) );
  INV_X1 U12256 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14946) );
  NAND2_X1 U12257 ( .A1(n22277), .A2(n14630), .ZN(n20728) );
  OR2_X1 U12258 ( .A1(n22289), .A2(n22468), .ZN(n17060) );
  INV_X1 U12259 ( .A(n17060), .ZN(n20762) );
  AOI21_X1 U12260 ( .B1(n16901), .B2(n17256), .A(n16911), .ZN(n16902) );
  NAND2_X1 U12261 ( .A1(n11491), .A2(n16919), .ZN(n16941) );
  NAND2_X1 U12262 ( .A1(n20748), .A2(n20747), .ZN(n20746) );
  NAND2_X1 U12263 ( .A1(n20740), .A2(n15583), .ZN(n20748) );
  NOR2_X1 U12264 ( .A1(n14931), .A2(n14856), .ZN(n14861) );
  INV_X1 U12265 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n14752) );
  NOR2_X1 U12266 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n17940) );
  OAI21_X1 U12267 ( .B1(n15036), .B2(n22391), .A(n15035), .ZN(n22698) );
  OAI21_X1 U12268 ( .B1(n15420), .B2(n22715), .A(n22480), .ZN(n22718) );
  OAI211_X1 U12269 ( .C1(n14188), .C2(n22744), .A(n15256), .B(n22410), .ZN(
        n22747) );
  AOI22_X1 U12270 ( .A1(n22475), .A2(n22485), .B1(n22474), .B2(n22473), .ZN(
        n22777) );
  INV_X1 U12271 ( .A(n15222), .ZN(n22490) );
  INV_X1 U12272 ( .A(n22546), .ZN(n22555) );
  INV_X1 U12273 ( .A(n22769), .ZN(n22792) );
  NOR2_X1 U12274 ( .A1(n16719), .A2(n14188), .ZN(n22296) );
  NOR2_X1 U12275 ( .A1(n15166), .A2(n19448), .ZN(n19074) );
  AND3_X1 U12276 ( .A1(n17963), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n19078) );
  AOI21_X1 U12277 ( .B1(n12227), .B2(n19348), .A(n12226), .ZN(n12228) );
  XNOR2_X1 U12278 ( .A(n12550), .B(n12549), .ZN(n19295) );
  NAND2_X1 U12279 ( .A1(n12542), .A2(n12547), .ZN(n12556) );
  INV_X1 U12280 ( .A(n19310), .ZN(n19349) );
  NAND2_X1 U12281 ( .A1(n15533), .A2(n11505), .ZN(n11504) );
  INV_X1 U12282 ( .A(n11507), .ZN(n11505) );
  INV_X1 U12283 ( .A(n17428), .ZN(n17417) );
  OR2_X1 U12284 ( .A1(n17423), .A2(n14581), .ZN(n17428) );
  OR2_X1 U12285 ( .A1(n16651), .A2(n16650), .ZN(n19337) );
  NAND2_X1 U12286 ( .A1(n16172), .A2(n16132), .ZN(n17768) );
  INV_X1 U12287 ( .A(n20164), .ZN(n15324) );
  INV_X1 U12288 ( .A(n17477), .ZN(n20321) );
  NOR2_X1 U12289 ( .A1(n18147), .A2(n18180), .ZN(n18159) );
  CLKBUF_X1 U12290 ( .A(n18168), .Z(n18180) );
  CLKBUF_X1 U12291 ( .A(n18159), .Z(n18179) );
  INV_X1 U12292 ( .A(n14549), .ZN(n14418) );
  NAND2_X1 U12293 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11322) );
  INV_X1 U12294 ( .A(n11323), .ZN(n17605) );
  NAND2_X1 U12295 ( .A1(n17898), .A2(n12684), .ZN(n18061) );
  INV_X1 U12296 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17641) );
  INV_X1 U12297 ( .A(n18070), .ZN(n18112) );
  NAND2_X1 U12298 ( .A1(n19451), .A2(n12766), .ZN(n18076) );
  AND2_X1 U12299 ( .A1(n18076), .A2(n16341), .ZN(n18070) );
  AOI21_X1 U12300 ( .B1(n19347), .B2(n19408), .A(n11416), .ZN(n11531) );
  NAND2_X1 U12301 ( .A1(n12735), .A2(n11417), .ZN(n11416) );
  INV_X1 U12302 ( .A(n16397), .ZN(n11417) );
  OR2_X1 U12303 ( .A1(n17793), .A2(n12726), .ZN(n17727) );
  NOR2_X1 U12304 ( .A1(n17556), .A2(n17550), .ZN(n17549) );
  NAND2_X1 U12305 ( .A1(n17639), .A2(n17638), .ZN(n17898) );
  INV_X1 U12306 ( .A(n18033), .ZN(n15133) );
  INV_X1 U12307 ( .A(n17928), .ZN(n19408) );
  INV_X1 U12308 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20094) );
  INV_X1 U12309 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20092) );
  INV_X1 U12310 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19998) );
  NAND2_X1 U12311 ( .A1(n11424), .A2(n11207), .ZN(n14567) );
  NAND2_X1 U12312 ( .A1(n14379), .A2(n14378), .ZN(n19929) );
  INV_X1 U12313 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20083) );
  XNOR2_X1 U12314 ( .A(n14716), .B(n14608), .ZN(n18127) );
  NAND2_X1 U12315 ( .A1(n16020), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19435) );
  OR2_X1 U12316 ( .A1(n14731), .A2(n14732), .ZN(n14734) );
  NOR2_X1 U12317 ( .A1(n20074), .A2(n20073), .ZN(n20524) );
  AND2_X1 U12318 ( .A1(n20028), .A2(n20015), .ZN(n20404) );
  NAND2_X1 U12319 ( .A1(n19982), .A2(n20027), .ZN(n20480) );
  OAI21_X1 U12320 ( .B1(n19978), .B2(n19977), .A(n19976), .ZN(n20468) );
  INV_X1 U12321 ( .A(n20478), .ZN(n20467) );
  INV_X1 U12322 ( .A(n20371), .ZN(n20375) );
  INV_X1 U12323 ( .A(n20455), .ZN(n20452) );
  NAND2_X1 U12324 ( .A1(n19941), .A2(n20015), .ZN(n20445) );
  INV_X1 U12325 ( .A(n20109), .ZN(n20107) );
  INV_X1 U12326 ( .A(n20537), .ZN(n20530) );
  INV_X1 U12327 ( .A(n20249), .ZN(n20270) );
  NAND2_X1 U12328 ( .A1(n19941), .A2(n19964), .ZN(n20439) );
  INV_X1 U12329 ( .A(n20216), .ZN(n20211) );
  INV_X1 U12330 ( .A(n20156), .ZN(n20153) );
  NAND2_X1 U12331 ( .A1(n19941), .A2(n20042), .ZN(n20540) );
  OAI22_X1 U12332 ( .A1(n22680), .A2(n20433), .B1(n19922), .B2(n20432), .ZN(
        n20109) );
  CLKBUF_X1 U12333 ( .A(n18207), .Z(n18202) );
  NAND2_X1 U12334 ( .A1(n20906), .A2(n20905), .ZN(n21162) );
  OR2_X1 U12335 ( .A1(n20946), .A2(P3_EBX_REG_4__SCAN_IN), .ZN(n20958) );
  INV_X1 U12336 ( .A(n20899), .ZN(n20897) );
  INV_X1 U12337 ( .A(n21287), .ZN(n21330) );
  INV_X1 U12338 ( .A(n21303), .ZN(n21331) );
  INV_X1 U12339 ( .A(n21119), .ZN(n21329) );
  INV_X1 U12340 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18563) );
  INV_X1 U12341 ( .A(n21474), .ZN(n21470) );
  NAND2_X1 U12342 ( .A1(n21470), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n21469) );
  INV_X1 U12343 ( .A(n21480), .ZN(n21444) );
  NAND2_X1 U12344 ( .A1(n21444), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n21449) );
  NOR2_X1 U12345 ( .A1(n21443), .A2(n21486), .ZN(n21481) );
  NOR2_X1 U12346 ( .A1(n21505), .A2(n21504), .ZN(n21503) );
  NOR2_X1 U12347 ( .A1(n13745), .A2(n13744), .ZN(n21391) );
  INV_X1 U12348 ( .A(n21527), .ZN(n21394) );
  INV_X1 U12349 ( .A(n13767), .ZN(n11450) );
  NOR2_X1 U12350 ( .A1(n21369), .A2(n21344), .ZN(n21527) );
  NOR2_X1 U12351 ( .A1(n19015), .A2(n19028), .ZN(n19037) );
  CLKBUF_X1 U12352 ( .A(n19037), .Z(n19044) );
  BUF_X1 U12353 ( .A(n20878), .Z(n20891) );
  CLKBUF_X1 U12355 ( .A(n20908), .Z(n21146) );
  INV_X1 U12356 ( .A(n18796), .ZN(n21794) );
  NOR2_X1 U12357 ( .A1(n18771), .A2(n21760), .ZN(n18793) );
  NAND2_X1 U12358 ( .A1(n18740), .A2(n11258), .ZN(n18771) );
  AND2_X1 U12359 ( .A1(n21756), .A2(n18741), .ZN(n11258) );
  NOR2_X1 U12360 ( .A1(n18643), .A2(n18590), .ZN(n18740) );
  AOI21_X1 U12361 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18682), .A(
        n19814), .ZN(n18726) );
  NOR2_X1 U12362 ( .A1(n18633), .A2(n18634), .ZN(n21074) );
  INV_X1 U12363 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18634) );
  OAI22_X1 U12364 ( .A1(n18839), .A2(n21870), .B1(n21670), .B2(n18974), .ZN(
        n18869) );
  AOI21_X1 U12365 ( .B1(n20833), .B2(n21960), .A(n14116), .ZN(n18957) );
  INV_X1 U12366 ( .A(n18957), .ZN(n18970) );
  OR2_X1 U12367 ( .A1(n21964), .A2(n20904), .ZN(n18974) );
  OAI21_X1 U12368 ( .B1(n14017), .B2(n18845), .A(n11432), .ZN(n11431) );
  NAND2_X1 U12369 ( .A1(n21780), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11432) );
  INV_X1 U12370 ( .A(n21899), .ZN(n21843) );
  NOR2_X1 U12371 ( .A1(n13966), .A2(n11254), .ZN(n13969) );
  NAND2_X1 U12372 ( .A1(n11255), .A2(n11257), .ZN(n11254) );
  AND2_X1 U12373 ( .A1(n11304), .A2(n21911), .ZN(n21899) );
  NOR2_X1 U12374 ( .A1(n21693), .A2(n18834), .ZN(n21724) );
  INV_X1 U12375 ( .A(n21927), .ZN(n21871) );
  NAND2_X1 U12376 ( .A1(n18915), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18914) );
  NAND2_X1 U12377 ( .A1(n11443), .A2(n11440), .ZN(n18915) );
  NAND2_X1 U12378 ( .A1(n21899), .A2(n20904), .ZN(n21614) );
  NAND2_X1 U12379 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21549) );
  INV_X2 U12380 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21559) );
  AND2_X1 U12381 ( .A1(n13702), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14775)
         );
  NAND2_X1 U12383 ( .A1(n16380), .A2(n13692), .ZN(n13709) );
  AND2_X1 U12384 ( .A1(n16693), .A2(n16692), .ZN(n11497) );
  AND2_X1 U12385 ( .A1(n16403), .A2(n16402), .ZN(n16404) );
  AOI21_X1 U12386 ( .B1(n16401), .B2(n18095), .A(n16400), .ZN(n16402) );
  AOI21_X1 U12387 ( .B1(n16411), .B2(n18095), .A(n16410), .ZN(n16412) );
  NAND2_X1 U12388 ( .A1(n11393), .A2(n11392), .ZN(n16707) );
  INV_X1 U12389 ( .A(n16706), .ZN(n11392) );
  OAI21_X1 U12390 ( .B1(n12788), .B2(n18103), .A(n12774), .ZN(n12775) );
  OR2_X1 U12391 ( .A1(n16686), .A2(n19416), .ZN(n12805) );
  OAI21_X1 U12392 ( .B1(n17656), .B2(n19416), .A(n17655), .ZN(n17657) );
  OAI21_X1 U12393 ( .B1(n12788), .B2(n19375), .A(n12787), .ZN(n12789) );
  AOI21_X1 U12394 ( .B1(n18797), .B2(n21803), .A(n11250), .ZN(n11249) );
  OR2_X1 U12395 ( .A1(n18816), .A2(n21803), .ZN(n11248) );
  OR2_X1 U12396 ( .A1(n21811), .A2(n18881), .ZN(n11252) );
  CLKBUF_X3 U12397 ( .A(n13916), .Z(n18388) );
  NAND2_X1 U12398 ( .A1(n11506), .A2(n15370), .ZN(n15446) );
  AND2_X1 U12399 ( .A1(n11203), .A2(n14108), .ZN(n11197) );
  AND2_X1 U12400 ( .A1(n11183), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12062) );
  NAND2_X1 U12401 ( .A1(n11185), .A2(n14319), .ZN(n11359) );
  NAND2_X1 U12402 ( .A1(n17410), .A2(n17411), .ZN(n17406) );
  NAND2_X1 U12403 ( .A1(n11387), .A2(n11385), .ZN(n15530) );
  OR2_X1 U12404 ( .A1(n16790), .A2(n11383), .ZN(n11198) );
  NAND2_X1 U12405 ( .A1(n16833), .A2(n11223), .ZN(n16826) );
  NAND2_X1 U12406 ( .A1(n14489), .A2(n20835), .ZN(n21911) );
  OAI21_X1 U12407 ( .B1(n17410), .B2(n11503), .A(n11498), .ZN(n17398) );
  XNOR2_X1 U12408 ( .A(n17398), .B(n16553), .ZN(n17393) );
  INV_X1 U12409 ( .A(n16031), .ZN(n11677) );
  AND2_X1 U12410 ( .A1(n11431), .A2(n21897), .ZN(n11199) );
  OR2_X1 U12411 ( .A1(n16770), .A2(n16771), .ZN(n11200) );
  NAND2_X1 U12412 ( .A1(n17740), .A2(n11197), .ZN(n14107) );
  INV_X1 U12413 ( .A(n11421), .ZN(n14084) );
  NAND2_X1 U12414 ( .A1(n13168), .A2(n13166), .ZN(n13176) );
  AND2_X1 U12415 ( .A1(n12449), .A2(n11470), .ZN(n11201) );
  NAND2_X1 U12416 ( .A1(n14623), .A2(n14622), .ZN(n14621) );
  AND2_X1 U12417 ( .A1(n14818), .A2(n11411), .ZN(n14995) );
  AND2_X1 U12418 ( .A1(n16129), .A2(n11233), .ZN(n16432) );
  OR2_X1 U12419 ( .A1(n15194), .A2(n11396), .ZN(n11202) );
  AND2_X1 U12420 ( .A1(n11409), .A2(n12781), .ZN(n11203) );
  OR2_X1 U12421 ( .A1(n13242), .A2(n13230), .ZN(n11204) );
  OR2_X1 U12422 ( .A1(n12038), .A2(n12037), .ZN(n14991) );
  OR2_X1 U12423 ( .A1(n12039), .A2(n11510), .ZN(n11205) );
  INV_X2 U12424 ( .A(n16497), .ZN(n11857) );
  NAND2_X2 U12425 ( .A1(n14297), .A2(n16710), .ZN(n14857) );
  NOR2_X1 U12426 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14151), .ZN(
        n18331) );
  INV_X1 U12427 ( .A(n12897), .ZN(n13560) );
  NAND2_X1 U12428 ( .A1(n12389), .A2(n12679), .ZN(n11475) );
  NAND3_X1 U12429 ( .A1(n14469), .A2(n11917), .A3(n11916), .ZN(n11207) );
  NAND2_X1 U12430 ( .A1(n12290), .A2(n12289), .ZN(n12288) );
  INV_X1 U12431 ( .A(n13821), .ZN(n13819) );
  NAND2_X2 U12432 ( .A1(n11494), .A2(n11492), .ZN(n11659) );
  NAND2_X1 U12433 ( .A1(n12500), .A2(n12501), .ZN(n12490) );
  AND2_X1 U12434 ( .A1(n16833), .A2(n11374), .ZN(n16823) );
  NOR2_X1 U12435 ( .A1(n16790), .A2(n11381), .ZN(n16756) );
  AND2_X1 U12436 ( .A1(n11430), .A2(n11429), .ZN(n11208) );
  NOR2_X1 U12437 ( .A1(n16790), .A2(n16791), .ZN(n16780) );
  AND2_X1 U12438 ( .A1(n12511), .A2(n12510), .ZN(n11210) );
  NOR2_X1 U12439 ( .A1(n16621), .A2(n16620), .ZN(n17373) );
  INV_X1 U12440 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11547) );
  NOR2_X1 U12441 ( .A1(n21337), .A2(n13937), .ZN(n13966) );
  AND2_X1 U12442 ( .A1(n14284), .A2(n14797), .ZN(n12940) );
  NAND2_X1 U12443 ( .A1(n16833), .A2(n16835), .ZN(n16800) );
  NAND2_X1 U12444 ( .A1(n16833), .A2(n11376), .ZN(n11211) );
  AND2_X1 U12445 ( .A1(n12312), .A2(n12308), .ZN(n12355) );
  XNOR2_X1 U12446 ( .A(n11309), .B(n12757), .ZN(n17548) );
  AND2_X1 U12447 ( .A1(n12315), .A2(n12303), .ZN(n12358) );
  NAND2_X1 U12448 ( .A1(n12947), .A2(n16710), .ZN(n16322) );
  INV_X1 U12449 ( .A(n12641), .ZN(n12581) );
  NAND2_X1 U12450 ( .A1(n12701), .A2(n12187), .ZN(n12800) );
  AND2_X1 U12451 ( .A1(n14714), .A2(n14720), .ZN(n14731) );
  NOR3_X1 U12452 ( .A1(n14031), .A2(n21868), .A3(n18745), .ZN(n11212) );
  NAND2_X1 U12453 ( .A1(n17394), .A2(n11534), .ZN(n16575) );
  XNOR2_X1 U12454 ( .A(n15584), .B(n13111), .ZN(n15593) );
  NAND2_X1 U12455 ( .A1(n12296), .A2(n12295), .ZN(n12367) );
  AND3_X1 U12456 ( .A1(n12758), .A2(n12755), .A3(n12522), .ZN(n11213) );
  NAND2_X1 U12457 ( .A1(n13614), .A2(n12933), .ZN(n12909) );
  AND2_X1 U12458 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11850) );
  AND2_X1 U12459 ( .A1(n14599), .A2(n14717), .ZN(n14716) );
  NAND2_X1 U12460 ( .A1(n11725), .A2(n11724), .ZN(n11726) );
  INV_X1 U12461 ( .A(n12684), .ZN(n11427) );
  AND2_X1 U12462 ( .A1(n12568), .A2(n17508), .ZN(n11214) );
  NOR2_X1 U12463 ( .A1(n16770), .A2(n11371), .ZN(n16746) );
  AND3_X1 U12464 ( .A1(n11544), .A2(n11545), .A3(n11496), .ZN(n11215) );
  NOR2_X1 U12465 ( .A1(n21404), .A2(n21405), .ZN(n13975) );
  INV_X1 U12466 ( .A(n13975), .ZN(n11300) );
  INV_X1 U12467 ( .A(n19727), .ZN(n14000) );
  NOR2_X1 U12468 ( .A1(n13905), .A2(n13904), .ZN(n19727) );
  AND4_X1 U12469 ( .A1(n11247), .A2(n11246), .A3(n11245), .A4(n11244), .ZN(
        n11216) );
  NAND2_X1 U12470 ( .A1(n12393), .A2(n12394), .ZN(n11217) );
  NAND2_X1 U12471 ( .A1(n17402), .A2(n17335), .ZN(n17334) );
  NAND2_X1 U12472 ( .A1(n11463), .A2(n11464), .ZN(n17611) );
  AND3_X1 U12473 ( .A1(n12759), .A2(n12537), .A3(n17561), .ZN(n11218) );
  OR2_X1 U12474 ( .A1(n13930), .A2(n19645), .ZN(n11219) );
  NAND2_X1 U12475 ( .A1(n12392), .A2(n19114), .ZN(n12416) );
  AND2_X1 U12476 ( .A1(n15592), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11220) );
  INV_X1 U12477 ( .A(n11601), .ZN(n11651) );
  INV_X1 U12478 ( .A(n11475), .ZN(n12668) );
  INV_X1 U12479 ( .A(n12685), .ZN(n12019) );
  INV_X1 U12480 ( .A(n21883), .ZN(n11304) );
  AND2_X1 U12481 ( .A1(n11876), .A2(n14377), .ZN(n11918) );
  INV_X1 U12482 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11287) );
  INV_X1 U12483 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11261) );
  NAND3_X1 U12484 ( .A1(n11476), .A2(n14183), .A3(n12949), .ZN(n13678) );
  AND2_X1 U12485 ( .A1(n13936), .A2(n14491), .ZN(n11221) );
  NOR2_X1 U12486 ( .A1(n15368), .A2(n11507), .ZN(n15534) );
  AND2_X2 U12487 ( .A1(n11639), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11905) );
  INV_X1 U12488 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11271) );
  INV_X1 U12489 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11358) );
  NOR2_X1 U12490 ( .A1(n15368), .A2(n11504), .ZN(n16115) );
  NAND2_X1 U12491 ( .A1(n12413), .A2(n12412), .ZN(n12390) );
  INV_X1 U12492 ( .A(n14761), .ZN(n13174) );
  NOR3_X1 U12493 ( .A1(n16195), .A2(n17424), .A3(n16216), .ZN(n12769) );
  AND2_X1 U12494 ( .A1(n16115), .A2(n16114), .ZN(n16129) );
  NOR2_X1 U12495 ( .A1(n15326), .A2(n11388), .ZN(n15529) );
  NAND2_X1 U12496 ( .A1(n15569), .A2(n15568), .ZN(n15567) );
  NAND2_X1 U12497 ( .A1(n11387), .A2(n13230), .ZN(n15619) );
  NOR2_X2 U12498 ( .A1(n12241), .A2(n12768), .ZN(n12242) );
  NAND2_X1 U12499 ( .A1(n16005), .A2(n15555), .ZN(n16155) );
  AND2_X1 U12500 ( .A1(n15568), .A2(n11402), .ZN(n11222) );
  AND2_X1 U12501 ( .A1(n16129), .A2(n16131), .ZN(n16210) );
  NAND2_X1 U12502 ( .A1(n16129), .A2(n11513), .ZN(n16233) );
  NOR2_X1 U12503 ( .A1(n15530), .A2(n16052), .ZN(n16051) );
  AND2_X1 U12504 ( .A1(n16711), .A2(n12942), .ZN(n14280) );
  AND2_X1 U12505 ( .A1(n13388), .A2(n11376), .ZN(n11223) );
  NAND2_X1 U12506 ( .A1(n17913), .A2(n12449), .ZN(n17634) );
  MUX2_X1 U12507 ( .A(n12626), .B(P2_EBX_REG_3__SCAN_IN), .S(n12211), .Z(
        n12407) );
  INV_X1 U12508 ( .A(n15326), .ZN(n11387) );
  NOR2_X2 U12509 ( .A1(n12239), .A2(n12232), .ZN(n12240) );
  XNOR2_X1 U12510 ( .A(n12416), .B(n16075), .ZN(n16081) );
  XNOR2_X1 U12511 ( .A(n16575), .B(n11533), .ZN(n17388) );
  OAI21_X1 U12512 ( .B1(n17406), .B2(n17407), .A(n11502), .ZN(n17397) );
  INV_X1 U12513 ( .A(n11370), .ZN(n17212) );
  NOR2_X1 U12514 ( .A1(n17210), .A2(n17209), .ZN(n11370) );
  NOR2_X1 U12515 ( .A1(n17336), .A2(n17442), .ZN(n11421) );
  INV_X1 U12516 ( .A(n15368), .ZN(n11506) );
  AND2_X1 U12517 ( .A1(n11222), .A2(n11401), .ZN(n11224) );
  OR2_X1 U12518 ( .A1(n12391), .A2(n11336), .ZN(n11225) );
  INV_X1 U12519 ( .A(n11400), .ZN(n16215) );
  NOR2_X1 U12520 ( .A1(n16195), .A2(n16216), .ZN(n11400) );
  AND2_X1 U12521 ( .A1(n17740), .A2(n11203), .ZN(n11226) );
  INV_X1 U12522 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11361) );
  AND2_X1 U12523 ( .A1(n11489), .A2(n16920), .ZN(n11227) );
  OR2_X1 U12524 ( .A1(n19420), .A2(n17786), .ZN(n11228) );
  AND2_X1 U12525 ( .A1(n11489), .A2(n16360), .ZN(n11229) );
  AND2_X1 U12526 ( .A1(n11410), .A2(n15319), .ZN(n11230) );
  AND2_X4 U12527 ( .A1(n12819), .A2(n12815), .ZN(n13244) );
  NOR2_X1 U12528 ( .A1(n12941), .A2(n22424), .ZN(n13156) );
  INV_X1 U12529 ( .A(n13156), .ZN(n13149) );
  INV_X1 U12530 ( .A(n21930), .ZN(n21897) );
  INV_X1 U12531 ( .A(n18755), .ZN(n18845) );
  INV_X1 U12532 ( .A(n18103), .ZN(n18095) );
  NAND2_X1 U12533 ( .A1(n12021), .A2(n12020), .ZN(n14623) );
  NAND2_X1 U12534 ( .A1(n11511), .A2(n11524), .ZN(n14989) );
  OR2_X1 U12535 ( .A1(n12746), .A2(n12745), .ZN(n19416) );
  INV_X1 U12536 ( .A(n19416), .ZN(n19398) );
  NAND2_X1 U12537 ( .A1(n14377), .A2(n20174), .ZN(n12152) );
  NAND2_X1 U12538 ( .A1(n14818), .A2(n14819), .ZN(n14820) );
  NOR2_X1 U12539 ( .A1(n14766), .A2(n11205), .ZN(n15191) );
  AND2_X2 U12540 ( .A1(n11848), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16226) );
  NAND2_X1 U12541 ( .A1(n14818), .A2(n11410), .ZN(n11231) );
  AND2_X2 U12542 ( .A1(n11848), .A2(n11571), .ZN(n16416) );
  NOR2_X1 U12543 ( .A1(n14769), .A2(n14863), .ZN(n14862) );
  NOR2_X1 U12544 ( .A1(n15194), .A2(n15195), .ZN(n15193) );
  AND2_X1 U12545 ( .A1(n14623), .A2(n11414), .ZN(n14643) );
  AND2_X1 U12546 ( .A1(n11420), .A2(n16132), .ZN(n11232) );
  AND2_X1 U12547 ( .A1(n13173), .A2(n13172), .ZN(n14867) );
  AND2_X1 U12548 ( .A1(n11513), .A2(n11512), .ZN(n11233) );
  AND2_X1 U12549 ( .A1(n11660), .A2(n11633), .ZN(n12709) );
  NAND2_X1 U12550 ( .A1(n14733), .A2(n14721), .ZN(n14739) );
  AND2_X1 U12551 ( .A1(n11511), .A2(n11509), .ZN(n11234) );
  NOR2_X1 U12552 ( .A1(n12554), .A2(n11343), .ZN(n11235) );
  AND2_X1 U12553 ( .A1(n11233), .A2(n17422), .ZN(n11236) );
  NOR2_X1 U12554 ( .A1(n15194), .A2(n11395), .ZN(n15447) );
  INV_X1 U12555 ( .A(n11503), .ZN(n11502) );
  NOR2_X1 U12556 ( .A1(n16532), .A2(n19079), .ZN(n11503) );
  AND2_X1 U12557 ( .A1(n16000), .A2(n15622), .ZN(n11237) );
  AND2_X1 U12558 ( .A1(n17399), .A2(n11501), .ZN(n11238) );
  AND2_X1 U12559 ( .A1(n11197), .A2(n11408), .ZN(n11239) );
  INV_X1 U12560 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11439) );
  NAND2_X1 U12561 ( .A1(n12179), .A2(n12178), .ZN(n11240) );
  NAND2_X1 U12562 ( .A1(n16287), .A2(n16286), .ZN(n11241) );
  INV_X1 U12563 ( .A(n11510), .ZN(n11509) );
  NAND2_X1 U12564 ( .A1(n11524), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11510) );
  INV_X1 U12565 ( .A(n15486), .ZN(n11508) );
  INV_X1 U12566 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11316) );
  NOR2_X1 U12567 ( .A1(n17198), .A2(n17244), .ZN(n11242) );
  INV_X1 U12568 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11267) );
  INV_X2 U12569 ( .A(U212), .ZN(n20812) );
  OAI22_X2 U12570 ( .A1(n22681), .A2(n22688), .B1(n22680), .B2(n22686), .ZN(
        n22786) );
  AOI22_X2 U12571 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n11143), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20424), .ZN(n20415) );
  NOR3_X2 U12572 ( .A1(n16139), .A2(n22310), .A3(n19985), .ZN(n20424) );
  NOR3_X2 U12573 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15215), .A3(
        n22441), .ZN(n22784) );
  NOR4_X4 U12574 ( .A1(n21537), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .A4(P3_STATEBS16_REG_SCAN_IN), .ZN(n21135)
         );
  NAND3_X1 U12575 ( .A1(n13809), .A2(n13810), .A3(n11216), .ZN(n11243) );
  NAND3_X1 U12576 ( .A1(n11252), .A2(n11249), .A3(n11248), .ZN(P3_U2800) );
  NAND2_X1 U12577 ( .A1(n18943), .A2(n18944), .ZN(n18942) );
  NAND4_X1 U12578 ( .A1(n20843), .A2(n11257), .A3(n14145), .A4(n11255), .ZN(
        n14140) );
  NOR2_X1 U12579 ( .A1(n14140), .A2(n13964), .ZN(n14147) );
  CLKBUF_X1 U12580 ( .A(n18254), .Z(n11259) );
  NOR2_X1 U12581 ( .A1(n13976), .A2(n21404), .ZN(n11296) );
  INV_X1 U12582 ( .A(n13933), .ZN(n11297) );
  NAND2_X1 U12583 ( .A1(n14142), .A2(n11299), .ZN(n11298) );
  OR2_X1 U12584 ( .A1(n13984), .A2(n13975), .ZN(n11303) );
  NAND2_X1 U12585 ( .A1(n17567), .A2(n17568), .ZN(n17559) );
  OR2_X1 U12586 ( .A1(n11309), .A2(n12757), .ZN(n11308) );
  AND2_X2 U12587 ( .A1(n12289), .A2(n12297), .ZN(n12300) );
  XNOR2_X2 U12588 ( .A(n12393), .B(n12394), .ZN(n15395) );
  OAI21_X2 U12589 ( .B1(n11314), .B2(n11315), .A(n11425), .ZN(n18059) );
  AND2_X2 U12590 ( .A1(n11317), .A2(n11318), .ZN(n12285) );
  NAND4_X1 U12591 ( .A1(n11317), .A2(n11318), .A3(n11728), .A4(n11729), .ZN(
        n11407) );
  NAND3_X1 U12592 ( .A1(n12294), .A2(n12293), .A3(n11716), .ZN(n11317) );
  INV_X1 U12593 ( .A(n11697), .ZN(n11319) );
  NAND2_X1 U12594 ( .A1(n12294), .A2(n12293), .ZN(n12289) );
  NAND2_X1 U12595 ( .A1(n11323), .A2(n11228), .ZN(n17790) );
  OAI22_X1 U12596 ( .A1(n11323), .A2(n19375), .B1(n17815), .B2(n17793), .ZN(
        n17803) );
  NAND3_X1 U12597 ( .A1(n11932), .A2(n11931), .A3(n11330), .ZN(n11329) );
  NAND2_X1 U12598 ( .A1(n11335), .A2(n11332), .ZN(n12450) );
  NAND3_X1 U12599 ( .A1(n11334), .A2(n12445), .A3(n12412), .ZN(n11333) );
  INV_X1 U12600 ( .A(n12407), .ZN(n11334) );
  NAND2_X1 U12601 ( .A1(n11862), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11496) );
  AOI22_X1 U12602 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11587) );
  AOI22_X1 U12603 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U12604 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U12605 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11642) );
  AOI22_X1 U12606 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U12607 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U12608 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U12609 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U12610 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11590) );
  AOI22_X1 U12611 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U12612 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11552) );
  AOI22_X1 U12613 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U12614 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11605) );
  AND2_X4 U12615 ( .A1(n11865), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11862) );
  NAND2_X1 U12616 ( .A1(n16918), .A2(n11227), .ZN(n11350) );
  OAI21_X1 U12617 ( .B1(n16359), .B2(n11351), .A(n11350), .ZN(n16940) );
  NOR2_X2 U12618 ( .A1(n16362), .A2(n16940), .ZN(n16933) );
  NAND2_X1 U12619 ( .A1(n16359), .A2(n16361), .ZN(n11491) );
  NAND2_X1 U12620 ( .A1(n16918), .A2(n16920), .ZN(n16361) );
  AND2_X1 U12621 ( .A1(n15585), .A2(n15602), .ZN(n11353) );
  NAND2_X2 U12622 ( .A1(n16092), .A2(n16091), .ZN(n17061) );
  AND2_X2 U12623 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14508) );
  AND2_X2 U12624 ( .A1(n11358), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12819) );
  AND3_X2 U12625 ( .A1(n12907), .A2(n12906), .A3(n11360), .ZN(n14319) );
  NAND2_X1 U12626 ( .A1(n15332), .A2(n15331), .ZN(n20699) );
  NAND2_X1 U12627 ( .A1(n11368), .A2(n11366), .ZN(n15328) );
  INV_X1 U12628 ( .A(n14931), .ZN(n11368) );
  NAND2_X1 U12629 ( .A1(n11369), .A2(n14684), .ZN(n14856) );
  NOR2_X2 U12630 ( .A1(n16839), .A2(n16805), .ZN(n16830) );
  NAND2_X2 U12631 ( .A1(n16747), .A2(n16305), .ZN(n16736) );
  AND2_X2 U12632 ( .A1(n16300), .A2(n16746), .ZN(n16747) );
  NAND3_X1 U12633 ( .A1(n12892), .A2(n12891), .A3(n11372), .ZN(n12893) );
  INV_X1 U12634 ( .A(n13166), .ZN(n13167) );
  NAND2_X2 U12635 ( .A1(n11373), .A2(n14748), .ZN(n22418) );
  NAND3_X1 U12636 ( .A1(n16711), .A2(n16710), .A3(n12942), .ZN(n13689) );
  NAND2_X1 U12637 ( .A1(n16263), .A2(n16264), .ZN(n16265) );
  NAND2_X1 U12638 ( .A1(n16263), .A2(n11389), .ZN(n16729) );
  INV_X1 U12639 ( .A(n12396), .ZN(n12646) );
  NAND2_X1 U12640 ( .A1(n11996), .A2(n12396), .ZN(n11875) );
  NAND2_X1 U12641 ( .A1(n14818), .A2(n11230), .ZN(n15316) );
  NAND2_X1 U12642 ( .A1(n14623), .A2(n11413), .ZN(n14668) );
  NOR2_X2 U12643 ( .A1(n14085), .A2(n14050), .ZN(n16649) );
  NAND2_X1 U12644 ( .A1(n11207), .A2(n11423), .ZN(n11422) );
  NAND2_X1 U12645 ( .A1(n16069), .A2(n16067), .ZN(n12677) );
  NAND2_X1 U12646 ( .A1(n11430), .A2(n11428), .ZN(n17497) );
  NAND2_X1 U12647 ( .A1(n18928), .A2(n11438), .ZN(n11434) );
  OAI211_X1 U12648 ( .C1(n18928), .C2(n13819), .A(n11434), .B(n11433), .ZN(
        n11436) );
  NAND2_X1 U12649 ( .A1(n18928), .A2(n11441), .ZN(n11440) );
  AOI21_X1 U12650 ( .B1(n18928), .B2(n13817), .A(n13821), .ZN(n11435) );
  NOR2_X1 U12651 ( .A1(n11441), .A2(n11442), .ZN(n11438) );
  NAND2_X1 U12652 ( .A1(n18928), .A2(n13817), .ZN(n13820) );
  INV_X1 U12653 ( .A(n13817), .ZN(n11442) );
  AND3_X2 U12654 ( .A1(n11445), .A2(n13841), .A3(n11515), .ZN(n13842) );
  NAND4_X1 U12655 ( .A1(n11450), .A2(n11448), .A3(n13769), .A4(n13768), .ZN(
        n21396) );
  NAND3_X1 U12656 ( .A1(n13830), .A2(n21688), .A3(n21697), .ZN(n11453) );
  OAI21_X1 U12657 ( .B1(n12564), .B2(n11461), .A(n11460), .ZN(n16697) );
  NAND3_X1 U12658 ( .A1(n11463), .A2(n11464), .A3(n11213), .ZN(n11462) );
  NAND4_X1 U12659 ( .A1(n11467), .A2(n11552), .A3(n11550), .A4(n11551), .ZN(
        n11466) );
  AND2_X1 U12660 ( .A1(n11549), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11467) );
  NAND4_X1 U12661 ( .A1(n11215), .A2(n11546), .A3(n11548), .A4(n11469), .ZN(
        n11468) );
  NAND2_X1 U12662 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11469) );
  NAND2_X1 U12663 ( .A1(n11471), .A2(n11677), .ZN(n11654) );
  OAI21_X2 U12664 ( .B1(n17519), .B2(n11473), .A(n11472), .ZN(n17499) );
  INV_X1 U12665 ( .A(n17520), .ZN(n11474) );
  NAND3_X1 U12666 ( .A1(n12389), .A2(n12679), .A3(n12685), .ZN(n12392) );
  NAND3_X1 U12667 ( .A1(n12393), .A2(n12394), .A3(n12354), .ZN(n12385) );
  NAND2_X1 U12668 ( .A1(n11476), .A2(n12885), .ZN(n12962) );
  AND2_X1 U12669 ( .A1(n11476), .A2(n14183), .ZN(n16722) );
  AND2_X2 U12670 ( .A1(n12883), .A2(n12884), .ZN(n11476) );
  AND2_X2 U12671 ( .A1(n12815), .A2(n11477), .ZN(n12876) );
  AND2_X2 U12672 ( .A1(n12818), .A2(n11477), .ZN(n12830) );
  NAND2_X1 U12673 ( .A1(n14437), .A2(n11477), .ZN(n14445) );
  NAND2_X1 U12674 ( .A1(n17061), .A2(n11479), .ZN(n11478) );
  NAND2_X1 U12675 ( .A1(n11480), .A2(n11478), .ZN(n16976) );
  NAND2_X1 U12676 ( .A1(n17061), .A2(n16345), .ZN(n17008) );
  INV_X1 U12677 ( .A(n16345), .ZN(n11484) );
  NAND2_X1 U12678 ( .A1(n20742), .A2(n20741), .ZN(n20740) );
  AOI21_X1 U12679 ( .B1(n20747), .B2(n11488), .A(n11220), .ZN(n11485) );
  NAND2_X1 U12680 ( .A1(n20742), .A2(n11487), .ZN(n11486) );
  AND2_X1 U12681 ( .A1(n20747), .A2(n20741), .ZN(n11487) );
  NAND4_X1 U12682 ( .A1(n11582), .A2(n11581), .A3(n11580), .A4(n11583), .ZN(
        n11493) );
  NAND4_X1 U12683 ( .A1(n11586), .A2(n11585), .A3(n11584), .A4(n11587), .ZN(
        n11495) );
  OAI21_X1 U12684 ( .B1(n16694), .B2(n20165), .A(n11497), .ZN(P2_U2889) );
  INV_X1 U12685 ( .A(n15312), .ZN(n13145) );
  OAI21_X1 U12686 ( .B1(n16686), .B2(n19310), .A(n12228), .ZN(n12229) );
  AOI21_X1 U12687 ( .B1(n11527), .B2(n18095), .A(n16707), .ZN(n16708) );
  AOI21_X1 U12688 ( .B1(n11527), .B2(n19420), .A(n17657), .ZN(n17658) );
  AND2_X2 U12689 ( .A1(n12819), .A2(n12818), .ZN(n12989) );
  AOI22_X1 U12690 ( .A1(n12357), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n19990), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12304) );
  NAND2_X1 U12691 ( .A1(n14639), .A2(n14638), .ZN(n14692) );
  INV_X1 U12692 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11543) );
  NAND2_X1 U12693 ( .A1(n16660), .A2(n16659), .ZN(n16661) );
  NAND2_X1 U12694 ( .A1(n15469), .A2(n16076), .ZN(n12662) );
  NAND2_X1 U12695 ( .A1(n13146), .A2(n13147), .ZN(n13023) );
  INV_X1 U12696 ( .A(n13146), .ZN(n13148) );
  AND2_X4 U12697 ( .A1(n12817), .A2(n12816), .ZN(n13441) );
  AOI22_X1 U12698 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11187), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11618) );
  OR2_X1 U12699 ( .A1(n13718), .A2(n14172), .ZN(n11514) );
  NOR2_X1 U12700 ( .A1(n13718), .A2(n13719), .ZN(n13845) );
  OR2_X1 U12701 ( .A1(n18755), .A2(n18718), .ZN(n11515) );
  NAND2_X1 U12702 ( .A1(n20727), .A2(n16150), .ZN(n16841) );
  AND2_X1 U12703 ( .A1(n17256), .A2(n17099), .ZN(n11516) );
  AND4_X1 U12704 ( .A1(n13752), .A2(n13751), .A3(n13750), .A4(n13749), .ZN(
        n11517) );
  NOR2_X1 U12705 ( .A1(n14672), .A2(n14626), .ZN(n11518) );
  AND2_X1 U12706 ( .A1(n11627), .A2(n12603), .ZN(n11519) );
  AND2_X1 U12707 ( .A1(n16903), .A2(n16902), .ZN(n11520) );
  NAND2_X1 U12708 ( .A1(n18776), .A2(n18734), .ZN(n18963) );
  INV_X1 U12709 ( .A(n14394), .ZN(n14522) );
  AND4_X1 U12710 ( .A1(n11948), .A2(n11947), .A3(n11946), .A4(n11945), .ZN(
        n11521) );
  AND4_X1 U12711 ( .A1(n11963), .A2(n11962), .A3(n11961), .A4(n11960), .ZN(
        n11523) );
  AND2_X1 U12712 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11524) );
  AND2_X1 U12713 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11525) );
  OR2_X1 U12714 ( .A1(n19225), .A2(n12507), .ZN(n12753) );
  AND4_X1 U12715 ( .A1(n12438), .A2(n12437), .A3(n12436), .A4(n12435), .ZN(
        n11526) );
  INV_X1 U12716 ( .A(n11873), .ZN(n12023) );
  INV_X1 U12717 ( .A(n19432), .ZN(n19316) );
  AND2_X1 U12718 ( .A1(n12643), .A2(n15153), .ZN(n19419) );
  INV_X1 U12719 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12231) );
  INV_X1 U12720 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12232) );
  NOR2_X1 U12721 ( .A1(n21559), .A2(n14151), .ZN(n13746) );
  NAND2_X1 U12722 ( .A1(n12303), .A2(n12316), .ZN(n12421) );
  AND2_X1 U12723 ( .A1(n16703), .A2(n16702), .ZN(n11527) );
  AND2_X1 U12724 ( .A1(n17492), .A2(n12695), .ZN(n11528) );
  INV_X1 U12725 ( .A(n15370), .ZN(n15369) );
  OR2_X1 U12726 ( .A1(n12068), .A2(n12067), .ZN(n15370) );
  OR2_X1 U12727 ( .A1(n19686), .A2(n19526), .ZN(n19813) );
  INV_X1 U12728 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19952) );
  INV_X1 U12729 ( .A(n11720), .ZN(n11745) );
  AND2_X1 U12730 ( .A1(n16054), .A2(n14366), .ZN(n15997) );
  AND2_X1 U12731 ( .A1(n13471), .A2(n13470), .ZN(n11529) );
  NOR2_X1 U12732 ( .A1(n15454), .A2(n15351), .ZN(n11530) );
  OR2_X1 U12733 ( .A1(n18027), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19380) );
  AND2_X1 U12734 ( .A1(n11913), .A2(n11874), .ZN(n11532) );
  INV_X1 U12735 ( .A(n11919), .ZN(n12120) );
  INV_X1 U12736 ( .A(n11918), .ZN(n12022) );
  NAND2_X1 U12737 ( .A1(n16071), .A2(n11997), .ZN(n14618) );
  AND2_X1 U12738 ( .A1(n16574), .A2(n16597), .ZN(n11533) );
  OR2_X1 U12739 ( .A1(n16556), .A2(n17398), .ZN(n11534) );
  AND2_X1 U12740 ( .A1(n12793), .A2(n16695), .ZN(n11535) );
  AND2_X1 U12741 ( .A1(n16031), .A2(n11658), .ZN(n11537) );
  NAND2_X1 U12742 ( .A1(n11651), .A2(n11658), .ZN(n11676) );
  AND4_X1 U12743 ( .A1(n12874), .A2(n12873), .A3(n12872), .A4(n12871), .ZN(
        n11538) );
  AND4_X1 U12744 ( .A1(n12868), .A2(n12867), .A3(n12866), .A4(n12865), .ZN(
        n11539) );
  AND3_X1 U12745 ( .A1(n14445), .A2(n14444), .A3(n14443), .ZN(n11542) );
  OR2_X1 U12746 ( .A1(n22406), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13633) );
  AND2_X1 U12747 ( .A1(n11359), .A2(n13615), .ZN(n13641) );
  OR2_X1 U12748 ( .A1(n13644), .A2(n13643), .ZN(n13646) );
  INV_X1 U12749 ( .A(n13184), .ZN(n13081) );
  NAND2_X1 U12750 ( .A1(n12317), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12318) );
  OR2_X1 U12751 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n15215), .ZN(
        n13653) );
  INV_X1 U12752 ( .A(n13203), .ZN(n13107) );
  AOI22_X1 U12753 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12840) );
  NAND2_X1 U12754 ( .A1(n12941), .A2(n14882), .ZN(n12870) );
  AND3_X1 U12755 ( .A1(n12956), .A2(n14428), .A3(n15070), .ZN(n12937) );
  AOI22_X1 U12756 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11187), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11623) );
  AOI22_X1 U12757 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11854), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11616) );
  AND2_X1 U12758 ( .A1(n16597), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14712) );
  AND4_X1 U12759 ( .A1(n11991), .A2(n11990), .A3(n11989), .A4(n11988), .ZN(
        n11994) );
  AOI22_X1 U12760 ( .A1(n11856), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11854), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U12761 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11186), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11643) );
  AOI22_X1 U12762 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20036), .B1(
        n19923), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12329) );
  AND2_X1 U12763 ( .A1(n14002), .A2(n14003), .ZN(n13987) );
  INV_X1 U12764 ( .A(n16828), .ZN(n13388) );
  INV_X1 U12765 ( .A(n16889), .ZN(n13339) );
  INV_X1 U12766 ( .A(n15620), .ZN(n13230) );
  INV_X1 U12767 ( .A(n12886), .ZN(n14284) );
  AND2_X1 U12768 ( .A1(n14291), .A2(n12936), .ZN(n14305) );
  NOR2_X1 U12769 ( .A1(n20174), .A2(n12198), .ZN(n12453) );
  OAI21_X1 U12770 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n14038), .ZN(n12563) );
  NAND2_X1 U12771 ( .A1(n11475), .A2(n16075), .ZN(n12665) );
  AOI22_X1 U12772 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11187), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11562) );
  INV_X1 U12773 ( .A(n13986), .ZN(n14003) );
  NAND2_X1 U12774 ( .A1(n13669), .A2(n13668), .ZN(n13683) );
  INV_X1 U12775 ( .A(n16144), .ZN(n13325) );
  OR2_X1 U12776 ( .A1(n16954), .A2(n13557), .ZN(n13495) );
  OR2_X1 U12777 ( .A1(n22258), .A2(n13557), .ZN(n13409) );
  OR2_X1 U12778 ( .A1(n17250), .A2(n16350), .ZN(n16354) );
  INV_X1 U12779 ( .A(n20722), .ZN(n15331) );
  AND2_X1 U12780 ( .A1(n14370), .A2(n11166), .ZN(n11680) );
  INV_X1 U12781 ( .A(n11939), .ZN(n16458) );
  INV_X1 U12782 ( .A(n12024), .ZN(n16452) );
  NAND2_X1 U12783 ( .A1(n11996), .A2(n12442), .ZN(n11997) );
  NAND2_X1 U12784 ( .A1(n12744), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11703) );
  AND2_X1 U12785 ( .A1(n17650), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17651) );
  NAND2_X1 U12786 ( .A1(n11875), .A2(n11532), .ZN(n14381) );
  NOR2_X1 U12787 ( .A1(n13717), .A2(n13716), .ZN(n13800) );
  NOR2_X1 U12788 ( .A1(n19027), .A2(n21337), .ZN(n13934) );
  INV_X1 U12789 ( .A(n19645), .ZN(n13977) );
  NOR2_X1 U12790 ( .A1(n21381), .A2(n13818), .ZN(n13791) );
  INV_X1 U12791 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13796) );
  NAND2_X1 U12792 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21535), .ZN(
        n14144) );
  AND4_X1 U12793 ( .A1(n12905), .A2(n12904), .A3(n12903), .A4(n12902), .ZN(
        n12906) );
  OR2_X1 U12794 ( .A1(n16936), .A2(n13557), .ZN(n13534) );
  NAND2_X1 U12795 ( .A1(n16899), .A2(n11541), .ZN(n16903) );
  AOI211_X1 U12796 ( .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n22424), .A(n17985), 
        .B(n22296), .ZN(n14757) );
  INV_X1 U12797 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22406) );
  NAND2_X1 U12798 ( .A1(n12225), .A2(n12224), .ZN(n12226) );
  OAI211_X1 U12799 ( .C1(n16598), .C2(n16599), .A(n17374), .B(n16597), .ZN(
        n16620) );
  NAND2_X1 U12800 ( .A1(n12240), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12237) );
  INV_X1 U12801 ( .A(n15447), .ZN(n15489) );
  AND2_X1 U12802 ( .A1(n12567), .A2(n17691), .ZN(n17507) );
  NOR2_X1 U12803 ( .A1(n17592), .A2(n12752), .ZN(n17582) );
  AND3_X1 U12804 ( .A1(n17874), .A2(n18063), .A3(n17873), .ZN(n17890) );
  NAND2_X1 U12805 ( .A1(n11669), .A2(n19080), .ZN(n11846) );
  NAND2_X1 U12806 ( .A1(n11606), .A2(n11571), .ZN(n11613) );
  NOR2_X2 U12808 ( .A1(n20943), .A2(n18916), .ZN(n18902) );
  INV_X1 U12809 ( .A(n21925), .ZN(n21731) );
  XNOR2_X1 U12810 ( .A(n13797), .B(n13796), .ZN(n18954) );
  INV_X1 U12811 ( .A(n12947), .ZN(n12949) );
  AOI21_X1 U12812 ( .B1(n16391), .B2(n22210), .A(n16390), .ZN(n16392) );
  NOR2_X1 U12813 ( .A1(n16776), .A2(n16952), .ZN(n16774) );
  NOR2_X1 U12814 ( .A1(n13389), .A2(n16993), .ZN(n13390) );
  NOR2_X1 U12815 ( .A1(n13222), .A2(n15457), .ZN(n13226) );
  OR2_X1 U12816 ( .A1(n13140), .A2(n15361), .ZN(n13222) );
  INV_X1 U12817 ( .A(n22264), .ZN(n22213) );
  AND3_X1 U12818 ( .A1(n13144), .A2(n13143), .A3(n13142), .ZN(n15351) );
  NAND2_X1 U12819 ( .A1(n13514), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13551) );
  AND2_X1 U12820 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n13322), .ZN(
        n13326) );
  AOI21_X1 U12821 ( .B1(n15585), .B2(n13299), .A(n13208), .ZN(n15281) );
  INV_X1 U12822 ( .A(n16324), .ZN(n16325) );
  NOR2_X2 U12823 ( .A1(n17322), .A2(n15552), .ZN(n16005) );
  AND2_X1 U12824 ( .A1(n15301), .A2(n15303), .ZN(n22053) );
  INV_X1 U12825 ( .A(n22401), .ZN(n22423) );
  OR2_X1 U12826 ( .A1(n14874), .A2(n14873), .ZN(n22728) );
  INV_X1 U12827 ( .A(n14939), .ZN(n15033) );
  AOI21_X1 U12828 ( .B1(n22457), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n22678), 
        .ZN(n15035) );
  OR2_X1 U12829 ( .A1(n11196), .A2(n14826), .ZN(n15002) );
  OR2_X1 U12830 ( .A1(n14841), .A2(n15415), .ZN(n22684) );
  INV_X1 U12831 ( .A(n12562), .ZN(n12560) );
  INV_X1 U12832 ( .A(n17420), .ZN(n14580) );
  NAND2_X1 U12833 ( .A1(n20429), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12597) );
  NOR2_X1 U12834 ( .A1(n17654), .A2(n17653), .ZN(n17655) );
  OR2_X1 U12835 ( .A1(n17825), .A2(n17602), .ZN(n17828) );
  AOI21_X1 U12836 ( .B1(n19105), .B2(n14704), .A(n14603), .ZN(n14611) );
  NAND2_X1 U12837 ( .A1(n12599), .A2(n12598), .ZN(n16020) );
  NAND2_X1 U12838 ( .A1(n20058), .A2(n16017), .ZN(n20074) );
  INV_X1 U12839 ( .A(n20028), .ZN(n20030) );
  NAND2_X1 U12840 ( .A1(n16022), .A2(n16021), .ZN(n20086) );
  INV_X1 U12841 ( .A(n20424), .ZN(n20432) );
  NOR3_X1 U12842 ( .A1(n13976), .A2(n14006), .A3(n14142), .ZN(n14489) );
  NOR2_X1 U12843 ( .A1(n21312), .A2(n21166), .ZN(n21167) );
  NOR2_X1 U12844 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n21044), .ZN(n21051) );
  NOR2_X1 U12845 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n20982), .ZN(n21004) );
  INV_X1 U12846 ( .A(n19605), .ZN(n21404) );
  INV_X1 U12847 ( .A(n21512), .ZN(n21461) );
  INV_X1 U12848 ( .A(n14129), .ZN(n17951) );
  CLKBUF_X1 U12849 ( .A(n11522), .Z(n18765) );
  NOR2_X1 U12850 ( .A1(n21720), .A2(n14025), .ZN(n21567) );
  AND2_X1 U12851 ( .A1(n21074), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18577) );
  INV_X1 U12852 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18916) );
  INV_X1 U12853 ( .A(n21964), .ZN(n14116) );
  NOR2_X2 U12854 ( .A1(n11145), .A2(n13825), .ZN(n18755) );
  NAND2_X1 U12855 ( .A1(n18845), .A2(n18824), .ZN(n18668) );
  NOR2_X1 U12856 ( .A1(n14122), .A2(n21656), .ZN(n21928) );
  INV_X1 U12857 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19524) );
  NOR2_X1 U12858 ( .A1(n13884), .A2(n13883), .ZN(n19605) );
  OAI21_X1 U12859 ( .B1(n17109), .B2(n22276), .A(n16392), .ZN(n16393) );
  AND2_X1 U12860 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n22273), .ZN(n16797) );
  NAND2_X1 U12861 ( .A1(n13390), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13424) );
  NAND2_X1 U12862 ( .A1(n13227), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13286) );
  XNOR2_X1 U12863 ( .A(n15065), .B(n16327), .ZN(n16378) );
  AND2_X1 U12864 ( .A1(n11192), .A2(n15072), .ZN(n22217) );
  INV_X1 U12865 ( .A(n22262), .ZN(n22236) );
  INV_X1 U12866 ( .A(n20698), .ZN(n20725) );
  INV_X1 U12867 ( .A(n16841), .ZN(n20724) );
  INV_X1 U12868 ( .A(n14328), .ZN(n22381) );
  AND2_X1 U12870 ( .A1(n16002), .A2(n15624), .ZN(n22168) );
  AND2_X1 U12871 ( .A1(n15352), .A2(n15313), .ZN(n22152) );
  NAND2_X1 U12872 ( .A1(n13188), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13196) );
  INV_X1 U12873 ( .A(n20759), .ZN(n20761) );
  INV_X1 U12874 ( .A(n22302), .ZN(n22807) );
  AND2_X1 U12875 ( .A1(n16983), .A2(n16982), .ZN(n16998) );
  AND2_X1 U12876 ( .A1(n17315), .A2(n17236), .ZN(n21976) );
  AND2_X1 U12877 ( .A1(n14295), .A2(n22807), .ZN(n14318) );
  INV_X1 U12878 ( .A(n22058), .ZN(n22075) );
  INV_X1 U12879 ( .A(n21999), .ZN(n22056) );
  AND2_X1 U12880 ( .A1(n14318), .A2(n14296), .ZN(n22043) );
  NOR2_X2 U12881 ( .A1(n22423), .A2(n15037), .ZN(n22697) );
  INV_X1 U12882 ( .A(n22701), .ZN(n22703) );
  AND2_X1 U12883 ( .A1(n22401), .A2(n22400), .ZN(n22709) );
  NOR2_X2 U12884 ( .A1(n22423), .A2(n15415), .ZN(n22717) );
  NOR2_X2 U12885 ( .A1(n14874), .A2(n15002), .ZN(n22730) );
  INV_X1 U12886 ( .A(n22728), .ZN(n22738) );
  INV_X1 U12887 ( .A(n22742), .ZN(n22746) );
  AND2_X1 U12888 ( .A1(n15020), .A2(n15034), .ZN(n22758) );
  AND2_X1 U12889 ( .A1(n11196), .A2(n14826), .ZN(n22400) );
  AND2_X1 U12890 ( .A1(n15020), .A2(n15019), .ZN(n22772) );
  OR2_X1 U12891 ( .A1(n11196), .A2(n22280), .ZN(n15037) );
  INV_X1 U12892 ( .A(n22513), .ZN(n22523) );
  INV_X1 U12893 ( .A(n22640), .ZN(n22649) );
  INV_X1 U12894 ( .A(n22684), .ZN(n22797) );
  INV_X1 U12895 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n22287) );
  INV_X1 U12896 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n22329) );
  NAND2_X1 U12897 ( .A1(n12278), .A2(n12277), .ZN(n12280) );
  NOR2_X1 U12898 ( .A1(n11181), .A2(n17357), .ZN(n14100) );
  OR2_X1 U12899 ( .A1(n19074), .A2(n12223), .ZN(n19338) );
  INV_X1 U12900 ( .A(n19342), .ZN(n19323) );
  INV_X1 U12901 ( .A(n19338), .ZN(n19307) );
  OR2_X1 U12902 ( .A1(n12102), .A2(n12101), .ZN(n15536) );
  INV_X1 U12903 ( .A(n14580), .ZN(n17423) );
  INV_X1 U12904 ( .A(n14618), .ZN(n14620) );
  INV_X1 U12905 ( .A(n20165), .ZN(n20322) );
  INV_X2 U12906 ( .A(n12188), .ZN(n19079) );
  INV_X1 U12907 ( .A(n18076), .ZN(n18102) );
  AND2_X1 U12908 ( .A1(n19411), .A2(n12723), .ZN(n17896) );
  NAND2_X1 U12909 ( .A1(n12640), .A2(n19078), .ZN(n12746) );
  OAI21_X1 U12910 ( .B1(n16028), .B2(n16027), .A(n16026), .ZN(n20543) );
  INV_X1 U12911 ( .A(n20536), .ZN(n20545) );
  AND2_X1 U12912 ( .A1(n20097), .A2(n20081), .ZN(n20532) );
  INV_X1 U12913 ( .A(n20515), .ZN(n20362) );
  OAI21_X1 U12914 ( .B1(n20054), .B2(n20053), .A(n20052), .ZN(n20509) );
  INV_X1 U12915 ( .A(n20507), .ZN(n20359) );
  NOR2_X1 U12916 ( .A1(n20030), .A2(n20073), .ZN(n20495) );
  OAI21_X1 U12917 ( .B1(n20347), .B2(n20001), .A(n20086), .ZN(n20483) );
  AND2_X1 U12918 ( .A1(n20058), .A2(n18127), .ZN(n20028) );
  NOR2_X1 U12919 ( .A1(n19944), .A2(n20081), .ZN(n20027) );
  INV_X1 U12920 ( .A(n20086), .ZN(n20426) );
  AND2_X1 U12921 ( .A1(n19982), .A2(n19964), .ZN(n20466) );
  NOR2_X1 U12922 ( .A1(n20058), .A2(n18127), .ZN(n19982) );
  AND2_X1 U12923 ( .A1(n19941), .A2(n20027), .ZN(n20455) );
  AOI21_X1 U12924 ( .B1(n20236), .B2(n20086), .A(n19934), .ZN(n20442) );
  AND2_X1 U12925 ( .A1(n19079), .A2(n20428), .ZN(n20418) );
  INV_X1 U12926 ( .A(n20540), .ZN(n20274) );
  AND3_X1 U12927 ( .A1(n15111), .A2(n15110), .A3(n15109), .ZN(n16063) );
  NAND2_X1 U12928 ( .A1(n17953), .A2(n20842), .ZN(n20899) );
  NAND2_X1 U12929 ( .A1(n21337), .A2(n21899), .ZN(n21847) );
  AND2_X1 U12930 ( .A1(n21179), .A2(n21178), .ZN(n21207) );
  NOR2_X1 U12931 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n21063), .ZN(n21088) );
  NOR2_X1 U12932 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n21019), .ZN(n21034) );
  NOR2_X1 U12933 ( .A1(n20899), .A2(n21336), .ZN(n20905) );
  INV_X1 U12934 ( .A(n21318), .ZN(n21301) );
  NOR3_X1 U12935 ( .A1(n21493), .A2(n21442), .A3(n21441), .ZN(n21487) );
  NAND2_X1 U12936 ( .A1(n21503), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n21493) );
  NAND2_X1 U12937 ( .A1(n21443), .A2(n21529), .ZN(n21512) );
  INV_X1 U12938 ( .A(n21461), .ZN(n21519) );
  INV_X1 U12939 ( .A(n21336), .ZN(n19027) );
  NOR2_X1 U12940 ( .A1(n20891), .A2(n20849), .ZN(n20860) );
  NOR2_X1 U12941 ( .A1(n20843), .A2(n21339), .ZN(n20878) );
  INV_X1 U12942 ( .A(n20893), .ZN(n20849) );
  NOR2_X1 U12943 ( .A1(n21961), .A2(n17951), .ZN(n20842) );
  INV_X1 U12944 ( .A(n18734), .ZN(n18808) );
  NOR3_X1 U12945 ( .A1(n18643), .A2(n21718), .A3(n21721), .ZN(n18826) );
  INV_X1 U12946 ( .A(n18839), .ZN(n18883) );
  NAND2_X1 U12947 ( .A1(n14147), .A2(n13938), .ZN(n21883) );
  INV_X1 U12948 ( .A(n21911), .ZN(n21875) );
  NOR2_X1 U12949 ( .A1(n11153), .A2(n21897), .ZN(n21835) );
  INV_X1 U12950 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n21537) );
  NOR2_X1 U12951 ( .A1(n21955), .A2(n14177), .ZN(n21944) );
  INV_X1 U12952 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n22361) );
  INV_X1 U12953 ( .A(n14191), .ZN(n22811) );
  INV_X1 U12954 ( .A(n22805), .ZN(n22803) );
  INV_X1 U12955 ( .A(n16393), .ZN(n16394) );
  OR2_X1 U12956 ( .A1(n16378), .A2(n15068), .ZN(n22269) );
  INV_X1 U12957 ( .A(n22217), .ZN(n22276) );
  NOR2_X1 U12958 ( .A1(n13707), .A2(n13706), .ZN(n13708) );
  OAI21_X1 U12959 ( .B1(n11529), .B2(n16780), .A(n11198), .ZN(n16963) );
  OR2_X1 U12960 ( .A1(n16890), .A2(n14366), .ZN(n16056) );
  INV_X1 U12961 ( .A(n20604), .ZN(n20635) );
  OR2_X1 U12962 ( .A1(n14191), .A2(n13690), .ZN(n14212) );
  INV_X1 U12963 ( .A(n22168), .ZN(n17059) );
  NAND2_X1 U12964 ( .A1(n20728), .A2(n14633), .ZN(n20759) );
  NAND2_X1 U12965 ( .A1(n14318), .A2(n14317), .ZN(n22058) );
  INV_X1 U12966 ( .A(n22030), .ZN(n22051) );
  INV_X1 U12967 ( .A(n22043), .ZN(n22082) );
  AOI22_X1 U12968 ( .A1(n22390), .A2(n22396), .B1(n22393), .B2(n22453), .ZN(
        n22693) );
  NAND2_X1 U12969 ( .A1(n22401), .A2(n15034), .ZN(n22701) );
  AOI22_X1 U12970 ( .A1(n22405), .A2(n22411), .B1(n22453), .B2(n22439), .ZN(
        n22707) );
  INV_X1 U12971 ( .A(n22425), .ZN(n22713) );
  OR2_X1 U12972 ( .A1(n15037), .A2(n14874), .ZN(n22726) );
  AOI22_X1 U12973 ( .A1(n22444), .A2(n22440), .B1(n22474), .B2(n22439), .ZN(
        n22734) );
  INV_X1 U12974 ( .A(n22739), .ZN(n14930) );
  NAND2_X1 U12975 ( .A1(n15020), .A2(n15000), .ZN(n22755) );
  AOI22_X1 U12976 ( .A1(n22455), .A2(n22463), .B1(n22454), .B2(n22453), .ZN(
        n22762) );
  NAND2_X1 U12977 ( .A1(n15020), .A2(n22400), .ZN(n22768) );
  INV_X1 U12978 ( .A(n15231), .ZN(n22583) );
  INV_X1 U12979 ( .A(n15248), .ZN(n22677) );
  OR2_X1 U12980 ( .A1(n15037), .A2(n14841), .ZN(n22783) );
  OR2_X1 U12981 ( .A1(n14841), .A2(n14873), .ZN(n22801) );
  AND2_X1 U12982 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n18017), .ZN(n22293) );
  OR2_X1 U12983 ( .A1(n15158), .A2(n12217), .ZN(n14198) );
  OR3_X1 U12984 ( .A1(n12215), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n22338), 
        .ZN(n19310) );
  OR3_X1 U12985 ( .A1(n12215), .A2(n12219), .A3(n12214), .ZN(n19342) );
  NAND2_X1 U12986 ( .A1(n14579), .A2(n19078), .ZN(n17420) );
  NAND2_X1 U12987 ( .A1(n14734), .A2(n14733), .ZN(n20058) );
  INV_X1 U12988 ( .A(n20319), .ZN(n17475) );
  NOR2_X1 U12989 ( .A1(n20322), .A2(n20321), .ZN(n20171) );
  OR2_X1 U12990 ( .A1(n20319), .A2(n11163), .ZN(n20165) );
  INV_X1 U12991 ( .A(n18147), .ZN(n18182) );
  OR2_X1 U12992 ( .A1(n19451), .A2(n19079), .ZN(n18103) );
  OR2_X1 U12993 ( .A1(n14060), .A2(n19375), .ZN(n14061) );
  INV_X1 U12994 ( .A(n19419), .ZN(n19388) );
  OR2_X1 U12995 ( .A1(n12746), .A2(n12696), .ZN(n19375) );
  AOI21_X1 U12996 ( .B1(n16025), .B2(n20538), .A(n20426), .ZN(n20548) );
  NAND2_X1 U12997 ( .A1(n20097), .A2(n19929), .ZN(n20536) );
  INV_X1 U12998 ( .A(n20532), .ZN(n20528) );
  INV_X1 U12999 ( .A(n20524), .ZN(n20521) );
  NAND2_X1 U13000 ( .A1(n20043), .A2(n20042), .ZN(n20515) );
  NAND2_X1 U13001 ( .A1(n20028), .A2(n20027), .ZN(n20507) );
  INV_X1 U13002 ( .A(n20404), .ZN(n20505) );
  INV_X1 U13003 ( .A(n20495), .ZN(n20402) );
  NAND2_X1 U13004 ( .A1(n20042), .A2(n20028), .ZN(n20492) );
  NAND2_X1 U13005 ( .A1(n19982), .A2(n20015), .ZN(n20478) );
  AOI211_X2 U13006 ( .C1(n19974), .C2(n19977), .A(n20426), .B(n19973), .ZN(
        n20471) );
  NAND2_X1 U13007 ( .A1(n20042), .A2(n19982), .ZN(n20464) );
  INV_X1 U13008 ( .A(n20368), .ZN(n20373) );
  INV_X1 U13009 ( .A(n20488), .ZN(n20539) );
  INV_X1 U13010 ( .A(n20147), .ZN(n20157) );
  INV_X1 U13011 ( .A(n20269), .ZN(n20266) );
  INV_X1 U13012 ( .A(n19078), .ZN(n19448) );
  AOI211_X1 U13013 ( .C1(n21331), .C2(P3_EBX_REG_31__SCAN_IN), .A(n21321), .B(
        n21320), .ZN(n21325) );
  NAND2_X1 U13014 ( .A1(n21329), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21318) );
  INV_X1 U13015 ( .A(n21135), .ZN(n21311) );
  AND2_X1 U13016 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n21363), .ZN(n21366) );
  NOR2_X1 U13017 ( .A1(n13735), .A2(n13734), .ZN(n21381) );
  INV_X1 U13018 ( .A(n21526), .ZN(n21522) );
  INV_X1 U13019 ( .A(n19028), .ZN(n19026) );
  INV_X1 U13020 ( .A(n20849), .ZN(n20889) );
  NAND3_X1 U13021 ( .A1(n18970), .A2(n22315), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n18734) );
  INV_X1 U13022 ( .A(n18869), .ZN(n18643) );
  INV_X1 U13023 ( .A(n18963), .ZN(n18955) );
  INV_X1 U13024 ( .A(n14124), .ZN(n18973) );
  NOR2_X1 U13025 ( .A1(n18729), .A2(n11212), .ZN(n14032) );
  INV_X1 U13026 ( .A(n21939), .ZN(n21868) );
  INV_X1 U13027 ( .A(n21835), .ZN(n21828) );
  INV_X1 U13028 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19523) );
  INV_X1 U13029 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17950) );
  INV_X1 U13030 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n21960) );
  INV_X1 U13031 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21949) );
  INV_X1 U13032 ( .A(n19062), .ZN(n19059) );
  NAND2_X1 U13033 ( .A1(n13709), .A2(n13708), .ZN(P1_U2873) );
  NAND2_X1 U13034 ( .A1(n14033), .A2(n14032), .ZN(P3_U2834) );
  OR4_X1 U13035 ( .A1(n21135), .A2(n21950), .A3(n17948), .A4(n14178), .ZN(
        P3_U2997) );
  AND2_X4 U13036 ( .A1(n11849), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11848) );
  AND2_X4 U13037 ( .A1(n11850), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11854) );
  AOI22_X1 U13038 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11854), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11546) );
  AND2_X4 U13039 ( .A1(n11850), .A2(n11830), .ZN(n11856) );
  NAND2_X1 U13040 ( .A1(n11186), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11544) );
  AOI22_X1 U13041 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11182), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11548) );
  NOR2_X4 U13042 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U13043 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11182), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U13044 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11186), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11550) );
  AOI22_X1 U13045 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11854), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11555) );
  AOI21_X1 U13046 ( .B1(n11187), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11554) );
  NAND2_X1 U13047 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11553) );
  AND3_X1 U13048 ( .A1(n11555), .A2(n11554), .A3(n11553), .ZN(n11558) );
  AOI22_X1 U13049 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U13050 ( .A1(n11639), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11556) );
  NAND3_X1 U13051 ( .A1(n11558), .A2(n11557), .A3(n11556), .ZN(n11566) );
  NOR2_X1 U13052 ( .A1(n11525), .A2(n11560), .ZN(n11564) );
  AOI22_X1 U13053 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11854), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11561) );
  NAND4_X1 U13054 ( .A1(n11564), .A2(n11563), .A3(n11562), .A4(n11561), .ZN(
        n11565) );
  NAND2_X1 U13055 ( .A1(n11649), .A2(n11601), .ZN(n11632) );
  AOI22_X1 U13056 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U13057 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11854), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U13058 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11187), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11568) );
  NAND4_X1 U13059 ( .A1(n11570), .A2(n11569), .A3(n11568), .A4(n11567), .ZN(
        n11572) );
  AOI22_X1 U13060 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11187), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11576) );
  AOI22_X1 U13061 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11854), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U13062 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11574) );
  NAND4_X1 U13063 ( .A1(n11576), .A2(n11575), .A3(n11574), .A4(n11573), .ZN(
        n11577) );
  NAND2_X1 U13064 ( .A1(n11577), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11578) );
  NAND2_X1 U13065 ( .A1(n11632), .A2(n11676), .ZN(n11600) );
  AOI22_X1 U13066 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11186), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U13067 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11854), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11581) );
  AOI22_X1 U13068 ( .A1(n11182), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11580) );
  AOI22_X1 U13069 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11187), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U13070 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11854), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11585) );
  AOI22_X1 U13071 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U13072 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11187), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11591) );
  AOI22_X1 U13073 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U13074 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11854), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11588) );
  NAND4_X1 U13075 ( .A1(n11591), .A2(n11590), .A3(n11589), .A4(n11588), .ZN(
        n11592) );
  AOI22_X1 U13076 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11187), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U13077 ( .A1(n11856), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11854), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11594) );
  NAND4_X1 U13078 ( .A1(n11596), .A2(n11595), .A3(n11594), .A4(n11593), .ZN(
        n11597) );
  NAND2_X1 U13079 ( .A1(n11652), .A2(n16031), .ZN(n11674) );
  NAND2_X1 U13080 ( .A1(n11600), .A2(n11674), .ZN(n11628) );
  AOI22_X1 U13081 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11186), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U13082 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11854), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11603) );
  AOI22_X1 U13083 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11602) );
  NAND4_X1 U13084 ( .A1(n11605), .A2(n11604), .A3(n11603), .A4(n11602), .ZN(
        n11606) );
  AOI22_X1 U13085 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11186), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U13086 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11608) );
  AOI22_X1 U13087 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11854), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11607) );
  NAND4_X1 U13088 ( .A1(n11610), .A2(n11609), .A3(n11608), .A4(n11607), .ZN(
        n11611) );
  NAND2_X1 U13089 ( .A1(n11611), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11612) );
  NAND2_X2 U13090 ( .A1(n11613), .A2(n11612), .ZN(n20330) );
  NAND4_X1 U13091 ( .A1(n20233), .A2(n20330), .A3(n11658), .A4(n11659), .ZN(
        n11614) );
  NOR2_X2 U13092 ( .A1(n11628), .A2(n11614), .ZN(n11669) );
  INV_X1 U13093 ( .A(n11669), .ZN(n11631) );
  AOI22_X1 U13094 ( .A1(n11182), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11615) );
  NAND2_X1 U13095 ( .A1(n11619), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11626) );
  AOI22_X1 U13096 ( .A1(n11182), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11621) );
  AOI22_X1 U13097 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11854), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11620) );
  NAND2_X1 U13098 ( .A1(n11624), .A2(n11571), .ZN(n11625) );
  NAND2_X1 U13099 ( .A1(n11649), .A2(n11659), .ZN(n11627) );
  INV_X1 U13100 ( .A(n11628), .ZN(n11629) );
  NAND2_X1 U13101 ( .A1(n11519), .A2(n11629), .ZN(n11630) );
  NAND3_X1 U13102 ( .A1(n11631), .A2(n19080), .A3(n11630), .ZN(n12707) );
  INV_X1 U13103 ( .A(n11632), .ZN(n11660) );
  NOR2_X1 U13104 ( .A1(n11658), .A2(n11659), .ZN(n11633) );
  AOI22_X1 U13105 ( .A1(n11182), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11848), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11637) );
  AOI22_X1 U13106 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11854), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U13107 ( .A1(n11187), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11634) );
  NAND4_X1 U13108 ( .A1(n11637), .A2(n11636), .A3(n11635), .A4(n11634), .ZN(
        n11638) );
  AOI22_X1 U13109 ( .A1(n11182), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11856), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11641) );
  AOI22_X1 U13110 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11854), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11640) );
  NAND4_X1 U13111 ( .A1(n11643), .A2(n11642), .A3(n11641), .A4(n11640), .ZN(
        n11644) );
  NAND2_X2 U13112 ( .A1(n11646), .A2(n11645), .ZN(n11872) );
  INV_X4 U13113 ( .A(n11872), .ZN(n12188) );
  AND2_X1 U13114 ( .A1(n11163), .A2(n12188), .ZN(n11647) );
  NAND2_X1 U13115 ( .A1(n11707), .A2(n19080), .ZN(n11648) );
  XNOR2_X1 U13116 ( .A(n11649), .B(n11659), .ZN(n12605) );
  INV_X1 U13117 ( .A(n12605), .ZN(n11650) );
  NAND2_X1 U13118 ( .A1(n11650), .A2(n20233), .ZN(n12609) );
  NAND2_X1 U13119 ( .A1(n11652), .A2(n11651), .ZN(n12604) );
  AND2_X1 U13120 ( .A1(n12604), .A2(n19921), .ZN(n11653) );
  NAND2_X1 U13121 ( .A1(n12609), .A2(n11653), .ZN(n12705) );
  NAND2_X1 U13122 ( .A1(n12705), .A2(n16031), .ZN(n11655) );
  NAND2_X1 U13123 ( .A1(n11655), .A2(n11654), .ZN(n11706) );
  NAND2_X1 U13124 ( .A1(n11706), .A2(n12581), .ZN(n11656) );
  NAND2_X1 U13125 ( .A1(n11708), .A2(n11656), .ZN(n11657) );
  NAND2_X1 U13126 ( .A1(n11657), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11667) );
  NAND3_X1 U13127 ( .A1(n11662), .A2(n11660), .A3(n11659), .ZN(n12642) );
  NAND3_X1 U13128 ( .A1(n12642), .A2(n12603), .A3(n19079), .ZN(n11665) );
  INV_X1 U13130 ( .A(n12601), .ZN(n11664) );
  NAND2_X1 U13131 ( .A1(n11665), .A2(n11664), .ZN(n12703) );
  NAND2_X1 U13132 ( .A1(n11698), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11673) );
  INV_X1 U13133 ( .A(n11699), .ZN(n11681) );
  INV_X1 U13134 ( .A(n12589), .ZN(n11668) );
  AND2_X1 U13135 ( .A1(n12192), .A2(n19921), .ZN(n11876) );
  NAND3_X1 U13136 ( .A1(n12710), .A2(n11876), .A3(n11649), .ZN(n11670) );
  NAND2_X1 U13137 ( .A1(n11670), .A2(n11846), .ZN(n11683) );
  INV_X1 U13138 ( .A(n11683), .ZN(n11671) );
  NAND2_X1 U13139 ( .A1(n11671), .A2(n12216), .ZN(n15115) );
  NOR2_X1 U13140 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11730) );
  AOI22_X1 U13141 ( .A1(n15115), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n11730), .ZN(n11672) );
  NAND2_X1 U13142 ( .A1(n11673), .A2(n11672), .ZN(n11695) );
  INV_X1 U13143 ( .A(n11695), .ZN(n11694) );
  INV_X1 U13144 ( .A(n11676), .ZN(n11675) );
  NAND2_X1 U13145 ( .A1(n11675), .A2(n12188), .ZN(n12717) );
  NAND2_X1 U13146 ( .A1(n16136), .A2(n12192), .ZN(n11678) );
  OAI22_X1 U13147 ( .A1(n12717), .A2(n11678), .B1(n11677), .B2(n11676), .ZN(
        n11679) );
  AND2_X2 U13148 ( .A1(n11680), .A2(n11679), .ZN(n15112) );
  NAND2_X1 U13149 ( .A1(n11719), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11692) );
  AND2_X1 U13150 ( .A1(n11872), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11685) );
  INV_X1 U13151 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n11689) );
  NOR2_X1 U13152 ( .A1(n11699), .A2(n12641), .ZN(n11686) );
  NAND2_X1 U13153 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11687) );
  OAI211_X1 U13154 ( .C1(n11733), .C2(n11689), .A(n11688), .B(n11687), .ZN(
        n11690) );
  INV_X1 U13155 ( .A(n11690), .ZN(n11691) );
  NAND2_X1 U13156 ( .A1(n11692), .A2(n11691), .ZN(n11696) );
  INV_X1 U13157 ( .A(n11696), .ZN(n11693) );
  NAND2_X2 U13158 ( .A1(n11694), .A2(n11693), .ZN(n11716) );
  NAND2_X1 U13159 ( .A1(n11696), .A2(n11695), .ZN(n11697) );
  NAND2_X1 U13160 ( .A1(n12581), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11700) );
  NOR2_X1 U13161 ( .A1(n11700), .A2(n11699), .ZN(n11701) );
  NAND2_X1 U13162 ( .A1(n11730), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11702) );
  AND2_X1 U13163 ( .A1(n11703), .A2(n11702), .ZN(n11704) );
  NAND2_X1 U13164 ( .A1(n11705), .A2(n11704), .ZN(n12294) );
  NAND2_X1 U13165 ( .A1(n11706), .A2(n11707), .ZN(n12715) );
  NAND2_X1 U13166 ( .A1(n11719), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11714) );
  INV_X1 U13167 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n16338) );
  OAI21_X1 U13168 ( .B1(n11733), .B2(n16338), .A(n11709), .ZN(n11712) );
  INV_X1 U13169 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n14582) );
  INV_X1 U13170 ( .A(n11730), .ZN(n19424) );
  NAND2_X1 U13171 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11710) );
  OAI211_X1 U13172 ( .C1(n11745), .C2(n14582), .A(n19424), .B(n11710), .ZN(
        n11711) );
  AOI21_X1 U13173 ( .B1(n19436), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11717) );
  NAND2_X1 U13174 ( .A1(n11719), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11725) );
  INV_X1 U13175 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n14569) );
  NAND2_X1 U13176 ( .A1(n11720), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n11722) );
  NAND2_X1 U13177 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11721) );
  OAI211_X1 U13178 ( .C1(n11733), .C2(n14569), .A(n11722), .B(n11721), .ZN(
        n11723) );
  INV_X1 U13179 ( .A(n11723), .ZN(n11724) );
  NAND2_X1 U13180 ( .A1(n11726), .A2(n11727), .ZN(n11728) );
  NAND2_X1 U13181 ( .A1(n11698), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11732) );
  NAND2_X1 U13182 ( .A1(n11730), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11731) );
  NAND2_X1 U13183 ( .A1(n11732), .A2(n11731), .ZN(n11740) );
  NAND2_X1 U13184 ( .A1(n11719), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11739) );
  BUF_X4 U13185 ( .A(n11733), .Z(n12741) );
  INV_X1 U13186 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n11736) );
  NAND2_X1 U13187 ( .A1(n11720), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n11735) );
  NAND2_X1 U13188 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11734) );
  OAI211_X1 U13189 ( .C1(n12741), .C2(n11736), .A(n11735), .B(n11734), .ZN(
        n11737) );
  INV_X1 U13190 ( .A(n11737), .ZN(n11738) );
  NAND2_X1 U13191 ( .A1(n11739), .A2(n11738), .ZN(n11741) );
  NAND2_X1 U13192 ( .A1(n11741), .A2(n11740), .ZN(n11742) );
  INV_X1 U13194 ( .A(n11743), .ZN(n11744) );
  INV_X1 U13195 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11748) );
  NAND2_X1 U13196 ( .A1(n12738), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11747) );
  INV_X2 U13197 ( .A(n11745), .ZN(n11791) );
  AOI22_X1 U13198 ( .A1(n11791), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11746) );
  OAI211_X1 U13199 ( .C1(n12741), .C2(n11748), .A(n11747), .B(n11746), .ZN(
        n14741) );
  NAND2_X1 U13200 ( .A1(n14742), .A2(n14741), .ZN(n14722) );
  INV_X1 U13201 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n16079) );
  NAND2_X1 U13202 ( .A1(n11791), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11750) );
  NAND2_X1 U13203 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11749) );
  OAI211_X1 U13204 ( .C1(n12741), .C2(n16079), .A(n11750), .B(n11749), .ZN(
        n11751) );
  AOI21_X1 U13205 ( .B1(n12738), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n11751), .ZN(n14723) );
  INV_X1 U13206 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n11754) );
  NAND2_X1 U13207 ( .A1(n12738), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11753) );
  AOI22_X1 U13208 ( .A1(n11791), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11752) );
  OAI211_X1 U13209 ( .C1(n12741), .C2(n11754), .A(n11753), .B(n11752), .ZN(
        n14768) );
  NAND2_X1 U13210 ( .A1(n14724), .A2(n14768), .ZN(n14769) );
  INV_X1 U13211 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n11757) );
  NAND2_X1 U13212 ( .A1(n11791), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11756) );
  NAND2_X1 U13213 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11755) );
  OAI211_X1 U13214 ( .C1(n12741), .C2(n11757), .A(n11756), .B(n11755), .ZN(
        n11758) );
  AOI21_X1 U13215 ( .B1(n12738), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n11758), .ZN(n14863) );
  INV_X1 U13216 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n11761) );
  NAND2_X1 U13217 ( .A1(n12738), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11760) );
  AOI22_X1 U13218 ( .A1(n11791), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11759) );
  OAI211_X1 U13219 ( .C1(n12741), .C2(n11761), .A(n11760), .B(n11759), .ZN(
        n14987) );
  NAND2_X1 U13220 ( .A1(n14862), .A2(n14987), .ZN(n15194) );
  INV_X1 U13221 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n11763) );
  AOI22_X1 U13222 ( .A1(n11791), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11762) );
  OAI21_X1 U13223 ( .B1(n12741), .B2(n11763), .A(n11762), .ZN(n11764) );
  AOI21_X1 U13224 ( .B1(n12738), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n11764), .ZN(n15195) );
  NAND2_X1 U13225 ( .A1(n12738), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11770) );
  INV_X1 U13226 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n11767) );
  NAND2_X1 U13227 ( .A1(n11791), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11766) );
  NAND2_X1 U13228 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11765) );
  OAI211_X1 U13229 ( .C1(n12741), .C2(n11767), .A(n11766), .B(n11765), .ZN(
        n11768) );
  INV_X1 U13230 ( .A(n11768), .ZN(n11769) );
  NAND2_X1 U13231 ( .A1(n11770), .A2(n11769), .ZN(n15366) );
  INV_X1 U13232 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n17624) );
  NAND2_X1 U13233 ( .A1(n11791), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11772) );
  NAND2_X1 U13234 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11771) );
  OAI211_X1 U13235 ( .C1(n12741), .C2(n17624), .A(n11772), .B(n11771), .ZN(
        n11773) );
  AOI21_X1 U13236 ( .B1(n12738), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n11773), .ZN(n15490) );
  INV_X1 U13237 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n11776) );
  NAND2_X1 U13238 ( .A1(n11791), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11775) );
  NAND2_X1 U13239 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11774) );
  OAI211_X1 U13240 ( .C1(n12741), .C2(n11776), .A(n11775), .B(n11774), .ZN(
        n11777) );
  AOI21_X1 U13241 ( .B1(n12738), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n11777), .ZN(n15448) );
  INV_X1 U13242 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19187) );
  NAND2_X1 U13243 ( .A1(n11791), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11779) );
  NAND2_X1 U13244 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11778) );
  OAI211_X1 U13245 ( .C1(n12741), .C2(n19187), .A(n11779), .B(n11778), .ZN(
        n11780) );
  AOI21_X1 U13246 ( .B1(n12738), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n11780), .ZN(n15538) );
  INV_X1 U13247 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n11783) );
  NAND2_X1 U13248 ( .A1(n12738), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11782) );
  AOI22_X1 U13249 ( .A1(n11791), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11781) );
  OAI211_X1 U13250 ( .C1(n12741), .C2(n11783), .A(n11782), .B(n11781), .ZN(
        n15568) );
  INV_X1 U13251 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n18193) );
  NAND2_X1 U13252 ( .A1(n11791), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11785) );
  NAND2_X1 U13253 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11784) );
  OAI211_X1 U13254 ( .C1(n12741), .C2(n18193), .A(n11785), .B(n11784), .ZN(
        n11786) );
  AOI21_X1 U13255 ( .B1(n12738), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n11786), .ZN(n16045) );
  INV_X1 U13256 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n11789) );
  NAND2_X1 U13257 ( .A1(n11791), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11788) );
  NAND2_X1 U13258 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n11787) );
  OAI211_X1 U13259 ( .C1(n12741), .C2(n11789), .A(n11788), .B(n11787), .ZN(
        n11790) );
  AOI21_X1 U13260 ( .B1(n12738), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11790), .ZN(n16186) );
  INV_X1 U13261 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n17585) );
  NAND2_X1 U13262 ( .A1(n11791), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11793) );
  NAND2_X1 U13263 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11792) );
  OAI211_X1 U13264 ( .C1(n12741), .C2(n17585), .A(n11793), .B(n11792), .ZN(
        n11794) );
  AOI21_X1 U13265 ( .B1(n12738), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n11794), .ZN(n16181) );
  INV_X1 U13266 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n17571) );
  NAND2_X1 U13267 ( .A1(n12738), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11796) );
  AOI22_X1 U13268 ( .A1(n11791), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11795) );
  OAI211_X1 U13269 ( .C1(n12741), .C2(n17571), .A(n11796), .B(n11795), .ZN(
        n16193) );
  NAND2_X1 U13270 ( .A1(n16194), .A2(n16193), .ZN(n16195) );
  INV_X1 U13271 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19260) );
  NAND2_X1 U13272 ( .A1(n11791), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11798) );
  NAND2_X1 U13273 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11797) );
  OAI211_X1 U13274 ( .C1(n12741), .C2(n19260), .A(n11798), .B(n11797), .ZN(
        n11799) );
  AOI21_X1 U13275 ( .B1(n12738), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n11799), .ZN(n16216) );
  INV_X1 U13276 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n17551) );
  NAND2_X1 U13277 ( .A1(n11791), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11801) );
  NAND2_X1 U13278 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11800) );
  OAI211_X1 U13279 ( .C1(n12741), .C2(n17551), .A(n11801), .B(n11800), .ZN(
        n11802) );
  AOI21_X1 U13280 ( .B1(n12738), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n11802), .ZN(n17424) );
  INV_X1 U13281 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n11805) );
  NAND2_X1 U13282 ( .A1(n12738), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11804) );
  AOI22_X1 U13283 ( .A1(n11791), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n11803) );
  OAI211_X1 U13284 ( .C1(n12741), .C2(n11805), .A(n11804), .B(n11803), .ZN(
        n12770) );
  INV_X1 U13285 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n18195) );
  NAND2_X1 U13286 ( .A1(n12738), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11807) );
  AOI22_X1 U13287 ( .A1(n11791), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11806) );
  OAI211_X1 U13288 ( .C1(n12741), .C2(n18195), .A(n11807), .B(n11806), .ZN(
        n17349) );
  NAND2_X1 U13289 ( .A1(n17350), .A2(n17349), .ZN(n14104) );
  INV_X1 U13290 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n18197) );
  NAND2_X1 U13291 ( .A1(n11791), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11809) );
  NAND2_X1 U13292 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n11808) );
  OAI211_X1 U13293 ( .C1(n12741), .C2(n18197), .A(n11809), .B(n11808), .ZN(
        n11810) );
  AOI21_X1 U13294 ( .B1(n12738), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n11810), .ZN(n14106) );
  INV_X1 U13295 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n18198) );
  NAND2_X1 U13296 ( .A1(n11791), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11812) );
  NAND2_X1 U13297 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11811) );
  OAI211_X1 U13298 ( .C1(n11733), .C2(n18198), .A(n11812), .B(n11811), .ZN(
        n11813) );
  AOI21_X1 U13299 ( .B1(n12738), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n11813), .ZN(n17400) );
  INV_X1 U13300 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n18199) );
  NAND2_X1 U13301 ( .A1(n12738), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11815) );
  AOI22_X1 U13302 ( .A1(n11791), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11814) );
  OAI211_X1 U13303 ( .C1(n11733), .C2(n18199), .A(n11815), .B(n11814), .ZN(
        n17335) );
  INV_X1 U13304 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n18200) );
  NAND2_X1 U13305 ( .A1(n11791), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11817) );
  NAND2_X1 U13306 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11816) );
  OAI211_X1 U13307 ( .C1(n11733), .C2(n18200), .A(n11817), .B(n11816), .ZN(
        n11818) );
  AOI21_X1 U13308 ( .B1(n12738), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11818), .ZN(n17387) );
  INV_X1 U13309 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n18201) );
  NAND2_X1 U13310 ( .A1(n11791), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11820) );
  NAND2_X1 U13311 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11819) );
  OAI211_X1 U13312 ( .C1(n11733), .C2(n18201), .A(n11820), .B(n11819), .ZN(
        n11821) );
  AOI21_X1 U13313 ( .B1(n12738), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n11821), .ZN(n14083) );
  INV_X1 U13314 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n14043) );
  NAND2_X1 U13315 ( .A1(n12738), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11823) );
  AOI22_X1 U13316 ( .A1(n11791), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11822) );
  OAI211_X1 U13317 ( .C1(n11733), .C2(n14043), .A(n11823), .B(n11822), .ZN(
        n14041) );
  INV_X1 U13318 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19326) );
  AOI22_X1 U13319 ( .A1(n11791), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11824) );
  OAI21_X1 U13320 ( .B1(n11733), .B2(n19326), .A(n11824), .ZN(n11825) );
  AOI21_X1 U13321 ( .B1(n12738), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n11825), .ZN(n16645) );
  INV_X1 U13322 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n18204) );
  NAND2_X1 U13323 ( .A1(n12738), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11827) );
  AOI22_X1 U13324 ( .A1(n11791), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11826) );
  OAI211_X1 U13325 ( .C1(n11733), .C2(n18204), .A(n11827), .B(n11826), .ZN(
        n12737) );
  NAND2_X1 U13326 ( .A1(n20092), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11829) );
  NAND2_X1 U13327 ( .A1(n11167), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11828) );
  NAND2_X1 U13328 ( .A1(n11829), .A2(n11828), .ZN(n12582) );
  NAND2_X1 U13329 ( .A1(n20094), .A2(n19360), .ZN(n12395) );
  NAND2_X1 U13330 ( .A1(n11836), .A2(n11829), .ZN(n11838) );
  NAND2_X1 U13331 ( .A1(n19998), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11833) );
  NAND2_X1 U13332 ( .A1(n11830), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11831) );
  NAND2_X1 U13333 ( .A1(n11833), .A2(n11831), .ZN(n11837) );
  INV_X1 U13334 ( .A(n11837), .ZN(n11832) );
  NAND2_X1 U13335 ( .A1(n11838), .A2(n11832), .ZN(n11834) );
  NAND2_X1 U13336 ( .A1(n11834), .A2(n11833), .ZN(n11840) );
  MUX2_X1 U13337 ( .A(n19952), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11839) );
  INV_X1 U13338 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19364) );
  INV_X1 U13339 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17967) );
  NOR2_X1 U13340 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17967), .ZN(
        n11835) );
  NAND2_X1 U13341 ( .A1(n12582), .A2(n12395), .ZN(n12624) );
  NAND2_X1 U13342 ( .A1(n11836), .A2(n12624), .ZN(n12583) );
  XNOR2_X1 U13343 ( .A(n11838), .B(n11837), .ZN(n12580) );
  NOR2_X1 U13344 ( .A1(n11840), .A2(n11839), .ZN(n11841) );
  OR2_X1 U13345 ( .A1(n11842), .A2(n11841), .ZN(n12194) );
  NAND3_X1 U13346 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n11843), .A3(
        n19364), .ZN(n12190) );
  INV_X1 U13347 ( .A(n12190), .ZN(n11844) );
  NAND2_X1 U13348 ( .A1(n12580), .A2(n12592), .ZN(n12615) );
  NOR2_X1 U13349 ( .A1(n12583), .A2(n12615), .ZN(n11845) );
  OR2_X1 U13350 ( .A1(n12631), .A2(n11845), .ZN(n15158) );
  AND2_X1 U13351 ( .A1(n12216), .A2(n11846), .ZN(n12702) );
  INV_X1 U13352 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n17963) );
  NAND2_X1 U13353 ( .A1(n19074), .A2(n12581), .ZN(n12215) );
  NAND2_X1 U13354 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19073) );
  INV_X1 U13355 ( .A(n19073), .ZN(n22338) );
  AOI22_X1 U13356 ( .A1(n16472), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16416), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11861) );
  NAND2_X1 U13357 ( .A1(n12024), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11852) );
  AND2_X1 U13358 ( .A1(n11849), .A2(n16489), .ZN(n16449) );
  AND2_X1 U13359 ( .A1(n16489), .A2(n11850), .ZN(n16448) );
  AOI22_X1 U13360 ( .A1(n16449), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16448), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11851) );
  AND2_X1 U13361 ( .A1(n11852), .A2(n11851), .ZN(n11860) );
  INV_X4 U13362 ( .A(n15126), .ZN(n16676) );
  AND2_X2 U13363 ( .A1(n16676), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11944) );
  AOI22_X1 U13364 ( .A1(n12062), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11944), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11859) );
  AND2_X2 U13365 ( .A1(n11855), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16418) );
  INV_X1 U13366 ( .A(n11856), .ZN(n16497) );
  AND2_X2 U13367 ( .A1(n11857), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11939) );
  AOI22_X1 U13368 ( .A1(n16418), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11939), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11858) );
  NAND4_X1 U13369 ( .A1(n11861), .A2(n11860), .A3(n11859), .A4(n11858), .ZN(
        n11871) );
  AND2_X1 U13370 ( .A1(n11862), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11978) );
  AOI22_X1 U13371 ( .A1(n11978), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11905), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U13372 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n16481), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11868) );
  AOI22_X1 U13373 ( .A1(n16482), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n16424), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11867) );
  NAND2_X1 U13374 ( .A1(n16217), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11866) );
  NAND4_X1 U13375 ( .A1(n11869), .A2(n11868), .A3(n11867), .A4(n11866), .ZN(
        n11870) );
  INV_X1 U13376 ( .A(n11163), .ZN(n14387) );
  AND2_X1 U13377 ( .A1(n11872), .A2(n20083), .ZN(n11873) );
  NAND2_X1 U13378 ( .A1(n14387), .A2(n11873), .ZN(n11913) );
  MUX2_X1 U13379 ( .A(n19921), .B(n20094), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11874) );
  NAND2_X1 U13380 ( .A1(n11918), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11879) );
  INV_X1 U13381 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n14417) );
  OAI21_X1 U13382 ( .B1(n19921), .B2(n14417), .A(n20083), .ZN(n11877) );
  AOI21_X1 U13383 ( .B1(n12086), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n11877), .ZN(n11878) );
  NAND2_X1 U13384 ( .A1(n11879), .A2(n11878), .ZN(n14382) );
  NAND2_X1 U13385 ( .A1(n11918), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11881) );
  NOR2_X1 U13386 ( .A1(n19921), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11919) );
  INV_X1 U13387 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14249) );
  AOI22_X1 U13388 ( .A1(n11919), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12086), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11880) );
  NAND2_X1 U13389 ( .A1(n11881), .A2(n11880), .ZN(n11898) );
  INV_X1 U13390 ( .A(n11898), .ZN(n11882) );
  NAND2_X1 U13391 ( .A1(n11163), .A2(n19921), .ZN(n11883) );
  MUX2_X1 U13392 ( .A(n11883), .B(n20092), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11897) );
  AOI22_X1 U13393 ( .A1(n16472), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n16416), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11889) );
  NAND2_X1 U13394 ( .A1(n12024), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11885) );
  AOI22_X1 U13395 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n16449), .B1(
        n16448), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11884) );
  AND2_X1 U13396 ( .A1(n11885), .A2(n11884), .ZN(n11888) );
  AOI22_X1 U13397 ( .A1(n12062), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11944), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11887) );
  AOI22_X1 U13398 ( .A1(n16418), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11939), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11886) );
  NAND4_X1 U13399 ( .A1(n11889), .A2(n11888), .A3(n11887), .A4(n11886), .ZN(
        n11895) );
  AOI22_X1 U13400 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11905), .B1(
        n11978), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U13401 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n16481), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11892) );
  AOI22_X1 U13402 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n16482), .B1(
        n16424), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11891) );
  NAND2_X1 U13403 ( .A1(n16217), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11890) );
  NAND4_X1 U13404 ( .A1(n11893), .A2(n11892), .A3(n11891), .A4(n11890), .ZN(
        n11894) );
  INV_X1 U13405 ( .A(n12647), .ZN(n12333) );
  OR2_X1 U13406 ( .A1(n12333), .A2(n12152), .ZN(n11896) );
  AOI22_X1 U13407 ( .A1(n16472), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16416), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11904) );
  NAND2_X1 U13408 ( .A1(n12024), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11900) );
  AOI22_X1 U13409 ( .A1(n16449), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n16448), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11899) );
  AND2_X1 U13410 ( .A1(n11900), .A2(n11899), .ZN(n11903) );
  AOI22_X1 U13411 ( .A1(n12062), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11944), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11902) );
  AOI22_X1 U13412 ( .A1(n16418), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11939), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11901) );
  NAND4_X1 U13413 ( .A1(n11904), .A2(n11903), .A3(n11902), .A4(n11901), .ZN(
        n11911) );
  AOI22_X1 U13414 ( .A1(n11978), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11905), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U13415 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n16481), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11908) );
  AOI22_X1 U13416 ( .A1(n16482), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n16424), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11907) );
  NAND2_X1 U13417 ( .A1(n16217), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n11906) );
  NAND4_X1 U13418 ( .A1(n11909), .A2(n11908), .A3(n11907), .A4(n11906), .ZN(
        n11910) );
  INV_X1 U13419 ( .A(n12645), .ZN(n11912) );
  OR2_X1 U13420 ( .A1(n11912), .A2(n12152), .ZN(n11914) );
  OAI211_X1 U13421 ( .C1(n19998), .C2(n20083), .A(n11914), .B(n11913), .ZN(
        n11916) );
  NAND2_X1 U13422 ( .A1(n12698), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11921) );
  INV_X2 U13423 ( .A(n12120), .ZN(n12697) );
  AOI22_X1 U13424 ( .A1(n12697), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12086), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11920) );
  NAND2_X1 U13425 ( .A1(n11921), .A2(n11920), .ZN(n14566) );
  AOI22_X1 U13426 ( .A1(n12024), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12062), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11929) );
  INV_X1 U13427 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11924) );
  NAND2_X1 U13428 ( .A1(n16449), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11923) );
  NAND2_X1 U13429 ( .A1(n16482), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11922) );
  OAI211_X1 U13430 ( .C1(n16454), .C2(n11924), .A(n11923), .B(n11922), .ZN(
        n11925) );
  INV_X1 U13431 ( .A(n11925), .ZN(n11928) );
  AOI22_X1 U13432 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16481), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11927) );
  AOI22_X1 U13433 ( .A1(n16416), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11944), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11926) );
  NAND4_X1 U13434 ( .A1(n11929), .A2(n11928), .A3(n11927), .A4(n11926), .ZN(
        n11933) );
  AOI22_X1 U13435 ( .A1(n11978), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11905), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11932) );
  AOI22_X1 U13436 ( .A1(n16418), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11939), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11931) );
  AOI22_X1 U13437 ( .A1(n16424), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n16448), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11930) );
  NAND2_X1 U13438 ( .A1(n12698), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11937) );
  AOI22_X1 U13439 ( .A1(n12086), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11935) );
  NAND2_X1 U13440 ( .A1(n12697), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11934) );
  AND2_X1 U13441 ( .A1(n11935), .A2(n11934), .ZN(n11936) );
  OAI211_X1 U13442 ( .C1(n12152), .C2(n12351), .A(n11937), .B(n11936), .ZN(
        n15198) );
  NAND2_X1 U13443 ( .A1(n15199), .A2(n15198), .ZN(n15200) );
  NAND2_X1 U13444 ( .A1(n12698), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U13445 ( .A1(n12697), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12086), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11957) );
  INV_X1 U13446 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11938) );
  OR2_X1 U13447 ( .A1(n16454), .A2(n11938), .ZN(n11943) );
  NAND2_X1 U13448 ( .A1(n16416), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11942) );
  NAND2_X1 U13449 ( .A1(n16418), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11941) );
  NAND2_X1 U13450 ( .A1(n11939), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11940) );
  AND4_X1 U13451 ( .A1(n11943), .A2(n11942), .A3(n11941), .A4(n11940), .ZN(
        n11955) );
  NAND2_X1 U13452 ( .A1(n12024), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11948) );
  NAND2_X1 U13453 ( .A1(n12062), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11947) );
  AOI22_X1 U13454 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n16449), .B1(
        n16448), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11946) );
  NAND2_X1 U13455 ( .A1(n11944), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11945) );
  AOI22_X1 U13456 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16481), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11954) );
  AOI22_X1 U13457 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n16482), .B1(
        n16424), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11952) );
  NAND2_X1 U13458 ( .A1(n11978), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11951) );
  NAND2_X1 U13459 ( .A1(n11905), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11950) );
  NAND2_X1 U13460 ( .A1(n16217), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11949) );
  AND4_X1 U13461 ( .A1(n11952), .A2(n11951), .A3(n11950), .A4(n11949), .ZN(
        n11953) );
  INV_X1 U13462 ( .A(n12354), .ZN(n12655) );
  OR2_X1 U13463 ( .A1(n12152), .A2(n12655), .ZN(n11956) );
  INV_X1 U13464 ( .A(n12022), .ZN(n12698) );
  INV_X1 U13465 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11959) );
  OR2_X1 U13466 ( .A1(n16454), .A2(n11959), .ZN(n11963) );
  AOI22_X1 U13467 ( .A1(n16482), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16449), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11962) );
  NAND2_X1 U13468 ( .A1(n16418), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11961) );
  NAND2_X1 U13469 ( .A1(n11944), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11960) );
  NAND2_X1 U13470 ( .A1(n12024), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11967) );
  NAND2_X1 U13471 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11966) );
  NAND2_X1 U13472 ( .A1(n16416), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11965) );
  NAND2_X1 U13473 ( .A1(n11939), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11964) );
  AND4_X1 U13474 ( .A1(n11967), .A2(n11966), .A3(n11965), .A4(n11964), .ZN(
        n11974) );
  AOI22_X1 U13475 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16481), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11973) );
  AOI22_X1 U13476 ( .A1(n16424), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n16448), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11971) );
  NAND2_X1 U13477 ( .A1(n11905), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11970) );
  NAND2_X1 U13478 ( .A1(n11978), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11969) );
  NAND2_X1 U13479 ( .A1(n16217), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11968) );
  AND4_X1 U13480 ( .A1(n11971), .A2(n11970), .A3(n11969), .A4(n11968), .ZN(
        n11972) );
  NAND4_X1 U13481 ( .A1(n11523), .A2(n11974), .A3(n11973), .A4(n11972), .ZN(
        n12381) );
  NAND2_X1 U13482 ( .A1(n12381), .A2(n20174), .ZN(n12195) );
  INV_X1 U13483 ( .A(n12195), .ZN(n11975) );
  AOI22_X1 U13484 ( .A1(n12698), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n14377), 
        .B2(n11975), .ZN(n11977) );
  AOI22_X1 U13485 ( .A1(n12697), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12086), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11976) );
  NAND2_X1 U13486 ( .A1(n11977), .A2(n11976), .ZN(n16072) );
  NAND2_X1 U13487 ( .A1(n16073), .A2(n16072), .ZN(n16071) );
  INV_X1 U13488 ( .A(n12152), .ZN(n11996) );
  AOI22_X1 U13489 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n16482), .B1(
        n16424), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11982) );
  NAND2_X1 U13490 ( .A1(n11978), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11981) );
  NAND2_X1 U13491 ( .A1(n11905), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11980) );
  NAND2_X1 U13492 ( .A1(n16217), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11979) );
  NAND4_X1 U13493 ( .A1(n11982), .A2(n11981), .A3(n11980), .A4(n11979), .ZN(
        n11986) );
  NAND2_X1 U13494 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11984) );
  NAND2_X1 U13495 ( .A1(n16481), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11983) );
  NAND2_X1 U13496 ( .A1(n11984), .A2(n11983), .ZN(n11985) );
  NOR2_X1 U13497 ( .A1(n11986), .A2(n11985), .ZN(n11995) );
  NAND2_X1 U13498 ( .A1(n12024), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11991) );
  NAND2_X1 U13499 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11990) );
  AOI22_X1 U13500 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n16449), .B1(
        n16448), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11989) );
  NAND2_X1 U13501 ( .A1(n11944), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11988) );
  AOI22_X1 U13502 ( .A1(n16472), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n16416), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U13503 ( .A1(n16418), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11939), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11992) );
  NAND4_X1 U13504 ( .A1(n11995), .A2(n11994), .A3(n11993), .A4(n11992), .ZN(
        n12442) );
  AOI222_X1 U13505 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n12698), .B1(n12086), 
        .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(P2_EAX_REG_6__SCAN_IN), 
        .C2(n12697), .ZN(n14619) );
  NAND2_X1 U13506 ( .A1(n14618), .A2(n11998), .ZN(n12021) );
  INV_X1 U13507 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16671) );
  OR2_X1 U13508 ( .A1(n16454), .A2(n16671), .ZN(n12002) );
  NAND2_X1 U13509 ( .A1(n16416), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12001) );
  NAND2_X1 U13510 ( .A1(n16418), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12000) );
  NAND2_X1 U13511 ( .A1(n11939), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11999) );
  NAND4_X1 U13512 ( .A1(n12002), .A2(n12001), .A3(n12000), .A4(n11999), .ZN(
        n12008) );
  NAND2_X1 U13513 ( .A1(n12024), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12006) );
  NAND2_X1 U13514 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12005) );
  AOI22_X1 U13515 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n16449), .B1(
        n16448), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12004) );
  NAND2_X1 U13516 ( .A1(n11944), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12003) );
  NAND4_X1 U13517 ( .A1(n12006), .A2(n12005), .A3(n12004), .A4(n12003), .ZN(
        n12007) );
  NOR2_X1 U13518 ( .A1(n12008), .A2(n12007), .ZN(n12018) );
  AOI22_X1 U13519 ( .A1(n16482), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n16424), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12012) );
  NAND2_X1 U13520 ( .A1(n11978), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12011) );
  NAND2_X1 U13521 ( .A1(n11905), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12010) );
  NAND2_X1 U13522 ( .A1(n16217), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12009) );
  NAND4_X1 U13523 ( .A1(n12012), .A2(n12011), .A3(n12010), .A4(n12009), .ZN(
        n12016) );
  NAND2_X1 U13524 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12014) );
  NAND2_X1 U13525 ( .A1(n16481), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12013) );
  NAND2_X1 U13526 ( .A1(n12014), .A2(n12013), .ZN(n12015) );
  NOR2_X1 U13527 ( .A1(n12016), .A2(n12015), .ZN(n12017) );
  INV_X1 U13528 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17904) );
  INV_X1 U13529 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n18163) );
  OAI222_X1 U13530 ( .A1(n17904), .A2(n12023), .B1(n12120), .B2(n18163), .C1(
        n12022), .C2(n11757), .ZN(n14622) );
  NAND2_X1 U13531 ( .A1(n12698), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U13532 ( .A1(n12697), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12086), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U13533 ( .A1(n12024), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n16418), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U13534 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16416), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12031) );
  INV_X1 U13535 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12027) );
  NAND2_X1 U13536 ( .A1(n16449), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12026) );
  NAND2_X1 U13537 ( .A1(n16482), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12025) );
  OAI211_X1 U13538 ( .C1(n16454), .C2(n12027), .A(n12026), .B(n12025), .ZN(
        n12028) );
  INV_X1 U13539 ( .A(n12028), .ZN(n12030) );
  AOI22_X1 U13540 ( .A1(n16481), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11944), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12029) );
  NAND4_X1 U13541 ( .A1(n12032), .A2(n12031), .A3(n12030), .A4(n12029), .ZN(
        n12038) );
  AOI22_X1 U13542 ( .A1(n11978), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16217), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U13543 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11939), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12035) );
  AOI22_X1 U13544 ( .A1(n16424), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n16448), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12034) );
  NAND2_X1 U13545 ( .A1(n11905), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12033) );
  NAND4_X1 U13546 ( .A1(n12036), .A2(n12035), .A3(n12034), .A4(n12033), .ZN(
        n12037) );
  INV_X1 U13547 ( .A(n14991), .ZN(n12039) );
  OR2_X1 U13548 ( .A1(n12152), .A2(n12039), .ZN(n12040) );
  AOI22_X1 U13549 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n16472), .B1(
        n16416), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12047) );
  INV_X1 U13550 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12320) );
  INV_X1 U13551 ( .A(n16449), .ZN(n16474) );
  INV_X1 U13552 ( .A(n16448), .ZN(n16473) );
  INV_X1 U13553 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n16117) );
  OAI22_X1 U13554 ( .A1(n12320), .A2(n16474), .B1(n16473), .B2(n16117), .ZN(
        n12043) );
  AOI21_X1 U13555 ( .B1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n12024), .A(
        n12043), .ZN(n12046) );
  AOI22_X1 U13556 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11944), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U13557 ( .A1(n16418), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11939), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12044) );
  NAND4_X1 U13558 ( .A1(n12047), .A2(n12046), .A3(n12045), .A4(n12044), .ZN(
        n12053) );
  AOI22_X1 U13559 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n11905), .B1(
        n11978), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12051) );
  AOI22_X1 U13560 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n16481), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U13561 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n16482), .B1(
        n16424), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12049) );
  NAND2_X1 U13562 ( .A1(n16217), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12048) );
  NAND4_X1 U13563 ( .A1(n12051), .A2(n12050), .A3(n12049), .A4(n12048), .ZN(
        n12052) );
  NOR2_X1 U13564 ( .A1(n12053), .A2(n12052), .ZN(n15190) );
  NAND2_X1 U13565 ( .A1(n12698), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12055) );
  AOI22_X1 U13566 ( .A1(n12697), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12086), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12054) );
  OAI211_X1 U13567 ( .C1(n12152), .C2(n15190), .A(n12055), .B(n12054), .ZN(
        n14667) );
  NAND2_X1 U13568 ( .A1(n12698), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U13569 ( .A1(n12697), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12086), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U13570 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n16418), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12059) );
  AOI22_X1 U13571 ( .A1(n11978), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16217), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12058) );
  AOI22_X1 U13572 ( .A1(n16482), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n16424), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12057) );
  NAND2_X1 U13573 ( .A1(n11905), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12056) );
  NAND4_X1 U13574 ( .A1(n12059), .A2(n12058), .A3(n12057), .A4(n12056), .ZN(
        n12068) );
  INV_X1 U13575 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12060) );
  INV_X1 U13576 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n16198) );
  OAI22_X1 U13577 ( .A1(n16474), .A2(n12060), .B1(n16473), .B2(n16198), .ZN(
        n12061) );
  AOI21_X1 U13578 ( .B1(n12024), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n12061), .ZN(n12066) );
  AOI22_X1 U13579 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16481), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U13580 ( .A1(n16416), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11944), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U13581 ( .A1(n16472), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11939), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12063) );
  NAND4_X1 U13582 ( .A1(n12066), .A2(n12065), .A3(n12064), .A4(n12063), .ZN(
        n12067) );
  OR2_X1 U13583 ( .A1(n12152), .A2(n15369), .ZN(n12069) );
  NOR2_X2 U13584 ( .A1(n14668), .A2(n14737), .ZN(n14818) );
  AOI22_X1 U13585 ( .A1(n16472), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16416), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12077) );
  INV_X1 U13586 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16558) );
  INV_X1 U13587 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12072) );
  OAI22_X1 U13588 ( .A1(n16474), .A2(n16558), .B1(n16473), .B2(n12072), .ZN(
        n12073) );
  AOI21_X1 U13589 ( .B1(n12024), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n12073), .ZN(n12076) );
  AOI22_X1 U13590 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11944), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12075) );
  AOI22_X1 U13591 ( .A1(n16418), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11939), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12074) );
  NAND4_X1 U13592 ( .A1(n12077), .A2(n12076), .A3(n12075), .A4(n12074), .ZN(
        n12083) );
  AOI22_X1 U13593 ( .A1(n11978), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11905), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12081) );
  AOI22_X1 U13594 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n16481), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U13595 ( .A1(n16482), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16424), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12079) );
  NAND2_X1 U13596 ( .A1(n16217), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12078) );
  NAND4_X1 U13597 ( .A1(n12081), .A2(n12080), .A3(n12079), .A4(n12078), .ZN(
        n12082) );
  NOR2_X1 U13598 ( .A1(n12083), .A2(n12082), .ZN(n15486) );
  NAND2_X1 U13599 ( .A1(n12698), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12085) );
  AOI22_X1 U13600 ( .A1(n12697), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12086), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12084) );
  OAI211_X1 U13601 ( .C1(n12152), .C2(n15486), .A(n12085), .B(n12084), .ZN(
        n14819) );
  NAND2_X1 U13602 ( .A1(n12698), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12106) );
  AOI22_X1 U13603 ( .A1(n12697), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12086), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U13604 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n16472), .B1(
        n16416), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12096) );
  INV_X1 U13605 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16426) );
  INV_X1 U13606 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12087) );
  OAI22_X1 U13607 ( .A1(n16426), .A2(n16474), .B1(n16473), .B2(n12087), .ZN(
        n12088) );
  AOI21_X1 U13608 ( .B1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B2(n12024), .A(
        n12088), .ZN(n12095) );
  INV_X1 U13609 ( .A(n11987), .ZN(n12091) );
  INV_X1 U13610 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12090) );
  INV_X1 U13611 ( .A(n11944), .ZN(n12124) );
  INV_X1 U13612 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12089) );
  OAI22_X1 U13613 ( .A1(n12091), .A2(n12090), .B1(n12124), .B2(n12089), .ZN(
        n12092) );
  INV_X1 U13614 ( .A(n12092), .ZN(n12094) );
  AOI22_X1 U13615 ( .A1(n16418), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11939), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12093) );
  NAND4_X1 U13616 ( .A1(n12096), .A2(n12095), .A3(n12094), .A4(n12093), .ZN(
        n12102) );
  AOI22_X1 U13617 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11978), .B1(
        n11905), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U13618 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n16481), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12099) );
  AOI22_X1 U13619 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n16482), .B1(
        n16424), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12098) );
  NAND2_X1 U13620 ( .A1(n16217), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12097) );
  NAND4_X1 U13621 ( .A1(n12100), .A2(n12099), .A3(n12098), .A4(n12097), .ZN(
        n12101) );
  INV_X1 U13622 ( .A(n15536), .ZN(n12103) );
  OR2_X1 U13623 ( .A1(n12152), .A2(n12103), .ZN(n12104) );
  AOI22_X1 U13624 ( .A1(n16472), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16416), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12113) );
  INV_X1 U13625 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12108) );
  INV_X1 U13626 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12107) );
  OAI22_X1 U13627 ( .A1(n16474), .A2(n12108), .B1(n16473), .B2(n12107), .ZN(
        n12109) );
  AOI21_X1 U13628 ( .B1(n12024), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n12109), .ZN(n12112) );
  AOI22_X1 U13629 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11944), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12111) );
  AOI22_X1 U13630 ( .A1(n16418), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11939), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12110) );
  NAND4_X1 U13631 ( .A1(n12113), .A2(n12112), .A3(n12111), .A4(n12110), .ZN(
        n12119) );
  AOI22_X1 U13632 ( .A1(n11978), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11905), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12117) );
  AOI22_X1 U13633 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n16481), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12116) );
  AOI22_X1 U13634 ( .A1(n16482), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16424), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12115) );
  NAND2_X1 U13635 ( .A1(n16217), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12114) );
  NAND4_X1 U13636 ( .A1(n12117), .A2(n12116), .A3(n12115), .A4(n12114), .ZN(
        n12118) );
  OR2_X1 U13637 ( .A1(n12119), .A2(n12118), .ZN(n15535) );
  INV_X1 U13638 ( .A(n15535), .ZN(n12123) );
  NAND2_X1 U13639 ( .A1(n12698), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U13640 ( .A1(n12697), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11873), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12121) );
  OAI211_X1 U13641 ( .C1(n12152), .C2(n12123), .A(n12122), .B(n12121), .ZN(
        n15188) );
  AOI22_X1 U13642 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n12024), .B1(
        n16418), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U13643 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n11987), .B1(
        n16416), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12130) );
  INV_X1 U13644 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12430) );
  INV_X1 U13645 ( .A(n16481), .ZN(n16441) );
  INV_X1 U13646 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16456) );
  OAI22_X1 U13647 ( .A1(n12430), .A2(n12124), .B1(n16441), .B2(n16456), .ZN(
        n12128) );
  INV_X1 U13648 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16459) );
  NAND2_X1 U13649 ( .A1(n16449), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12126) );
  NAND2_X1 U13650 ( .A1(n16482), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12125) );
  OAI211_X1 U13651 ( .C1(n16458), .C2(n16459), .A(n12126), .B(n12125), .ZN(
        n12127) );
  NOR2_X1 U13652 ( .A1(n12128), .A2(n12127), .ZN(n12129) );
  NAND3_X1 U13653 ( .A1(n12131), .A2(n12130), .A3(n12129), .ZN(n12137) );
  AOI22_X1 U13654 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n16472), .B1(
        n16226), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12135) );
  AOI22_X1 U13655 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n16217), .B1(
        n11978), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U13656 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n16448), .B1(
        n16424), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12133) );
  NAND2_X1 U13657 ( .A1(n11905), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12132) );
  NAND4_X1 U13658 ( .A1(n12135), .A2(n12134), .A3(n12133), .A4(n12132), .ZN(
        n12136) );
  OR2_X1 U13659 ( .A1(n12137), .A2(n12136), .ZN(n16112) );
  INV_X1 U13660 ( .A(n16112), .ZN(n12140) );
  NAND2_X1 U13661 ( .A1(n12698), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U13662 ( .A1(n12697), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11873), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12138) );
  OAI211_X1 U13663 ( .C1(n12152), .C2(n12140), .A(n12139), .B(n12138), .ZN(
        n15319) );
  NAND2_X1 U13664 ( .A1(n12698), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12155) );
  AOI22_X1 U13665 ( .A1(n12697), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11873), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U13666 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n16472), .B1(
        n16416), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12145) );
  INV_X1 U13667 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16670) );
  INV_X1 U13668 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16475) );
  OAI22_X1 U13669 ( .A1(n16670), .A2(n16474), .B1(n16473), .B2(n16475), .ZN(
        n12141) );
  AOI21_X1 U13670 ( .B1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n12024), .A(
        n12141), .ZN(n12144) );
  AOI22_X1 U13671 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11944), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12143) );
  AOI22_X1 U13672 ( .A1(n16418), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11939), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12142) );
  NAND4_X1 U13673 ( .A1(n12145), .A2(n12144), .A3(n12143), .A4(n12142), .ZN(
        n12151) );
  AOI22_X1 U13674 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n11905), .B1(
        n11978), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U13675 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n16481), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U13676 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n16482), .B1(
        n16424), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12147) );
  NAND2_X1 U13677 ( .A1(n16217), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12146) );
  NAND4_X1 U13678 ( .A1(n12149), .A2(n12148), .A3(n12147), .A4(n12146), .ZN(
        n12150) );
  NOR2_X1 U13679 ( .A1(n12151), .A2(n12150), .ZN(n16111) );
  OR2_X1 U13680 ( .A1(n12152), .A2(n16111), .ZN(n12153) );
  NAND2_X1 U13681 ( .A1(n12698), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U13682 ( .A1(n12697), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11873), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12156) );
  NOR2_X4 U13683 ( .A1(n16171), .A2(n16170), .ZN(n16172) );
  NAND2_X1 U13684 ( .A1(n12698), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U13685 ( .A1(n12697), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11873), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12158) );
  NAND2_X1 U13686 ( .A1(n12159), .A2(n12158), .ZN(n16132) );
  NAND2_X1 U13687 ( .A1(n12698), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12161) );
  AOI22_X1 U13688 ( .A1(n12697), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11873), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12160) );
  AND2_X1 U13689 ( .A1(n12161), .A2(n12160), .ZN(n17767) );
  NAND2_X1 U13690 ( .A1(n11918), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12163) );
  AOI22_X1 U13691 ( .A1(n12697), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11873), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12162) );
  NAND2_X1 U13692 ( .A1(n11918), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12165) );
  AOI22_X1 U13693 ( .A1(n12697), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11873), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12164) );
  NAND2_X1 U13694 ( .A1(n12165), .A2(n12164), .ZN(n17742) );
  AND2_X2 U13695 ( .A1(n17743), .A2(n17742), .ZN(n17740) );
  NAND2_X1 U13696 ( .A1(n11918), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U13697 ( .A1(n12697), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11873), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12166) );
  NAND2_X1 U13698 ( .A1(n12167), .A2(n12166), .ZN(n12781) );
  NAND2_X1 U13699 ( .A1(n12698), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U13700 ( .A1(n12697), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11873), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12168) );
  AND2_X1 U13701 ( .A1(n12169), .A2(n12168), .ZN(n17353) );
  NAND2_X1 U13702 ( .A1(n11918), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12171) );
  AOI22_X1 U13703 ( .A1(n12697), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11873), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12170) );
  NAND2_X1 U13704 ( .A1(n12171), .A2(n12170), .ZN(n14108) );
  NAND2_X1 U13705 ( .A1(n11918), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12173) );
  AOI22_X1 U13706 ( .A1(n12697), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11873), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12172) );
  AND2_X1 U13707 ( .A1(n12173), .A2(n12172), .ZN(n17456) );
  NAND2_X1 U13708 ( .A1(n11918), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12175) );
  AOI22_X1 U13709 ( .A1(n12697), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11873), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12174) );
  NAND2_X1 U13710 ( .A1(n12175), .A2(n12174), .ZN(n17338) );
  NAND2_X1 U13711 ( .A1(n17337), .A2(n17338), .ZN(n17336) );
  NAND2_X1 U13712 ( .A1(n11918), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12177) );
  AOI22_X1 U13713 ( .A1(n12697), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11873), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12176) );
  AND2_X1 U13714 ( .A1(n12177), .A2(n12176), .ZN(n17442) );
  NAND2_X1 U13715 ( .A1(n11918), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U13716 ( .A1(n12697), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11873), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12178) );
  NAND2_X1 U13717 ( .A1(n11918), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U13718 ( .A1(n12697), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11873), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12180) );
  AND2_X1 U13719 ( .A1(n12181), .A2(n12180), .ZN(n14050) );
  NAND2_X1 U13720 ( .A1(n11918), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12183) );
  AOI22_X1 U13721 ( .A1(n11919), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11873), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12182) );
  NAND2_X1 U13722 ( .A1(n12183), .A2(n12182), .ZN(n16648) );
  NAND2_X1 U13723 ( .A1(n11918), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12185) );
  AOI22_X1 U13724 ( .A1(n11919), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11873), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12184) );
  NAND2_X1 U13725 ( .A1(n12185), .A2(n12184), .ZN(n12186) );
  INV_X1 U13726 ( .A(n12800), .ZN(n12227) );
  AND2_X1 U13727 ( .A1(n12188), .A2(n20429), .ZN(n12633) );
  INV_X1 U13728 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n22310) );
  INV_X1 U13729 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n18185) );
  NAND2_X1 U13730 ( .A1(n18185), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n22341) );
  INV_X2 U13731 ( .A(n22341), .ZN(n18205) );
  INV_X1 U13732 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n22354) );
  NAND2_X1 U13733 ( .A1(n18205), .A2(n22354), .ZN(n18207) );
  NOR2_X1 U13734 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_0__SCAN_IN), 
        .ZN(n17957) );
  NAND2_X1 U13735 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n17957), .ZN(n18184) );
  NAND2_X1 U13736 ( .A1(n18202), .A2(n18184), .ZN(n19084) );
  INV_X1 U13737 ( .A(n19084), .ZN(n22347) );
  NOR2_X1 U13738 ( .A1(n22338), .A2(n22347), .ZN(n15164) );
  NAND2_X1 U13739 ( .A1(n22310), .A2(n15164), .ZN(n12218) );
  INV_X1 U13740 ( .A(n12218), .ZN(n12189) );
  AND2_X1 U13741 ( .A1(n12633), .A2(n12189), .ZN(n15176) );
  NAND2_X1 U13742 ( .A1(n19074), .A2(n15176), .ZN(n19336) );
  INV_X1 U13743 ( .A(n19336), .ZN(n19348) );
  MUX2_X1 U13744 ( .A(n12190), .B(n12354), .S(n12581), .Z(n12628) );
  INV_X1 U13745 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n12191) );
  MUX2_X1 U13746 ( .A(n12628), .B(n12191), .S(n12211), .Z(n12412) );
  MUX2_X1 U13747 ( .A(n12645), .B(n12580), .S(n12641), .Z(n12623) );
  INV_X1 U13748 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n14609) );
  MUX2_X1 U13749 ( .A(n12623), .B(n14609), .S(n12211), .Z(n12402) );
  NOR2_X1 U13750 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n12193) );
  MUX2_X1 U13751 ( .A(n12647), .B(n12193), .S(n12211), .Z(n12401) );
  NAND2_X1 U13752 ( .A1(n12402), .A2(n12401), .ZN(n12408) );
  OAI21_X1 U13753 ( .B1(n20174), .B2(P2_EBX_REG_5__SCAN_IN), .A(n12195), .ZN(
        n12196) );
  INV_X1 U13754 ( .A(n12196), .ZN(n12391) );
  INV_X1 U13755 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n12197) );
  MUX2_X1 U13756 ( .A(n12197), .B(n12442), .S(n20174), .Z(n12445) );
  MUX2_X1 U13757 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n12685), .S(n20174), .Z(
        n12451) );
  OR2_X2 U13758 ( .A1(n12450), .A2(n12451), .ZN(n12455) );
  INV_X1 U13759 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n12198) );
  NAND2_X1 U13760 ( .A1(n12211), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12458) );
  NAND2_X1 U13761 ( .A1(n12211), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12456) );
  INV_X1 U13762 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n12199) );
  NAND2_X1 U13763 ( .A1(n12211), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12472) );
  INV_X1 U13764 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n12200) );
  NOR2_X1 U13765 ( .A1(n20174), .A2(n12200), .ZN(n12512) );
  INV_X1 U13766 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n12201) );
  NOR2_X1 U13767 ( .A1(n20174), .A2(n12201), .ZN(n12516) );
  INV_X1 U13768 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n12202) );
  NOR2_X1 U13769 ( .A1(n20174), .A2(n12202), .ZN(n12509) );
  INV_X1 U13770 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n12203) );
  NOR2_X1 U13771 ( .A1(n20174), .A2(n12203), .ZN(n12504) );
  NAND2_X1 U13772 ( .A1(n12211), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12501) );
  INV_X1 U13773 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n12204) );
  NOR2_X1 U13774 ( .A1(n20174), .A2(n12204), .ZN(n12491) );
  INV_X1 U13775 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n12205) );
  NOR2_X1 U13776 ( .A1(n20174), .A2(n12205), .ZN(n12487) );
  NAND2_X1 U13777 ( .A1(n12211), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12495) );
  INV_X1 U13778 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n12206) );
  NOR2_X1 U13779 ( .A1(n20174), .A2(n12206), .ZN(n12485) );
  NAND2_X1 U13780 ( .A1(n12211), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12538) );
  INV_X1 U13781 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n12207) );
  NOR2_X1 U13782 ( .A1(n20174), .A2(n12207), .ZN(n12543) );
  NAND2_X1 U13783 ( .A1(n12211), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12547) );
  INV_X1 U13784 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n12208) );
  NOR2_X1 U13785 ( .A1(n20174), .A2(n12208), .ZN(n12554) );
  INV_X1 U13786 ( .A(n12550), .ZN(n12209) );
  NAND2_X1 U13787 ( .A1(n12211), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12549) );
  INV_X1 U13788 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n12210) );
  NOR2_X1 U13789 ( .A1(n20174), .A2(n12210), .ZN(n12557) );
  NAND2_X1 U13790 ( .A1(n12211), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12561) );
  INV_X1 U13791 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n12212) );
  NOR2_X1 U13792 ( .A1(n20174), .A2(n12212), .ZN(n12569) );
  NAND2_X1 U13793 ( .A1(n12211), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12213) );
  INV_X1 U13794 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n12219) );
  NAND2_X1 U13795 ( .A1(n22310), .A2(n19073), .ZN(n12220) );
  INV_X1 U13796 ( .A(n12220), .ZN(n12214) );
  NAND2_X1 U13797 ( .A1(n12572), .A2(n19323), .ZN(n12225) );
  OR2_X1 U13798 ( .A1(n12216), .A2(n19448), .ZN(n12217) );
  NOR2_X2 U13799 ( .A1(n14198), .A2(n19079), .ZN(n14549) );
  NAND2_X1 U13800 ( .A1(n14549), .A2(n12218), .ZN(n19341) );
  INV_X1 U13801 ( .A(n14198), .ZN(n14199) );
  NAND3_X1 U13802 ( .A1(n14199), .A2(n12220), .A3(n12219), .ZN(n12221) );
  NAND2_X2 U13803 ( .A1(n19341), .A2(n12221), .ZN(n19328) );
  NOR2_X1 U13804 ( .A1(n19436), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19441) );
  INV_X1 U13805 ( .A(n19441), .ZN(n19428) );
  NOR3_X1 U13806 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n20083), .A3(n19428), 
        .ZN(n19440) );
  NOR2_X2 U13807 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20100) );
  NAND2_X1 U13808 ( .A1(n20100), .A2(n17963), .ZN(n18027) );
  INV_X1 U13809 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19999) );
  NAND4_X1 U13810 ( .A1(n19436), .A2(n19999), .A3(n22310), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19432) );
  NAND2_X1 U13811 ( .A1(n19380), .A2(n19432), .ZN(n12222) );
  OR2_X1 U13812 ( .A1(n19440), .A2(n12222), .ZN(n12223) );
  NAND2_X1 U13813 ( .A1(n19338), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19237) );
  INV_X2 U13814 ( .A(n19237), .ZN(n19346) );
  AOI22_X1 U13815 ( .A1(n19328), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n19346), .ZN(n12224) );
  INV_X1 U13816 ( .A(n12229), .ZN(n12283) );
  OR2_X1 U13817 ( .A1(n19338), .A2(n18204), .ZN(n12282) );
  INV_X1 U13818 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12732) );
  AND2_X1 U13819 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12230) );
  AND2_X2 U13820 ( .A1(n12254), .A2(n12230), .ZN(n12255) );
  NAND2_X2 U13821 ( .A1(n12255), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12259) );
  NOR2_X4 U13822 ( .A1(n12259), .A2(n17641), .ZN(n12253) );
  NAND2_X1 U13823 ( .A1(n12253), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12260) );
  INV_X1 U13824 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18077) );
  INV_X1 U13825 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n19177) );
  INV_X1 U13826 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17616) );
  INV_X1 U13827 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12246) );
  INV_X1 U13828 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17558) );
  INV_X1 U13829 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12768) );
  INV_X1 U13830 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17512) );
  NOR2_X2 U13831 ( .A1(n12237), .A2(n17512), .ZN(n12238) );
  NAND2_X1 U13832 ( .A1(n12238), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12235) );
  INV_X1 U13833 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17489) );
  OR2_X2 U13834 ( .A1(n12235), .A2(n17489), .ZN(n12273) );
  INV_X1 U13835 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12272) );
  INV_X1 U13836 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16705) );
  NOR2_X4 U13837 ( .A1(n12275), .A2(n16705), .ZN(n12276) );
  NAND2_X1 U13838 ( .A1(n12276), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12234) );
  INV_X1 U13839 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12233) );
  INV_X1 U13840 ( .A(n12273), .ZN(n12236) );
  AOI21_X1 U13841 ( .B1(n17489), .B2(n12271), .A(n12236), .ZN(n17487) );
  AOI21_X1 U13842 ( .B1(n17512), .B2(n12237), .A(n12238), .ZN(n17515) );
  AOI21_X1 U13843 ( .B1(n12239), .B2(n12232), .A(n12240), .ZN(n17532) );
  CLKBUF_X1 U13844 ( .A(n12241), .Z(n12268) );
  AOI21_X1 U13845 ( .B1(n12768), .B2(n12268), .A(n12242), .ZN(n14091) );
  AOI21_X1 U13846 ( .B1(n17558), .B2(n12266), .A(n12243), .ZN(n19264) );
  CLKBUF_X1 U13847 ( .A(n12244), .Z(n12264) );
  AOI21_X1 U13848 ( .B1(n12264), .B2(n12231), .A(n12245), .ZN(n19236) );
  NAND2_X1 U13849 ( .A1(n12246), .A2(n12263), .ZN(n12248) );
  INV_X1 U13850 ( .A(n12265), .ZN(n12247) );
  AND2_X1 U13851 ( .A1(n12248), .A2(n12247), .ZN(n17606) );
  AOI21_X1 U13852 ( .B1(n12262), .B2(n17616), .A(n12249), .ZN(n19193) );
  CLKBUF_X1 U13853 ( .A(n12250), .Z(n12261) );
  AOI21_X1 U13854 ( .B1(n19177), .B2(n12261), .A(n12251), .ZN(n17625) );
  AOI21_X1 U13855 ( .B1(n18077), .B2(n12260), .A(n12252), .ZN(n19156) );
  AOI21_X1 U13856 ( .B1(n17641), .B2(n12259), .A(n12253), .ZN(n19140) );
  INV_X1 U13857 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12256) );
  NAND2_X1 U13858 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n11175), .ZN(
        n12258) );
  AOI21_X1 U13859 ( .B1(n12256), .B2(n12258), .A(n12255), .ZN(n19121) );
  AOI21_X1 U13860 ( .B1(n15402), .B2(n12257), .A(n11175), .ZN(n15400) );
  OAI22_X1 U13861 ( .A1(n19436), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n19100) );
  INV_X1 U13862 ( .A(n19100), .ZN(n16060) );
  AOI22_X1 U13863 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14249), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19436), .ZN(n16059) );
  NOR2_X1 U13864 ( .A1(n16060), .A2(n16059), .ZN(n16058) );
  OAI21_X1 U13865 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n12257), .ZN(n18031) );
  NAND2_X1 U13866 ( .A1(n16058), .A2(n18031), .ZN(n15383) );
  NOR2_X1 U13867 ( .A1(n15400), .A2(n15383), .ZN(n15494) );
  OAI21_X1 U13868 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n11175), .A(
        n12258), .ZN(n18039) );
  NAND2_X1 U13869 ( .A1(n15494), .A2(n18039), .ZN(n19119) );
  NOR2_X1 U13870 ( .A1(n19121), .A2(n19119), .ZN(n19127) );
  OAI21_X1 U13871 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12255), .A(
        n12259), .ZN(n19129) );
  NAND2_X1 U13872 ( .A1(n19127), .A2(n19129), .ZN(n19139) );
  NOR2_X1 U13873 ( .A1(n19140), .A2(n19139), .ZN(n17363) );
  OAI21_X1 U13874 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12253), .A(
        n12260), .ZN(n18069) );
  NAND2_X1 U13875 ( .A1(n17363), .A2(n18069), .ZN(n19154) );
  NOR2_X1 U13876 ( .A1(n19156), .A2(n19154), .ZN(n19165) );
  OAI21_X1 U13877 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12252), .A(
        n12261), .ZN(n19166) );
  NAND2_X1 U13878 ( .A1(n19165), .A2(n19166), .ZN(n19181) );
  NOR2_X1 U13879 ( .A1(n17625), .A2(n19181), .ZN(n15519) );
  OAI21_X1 U13880 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12251), .A(
        n12262), .ZN(n18101) );
  NAND2_X1 U13881 ( .A1(n15519), .A2(n18101), .ZN(n19192) );
  NOR2_X1 U13882 ( .A1(n19193), .A2(n19192), .ZN(n19200) );
  OAI21_X1 U13883 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n12249), .A(
        n12263), .ZN(n19201) );
  NAND2_X1 U13884 ( .A1(n19200), .A2(n19201), .ZN(n19217) );
  NOR2_X1 U13885 ( .A1(n17606), .A2(n19217), .ZN(n19218) );
  OAI21_X1 U13886 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12265), .A(
        n12264), .ZN(n19227) );
  NAND2_X1 U13887 ( .A1(n19218), .A2(n19227), .ZN(n19234) );
  NOR2_X1 U13888 ( .A1(n19236), .A2(n19234), .ZN(n19247) );
  OAI21_X1 U13889 ( .B1(n12245), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n12266), .ZN(n19248) );
  NAND2_X1 U13890 ( .A1(n19247), .A2(n19248), .ZN(n19262) );
  NOR2_X1 U13891 ( .A1(n19264), .A2(n19262), .ZN(n19278) );
  OR2_X1 U13892 ( .A1(n12243), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12267) );
  NAND2_X1 U13893 ( .A1(n12268), .A2(n12267), .ZN(n19281) );
  INV_X1 U13894 ( .A(n16057), .ZN(n12269) );
  AOI21_X2 U13895 ( .B1(n19278), .B2(n19281), .A(n12269), .ZN(n19277) );
  OAI21_X1 U13896 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12242), .A(
        n12239), .ZN(n17543) );
  INV_X1 U13897 ( .A(n17543), .ZN(n17358) );
  NOR2_X1 U13898 ( .A1(n17359), .A2(n17358), .ZN(n17357) );
  NOR2_X1 U13899 ( .A1(n17532), .A2(n14100), .ZN(n14099) );
  OAI21_X1 U13900 ( .B1(n12240), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n12237), .ZN(n17522) );
  INV_X1 U13901 ( .A(n17522), .ZN(n19288) );
  NOR2_X1 U13902 ( .A1(n11181), .A2(n19287), .ZN(n17344) );
  NOR2_X1 U13903 ( .A1(n17515), .A2(n17344), .ZN(n17343) );
  NOR2_X2 U13904 ( .A1(n17343), .A2(n11181), .ZN(n19300) );
  OR2_X1 U13905 ( .A1(n12238), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12270) );
  NAND2_X1 U13906 ( .A1(n12271), .A2(n12270), .ZN(n17504) );
  INV_X1 U13907 ( .A(n17504), .ZN(n19299) );
  NOR2_X1 U13908 ( .A1(n19300), .A2(n19299), .ZN(n19298) );
  NOR2_X1 U13909 ( .A1(n11181), .A2(n19298), .ZN(n14079) );
  NOR2_X1 U13910 ( .A1(n17487), .A2(n14079), .ZN(n14078) );
  NAND2_X1 U13911 ( .A1(n12273), .A2(n12272), .ZN(n12274) );
  NAND2_X1 U13912 ( .A1(n12275), .A2(n12274), .ZN(n19313) );
  AOI21_X1 U13913 ( .B1(n14078), .B2(n19313), .A(n11181), .ZN(n19330) );
  AOI21_X1 U13914 ( .B1(n16705), .B2(n12275), .A(n12276), .ZN(n19329) );
  NAND2_X1 U13915 ( .A1(n16057), .A2(n19332), .ZN(n12279) );
  INV_X1 U13916 ( .A(n12279), .ZN(n12278) );
  XNOR2_X1 U13917 ( .A(n12276), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16406) );
  INV_X1 U13918 ( .A(n16406), .ZN(n12277) );
  NAND3_X1 U13919 ( .A1(n12280), .A2(n19354), .A3(n19316), .ZN(n12281) );
  NAND3_X1 U13920 ( .A1(n12283), .A2(n12282), .A3(n12281), .ZN(P2_U2825) );
  XNOR2_X2 U13921 ( .A(n12285), .B(n12284), .ZN(n14592) );
  BUF_X2 U13922 ( .A(n14592), .Z(n18033) );
  XNOR2_X2 U13923 ( .A(n12287), .B(n12286), .ZN(n14705) );
  NAND2_X1 U13924 ( .A1(n18033), .A2(n14705), .ZN(n12328) );
  INV_X1 U13925 ( .A(n12328), .ZN(n12296) );
  INV_X1 U13926 ( .A(n12289), .ZN(n12291) );
  INV_X1 U13927 ( .A(n12290), .ZN(n12299) );
  NAND2_X1 U13928 ( .A1(n12291), .A2(n12299), .ZN(n12292) );
  NAND2_X1 U13929 ( .A1(n19954), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12306) );
  OR2_X2 U13930 ( .A1(n14592), .A2(n12300), .ZN(n12307) );
  INV_X1 U13931 ( .A(n19105), .ZN(n14664) );
  NOR2_X1 U13932 ( .A1(n12307), .A2(n14664), .ZN(n12308) );
  INV_X1 U13933 ( .A(n12288), .ZN(n12298) );
  NAND2_X1 U13934 ( .A1(n12298), .A2(n12297), .ZN(n12327) );
  NOR2_X1 U13935 ( .A1(n12303), .A2(n12314), .ZN(n12359) );
  AOI22_X1 U13936 ( .A1(n12355), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12359), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12305) );
  INV_X1 U13937 ( .A(n12301), .ZN(n12302) );
  AND2_X2 U13938 ( .A1(n12303), .A2(n12302), .ZN(n19990) );
  NAND3_X1 U13939 ( .A1(n12306), .A2(n12305), .A3(n12304), .ZN(n12311) );
  NOR2_X1 U13940 ( .A1(n12307), .A2(n19105), .ZN(n12316) );
  INV_X1 U13941 ( .A(n12309), .ZN(n12310) );
  NAND2_X2 U13942 ( .A1(n12312), .A2(n18033), .ZN(n12326) );
  INV_X1 U13943 ( .A(n12314), .ZN(n12315) );
  OAI211_X1 U13944 ( .C1(n12346), .C2(n12320), .A(n12319), .B(n12318), .ZN(
        n12323) );
  NAND2_X1 U13945 ( .A1(n19105), .A2(n16344), .ZN(n12324) );
  NOR2_X2 U13946 ( .A1(n12326), .A2(n12324), .ZN(n12364) );
  INV_X1 U13947 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n16116) );
  NOR2_X2 U13948 ( .A1(n12326), .A2(n12327), .ZN(n12365) );
  NAND2_X1 U13949 ( .A1(n12365), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12321) );
  OAI21_X1 U13950 ( .B1(n20021), .B2(n16116), .A(n12321), .ZN(n12322) );
  NOR2_X1 U13951 ( .A1(n12323), .A2(n12322), .ZN(n12331) );
  INV_X1 U13952 ( .A(n12371), .ZN(n19942) );
  NAND4_X1 U13953 ( .A1(n12332), .A2(n12331), .A3(n12330), .A4(n12329), .ZN(
        n12335) );
  NAND2_X1 U13954 ( .A1(n12188), .A2(n12396), .ZN(n16337) );
  NOR2_X1 U13955 ( .A1(n16337), .A2(n12333), .ZN(n12644) );
  OR2_X1 U13956 ( .A1(n12644), .A2(n12645), .ZN(n12334) );
  AND2_X2 U13957 ( .A1(n12335), .A2(n12334), .ZN(n12393) );
  AOI22_X1 U13958 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19975), .B1(
        n12355), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U13959 ( .A1(n12359), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12358), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U13960 ( .A1(n12357), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n19990), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12337) );
  AOI22_X1 U13961 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12356), .B1(
        n12317), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12336) );
  INV_X1 U13962 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12341) );
  INV_X1 U13963 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12340) );
  INV_X1 U13964 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12343) );
  INV_X1 U13965 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12342) );
  NOR2_X1 U13966 ( .A1(n12345), .A2(n12344), .ZN(n12349) );
  AOI22_X1 U13967 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12364), .B1(
        n20036), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12348) );
  INV_X1 U13968 ( .A(n12346), .ZN(n12366) );
  NAND4_X1 U13969 ( .A1(n12350), .A2(n12349), .A3(n12348), .A4(n12347), .ZN(
        n12353) );
  NAND2_X1 U13970 ( .A1(n12351), .A2(n12188), .ZN(n12352) );
  AND2_X2 U13971 ( .A1(n12353), .A2(n12352), .ZN(n12394) );
  AOI22_X1 U13972 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19975), .B1(
        n12355), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12363) );
  AOI22_X1 U13973 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n12317), .B1(
        n12356), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12362) );
  AOI22_X1 U13974 ( .A1(n12357), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12358), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U13975 ( .A1(n20070), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n19990), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U13976 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n12364), .B1(
        n20036), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12379) );
  AOI22_X1 U13977 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n12365), .B1(
        n12366), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12378) );
  INV_X1 U13978 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12370) );
  INV_X1 U13979 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12369) );
  OAI22_X1 U13980 ( .A1(n12370), .A2(n12367), .B1(n12368), .B2(n12369), .ZN(
        n12376) );
  INV_X1 U13981 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12374) );
  INV_X1 U13982 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12372) );
  OAI22_X1 U13983 ( .A1(n12374), .A2(n12373), .B1(n12371), .B2(n12372), .ZN(
        n12375) );
  NOR2_X1 U13984 ( .A1(n12376), .A2(n12375), .ZN(n12377) );
  NAND4_X1 U13985 ( .A1(n12380), .A2(n12379), .A3(n12378), .A4(n12377), .ZN(
        n12384) );
  INV_X1 U13986 ( .A(n12381), .ZN(n12382) );
  NAND2_X1 U13987 ( .A1(n12382), .A2(n12188), .ZN(n12383) );
  NAND2_X1 U13988 ( .A1(n12384), .A2(n12383), .ZN(n12386) );
  NAND2_X1 U13989 ( .A1(n12657), .A2(n12386), .ZN(n12389) );
  INV_X1 U13990 ( .A(n12385), .ZN(n12388) );
  INV_X1 U13991 ( .A(n12386), .ZN(n12387) );
  NAND2_X2 U13992 ( .A1(n12388), .A2(n12387), .ZN(n12679) );
  XNOR2_X1 U13993 ( .A(n12390), .B(n12391), .ZN(n19114) );
  INV_X1 U13994 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16075) );
  OAI21_X1 U13995 ( .B1(n20094), .B2(n19360), .A(n12395), .ZN(n12616) );
  INV_X1 U13996 ( .A(n12616), .ZN(n12585) );
  MUX2_X1 U13997 ( .A(n12396), .B(n12585), .S(n12641), .Z(n12625) );
  MUX2_X1 U13998 ( .A(n12625), .B(P2_EBX_REG_0__SCAN_IN), .S(n12211), .Z(
        n19091) );
  INV_X1 U13999 ( .A(n19091), .ZN(n12398) );
  INV_X1 U14000 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12397) );
  NOR2_X1 U14001 ( .A1(n12398), .A2(n12397), .ZN(n16334) );
  NAND2_X1 U14002 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n12399) );
  NOR2_X1 U14003 ( .A1(n20174), .A2(n12399), .ZN(n12400) );
  NOR2_X1 U14004 ( .A1(n12401), .A2(n12400), .ZN(n19101) );
  NOR2_X1 U14005 ( .A1(n16334), .A2(n19101), .ZN(n14244) );
  INV_X1 U14006 ( .A(n14244), .ZN(n14245) );
  NAND2_X1 U14007 ( .A1(n16334), .A2(n19101), .ZN(n14246) );
  NAND2_X1 U14008 ( .A1(n14249), .A2(n14246), .ZN(n14243) );
  NAND2_X1 U14009 ( .A1(n14245), .A2(n14243), .ZN(n14560) );
  INV_X1 U14010 ( .A(n14560), .ZN(n12404) );
  OR2_X1 U14011 ( .A1(n12402), .A2(n12401), .ZN(n12403) );
  NAND2_X1 U14012 ( .A1(n12408), .A2(n12403), .ZN(n15512) );
  XNOR2_X1 U14013 ( .A(n15512), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14558) );
  NAND2_X1 U14014 ( .A1(n12404), .A2(n14558), .ZN(n14562) );
  INV_X1 U14015 ( .A(n15512), .ZN(n12405) );
  NAND2_X1 U14016 ( .A1(n12405), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12406) );
  NAND2_X1 U14017 ( .A1(n14562), .A2(n12406), .ZN(n15399) );
  XNOR2_X1 U14018 ( .A(n12408), .B(n11334), .ZN(n15397) );
  AOI21_X1 U14019 ( .B1(n15399), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n15397), .ZN(n12409) );
  OAI21_X1 U14020 ( .B1(n15395), .B2(n12019), .A(n12409), .ZN(n12411) );
  OR2_X1 U14021 ( .A1(n15399), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12410) );
  NAND2_X1 U14022 ( .A1(n12411), .A2(n12410), .ZN(n15471) );
  OAI21_X1 U14023 ( .B1(n12413), .B2(n12412), .A(n12390), .ZN(n15502) );
  INV_X1 U14024 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16076) );
  XNOR2_X1 U14025 ( .A(n15502), .B(n16076), .ZN(n15470) );
  INV_X1 U14026 ( .A(n15502), .ZN(n12414) );
  NAND2_X1 U14027 ( .A1(n12414), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12415) );
  NAND2_X1 U14028 ( .A1(n15473), .A2(n12415), .ZN(n16083) );
  NAND2_X1 U14029 ( .A1(n12416), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12417) );
  NAND2_X1 U14030 ( .A1(n16082), .A2(n12417), .ZN(n17915) );
  INV_X1 U14031 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12420) );
  INV_X1 U14032 ( .A(n12355), .ZN(n12419) );
  INV_X1 U14033 ( .A(n19975), .ZN(n12418) );
  INV_X1 U14034 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16626) );
  OAI22_X1 U14035 ( .A1(n12420), .A2(n12419), .B1(n12418), .B2(n16626), .ZN(
        n12423) );
  INV_X1 U14036 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20162) );
  INV_X1 U14037 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16453) );
  OAI22_X1 U14038 ( .A1(n20162), .A2(n16023), .B1(n12421), .B2(n16453), .ZN(
        n12422) );
  NOR2_X1 U14039 ( .A1(n12423), .A2(n12422), .ZN(n12441) );
  INV_X1 U14040 ( .A(n20036), .ZN(n20033) );
  INV_X1 U14041 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12424) );
  INV_X1 U14042 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16457) );
  OAI22_X1 U14043 ( .A1(n20033), .A2(n12424), .B1(n12368), .B2(n16457), .ZN(
        n12427) );
  INV_X1 U14044 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12425) );
  OAI22_X1 U14045 ( .A1(n12425), .A2(n12367), .B1(n12371), .B2(n16459), .ZN(
        n12426) );
  NOR2_X1 U14046 ( .A1(n12427), .A2(n12426), .ZN(n12440) );
  INV_X1 U14047 ( .A(n12358), .ZN(n12429) );
  INV_X1 U14048 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12428) );
  OAI22_X1 U14049 ( .A1(n11176), .A2(n12430), .B1(n12429), .B2(n12428), .ZN(
        n12434) );
  INV_X1 U14050 ( .A(n20070), .ZN(n12432) );
  INV_X1 U14051 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n20150) );
  INV_X1 U14052 ( .A(n19990), .ZN(n12431) );
  OAI22_X1 U14053 ( .A1(n12432), .A2(n20150), .B1(n12431), .B2(n16456), .ZN(
        n12433) );
  NOR2_X1 U14054 ( .A1(n12434), .A2(n12433), .ZN(n12439) );
  NAND2_X1 U14055 ( .A1(n12364), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12438) );
  NAND2_X1 U14056 ( .A1(n12365), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12437) );
  NAND2_X1 U14057 ( .A1(n12366), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12436) );
  NAND2_X1 U14058 ( .A1(n19923), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12435) );
  NAND4_X1 U14059 ( .A1(n12441), .A2(n12440), .A3(n12439), .A4(n11526), .ZN(
        n12444) );
  OR2_X1 U14060 ( .A1(n19079), .A2(n12442), .ZN(n12443) );
  XNOR2_X2 U14061 ( .A(n12679), .B(n12680), .ZN(n12676) );
  NAND2_X1 U14062 ( .A1(n12676), .A2(n12685), .ZN(n12447) );
  XNOR2_X1 U14063 ( .A(n12446), .B(n12445), .ZN(n19130) );
  NAND2_X1 U14064 ( .A1(n12447), .A2(n19130), .ZN(n12448) );
  NAND2_X1 U14065 ( .A1(n12448), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12449) );
  INV_X1 U14066 ( .A(n12451), .ZN(n12452) );
  XNOR2_X1 U14067 ( .A(n12450), .B(n12452), .ZN(n19142) );
  AND2_X1 U14068 ( .A1(n19142), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17635) );
  INV_X1 U14069 ( .A(n12453), .ZN(n12454) );
  XNOR2_X1 U14070 ( .A(n12455), .B(n12454), .ZN(n17366) );
  NAND2_X1 U14071 ( .A1(n17366), .A2(n12019), .ZN(n18064) );
  INV_X1 U14072 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12463) );
  NOR2_X1 U14073 ( .A1(n18064), .A2(n12463), .ZN(n12467) );
  OR2_X1 U14074 ( .A1(n12461), .A2(n12456), .ZN(n12457) );
  AND2_X1 U14075 ( .A1(n12470), .A2(n12457), .ZN(n12479) );
  INV_X1 U14076 ( .A(n12479), .ZN(n19163) );
  INV_X1 U14077 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17865) );
  OAI21_X1 U14078 ( .B1(n19163), .B2(n12685), .A(n17865), .ZN(n17876) );
  NOR2_X1 U14079 ( .A1(n12459), .A2(n12458), .ZN(n12460) );
  OR2_X1 U14080 ( .A1(n12461), .A2(n12460), .ZN(n19151) );
  NOR2_X1 U14081 ( .A1(n19151), .A2(n12685), .ZN(n12477) );
  INV_X1 U14082 ( .A(n12477), .ZN(n12462) );
  INV_X1 U14083 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17895) );
  NAND2_X1 U14084 ( .A1(n12462), .A2(n17895), .ZN(n17887) );
  NAND2_X1 U14085 ( .A1(n18064), .A2(n12463), .ZN(n12465) );
  INV_X1 U14086 ( .A(n19142), .ZN(n12464) );
  NAND2_X1 U14087 ( .A1(n12464), .A2(n17904), .ZN(n18063) );
  AND4_X1 U14088 ( .A1(n17876), .A2(n17887), .A3(n12465), .A4(n18063), .ZN(
        n12466) );
  INV_X1 U14089 ( .A(n12468), .ZN(n12469) );
  XNOR2_X1 U14090 ( .A(n12470), .B(n12469), .ZN(n19180) );
  INV_X1 U14091 ( .A(n12471), .ZN(n12474) );
  INV_X1 U14092 ( .A(n12472), .ZN(n12473) );
  NAND2_X1 U14093 ( .A1(n12474), .A2(n12473), .ZN(n12475) );
  NAND2_X1 U14094 ( .A1(n12513), .A2(n12475), .ZN(n15528) );
  OR2_X1 U14095 ( .A1(n15528), .A2(n12685), .ZN(n12483) );
  INV_X1 U14096 ( .A(n12483), .ZN(n12476) );
  NAND2_X1 U14097 ( .A1(n12476), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18088) );
  NAND2_X1 U14098 ( .A1(n12477), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17888) );
  NOR2_X1 U14099 ( .A1(n12685), .A2(n17865), .ZN(n12478) );
  NAND2_X1 U14100 ( .A1(n12479), .A2(n12478), .ZN(n17875) );
  NAND2_X1 U14101 ( .A1(n17888), .A2(n17875), .ZN(n17630) );
  INV_X1 U14102 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17853) );
  NOR2_X1 U14103 ( .A1(n12685), .A2(n17853), .ZN(n12480) );
  AND2_X1 U14104 ( .A1(n19180), .A2(n12480), .ZN(n17627) );
  OR2_X1 U14105 ( .A1(n17630), .A2(n17627), .ZN(n18085) );
  INV_X1 U14106 ( .A(n18085), .ZN(n12481) );
  AND2_X1 U14107 ( .A1(n18088), .A2(n12481), .ZN(n12482) );
  INV_X1 U14108 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n19393) );
  NAND2_X1 U14109 ( .A1(n12483), .A2(n19393), .ZN(n18087) );
  NAND2_X1 U14110 ( .A1(n12499), .A2(n12485), .ZN(n12486) );
  AND2_X1 U14111 ( .A1(n12539), .A2(n12486), .ZN(n14092) );
  NAND2_X1 U14112 ( .A1(n14092), .A2(n12019), .ZN(n12523) );
  INV_X1 U14113 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12780) );
  NAND2_X1 U14114 ( .A1(n12523), .A2(n12780), .ZN(n12758) );
  INV_X1 U14115 ( .A(n12487), .ZN(n12488) );
  XNOR2_X1 U14116 ( .A(n12489), .B(n12488), .ZN(n19257) );
  NAND2_X1 U14117 ( .A1(n19257), .A2(n12019), .ZN(n12535) );
  INV_X1 U14118 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17761) );
  NAND2_X1 U14119 ( .A1(n12535), .A2(n17761), .ZN(n17560) );
  INV_X1 U14120 ( .A(n12491), .ZN(n12492) );
  XNOR2_X1 U14121 ( .A(n12490), .B(n12492), .ZN(n19250) );
  NAND2_X1 U14122 ( .A1(n19250), .A2(n12019), .ZN(n12493) );
  INV_X1 U14123 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17756) );
  NAND2_X1 U14124 ( .A1(n12493), .A2(n17756), .ZN(n17569) );
  AND2_X1 U14125 ( .A1(n17560), .A2(n17569), .ZN(n12755) );
  INV_X1 U14126 ( .A(n12494), .ZN(n12497) );
  INV_X1 U14127 ( .A(n12495), .ZN(n12496) );
  NAND2_X1 U14128 ( .A1(n12497), .A2(n12496), .ZN(n12498) );
  NAND2_X1 U14129 ( .A1(n12499), .A2(n12498), .ZN(n19272) );
  INV_X1 U14130 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17550) );
  INV_X1 U14131 ( .A(n12500), .ZN(n12506) );
  INV_X1 U14132 ( .A(n12501), .ZN(n12502) );
  NAND2_X1 U14133 ( .A1(n12506), .A2(n12502), .ZN(n12503) );
  NAND2_X1 U14134 ( .A1(n12490), .A2(n12503), .ZN(n19238) );
  INV_X1 U14135 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17794) );
  NAND2_X1 U14136 ( .A1(n12525), .A2(n17794), .ZN(n17579) );
  NAND2_X1 U14137 ( .A1(n12511), .A2(n12504), .ZN(n12505) );
  NAND2_X1 U14138 ( .A1(n12506), .A2(n12505), .ZN(n19225) );
  NAND2_X1 U14139 ( .A1(n12019), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12507) );
  INV_X1 U14140 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17806) );
  OAI21_X1 U14141 ( .B1(n19225), .B2(n12685), .A(n17806), .ZN(n12508) );
  NAND2_X1 U14142 ( .A1(n12519), .A2(n12509), .ZN(n12510) );
  NAND2_X1 U14143 ( .A1(n11210), .A2(n12019), .ZN(n12527) );
  INV_X1 U14144 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17815) );
  NAND2_X1 U14145 ( .A1(n12527), .A2(n17815), .ZN(n17599) );
  NAND2_X1 U14146 ( .A1(n12513), .A2(n12512), .ZN(n12514) );
  NAND2_X1 U14147 ( .A1(n12517), .A2(n12514), .ZN(n19189) );
  OR2_X1 U14148 ( .A1(n19189), .A2(n12685), .ZN(n12515) );
  INV_X1 U14149 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17842) );
  NAND2_X1 U14150 ( .A1(n12515), .A2(n17842), .ZN(n17613) );
  NAND2_X1 U14151 ( .A1(n12517), .A2(n12516), .ZN(n12518) );
  NAND2_X1 U14152 ( .A1(n12519), .A2(n12518), .ZN(n19204) );
  NOR2_X1 U14153 ( .A1(n19204), .A2(n12685), .ZN(n12529) );
  NOR2_X1 U14154 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n12529), .ZN(
        n17602) );
  INV_X1 U14155 ( .A(n17602), .ZN(n17822) );
  AND2_X1 U14156 ( .A1(n17613), .A2(n17822), .ZN(n12520) );
  AND2_X1 U14157 ( .A1(n17599), .A2(n12520), .ZN(n12751) );
  NAND3_X1 U14158 ( .A1(n17579), .A2(n17591), .A3(n12751), .ZN(n12521) );
  AOI21_X1 U14159 ( .B1(n12757), .B2(n17550), .A(n12521), .ZN(n12522) );
  INV_X1 U14160 ( .A(n12523), .ZN(n12524) );
  NAND2_X1 U14161 ( .A1(n12524), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12759) );
  INV_X1 U14162 ( .A(n12757), .ZN(n12534) );
  INV_X1 U14163 ( .A(n12525), .ZN(n12526) );
  NAND2_X1 U14164 ( .A1(n12526), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17580) );
  INV_X1 U14165 ( .A(n12527), .ZN(n12528) );
  NAND2_X1 U14166 ( .A1(n12528), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17600) );
  NAND2_X1 U14167 ( .A1(n12529), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17823) );
  NAND2_X1 U14168 ( .A1(n17600), .A2(n17823), .ZN(n12750) );
  OR3_X1 U14169 ( .A1(n19189), .A2(n12685), .A3(n17842), .ZN(n17612) );
  NAND2_X1 U14170 ( .A1(n12753), .A2(n17612), .ZN(n12530) );
  NOR2_X1 U14171 ( .A1(n12750), .A2(n12530), .ZN(n12532) );
  NOR2_X1 U14172 ( .A1(n12685), .A2(n17756), .ZN(n12531) );
  NAND2_X1 U14173 ( .A1(n19250), .A2(n12531), .ZN(n17568) );
  NAND3_X1 U14174 ( .A1(n17580), .A2(n12532), .A3(n17568), .ZN(n12533) );
  AOI21_X1 U14175 ( .B1(n12534), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n12533), .ZN(n12537) );
  INV_X1 U14176 ( .A(n12535), .ZN(n12536) );
  NAND2_X1 U14177 ( .A1(n12536), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17561) );
  XNOR2_X1 U14178 ( .A(n12539), .B(n12538), .ZN(n17354) );
  NAND2_X1 U14179 ( .A1(n17354), .A2(n12019), .ZN(n12540) );
  XNOR2_X1 U14180 ( .A(n12540), .B(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17542) );
  NAND2_X1 U14181 ( .A1(n17540), .A2(n17542), .ZN(n17541) );
  INV_X1 U14182 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17708) );
  NAND2_X1 U14183 ( .A1(n12540), .A2(n17708), .ZN(n12541) );
  INV_X1 U14184 ( .A(n12542), .ZN(n12548) );
  NAND2_X1 U14185 ( .A1(n12544), .A2(n12543), .ZN(n12545) );
  AND2_X1 U14186 ( .A1(n12548), .A2(n12545), .ZN(n14101) );
  AOI21_X1 U14187 ( .B1(n14101), .B2(n12019), .A(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17528) );
  AND2_X1 U14188 ( .A1(n12019), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12546) );
  NAND2_X1 U14189 ( .A1(n14101), .A2(n12546), .ZN(n17529) );
  XNOR2_X1 U14190 ( .A(n12548), .B(n12547), .ZN(n19283) );
  INV_X1 U14191 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17671) );
  NAND2_X1 U14192 ( .A1(n12551), .A2(n17671), .ZN(n12553) );
  NOR2_X1 U14193 ( .A1(n12685), .A2(n17671), .ZN(n12552) );
  NAND2_X1 U14194 ( .A1(n19295), .A2(n12552), .ZN(n12568) );
  NAND2_X1 U14195 ( .A1(n12553), .A2(n12568), .ZN(n17500) );
  INV_X1 U14196 ( .A(n12554), .ZN(n12555) );
  XNOR2_X1 U14197 ( .A(n12556), .B(n12555), .ZN(n17347) );
  NAND2_X1 U14198 ( .A1(n17347), .A2(n12019), .ZN(n12567) );
  INV_X1 U14199 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17691) );
  NAND2_X1 U14200 ( .A1(n12558), .A2(n12557), .ZN(n12559) );
  NAND2_X1 U14201 ( .A1(n12560), .A2(n12559), .ZN(n14080) );
  NAND2_X1 U14202 ( .A1(n14034), .A2(n11536), .ZN(n12564) );
  XNOR2_X1 U14203 ( .A(n12562), .B(n12561), .ZN(n19306) );
  INV_X1 U14204 ( .A(n14038), .ZN(n12565) );
  INV_X1 U14205 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16700) );
  NAND2_X1 U14206 ( .A1(n12565), .A2(n16700), .ZN(n12566) );
  XNOR2_X1 U14207 ( .A(n12570), .B(n12569), .ZN(n12573) );
  INV_X1 U14208 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16699) );
  OAI21_X1 U14209 ( .B1(n12573), .B2(n12685), .A(n16699), .ZN(n16696) );
  INV_X1 U14210 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12804) );
  NOR2_X1 U14211 ( .A1(n12685), .A2(n12804), .ZN(n12571) );
  NAND2_X1 U14212 ( .A1(n12572), .A2(n12571), .ZN(n12793) );
  INV_X1 U14213 ( .A(n12573), .ZN(n19324) );
  NAND3_X1 U14214 ( .A1(n19324), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12019), .ZN(n16695) );
  NOR2_X1 U14215 ( .A1(n12574), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12575) );
  MUX2_X1 U14216 ( .A(n12450), .B(n12575), .S(n12211), .Z(n19340) );
  NAND2_X1 U14217 ( .A1(n19340), .A2(n12019), .ZN(n12576) );
  XNOR2_X1 U14218 ( .A(n12578), .B(n12577), .ZN(n16405) );
  INV_X1 U14219 ( .A(n12631), .ZN(n12595) );
  NAND2_X1 U14220 ( .A1(n12597), .A2(n19079), .ZN(n12579) );
  MUX2_X1 U14221 ( .A(n12579), .B(n12641), .S(n12580), .Z(n12591) );
  INV_X1 U14222 ( .A(n12580), .ZN(n12588) );
  OAI21_X1 U14223 ( .B1(n12616), .B2(n12582), .A(n12581), .ZN(n12587) );
  INV_X1 U14224 ( .A(n12583), .ZN(n12584) );
  OAI211_X1 U14225 ( .C1(n19079), .C2(n12585), .A(n19080), .B(n12584), .ZN(
        n12586) );
  OAI211_X1 U14226 ( .C1(n12589), .C2(n12588), .A(n12587), .B(n12586), .ZN(
        n12590) );
  NAND2_X1 U14227 ( .A1(n12591), .A2(n12590), .ZN(n12593) );
  MUX2_X1 U14228 ( .A(n12641), .B(n12593), .S(n12592), .Z(n12594) );
  NAND2_X1 U14229 ( .A1(n12595), .A2(n12594), .ZN(n12596) );
  MUX2_X1 U14230 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n12596), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n12599) );
  INV_X1 U14231 ( .A(n12597), .ZN(n14267) );
  NAND2_X1 U14232 ( .A1(n12631), .A2(n14267), .ZN(n12598) );
  NAND2_X1 U14233 ( .A1(n16020), .A2(n19079), .ZN(n12639) );
  NAND2_X1 U14234 ( .A1(n20330), .A2(n15164), .ZN(n12638) );
  AOI21_X1 U14235 ( .B1(n12599), .B2(n19080), .A(n20233), .ZN(n12600) );
  NAND2_X1 U14236 ( .A1(n12639), .A2(n12600), .ZN(n12637) );
  NAND2_X1 U14237 ( .A1(n12601), .A2(n15164), .ZN(n12602) );
  OR2_X1 U14238 ( .A1(n15158), .A2(n12602), .ZN(n12612) );
  NAND2_X1 U14239 ( .A1(n12604), .A2(n12603), .ZN(n12611) );
  NAND2_X1 U14240 ( .A1(n12605), .A2(n19921), .ZN(n12606) );
  NAND2_X1 U14241 ( .A1(n12606), .A2(n12633), .ZN(n12706) );
  AOI21_X1 U14242 ( .B1(n19921), .B2(n20429), .A(n20330), .ZN(n12607) );
  NAND2_X1 U14243 ( .A1(n12717), .A2(n12607), .ZN(n12608) );
  NAND4_X1 U14244 ( .A1(n12706), .A2(n11699), .A3(n12609), .A4(n12608), .ZN(
        n12610) );
  AOI21_X1 U14245 ( .B1(n11846), .B2(n12611), .A(n12610), .ZN(n12719) );
  AND2_X1 U14246 ( .A1(n12612), .A2(n12719), .ZN(n15104) );
  MUX2_X1 U14247 ( .A(n12601), .B(n20330), .S(n12188), .Z(n12613) );
  NAND2_X1 U14248 ( .A1(n12613), .A2(n19073), .ZN(n12621) );
  INV_X1 U14249 ( .A(n15158), .ZN(n12614) );
  OAI21_X1 U14250 ( .B1(n12616), .B2(n12615), .A(n12614), .ZN(n12617) );
  INV_X1 U14251 ( .A(n12617), .ZN(n12619) );
  NAND2_X1 U14252 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16490) );
  OAI21_X1 U14253 ( .B1(n16490), .B2(n11167), .A(n19364), .ZN(n15167) );
  INV_X1 U14254 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12618) );
  OAI21_X1 U14255 ( .B1(n12024), .B2(n15167), .A(n12618), .ZN(n18113) );
  MUX2_X1 U14256 ( .A(n12619), .B(n18113), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n17965) );
  NAND2_X1 U14257 ( .A1(n17965), .A2(n19079), .ZN(n12620) );
  OAI22_X1 U14258 ( .A1(n15158), .A2(n12621), .B1(n12642), .B2(n12620), .ZN(
        n12622) );
  INV_X1 U14259 ( .A(n12622), .ZN(n12635) );
  AOI21_X1 U14260 ( .B1(n12625), .B2(n12624), .A(n12623), .ZN(n12630) );
  INV_X1 U14261 ( .A(n12626), .ZN(n12627) );
  NAND2_X1 U14262 ( .A1(n12628), .A2(n12627), .ZN(n12629) );
  NOR2_X1 U14263 ( .A1(n12630), .A2(n12629), .ZN(n12632) );
  OR2_X1 U14264 ( .A1(n12632), .A2(n12631), .ZN(n15156) );
  INV_X1 U14265 ( .A(n15156), .ZN(n12634) );
  INV_X1 U14266 ( .A(n12633), .ZN(n19083) );
  NOR2_X1 U14267 ( .A1(n12642), .A2(n19083), .ZN(n15155) );
  NAND2_X1 U14268 ( .A1(n12634), .A2(n15155), .ZN(n12763) );
  AND3_X1 U14269 ( .A1(n15104), .A2(n12635), .A3(n12763), .ZN(n12636) );
  OAI211_X1 U14270 ( .C1(n12639), .C2(n12638), .A(n12637), .B(n12636), .ZN(
        n12640) );
  INV_X1 U14271 ( .A(n12746), .ZN(n12643) );
  NOR2_X1 U14272 ( .A1(n12642), .A2(n12641), .ZN(n15153) );
  XOR2_X1 U14273 ( .A(n12645), .B(n12644), .Z(n14565) );
  XOR2_X1 U14274 ( .A(n12647), .B(n12646), .Z(n12648) );
  NAND2_X1 U14275 ( .A1(n16337), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16336) );
  NOR2_X1 U14276 ( .A1(n12648), .A2(n16336), .ZN(n12649) );
  XNOR2_X1 U14277 ( .A(n12648), .B(n16336), .ZN(n14248) );
  NOR2_X1 U14278 ( .A1(n14249), .A2(n14248), .ZN(n14247) );
  NOR2_X1 U14279 ( .A1(n12649), .A2(n14247), .ZN(n12650) );
  XOR2_X1 U14280 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12650), .Z(
        n14564) );
  NOR2_X1 U14281 ( .A1(n14565), .A2(n14564), .ZN(n14563) );
  INV_X1 U14282 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14557) );
  NOR2_X1 U14283 ( .A1(n12650), .A2(n14557), .ZN(n12651) );
  OR2_X1 U14284 ( .A1(n14563), .A2(n12651), .ZN(n12653) );
  XNOR2_X1 U14285 ( .A(n12653), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15396) );
  NAND2_X1 U14286 ( .A1(n12653), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12654) );
  NAND2_X1 U14287 ( .A1(n11217), .A2(n12655), .ZN(n12656) );
  INV_X1 U14288 ( .A(n12658), .ZN(n12660) );
  NAND2_X1 U14289 ( .A1(n12660), .A2(n12659), .ZN(n12661) );
  INV_X1 U14290 ( .A(n12663), .ZN(n12671) );
  NAND2_X1 U14291 ( .A1(n16069), .A2(n12664), .ZN(n12675) );
  OAI21_X1 U14292 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n12676), .A(
        n12666), .ZN(n12673) );
  INV_X1 U14293 ( .A(n12676), .ZN(n12667) );
  OAI21_X1 U14294 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n12668), .A(
        n12667), .ZN(n12669) );
  INV_X1 U14295 ( .A(n12669), .ZN(n12670) );
  NAND2_X1 U14296 ( .A1(n12671), .A2(n12670), .ZN(n12672) );
  NAND2_X1 U14297 ( .A1(n12677), .A2(n12676), .ZN(n12678) );
  XNOR2_X1 U14298 ( .A(n12686), .B(n12685), .ZN(n12682) );
  XNOR2_X1 U14299 ( .A(n12682), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17638) );
  INV_X1 U14300 ( .A(n12682), .ZN(n12683) );
  NAND2_X1 U14301 ( .A1(n12683), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12684) );
  INV_X1 U14302 ( .A(n12687), .ZN(n12688) );
  NAND2_X1 U14303 ( .A1(n12688), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12689) );
  NAND2_X1 U14304 ( .A1(n18059), .A2(n12689), .ZN(n17615) );
  NAND3_X1 U14305 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n19379) );
  NAND2_X1 U14306 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12690) );
  NOR2_X1 U14307 ( .A1(n19379), .A2(n12690), .ZN(n17830) );
  AND2_X1 U14308 ( .A1(n17830), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17734) );
  NAND2_X1 U14309 ( .A1(n17615), .A2(n17734), .ZN(n12764) );
  NAND2_X1 U14310 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12779) );
  NAND2_X1 U14311 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12691) );
  NOR2_X1 U14312 ( .A1(n12779), .A2(n12691), .ZN(n12692) );
  AND3_X1 U14313 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17738) );
  NAND2_X1 U14314 ( .A1(n12692), .A2(n17738), .ZN(n12726) );
  INV_X1 U14315 ( .A(n12726), .ZN(n12693) );
  INV_X1 U14316 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17709) );
  OR2_X1 U14317 ( .A1(n17709), .A2(n17708), .ZN(n12694) );
  NAND2_X1 U14318 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17674) );
  NOR2_X2 U14319 ( .A1(n17497), .A2(n17674), .ZN(n17492) );
  NAND4_X1 U14320 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A4(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12731) );
  INV_X1 U14321 ( .A(n12731), .ZN(n12695) );
  XNOR2_X1 U14322 ( .A(n11528), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16396) );
  INV_X1 U14323 ( .A(n15155), .ZN(n12696) );
  AOI222_X1 U14324 ( .A1(n12698), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12697), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n11873), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12699) );
  INV_X1 U14325 ( .A(n12699), .ZN(n12700) );
  INV_X1 U14326 ( .A(n12702), .ZN(n15157) );
  AND2_X1 U14327 ( .A1(n12703), .A2(n15112), .ZN(n15163) );
  AOI21_X1 U14328 ( .B1(n15157), .B2(n19079), .A(n15163), .ZN(n12704) );
  INV_X1 U14329 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19339) );
  NOR2_X1 U14330 ( .A1(n19380), .A2(n19339), .ZN(n16397) );
  NAND2_X1 U14331 ( .A1(n12705), .A2(n19079), .ZN(n15113) );
  AOI21_X1 U14332 ( .B1(n15113), .B2(n12706), .A(n11677), .ZN(n12713) );
  INV_X1 U14333 ( .A(n14370), .ZN(n14181) );
  NAND2_X1 U14334 ( .A1(n11699), .A2(n20233), .ZN(n12708) );
  AOI22_X1 U14335 ( .A1(n14181), .A2(n12708), .B1(n20330), .B2(n20429), .ZN(
        n12711) );
  NAND2_X1 U14336 ( .A1(n12710), .A2(n12709), .ZN(n14368) );
  NAND3_X1 U14337 ( .A1(n12707), .A2(n12711), .A3(n14368), .ZN(n12712) );
  NOR2_X1 U14338 ( .A1(n12713), .A2(n12712), .ZN(n12714) );
  OAI21_X1 U14339 ( .B1(n12715), .B2(n11699), .A(n12714), .ZN(n15150) );
  NOR2_X1 U14340 ( .A1(n15150), .A2(n15127), .ZN(n12716) );
  NOR2_X1 U14341 ( .A1(n12397), .A2(n14249), .ZN(n14556) );
  NAND2_X1 U14342 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14556), .ZN(
        n14568) );
  INV_X1 U14343 ( .A(n12717), .ZN(n12718) );
  AND2_X1 U14344 ( .A1(n12719), .A2(n12718), .ZN(n14367) );
  INV_X1 U14345 ( .A(n14367), .ZN(n15161) );
  OAI21_X1 U14346 ( .B1(n17787), .B2(n14568), .A(n17923), .ZN(n19411) );
  INV_X1 U14347 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12720) );
  NOR2_X1 U14348 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14556), .ZN(
        n15474) );
  NOR4_X1 U14349 ( .A1(n16076), .A2(n12720), .A3(n16075), .A4(n15474), .ZN(
        n17924) );
  NAND2_X1 U14350 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17924), .ZN(
        n17900) );
  NAND2_X1 U14351 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19401) );
  NOR2_X1 U14352 ( .A1(n17900), .A2(n19401), .ZN(n12723) );
  NAND2_X1 U14353 ( .A1(n17896), .A2(n17734), .ZN(n17793) );
  NOR2_X1 U14354 ( .A1(n17709), .A2(n17708), .ZN(n17707) );
  NAND2_X1 U14355 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17707), .ZN(
        n12721) );
  NOR2_X1 U14356 ( .A1(n17727), .A2(n12721), .ZN(n17692) );
  INV_X1 U14357 ( .A(n17674), .ZN(n12722) );
  NAND2_X1 U14358 ( .A1(n17692), .A2(n12722), .ZN(n14052) );
  NOR3_X1 U14359 ( .A1(n14052), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12731), .ZN(n12734) );
  NAND2_X1 U14360 ( .A1(n17923), .A2(n17787), .ZN(n19378) );
  INV_X1 U14361 ( .A(n19378), .ZN(n17791) );
  NAND2_X1 U14362 ( .A1(n12746), .A2(n19380), .ZN(n14555) );
  NAND2_X1 U14363 ( .A1(n17791), .A2(n14555), .ZN(n12729) );
  NAND2_X1 U14364 ( .A1(n12729), .A2(n17674), .ZN(n12730) );
  INV_X1 U14365 ( .A(n12729), .ZN(n17851) );
  OAI21_X1 U14366 ( .B1(n17923), .B2(n12723), .A(n14555), .ZN(n17735) );
  OR2_X1 U14367 ( .A1(n17900), .A2(n14568), .ZN(n17901) );
  NOR2_X1 U14368 ( .A1(n19401), .A2(n17901), .ZN(n17732) );
  NOR2_X1 U14369 ( .A1(n17787), .A2(n17732), .ZN(n12724) );
  OR2_X1 U14370 ( .A1(n17735), .A2(n12724), .ZN(n19377) );
  INV_X1 U14371 ( .A(n17734), .ZN(n12725) );
  NOR3_X1 U14372 ( .A1(n19377), .A2(n12726), .A3(n12725), .ZN(n12727) );
  NOR2_X1 U14373 ( .A1(n12727), .A2(n17851), .ZN(n17724) );
  INV_X1 U14374 ( .A(n17724), .ZN(n12728) );
  OAI211_X1 U14375 ( .C1(n17707), .C2(n17851), .A(n12728), .B(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17698) );
  NAND2_X1 U14376 ( .A1(n12729), .A2(n17698), .ZN(n17687) );
  NAND2_X1 U14377 ( .A1(n12730), .A2(n17687), .ZN(n17663) );
  AOI21_X1 U14378 ( .B1(n12731), .B2(n19378), .A(n17663), .ZN(n12799) );
  NOR2_X1 U14379 ( .A1(n12799), .A2(n12732), .ZN(n12733) );
  NOR2_X1 U14380 ( .A1(n12734), .A2(n12733), .ZN(n12735) );
  NAND2_X1 U14381 ( .A1(n16643), .A2(n12737), .ZN(n12743) );
  NAND2_X1 U14382 ( .A1(n12738), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12740) );
  AOI22_X1 U14383 ( .A1(n11791), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12739) );
  OAI211_X1 U14384 ( .C1(n12741), .C2(n19339), .A(n12740), .B(n12739), .ZN(
        n12742) );
  AOI21_X1 U14385 ( .B1(n15115), .B2(n12188), .A(n11164), .ZN(n12745) );
  NAND2_X1 U14386 ( .A1(n19350), .A2(n19398), .ZN(n12747) );
  OAI21_X1 U14387 ( .B1(n16405), .B2(n19388), .A(n12749), .ZN(P2_U3015) );
  INV_X1 U14388 ( .A(n17591), .ZN(n12752) );
  INV_X1 U14389 ( .A(n12753), .ZN(n17581) );
  INV_X1 U14390 ( .A(n17561), .ZN(n12756) );
  NAND2_X1 U14391 ( .A1(n12759), .A2(n12758), .ZN(n12760) );
  XNOR2_X1 U14392 ( .A(n12761), .B(n12760), .ZN(n12778) );
  NAND2_X1 U14393 ( .A1(n15153), .A2(n17965), .ZN(n12762) );
  NAND2_X1 U14394 ( .A1(n12763), .A2(n12762), .ZN(n15169) );
  NAND2_X1 U14395 ( .A1(n15169), .A2(n19078), .ZN(n19451) );
  OR2_X1 U14396 ( .A1(n19451), .A2(n12188), .ZN(n18106) );
  NAND2_X1 U14397 ( .A1(n12778), .A2(n18079), .ZN(n12777) );
  NAND2_X1 U14398 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12765) );
  NAND2_X1 U14399 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n18114) );
  NAND2_X1 U14400 ( .A1(n20083), .A2(n18114), .ZN(n19077) );
  OR2_X1 U14401 ( .A1(n19077), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12766) );
  INV_X1 U14402 ( .A(n14704), .ZN(n15178) );
  NAND2_X1 U14403 ( .A1(n22310), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12767) );
  NAND2_X1 U14404 ( .A1(n15178), .A2(n12767), .ZN(n16341) );
  INV_X2 U14405 ( .A(n19380), .ZN(n19407) );
  NAND2_X1 U14406 ( .A1(n19407), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12783) );
  OAI21_X1 U14407 ( .B1(n18076), .B2(n12768), .A(n12783), .ZN(n12773) );
  NOR2_X1 U14408 ( .A1(n12769), .A2(n12770), .ZN(n12771) );
  OR2_X1 U14409 ( .A1(n17350), .A2(n12771), .ZN(n17421) );
  AND2_X1 U14410 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n17961) );
  NOR2_X1 U14411 ( .A1(n17421), .A2(n18105), .ZN(n12772) );
  AOI211_X1 U14412 ( .C1(n18070), .C2(n14091), .A(n12773), .B(n12772), .ZN(
        n12774) );
  INV_X1 U14413 ( .A(n12775), .ZN(n12776) );
  NAND2_X1 U14414 ( .A1(n12777), .A2(n12776), .ZN(P2_U2993) );
  NAND2_X1 U14415 ( .A1(n12778), .A2(n19419), .ZN(n12791) );
  INV_X1 U14416 ( .A(n17793), .ZN(n17816) );
  NAND2_X1 U14417 ( .A1(n17816), .A2(n17738), .ZN(n17757) );
  OR2_X1 U14418 ( .A1(n17757), .A2(n12779), .ZN(n17748) );
  OAI21_X1 U14419 ( .B1(n17748), .B2(n17550), .A(n12780), .ZN(n12786) );
  OR2_X1 U14420 ( .A1(n17740), .A2(n12781), .ZN(n12782) );
  NAND2_X1 U14421 ( .A1(n12782), .A2(n17352), .ZN(n17476) );
  OAI21_X1 U14422 ( .B1(n17928), .B2(n17476), .A(n12783), .ZN(n12785) );
  NOR2_X1 U14423 ( .A1(n17421), .A2(n19416), .ZN(n12784) );
  AOI211_X1 U14424 ( .C1(n17724), .C2(n12786), .A(n12785), .B(n12784), .ZN(
        n12787) );
  INV_X1 U14425 ( .A(n12789), .ZN(n12790) );
  NAND2_X1 U14426 ( .A1(n12791), .A2(n12790), .ZN(P2_U3025) );
  NAND2_X1 U14427 ( .A1(n12792), .A2(n16695), .ZN(n12797) );
  INV_X1 U14428 ( .A(n12793), .ZN(n12794) );
  NOR2_X1 U14429 ( .A1(n12795), .A2(n12794), .ZN(n12796) );
  XNOR2_X1 U14430 ( .A(n12797), .B(n12796), .ZN(n16413) );
  NAND3_X1 U14431 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12798) );
  OAI21_X1 U14432 ( .B1(n14052), .B2(n12798), .A(n12804), .ZN(n12803) );
  INV_X1 U14433 ( .A(n12799), .ZN(n12802) );
  NOR2_X1 U14434 ( .A1(n12800), .A2(n17928), .ZN(n12801) );
  NOR2_X1 U14435 ( .A1(n19380), .A2(n18204), .ZN(n16408) );
  INV_X1 U14436 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17494) );
  NAND3_X1 U14437 ( .A1(n17493), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16702) );
  AOI21_X2 U14438 ( .B1(n16702), .B2(n12804), .A(n11528), .ZN(n16411) );
  NAND2_X1 U14439 ( .A1(n16411), .A2(n19420), .ZN(n12806) );
  OAI21_X1 U14440 ( .B1(n16413), .B2(n19388), .A(n12808), .ZN(P2_U3016) );
  AND2_X2 U14441 ( .A1(n12819), .A2(n12817), .ZN(n13115) );
  AOI22_X1 U14442 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11178), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12814) );
  AOI22_X1 U14443 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12860), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12813) );
  AOI22_X1 U14444 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11189), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12812) );
  AOI22_X1 U14445 ( .A1(n12830), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12811) );
  NAND4_X1 U14446 ( .A1(n12814), .A2(n12813), .A3(n12812), .A4(n12811), .ZN(
        n12825) );
  AOI22_X1 U14447 ( .A1(n12847), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13453), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12823) );
  AOI22_X1 U14448 ( .A1(n13441), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12969), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12822) );
  AND2_X2 U14449 ( .A1(n12817), .A2(n14746), .ZN(n12984) );
  AOI22_X1 U14450 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12821) );
  AND2_X2 U14451 ( .A1(n14508), .A2(n14746), .ZN(n12990) );
  AOI22_X1 U14452 ( .A1(n12989), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12990), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12820) );
  NAND4_X1 U14453 ( .A1(n12823), .A2(n12822), .A3(n12821), .A4(n12820), .ZN(
        n12824) );
  OR2_X2 U14454 ( .A1(n12825), .A2(n12824), .ZN(n12941) );
  AOI22_X1 U14455 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13453), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12829) );
  AOI22_X1 U14456 ( .A1(n13560), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12828) );
  AOI22_X1 U14457 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12969), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12827) );
  AOI22_X1 U14458 ( .A1(n12847), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12826) );
  AOI22_X1 U14459 ( .A1(n12989), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12860), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12833) );
  AOI22_X1 U14460 ( .A1(n11178), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13441), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12832) );
  AOI22_X1 U14461 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12990), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12831) );
  INV_X1 U14462 ( .A(n12870), .ZN(n12859) );
  AOI22_X1 U14463 ( .A1(n12860), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11189), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12839) );
  AOI22_X1 U14464 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12983), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12838) );
  AOI22_X1 U14465 ( .A1(n12989), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12990), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12837) );
  NAND4_X1 U14466 ( .A1(n12840), .A2(n12839), .A3(n12838), .A4(n12837), .ZN(
        n12841) );
  INV_X1 U14467 ( .A(n12841), .ZN(n12846) );
  AOI22_X1 U14468 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12845) );
  AOI22_X1 U14469 ( .A1(n12830), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13453), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12844) );
  AOI22_X1 U14470 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12969), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12843) );
  AOI22_X1 U14471 ( .A1(n13441), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12842) );
  AOI22_X1 U14472 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11189), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12851) );
  AOI22_X1 U14473 ( .A1(n12830), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12850) );
  AOI22_X1 U14474 ( .A1(n12860), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13453), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12849) );
  AOI22_X1 U14475 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11179), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12848) );
  AOI22_X1 U14476 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13441), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12855) );
  AOI22_X1 U14477 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12969), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12854) );
  AOI22_X1 U14478 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12853) );
  AOI22_X1 U14479 ( .A1(n12989), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12990), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12852) );
  AND2_X4 U14480 ( .A1(n12856), .A2(n12857), .ZN(n12933) );
  INV_X1 U14481 ( .A(n12909), .ZN(n12858) );
  NAND2_X1 U14482 ( .A1(n12859), .A2(n12858), .ZN(n12911) );
  AOI22_X1 U14483 ( .A1(n12830), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12864) );
  AOI22_X1 U14484 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12847), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12863) );
  AOI22_X1 U14485 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12862) );
  AOI22_X1 U14486 ( .A1(n12860), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13453), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12861) );
  AOI22_X1 U14487 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12969), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12868) );
  AOI22_X1 U14488 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13441), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12867) );
  AOI22_X1 U14489 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12866) );
  AOI22_X1 U14490 ( .A1(n12989), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12990), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12865) );
  NAND2_X2 U14491 ( .A1(n12869), .A2(n11539), .ZN(n14797) );
  NAND2_X1 U14492 ( .A1(n12911), .A2(n14797), .ZN(n12884) );
  NAND2_X1 U14493 ( .A1(n12948), .A2(n12870), .ZN(n12882) );
  AOI22_X1 U14494 ( .A1(n12830), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12860), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12874) );
  AOI22_X1 U14495 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11177), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12873) );
  AOI22_X1 U14496 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13441), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12872) );
  AOI22_X1 U14497 ( .A1(n12847), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12990), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12871) );
  AOI22_X1 U14498 ( .A1(n13453), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13560), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12880) );
  AOI22_X1 U14499 ( .A1(n12989), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12876), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12879) );
  AOI22_X1 U14500 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12878) );
  AOI22_X1 U14501 ( .A1(n12969), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12984), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12877) );
  NAND2_X2 U14502 ( .A1(n11538), .A2(n11209), .ZN(n12886) );
  NAND3_X1 U14503 ( .A1(n14284), .A2(n13614), .A3(n12957), .ZN(n12881) );
  NAND2_X1 U14504 ( .A1(n14310), .A2(n12886), .ZN(n12885) );
  NAND2_X1 U14505 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12890) );
  NAND2_X1 U14506 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12889) );
  NAND2_X1 U14507 ( .A1(n12969), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12888) );
  NAND2_X1 U14508 ( .A1(n13441), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12887) );
  NAND4_X1 U14509 ( .A1(n12890), .A2(n12889), .A3(n12888), .A4(n12887), .ZN(
        n12894) );
  NAND2_X1 U14510 ( .A1(n12984), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12891) );
  NAND2_X1 U14511 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12892) );
  CLKBUF_X1 U14512 ( .A(n13244), .Z(n12895) );
  NAND2_X1 U14513 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12901) );
  NAND2_X1 U14514 ( .A1(n13560), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12900) );
  NAND2_X1 U14515 ( .A1(n12830), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12899) );
  NAND2_X1 U14516 ( .A1(n12968), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12898) );
  NAND2_X1 U14517 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12905) );
  NAND2_X1 U14518 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12904) );
  NAND2_X1 U14519 ( .A1(n12860), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12903) );
  NAND2_X1 U14520 ( .A1(n13453), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12902) );
  OAI21_X1 U14521 ( .B1(n13614), .B2(n12933), .A(n12941), .ZN(n12908) );
  INV_X1 U14522 ( .A(n12908), .ZN(n14289) );
  INV_X1 U14523 ( .A(n12961), .ZN(n12910) );
  NAND2_X1 U14524 ( .A1(n12910), .A2(n12909), .ZN(n12934) );
  NAND2_X1 U14525 ( .A1(n12934), .A2(n14462), .ZN(n12956) );
  NAND2_X1 U14526 ( .A1(n12876), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12915) );
  NAND2_X1 U14527 ( .A1(n11179), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12914) );
  NAND2_X1 U14528 ( .A1(n12860), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12913) );
  NAND2_X1 U14529 ( .A1(n13453), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12912) );
  NAND2_X1 U14530 ( .A1(n11191), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12919) );
  NAND2_X1 U14531 ( .A1(n11189), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12918) );
  NAND2_X1 U14532 ( .A1(n12830), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12917) );
  NAND2_X1 U14533 ( .A1(n12968), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12916) );
  NAND2_X1 U14534 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12924) );
  NAND2_X1 U14535 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12923) );
  NAND2_X1 U14536 ( .A1(n12969), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12922) );
  NAND2_X1 U14537 ( .A1(n13441), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12921) );
  NAND2_X1 U14538 ( .A1(n12989), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12928) );
  NAND2_X1 U14539 ( .A1(n12983), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12927) );
  NAND2_X1 U14540 ( .A1(n12984), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12926) );
  NAND2_X1 U14541 ( .A1(n12990), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12925) );
  NAND4_X4 U14542 ( .A1(n12932), .A2(n12931), .A3(n12930), .A4(n12929), .ZN(
        n12947) );
  NAND2_X2 U14543 ( .A1(n14797), .A2(n12947), .ZN(n16321) );
  NAND2_X1 U14544 ( .A1(n14319), .A2(n12947), .ZN(n15070) );
  AND2_X1 U14545 ( .A1(n12947), .A2(n13614), .ZN(n13617) );
  NAND2_X1 U14546 ( .A1(n13617), .A2(n12933), .ZN(n14287) );
  NAND2_X1 U14547 ( .A1(n12935), .A2(n12934), .ZN(n14291) );
  NAND3_X1 U14548 ( .A1(n12938), .A2(n12937), .A3(n14305), .ZN(n12951) );
  NOR2_X1 U14549 ( .A1(n11160), .A2(n14882), .ZN(n12939) );
  NAND2_X1 U14550 ( .A1(n22329), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n22323) );
  INV_X1 U14551 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n12943) );
  NAND2_X1 U14552 ( .A1(n12943), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n12944) );
  NAND2_X1 U14553 ( .A1(n22323), .A2(n12944), .ZN(n14278) );
  NOR2_X1 U14554 ( .A1(n12947), .A2(n14278), .ZN(n12950) );
  INV_X1 U14555 ( .A(n13614), .ZN(n12945) );
  NAND2_X1 U14557 ( .A1(n14421), .A2(n16724), .ZN(n13687) );
  NAND2_X1 U14558 ( .A1(n17940), .A2(n22287), .ZN(n14629) );
  XNOR2_X1 U14559 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n22404) );
  OR2_X1 U14560 ( .A1(n17985), .A2(n22406), .ZN(n13024) );
  OAI21_X1 U14561 ( .B1(n14629), .B2(n22404), .A(n13024), .ZN(n12952) );
  INV_X1 U14562 ( .A(n12952), .ZN(n12953) );
  MUX2_X1 U14563 ( .A(n14629), .B(n17985), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n13013) );
  AND2_X1 U14564 ( .A1(n12949), .A2(n16710), .ZN(n15607) );
  INV_X1 U14565 ( .A(n12946), .ZN(n12958) );
  OR2_X1 U14566 ( .A1(n12958), .A2(n12957), .ZN(n14306) );
  NAND2_X1 U14567 ( .A1(n17940), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20768) );
  AOI21_X1 U14568 ( .B1(n12886), .B2(n16710), .A(n20768), .ZN(n12959) );
  NAND3_X1 U14569 ( .A1(n14306), .A2(n12959), .A3(n15070), .ZN(n12960) );
  AOI21_X1 U14570 ( .B1(n15607), .B2(n12961), .A(n12960), .ZN(n12965) );
  NAND3_X1 U14571 ( .A1(n12909), .A2(n11359), .A3(n14797), .ZN(n12963) );
  NAND2_X1 U14572 ( .A1(n12962), .A2(n12963), .ZN(n12964) );
  OAI211_X1 U14573 ( .C1(n12956), .C2(n12949), .A(n12965), .B(n12964), .ZN(
        n13153) );
  NAND2_X1 U14574 ( .A1(n13155), .A2(n13153), .ZN(n12967) );
  INV_X1 U14575 ( .A(n12967), .ZN(n12966) );
  NAND2_X1 U14576 ( .A1(n22416), .A2(n12966), .ZN(n13028) );
  NAND2_X1 U14577 ( .A1(n11154), .A2(n12967), .ZN(n14824) );
  NAND2_X1 U14578 ( .A1(n14824), .A2(n13028), .ZN(n14461) );
  NAND2_X1 U14579 ( .A1(n14461), .A2(n22287), .ZN(n12982) );
  AOI22_X1 U14580 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13595), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12973) );
  AOI22_X1 U14581 ( .A1(n13583), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12972) );
  BUF_X1 U14582 ( .A(n12968), .Z(n13586) );
  AOI22_X1 U14583 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12971) );
  AOI22_X1 U14584 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12970) );
  NAND4_X1 U14585 ( .A1(n12973), .A2(n12972), .A3(n12971), .A4(n12970), .ZN(
        n12979) );
  INV_X1 U14586 ( .A(n12875), .ZN(n13479) );
  AOI22_X1 U14587 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12977) );
  AOI22_X1 U14588 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12976) );
  AOI22_X1 U14589 ( .A1(n11178), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13441), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12975) );
  AOI22_X1 U14590 ( .A1(n13594), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12974) );
  NAND4_X1 U14591 ( .A1(n12977), .A2(n12976), .A3(n12975), .A4(n12974), .ZN(
        n12978) );
  NAND2_X1 U14592 ( .A1(n14314), .A2(n14635), .ZN(n12980) );
  INV_X1 U14593 ( .A(n14635), .ZN(n12999) );
  NAND2_X1 U14594 ( .A1(n14319), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12998) );
  NOR2_X1 U14595 ( .A1(n14882), .A2(n22287), .ZN(n13014) );
  AOI22_X1 U14596 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13593), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12988) );
  AOI22_X1 U14597 ( .A1(n13583), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12987) );
  AOI22_X1 U14598 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12986) );
  AOI22_X1 U14599 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12985) );
  NAND4_X1 U14600 ( .A1(n12988), .A2(n12987), .A3(n12986), .A4(n12985), .ZN(
        n12996) );
  AOI22_X1 U14601 ( .A1(n11152), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13453), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12994) );
  AOI22_X1 U14602 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12993) );
  AOI22_X1 U14603 ( .A1(n13592), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12992) );
  AOI22_X1 U14604 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12991) );
  NAND4_X1 U14605 ( .A1(n12994), .A2(n12993), .A3(n12992), .A4(n12991), .ZN(
        n12995) );
  INV_X1 U14606 ( .A(n15606), .ZN(n13110) );
  NAND2_X1 U14607 ( .A1(n13014), .A2(n13110), .ZN(n13015) );
  AND3_X2 U14608 ( .A1(n16710), .A2(n14882), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n13637) );
  NAND2_X1 U14609 ( .A1(n13637), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12997) );
  OAI211_X1 U14610 ( .C1(n12999), .C2(n12998), .A(n13015), .B(n12997), .ZN(
        n13020) );
  AOI22_X1 U14611 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n13453), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13003) );
  AOI22_X1 U14612 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n12860), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13002) );
  AOI22_X1 U14613 ( .A1(n11178), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13001) );
  AOI22_X1 U14614 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13441), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13000) );
  NAND4_X1 U14615 ( .A1(n13003), .A2(n13002), .A3(n13001), .A4(n13000), .ZN(
        n13009) );
  AOI22_X1 U14616 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n13244), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13007) );
  AOI22_X1 U14617 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n13561), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13006) );
  AOI22_X1 U14618 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13005) );
  AOI22_X1 U14619 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13004) );
  NAND4_X1 U14620 ( .A1(n13007), .A2(n13006), .A3(n13005), .A4(n13004), .ZN(
        n13008) );
  INV_X1 U14621 ( .A(n14636), .ZN(n13012) );
  NAND2_X1 U14622 ( .A1(n13637), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13011) );
  AOI21_X1 U14623 ( .B1(n14314), .B2(n15606), .A(n22287), .ZN(n13010) );
  OAI211_X1 U14624 ( .C1(n13012), .C2(n16710), .A(n13011), .B(n13010), .ZN(
        n13163) );
  NAND2_X1 U14625 ( .A1(n13013), .A2(n22287), .ZN(n13017) );
  NAND2_X1 U14626 ( .A1(n13014), .A2(n15606), .ZN(n15603) );
  MUX2_X1 U14627 ( .A(n15603), .B(n13015), .S(n14636), .Z(n13016) );
  NAND2_X1 U14628 ( .A1(n13017), .A2(n13016), .ZN(n13161) );
  NAND2_X1 U14629 ( .A1(n13163), .A2(n13161), .ZN(n13018) );
  NAND2_X1 U14630 ( .A1(n13018), .A2(n15603), .ZN(n13147) );
  INV_X1 U14631 ( .A(n13019), .ZN(n13021) );
  NAND2_X1 U14632 ( .A1(n13021), .A2(n13020), .ZN(n13022) );
  INV_X1 U14633 ( .A(n13024), .ZN(n13026) );
  NAND2_X1 U14634 ( .A1(n13028), .A2(n13027), .ZN(n13039) );
  INV_X1 U14635 ( .A(n13039), .ZN(n13037) );
  NAND2_X1 U14636 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n13030) );
  NAND2_X1 U14637 ( .A1(n18000), .A2(n13030), .ZN(n13032) );
  NAND2_X1 U14638 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22441) );
  INV_X1 U14639 ( .A(n22441), .ZN(n13031) );
  NAND2_X1 U14640 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13031), .ZN(
        n13053) );
  NAND2_X1 U14641 ( .A1(n13032), .A2(n13053), .ZN(n15219) );
  OAI22_X1 U14642 ( .A1(n14629), .A2(n15219), .B1(n17985), .B2(n18000), .ZN(
        n13033) );
  INV_X1 U14643 ( .A(n13033), .ZN(n13034) );
  INV_X1 U14644 ( .A(n13038), .ZN(n13036) );
  NAND2_X1 U14645 ( .A1(n14882), .A2(n16710), .ZN(n13040) );
  AOI22_X1 U14646 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11188), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13045) );
  AOI22_X1 U14647 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13044) );
  AOI22_X1 U14648 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13043) );
  AOI22_X1 U14649 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13042) );
  NAND4_X1 U14650 ( .A1(n13045), .A2(n13044), .A3(n13043), .A4(n13042), .ZN(
        n13051) );
  AOI22_X1 U14651 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13049) );
  AOI22_X1 U14652 ( .A1(n11178), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13048) );
  AOI22_X1 U14653 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13441), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13047) );
  AOI22_X1 U14654 ( .A1(n13583), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13046) );
  NAND4_X1 U14655 ( .A1(n13049), .A2(n13048), .A3(n13047), .A4(n13046), .ZN(
        n13050) );
  OR2_X1 U14656 ( .A1(n13051), .A2(n13050), .ZN(n14694) );
  AOI22_X1 U14657 ( .A1(n13674), .A2(n14694), .B1(n13637), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13052) );
  OR2_X1 U14658 ( .A1(n13029), .A2(n11358), .ZN(n13058) );
  INV_X1 U14659 ( .A(n14629), .ZN(n13056) );
  INV_X1 U14660 ( .A(n13053), .ZN(n14782) );
  NAND2_X1 U14661 ( .A1(n14782), .A2(n15215), .ZN(n22735) );
  NAND2_X1 U14662 ( .A1(n13053), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13054) );
  NAND2_X1 U14663 ( .A1(n22735), .A2(n13054), .ZN(n15422) );
  INV_X1 U14664 ( .A(n17985), .ZN(n13055) );
  AOI22_X1 U14665 ( .A1(n13056), .A2(n15422), .B1(n13055), .B2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13057) );
  AOI22_X1 U14666 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13062) );
  AOI22_X1 U14667 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13061) );
  AOI22_X1 U14668 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13060) );
  AOI22_X1 U14669 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13059) );
  NAND4_X1 U14670 ( .A1(n13062), .A2(n13061), .A3(n13060), .A4(n13059), .ZN(
        n13068) );
  AOI22_X1 U14671 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13066) );
  AOI22_X1 U14672 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13441), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13065) );
  AOI22_X1 U14673 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13064) );
  AOI22_X1 U14674 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13063) );
  NAND4_X1 U14675 ( .A1(n13066), .A2(n13065), .A3(n13064), .A4(n13063), .ZN(
        n13067) );
  AOI22_X1 U14676 ( .A1(n13674), .A2(n15289), .B1(n13637), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13069) );
  AOI22_X1 U14677 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13073) );
  AOI22_X1 U14678 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13072) );
  AOI22_X1 U14679 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13071) );
  AOI22_X1 U14680 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13070) );
  NAND4_X1 U14681 ( .A1(n13073), .A2(n13072), .A3(n13071), .A4(n13070), .ZN(
        n13079) );
  AOI22_X1 U14682 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13077) );
  AOI22_X1 U14683 ( .A1(n11178), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13441), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13076) );
  AOI22_X1 U14684 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13075) );
  AOI22_X1 U14685 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13074) );
  NAND4_X1 U14686 ( .A1(n13077), .A2(n13076), .A3(n13075), .A4(n13074), .ZN(
        n13078) );
  NOR2_X1 U14687 ( .A1(n13079), .A2(n13078), .ZN(n15577) );
  NAND2_X1 U14688 ( .A1(n13637), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13080) );
  OAI21_X1 U14689 ( .B1(n13624), .B2(n15577), .A(n13080), .ZN(n13184) );
  AOI22_X1 U14690 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13595), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13086) );
  AOI22_X1 U14691 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13593), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13085) );
  AOI22_X1 U14692 ( .A1(n13583), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13084) );
  AOI22_X1 U14693 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13083) );
  NAND4_X1 U14694 ( .A1(n13086), .A2(n13085), .A3(n13084), .A4(n13083), .ZN(
        n13092) );
  AOI22_X1 U14695 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13090) );
  AOI22_X1 U14696 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13089) );
  AOI22_X1 U14697 ( .A1(n13586), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13088) );
  AOI22_X1 U14698 ( .A1(n13592), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13087) );
  NAND4_X1 U14699 ( .A1(n13090), .A2(n13089), .A3(n13088), .A4(n13087), .ZN(
        n13091) );
  INV_X1 U14700 ( .A(n15587), .ZN(n13094) );
  NAND2_X1 U14701 ( .A1(n13637), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n13093) );
  OAI21_X1 U14702 ( .B1(n13624), .B2(n13094), .A(n13093), .ZN(n13194) );
  AOI22_X1 U14703 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13098) );
  AOI22_X1 U14704 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13097) );
  AOI22_X1 U14705 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13096) );
  AOI22_X1 U14706 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13095) );
  NAND4_X1 U14707 ( .A1(n13098), .A2(n13097), .A3(n13096), .A4(n13095), .ZN(
        n13104) );
  AOI22_X1 U14708 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13102) );
  AOI22_X1 U14709 ( .A1(n11177), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13441), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13101) );
  AOI22_X1 U14710 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13100) );
  AOI22_X1 U14711 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13099) );
  NAND4_X1 U14712 ( .A1(n13102), .A2(n13101), .A3(n13100), .A4(n13099), .ZN(
        n13103) );
  NOR2_X1 U14713 ( .A1(n13104), .A2(n13103), .ZN(n15589) );
  OR2_X1 U14714 ( .A1(n13624), .A2(n15589), .ZN(n13106) );
  NAND2_X1 U14715 ( .A1(n13637), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n13105) );
  NAND2_X1 U14716 ( .A1(n13637), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13109) );
  OAI21_X1 U14717 ( .B1(n13624), .B2(n13110), .A(n13109), .ZN(n13111) );
  NOR2_X2 U14718 ( .A1(n12957), .A2(n22424), .ZN(n13299) );
  INV_X1 U14719 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n15314) );
  NOR2_X2 U14720 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13582) );
  OAI21_X1 U14721 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n13112), .A(
        n13140), .ZN(n22142) );
  AOI22_X1 U14722 ( .A1(n13582), .A2(n22142), .B1(n13611), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13113) );
  OAI21_X1 U14723 ( .B1(n13149), .B2(n15314), .A(n13113), .ZN(n13114) );
  AOI21_X1 U14724 ( .B1(n15593), .B2(n13299), .A(n13114), .ZN(n15312) );
  XOR2_X1 U14725 ( .A(n15457), .B(n13222), .Z(n15466) );
  INV_X1 U14726 ( .A(n15466), .ZN(n16094) );
  AOI22_X1 U14727 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13119) );
  AOI22_X1 U14728 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13118) );
  AOI22_X1 U14729 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13117) );
  AOI22_X1 U14730 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13116) );
  NAND4_X1 U14731 ( .A1(n13119), .A2(n13118), .A3(n13117), .A4(n13116), .ZN(
        n13125) );
  AOI22_X1 U14732 ( .A1(n13479), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13123) );
  AOI22_X1 U14733 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U14734 ( .A1(n11178), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13441), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13121) );
  AOI22_X1 U14735 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13120) );
  NAND4_X1 U14736 ( .A1(n13123), .A2(n13122), .A3(n13121), .A4(n13120), .ZN(
        n13124) );
  OAI21_X1 U14737 ( .B1(n13125), .B2(n13124), .A(n13299), .ZN(n13128) );
  NAND2_X1 U14738 ( .A1(n13612), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n13127) );
  NAND2_X1 U14739 ( .A1(n13611), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13126) );
  NAND3_X1 U14740 ( .A1(n13128), .A2(n13127), .A3(n13126), .ZN(n13129) );
  AOI21_X1 U14741 ( .B1(n16094), .B2(n13582), .A(n13129), .ZN(n15454) );
  AOI22_X1 U14742 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n13479), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13133) );
  AOI22_X1 U14743 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n13561), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13132) );
  AOI22_X1 U14744 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n13593), .B1(
        n13441), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13131) );
  AOI22_X1 U14745 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13130) );
  NAND4_X1 U14746 ( .A1(n13133), .A2(n13132), .A3(n13131), .A4(n13130), .ZN(
        n13139) );
  AOI22_X1 U14747 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n11188), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13137) );
  AOI22_X1 U14748 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13136) );
  AOI22_X1 U14749 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13135) );
  AOI22_X1 U14750 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13134) );
  NAND4_X1 U14751 ( .A1(n13137), .A2(n13136), .A3(n13135), .A4(n13134), .ZN(
        n13138) );
  OAI21_X1 U14752 ( .B1(n13139), .B2(n13138), .A(n13299), .ZN(n13144) );
  INV_X1 U14753 ( .A(n13140), .ZN(n13141) );
  XNOR2_X1 U14754 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n13141), .ZN(
        n15615) );
  AOI22_X1 U14755 ( .A1(n13582), .A2(n15615), .B1(n13611), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13143) );
  NAND2_X1 U14756 ( .A1(n13612), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n13142) );
  NAND2_X1 U14757 ( .A1(n13145), .A2(n11530), .ZN(n13211) );
  NAND2_X1 U14758 ( .A1(n14759), .A2(n13299), .ZN(n14625) );
  INV_X1 U14759 ( .A(n13149), .ZN(n13612) );
  AOI22_X1 U14760 ( .A1(n13612), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n22424), .ZN(n13151) );
  INV_X1 U14761 ( .A(n12948), .ZN(n13705) );
  NAND2_X1 U14762 ( .A1(n13705), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13181) );
  INV_X1 U14763 ( .A(n13181), .ZN(n13186) );
  NAND2_X1 U14764 ( .A1(n13186), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13150) );
  AND2_X1 U14765 ( .A1(n13151), .A2(n13150), .ZN(n14624) );
  NAND2_X1 U14766 ( .A1(n13611), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13152) );
  AND2_X1 U14767 ( .A1(n14624), .A2(n13152), .ZN(n13165) );
  INV_X1 U14768 ( .A(n13152), .ZN(n14672) );
  INV_X1 U14769 ( .A(n13153), .ZN(n13154) );
  XNOR2_X1 U14770 ( .A(n13155), .B(n13154), .ZN(n22417) );
  NAND2_X1 U14771 ( .A1(n22417), .A2(n13299), .ZN(n13160) );
  AOI22_X1 U14772 ( .A1(n13156), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n22424), .ZN(n13158) );
  NAND2_X1 U14773 ( .A1(n13186), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13157) );
  AND2_X1 U14774 ( .A1(n13158), .A2(n13157), .ZN(n13159) );
  NAND2_X1 U14775 ( .A1(n13160), .A2(n13159), .ZN(n14365) );
  INV_X1 U14776 ( .A(n13161), .ZN(n13162) );
  XNOR2_X1 U14777 ( .A(n13163), .B(n13162), .ZN(n22280) );
  INV_X1 U14778 ( .A(n22280), .ZN(n14826) );
  AOI21_X1 U14779 ( .B1(n14826), .B2(n12933), .A(n22424), .ZN(n14364) );
  NAND2_X1 U14780 ( .A1(n14365), .A2(n14364), .ZN(n14363) );
  OR2_X1 U14781 ( .A1(n14365), .A2(n13557), .ZN(n13164) );
  NAND2_X1 U14782 ( .A1(n14363), .A2(n13164), .ZN(n14626) );
  NAND2_X1 U14783 ( .A1(n11194), .A2(n13299), .ZN(n14674) );
  XNOR2_X1 U14784 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15101) );
  AOI21_X1 U14785 ( .B1(n13582), .B2(n15101), .A(n13611), .ZN(n13170) );
  NAND2_X1 U14786 ( .A1(n13612), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n13169) );
  OAI211_X1 U14787 ( .C1(n13181), .C2(n12809), .A(n13170), .B(n13169), .ZN(
        n13171) );
  INV_X1 U14788 ( .A(n13171), .ZN(n14671) );
  NAND2_X1 U14789 ( .A1(n14674), .A2(n14671), .ZN(n13172) );
  NAND2_X1 U14790 ( .A1(n13176), .A2(n14761), .ZN(n13177) );
  INV_X1 U14791 ( .A(n13299), .ZN(n13289) );
  AOI21_X1 U14792 ( .B1(n14946), .B2(n13178), .A(n13188), .ZN(n22097) );
  INV_X1 U14793 ( .A(n13611), .ZN(n13228) );
  OAI22_X1 U14794 ( .A1(n22097), .A2(n13557), .B1(n13228), .B2(n14946), .ZN(
        n13179) );
  AOI21_X1 U14795 ( .B1(n13612), .B2(P1_EAX_REG_3__SCAN_IN), .A(n13179), .ZN(
        n13180) );
  OAI21_X1 U14796 ( .B1(n11358), .B2(n13181), .A(n13180), .ZN(n13182) );
  INV_X1 U14797 ( .A(n13182), .ZN(n13183) );
  NAND2_X1 U14798 ( .A1(n14867), .A2(n14868), .ZN(n14815) );
  NAND2_X1 U14799 ( .A1(n13186), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13191) );
  INV_X1 U14800 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n22110) );
  AOI21_X1 U14801 ( .B1(n22110), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13187) );
  AOI21_X1 U14802 ( .B1(n13612), .B2(P1_EAX_REG_4__SCAN_IN), .A(n13187), .ZN(
        n13190) );
  OAI21_X1 U14803 ( .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13188), .A(
        n13196), .ZN(n22118) );
  NOR2_X1 U14804 ( .A1(n22118), .A2(n13557), .ZN(n13189) );
  AOI21_X1 U14805 ( .B1(n13191), .B2(n13190), .A(n13189), .ZN(n13192) );
  AOI21_X1 U14806 ( .B1(n15288), .B2(n13299), .A(n13192), .ZN(n14816) );
  INV_X1 U14807 ( .A(n13193), .ZN(n13195) );
  NAND2_X1 U14808 ( .A1(n15576), .A2(n13299), .ZN(n13202) );
  INV_X1 U14809 ( .A(n13196), .ZN(n13198) );
  INV_X1 U14810 ( .A(n13206), .ZN(n13197) );
  OAI21_X1 U14811 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n13198), .A(
        n13197), .ZN(n22129) );
  NAND2_X1 U14812 ( .A1(n22129), .A2(n13582), .ZN(n13199) );
  OAI21_X1 U14813 ( .B1(n22119), .B2(n13228), .A(n13199), .ZN(n13200) );
  AOI21_X1 U14814 ( .B1(n13612), .B2(P1_EAX_REG_5__SCAN_IN), .A(n13200), .ZN(
        n13201) );
  NAND2_X1 U14815 ( .A1(n13202), .A2(n13201), .ZN(n14982) );
  NAND2_X1 U14816 ( .A1(n14814), .A2(n14982), .ZN(n14980) );
  INV_X1 U14817 ( .A(n14980), .ZN(n13210) );
  NAND2_X1 U14818 ( .A1(n13204), .A2(n13203), .ZN(n15585) );
  INV_X1 U14819 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n15284) );
  OAI21_X1 U14820 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13206), .A(
        n13205), .ZN(n22141) );
  AOI22_X1 U14821 ( .A1(n13582), .A2(n22141), .B1(n13611), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13207) );
  OAI21_X1 U14822 ( .B1(n13149), .B2(n15284), .A(n13207), .ZN(n13208) );
  INV_X1 U14823 ( .A(n15281), .ZN(n13209) );
  NAND2_X1 U14824 ( .A1(n13210), .A2(n13209), .ZN(n15311) );
  AOI22_X1 U14825 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11178), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13215) );
  AOI22_X1 U14826 ( .A1(n13479), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13214) );
  AOI22_X1 U14827 ( .A1(n12895), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13213) );
  AOI22_X1 U14828 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13441), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13212) );
  NAND4_X1 U14829 ( .A1(n13215), .A2(n13214), .A3(n13213), .A4(n13212), .ZN(
        n13221) );
  AOI22_X1 U14830 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13219) );
  AOI22_X1 U14831 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13218) );
  AOI22_X1 U14832 ( .A1(n13591), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13217) );
  AOI22_X1 U14833 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13216) );
  NAND4_X1 U14834 ( .A1(n13219), .A2(n13218), .A3(n13217), .A4(n13216), .ZN(
        n13220) );
  NOR2_X1 U14835 ( .A1(n13221), .A2(n13220), .ZN(n13225) );
  XNOR2_X1 U14836 ( .A(n13226), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17071) );
  NAND2_X1 U14837 ( .A1(n17071), .A2(n13582), .ZN(n13224) );
  AOI22_X1 U14838 ( .A1(n13156), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n13611), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13223) );
  OAI211_X1 U14839 ( .C1(n13225), .C2(n13289), .A(n13224), .B(n13223), .ZN(
        n15327) );
  NAND2_X1 U14840 ( .A1(n15325), .A2(n15327), .ZN(n15326) );
  OAI21_X1 U14841 ( .B1(n13227), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n13286), .ZN(n22167) );
  INV_X1 U14842 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n16041) );
  INV_X1 U14843 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n22159) );
  OAI22_X1 U14844 ( .A1(n13149), .A2(n16041), .B1(n13228), .B2(n22159), .ZN(
        n13229) );
  AOI21_X1 U14845 ( .B1(n22167), .B2(n13582), .A(n13229), .ZN(n15620) );
  AOI22_X1 U14846 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13595), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13234) );
  AOI22_X1 U14847 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13233) );
  AOI22_X1 U14848 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13232) );
  AOI22_X1 U14849 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13231) );
  NAND4_X1 U14850 ( .A1(n13234), .A2(n13233), .A3(n13232), .A4(n13231), .ZN(
        n13240) );
  AOI22_X1 U14851 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13238) );
  AOI22_X1 U14852 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13237) );
  AOI22_X1 U14853 ( .A1(n13592), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13236) );
  AOI22_X1 U14854 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13235) );
  NAND4_X1 U14855 ( .A1(n13238), .A2(n13237), .A3(n13236), .A4(n13235), .ZN(
        n13239) );
  OR2_X1 U14856 ( .A1(n13240), .A2(n13239), .ZN(n13241) );
  NAND2_X1 U14857 ( .A1(n13299), .A2(n13241), .ZN(n16040) );
  INV_X1 U14858 ( .A(n16040), .ZN(n13242) );
  INV_X1 U14859 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n22175) );
  OR2_X1 U14860 ( .A1(n13286), .A2(n22175), .ZN(n13243) );
  INV_X1 U14861 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16012) );
  XNOR2_X1 U14862 ( .A(n13243), .B(n16012), .ZN(n17049) );
  NAND2_X1 U14863 ( .A1(n17049), .A2(n13582), .ZN(n13259) );
  AOI22_X1 U14864 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11188), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13248) );
  AOI22_X1 U14865 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13247) );
  AOI22_X1 U14866 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13246) );
  AOI22_X1 U14867 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13245) );
  NAND4_X1 U14868 ( .A1(n13248), .A2(n13247), .A3(n13246), .A4(n13245), .ZN(
        n13254) );
  AOI22_X1 U14869 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13252) );
  AOI22_X1 U14870 ( .A1(n11177), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13441), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13251) );
  AOI22_X1 U14871 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13250) );
  AOI22_X1 U14872 ( .A1(n13583), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13249) );
  NAND4_X1 U14873 ( .A1(n13252), .A2(n13251), .A3(n13250), .A4(n13249), .ZN(
        n13253) );
  OAI21_X1 U14874 ( .B1(n13254), .B2(n13253), .A(n13299), .ZN(n13257) );
  NAND2_X1 U14875 ( .A1(n13612), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n13256) );
  NAND2_X1 U14876 ( .A1(n13611), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13255) );
  AND3_X1 U14877 ( .A1(n13257), .A2(n13256), .A3(n13255), .ZN(n13258) );
  NAND2_X1 U14878 ( .A1(n13259), .A2(n13258), .ZN(n16000) );
  XNOR2_X1 U14879 ( .A(n13286), .B(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n22169) );
  OR2_X1 U14880 ( .A1(n22169), .A2(n13557), .ZN(n13274) );
  AOI22_X1 U14881 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13263) );
  AOI22_X1 U14882 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13262) );
  AOI22_X1 U14883 ( .A1(n13592), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13261) );
  AOI22_X1 U14884 ( .A1(n13583), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13260) );
  NAND4_X1 U14885 ( .A1(n13263), .A2(n13262), .A3(n13261), .A4(n13260), .ZN(
        n13269) );
  AOI22_X1 U14886 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11178), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13267) );
  AOI22_X1 U14887 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11188), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13266) );
  AOI22_X1 U14888 ( .A1(n13244), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13265) );
  AOI22_X1 U14889 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13264) );
  NAND4_X1 U14890 ( .A1(n13267), .A2(n13266), .A3(n13265), .A4(n13264), .ZN(
        n13268) );
  OAI21_X1 U14891 ( .B1(n13269), .B2(n13268), .A(n13299), .ZN(n13272) );
  NAND2_X1 U14892 ( .A1(n13612), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n13271) );
  NAND2_X1 U14893 ( .A1(n13611), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13270) );
  AND3_X1 U14894 ( .A1(n13272), .A2(n13271), .A3(n13270), .ZN(n13273) );
  NAND2_X1 U14895 ( .A1(n13274), .A2(n13273), .ZN(n15622) );
  AOI22_X1 U14896 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13278) );
  AOI22_X1 U14897 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13277) );
  AOI22_X1 U14898 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13276) );
  AOI22_X1 U14899 ( .A1(n13594), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13275) );
  NAND4_X1 U14900 ( .A1(n13278), .A2(n13277), .A3(n13276), .A4(n13275), .ZN(
        n13284) );
  AOI22_X1 U14901 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13595), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13282) );
  AOI22_X1 U14902 ( .A1(n12895), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13281) );
  AOI22_X1 U14903 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13280) );
  AOI22_X1 U14904 ( .A1(n11178), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13441), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13279) );
  NAND4_X1 U14905 ( .A1(n13282), .A2(n13281), .A3(n13280), .A4(n13279), .ZN(
        n13283) );
  NOR2_X1 U14906 ( .A1(n13284), .A2(n13283), .ZN(n13290) );
  NAND2_X1 U14907 ( .A1(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n13285) );
  XNOR2_X1 U14908 ( .A(n13302), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17034) );
  NAND2_X1 U14909 ( .A1(n17034), .A2(n13582), .ZN(n13288) );
  AOI22_X1 U14910 ( .A1(n13156), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n13611), 
        .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n13287) );
  OAI211_X1 U14911 ( .C1(n13290), .C2(n13289), .A(n13288), .B(n13287), .ZN(
        n15531) );
  AOI22_X1 U14912 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13294) );
  AOI22_X1 U14913 ( .A1(n12895), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13293) );
  AOI22_X1 U14914 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13292) );
  AOI22_X1 U14915 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13291) );
  NAND4_X1 U14916 ( .A1(n13294), .A2(n13293), .A3(n13292), .A4(n13291), .ZN(
        n13301) );
  AOI22_X1 U14917 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11188), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13298) );
  AOI22_X1 U14918 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13297) );
  AOI22_X1 U14919 ( .A1(n11178), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13441), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13296) );
  AOI22_X1 U14920 ( .A1(n13594), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13295) );
  NAND4_X1 U14921 ( .A1(n13298), .A2(n13297), .A3(n13296), .A4(n13295), .ZN(
        n13300) );
  OAI21_X1 U14922 ( .B1(n13301), .B2(n13300), .A(n13299), .ZN(n13306) );
  NAND2_X1 U14923 ( .A1(n13156), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n13305) );
  INV_X1 U14924 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n22184) );
  XOR2_X1 U14925 ( .A(n22184), .B(n13321), .Z(n22187) );
  INV_X1 U14926 ( .A(n22187), .ZN(n13303) );
  AOI22_X1 U14927 ( .A1(n13611), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n13582), .B2(n13303), .ZN(n13304) );
  INV_X1 U14928 ( .A(n14462), .ZN(n14481) );
  AOI22_X1 U14929 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13595), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13310) );
  AOI22_X1 U14930 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n11188), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13309) );
  AOI22_X1 U14931 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n13586), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13308) );
  AOI22_X1 U14932 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n13592), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13307) );
  NAND4_X1 U14933 ( .A1(n13310), .A2(n13309), .A3(n13308), .A4(n13307), .ZN(
        n13316) );
  AOI22_X1 U14934 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n12895), .B1(
        n13561), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13314) );
  AOI22_X1 U14935 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n13453), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13313) );
  AOI22_X1 U14936 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13312) );
  AOI22_X1 U14937 ( .A1(n11178), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13311) );
  NAND4_X1 U14938 ( .A1(n13314), .A2(n13313), .A3(n13312), .A4(n13311), .ZN(
        n13315) );
  NOR2_X1 U14939 ( .A1(n13316), .A2(n13315), .ZN(n13320) );
  NAND2_X1 U14940 ( .A1(n22424), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13317) );
  NAND2_X1 U14941 ( .A1(n13557), .A2(n13317), .ZN(n13318) );
  AOI21_X1 U14942 ( .B1(n13156), .B2(P1_EAX_REG_16__SCAN_IN), .A(n13318), .ZN(
        n13319) );
  OAI21_X1 U14943 ( .B1(n13607), .B2(n13320), .A(n13319), .ZN(n13324) );
  INV_X1 U14944 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17017) );
  XNOR2_X1 U14945 ( .A(n13326), .B(n17017), .ZN(n22197) );
  NAND2_X1 U14946 ( .A1(n22197), .A2(n13582), .ZN(n13323) );
  NAND2_X1 U14947 ( .A1(n13324), .A2(n13323), .ZN(n16144) );
  NAND2_X1 U14948 ( .A1(n16051), .A2(n13325), .ZN(n16146) );
  INV_X1 U14949 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n22212) );
  XOR2_X1 U14950 ( .A(n22212), .B(n13340), .Z(n22215) );
  AOI22_X1 U14951 ( .A1(n13156), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n13611), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13338) );
  AOI22_X1 U14952 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13593), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13330) );
  AOI22_X1 U14953 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13329) );
  AOI22_X1 U14954 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13328) );
  AOI22_X1 U14955 ( .A1(n13594), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13327) );
  NAND4_X1 U14956 ( .A1(n13330), .A2(n13329), .A3(n13328), .A4(n13327), .ZN(
        n13336) );
  AOI22_X1 U14957 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13595), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13334) );
  AOI22_X1 U14958 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13333) );
  AOI22_X1 U14959 ( .A1(n12895), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13332) );
  AOI22_X1 U14960 ( .A1(n13592), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13331) );
  NAND4_X1 U14961 ( .A1(n13334), .A2(n13333), .A3(n13332), .A4(n13331), .ZN(
        n13335) );
  OAI21_X1 U14962 ( .B1(n13336), .B2(n13335), .A(n13573), .ZN(n13337) );
  OAI211_X1 U14963 ( .C1(n22215), .C2(n13557), .A(n13338), .B(n13337), .ZN(
        n16889) );
  NOR2_X2 U14964 ( .A1(n16146), .A2(n13339), .ZN(n16833) );
  XNOR2_X1 U14965 ( .A(n13356), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n22222) );
  NAND2_X1 U14966 ( .A1(n22222), .A2(n13582), .ZN(n13355) );
  AOI22_X1 U14967 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11177), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13344) );
  AOI22_X1 U14968 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13595), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13343) );
  AOI22_X1 U14969 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13342) );
  AOI22_X1 U14970 ( .A1(n12895), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13341) );
  NAND4_X1 U14971 ( .A1(n13344), .A2(n13343), .A3(n13342), .A4(n13341), .ZN(
        n13350) );
  AOI22_X1 U14972 ( .A1(n13583), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13348) );
  AOI22_X1 U14973 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13347) );
  AOI22_X1 U14974 ( .A1(n13592), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13346) );
  AOI22_X1 U14975 ( .A1(n13594), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13345) );
  NAND4_X1 U14976 ( .A1(n13348), .A2(n13347), .A3(n13346), .A4(n13345), .ZN(
        n13349) );
  NOR2_X1 U14977 ( .A1(n13350), .A2(n13349), .ZN(n13352) );
  AOI22_X1 U14978 ( .A1(n13156), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n22424), .ZN(n13351) );
  OAI21_X1 U14979 ( .B1(n13607), .B2(n13352), .A(n13351), .ZN(n13353) );
  NAND2_X1 U14980 ( .A1(n13353), .A2(n13557), .ZN(n13354) );
  NAND2_X1 U14981 ( .A1(n13355), .A2(n13354), .ZN(n16835) );
  OAI21_X1 U14982 ( .B1(n13357), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n13389), .ZN(n17000) );
  OR2_X1 U14983 ( .A1(n17000), .A2(n13557), .ZN(n13372) );
  AOI22_X1 U14984 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13361) );
  AOI22_X1 U14985 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13360) );
  AOI22_X1 U14986 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13359) );
  AOI22_X1 U14987 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13358) );
  NAND4_X1 U14988 ( .A1(n13361), .A2(n13360), .A3(n13359), .A4(n13358), .ZN(
        n13367) );
  AOI22_X1 U14989 ( .A1(n13583), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13365) );
  AOI22_X1 U14990 ( .A1(n12895), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13364) );
  AOI22_X1 U14991 ( .A1(n11177), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13592), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13363) );
  AOI22_X1 U14992 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13362) );
  NAND4_X1 U14993 ( .A1(n13365), .A2(n13364), .A3(n13363), .A4(n13362), .ZN(
        n13366) );
  NOR2_X1 U14994 ( .A1(n13367), .A2(n13366), .ZN(n13370) );
  INV_X1 U14995 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n22305) );
  OAI21_X1 U14996 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n22305), .A(
        n22424), .ZN(n13369) );
  NAND2_X1 U14997 ( .A1(n13156), .A2(P1_EAX_REG_19__SCAN_IN), .ZN(n13368) );
  OAI211_X1 U14998 ( .C1(n13607), .C2(n13370), .A(n13369), .B(n13368), .ZN(
        n13371) );
  NAND2_X1 U14999 ( .A1(n13372), .A2(n13371), .ZN(n16801) );
  XNOR2_X1 U15000 ( .A(n13389), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n22240) );
  NAND2_X1 U15001 ( .A1(n22240), .A2(n13582), .ZN(n13387) );
  AOI22_X1 U15002 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13376) );
  AOI22_X1 U15003 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13375) );
  AOI22_X1 U15004 ( .A1(n12895), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13374) );
  AOI22_X1 U15005 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13373) );
  NAND4_X1 U15006 ( .A1(n13376), .A2(n13375), .A3(n13374), .A4(n13373), .ZN(
        n13382) );
  AOI22_X1 U15007 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13380) );
  AOI22_X1 U15008 ( .A1(n11177), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13592), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13379) );
  AOI22_X1 U15009 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13378) );
  AOI22_X1 U15010 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13377) );
  NAND4_X1 U15011 ( .A1(n13380), .A2(n13379), .A3(n13378), .A4(n13377), .ZN(
        n13381) );
  NOR2_X1 U15012 ( .A1(n13382), .A2(n13381), .ZN(n13385) );
  INV_X1 U15013 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16993) );
  AOI21_X1 U15014 ( .B1(n16993), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13383) );
  AOI21_X1 U15015 ( .B1(n13156), .B2(P1_EAX_REG_20__SCAN_IN), .A(n13383), .ZN(
        n13384) );
  OAI21_X1 U15016 ( .B1(n13607), .B2(n13385), .A(n13384), .ZN(n13386) );
  NAND2_X1 U15017 ( .A1(n13387), .A2(n13386), .ZN(n16828) );
  INV_X1 U15018 ( .A(n13390), .ZN(n13392) );
  INV_X1 U15019 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n13391) );
  NAND2_X1 U15020 ( .A1(n13392), .A2(n13391), .ZN(n13393) );
  NAND2_X1 U15021 ( .A1(n13424), .A2(n13393), .ZN(n22258) );
  AOI22_X1 U15022 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13397) );
  AOI22_X1 U15023 ( .A1(n12896), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13396) );
  AOI22_X1 U15024 ( .A1(n11178), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13395) );
  AOI22_X1 U15025 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13394) );
  NAND4_X1 U15026 ( .A1(n13397), .A2(n13396), .A3(n13395), .A4(n13394), .ZN(
        n13403) );
  AOI22_X1 U15027 ( .A1(n12895), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13561), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13401) );
  AOI22_X1 U15028 ( .A1(n13583), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13400) );
  AOI22_X1 U15029 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13592), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13399) );
  AOI22_X1 U15030 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13398) );
  NAND4_X1 U15031 ( .A1(n13401), .A2(n13400), .A3(n13399), .A4(n13398), .ZN(
        n13402) );
  NOR2_X1 U15032 ( .A1(n13403), .A2(n13402), .ZN(n13407) );
  NAND2_X1 U15033 ( .A1(n22424), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13404) );
  NAND2_X1 U15034 ( .A1(n13557), .A2(n13404), .ZN(n13405) );
  AOI21_X1 U15035 ( .B1(n13156), .B2(P1_EAX_REG_21__SCAN_IN), .A(n13405), .ZN(
        n13406) );
  OAI21_X1 U15036 ( .B1(n13607), .B2(n13407), .A(n13406), .ZN(n13408) );
  NAND2_X1 U15037 ( .A1(n13409), .A2(n13408), .ZN(n16872) );
  XNOR2_X1 U15038 ( .A(n13424), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n22265) );
  AOI22_X1 U15039 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13413) );
  AOI22_X1 U15040 ( .A1(n12860), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13453), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13412) );
  AOI22_X1 U15041 ( .A1(n12895), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13411) );
  AOI22_X1 U15042 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13410) );
  NAND4_X1 U15043 ( .A1(n13413), .A2(n13412), .A3(n13411), .A4(n13410), .ZN(
        n13419) );
  AOI22_X1 U15044 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13417) );
  AOI22_X1 U15045 ( .A1(n11177), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13592), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13416) );
  AOI22_X1 U15046 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13415) );
  AOI22_X1 U15047 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13414) );
  NAND4_X1 U15048 ( .A1(n13417), .A2(n13416), .A3(n13415), .A4(n13414), .ZN(
        n13418) );
  OR2_X1 U15049 ( .A1(n13419), .A2(n13418), .ZN(n13422) );
  INV_X1 U15050 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14964) );
  OAI21_X1 U15051 ( .B1(n22305), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n22424), .ZN(n13420) );
  OAI21_X1 U15052 ( .B1(n13149), .B2(n14964), .A(n13420), .ZN(n13421) );
  AOI21_X1 U15053 ( .B1(n13573), .B2(n13422), .A(n13421), .ZN(n13423) );
  AOI21_X1 U15054 ( .B1(n22265), .B2(n13582), .A(n13423), .ZN(n16824) );
  NAND2_X1 U15055 ( .A1(n16823), .A2(n16824), .ZN(n16790) );
  INV_X1 U15056 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16978) );
  INV_X1 U15057 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n13448) );
  NAND2_X1 U15058 ( .A1(n13425), .A2(n13448), .ZN(n13426) );
  NAND2_X1 U15059 ( .A1(n13472), .A2(n13426), .ZN(n16971) );
  AOI22_X1 U15060 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13430) );
  AOI22_X1 U15061 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13453), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13429) );
  AOI22_X1 U15062 ( .A1(n12895), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13428) );
  AOI22_X1 U15063 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13427) );
  NAND4_X1 U15064 ( .A1(n13430), .A2(n13429), .A3(n13428), .A4(n13427), .ZN(
        n13436) );
  AOI22_X1 U15065 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13434) );
  AOI22_X1 U15066 ( .A1(n11178), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13441), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13433) );
  AOI22_X1 U15067 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13432) );
  AOI22_X1 U15068 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13431) );
  NAND4_X1 U15069 ( .A1(n13434), .A2(n13433), .A3(n13432), .A4(n13431), .ZN(
        n13435) );
  OR2_X1 U15070 ( .A1(n13436), .A2(n13435), .ZN(n13464) );
  AOI22_X1 U15071 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13440) );
  AOI22_X1 U15072 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n12860), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13439) );
  AOI22_X1 U15073 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n12895), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13438) );
  AOI22_X1 U15074 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n13561), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13437) );
  NAND4_X1 U15075 ( .A1(n13440), .A2(n13439), .A3(n13438), .A4(n13437), .ZN(
        n13447) );
  AOI22_X1 U15076 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13445) );
  AOI22_X1 U15077 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13441), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13444) );
  AOI22_X1 U15078 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13443) );
  AOI22_X1 U15079 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13442) );
  NAND4_X1 U15080 ( .A1(n13445), .A2(n13444), .A3(n13443), .A4(n13442), .ZN(
        n13446) );
  OR2_X1 U15081 ( .A1(n13447), .A2(n13446), .ZN(n13465) );
  XNOR2_X1 U15082 ( .A(n13464), .B(n13465), .ZN(n13451) );
  AOI21_X1 U15083 ( .B1(n13448), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13449) );
  AOI21_X1 U15084 ( .B1(n13612), .B2(P1_EAX_REG_23__SCAN_IN), .A(n13449), .ZN(
        n13450) );
  OAI21_X1 U15085 ( .B1(n13607), .B2(n13451), .A(n13450), .ZN(n13452) );
  OAI21_X1 U15086 ( .B1(n16971), .B2(n13557), .A(n13452), .ZN(n16791) );
  XNOR2_X1 U15087 ( .A(n13472), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16966) );
  NAND2_X1 U15088 ( .A1(n16966), .A2(n13582), .ZN(n13471) );
  AOI22_X1 U15089 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13457) );
  AOI22_X1 U15090 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13453), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13456) );
  AOI22_X1 U15091 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13455) );
  AOI22_X1 U15092 ( .A1(n13592), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13454) );
  NAND4_X1 U15093 ( .A1(n13457), .A2(n13456), .A3(n13455), .A4(n13454), .ZN(
        n13463) );
  AOI22_X1 U15094 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13595), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13461) );
  AOI22_X1 U15095 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13460) );
  AOI22_X1 U15096 ( .A1(n12895), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13459) );
  AOI22_X1 U15097 ( .A1(n11178), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13458) );
  NAND4_X1 U15098 ( .A1(n13461), .A2(n13460), .A3(n13459), .A4(n13458), .ZN(
        n13462) );
  NOR2_X1 U15099 ( .A1(n13463), .A2(n13462), .ZN(n13478) );
  NAND2_X1 U15100 ( .A1(n13465), .A2(n13464), .ZN(n13477) );
  XOR2_X1 U15101 ( .A(n13478), .B(n13477), .Z(n13466) );
  NAND2_X1 U15102 ( .A1(n13466), .A2(n13573), .ZN(n13469) );
  INV_X1 U15103 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16962) );
  AOI21_X1 U15104 ( .B1(n16962), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13467) );
  AOI21_X1 U15105 ( .B1(n13612), .B2(P1_EAX_REG_24__SCAN_IN), .A(n13467), .ZN(
        n13468) );
  NAND2_X1 U15106 ( .A1(n13469), .A2(n13468), .ZN(n13470) );
  INV_X1 U15107 ( .A(n13473), .ZN(n13475) );
  INV_X1 U15108 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n13474) );
  NAND2_X1 U15109 ( .A1(n13475), .A2(n13474), .ZN(n13476) );
  NAND2_X1 U15110 ( .A1(n13512), .A2(n13476), .ZN(n16954) );
  NOR2_X1 U15111 ( .A1(n13478), .A2(n13477), .ZN(n13507) );
  AOI22_X1 U15112 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13483) );
  AOI22_X1 U15113 ( .A1(n12860), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13482) );
  AOI22_X1 U15114 ( .A1(n12895), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13481) );
  AOI22_X1 U15115 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13480) );
  NAND4_X1 U15116 ( .A1(n13483), .A2(n13482), .A3(n13481), .A4(n13480), .ZN(
        n13489) );
  AOI22_X1 U15117 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13487) );
  AOI22_X1 U15118 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13592), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13486) );
  AOI22_X1 U15119 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13485) );
  AOI22_X1 U15120 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13484) );
  NAND4_X1 U15121 ( .A1(n13487), .A2(n13486), .A3(n13485), .A4(n13484), .ZN(
        n13488) );
  OR2_X1 U15122 ( .A1(n13489), .A2(n13488), .ZN(n13506) );
  XNOR2_X1 U15123 ( .A(n13507), .B(n13506), .ZN(n13493) );
  NAND2_X1 U15124 ( .A1(n22424), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13490) );
  NAND2_X1 U15125 ( .A1(n13557), .A2(n13490), .ZN(n13491) );
  AOI21_X1 U15126 ( .B1(n13612), .B2(P1_EAX_REG_25__SCAN_IN), .A(n13491), .ZN(
        n13492) );
  OAI21_X1 U15127 ( .B1(n13493), .B2(n13607), .A(n13492), .ZN(n13494) );
  XNOR2_X1 U15128 ( .A(n13512), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16944) );
  AOI22_X1 U15129 ( .A1(n13583), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13499) );
  AOI22_X1 U15130 ( .A1(n12895), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13498) );
  AOI22_X1 U15131 ( .A1(n13591), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13497) );
  AOI22_X1 U15132 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13496) );
  NAND4_X1 U15133 ( .A1(n13499), .A2(n13498), .A3(n13497), .A4(n13496), .ZN(
        n13505) );
  AOI22_X1 U15134 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11177), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13503) );
  AOI22_X1 U15135 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13585), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13502) );
  AOI22_X1 U15136 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13501) );
  AOI22_X1 U15137 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13592), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13500) );
  NAND4_X1 U15138 ( .A1(n13503), .A2(n13502), .A3(n13501), .A4(n13500), .ZN(
        n13504) );
  NOR2_X1 U15139 ( .A1(n13505), .A2(n13504), .ZN(n13518) );
  NAND2_X1 U15140 ( .A1(n13507), .A2(n13506), .ZN(n13517) );
  XOR2_X1 U15141 ( .A(n13518), .B(n13517), .Z(n13510) );
  INV_X1 U15142 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14972) );
  OAI21_X1 U15143 ( .B1(n22305), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n22424), .ZN(n13508) );
  OAI21_X1 U15144 ( .B1(n13149), .B2(n14972), .A(n13508), .ZN(n13509) );
  AOI21_X1 U15145 ( .B1(n13510), .B2(n13573), .A(n13509), .ZN(n13511) );
  AOI21_X1 U15146 ( .B1(n16944), .B2(n13582), .A(n13511), .ZN(n16758) );
  INV_X1 U15147 ( .A(n13512), .ZN(n13513) );
  INV_X1 U15148 ( .A(n13514), .ZN(n13515) );
  INV_X1 U15149 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n13529) );
  NAND2_X1 U15150 ( .A1(n13515), .A2(n13529), .ZN(n13516) );
  NAND2_X1 U15151 ( .A1(n13551), .A2(n13516), .ZN(n16936) );
  NOR2_X1 U15152 ( .A1(n13518), .A2(n13517), .ZN(n13546) );
  AOI22_X1 U15153 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13522) );
  AOI22_X1 U15154 ( .A1(n12860), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13453), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13521) );
  AOI22_X1 U15155 ( .A1(n12895), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13520) );
  AOI22_X1 U15156 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13519) );
  NAND4_X1 U15157 ( .A1(n13522), .A2(n13521), .A3(n13520), .A4(n13519), .ZN(
        n13528) );
  AOI22_X1 U15158 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13526) );
  AOI22_X1 U15159 ( .A1(n11177), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13592), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13525) );
  AOI22_X1 U15160 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13524) );
  AOI22_X1 U15161 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13523) );
  NAND4_X1 U15162 ( .A1(n13526), .A2(n13525), .A3(n13524), .A4(n13523), .ZN(
        n13527) );
  OR2_X1 U15163 ( .A1(n13528), .A2(n13527), .ZN(n13545) );
  XNOR2_X1 U15164 ( .A(n13546), .B(n13545), .ZN(n13532) );
  AOI21_X1 U15165 ( .B1(n13529), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13530) );
  AOI21_X1 U15166 ( .B1(n13612), .B2(P1_EAX_REG_27__SCAN_IN), .A(n13530), .ZN(
        n13531) );
  OAI21_X1 U15167 ( .B1(n13532), .B2(n13607), .A(n13531), .ZN(n13533) );
  NAND2_X1 U15168 ( .A1(n13534), .A2(n13533), .ZN(n16745) );
  XNOR2_X1 U15169 ( .A(n13551), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16930) );
  AOI22_X1 U15170 ( .A1(n12895), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13561), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13538) );
  AOI22_X1 U15171 ( .A1(n12860), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13537) );
  AOI22_X1 U15172 ( .A1(n11177), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13592), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13536) );
  AOI22_X1 U15173 ( .A1(n13453), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13535) );
  NAND4_X1 U15174 ( .A1(n13538), .A2(n13537), .A3(n13536), .A4(n13535), .ZN(
        n13544) );
  AOI22_X1 U15175 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13542) );
  AOI22_X1 U15176 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13541) );
  AOI22_X1 U15177 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13540) );
  AOI22_X1 U15178 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13539) );
  NAND4_X1 U15179 ( .A1(n13542), .A2(n13541), .A3(n13540), .A4(n13539), .ZN(
        n13543) );
  NOR2_X1 U15180 ( .A1(n13544), .A2(n13543), .ZN(n13559) );
  NAND2_X1 U15181 ( .A1(n13546), .A2(n13545), .ZN(n13558) );
  XOR2_X1 U15182 ( .A(n13559), .B(n13558), .Z(n13549) );
  INV_X1 U15183 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14958) );
  OAI21_X1 U15184 ( .B1(n22305), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n22424), .ZN(n13547) );
  OAI21_X1 U15185 ( .B1(n13149), .B2(n14958), .A(n13547), .ZN(n13548) );
  AOI21_X1 U15186 ( .B1(n13549), .B2(n13573), .A(n13548), .ZN(n13550) );
  AOI21_X1 U15187 ( .B1(n16930), .B2(n13582), .A(n13550), .ZN(n16264) );
  INV_X1 U15188 ( .A(n13551), .ZN(n13552) );
  INV_X1 U15189 ( .A(n13553), .ZN(n13555) );
  INV_X1 U15190 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13554) );
  NAND2_X1 U15191 ( .A1(n13555), .A2(n13554), .ZN(n13556) );
  NAND2_X1 U15192 ( .A1(n15064), .A2(n13556), .ZN(n16914) );
  NOR2_X1 U15193 ( .A1(n13559), .A2(n13558), .ZN(n13575) );
  AOI22_X1 U15194 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13565) );
  AOI22_X1 U15195 ( .A1(n12860), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13564) );
  AOI22_X1 U15196 ( .A1(n12895), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13563) );
  AOI22_X1 U15197 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12968), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13562) );
  NAND4_X1 U15198 ( .A1(n13565), .A2(n13564), .A3(n13563), .A4(n13562), .ZN(
        n13572) );
  AOI22_X1 U15199 ( .A1(n13115), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13570) );
  AOI22_X1 U15200 ( .A1(n11177), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13592), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13569) );
  AOI22_X1 U15201 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13568) );
  AOI22_X1 U15202 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13567) );
  NAND4_X1 U15203 ( .A1(n13570), .A2(n13569), .A3(n13568), .A4(n13567), .ZN(
        n13571) );
  OR2_X1 U15204 ( .A1(n13572), .A2(n13571), .ZN(n13574) );
  NAND2_X1 U15205 ( .A1(n13575), .A2(n13574), .ZN(n13604) );
  OAI211_X1 U15206 ( .C1(n13575), .C2(n13574), .A(n13604), .B(n13573), .ZN(
        n13579) );
  NOR2_X1 U15207 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n22305), .ZN(
        n13576) );
  NOR2_X1 U15208 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n13576), .ZN(n13577) );
  AOI21_X1 U15209 ( .B1(n13612), .B2(P1_EAX_REG_29__SCAN_IN), .A(n13577), .ZN(
        n13578) );
  NAND2_X1 U15210 ( .A1(n13579), .A2(n13578), .ZN(n13580) );
  NAND2_X1 U15211 ( .A1(n13581), .A2(n13580), .ZN(n16731) );
  XNOR2_X1 U15212 ( .A(n15064), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16904) );
  NAND2_X1 U15213 ( .A1(n16904), .A2(n13582), .ZN(n13610) );
  AOI22_X1 U15214 ( .A1(n11188), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13583), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13590) );
  AOI22_X1 U15215 ( .A1(n13585), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13479), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13589) );
  AOI22_X1 U15216 ( .A1(n12895), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12896), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13588) );
  AOI22_X1 U15217 ( .A1(n13561), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13586), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13587) );
  NAND4_X1 U15218 ( .A1(n13590), .A2(n13589), .A3(n13588), .A4(n13587), .ZN(
        n13602) );
  AOI22_X1 U15219 ( .A1(n12920), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13591), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13600) );
  AOI22_X1 U15220 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13592), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13599) );
  AOI22_X1 U15221 ( .A1(n13595), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13594), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13598) );
  AOI22_X1 U15222 ( .A1(n13566), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13596), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13597) );
  NAND4_X1 U15223 ( .A1(n13600), .A2(n13599), .A3(n13598), .A4(n13597), .ZN(
        n13601) );
  NOR2_X1 U15224 ( .A1(n13602), .A2(n13601), .ZN(n13603) );
  XNOR2_X1 U15225 ( .A(n13604), .B(n13603), .ZN(n13608) );
  INV_X1 U15226 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16906) );
  AOI21_X1 U15227 ( .B1(n16906), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13605) );
  AOI21_X1 U15228 ( .B1(n13612), .B2(P1_EAX_REG_30__SCAN_IN), .A(n13605), .ZN(
        n13606) );
  OAI21_X1 U15229 ( .B1(n13608), .B2(n13607), .A(n13606), .ZN(n13609) );
  NAND2_X1 U15230 ( .A1(n13610), .A2(n13609), .ZN(n16383) );
  AOI22_X1 U15231 ( .A1(n13612), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13611), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13613) );
  NAND2_X1 U15232 ( .A1(n12949), .A2(n11160), .ZN(n13615) );
  NAND2_X1 U15233 ( .A1(n22457), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13632) );
  OAI21_X1 U15234 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n22457), .A(
        n13632), .ZN(n13618) );
  INV_X1 U15235 ( .A(n13618), .ZN(n13616) );
  OAI211_X1 U15236 ( .C1(n14319), .C2(n14310), .A(n13641), .B(n13616), .ZN(
        n13622) );
  NAND2_X1 U15237 ( .A1(n13637), .A2(n15602), .ZN(n13670) );
  OAI21_X1 U15238 ( .B1(n13618), .B2(n13624), .A(n13670), .ZN(n13621) );
  OR2_X1 U15239 ( .A1(n11160), .A2(n22287), .ZN(n13623) );
  XNOR2_X1 U15240 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n13632), .ZN(
        n13619) );
  XNOR2_X1 U15241 ( .A(n13619), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13679) );
  INV_X1 U15242 ( .A(n13679), .ZN(n13625) );
  NAND3_X1 U15243 ( .A1(n13623), .A2(n12949), .A3(n13625), .ZN(n13620) );
  NAND3_X1 U15244 ( .A1(n13622), .A2(n13621), .A3(n13620), .ZN(n13630) );
  OAI211_X1 U15245 ( .C1(n13624), .C2(n12949), .A(n13679), .B(n13623), .ZN(
        n13628) );
  NAND2_X1 U15246 ( .A1(n13624), .A2(n15602), .ZN(n13626) );
  NAND2_X1 U15247 ( .A1(n13626), .A2(n13625), .ZN(n13627) );
  NAND2_X1 U15248 ( .A1(n13628), .A2(n13627), .ZN(n13629) );
  NAND2_X1 U15249 ( .A1(n13630), .A2(n13629), .ZN(n13639) );
  NAND2_X1 U15250 ( .A1(n18000), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13645) );
  NAND2_X1 U15251 ( .A1(n12809), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13631) );
  NAND2_X1 U15252 ( .A1(n13645), .A2(n13631), .ZN(n13643) );
  NAND2_X1 U15253 ( .A1(n22406), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13636) );
  INV_X1 U15254 ( .A(n13632), .ZN(n13634) );
  NAND2_X1 U15255 ( .A1(n13634), .A2(n13633), .ZN(n13635) );
  NAND2_X1 U15256 ( .A1(n13636), .A2(n13635), .ZN(n13642) );
  XNOR2_X1 U15257 ( .A(n13643), .B(n13642), .ZN(n13680) );
  INV_X1 U15258 ( .A(n13637), .ZN(n13658) );
  NAND2_X1 U15259 ( .A1(n13674), .A2(n13680), .ZN(n13640) );
  OAI211_X1 U15260 ( .C1(n13680), .C2(n13658), .A(n13641), .B(n13640), .ZN(
        n13638) );
  NAND2_X1 U15261 ( .A1(n13639), .A2(n13638), .ZN(n13651) );
  INV_X1 U15262 ( .A(n13640), .ZN(n13649) );
  INV_X1 U15263 ( .A(n13641), .ZN(n13648) );
  INV_X1 U15264 ( .A(n13642), .ZN(n13644) );
  NAND2_X1 U15265 ( .A1(n13646), .A2(n13645), .ZN(n13654) );
  XNOR2_X1 U15266 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13647) );
  XNOR2_X1 U15267 ( .A(n13654), .B(n13647), .ZN(n13656) );
  AOI22_X1 U15268 ( .A1(n13649), .A2(n13648), .B1(n15602), .B2(n13656), .ZN(
        n13650) );
  NAND2_X1 U15269 ( .A1(n13651), .A2(n13650), .ZN(n13660) );
  NOR2_X1 U15270 ( .A1(n11358), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13652) );
  AOI21_X1 U15271 ( .B1(n13654), .B2(n13653), .A(n13652), .ZN(n13667) );
  INV_X1 U15272 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18024) );
  NOR2_X1 U15273 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18024), .ZN(
        n13655) );
  NAND2_X1 U15274 ( .A1(n13667), .A2(n13655), .ZN(n13661) );
  INV_X1 U15275 ( .A(n13656), .ZN(n13657) );
  NAND2_X1 U15276 ( .A1(n13661), .A2(n13657), .ZN(n13682) );
  NAND2_X1 U15277 ( .A1(n13658), .A2(n13682), .ZN(n13659) );
  NAND2_X1 U15278 ( .A1(n13660), .A2(n13659), .ZN(n13665) );
  INV_X1 U15279 ( .A(n13670), .ZN(n13663) );
  INV_X1 U15280 ( .A(n13661), .ZN(n13662) );
  AOI22_X1 U15281 ( .A1(n13663), .A2(n13662), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n22287), .ZN(n13664) );
  NAND2_X1 U15282 ( .A1(n13665), .A2(n13664), .ZN(n13672) );
  NAND2_X1 U15283 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18024), .ZN(
        n13666) );
  NAND2_X1 U15284 ( .A1(n13667), .A2(n13666), .ZN(n13669) );
  INV_X1 U15285 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17942) );
  NAND2_X1 U15286 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n17942), .ZN(
        n13668) );
  INV_X1 U15287 ( .A(n13683), .ZN(n13673) );
  INV_X1 U15288 ( .A(n12940), .ZN(n13677) );
  NOR2_X1 U15289 ( .A1(n13677), .A2(n14462), .ZN(n14436) );
  NAND2_X1 U15290 ( .A1(n14436), .A2(n16724), .ZN(n14313) );
  OR2_X1 U15291 ( .A1(n16719), .A2(n14313), .ZN(n13686) );
  NAND2_X1 U15292 ( .A1(n13680), .A2(n13679), .ZN(n13681) );
  OR2_X1 U15293 ( .A1(n13682), .A2(n13681), .ZN(n13684) );
  NAND2_X1 U15294 ( .A1(n13684), .A2(n13683), .ZN(n16715) );
  NOR2_X1 U15295 ( .A1(n13678), .A2(n16715), .ZN(n14184) );
  NAND2_X1 U15296 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n22322) );
  NAND2_X1 U15297 ( .A1(n14184), .A2(n22322), .ZN(n13685) );
  NAND2_X1 U15298 ( .A1(n13686), .A2(n13685), .ZN(n14457) );
  INV_X1 U15299 ( .A(n12941), .ZN(n16150) );
  NAND3_X1 U15300 ( .A1(n16150), .A2(n14314), .A3(n12957), .ZN(n14419) );
  NOR2_X1 U15301 ( .A1(n13687), .A2(n14419), .ZN(n13688) );
  NAND2_X1 U15302 ( .A1(n17985), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n22302) );
  OAI21_X1 U15303 ( .B1(n14457), .B2(n13688), .A(n22807), .ZN(n13691) );
  NAND2_X1 U15304 ( .A1(n12947), .A2(n22322), .ZN(n13690) );
  AND2_X1 U15305 ( .A1(n16054), .A2(n16150), .ZN(n13692) );
  NOR4_X1 U15306 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13696) );
  NOR4_X1 U15307 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n13695) );
  NOR4_X1 U15308 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13694) );
  NOR4_X1 U15309 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13693) );
  AND4_X1 U15310 ( .A1(n13696), .A2(n13695), .A3(n13694), .A4(n13693), .ZN(
        n13701) );
  NOR4_X1 U15311 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13699) );
  NOR4_X1 U15312 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13698) );
  NOR4_X1 U15313 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13697) );
  INV_X1 U15314 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20636) );
  AND4_X1 U15315 ( .A1(n13699), .A2(n13698), .A3(n13697), .A4(n20636), .ZN(
        n13700) );
  NAND2_X1 U15316 ( .A1(n13701), .A2(n13700), .ZN(n13702) );
  NOR3_X1 U15317 ( .A1(n16890), .A2(n14775), .A3(n12948), .ZN(n13703) );
  AOI22_X1 U15318 ( .A1(n16892), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n16890), .ZN(n13704) );
  INV_X1 U15319 ( .A(n13704), .ZN(n13707) );
  NAND3_X1 U15320 ( .A1(n16054), .A2(n13705), .A3(n14775), .ZN(n16149) );
  INV_X1 U15321 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n22680) );
  NOR2_X1 U15322 ( .A1(n16149), .A2(n22680), .ZN(n13706) );
  AOI22_X1 U15323 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18545), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13714) );
  AOI22_X1 U15324 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13712) );
  INV_X2 U15325 ( .A(n18414), .ZN(n18547) );
  INV_X2 U15326 ( .A(n13843), .ZN(n20948) );
  AOI22_X1 U15327 ( .A1(n18547), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n20948), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13711) );
  NAND4_X1 U15328 ( .A1(n13714), .A2(n13713), .A3(n13712), .A4(n13711), .ZN(
        n13725) );
  NOR2_X2 U15329 ( .A1(n14159), .A2(n13717), .ZN(n13916) );
  NOR3_X4 U15330 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n14144), .ZN(n13798) );
  AOI22_X1 U15331 ( .A1(n13916), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13798), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13723) );
  AOI22_X1 U15332 ( .A1(n18540), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13722) );
  AOI22_X1 U15333 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11156), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13721) );
  INV_X2 U15334 ( .A(n11514), .ZN(n18480) );
  BUF_X1 U15335 ( .A(n13801), .Z(n18528) );
  AOI22_X1 U15336 ( .A1(n18480), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13720) );
  NAND4_X1 U15337 ( .A1(n13723), .A2(n13722), .A3(n13721), .A4(n13720), .ZN(
        n13724) );
  AOI22_X1 U15338 ( .A1(n18480), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13899), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13729) );
  AOI22_X1 U15339 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13728) );
  AOI22_X1 U15340 ( .A1(n13916), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13727) );
  AOI22_X1 U15341 ( .A1(n13798), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n20948), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13726) );
  NAND4_X1 U15342 ( .A1(n13729), .A2(n13728), .A3(n13727), .A4(n13726), .ZN(
        n13735) );
  INV_X2 U15343 ( .A(n18254), .ZN(n18546) );
  AOI22_X1 U15344 ( .A1(n18547), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18546), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13733) );
  AOI22_X1 U15345 ( .A1(n18540), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11157), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13732) );
  AOI22_X1 U15346 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13731) );
  AOI22_X1 U15347 ( .A1(n18545), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13730) );
  NAND4_X1 U15348 ( .A1(n13733), .A2(n13732), .A3(n13731), .A4(n13730), .ZN(
        n13734) );
  AOI22_X1 U15349 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13739) );
  BUF_X4 U15350 ( .A(n13798), .Z(n18514) );
  AOI22_X1 U15351 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18538), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13738) );
  AOI22_X1 U15352 ( .A1(n18546), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13737) );
  AOI22_X1 U15353 ( .A1(n18393), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n20948), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13736) );
  NAND4_X1 U15354 ( .A1(n13739), .A2(n13738), .A3(n13737), .A4(n13736), .ZN(
        n13745) );
  AOI22_X1 U15355 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13899), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13743) );
  AOI22_X1 U15356 ( .A1(n18547), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18540), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13742) );
  AOI22_X1 U15357 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13741) );
  AOI22_X1 U15358 ( .A1(n13916), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11156), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13740) );
  NAND4_X1 U15359 ( .A1(n13743), .A2(n13742), .A3(n13741), .A4(n13740), .ZN(
        n13744) );
  INV_X1 U15360 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13755) );
  INV_X1 U15361 ( .A(n11151), .ZN(n13754) );
  AOI22_X1 U15362 ( .A1(n18393), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n18538), .ZN(n13747) );
  OAI21_X1 U15363 ( .B1(n13843), .B2(n18563), .A(n13747), .ZN(n13748) );
  INV_X1 U15364 ( .A(n13748), .ZN(n13753) );
  INV_X2 U15365 ( .A(n18414), .ZN(n18498) );
  AOI22_X1 U15366 ( .A1(n13798), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18498), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13752) );
  AOI22_X1 U15367 ( .A1(n13916), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n13808), .ZN(n13751) );
  AOI22_X1 U15368 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n13799), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n13801), .ZN(n13750) );
  AOI22_X1 U15369 ( .A1(n13806), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n13845), .ZN(n13749) );
  INV_X1 U15370 ( .A(n13756), .ZN(n13760) );
  AOI22_X1 U15371 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n18546), .ZN(n13758) );
  AOI22_X1 U15372 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13771), .B1(
        n11156), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13757) );
  AOI22_X1 U15373 ( .A1(n18480), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13771), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13769) );
  AOI22_X1 U15374 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18546), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13768) );
  AOI22_X1 U15375 ( .A1(n18523), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13761) );
  OAI21_X1 U15376 ( .B1(n13843), .B2(n11287), .A(n13761), .ZN(n13767) );
  AOI22_X1 U15377 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13801), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13765) );
  AOI22_X1 U15378 ( .A1(n18393), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11156), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13764) );
  AOI22_X1 U15379 ( .A1(n13798), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13799), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13763) );
  AOI22_X1 U15380 ( .A1(n18498), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13808), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13762) );
  NAND4_X1 U15381 ( .A1(n13765), .A2(n13764), .A3(n13763), .A4(n13762), .ZN(
        n13766) );
  AOI22_X1 U15382 ( .A1(n13916), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11157), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13780) );
  AOI22_X1 U15383 ( .A1(n18540), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18538), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13779) );
  AOI22_X1 U15384 ( .A1(n13899), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13770) );
  OAI21_X1 U15385 ( .B1(n13843), .B2(n11271), .A(n13770), .ZN(n13777) );
  AOI22_X1 U15386 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11156), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13775) );
  AOI22_X1 U15387 ( .A1(n18545), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18546), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13774) );
  AOI22_X1 U15388 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13773) );
  AOI22_X1 U15389 ( .A1(n18547), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13772) );
  NAND4_X1 U15390 ( .A1(n13775), .A2(n13774), .A3(n13773), .A4(n13772), .ZN(
        n13776) );
  AOI211_X1 U15391 ( .C1(n11159), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n13777), .B(n13776), .ZN(n13778) );
  NAND3_X1 U15392 ( .A1(n13780), .A2(n13779), .A3(n13778), .ZN(n21386) );
  NAND2_X1 U15393 ( .A1(n13792), .A2(n21386), .ZN(n13818) );
  AOI22_X1 U15394 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13790) );
  AOI22_X1 U15395 ( .A1(n13916), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13789) );
  AOI22_X1 U15396 ( .A1(n18522), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13781) );
  OAI21_X1 U15397 ( .B1(n13843), .B2(n11261), .A(n13781), .ZN(n13787) );
  AOI22_X1 U15398 ( .A1(n18540), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18538), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13785) );
  AOI22_X1 U15399 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18545), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13784) );
  AOI22_X1 U15400 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18546), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13783) );
  AOI22_X1 U15401 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11157), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13782) );
  NAND4_X1 U15402 ( .A1(n13785), .A2(n13784), .A3(n13783), .A4(n13782), .ZN(
        n13786) );
  AOI211_X1 U15403 ( .C1(n18498), .C2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n13787), .B(n13786), .ZN(n13788) );
  NAND3_X1 U15404 ( .A1(n13790), .A2(n13789), .A3(n13788), .ZN(n21376) );
  NOR2_X1 U15405 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18755), .ZN(
        n18801) );
  AOI21_X1 U15406 ( .B1(n18755), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n18801), .ZN(n18745) );
  NOR2_X1 U15407 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18851) );
  INV_X1 U15408 ( .A(n18851), .ZN(n18858) );
  NOR4_X1 U15409 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A4(n18858), .ZN(n13830) );
  XOR2_X1 U15410 ( .A(n21376), .B(n13791), .Z(n13823) );
  NAND2_X1 U15411 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13823), .ZN(
        n13824) );
  XOR2_X1 U15412 ( .A(n21386), .B(n13792), .Z(n13816) );
  XOR2_X1 U15413 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n13816), .Z(
        n18930) );
  NOR2_X1 U15414 ( .A1(n21396), .A2(n13949), .ZN(n13794) );
  NAND2_X1 U15415 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13797), .ZN(
        n13813) );
  INV_X1 U15416 ( .A(n13949), .ZN(n21523) );
  NAND2_X1 U15417 ( .A1(n21523), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13812) );
  AOI22_X1 U15418 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13805) );
  AOI22_X1 U15419 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18545), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13804) );
  AOI22_X1 U15420 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13899), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13803) );
  AOI22_X1 U15421 ( .A1(n13746), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13802) );
  NAND4_X1 U15422 ( .A1(n13805), .A2(n13804), .A3(n13803), .A4(n13802), .ZN(
        n13811) );
  AOI22_X1 U15423 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13710), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13810) );
  AOI22_X1 U15424 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18381), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13809) );
  INV_X1 U15425 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21732) );
  NOR2_X1 U15426 ( .A1(n18968), .A2(n21732), .ZN(n18967) );
  XNOR2_X1 U15427 ( .A(n13949), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18960) );
  NAND2_X1 U15428 ( .A1(n18967), .A2(n18960), .ZN(n18959) );
  NAND2_X1 U15429 ( .A1(n13812), .A2(n18959), .ZN(n18953) );
  NAND2_X1 U15430 ( .A1(n18954), .A2(n18953), .ZN(n18952) );
  NAND2_X1 U15431 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13814), .ZN(
        n13815) );
  INV_X1 U15432 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21626) );
  XOR2_X1 U15433 ( .A(n21391), .B(n13793), .Z(n18939) );
  NAND2_X1 U15434 ( .A1(n18930), .A2(n18929), .ZN(n18928) );
  NAND2_X1 U15435 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13816), .ZN(
        n13817) );
  XOR2_X1 U15436 ( .A(n21381), .B(n13818), .Z(n13821) );
  NAND2_X1 U15437 ( .A1(n13821), .A2(n13820), .ZN(n13822) );
  XOR2_X1 U15438 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n13823), .Z(
        n18905) );
  AOI21_X1 U15439 ( .B1(n11147), .B2(n13825), .A(n18755), .ZN(n13827) );
  NAND2_X1 U15440 ( .A1(n13827), .A2(n13826), .ZN(n13828) );
  INV_X1 U15441 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21656) );
  AOI22_X1 U15442 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18845), .B1(
        n18755), .B2(n21656), .ZN(n18878) );
  NAND2_X1 U15443 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18845), .ZN(
        n13829) );
  INV_X1 U15444 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21721) );
  NAND2_X1 U15445 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21675) );
  INV_X1 U15446 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18622) );
  INV_X1 U15447 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21688) );
  NOR3_X1 U15448 ( .A1(n21675), .A2(n18622), .A3(n21688), .ZN(n21681) );
  INV_X1 U15449 ( .A(n21681), .ZN(n21684) );
  INV_X1 U15450 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21697) );
  NOR2_X1 U15451 ( .A1(n21684), .A2(n21697), .ZN(n21700) );
  NAND2_X1 U15452 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21700), .ZN(
        n21718) );
  NOR2_X1 U15453 ( .A1(n21721), .A2(n21718), .ZN(n14023) );
  NAND2_X1 U15454 ( .A1(n14023), .A2(n18847), .ZN(n13834) );
  INV_X1 U15455 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21902) );
  NAND2_X1 U15456 ( .A1(n18755), .A2(n21902), .ZN(n13831) );
  NOR2_X1 U15457 ( .A1(n13836), .A2(n13833), .ZN(n18825) );
  INV_X1 U15458 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21882) );
  NOR2_X1 U15459 ( .A1(n18755), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18670) );
  INV_X1 U15460 ( .A(n18670), .ZN(n18588) );
  NOR4_X1 U15461 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A4(n18588), .ZN(n18646) );
  INV_X1 U15462 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21737) );
  NAND2_X1 U15463 ( .A1(n18646), .A2(n21737), .ZN(n18695) );
  INV_X1 U15464 ( .A(n13834), .ZN(n13835) );
  NOR2_X1 U15465 ( .A1(n13836), .A2(n13835), .ZN(n18616) );
  NAND2_X1 U15466 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21877) );
  NOR2_X1 U15467 ( .A1(n18616), .A2(n21877), .ZN(n13838) );
  NAND2_X1 U15468 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n13838), .ZN(
        n18586) );
  INV_X1 U15469 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21854) );
  INV_X1 U15470 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21863) );
  NOR2_X1 U15471 ( .A1(n21854), .A2(n21863), .ZN(n21570) );
  NAND2_X1 U15472 ( .A1(n21570), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n18644) );
  INV_X1 U15473 ( .A(n18644), .ZN(n18741) );
  INV_X1 U15474 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21833) );
  NOR2_X1 U15475 ( .A1(n21737), .A2(n21833), .ZN(n18705) );
  NAND2_X1 U15476 ( .A1(n18741), .A2(n18705), .ZN(n21739) );
  OAI22_X1 U15477 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18695), .B1(
        n18586), .B2(n21739), .ZN(n13837) );
  INV_X1 U15478 ( .A(n13838), .ZN(n13839) );
  NAND2_X1 U15479 ( .A1(n18668), .A2(n13839), .ZN(n18587) );
  NAND2_X1 U15480 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18587), .ZN(
        n18645) );
  INV_X1 U15481 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21760) );
  INV_X1 U15482 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21762) );
  NOR2_X1 U15483 ( .A1(n21760), .A2(n21762), .ZN(n18738) );
  AOI21_X1 U15484 ( .B1(n21760), .B2(n21762), .A(n18755), .ZN(n13840) );
  INV_X1 U15485 ( .A(n13840), .ZN(n13841) );
  INV_X1 U15486 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21778) );
  NAND2_X1 U15487 ( .A1(n13842), .A2(n21778), .ZN(n14031) );
  NOR2_X1 U15488 ( .A1(n13842), .A2(n21778), .ZN(n14016) );
  NAND2_X1 U15489 ( .A1(n18745), .A2(n18744), .ZN(n18743) );
  AOI22_X1 U15490 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13854) );
  AOI22_X1 U15491 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n18432), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13853) );
  AOI22_X1 U15492 ( .A1(n18522), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13844) );
  OAI21_X1 U15493 ( .B1(n18254), .B2(n18563), .A(n13844), .ZN(n13851) );
  AOI22_X1 U15494 ( .A1(n18547), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18381), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13849) );
  INV_X2 U15495 ( .A(n11206), .ZN(n18393) );
  AOI22_X1 U15496 ( .A1(n18393), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11156), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13848) );
  AOI22_X1 U15497 ( .A1(n18480), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13899), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13847) );
  AOI22_X1 U15498 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13846) );
  NAND4_X1 U15499 ( .A1(n13849), .A2(n13848), .A3(n13847), .A4(n13846), .ZN(
        n13850) );
  AOI22_X1 U15500 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18540), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13858) );
  AOI22_X1 U15501 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11156), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13857) );
  AOI22_X1 U15502 ( .A1(n18547), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18480), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13856) );
  AOI22_X1 U15503 ( .A1(n18279), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13855) );
  NAND4_X1 U15504 ( .A1(n13858), .A2(n13857), .A3(n13856), .A4(n13855), .ZN(
        n13864) );
  AOI22_X1 U15505 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13861) );
  AOI22_X1 U15506 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11157), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13860) );
  AOI22_X1 U15507 ( .A1(n18528), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13859) );
  NAND4_X1 U15508 ( .A1(n13862), .A2(n13861), .A3(n13860), .A4(n13859), .ZN(
        n13863) );
  AOI22_X1 U15509 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18540), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13868) );
  AOI22_X1 U15510 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18546), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13867) );
  AOI22_X1 U15511 ( .A1(n13916), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13798), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13866) );
  AOI22_X1 U15512 ( .A1(n18279), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13865) );
  NAND4_X1 U15513 ( .A1(n13868), .A2(n13867), .A3(n13866), .A4(n13865), .ZN(
        n13874) );
  AOI22_X1 U15514 ( .A1(n18523), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18538), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13872) );
  AOI22_X1 U15515 ( .A1(n18393), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13871) );
  AOI22_X1 U15516 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18498), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13870) );
  AOI22_X1 U15517 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13899), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13869) );
  NAND4_X1 U15518 ( .A1(n13872), .A2(n13871), .A3(n13870), .A4(n13869), .ZN(
        n13873) );
  AOI22_X1 U15519 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13878) );
  AOI22_X1 U15520 ( .A1(n18393), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18480), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13877) );
  AOI22_X1 U15521 ( .A1(n18547), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18381), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13876) );
  AOI22_X1 U15522 ( .A1(n18279), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13875) );
  NAND4_X1 U15523 ( .A1(n13878), .A2(n13877), .A3(n13876), .A4(n13875), .ZN(
        n13884) );
  AOI22_X1 U15524 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13899), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13882) );
  AOI22_X1 U15525 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13881) );
  AOI22_X1 U15526 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13880) );
  NAND4_X1 U15527 ( .A1(n13882), .A2(n13881), .A3(n13880), .A4(n13879), .ZN(
        n13883) );
  AOI22_X1 U15528 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13888) );
  AOI22_X1 U15529 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13899), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13887) );
  AOI22_X1 U15530 ( .A1(n18523), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13886) );
  AOI22_X1 U15531 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n20948), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13885) );
  NAND4_X1 U15532 ( .A1(n13888), .A2(n13887), .A3(n13886), .A4(n13885), .ZN(
        n13894) );
  AOI22_X1 U15533 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18540), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13891) );
  AOI22_X1 U15534 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18480), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13890) );
  AOI22_X1 U15535 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18545), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13889) );
  NAND4_X1 U15536 ( .A1(n13892), .A2(n13891), .A3(n13890), .A4(n13889), .ZN(
        n13893) );
  NOR2_X1 U15537 ( .A1(n19605), .A2(n21405), .ZN(n14010) );
  NOR2_X1 U15538 ( .A1(n21524), .A2(n14010), .ZN(n13930) );
  INV_X1 U15539 ( .A(n14010), .ZN(n13931) );
  AOI22_X1 U15540 ( .A1(n18480), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13898) );
  AOI22_X1 U15541 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13897) );
  AOI22_X1 U15542 ( .A1(n18540), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13896) );
  NAND4_X1 U15543 ( .A1(n13898), .A2(n13897), .A3(n13896), .A4(n13895), .ZN(
        n13905) );
  AOI22_X1 U15544 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18547), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13903) );
  AOI22_X1 U15545 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11157), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13902) );
  AOI22_X1 U15546 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13899), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13901) );
  AOI22_X1 U15547 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18545), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13900) );
  NAND4_X1 U15548 ( .A1(n13903), .A2(n13902), .A3(n13901), .A4(n13900), .ZN(
        n13904) );
  AOI22_X1 U15549 ( .A1(n13899), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13909) );
  AOI22_X1 U15550 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18498), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13908) );
  AOI22_X1 U15551 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18545), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13907) );
  AOI22_X1 U15552 ( .A1(n18279), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13906) );
  NAND4_X1 U15553 ( .A1(n13909), .A2(n13908), .A3(n13907), .A4(n13906), .ZN(
        n13915) );
  AOI22_X1 U15554 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18381), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13912) );
  AOI22_X1 U15555 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18432), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13911) );
  AOI22_X1 U15556 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13910) );
  NAND4_X1 U15557 ( .A1(n13913), .A2(n13912), .A3(n13911), .A4(n13910), .ZN(
        n13914) );
  INV_X2 U15558 ( .A(n20904), .ZN(n21337) );
  OR2_X1 U15559 ( .A1(n14000), .A2(n13934), .ZN(n13981) );
  NAND2_X1 U15560 ( .A1(n21336), .A2(n21443), .ZN(n13932) );
  NOR2_X1 U15561 ( .A1(n20904), .A2(n13932), .ZN(n13936) );
  AOI22_X1 U15562 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18545), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13926) );
  AOI22_X1 U15563 ( .A1(n18547), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18381), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13925) );
  INV_X1 U15564 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18213) );
  AOI22_X1 U15565 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11157), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13917) );
  OAI21_X1 U15566 ( .B1(n18254), .B2(n18213), .A(n13917), .ZN(n13923) );
  AOI22_X1 U15567 ( .A1(n13899), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13921) );
  AOI22_X1 U15568 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18480), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13920) );
  AOI22_X1 U15569 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13919) );
  AOI22_X1 U15570 ( .A1(n18279), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13918) );
  NAND4_X1 U15571 ( .A1(n13921), .A2(n13920), .A3(n13919), .A4(n13918), .ZN(
        n13922) );
  AOI211_X1 U15572 ( .C1(n18388), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n13923), .B(n13922), .ZN(n13924) );
  NAND3_X1 U15573 ( .A1(n13926), .A2(n13925), .A3(n13924), .ZN(n13935) );
  NOR3_X1 U15574 ( .A1(n13934), .A2(n13936), .A3(n13935), .ZN(n13928) );
  NAND2_X1 U15575 ( .A1(n21405), .A2(n13977), .ZN(n14142) );
  NAND2_X1 U15576 ( .A1(n19727), .A2(n19645), .ZN(n13984) );
  NAND2_X1 U15577 ( .A1(n21404), .A2(n19727), .ZN(n14006) );
  AND2_X1 U15578 ( .A1(n13935), .A2(n14006), .ZN(n13927) );
  AOI211_X1 U15579 ( .C1(n13931), .C2(n13981), .A(n13928), .B(n13933), .ZN(
        n13929) );
  NAND2_X1 U15580 ( .A1(n21443), .A2(n21345), .ZN(n21344) );
  NAND3_X1 U15581 ( .A1(n21337), .A2(n19027), .A3(n21344), .ZN(n13983) );
  NOR4_X2 U15582 ( .A1(n13935), .A2(n13977), .A3(n13932), .A4(n13931), .ZN(
        n13964) );
  NAND2_X1 U15583 ( .A1(n13964), .A2(n14000), .ZN(n13979) );
  NAND2_X1 U15584 ( .A1(n13979), .A2(n13937), .ZN(n14130) );
  INV_X1 U15585 ( .A(n13935), .ZN(n19687) );
  NAND2_X1 U15586 ( .A1(n19727), .A2(n19687), .ZN(n14141) );
  NOR2_X1 U15587 ( .A1(n11300), .A2(n14141), .ZN(n14491) );
  INV_X1 U15588 ( .A(n13966), .ZN(n20843) );
  NAND2_X1 U15589 ( .A1(n20904), .A2(n13976), .ZN(n14139) );
  NAND2_X1 U15590 ( .A1(n14141), .A2(n14139), .ZN(n13968) );
  INV_X1 U15591 ( .A(n13968), .ZN(n13938) );
  XOR2_X1 U15592 ( .A(n20904), .B(n21336), .Z(n20835) );
  INV_X1 U15593 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18585) );
  NOR2_X1 U15594 ( .A1(n21877), .A2(n18585), .ZN(n18591) );
  NAND2_X1 U15595 ( .A1(n14023), .A2(n18591), .ZN(n18590) );
  INV_X1 U15596 ( .A(n18590), .ZN(n13973) );
  AOI21_X1 U15597 ( .B1(n13949), .B2(n21525), .A(n21396), .ZN(n13944) );
  NOR2_X1 U15598 ( .A1(n21391), .A2(n13944), .ZN(n13953) );
  NAND2_X1 U15599 ( .A1(n13953), .A2(n21386), .ZN(n13941) );
  NOR2_X1 U15600 ( .A1(n21381), .A2(n13941), .ZN(n13940) );
  NAND2_X1 U15601 ( .A1(n13940), .A2(n21376), .ZN(n13939) );
  NOR2_X1 U15602 ( .A1(n11148), .A2(n13939), .ZN(n13962) );
  XOR2_X1 U15603 ( .A(n11147), .B(n13939), .Z(n18891) );
  XOR2_X1 U15604 ( .A(n21376), .B(n13940), .Z(n13956) );
  XOR2_X1 U15605 ( .A(n21381), .B(n13941), .Z(n13942) );
  NAND2_X1 U15606 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13942), .ZN(
        n13955) );
  XOR2_X1 U15607 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n13942), .Z(
        n18920) );
  XOR2_X1 U15608 ( .A(n21391), .B(n13944), .Z(n13943) );
  NAND2_X1 U15609 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13943), .ZN(
        n13951) );
  XOR2_X1 U15610 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n13943), .Z(
        n18944) );
  INV_X1 U15611 ( .A(n13944), .ZN(n13945) );
  OAI21_X1 U15612 ( .B1(n18968), .B2(n13793), .A(n13945), .ZN(n13946) );
  NAND2_X1 U15613 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13946), .ZN(
        n13950) );
  XNOR2_X1 U15614 ( .A(n13796), .B(n13946), .ZN(n18951) );
  AOI21_X1 U15615 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13949), .A(
        n21525), .ZN(n13948) );
  NOR2_X1 U15616 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13949), .ZN(
        n13947) );
  AOI221_X1 U15617 ( .B1(n21525), .B2(n13949), .C1(n13948), .C2(n21732), .A(
        n13947), .ZN(n18950) );
  NAND2_X1 U15618 ( .A1(n18951), .A2(n18950), .ZN(n18949) );
  NAND2_X1 U15619 ( .A1(n13950), .A2(n18949), .ZN(n18943) );
  NAND2_X1 U15620 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13952), .ZN(
        n13954) );
  INV_X1 U15621 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21625) );
  XOR2_X1 U15622 ( .A(n21386), .B(n13953), .Z(n18926) );
  NAND2_X1 U15623 ( .A1(n13954), .A2(n18925), .ZN(n18919) );
  NAND2_X1 U15624 ( .A1(n18920), .A2(n18919), .ZN(n18918) );
  NAND2_X1 U15625 ( .A1(n13955), .A2(n18918), .ZN(n13957) );
  NAND2_X1 U15626 ( .A1(n13956), .A2(n13957), .ZN(n13958) );
  XOR2_X1 U15627 ( .A(n13957), .B(n13956), .Z(n18901) );
  NAND2_X1 U15628 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18901), .ZN(
        n18900) );
  INV_X1 U15629 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21655) );
  NAND2_X1 U15630 ( .A1(n13962), .A2(n13959), .ZN(n13963) );
  NAND2_X1 U15631 ( .A1(n18891), .A2(n18892), .ZN(n18890) );
  NAND2_X1 U15632 ( .A1(n13962), .A2(n13961), .ZN(n13960) );
  OAI211_X1 U15633 ( .C1(n13962), .C2(n13961), .A(n18890), .B(n13960), .ZN(
        n18880) );
  NAND2_X1 U15634 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18880), .ZN(
        n18879) );
  NAND2_X1 U15635 ( .A1(n13963), .A2(n18879), .ZN(n14024) );
  INV_X1 U15636 ( .A(n14024), .ZN(n21670) );
  NAND2_X1 U15637 ( .A1(n14137), .A2(n11148), .ZN(n21927) );
  INV_X1 U15638 ( .A(n21928), .ZN(n21870) );
  OAI22_X1 U15639 ( .A1(n21670), .A2(n21847), .B1(n21927), .B2(n21870), .ZN(
        n21686) );
  INV_X1 U15640 ( .A(n18591), .ZN(n13972) );
  INV_X1 U15641 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21536) );
  NOR2_X1 U15642 ( .A1(n13796), .A2(n21536), .ZN(n21601) );
  INV_X1 U15643 ( .A(n21601), .ZN(n21603) );
  NOR3_X1 U15644 ( .A1(n21625), .A2(n21626), .A3(n11439), .ZN(n13967) );
  INV_X1 U15645 ( .A(n13967), .ZN(n21633) );
  NOR2_X1 U15646 ( .A1(n21603), .A2(n21633), .ZN(n21622) );
  NAND2_X1 U15647 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21622), .ZN(
        n21647) );
  NOR2_X1 U15648 ( .A1(n21655), .A2(n21647), .ZN(n21935) );
  NAND2_X1 U15649 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21935), .ZN(
        n21674) );
  INV_X1 U15650 ( .A(n21674), .ZN(n21699) );
  NAND2_X1 U15651 ( .A1(n14023), .A2(n21699), .ZN(n21563) );
  INV_X1 U15652 ( .A(n21563), .ZN(n21873) );
  INV_X1 U15653 ( .A(n13964), .ZN(n13965) );
  NOR2_X1 U15654 ( .A1(n13965), .A2(n14140), .ZN(n14173) );
  NOR2_X2 U15655 ( .A1(n13966), .A2(n14173), .ZN(n21340) );
  NAND2_X1 U15656 ( .A1(n14133), .A2(n21340), .ZN(n17953) );
  NAND2_X1 U15657 ( .A1(n21873), .A2(n21746), .ZN(n13971) );
  INV_X1 U15658 ( .A(n14023), .ZN(n21884) );
  INV_X1 U15659 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21642) );
  OAI21_X1 U15660 ( .B1(n21536), .B2(n21732), .A(n13796), .ZN(n21605) );
  NAND2_X1 U15661 ( .A1(n13967), .A2(n21605), .ZN(n21623) );
  NOR2_X1 U15662 ( .A1(n21642), .A2(n21623), .ZN(n21645) );
  NAND3_X1 U15663 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n21645), .ZN(n21673) );
  NOR2_X1 U15664 ( .A1(n21884), .A2(n21673), .ZN(n14019) );
  INV_X1 U15665 ( .A(n14019), .ZN(n21876) );
  NOR2_X1 U15666 ( .A1(n13972), .A2(n21876), .ZN(n21565) );
  NAND2_X1 U15667 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21699), .ZN(
        n21931) );
  NOR2_X1 U15668 ( .A1(n18590), .A2(n21931), .ZN(n21561) );
  AOI21_X1 U15669 ( .B1(n13969), .B2(n13968), .A(n14153), .ZN(n21925) );
  AOI22_X1 U15670 ( .A1(n21875), .A2(n21565), .B1(n21561), .B2(n21731), .ZN(
        n13970) );
  OAI21_X1 U15671 ( .B1(n13972), .B2(n13971), .A(n13970), .ZN(n21738) );
  AOI21_X1 U15672 ( .B1(n13973), .B2(n21686), .A(n21738), .ZN(n21572) );
  NOR2_X1 U15673 ( .A1(n21572), .A2(n18644), .ZN(n21757) );
  NAND2_X1 U15674 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n21757), .ZN(
        n21834) );
  NAND3_X1 U15675 ( .A1(n18738), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21772) );
  NOR2_X1 U15676 ( .A1(n21834), .A2(n21772), .ZN(n21780) );
  INV_X1 U15677 ( .A(n13974), .ZN(n13985) );
  AOI211_X1 U15678 ( .C1(n21345), .C2(n13977), .A(n13976), .B(n13975), .ZN(
        n13978) );
  INV_X1 U15679 ( .A(n13978), .ZN(n13980) );
  OAI21_X1 U15680 ( .B1(n13981), .B2(n13980), .A(n13979), .ZN(n13982) );
  OAI211_X1 U15681 ( .C1(n13985), .C2(n13984), .A(n13983), .B(n13982), .ZN(
        n14134) );
  NAND2_X1 U15682 ( .A1(n19530), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13986) );
  OAI21_X1 U15683 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19530), .A(
        n13986), .ZN(n14008) );
  AOI22_X1 U15684 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19524), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n21541), .ZN(n14002) );
  OAI22_X1 U15685 ( .A1(n21550), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n19523), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13993) );
  OAI21_X1 U15686 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n21550), .A(
        n13988), .ZN(n13989) );
  OAI22_X1 U15687 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17950), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13989), .ZN(n13996) );
  NOR2_X1 U15688 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17950), .ZN(
        n13990) );
  NAND2_X1 U15689 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13989), .ZN(
        n13995) );
  AOI22_X1 U15690 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13996), .B1(
        n13990), .B2(n13995), .ZN(n13991) );
  NAND2_X1 U15691 ( .A1(n14002), .A2(n13991), .ZN(n13999) );
  OAI21_X1 U15692 ( .B1(n13994), .B2(n13993), .A(n13991), .ZN(n13992) );
  AOI21_X1 U15693 ( .B1(n13994), .B2(n13993), .A(n13992), .ZN(n14007) );
  INV_X1 U15694 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14171) );
  AND2_X1 U15695 ( .A1(n13995), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13997) );
  OAI22_X1 U15696 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n14171), .B1(
        n13997), .B2(n13996), .ZN(n14004) );
  NOR2_X1 U15697 ( .A1(n14007), .A2(n14004), .ZN(n13998) );
  OAI21_X1 U15698 ( .B1(n14008), .B2(n13999), .A(n13998), .ZN(n14114) );
  XOR2_X1 U15699 ( .A(n14000), .B(n21337), .Z(n14001) );
  INV_X1 U15700 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n22356) );
  NAND2_X1 U15701 ( .A1(n22361), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19068) );
  NOR2_X1 U15702 ( .A1(n22356), .A2(n19068), .ZN(n19062) );
  OAI211_X1 U15703 ( .C1(P3_STATE_REG_2__SCAN_IN), .C2(P3_STATE_REG_1__SCAN_IN), .A(n22359), .B(n22361), .ZN(n20834) );
  NAND2_X1 U15704 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n22363) );
  INV_X1 U15705 ( .A(n22363), .ZN(n22367) );
  AOI21_X1 U15706 ( .B1(n14001), .B2(n20834), .A(n22367), .ZN(n14131) );
  XOR2_X1 U15707 ( .A(n14003), .B(n14002), .Z(n14005) );
  NAND3_X1 U15708 ( .A1(n14131), .A2(n14129), .A3(n14006), .ZN(n14013) );
  INV_X1 U15709 ( .A(n14007), .ZN(n14009) );
  OAI21_X1 U15710 ( .B1(n14009), .B2(n14008), .A(n14129), .ZN(n14136) );
  NOR2_X1 U15711 ( .A1(n21337), .A2(n14136), .ZN(n14011) );
  INV_X1 U15712 ( .A(n14114), .ZN(n14490) );
  OAI211_X1 U15713 ( .C1(n14011), .C2(n14490), .A(n14010), .B(n19727), .ZN(
        n14012) );
  OAI211_X1 U15714 ( .C1(n19645), .C2(n14114), .A(n14013), .B(n14012), .ZN(
        n14014) );
  NOR2_X1 U15715 ( .A1(n21960), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n20895) );
  NAND2_X1 U15716 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n20895), .ZN(n21961) );
  INV_X1 U15717 ( .A(n21961), .ZN(n21956) );
  OAI21_X2 U15718 ( .B1(n14134), .B2(n14014), .A(n21956), .ZN(n21930) );
  INV_X1 U15719 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n18742) );
  NOR2_X1 U15720 ( .A1(n18742), .A2(n18845), .ZN(n14015) );
  NAND2_X1 U15721 ( .A1(n14016), .A2(n14015), .ZN(n18788) );
  INV_X1 U15722 ( .A(n18788), .ZN(n18799) );
  AOI221_X1 U15723 ( .B1(n11145), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), 
        .C1(n14017), .C2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(n18799), .ZN(
        n14028) );
  NAND2_X1 U15724 ( .A1(n18591), .A2(n18741), .ZN(n14025) );
  NOR2_X1 U15725 ( .A1(n21737), .A2(n14025), .ZN(n14018) );
  NAND2_X1 U15726 ( .A1(n21873), .A2(n14018), .ZN(n21745) );
  NOR3_X1 U15727 ( .A1(n21772), .A2(n21778), .A3(n21745), .ZN(n14020) );
  NOR2_X1 U15728 ( .A1(n21936), .A2(n14020), .ZN(n14022) );
  NAND2_X1 U15729 ( .A1(n14019), .A2(n14018), .ZN(n21742) );
  OAI21_X1 U15730 ( .B1(n21772), .B2(n21742), .A(n21875), .ZN(n21773) );
  OAI221_X1 U15731 ( .B1(n21925), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C1(
        n21925), .C2(n14020), .A(n21773), .ZN(n14021) );
  NOR2_X1 U15732 ( .A1(n14022), .A2(n14021), .ZN(n21786) );
  INV_X1 U15733 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n21740) );
  NAND2_X1 U15734 ( .A1(n21928), .A2(n14023), .ZN(n21720) );
  NAND2_X1 U15735 ( .A1(n18705), .A2(n21567), .ZN(n21827) );
  AND3_X1 U15736 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18738), .A3(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21796) );
  NAND2_X1 U15737 ( .A1(n18737), .A2(n21796), .ZN(n18796) );
  INV_X1 U15738 ( .A(n21847), .ZN(n21826) );
  INV_X1 U15739 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21693) );
  NAND2_X1 U15740 ( .A1(n21700), .A2(n14024), .ZN(n18834) );
  NAND2_X1 U15741 ( .A1(n21796), .A2(n18736), .ZN(n18795) );
  AOI22_X1 U15742 ( .A1(n21871), .A2(n18796), .B1(n21826), .B2(n18795), .ZN(
        n14026) );
  NOR2_X1 U15743 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n21952) );
  NAND2_X1 U15744 ( .A1(n21952), .A2(n21949), .ZN(n18571) );
  NAND2_X1 U15745 ( .A1(n21875), .A2(n21778), .ZN(n21787) );
  NAND4_X1 U15746 ( .A1(n21786), .A2(n14026), .A3(n21828), .A4(n21787), .ZN(
        n14027) );
  OR2_X1 U15747 ( .A1(n14028), .A2(n14027), .ZN(n14029) );
  OAI211_X1 U15748 ( .C1(n11199), .C2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14029), .B(n14030), .ZN(n14033) );
  INV_X1 U15749 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n21275) );
  NOR2_X1 U15750 ( .A1(n14030), .A2(n21275), .ZN(n18729) );
  NAND2_X1 U15751 ( .A1(n21897), .A2(n14137), .ZN(n21653) );
  NAND2_X1 U15752 ( .A1(n14035), .A2(n11214), .ZN(n14037) );
  NAND2_X1 U15753 ( .A1(n14037), .A2(n14036), .ZN(n17484) );
  OAI21_X1 U15754 ( .B1(n17483), .B2(n17494), .A(n17484), .ZN(n14040) );
  XNOR2_X1 U15755 ( .A(n14038), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14039) );
  XNOR2_X1 U15756 ( .A(n14040), .B(n14039), .ZN(n14059) );
  OR2_X1 U15757 ( .A1(n14082), .A2(n14041), .ZN(n14042) );
  NAND2_X1 U15758 ( .A1(n16644), .A2(n14042), .ZN(n19311) );
  NOR2_X1 U15759 ( .A1(n19380), .A2(n14043), .ZN(n14054) );
  NOR2_X1 U15760 ( .A1(n18112), .A2(n19313), .ZN(n14044) );
  AOI211_X1 U15761 ( .C1(n18102), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14054), .B(n14044), .ZN(n14045) );
  OAI21_X1 U15762 ( .B1(n19311), .B2(n18105), .A(n14045), .ZN(n14046) );
  AOI21_X1 U15763 ( .B1(n14059), .B2(n18079), .A(n14046), .ZN(n14048) );
  XNOR2_X1 U15764 ( .A(n17493), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14060) );
  NAND2_X1 U15765 ( .A1(n14048), .A2(n14047), .ZN(P2_U2986) );
  OR2_X1 U15766 ( .A1(n14052), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17664) );
  INV_X1 U15767 ( .A(n17663), .ZN(n14049) );
  NAND2_X1 U15768 ( .A1(n17664), .A2(n14049), .ZN(n17650) );
  AND2_X1 U15769 ( .A1(n14085), .A2(n14050), .ZN(n14051) );
  OR2_X1 U15770 ( .A1(n14051), .A2(n16649), .ZN(n19309) );
  OR2_X1 U15771 ( .A1(n17494), .A2(n14052), .ZN(n17649) );
  NOR2_X1 U15772 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17649), .ZN(
        n14053) );
  NOR2_X1 U15773 ( .A1(n14054), .A2(n14053), .ZN(n14055) );
  OAI21_X1 U15774 ( .B1(n17928), .B2(n19309), .A(n14055), .ZN(n14056) );
  AOI21_X1 U15775 ( .B1(n17650), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14056), .ZN(n14057) );
  OAI21_X1 U15776 ( .B1(n19311), .B2(n19416), .A(n14057), .ZN(n14058) );
  AOI21_X1 U15777 ( .B1(n14059), .B2(n19419), .A(n14058), .ZN(n14062) );
  NAND2_X1 U15778 ( .A1(n14062), .A2(n14061), .ZN(P2_U3018) );
  INV_X1 U15779 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20830) );
  NOR3_X1 U15780 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20830), .ZN(n14064) );
  NOR4_X1 U15781 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n14063) );
  NAND4_X1 U15782 ( .A1(n14775), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n14064), .A4(
        n14063), .ZN(U214) );
  NOR4_X1 U15783 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n14068) );
  NOR4_X1 U15784 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n14067) );
  NOR4_X1 U15785 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n14066) );
  NOR4_X1 U15786 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n14065) );
  AND4_X1 U15787 ( .A1(n14068), .A2(n14067), .A3(n14066), .A4(n14065), .ZN(
        n14073) );
  NOR4_X1 U15788 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n14071) );
  NOR4_X1 U15789 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n14070) );
  NOR4_X1 U15790 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n14069) );
  INV_X1 U15791 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20551) );
  AND4_X1 U15792 ( .A1(n14071), .A2(n14070), .A3(n14069), .A4(n20551), .ZN(
        n14072) );
  NAND2_X1 U15793 ( .A1(n14073), .A2(n14072), .ZN(n14074) );
  NAND2_X2 U15794 ( .A1(n14074), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n16030)
         );
  NOR2_X1 U15795 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n14076) );
  NOR4_X1 U15796 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n14075) );
  NAND4_X1 U15797 ( .A1(n14076), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n14075), .ZN(n14077) );
  NOR2_X1 U15798 ( .A1(n16030), .A2(n14077), .ZN(n20771) );
  NAND2_X1 U15799 ( .A1(n20771), .A2(U214), .ZN(U212) );
  NOR2_X1 U15800 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n14077), .ZN(n19476)
         );
  AOI211_X1 U15801 ( .C1(n14079), .C2(n17487), .A(n19318), .B(n19432), .ZN(
        n14089) );
  OAI22_X1 U15802 ( .A1(n14080), .A2(n19342), .B1(n18201), .B2(n19338), .ZN(
        n14088) );
  AOI22_X1 U15803 ( .A1(n19328), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n19346), .ZN(n14081) );
  INV_X1 U15804 ( .A(n14081), .ZN(n14087) );
  AOI21_X1 U15805 ( .B1(n14083), .B2(n17385), .A(n14082), .ZN(n17491) );
  INV_X1 U15806 ( .A(n17491), .ZN(n17666) );
  OAI21_X1 U15807 ( .B1(n11421), .B2(n11240), .A(n14085), .ZN(n17661) );
  OAI22_X1 U15808 ( .A1(n17666), .A2(n19310), .B1(n17661), .B2(n19336), .ZN(
        n14086) );
  OR4_X1 U15809 ( .A1(n14089), .A2(n14088), .A3(n14087), .A4(n14086), .ZN(
        P2_U2828) );
  AOI211_X1 U15810 ( .C1(n19277), .C2(n14091), .A(n14090), .B(n19432), .ZN(
        n14098) );
  INV_X1 U15811 ( .A(n14092), .ZN(n14093) );
  OAI22_X1 U15812 ( .A1(n14093), .A2(n19342), .B1(n11805), .B2(n19338), .ZN(
        n14097) );
  AOI22_X1 U15813 ( .A1(n19328), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n19346), .ZN(n14094) );
  INV_X1 U15814 ( .A(n14094), .ZN(n14096) );
  OAI22_X1 U15815 ( .A1(n17421), .A2(n19310), .B1(n17476), .B2(n19336), .ZN(
        n14095) );
  OR4_X1 U15816 ( .A1(n14098), .A2(n14097), .A3(n14096), .A4(n14095), .ZN(
        P2_U2834) );
  AOI211_X1 U15817 ( .C1(n14100), .C2(n17532), .A(n14099), .B(n19432), .ZN(
        n14113) );
  INV_X1 U15818 ( .A(n14101), .ZN(n14102) );
  OAI22_X1 U15819 ( .A1(n14102), .A2(n19342), .B1(n19237), .B2(n12232), .ZN(
        n14112) );
  AOI22_X1 U15820 ( .A1(n19328), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19307), .ZN(n14103) );
  INV_X1 U15821 ( .A(n14103), .ZN(n14111) );
  INV_X1 U15822 ( .A(n17401), .ZN(n14105) );
  AOI21_X1 U15823 ( .B1(n14106), .B2(n14104), .A(n14105), .ZN(n17715) );
  INV_X1 U15824 ( .A(n17715), .ZN(n14109) );
  OAI21_X1 U15825 ( .B1(n14108), .B2(n11226), .A(n14107), .ZN(n17712) );
  OAI22_X1 U15826 ( .A1(n14109), .A2(n19310), .B1(n17712), .B2(n19336), .ZN(
        n14110) );
  OR4_X1 U15827 ( .A1(n14113), .A2(n14112), .A3(n14111), .A4(n14110), .ZN(
        P2_U2832) );
  INV_X1 U15828 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19054) );
  NOR2_X1 U15829 ( .A1(n14030), .A2(n19054), .ZN(n14128) );
  NOR2_X1 U15830 ( .A1(n21675), .A2(n18622), .ZN(n21685) );
  NAND2_X1 U15831 ( .A1(n11145), .A2(n14124), .ZN(n18839) );
  AOI211_X1 U15832 ( .C1(n21675), .C2(n18622), .A(n21685), .B(n18643), .ZN(
        n14127) );
  AND2_X2 U15833 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18934) );
  INV_X2 U15834 ( .A(n18886), .ZN(n20970) );
  INV_X1 U15835 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n21007) );
  INV_X1 U15836 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20984) );
  INV_X1 U15837 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n21030) );
  NOR4_X2 U15838 ( .A1(n21007), .A2(n20984), .A3(n18862), .A4(n21030), .ZN(
        n14117) );
  AND2_X1 U15839 ( .A1(n14117), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n14115) );
  INV_X1 U15840 ( .A(n18624), .ZN(n14119) );
  INV_X1 U15841 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n21858) );
  NOR2_X1 U15842 ( .A1(n21537), .A2(n21858), .ZN(n18572) );
  NAND2_X1 U15843 ( .A1(n14171), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21532) );
  OAI21_X1 U15844 ( .B1(n21952), .B2(n18572), .A(n21532), .ZN(n19478) );
  NAND2_X1 U15845 ( .A1(n21960), .A2(n19478), .ZN(n19686) );
  NAND3_X1 U15846 ( .A1(n21858), .A2(n21949), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n19526) );
  NOR2_X1 U15847 ( .A1(n14119), .A2(n19813), .ZN(n18830) );
  NOR2_X1 U15848 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18572), .ZN(n20833) );
  NAND2_X1 U15849 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18933) );
  INV_X1 U15850 ( .A(n18933), .ZN(n18728) );
  NOR2_X1 U15851 ( .A1(n18957), .A2(n18728), .ZN(n18908) );
  INV_X1 U15852 ( .A(n18908), .ZN(n18964) );
  INV_X1 U15853 ( .A(n14117), .ZN(n21041) );
  NOR3_X1 U15854 ( .A1(n18886), .A2(n21041), .A3(n19813), .ZN(n18855) );
  AOI21_X1 U15855 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18964), .A(
        n18855), .ZN(n14120) );
  NAND2_X1 U15856 ( .A1(n21960), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18969) );
  INV_X1 U15857 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n22315) );
  NAND2_X1 U15858 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14118) );
  INV_X1 U15859 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20902) );
  NAND2_X1 U15860 ( .A1(n20970), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n21000) );
  NOR2_X1 U15861 ( .A1(n20902), .A2(n21000), .ZN(n18887) );
  NAND2_X1 U15862 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18887), .ZN(
        n18874) );
  NOR2_X1 U15863 ( .A1(n14118), .A2(n18874), .ZN(n18852) );
  NOR2_X1 U15864 ( .A1(n14119), .A2(n20902), .ZN(n21053) );
  INV_X1 U15865 ( .A(n21053), .ZN(n18626) );
  OAI21_X1 U15866 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18852), .A(
        n18626), .ZN(n21043) );
  OAI22_X1 U15867 ( .A1(n18830), .A2(n14120), .B1(n18955), .B2(n21043), .ZN(
        n14126) );
  NAND2_X1 U15868 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21668) );
  NOR3_X1 U15869 ( .A1(n18845), .A2(n21668), .A3(n14121), .ZN(n18848) );
  INV_X1 U15870 ( .A(n21675), .ZN(n21671) );
  NAND2_X1 U15871 ( .A1(n14122), .A2(n21656), .ZN(n18867) );
  NOR2_X1 U15872 ( .A1(n18858), .A2(n18867), .ZN(n18601) );
  AOI21_X1 U15873 ( .B1(n18848), .B2(n21671), .A(n18601), .ZN(n14123) );
  XOR2_X1 U15874 ( .A(n14123), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n21679) );
  NOR2_X2 U15875 ( .A1(n11148), .A2(n18973), .ZN(n18870) );
  AOI22_X1 U15876 ( .A1(n18962), .A2(n21670), .B1(n18883), .B2(n21870), .ZN(
        n18873) );
  OAI22_X1 U15877 ( .A1(n21679), .A2(n18881), .B1(n18873), .B2(n18622), .ZN(
        n14125) );
  OR4_X1 U15878 ( .A1(n14128), .A2(n14127), .A3(n14126), .A4(n14125), .ZN(
        P3_U2819) );
  OR2_X1 U15879 ( .A1(n21537), .A2(n18969), .ZN(n20831) );
  NOR2_X1 U15880 ( .A1(n22363), .A2(n20831), .ZN(n21950) );
  NOR4_X1 U15881 ( .A1(n21537), .A2(n21960), .A3(n22363), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n17948) );
  INV_X1 U15882 ( .A(n14130), .ZN(n18569) );
  NOR3_X1 U15883 ( .A1(n17951), .A2(n14131), .A3(n18569), .ZN(n21962) );
  AOI221_X1 U15884 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n21962), .C1(
        P3_MORE_REG_SCAN_IN), .C2(n21962), .A(n14132), .ZN(n14175) );
  OR2_X1 U15885 ( .A1(n20834), .A2(n14133), .ZN(n17952) );
  AOI211_X1 U15886 ( .C1(n21340), .C2(n17952), .A(n17951), .B(n22367), .ZN(
        n14135) );
  AOI211_X1 U15887 ( .C1(n14490), .C2(n14489), .A(n14135), .B(n14134), .ZN(
        n16260) );
  AOI22_X1 U15888 ( .A1(n17951), .A2(n17953), .B1(n14137), .B2(n14136), .ZN(
        n14138) );
  OAI221_X1 U15889 ( .B1(n14490), .B2(n21911), .C1(n14490), .C2(n21847), .A(
        n14138), .ZN(n21963) );
  OAI22_X1 U15890 ( .A1(n14142), .A2(n14141), .B1(n14140), .B2(n14139), .ZN(
        n14152) );
  AOI21_X1 U15891 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14155), .A(
        n21559), .ZN(n20933) );
  NAND2_X1 U15892 ( .A1(n21550), .A2(n21549), .ZN(n14150) );
  XOR2_X1 U15893 ( .A(n21559), .B(n14150), .Z(n14143) );
  OAI22_X1 U15894 ( .A1(n14145), .A2(n14144), .B1(n21911), .B2(n14143), .ZN(
        n14149) );
  OAI21_X1 U15895 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21746), .A(
        n21883), .ZN(n14160) );
  OAI33_X1 U15896 ( .A1(n14155), .A2(n14147), .A3(n21559), .B1(n14146), .B2(
        n14160), .B3(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14148) );
  AOI211_X1 U15897 ( .C1(n14152), .C2(n20933), .A(n14149), .B(n14148), .ZN(
        n21553) );
  INV_X1 U15898 ( .A(n16260), .ZN(n14158) );
  MUX2_X1 U15899 ( .A(n21559), .B(n21553), .S(n14158), .Z(n14169) );
  NAND2_X1 U15900 ( .A1(n14151), .A2(n14150), .ZN(n20914) );
  NAND2_X1 U15901 ( .A1(n21541), .A2(n21550), .ZN(n14157) );
  OAI211_X1 U15902 ( .C1(n14153), .C2(n14152), .A(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n21549), .ZN(n14154) );
  OAI21_X1 U15903 ( .B1(n14155), .B2(n14160), .A(n14154), .ZN(n14156) );
  AOI22_X1 U15904 ( .A1(n21875), .A2(n20914), .B1(n14157), .B2(n14156), .ZN(
        n21546) );
  AOI22_X1 U15905 ( .A1(n16260), .A2(n21550), .B1(n21546), .B2(n14158), .ZN(
        n14166) );
  AND2_X1 U15906 ( .A1(n21345), .A2(n21925), .ZN(n14161) );
  AOI22_X1 U15907 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21936), .B1(
        n14161), .B2(n21535), .ZN(n21533) );
  NAND2_X1 U15908 ( .A1(n14159), .A2(n21549), .ZN(n20898) );
  OAI22_X1 U15909 ( .A1(n14161), .A2(n20898), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n14160), .ZN(n21539) );
  OR3_X1 U15910 ( .A1(n21533), .A2(n19524), .A3(n19530), .ZN(n14162) );
  AOI22_X1 U15911 ( .A1(n21533), .A2(n19524), .B1(n21539), .B2(n14162), .ZN(
        n14163) );
  NAND2_X1 U15912 ( .A1(n19524), .A2(n19530), .ZN(n19542) );
  OAI21_X1 U15913 ( .B1(n16260), .B2(n14163), .A(n19542), .ZN(n14165) );
  AND2_X1 U15914 ( .A1(n14166), .A2(n14165), .ZN(n14164) );
  OAI221_X1 U15915 ( .B1(n14166), .B2(n14165), .C1(n19523), .C2(n14164), .A(
        n17950), .ZN(n14168) );
  INV_X1 U15916 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19522) );
  AOI21_X1 U15917 ( .B1(n17950), .B2(n19522), .A(n14166), .ZN(n14167) );
  AOI222_X1 U15918 ( .A1(n14169), .A2(n14168), .B1(n14169), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n14168), .C2(n14167), .ZN(
        n14170) );
  OAI21_X1 U15919 ( .B1(n14172), .B2(n21541), .A(n14171), .ZN(n17934) );
  NAND2_X1 U15920 ( .A1(n14173), .A2(n17934), .ZN(n16259) );
  NAND3_X1 U15921 ( .A1(n14175), .A2(n14174), .A3(n16259), .ZN(n21955) );
  AOI211_X1 U15922 ( .C1(n20834), .C2(n21337), .A(n22367), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n20906) );
  NAND2_X1 U15923 ( .A1(n20841), .A2(n20906), .ZN(n14176) );
  NAND2_X1 U15924 ( .A1(n14176), .A2(n21956), .ZN(n14177) );
  AOI21_X1 U15925 ( .B1(n21858), .B2(n22367), .A(n21944), .ZN(n21959) );
  NOR2_X1 U15926 ( .A1(n21949), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n20894) );
  INV_X1 U15927 ( .A(n20894), .ZN(n19555) );
  AND3_X1 U15928 ( .A1(n20895), .A2(n21959), .A3(n19555), .ZN(n14178) );
  OR2_X1 U15929 ( .A1(n11846), .A2(n19448), .ZN(n14179) );
  NOR2_X1 U15930 ( .A1(n15158), .A2(n14179), .ZN(n19110) );
  INV_X1 U15931 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n14180) );
  OAI211_X1 U15932 ( .C1(n19110), .C2(n14180), .A(n18027), .B(n14198), .ZN(
        P2_U2814) );
  NOR2_X1 U15933 ( .A1(n19074), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n14182)
         );
  AOI22_X1 U15934 ( .A1(n14182), .A2(n18027), .B1(n14181), .B2(n19074), .ZN(
        P2_U3612) );
  INV_X1 U15935 ( .A(n14584), .ZN(n14186) );
  INV_X1 U15936 ( .A(n14184), .ZN(n14185) );
  OAI21_X1 U15937 ( .B1(n16719), .B2(n14186), .A(n14185), .ZN(n14187) );
  NOR2_X1 U15938 ( .A1(n16724), .A2(n16320), .ZN(n14190) );
  INV_X1 U15939 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n14188) );
  NAND2_X1 U15940 ( .A1(n22424), .A2(n14188), .ZN(n22468) );
  NOR2_X1 U15941 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n22468), .ZN(n22810) );
  OAI21_X1 U15942 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(n22810), .A(n21967), 
        .ZN(n14189) );
  OAI21_X1 U15943 ( .B1(n21967), .B2(n14190), .A(n14189), .ZN(P1_U3487) );
  OR2_X1 U15944 ( .A1(n14191), .A2(n12947), .ZN(n14587) );
  INV_X1 U15945 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n14956) );
  MUX2_X1 U15946 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n14775), .Z(
        n16858) );
  NAND2_X1 U15947 ( .A1(n14357), .A2(n16858), .ZN(n22375) );
  OAI21_X2 U15948 ( .B1(n15607), .B2(n22322), .A(n22811), .ZN(n22385) );
  NAND2_X1 U15949 ( .A1(n22385), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n14192) );
  OAI211_X1 U15950 ( .C1(n14587), .C2(n14956), .A(n22375), .B(n14192), .ZN(
        P1_U2946) );
  MUX2_X1 U15951 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n14775), .Z(
        n16267) );
  NAND2_X1 U15952 ( .A1(n14357), .A2(n16267), .ZN(n22379) );
  NAND2_X1 U15953 ( .A1(n22385), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n14193) );
  OAI211_X1 U15954 ( .C1(n14587), .C2(n14958), .A(n22379), .B(n14193), .ZN(
        P1_U2949) );
  INV_X1 U15955 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14954) );
  MUX2_X1 U15956 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n14775), .Z(
        n16847) );
  NAND2_X1 U15957 ( .A1(n14357), .A2(n16847), .ZN(n22382) );
  NAND2_X1 U15958 ( .A1(n22385), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n14194) );
  OAI211_X1 U15959 ( .C1(n14587), .C2(n14954), .A(n22382), .B(n14194), .ZN(
        P1_U2950) );
  INV_X1 U15960 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14962) );
  MUX2_X1 U15961 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n14775), .Z(
        n16851) );
  NAND2_X1 U15962 ( .A1(n14357), .A2(n16851), .ZN(n22377) );
  NAND2_X1 U15963 ( .A1(n22385), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n14195) );
  OAI211_X1 U15964 ( .C1(n14587), .C2(n14962), .A(n22377), .B(n14195), .ZN(
        P1_U2948) );
  INV_X1 U15965 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14952) );
  MUX2_X1 U15966 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n14775), .Z(
        n16843) );
  NAND2_X1 U15967 ( .A1(n14357), .A2(n16843), .ZN(n22386) );
  NAND2_X1 U15968 ( .A1(n22385), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n14196) );
  OAI211_X1 U15969 ( .C1(n14952), .C2(n14587), .A(n22386), .B(n14196), .ZN(
        P1_U2951) );
  INV_X1 U15970 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20619) );
  MUX2_X1 U15971 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n14775), .Z(
        n16862) );
  NAND2_X1 U15972 ( .A1(n14357), .A2(n16862), .ZN(n14346) );
  NAND2_X1 U15973 ( .A1(n22385), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n14197) );
  OAI211_X1 U15974 ( .C1(n20619), .C2(n14587), .A(n14346), .B(n14197), .ZN(
        P1_U2960) );
  OAI21_X2 U15975 ( .B1(n22338), .B2(n14198), .A(n14418), .ZN(n14394) );
  INV_X1 U15976 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n14201) );
  NAND3_X1 U15977 ( .A1(n14199), .A2(n19079), .A3(n19073), .ZN(n14536) );
  MUX2_X1 U15978 ( .A(BUF1_REG_9__SCAN_IN), .B(BUF2_REG_9__SCAN_IN), .S(n16030), .Z(n17452) );
  INV_X1 U15979 ( .A(n17452), .ZN(n14670) );
  NOR2_X1 U15980 ( .A1(n14536), .A2(n14670), .ZN(n14207) );
  AOI21_X1 U15981 ( .B1(n14549), .B2(P2_EAX_REG_9__SCAN_IN), .A(n14207), .ZN(
        n14200) );
  OAI21_X1 U15982 ( .B1(n14394), .B2(n14201), .A(n14200), .ZN(P2_U2976) );
  INV_X1 U15983 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n14206) );
  INV_X1 U15984 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n14202) );
  OR2_X1 U15985 ( .A1(n16030), .A2(n14202), .ZN(n14204) );
  NAND2_X1 U15986 ( .A1(n16030), .A2(BUF2_REG_4__SCAN_IN), .ZN(n14203) );
  AND2_X1 U15987 ( .A1(n14204), .A2(n14203), .ZN(n20230) );
  NOR2_X1 U15988 ( .A1(n14536), .A2(n20230), .ZN(n14545) );
  AOI21_X1 U15989 ( .B1(n14549), .B2(P2_EAX_REG_20__SCAN_IN), .A(n14545), .ZN(
        n14205) );
  OAI21_X1 U15990 ( .B1(n14394), .B2(n14206), .A(n14205), .ZN(P2_U2956) );
  INV_X1 U15991 ( .A(P2_UWORD_REG_9__SCAN_IN), .ZN(n14209) );
  AOI21_X1 U15992 ( .B1(n14549), .B2(P2_EAX_REG_25__SCAN_IN), .A(n14207), .ZN(
        n14208) );
  OAI21_X1 U15993 ( .B1(n14394), .B2(n14209), .A(n14208), .ZN(P2_U2961) );
  INV_X1 U15994 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14214) );
  INV_X1 U15995 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n14213) );
  INV_X1 U15996 ( .A(n22385), .ZN(n14328) );
  INV_X1 U15997 ( .A(DATAI_15_), .ZN(n14210) );
  NOR2_X1 U15998 ( .A1(n14775), .A2(n14210), .ZN(n14211) );
  AOI21_X1 U15999 ( .B1(n14775), .B2(BUF1_REG_15__SCAN_IN), .A(n14211), .ZN(
        n16055) );
  OAI222_X1 U16000 ( .A1(n14587), .A2(n14214), .B1(n14213), .B2(n14328), .C1(
        n14212), .C2(n16055), .ZN(P1_U2967) );
  INV_X1 U16001 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n14219) );
  INV_X1 U16002 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n14215) );
  OR2_X1 U16003 ( .A1(n16030), .A2(n14215), .ZN(n14217) );
  NAND2_X1 U16004 ( .A1(n16030), .A2(BUF2_REG_6__SCAN_IN), .ZN(n14216) );
  AND2_X1 U16005 ( .A1(n14217), .A2(n14216), .ZN(n20114) );
  INV_X1 U16006 ( .A(n20114), .ZN(n17471) );
  NAND2_X1 U16007 ( .A1(n14413), .A2(n17471), .ZN(n14409) );
  NAND2_X1 U16008 ( .A1(n14549), .A2(P2_EAX_REG_6__SCAN_IN), .ZN(n14218) );
  OAI211_X1 U16009 ( .C1(n14394), .C2(n14219), .A(n14409), .B(n14218), .ZN(
        P2_U2973) );
  INV_X1 U16010 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n14224) );
  INV_X1 U16011 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n14220) );
  OR2_X1 U16012 ( .A1(n16030), .A2(n14220), .ZN(n14222) );
  NAND2_X1 U16013 ( .A1(n16030), .A2(BUF2_REG_5__SCAN_IN), .ZN(n14221) );
  AND2_X1 U16014 ( .A1(n14222), .A2(n14221), .ZN(n20172) );
  INV_X1 U16015 ( .A(n20172), .ZN(n20163) );
  NAND2_X1 U16016 ( .A1(n14413), .A2(n20163), .ZN(n14405) );
  NAND2_X1 U16017 ( .A1(n14549), .A2(P2_EAX_REG_5__SCAN_IN), .ZN(n14223) );
  OAI211_X1 U16018 ( .C1(n14394), .C2(n14224), .A(n14405), .B(n14223), .ZN(
        P2_U2972) );
  INV_X1 U16019 ( .A(P2_LWORD_REG_10__SCAN_IN), .ZN(n14226) );
  MUX2_X1 U16020 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n16030), .Z(n17444) );
  NAND2_X1 U16021 ( .A1(n14413), .A2(n17444), .ZN(n14395) );
  NAND2_X1 U16022 ( .A1(n14549), .A2(P2_EAX_REG_10__SCAN_IN), .ZN(n14225) );
  OAI211_X1 U16023 ( .C1(n14394), .C2(n14226), .A(n14395), .B(n14225), .ZN(
        P2_U2977) );
  INV_X1 U16024 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n14228) );
  MUX2_X1 U16025 ( .A(BUF1_REG_11__SCAN_IN), .B(BUF2_REG_11__SCAN_IN), .S(
        n16030), .Z(n17437) );
  NAND2_X1 U16026 ( .A1(n14413), .A2(n17437), .ZN(n14400) );
  NAND2_X1 U16027 ( .A1(n14549), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n14227) );
  OAI211_X1 U16028 ( .C1(n14394), .C2(n14228), .A(n14400), .B(n14227), .ZN(
        P2_U2978) );
  INV_X1 U16029 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n14230) );
  MUX2_X1 U16030 ( .A(BUF1_REG_13__SCAN_IN), .B(BUF2_REG_13__SCAN_IN), .S(
        n16030), .Z(n16654) );
  NAND2_X1 U16031 ( .A1(n14413), .A2(n16654), .ZN(n14411) );
  NAND2_X1 U16032 ( .A1(n14549), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n14229) );
  OAI211_X1 U16033 ( .C1(n14394), .C2(n14230), .A(n14411), .B(n14229), .ZN(
        P2_U2980) );
  INV_X1 U16034 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n14232) );
  MUX2_X1 U16035 ( .A(BUF1_REG_8__SCAN_IN), .B(BUF2_REG_8__SCAN_IN), .S(n16030), .Z(n17459) );
  NAND2_X1 U16036 ( .A1(n14413), .A2(n17459), .ZN(n14407) );
  NAND2_X1 U16037 ( .A1(n14549), .A2(P2_EAX_REG_8__SCAN_IN), .ZN(n14231) );
  OAI211_X1 U16038 ( .C1(n14394), .C2(n14232), .A(n14407), .B(n14231), .ZN(
        P2_U2975) );
  INV_X1 U16039 ( .A(P2_LWORD_REG_12__SCAN_IN), .ZN(n14234) );
  MUX2_X1 U16040 ( .A(BUF1_REG_12__SCAN_IN), .B(BUF2_REG_12__SCAN_IN), .S(
        n16030), .Z(n17431) );
  NAND2_X1 U16041 ( .A1(n14413), .A2(n17431), .ZN(n14402) );
  NAND2_X1 U16042 ( .A1(n14549), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n14233) );
  OAI211_X1 U16043 ( .C1(n14394), .C2(n14234), .A(n14402), .B(n14233), .ZN(
        P2_U2979) );
  INV_X1 U16044 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n14239) );
  INV_X1 U16045 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n14235) );
  OR2_X1 U16046 ( .A1(n16030), .A2(n14235), .ZN(n14237) );
  NAND2_X1 U16047 ( .A1(n16030), .A2(BUF2_REG_7__SCAN_IN), .ZN(n14236) );
  AND2_X1 U16048 ( .A1(n14237), .A2(n14236), .ZN(n19919) );
  INV_X1 U16049 ( .A(n19919), .ZN(n17464) );
  NAND2_X1 U16050 ( .A1(n14413), .A2(n17464), .ZN(n14398) );
  NAND2_X1 U16051 ( .A1(n14549), .A2(P2_EAX_REG_7__SCAN_IN), .ZN(n14238) );
  OAI211_X1 U16052 ( .C1(n14394), .C2(n14239), .A(n14398), .B(n14238), .ZN(
        P2_U2974) );
  INV_X1 U16053 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n14242) );
  INV_X1 U16054 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n14240) );
  NOR2_X1 U16055 ( .A1(n16139), .A2(n14240), .ZN(n14241) );
  AOI21_X1 U16056 ( .B1(BUF1_REG_15__SCAN_IN), .B2(n16139), .A(n14241), .ZN(
        n15318) );
  INV_X1 U16057 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n18183) );
  OAI222_X1 U16058 ( .A1(n14394), .A2(n14242), .B1(n14536), .B2(n15318), .C1(
        n14418), .C2(n18183), .ZN(P2_U2982) );
  OAI222_X1 U16059 ( .A1(n14249), .A2(n14246), .B1(n14249), .B2(n14245), .C1(
        n14244), .C2(n14243), .ZN(n14475) );
  AOI21_X1 U16060 ( .B1(n14249), .B2(n14248), .A(n14247), .ZN(n14472) );
  INV_X1 U16061 ( .A(n14472), .ZN(n14250) );
  NAND2_X1 U16062 ( .A1(n19407), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n14476) );
  OAI21_X1 U16063 ( .B1(n18103), .B2(n14250), .A(n14476), .ZN(n14252) );
  MUX2_X1 U16064 ( .A(n18070), .B(n18102), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n14251) );
  AOI211_X1 U16065 ( .C1(n14475), .C2(n18079), .A(n14252), .B(n14251), .ZN(
        n14253) );
  OAI21_X1 U16066 ( .B1(n14664), .B2(n18105), .A(n14253), .ZN(P2_U3013) );
  AOI22_X1 U16067 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n22385), .B1(n22384), 
        .B2(P1_EAX_REG_18__SCAN_IN), .ZN(n14256) );
  INV_X1 U16068 ( .A(n14775), .ZN(n14354) );
  NAND2_X1 U16069 ( .A1(n14354), .A2(DATAI_2_), .ZN(n14255) );
  NAND2_X1 U16070 ( .A1(n14775), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14254) );
  AND2_X1 U16071 ( .A1(n14255), .A2(n14254), .ZN(n14894) );
  INV_X1 U16072 ( .A(n14894), .ZN(n16885) );
  NAND2_X1 U16073 ( .A1(n14357), .A2(n16885), .ZN(n14329) );
  NAND2_X1 U16074 ( .A1(n14256), .A2(n14329), .ZN(P1_U2939) );
  AOI22_X1 U16075 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n22385), .B1(n22384), 
        .B2(P1_EAX_REG_16__SCAN_IN), .ZN(n14259) );
  NAND2_X1 U16076 ( .A1(n14354), .A2(DATAI_0_), .ZN(n14258) );
  NAND2_X1 U16077 ( .A1(n14775), .A2(BUF1_REG_0__SCAN_IN), .ZN(n14257) );
  AND2_X1 U16078 ( .A1(n14258), .A2(n14257), .ZN(n14806) );
  INV_X1 U16079 ( .A(n14806), .ZN(n16152) );
  NAND2_X1 U16080 ( .A1(n14357), .A2(n16152), .ZN(n14331) );
  NAND2_X1 U16081 ( .A1(n14259), .A2(n14331), .ZN(P1_U2937) );
  AOI22_X1 U16082 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n22385), .B1(n22384), 
        .B2(P1_EAX_REG_19__SCAN_IN), .ZN(n14262) );
  NAND2_X1 U16083 ( .A1(n14354), .A2(DATAI_3_), .ZN(n14261) );
  NAND2_X1 U16084 ( .A1(n14775), .A2(BUF1_REG_3__SCAN_IN), .ZN(n14260) );
  AND2_X1 U16085 ( .A1(n14261), .A2(n14260), .ZN(n14869) );
  INV_X1 U16086 ( .A(n14869), .ZN(n16881) );
  NAND2_X1 U16087 ( .A1(n14357), .A2(n16881), .ZN(n14263) );
  NAND2_X1 U16088 ( .A1(n14262), .A2(n14263), .ZN(P1_U2940) );
  AOI22_X1 U16089 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n22385), .B1(n22384), 
        .B2(P1_EAX_REG_3__SCAN_IN), .ZN(n14264) );
  NAND2_X1 U16090 ( .A1(n14264), .A2(n14263), .ZN(P1_U2955) );
  INV_X1 U16091 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14269) );
  NOR2_X1 U16092 ( .A1(n11846), .A2(n12188), .ZN(n14265) );
  NAND2_X1 U16093 ( .A1(n16020), .A2(n14265), .ZN(n15102) );
  OAI21_X1 U16094 ( .B1(n15102), .B2(n19448), .A(n14418), .ZN(n14266) );
  NAND2_X1 U16095 ( .A1(n18147), .A2(n14267), .ZN(n14662) );
  NOR2_X1 U16096 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18114), .ZN(n18168) );
  AOI22_X1 U16097 ( .A1(n18180), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n18159), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n14268) );
  OAI21_X1 U16098 ( .B1(n14269), .B2(n14662), .A(n14268), .ZN(P2_U2930) );
  INV_X1 U16099 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14271) );
  AOI22_X1 U16100 ( .A1(n18180), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n18159), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n14270) );
  OAI21_X1 U16101 ( .B1(n14271), .B2(n14662), .A(n14270), .ZN(P2_U2929) );
  INV_X1 U16102 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14273) );
  AOI22_X1 U16103 ( .A1(n18168), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n18159), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n14272) );
  OAI21_X1 U16104 ( .B1(n14273), .B2(n14662), .A(n14272), .ZN(P2_U2932) );
  INV_X1 U16105 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n14275) );
  AOI22_X1 U16106 ( .A1(n18180), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n18159), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n14274) );
  OAI21_X1 U16107 ( .B1(n14275), .B2(n14662), .A(n14274), .ZN(P2_U2928) );
  INV_X1 U16108 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n14277) );
  AOI22_X1 U16109 ( .A1(n18180), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n18159), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n14276) );
  OAI21_X1 U16110 ( .B1(n14277), .B2(n14662), .A(n14276), .ZN(P2_U2927) );
  INV_X1 U16111 ( .A(n16715), .ZN(n16721) );
  INV_X1 U16112 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n22335) );
  NAND2_X1 U16113 ( .A1(n14278), .A2(n22335), .ZN(n22331) );
  INV_X1 U16114 ( .A(n22322), .ZN(n22330) );
  AOI21_X1 U16115 ( .B1(n12947), .B2(n22331), .A(n22330), .ZN(n14279) );
  NAND2_X1 U16116 ( .A1(n16721), .A2(n14279), .ZN(n14286) );
  INV_X1 U16117 ( .A(n22331), .ZN(n14448) );
  OAI21_X1 U16118 ( .B1(n12947), .B2(n14448), .A(n22322), .ZN(n15073) );
  INV_X1 U16119 ( .A(n15073), .ZN(n14282) );
  NAND2_X1 U16120 ( .A1(n12948), .A2(n16710), .ZN(n14281) );
  AOI21_X1 U16121 ( .B1(n14280), .B2(n14282), .A(n14281), .ZN(n14283) );
  OR2_X1 U16122 ( .A1(n16719), .A2(n14283), .ZN(n14285) );
  MUX2_X1 U16123 ( .A(n14286), .B(n14285), .S(n14284), .Z(n14294) );
  INV_X1 U16124 ( .A(n14287), .ZN(n14292) );
  OR2_X1 U16125 ( .A1(n14310), .A2(n12957), .ZN(n14288) );
  AND2_X1 U16126 ( .A1(n14289), .A2(n14288), .ZN(n14301) );
  NAND2_X1 U16127 ( .A1(n14462), .A2(n14319), .ZN(n14290) );
  AND3_X1 U16128 ( .A1(n14301), .A2(n12940), .A3(n14290), .ZN(n14312) );
  OAI21_X1 U16129 ( .B1(n16722), .B2(n14312), .A(n14291), .ZN(n14453) );
  AOI21_X1 U16130 ( .B1(n16719), .B2(n14292), .A(n14453), .ZN(n14293) );
  NAND2_X1 U16131 ( .A1(n14294), .A2(n14293), .ZN(n14295) );
  OAI22_X1 U16132 ( .A1(n13689), .A2(n12947), .B1(n14315), .B2(n14882), .ZN(
        n14296) );
  INV_X1 U16133 ( .A(n14797), .ZN(n14297) );
  MUX2_X1 U16134 ( .A(n16321), .B(n14857), .S(P1_EBX_REG_0__SCAN_IN), .Z(
        n14649) );
  OR2_X1 U16135 ( .A1(n16323), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14298) );
  NAND2_X1 U16136 ( .A1(n14649), .A2(n14298), .ZN(n15181) );
  INV_X1 U16137 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21986) );
  AND2_X1 U16138 ( .A1(n14436), .A2(n11192), .ZN(n16709) );
  NAND2_X1 U16139 ( .A1(n14318), .A2(n16709), .ZN(n21999) );
  AOI21_X1 U16140 ( .B1(n12933), .B2(n12886), .A(n16150), .ZN(n14300) );
  INV_X1 U16141 ( .A(n15070), .ZN(n14435) );
  OAI21_X1 U16142 ( .B1(n12946), .B2(n14310), .A(n14435), .ZN(n14299) );
  OAI211_X1 U16143 ( .C1(n14301), .C2(n16385), .A(n14300), .B(n14299), .ZN(
        n14302) );
  INV_X1 U16144 ( .A(n14302), .ZN(n14304) );
  NAND2_X1 U16145 ( .A1(n12962), .A2(n16724), .ZN(n14303) );
  AND3_X1 U16146 ( .A1(n14305), .A2(n14304), .A3(n14303), .ZN(n14432) );
  OAI211_X1 U16147 ( .C1(n14428), .C2(n16710), .A(n14432), .B(n14306), .ZN(
        n14307) );
  NAND2_X1 U16148 ( .A1(n14318), .A2(n14307), .ZN(n15301) );
  NAND2_X1 U16149 ( .A1(n21999), .A2(n15301), .ZN(n14308) );
  OR2_X1 U16150 ( .A1(n14629), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22066) );
  INV_X1 U16151 ( .A(n22066), .ZN(n22021) );
  NOR2_X1 U16152 ( .A1(n14318), .A2(n22021), .ZN(n15298) );
  AOI21_X1 U16153 ( .B1(n21986), .B2(n14308), .A(n15298), .ZN(n22088) );
  INV_X1 U16154 ( .A(n22088), .ZN(n14309) );
  NAND2_X1 U16155 ( .A1(n14318), .A2(n14584), .ZN(n15303) );
  INV_X1 U16156 ( .A(n15303), .ZN(n22079) );
  OAI22_X1 U16157 ( .A1(n14309), .A2(n22079), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n14308), .ZN(n14327) );
  INV_X1 U16158 ( .A(n14310), .ZN(n14311) );
  NAND2_X1 U16159 ( .A1(n14312), .A2(n14311), .ZN(n14628) );
  AND2_X1 U16160 ( .A1(n14628), .A2(n14313), .ZN(n16713) );
  OR2_X1 U16161 ( .A1(n13689), .A2(n12949), .ZN(n14449) );
  OR2_X1 U16162 ( .A1(n14315), .A2(n14314), .ZN(n14316) );
  NAND4_X1 U16163 ( .A1(n13678), .A2(n16713), .A3(n14449), .A4(n14316), .ZN(
        n14317) );
  NAND2_X1 U16164 ( .A1(n22280), .A2(n15602), .ZN(n14322) );
  INV_X1 U16165 ( .A(n15607), .ZN(n21971) );
  NAND2_X1 U16166 ( .A1(n14319), .A2(n14797), .ZN(n14695) );
  OAI21_X1 U16167 ( .B1(n21971), .B2(n14636), .A(n14695), .ZN(n14320) );
  INV_X1 U16168 ( .A(n14320), .ZN(n14321) );
  NAND2_X1 U16169 ( .A1(n14322), .A2(n14321), .ZN(n14323) );
  NAND2_X1 U16170 ( .A1(n14323), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14690) );
  OR2_X1 U16171 ( .A1(n14323), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14324) );
  NAND2_X1 U16172 ( .A1(n14690), .A2(n14324), .ZN(n20735) );
  INV_X1 U16173 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n20696) );
  OAI22_X1 U16174 ( .A1(n22058), .A2(n20735), .B1(n20696), .B2(n22066), .ZN(
        n14325) );
  INV_X1 U16175 ( .A(n14325), .ZN(n14326) );
  OAI211_X1 U16176 ( .C1(n22082), .C2(n15181), .A(n14327), .B(n14326), .ZN(
        P1_U3031) );
  AOI22_X1 U16177 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n22381), .B1(n22384), 
        .B2(P1_EAX_REG_2__SCAN_IN), .ZN(n14330) );
  NAND2_X1 U16178 ( .A1(n14330), .A2(n14329), .ZN(P1_U2954) );
  AOI22_X1 U16179 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n22381), .B1(n22384), 
        .B2(P1_EAX_REG_0__SCAN_IN), .ZN(n14332) );
  NAND2_X1 U16180 ( .A1(n14332), .A2(n14331), .ZN(P1_U2952) );
  AOI22_X1 U16181 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n22381), .B1(n22384), 
        .B2(P1_EAX_REG_7__SCAN_IN), .ZN(n14333) );
  MUX2_X1 U16182 ( .A(DATAI_7_), .B(BUF1_REG_7__SCAN_IN), .S(n14775), .Z(
        n16865) );
  NAND2_X1 U16183 ( .A1(n14357), .A2(n16865), .ZN(n14335) );
  NAND2_X1 U16184 ( .A1(n14333), .A2(n14335), .ZN(P1_U2959) );
  AOI22_X1 U16185 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n22381), .B1(n22384), 
        .B2(P1_EAX_REG_26__SCAN_IN), .ZN(n14334) );
  MUX2_X1 U16186 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n14775), .Z(
        n16855) );
  NAND2_X1 U16187 ( .A1(n14357), .A2(n16855), .ZN(n14350) );
  NAND2_X1 U16188 ( .A1(n14334), .A2(n14350), .ZN(P1_U2947) );
  AOI22_X1 U16189 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n22381), .B1(n22384), 
        .B2(P1_EAX_REG_23__SCAN_IN), .ZN(n14336) );
  NAND2_X1 U16190 ( .A1(n14336), .A2(n14335), .ZN(P1_U2944) );
  AOI22_X1 U16191 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n22381), .B1(n22384), 
        .B2(P1_EAX_REG_1__SCAN_IN), .ZN(n14339) );
  NAND2_X1 U16192 ( .A1(n14354), .A2(DATAI_1_), .ZN(n14338) );
  NAND2_X1 U16193 ( .A1(n14775), .A2(BUF1_REG_1__SCAN_IN), .ZN(n14337) );
  AND2_X1 U16194 ( .A1(n14338), .A2(n14337), .ZN(n14914) );
  INV_X1 U16195 ( .A(n14914), .ZN(n16893) );
  NAND2_X1 U16196 ( .A1(n14357), .A2(n16893), .ZN(n14361) );
  NAND2_X1 U16197 ( .A1(n14339), .A2(n14361), .ZN(P1_U2953) );
  AOI22_X1 U16198 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n22381), .B1(n22384), 
        .B2(P1_EAX_REG_4__SCAN_IN), .ZN(n14342) );
  NAND2_X1 U16199 ( .A1(n14354), .A2(DATAI_4_), .ZN(n14341) );
  NAND2_X1 U16200 ( .A1(n14775), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14340) );
  AND2_X1 U16201 ( .A1(n14341), .A2(n14340), .ZN(n14881) );
  INV_X1 U16202 ( .A(n14881), .ZN(n16878) );
  NAND2_X1 U16203 ( .A1(n14357), .A2(n16878), .ZN(n14348) );
  NAND2_X1 U16204 ( .A1(n14342), .A2(n14348), .ZN(P1_U2956) );
  AOI22_X1 U16205 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n22381), .B1(n22384), 
        .B2(P1_EAX_REG_21__SCAN_IN), .ZN(n14345) );
  NAND2_X1 U16206 ( .A1(n14354), .A2(DATAI_5_), .ZN(n14344) );
  NAND2_X1 U16207 ( .A1(n14775), .A2(BUF1_REG_5__SCAN_IN), .ZN(n14343) );
  AND2_X1 U16208 ( .A1(n14344), .A2(n14343), .ZN(n14985) );
  INV_X1 U16209 ( .A(n14985), .ZN(n16874) );
  NAND2_X1 U16210 ( .A1(n14357), .A2(n16874), .ZN(n14352) );
  NAND2_X1 U16211 ( .A1(n14345), .A2(n14352), .ZN(P1_U2942) );
  AOI22_X1 U16212 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n22381), .B1(n22384), 
        .B2(P1_EAX_REG_24__SCAN_IN), .ZN(n14347) );
  NAND2_X1 U16213 ( .A1(n14347), .A2(n14346), .ZN(P1_U2945) );
  AOI22_X1 U16214 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n22381), .B1(n22384), 
        .B2(P1_EAX_REG_20__SCAN_IN), .ZN(n14349) );
  NAND2_X1 U16215 ( .A1(n14349), .A2(n14348), .ZN(P1_U2941) );
  AOI22_X1 U16216 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n22381), .B1(n22384), 
        .B2(P1_EAX_REG_10__SCAN_IN), .ZN(n14351) );
  NAND2_X1 U16217 ( .A1(n14351), .A2(n14350), .ZN(P1_U2962) );
  AOI22_X1 U16218 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n22381), .B1(n22384), 
        .B2(P1_EAX_REG_5__SCAN_IN), .ZN(n14353) );
  NAND2_X1 U16219 ( .A1(n14353), .A2(n14352), .ZN(P1_U2957) );
  AOI22_X1 U16220 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n22381), .B1(n22384), 
        .B2(P1_EAX_REG_22__SCAN_IN), .ZN(n14358) );
  NAND2_X1 U16221 ( .A1(n14354), .A2(DATAI_6_), .ZN(n14356) );
  NAND2_X1 U16222 ( .A1(n14775), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14355) );
  AND2_X1 U16223 ( .A1(n14356), .A2(n14355), .ZN(n15283) );
  INV_X1 U16224 ( .A(n15283), .ZN(n16869) );
  NAND2_X1 U16225 ( .A1(n14357), .A2(n16869), .ZN(n14359) );
  NAND2_X1 U16226 ( .A1(n14358), .A2(n14359), .ZN(P1_U2943) );
  AOI22_X1 U16227 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n22381), .B1(n22384), 
        .B2(P1_EAX_REG_6__SCAN_IN), .ZN(n14360) );
  NAND2_X1 U16228 ( .A1(n14360), .A2(n14359), .ZN(P1_U2958) );
  AOI22_X1 U16229 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n22381), .B1(n22384), 
        .B2(P1_EAX_REG_17__SCAN_IN), .ZN(n14362) );
  NAND2_X1 U16230 ( .A1(n14362), .A2(n14361), .ZN(P1_U2938) );
  OAI21_X1 U16231 ( .B1(n14365), .B2(n14364), .A(n14363), .ZN(n20730) );
  NAND2_X1 U16232 ( .A1(n12909), .A2(n12941), .ZN(n14366) );
  INV_X2 U16233 ( .A(n15997), .ZN(n16897) );
  INV_X1 U16234 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20606) );
  OAI222_X1 U16235 ( .A1(n20730), .A2(n16897), .B1(n16056), .B2(n14806), .C1(
        n16054), .C2(n20606), .ZN(P1_U2904) );
  NAND2_X1 U16236 ( .A1(n16020), .A2(n14367), .ZN(n15108) );
  NAND2_X1 U16237 ( .A1(n15108), .A2(n14368), .ZN(n14369) );
  NAND2_X1 U16238 ( .A1(n14369), .A2(n19078), .ZN(n14372) );
  AND2_X1 U16239 ( .A1(n14370), .A2(n19073), .ZN(n15165) );
  NAND2_X1 U16240 ( .A1(n19074), .A2(n15165), .ZN(n14371) );
  NAND2_X1 U16241 ( .A1(n11649), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14373) );
  NAND2_X1 U16242 ( .A1(n14373), .A2(n20083), .ZN(n14709) );
  NOR2_X1 U16243 ( .A1(n20096), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n14374) );
  AOI21_X1 U16244 ( .B1(n14709), .B2(n19360), .A(n14374), .ZN(n14375) );
  INV_X1 U16245 ( .A(n14606), .ZN(n14379) );
  NOR2_X1 U16246 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14376) );
  NOR2_X1 U16247 ( .A1(n11649), .A2(n19436), .ZN(n14596) );
  OAI21_X1 U16248 ( .B1(n14377), .B2(n14376), .A(n14596), .ZN(n14378) );
  INV_X1 U16249 ( .A(n14380), .ZN(n14386) );
  INV_X1 U16250 ( .A(n14381), .ZN(n14384) );
  INV_X1 U16251 ( .A(n14382), .ZN(n14383) );
  NAND2_X1 U16252 ( .A1(n14384), .A2(n14383), .ZN(n14385) );
  NAND2_X1 U16253 ( .A1(n14386), .A2(n14385), .ZN(n19366) );
  XNOR2_X1 U16254 ( .A(n19929), .B(n19366), .ZN(n14393) );
  INV_X1 U16255 ( .A(n19921), .ZN(n14581) );
  NOR2_X1 U16256 ( .A1(n16141), .A2(n14387), .ZN(n20164) );
  INV_X1 U16257 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n14388) );
  OR2_X1 U16258 ( .A1(n16030), .A2(n14388), .ZN(n14390) );
  NAND2_X1 U16259 ( .A1(n16030), .A2(BUF2_REG_0__SCAN_IN), .ZN(n14389) );
  AND2_X1 U16260 ( .A1(n14390), .A2(n14389), .ZN(n20427) );
  INV_X1 U16261 ( .A(n20427), .ZN(n16178) );
  OR2_X1 U16262 ( .A1(n20319), .A2(n19921), .ZN(n17477) );
  OAI22_X1 U16263 ( .A1(n17477), .A2(n19366), .B1(n17475), .B2(n14417), .ZN(
        n14391) );
  AOI21_X1 U16264 ( .B1(n20164), .B2(n16178), .A(n14391), .ZN(n14392) );
  OAI21_X1 U16265 ( .B1(n20165), .B2(n14393), .A(n14392), .ZN(P2_U2919) );
  INV_X1 U16266 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14397) );
  NAND2_X1 U16267 ( .A1(n14522), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n14396) );
  OAI211_X1 U16268 ( .C1(n14418), .C2(n14397), .A(n14396), .B(n14395), .ZN(
        P2_U2962) );
  NAND2_X1 U16269 ( .A1(n14522), .A2(P2_UWORD_REG_7__SCAN_IN), .ZN(n14399) );
  OAI211_X1 U16270 ( .C1(n14418), .C2(n14275), .A(n14399), .B(n14398), .ZN(
        P2_U2959) );
  INV_X1 U16271 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n17435) );
  NAND2_X1 U16272 ( .A1(n14522), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n14401) );
  OAI211_X1 U16273 ( .C1(n14418), .C2(n17435), .A(n14401), .B(n14400), .ZN(
        P2_U2963) );
  INV_X1 U16274 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n17429) );
  NAND2_X1 U16275 ( .A1(n14522), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n14403) );
  OAI211_X1 U16276 ( .C1(n14418), .C2(n17429), .A(n14403), .B(n14402), .ZN(
        P2_U2964) );
  INV_X1 U16277 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n16174) );
  NAND2_X1 U16278 ( .A1(n14522), .A2(P2_UWORD_REG_0__SCAN_IN), .ZN(n14404) );
  NAND2_X1 U16279 ( .A1(n14413), .A2(n16178), .ZN(n14415) );
  OAI211_X1 U16280 ( .C1(n14418), .C2(n16174), .A(n14404), .B(n14415), .ZN(
        P2_U2952) );
  NAND2_X1 U16281 ( .A1(n14522), .A2(P2_UWORD_REG_5__SCAN_IN), .ZN(n14406) );
  OAI211_X1 U16282 ( .C1(n14418), .C2(n14269), .A(n14406), .B(n14405), .ZN(
        P2_U2957) );
  NAND2_X1 U16283 ( .A1(n14522), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n14408) );
  OAI211_X1 U16284 ( .C1(n14418), .C2(n14277), .A(n14408), .B(n14407), .ZN(
        P2_U2960) );
  NAND2_X1 U16285 ( .A1(n14522), .A2(P2_UWORD_REG_6__SCAN_IN), .ZN(n14410) );
  OAI211_X1 U16286 ( .C1(n14418), .C2(n14271), .A(n14410), .B(n14409), .ZN(
        P2_U2958) );
  INV_X1 U16287 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n16652) );
  NAND2_X1 U16288 ( .A1(n14522), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n14412) );
  OAI211_X1 U16289 ( .C1(n14418), .C2(n16652), .A(n14412), .B(n14411), .ZN(
        P2_U2965) );
  INV_X1 U16290 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n16689) );
  NAND2_X1 U16291 ( .A1(n14522), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n14414) );
  MUX2_X1 U16292 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n16030), .Z(n16691) );
  NAND2_X1 U16293 ( .A1(n14413), .A2(n16691), .ZN(n14553) );
  OAI211_X1 U16294 ( .C1(n14418), .C2(n16689), .A(n14414), .B(n14553), .ZN(
        P2_U2966) );
  NAND2_X1 U16295 ( .A1(n14522), .A2(P2_LWORD_REG_0__SCAN_IN), .ZN(n14416) );
  OAI211_X1 U16296 ( .C1(n14418), .C2(n14417), .A(n14416), .B(n14415), .ZN(
        P2_U2967) );
  NAND2_X1 U16297 ( .A1(n16719), .A2(n14436), .ZN(n14423) );
  INV_X1 U16298 ( .A(n14419), .ZN(n14420) );
  NAND2_X1 U16299 ( .A1(n14421), .A2(n14420), .ZN(n14422) );
  NAND2_X1 U16300 ( .A1(n14423), .A2(n14422), .ZN(n14425) );
  AND2_X1 U16301 ( .A1(n11192), .A2(n22807), .ZN(n14424) );
  INV_X1 U16302 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14426) );
  NAND2_X1 U16303 ( .A1(n20727), .A2(n12941), .ZN(n20698) );
  OAI222_X1 U16304 ( .A1(n15181), .A2(n16841), .B1(n14426), .B2(n20727), .C1(
        n20730), .C2(n20698), .ZN(P1_U2872) );
  NAND2_X1 U16305 ( .A1(n13687), .A2(n14428), .ZN(n14429) );
  NOR2_X1 U16306 ( .A1(n14280), .A2(n14429), .ZN(n14430) );
  AND2_X1 U16307 ( .A1(n13678), .A2(n14430), .ZN(n14431) );
  NAND2_X1 U16308 ( .A1(n14432), .A2(n14431), .ZN(n14480) );
  NAND2_X1 U16309 ( .A1(n14427), .A2(n14480), .ZN(n14446) );
  INV_X1 U16310 ( .A(n14508), .ZN(n14437) );
  INV_X1 U16311 ( .A(n14480), .ZN(n14514) );
  NAND2_X1 U16312 ( .A1(n14508), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14433) );
  NAND2_X1 U16313 ( .A1(n14433), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14434) );
  NAND2_X1 U16314 ( .A1(n11190), .A2(n14434), .ZN(n14447) );
  NAND3_X1 U16315 ( .A1(n14514), .A2(n12946), .A3(n14447), .ZN(n14444) );
  NAND2_X1 U16316 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14440) );
  INV_X1 U16317 ( .A(n14440), .ZN(n14439) );
  NOR2_X1 U16318 ( .A1(n14435), .A2(n15607), .ZN(n16726) );
  AND2_X1 U16319 ( .A1(n14436), .A2(n16726), .ZN(n14510) );
  NAND2_X1 U16320 ( .A1(n14437), .A2(n12809), .ZN(n14438) );
  AOI22_X1 U16321 ( .A1(n14584), .A2(n14439), .B1(n14510), .B2(n14438), .ZN(
        n14442) );
  NAND2_X1 U16322 ( .A1(n14584), .A2(n14440), .ZN(n14441) );
  MUX2_X1 U16323 ( .A(n14442), .B(n14441), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n14443) );
  NAND2_X1 U16324 ( .A1(n14446), .A2(n11542), .ZN(n17988) );
  AOI22_X1 U16325 ( .A1(n17988), .A2(n17940), .B1(n22296), .B2(n14447), .ZN(
        n14460) );
  OAI21_X1 U16326 ( .B1(n14584), .B2(n14280), .A(n14448), .ZN(n14450) );
  AOI21_X1 U16327 ( .B1(n14450), .B2(n14449), .A(n22330), .ZN(n14451) );
  INV_X1 U16328 ( .A(n16719), .ZN(n16725) );
  NAND2_X1 U16329 ( .A1(n14451), .A2(n16725), .ZN(n14456) );
  NOR2_X1 U16330 ( .A1(n15070), .A2(n12886), .ZN(n14452) );
  OR2_X1 U16331 ( .A1(n14453), .A2(n14452), .ZN(n14454) );
  AOI21_X1 U16332 ( .B1(n16719), .B2(n16709), .A(n14454), .ZN(n14455) );
  NAND2_X1 U16333 ( .A1(n14456), .A2(n14455), .ZN(n14458) );
  INV_X1 U16334 ( .A(n17994), .ZN(n14750) );
  NOR2_X1 U16335 ( .A1(n14752), .A2(n22424), .ZN(n22290) );
  NAND2_X1 U16336 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n22290), .ZN(n22292) );
  INV_X1 U16337 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n22278) );
  OAI22_X1 U16338 ( .A1(n14750), .A2(n22302), .B1(n22292), .B2(n22278), .ZN(
        n17938) );
  AOI21_X1 U16339 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22287), .A(n17938), 
        .ZN(n14519) );
  NAND2_X1 U16340 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14519), .ZN(
        n14459) );
  OAI21_X1 U16341 ( .B1(n14460), .B2(n14519), .A(n14459), .ZN(P1_U3469) );
  NOR3_X1 U16342 ( .A1(n14462), .A2(n12817), .A3(n14508), .ZN(n14463) );
  AOI21_X1 U16343 ( .B1(n14584), .B2(n12810), .A(n14463), .ZN(n14464) );
  OAI21_X1 U16344 ( .B1(n11193), .B2(n14514), .A(n14464), .ZN(n17995) );
  NOR2_X1 U16345 ( .A1(n14752), .A2(n21986), .ZN(n14518) );
  INV_X1 U16346 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n22087) );
  INV_X1 U16347 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17100) );
  OAI22_X1 U16348 ( .A1(n22087), .A2(n17100), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14515) );
  AND2_X1 U16349 ( .A1(n14518), .A2(n14515), .ZN(n14466) );
  INV_X1 U16350 ( .A(n22296), .ZN(n14484) );
  NOR3_X1 U16351 ( .A1(n12817), .A2(n14508), .A3(n14484), .ZN(n14465) );
  AOI211_X1 U16352 ( .C1(n17995), .C2(n17940), .A(n14466), .B(n14465), .ZN(
        n14468) );
  NAND2_X1 U16353 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n14519), .ZN(
        n14467) );
  OAI21_X1 U16354 ( .B1(n14468), .B2(n14519), .A(n14467), .ZN(P1_U3473) );
  OAI21_X1 U16355 ( .B1(n14471), .B2(n14470), .A(n14469), .ZN(n18125) );
  INV_X1 U16356 ( .A(n18125), .ZN(n19103) );
  INV_X1 U16357 ( .A(n14556), .ZN(n14574) );
  OAI211_X1 U16358 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n19378), .B(n14574), .ZN(n14474) );
  NAND2_X1 U16359 ( .A1(n19420), .A2(n14472), .ZN(n14473) );
  OAI211_X1 U16360 ( .C1(n19103), .C2(n17928), .A(n14474), .B(n14473), .ZN(
        n14479) );
  INV_X1 U16361 ( .A(n14555), .ZN(n19367) );
  AOI22_X1 U16362 ( .A1(n19419), .A2(n14475), .B1(n19367), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14477) );
  OAI211_X1 U16363 ( .C1(n14664), .C2(n19416), .A(n14477), .B(n14476), .ZN(
        n14478) );
  OR2_X1 U16364 ( .A1(n14479), .A2(n14478), .ZN(P2_U3045) );
  NAND2_X1 U16365 ( .A1(n22417), .A2(n14480), .ZN(n14483) );
  NAND2_X1 U16366 ( .A1(n14481), .A2(n11361), .ZN(n14482) );
  NAND2_X1 U16367 ( .A1(n14483), .A2(n14482), .ZN(n17992) );
  OAI22_X1 U16368 ( .A1(n14752), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14484), .ZN(n14485) );
  AOI21_X1 U16369 ( .B1(n17992), .B2(n17940), .A(n14485), .ZN(n14488) );
  NAND2_X1 U16370 ( .A1(n14584), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n17990) );
  INV_X1 U16371 ( .A(n17990), .ZN(n14486) );
  AOI22_X1 U16372 ( .A1(n14486), .A2(n17940), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14519), .ZN(n14487) );
  OAI21_X1 U16373 ( .B1(n14488), .B2(n14519), .A(n14487), .ZN(P1_U3474) );
  NAND2_X1 U16374 ( .A1(n14490), .A2(n14489), .ZN(n14493) );
  NAND3_X1 U16375 ( .A1(n21524), .A2(n19645), .A3(n14491), .ZN(n14492) );
  AOI21_X1 U16376 ( .B1(n14493), .B2(n14492), .A(n21961), .ZN(n21335) );
  NAND3_X1 U16377 ( .A1(n21335), .A2(n20904), .A3(n19027), .ZN(n18564) );
  NOR2_X2 U16378 ( .A1(n18564), .A2(n21524), .ZN(n18565) );
  NAND4_X1 U16379 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(P3_EBX_REG_9__SCAN_IN), .A4(P3_EBX_REG_8__SCAN_IN), .ZN(n18320) );
  INV_X1 U16380 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n20926) );
  NAND2_X1 U16381 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n18216) );
  NOR2_X1 U16382 ( .A1(n20926), .A2(n18216), .ZN(n18211) );
  NAND3_X1 U16383 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n18211), .ZN(n18321) );
  NOR2_X1 U16384 ( .A1(n18564), .A2(n18321), .ZN(n18237) );
  NAND4_X1 U16385 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .A4(n18237), .ZN(n18316) );
  NOR2_X1 U16386 ( .A1(n18320), .A2(n18316), .ZN(n18290) );
  INV_X1 U16387 ( .A(n18290), .ZN(n18291) );
  INV_X2 U16388 ( .A(n18565), .ZN(n18562) );
  AOI22_X1 U16389 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18480), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14503) );
  AOI22_X1 U16390 ( .A1(n18546), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14502) );
  AOI22_X1 U16391 ( .A1(n18540), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14494) );
  OAI21_X1 U16392 ( .B1(n11206), .B2(n18213), .A(n14494), .ZN(n14500) );
  AOI22_X1 U16393 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18432), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14498) );
  AOI22_X1 U16394 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14497) );
  AOI22_X1 U16395 ( .A1(n18547), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14496) );
  AOI22_X1 U16396 ( .A1(n18279), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14495) );
  NAND4_X1 U16397 ( .A1(n14498), .A2(n14497), .A3(n14496), .A4(n14495), .ZN(
        n14499) );
  AOI211_X1 U16398 ( .C1(n11156), .C2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n14500), .B(n14499), .ZN(n14501) );
  NAND3_X1 U16399 ( .A1(n14503), .A2(n14502), .A3(n14501), .ZN(n21356) );
  OAI222_X1 U16400 ( .A1(n18565), .A2(P3_EBX_REG_11__SCAN_IN), .B1(n18565), 
        .B2(n18291), .C1(n18562), .C2(n21356), .ZN(n14507) );
  INV_X1 U16401 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n14505) );
  INV_X1 U16402 ( .A(n18316), .ZN(n18229) );
  AND3_X1 U16403 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(n18229), .ZN(n18293) );
  NAND2_X1 U16404 ( .A1(n21524), .A2(n18293), .ZN(n18305) );
  INV_X1 U16405 ( .A(n18305), .ZN(n14504) );
  NAND3_X1 U16406 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n14505), .A3(n14504), 
        .ZN(n14506) );
  NAND2_X1 U16407 ( .A1(n14507), .A2(n14506), .ZN(P3_U2692) );
  XNOR2_X1 U16408 ( .A(n12810), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14511) );
  XNOR2_X1 U16409 ( .A(n14508), .B(n12809), .ZN(n14516) );
  INV_X1 U16410 ( .A(n14516), .ZN(n14509) );
  AOI22_X1 U16411 ( .A1(n14584), .A2(n14511), .B1(n14510), .B2(n14509), .ZN(
        n14513) );
  NAND3_X1 U16412 ( .A1(n14514), .A2(n12946), .A3(n14516), .ZN(n14512) );
  OAI211_X1 U16413 ( .C1(n22418), .C2(n14514), .A(n14513), .B(n14512), .ZN(
        n17989) );
  INV_X1 U16414 ( .A(n14515), .ZN(n14517) );
  AOI222_X1 U16415 ( .A1(n17989), .A2(n17940), .B1(n14518), .B2(n14517), .C1(
        n14516), .C2(n22296), .ZN(n14520) );
  INV_X1 U16416 ( .A(n14519), .ZN(n17943) );
  MUX2_X1 U16417 ( .A(n12809), .B(n14520), .S(n17943), .Z(n14521) );
  INV_X1 U16418 ( .A(n14521), .ZN(P1_U3472) );
  INV_X1 U16419 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n14527) );
  INV_X1 U16420 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n14523) );
  OR2_X1 U16421 ( .A1(n16030), .A2(n14523), .ZN(n14525) );
  NAND2_X1 U16422 ( .A1(n16030), .A2(BUF2_REG_2__SCAN_IN), .ZN(n14524) );
  AND2_X1 U16423 ( .A1(n14525), .A2(n14524), .ZN(n20328) );
  NOR2_X1 U16424 ( .A1(n14536), .A2(n20328), .ZN(n14539) );
  AOI21_X1 U16425 ( .B1(n14549), .B2(P2_EAX_REG_18__SCAN_IN), .A(n14539), .ZN(
        n14526) );
  OAI21_X1 U16426 ( .B1(n14394), .B2(n14527), .A(n14526), .ZN(P2_U2954) );
  INV_X1 U16427 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n14532) );
  INV_X1 U16428 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n14528) );
  OR2_X1 U16429 ( .A1(n16030), .A2(n14528), .ZN(n14530) );
  NAND2_X1 U16430 ( .A1(n16030), .A2(BUF2_REG_3__SCAN_IN), .ZN(n14529) );
  AND2_X1 U16431 ( .A1(n14530), .A2(n14529), .ZN(n16241) );
  NOR2_X1 U16432 ( .A1(n14536), .A2(n16241), .ZN(n14542) );
  AOI21_X1 U16433 ( .B1(n14549), .B2(P2_EAX_REG_19__SCAN_IN), .A(n14542), .ZN(
        n14531) );
  OAI21_X1 U16434 ( .B1(n14394), .B2(n14532), .A(n14531), .ZN(P2_U2955) );
  INV_X1 U16435 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n14538) );
  INV_X1 U16436 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n14533) );
  OR2_X1 U16437 ( .A1(n16030), .A2(n14533), .ZN(n14535) );
  NAND2_X1 U16438 ( .A1(n16030), .A2(BUF2_REG_1__SCAN_IN), .ZN(n14534) );
  AND2_X1 U16439 ( .A1(n14535), .A2(n14534), .ZN(n16035) );
  NOR2_X1 U16440 ( .A1(n14536), .A2(n16035), .ZN(n14548) );
  AOI21_X1 U16441 ( .B1(n14549), .B2(P2_EAX_REG_17__SCAN_IN), .A(n14548), .ZN(
        n14537) );
  OAI21_X1 U16442 ( .B1(n14394), .B2(n14538), .A(n14537), .ZN(P2_U2953) );
  INV_X1 U16443 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n14541) );
  AOI21_X1 U16444 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(n14549), .A(n14539), .ZN(
        n14540) );
  OAI21_X1 U16445 ( .B1(n14394), .B2(n14541), .A(n14540), .ZN(P2_U2969) );
  INV_X1 U16446 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n14544) );
  AOI21_X1 U16447 ( .B1(n14549), .B2(P2_EAX_REG_3__SCAN_IN), .A(n14542), .ZN(
        n14543) );
  OAI21_X1 U16448 ( .B1(n14394), .B2(n14544), .A(n14543), .ZN(P2_U2970) );
  INV_X1 U16449 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n14547) );
  AOI21_X1 U16450 ( .B1(n14549), .B2(P2_EAX_REG_4__SCAN_IN), .A(n14545), .ZN(
        n14546) );
  OAI21_X1 U16451 ( .B1(n14394), .B2(n14547), .A(n14546), .ZN(P2_U2971) );
  INV_X1 U16452 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n14551) );
  AOI21_X1 U16453 ( .B1(P2_EAX_REG_1__SCAN_IN), .B2(n14549), .A(n14548), .ZN(
        n14550) );
  OAI21_X1 U16454 ( .B1(n14394), .B2(n14551), .A(n14550), .ZN(P2_U2968) );
  INV_X1 U16455 ( .A(P2_LWORD_REG_14__SCAN_IN), .ZN(n14554) );
  NAND2_X1 U16456 ( .A1(n14549), .A2(P2_EAX_REG_14__SCAN_IN), .ZN(n14552) );
  OAI211_X1 U16457 ( .C1(n14394), .C2(n14554), .A(n14553), .B(n14552), .ZN(
        P2_U2981) );
  OAI21_X1 U16458 ( .B1(n17787), .B2(n14556), .A(n14555), .ZN(n15477) );
  INV_X1 U16459 ( .A(n17787), .ZN(n17902) );
  NAND2_X1 U16460 ( .A1(n17902), .A2(n14557), .ZN(n15476) );
  INV_X1 U16461 ( .A(n14558), .ZN(n14559) );
  NAND2_X1 U16462 ( .A1(n14560), .A2(n14559), .ZN(n14561) );
  AND2_X1 U16463 ( .A1(n14562), .A2(n14561), .ZN(n18030) );
  AOI21_X1 U16464 ( .B1(n14565), .B2(n14564), .A(n14563), .ZN(n18029) );
  AOI22_X1 U16465 ( .A1(n19419), .A2(n18030), .B1(n19420), .B2(n18029), .ZN(
        n14573) );
  XNOR2_X1 U16466 ( .A(n14567), .B(n14566), .ZN(n18120) );
  INV_X1 U16467 ( .A(n15474), .ZN(n19410) );
  AOI21_X1 U16468 ( .B1(n19410), .B2(n14568), .A(n17923), .ZN(n14571) );
  NOR2_X1 U16469 ( .A1(n19380), .A2(n14569), .ZN(n14570) );
  AOI211_X1 U16470 ( .C1(n19408), .C2(n18120), .A(n14571), .B(n14570), .ZN(
        n14572) );
  OAI211_X1 U16471 ( .C1(n14574), .C2(n15476), .A(n14573), .B(n14572), .ZN(
        n14575) );
  AOI21_X1 U16472 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n15477), .A(
        n14575), .ZN(n14576) );
  OAI21_X1 U16473 ( .B1(n15133), .B2(n19416), .A(n14576), .ZN(P2_U3044) );
  INV_X1 U16474 ( .A(n16020), .ZN(n14577) );
  NAND2_X1 U16475 ( .A1(n14577), .A2(n15163), .ZN(n15109) );
  INV_X1 U16476 ( .A(n15127), .ZN(n14578) );
  NAND2_X1 U16477 ( .A1(n15109), .A2(n14578), .ZN(n14579) );
  MUX2_X1 U16478 ( .A(n16344), .B(n14582), .S(n17423), .Z(n14583) );
  OAI21_X1 U16479 ( .B1(n19929), .B2(n17428), .A(n14583), .ZN(P2_U2887) );
  INV_X1 U16480 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14589) );
  NAND2_X1 U16481 ( .A1(n14584), .A2(n22807), .ZN(n14585) );
  OR2_X1 U16482 ( .A1(n14585), .A2(n16719), .ZN(n14586) );
  NAND2_X1 U16483 ( .A1(n20604), .A2(n16710), .ZN(n14974) );
  AND2_X2 U16484 ( .A1(n22287), .A2(n22290), .ZN(n20633) );
  AOI22_X1 U16485 ( .A1(n20633), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20620), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14588) );
  OAI21_X1 U16486 ( .B1(n14589), .B2(n14974), .A(n14588), .ZN(P1_U2918) );
  INV_X1 U16487 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14591) );
  AOI22_X1 U16488 ( .A1(n20633), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20620), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14590) );
  OAI21_X1 U16489 ( .B1(n14591), .B2(n14974), .A(n14590), .ZN(P1_U2919) );
  NAND2_X1 U16490 ( .A1(n14592), .A2(n14704), .ZN(n14595) );
  AND2_X1 U16491 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20061) );
  NAND2_X1 U16492 ( .A1(n20061), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14706) );
  INV_X1 U16493 ( .A(n20061), .ZN(n15121) );
  NAND2_X1 U16494 ( .A1(n15121), .A2(n19998), .ZN(n14593) );
  AND2_X1 U16495 ( .A1(n14706), .A2(n14593), .ZN(n19951) );
  AOI22_X1 U16496 ( .A1(n14709), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n20100), .B2(n19951), .ZN(n14594) );
  NAND2_X1 U16497 ( .A1(n14595), .A2(n14594), .ZN(n14598) );
  OR2_X1 U16498 ( .A1(n14598), .A2(n14597), .ZN(n14599) );
  NAND2_X1 U16499 ( .A1(n14598), .A2(n14597), .ZN(n14717) );
  INV_X1 U16500 ( .A(n16597), .ZN(n14600) );
  INV_X1 U16501 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n16516) );
  NAND2_X1 U16502 ( .A1(n14709), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14602) );
  NOR2_X1 U16503 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20045) );
  INV_X1 U16504 ( .A(n20045), .ZN(n14601) );
  NAND2_X1 U16505 ( .A1(n15121), .A2(n14601), .ZN(n20017) );
  OR2_X1 U16506 ( .A1(n20017), .A2(n20096), .ZN(n20079) );
  NAND2_X1 U16507 ( .A1(n14602), .A2(n20079), .ZN(n14603) );
  INV_X1 U16508 ( .A(n14604), .ZN(n14605) );
  NOR2_X1 U16509 ( .A1(n14606), .A2(n14605), .ZN(n14607) );
  INV_X1 U16510 ( .A(n14715), .ZN(n14608) );
  MUX2_X1 U16511 ( .A(n15133), .B(n14609), .S(n17423), .Z(n14610) );
  OAI21_X1 U16512 ( .B1(n16017), .B2(n17428), .A(n14610), .ZN(P2_U2885) );
  XNOR2_X1 U16513 ( .A(n19944), .B(n18125), .ZN(n14614) );
  NOR2_X1 U16514 ( .A1(n19929), .A2(n19366), .ZN(n14613) );
  NOR2_X1 U16515 ( .A1(n14614), .A2(n14613), .ZN(n14976) );
  AOI21_X1 U16516 ( .B1(n14614), .B2(n14613), .A(n14976), .ZN(n14617) );
  AOI22_X1 U16517 ( .A1(n20321), .A2(n18125), .B1(n20319), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n14616) );
  INV_X1 U16518 ( .A(n16035), .ZN(n16135) );
  NAND2_X1 U16519 ( .A1(n20164), .A2(n16135), .ZN(n14615) );
  OAI211_X1 U16520 ( .C1(n14617), .C2(n20165), .A(n14616), .B(n14615), .ZN(
        P2_U2918) );
  XNOR2_X1 U16521 ( .A(n14620), .B(n14619), .ZN(n19134) );
  INV_X1 U16522 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n18161) );
  OAI222_X1 U16523 ( .A1(n15324), .A2(n20114), .B1(n19134), .B2(n20171), .C1(
        n17475), .C2(n18161), .ZN(P2_U2913) );
  OAI21_X1 U16524 ( .B1(n14623), .B2(n14622), .A(n14621), .ZN(n19145) );
  OAI222_X1 U16525 ( .A1(n15324), .A2(n19919), .B1(n19145), .B2(n20171), .C1(
        n17475), .C2(n18163), .ZN(P2_U2912) );
  NAND2_X1 U16526 ( .A1(n14625), .A2(n14624), .ZN(n14627) );
  NAND2_X1 U16527 ( .A1(n14627), .A2(n14626), .ZN(n14675) );
  OAI21_X1 U16528 ( .B1(n14627), .B2(n14626), .A(n14675), .ZN(n15090) );
  NAND3_X1 U16529 ( .A1(n22287), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n22289) );
  NOR2_X1 U16530 ( .A1(n16719), .A2(n14628), .ZN(n18014) );
  NAND2_X1 U16531 ( .A1(n14629), .A2(n22468), .ZN(n21969) );
  NAND2_X1 U16532 ( .A1(n21969), .A2(n22287), .ZN(n14630) );
  NAND2_X1 U16533 ( .A1(n22287), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14632) );
  NAND2_X1 U16534 ( .A1(n22305), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14631) );
  AND2_X1 U16535 ( .A1(n14632), .A2(n14631), .ZN(n20729) );
  INV_X1 U16536 ( .A(n20729), .ZN(n14633) );
  INV_X1 U16537 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15088) );
  NAND2_X1 U16538 ( .A1(n22021), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n22080) );
  OAI21_X1 U16539 ( .B1(n20728), .B2(n15088), .A(n22080), .ZN(n14634) );
  AOI21_X1 U16540 ( .B1(n20761), .B2(n15088), .A(n14634), .ZN(n14642) );
  NAND2_X1 U16541 ( .A1(n13019), .A2(n12947), .ZN(n14639) );
  NAND2_X1 U16542 ( .A1(n14636), .A2(n14635), .ZN(n14934) );
  OAI211_X1 U16543 ( .C1(n14636), .C2(n14635), .A(n15607), .B(n14934), .ZN(
        n14637) );
  AND3_X1 U16544 ( .A1(n14637), .A2(n12940), .A3(n11160), .ZN(n14638) );
  XNOR2_X1 U16545 ( .A(n14692), .B(n14690), .ZN(n14640) );
  OR2_X1 U16546 ( .A1(n14640), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n22077) );
  NAND2_X1 U16547 ( .A1(n14640), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n22076) );
  INV_X1 U16548 ( .A(n22277), .ZN(n20756) );
  NAND3_X1 U16549 ( .A1(n22077), .A2(n22076), .A3(n20756), .ZN(n14641) );
  OAI211_X1 U16550 ( .C1(n15090), .C2(n17060), .A(n14642), .B(n14641), .ZN(
        P1_U2998) );
  INV_X1 U16551 ( .A(n17459), .ZN(n14646) );
  AOI21_X1 U16552 ( .B1(n14644), .B2(n14621), .A(n14643), .ZN(n19395) );
  INV_X1 U16553 ( .A(n19395), .ZN(n14645) );
  INV_X1 U16554 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n18165) );
  OAI222_X1 U16555 ( .A1(n15324), .A2(n14646), .B1(n14645), .B2(n20171), .C1(
        n17475), .C2(n18165), .ZN(P2_U2911) );
  INV_X1 U16556 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20608) );
  OAI222_X1 U16557 ( .A1(n15090), .A2(n16897), .B1(n16056), .B2(n14914), .C1(
        n16054), .C2(n20608), .ZN(P1_U2903) );
  INV_X1 U16558 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n15080) );
  NAND2_X1 U16559 ( .A1(n14857), .A2(n22087), .ZN(n14647) );
  OAI211_X1 U16560 ( .C1(P1_EBX_REG_1__SCAN_IN), .C2(n11150), .A(n14647), .B(
        n16385), .ZN(n14648) );
  XNOR2_X1 U16561 ( .A(n14679), .B(n14649), .ZN(n14650) );
  NAND2_X1 U16562 ( .A1(n14650), .A2(n11192), .ZN(n14680) );
  OAI21_X1 U16563 ( .B1(n14650), .B2(n11192), .A(n14680), .ZN(n15082) );
  INV_X1 U16564 ( .A(n15082), .ZN(n22083) );
  OAI222_X1 U16565 ( .A1(n20698), .A2(n15090), .B1(n15080), .B2(n20727), .C1(
        n16841), .C2(n22083), .ZN(P1_U2871) );
  AOI22_X1 U16566 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n18179), .B1(n18180), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n14651) );
  OAI21_X1 U16567 ( .B1(n16174), .B2(n14662), .A(n14651), .ZN(P2_U2935) );
  AOI22_X1 U16568 ( .A1(n18180), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n14652) );
  OAI21_X1 U16569 ( .B1(n16652), .B2(n14662), .A(n14652), .ZN(P2_U2922) );
  INV_X1 U16570 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n17449) );
  AOI22_X1 U16571 ( .A1(n18180), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n14653) );
  OAI21_X1 U16572 ( .B1(n17449), .B2(n14662), .A(n14653), .ZN(P2_U2926) );
  AOI22_X1 U16573 ( .A1(n18180), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n14654) );
  OAI21_X1 U16574 ( .B1(n14397), .B2(n14662), .A(n14654), .ZN(P2_U2925) );
  AOI22_X1 U16575 ( .A1(n18180), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n14655) );
  OAI21_X1 U16576 ( .B1(n17435), .B2(n14662), .A(n14655), .ZN(P2_U2924) );
  AOI22_X1 U16577 ( .A1(n18180), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n14656) );
  OAI21_X1 U16578 ( .B1(n17429), .B2(n14662), .A(n14656), .ZN(P2_U2923) );
  INV_X1 U16579 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n14658) );
  AOI22_X1 U16580 ( .A1(n18180), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n14657) );
  OAI21_X1 U16581 ( .B1(n14658), .B2(n14662), .A(n14657), .ZN(P2_U2931) );
  AOI22_X1 U16582 ( .A1(n18168), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n14659) );
  OAI21_X1 U16583 ( .B1(n16689), .B2(n14662), .A(n14659), .ZN(P2_U2921) );
  INV_X1 U16584 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n16133) );
  AOI22_X1 U16585 ( .A1(n18168), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n14660) );
  OAI21_X1 U16586 ( .B1(n16133), .B2(n14662), .A(n14660), .ZN(P2_U2934) );
  INV_X1 U16587 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n14663) );
  AOI22_X1 U16588 ( .A1(n18168), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n14661) );
  OAI21_X1 U16589 ( .B1(n14663), .B2(n14662), .A(n14661), .ZN(P2_U2933) );
  INV_X1 U16590 ( .A(n19944), .ZN(n18128) );
  NOR2_X1 U16591 ( .A1(n14664), .A2(n17420), .ZN(n14665) );
  AOI21_X1 U16592 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n17420), .A(n14665), .ZN(
        n14666) );
  OAI21_X1 U16593 ( .B1(n18128), .B2(n17428), .A(n14666), .ZN(P2_U2886) );
  OR2_X1 U16594 ( .A1(n14667), .A2(n14643), .ZN(n14669) );
  NAND2_X1 U16595 ( .A1(n14669), .A2(n14668), .ZN(n19161) );
  INV_X1 U16596 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n18167) );
  OAI222_X1 U16597 ( .A1(n19161), .A2(n20171), .B1(n15324), .B2(n14670), .C1(
        n17475), .C2(n18167), .ZN(P2_U2910) );
  OR2_X1 U16598 ( .A1(n14672), .A2(n14671), .ZN(n14673) );
  AND2_X1 U16599 ( .A1(n14674), .A2(n14673), .ZN(n14676) );
  OR2_X1 U16600 ( .A1(n14676), .A2(n14675), .ZN(n14678) );
  NAND2_X1 U16601 ( .A1(n14676), .A2(n14675), .ZN(n14677) );
  AND2_X1 U16602 ( .A1(n14678), .A2(n14677), .ZN(n15098) );
  INV_X1 U16603 ( .A(n15098), .ZN(n14730) );
  NAND2_X1 U16604 ( .A1(n14680), .A2(n14679), .ZN(n14686) );
  INV_X1 U16605 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n15971) );
  NAND2_X1 U16606 ( .A1(n16293), .A2(n15971), .ZN(n14683) );
  INV_X1 U16607 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n22003) );
  NAND2_X1 U16608 ( .A1(n14857), .A2(n22003), .ZN(n14681) );
  OAI211_X1 U16609 ( .C1(P1_EBX_REG_2__SCAN_IN), .C2(n11150), .A(n14681), .B(
        n16385), .ZN(n14682) );
  NAND2_X1 U16610 ( .A1(n14686), .A2(n14685), .ZN(n14687) );
  AND2_X1 U16611 ( .A1(n14856), .A2(n14687), .ZN(n21995) );
  INV_X1 U16612 ( .A(n20727), .ZN(n16821) );
  AOI22_X1 U16613 ( .A1(n20724), .A2(n21995), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n16821), .ZN(n14688) );
  OAI21_X1 U16614 ( .B1(n14730), .B2(n20698), .A(n14688), .ZN(P1_U2870) );
  INV_X1 U16615 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n22099) );
  NOR2_X1 U16616 ( .A1(n22066), .A2(n22099), .ZN(n21994) );
  NOR2_X1 U16617 ( .A1(n20759), .A2(n15101), .ZN(n14689) );
  AOI211_X1 U16618 ( .C1(n20760), .C2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n21994), .B(n14689), .ZN(n14703) );
  INV_X1 U16619 ( .A(n14690), .ZN(n14691) );
  NAND2_X1 U16620 ( .A1(n14692), .A2(n14691), .ZN(n14693) );
  NAND2_X1 U16621 ( .A1(n22076), .A2(n14693), .ZN(n14940) );
  XNOR2_X1 U16622 ( .A(n14940), .B(n22003), .ZN(n14701) );
  NAND2_X1 U16623 ( .A1(n11195), .A2(n15602), .ZN(n14699) );
  INV_X1 U16624 ( .A(n14694), .ZN(n14933) );
  XNOR2_X1 U16625 ( .A(n14934), .B(n14933), .ZN(n14697) );
  INV_X1 U16626 ( .A(n14695), .ZN(n14696) );
  AOI21_X1 U16627 ( .B1(n14697), .B2(n15607), .A(n14696), .ZN(n14698) );
  NAND2_X1 U16628 ( .A1(n14699), .A2(n14698), .ZN(n14700) );
  OR2_X1 U16629 ( .A1(n14701), .A2(n14700), .ZN(n21991) );
  NAND2_X1 U16630 ( .A1(n14701), .A2(n14700), .ZN(n21990) );
  NAND3_X1 U16631 ( .A1(n21991), .A2(n21990), .A3(n20756), .ZN(n14702) );
  OAI211_X1 U16632 ( .C1(n14730), .C2(n17060), .A(n14703), .B(n14702), .ZN(
        P1_U2997) );
  NAND2_X1 U16633 ( .A1(n14705), .A2(n14704), .ZN(n14711) );
  AOI21_X1 U16634 ( .B1(n14706), .B2(n19952), .A(n20096), .ZN(n14708) );
  INV_X1 U16635 ( .A(n14706), .ZN(n14707) );
  NAND2_X1 U16636 ( .A1(n14707), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16019) );
  AOI22_X1 U16637 ( .A1(n14709), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n14708), .B2(n16019), .ZN(n14710) );
  NAND2_X1 U16638 ( .A1(n14711), .A2(n14710), .ZN(n14713) );
  OR2_X1 U16639 ( .A1(n14713), .A2(n14712), .ZN(n14714) );
  NAND2_X1 U16640 ( .A1(n14713), .A2(n14712), .ZN(n14720) );
  NAND2_X1 U16641 ( .A1(n14716), .A2(n14715), .ZN(n14718) );
  NAND2_X1 U16642 ( .A1(n14731), .A2(n14732), .ZN(n14733) );
  NAND2_X1 U16643 ( .A1(n11649), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14719) );
  NAND2_X1 U16644 ( .A1(n14739), .A2(n14740), .ZN(n14766) );
  XOR2_X1 U16645 ( .A(n14766), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n14729)
         );
  NAND2_X1 U16646 ( .A1(n14723), .A2(n14722), .ZN(n14726) );
  INV_X1 U16647 ( .A(n14724), .ZN(n14725) );
  NAND2_X1 U16648 ( .A1(n14726), .A2(n14725), .ZN(n19122) );
  NOR2_X1 U16649 ( .A1(n17423), .A2(n19122), .ZN(n14727) );
  AOI21_X1 U16650 ( .B1(P2_EBX_REG_5__SCAN_IN), .B2(n17420), .A(n14727), .ZN(
        n14728) );
  OAI21_X1 U16651 ( .B1(n14729), .B2(n17428), .A(n14728), .ZN(P2_U2882) );
  INV_X1 U16652 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20610) );
  OAI222_X1 U16653 ( .A1(n14730), .A2(n16897), .B1(n16056), .B2(n14894), .C1(
        n16054), .C2(n20610), .ZN(P1_U2902) );
  NOR2_X1 U16654 ( .A1(n12312), .A2(n17420), .ZN(n14735) );
  AOI21_X1 U16655 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n17420), .A(n14735), .ZN(
        n14736) );
  OAI21_X1 U16656 ( .B1(n20058), .B2(n17428), .A(n14736), .ZN(P2_U2884) );
  INV_X1 U16657 ( .A(n17444), .ZN(n14738) );
  XNOR2_X1 U16658 ( .A(n14668), .B(n14737), .ZN(n19172) );
  INV_X1 U16659 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n18170) );
  OAI222_X1 U16660 ( .A1(n15324), .A2(n14738), .B1(n19172), .B2(n20171), .C1(
        n17475), .C2(n18170), .ZN(P2_U2909) );
  OAI21_X1 U16661 ( .B1(n14739), .B2(n14740), .A(n14766), .ZN(n20166) );
  OR2_X1 U16662 ( .A1(n14742), .A2(n14741), .ZN(n14743) );
  NAND2_X1 U16663 ( .A1(n14743), .A2(n14722), .ZN(n18045) );
  NOR2_X1 U16664 ( .A1(n18045), .A2(n17420), .ZN(n14744) );
  AOI21_X1 U16665 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n17423), .A(n14744), .ZN(
        n14745) );
  OAI21_X1 U16666 ( .B1(n20166), .B2(n17428), .A(n14745), .ZN(P2_U2883) );
  NAND2_X1 U16667 ( .A1(n14746), .A2(n22278), .ZN(n14747) );
  NOR2_X1 U16668 ( .A1(n14747), .A2(n12817), .ZN(n14755) );
  INV_X1 U16669 ( .A(n14823), .ZN(n14780) );
  OR2_X1 U16670 ( .A1(n14748), .A2(n14780), .ZN(n14749) );
  XNOR2_X1 U16671 ( .A(n14749), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n22107) );
  INV_X1 U16672 ( .A(n13678), .ZN(n17939) );
  AOI21_X1 U16673 ( .B1(n22107), .B2(n17939), .A(n14750), .ZN(n14751) );
  MUX2_X1 U16674 ( .A(P1_FLUSH_REG_SCAN_IN), .B(n14751), .S(n14752), .Z(n14754) );
  AOI21_X1 U16675 ( .B1(n14752), .B2(n17994), .A(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14753) );
  NOR2_X1 U16676 ( .A1(n14754), .A2(n14753), .ZN(n18005) );
  OR2_X1 U16677 ( .A1(n14755), .A2(n18005), .ZN(n22283) );
  INV_X1 U16678 ( .A(n22292), .ZN(n14756) );
  OAI21_X1 U16679 ( .B1(n22283), .B2(P1_FLUSH_REG_SCAN_IN), .A(n14756), .ZN(
        n14758) );
  NAND2_X1 U16680 ( .A1(n14758), .A2(n22678), .ZN(n18023) );
  INV_X1 U16681 ( .A(n18023), .ZN(n22286) );
  NAND2_X1 U16682 ( .A1(n11196), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22422) );
  OAI21_X1 U16683 ( .B1(n14841), .B2(n22422), .A(n15033), .ZN(n14762) );
  OAI21_X1 U16684 ( .B1(n22422), .B2(n14874), .A(n14762), .ZN(n14763) );
  INV_X1 U16685 ( .A(n22468), .ZN(n22434) );
  NAND2_X1 U16686 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n14188), .ZN(n22281) );
  AOI22_X1 U16687 ( .A1(n14763), .A2(n22434), .B1(n22281), .B2(n14427), .ZN(
        n14765) );
  NAND2_X1 U16688 ( .A1(n22286), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14764) );
  OAI21_X1 U16689 ( .B1(n22286), .B2(n14765), .A(n14764), .ZN(P1_U3475) );
  INV_X1 U16690 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16601) );
  NOR2_X1 U16691 ( .A1(n14766), .A2(n16601), .ZN(n14767) );
  OAI211_X1 U16692 ( .C1(n14767), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n17417), .B(n14989), .ZN(n14772) );
  OR2_X1 U16693 ( .A1(n14768), .A2(n14724), .ZN(n14770) );
  NAND2_X1 U16694 ( .A1(n14770), .A2(n14769), .ZN(n19133) );
  INV_X1 U16695 ( .A(n19133), .ZN(n17921) );
  NAND2_X1 U16696 ( .A1(n14580), .A2(n17921), .ZN(n14771) );
  OAI211_X1 U16697 ( .C1(n14580), .C2(n12197), .A(n14772), .B(n14771), .ZN(
        P2_U2881) );
  INV_X1 U16698 ( .A(n22422), .ZN(n14773) );
  NAND2_X1 U16699 ( .A1(n14773), .A2(n22434), .ZN(n17330) );
  OR2_X1 U16700 ( .A1(n15215), .A2(n22441), .ZN(n14783) );
  OAI21_X1 U16701 ( .B1(n17330), .B2(n14841), .A(n14783), .ZN(n14774) );
  INV_X1 U16702 ( .A(n15035), .ZN(n22427) );
  NAND2_X1 U16703 ( .A1(n14774), .A2(n15035), .ZN(n22798) );
  INV_X1 U16704 ( .A(n22798), .ZN(n14813) );
  INV_X1 U16705 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14792) );
  INV_X1 U16706 ( .A(n22400), .ZN(n14873) );
  INV_X1 U16707 ( .A(n22801), .ZN(n15212) );
  INV_X1 U16708 ( .A(DATAI_30_), .ZN(n14777) );
  NAND2_X1 U16709 ( .A1(n14775), .A2(n20762), .ZN(n22686) );
  INV_X1 U16710 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20827) );
  OR2_X1 U16711 ( .A1(n22686), .A2(n20827), .ZN(n14776) );
  OAI21_X1 U16712 ( .B1(n22688), .B2(n14777), .A(n14776), .ZN(n22674) );
  INV_X1 U16713 ( .A(n22688), .ZN(n14904) );
  NAND2_X1 U16714 ( .A1(n14904), .A2(DATAI_22_), .ZN(n14779) );
  INV_X1 U16715 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20809) );
  OR2_X1 U16716 ( .A1(n22686), .A2(n20809), .ZN(n14778) );
  AND2_X1 U16717 ( .A1(n14779), .A2(n14778), .ZN(n22672) );
  OR2_X1 U16718 ( .A1(n22418), .A2(n14780), .ZN(n22472) );
  NOR2_X1 U16719 ( .A1(n11154), .A2(n22468), .ZN(n14781) );
  AND2_X1 U16720 ( .A1(n14781), .A2(n22417), .ZN(n15022) );
  INV_X1 U16721 ( .A(n15022), .ZN(n14786) );
  NAND2_X1 U16722 ( .A1(n14782), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14807) );
  OAI22_X1 U16723 ( .A1(n14807), .A2(n22468), .B1(n14783), .B2(n22424), .ZN(
        n14784) );
  INV_X1 U16724 ( .A(n14784), .ZN(n14785) );
  OAI21_X1 U16725 ( .B1(n22472), .B2(n14786), .A(n14785), .ZN(n22795) );
  NOR2_X1 U16726 ( .A1(n22678), .A2(n15283), .ZN(n15248) );
  NAND2_X1 U16727 ( .A1(n12957), .A2(n22682), .ZN(n22671) );
  NOR2_X1 U16728 ( .A1(n22671), .A2(n14807), .ZN(n14788) );
  AOI21_X1 U16729 ( .B1(n22795), .B2(n15248), .A(n14788), .ZN(n14789) );
  OAI21_X1 U16730 ( .B1(n22684), .B2(n22672), .A(n14789), .ZN(n14790) );
  AOI21_X1 U16731 ( .B1(n15212), .B2(n22674), .A(n14790), .ZN(n14791) );
  OAI21_X1 U16732 ( .B1(n14813), .B2(n14792), .A(n14791), .ZN(P1_U3159) );
  INV_X1 U16733 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14801) );
  INV_X1 U16734 ( .A(DATAI_27_), .ZN(n14794) );
  INV_X1 U16735 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20820) );
  OR2_X1 U16736 ( .A1(n22686), .A2(n20820), .ZN(n14793) );
  OAI21_X1 U16737 ( .B1(n22688), .B2(n14794), .A(n14793), .ZN(n22580) );
  INV_X1 U16738 ( .A(DATAI_19_), .ZN(n14796) );
  INV_X1 U16739 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20803) );
  OR2_X1 U16740 ( .A1(n22686), .A2(n20803), .ZN(n14795) );
  OAI21_X1 U16741 ( .B1(n22688), .B2(n14796), .A(n14795), .ZN(n22571) );
  INV_X1 U16742 ( .A(n22571), .ZN(n22578) );
  NOR2_X1 U16743 ( .A1(n22678), .A2(n14869), .ZN(n15231) );
  NAND2_X1 U16744 ( .A1(n14797), .A2(n22682), .ZN(n22577) );
  INV_X1 U16745 ( .A(n22577), .ZN(n22570) );
  INV_X1 U16746 ( .A(n14807), .ZN(n22793) );
  AOI22_X1 U16747 ( .A1(n22795), .A2(n15231), .B1(n22570), .B2(n22793), .ZN(
        n14798) );
  OAI21_X1 U16748 ( .B1(n22684), .B2(n22578), .A(n14798), .ZN(n14799) );
  AOI21_X1 U16749 ( .B1(n15212), .B2(n22580), .A(n14799), .ZN(n14800) );
  OAI21_X1 U16750 ( .B1(n14813), .B2(n14801), .A(n14800), .ZN(P1_U3156) );
  INV_X1 U16751 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14812) );
  INV_X1 U16752 ( .A(DATAI_16_), .ZN(n14803) );
  INV_X1 U16753 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20797) );
  OR2_X1 U16754 ( .A1(n22686), .A2(n20797), .ZN(n14802) );
  OAI21_X1 U16755 ( .B1(n22688), .B2(n14803), .A(n14802), .ZN(n22465) );
  INV_X1 U16756 ( .A(DATAI_24_), .ZN(n14805) );
  INV_X1 U16757 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20814) );
  OR2_X1 U16758 ( .A1(n22686), .A2(n20814), .ZN(n14804) );
  OAI21_X1 U16759 ( .B1(n22688), .B2(n14805), .A(n14804), .ZN(n22487) );
  INV_X1 U16760 ( .A(n22487), .ZN(n22407) );
  NOR2_X1 U16761 ( .A1(n22678), .A2(n14806), .ZN(n15222) );
  NAND2_X1 U16762 ( .A1(n16710), .A2(n22682), .ZN(n22477) );
  NOR2_X1 U16763 ( .A1(n22477), .A2(n14807), .ZN(n14808) );
  AOI21_X1 U16764 ( .B1(n22795), .B2(n15222), .A(n14808), .ZN(n14809) );
  OAI21_X1 U16765 ( .B1(n22801), .B2(n22407), .A(n14809), .ZN(n14810) );
  AOI21_X1 U16766 ( .B1(n22797), .B2(n22465), .A(n14810), .ZN(n14811) );
  OAI21_X1 U16767 ( .B1(n14813), .B2(n14812), .A(n14811), .ZN(P1_U3153) );
  AND2_X1 U16768 ( .A1(n14816), .A2(n14815), .ZN(n14817) );
  OR2_X1 U16769 ( .A1(n14814), .A2(n14817), .ZN(n20736) );
  INV_X1 U16770 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20614) );
  OAI222_X1 U16771 ( .A1(n20736), .A2(n16897), .B1(n16056), .B2(n14881), .C1(
        n20614), .C2(n16054), .ZN(P1_U2900) );
  INV_X1 U16772 ( .A(n17437), .ZN(n14822) );
  OR2_X1 U16773 ( .A1(n14819), .A2(n14818), .ZN(n14821) );
  NAND2_X1 U16774 ( .A1(n14821), .A2(n14820), .ZN(n19176) );
  INV_X1 U16775 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n18172) );
  OAI222_X1 U16776 ( .A1(n15324), .A2(n14822), .B1(n19176), .B2(n20171), .C1(
        n17475), .C2(n18172), .ZN(P2_U2908) );
  INV_X1 U16777 ( .A(n22580), .ZN(n22564) );
  NOR3_X1 U16778 ( .A1(n18000), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14828) );
  NOR2_X1 U16779 ( .A1(n22418), .A2(n14823), .ZN(n22438) );
  INV_X1 U16780 ( .A(n14824), .ZN(n15038) );
  INV_X1 U16781 ( .A(n14828), .ZN(n15419) );
  NOR2_X1 U16782 ( .A1(n22457), .A2(n15419), .ZN(n22721) );
  AOI21_X1 U16783 ( .B1(n22438), .B2(n15038), .A(n22721), .ZN(n14827) );
  OAI211_X1 U16784 ( .C1(n14874), .C2(n22305), .A(n22434), .B(n14827), .ZN(
        n14825) );
  OAI211_X1 U16785 ( .C1(n22434), .C2(n14828), .A(n14825), .B(n15035), .ZN(
        n22723) );
  NAND2_X1 U16786 ( .A1(n22723), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n14832) );
  INV_X1 U16787 ( .A(n14827), .ZN(n14829) );
  AOI22_X1 U16788 ( .A1(n14829), .A2(n22434), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14828), .ZN(n22499) );
  INV_X1 U16789 ( .A(n22721), .ZN(n14836) );
  OAI22_X1 U16790 ( .A1(n22499), .A2(n22583), .B1(n22577), .B2(n14836), .ZN(
        n14830) );
  AOI21_X1 U16791 ( .B1(n22730), .B2(n22571), .A(n14830), .ZN(n14831) );
  OAI211_X1 U16792 ( .C1(n22564), .C2(n22726), .A(n14832), .B(n14831), .ZN(
        P1_U3076) );
  INV_X1 U16793 ( .A(n22674), .ZN(n22655) );
  NAND2_X1 U16794 ( .A1(n22723), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n14835) );
  INV_X1 U16795 ( .A(n22672), .ZN(n22665) );
  OAI22_X1 U16796 ( .A1(n22499), .A2(n22677), .B1(n22671), .B2(n14836), .ZN(
        n14833) );
  AOI21_X1 U16797 ( .B1(n22730), .B2(n22665), .A(n14833), .ZN(n14834) );
  OAI211_X1 U16798 ( .C1(n22655), .C2(n22726), .A(n14835), .B(n14834), .ZN(
        P1_U3079) );
  NAND2_X1 U16799 ( .A1(n22723), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n14839) );
  OAI22_X1 U16800 ( .A1(n22499), .A2(n22490), .B1(n22477), .B2(n14836), .ZN(
        n14837) );
  AOI21_X1 U16801 ( .B1(n22730), .B2(n22465), .A(n14837), .ZN(n14838) );
  OAI211_X1 U16802 ( .C1(n22407), .C2(n22726), .A(n14839), .B(n14838), .ZN(
        P1_U3073) );
  NOR3_X1 U16803 ( .A1(n18000), .A2(n15215), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14843) );
  INV_X1 U16804 ( .A(n22472), .ZN(n15213) );
  INV_X1 U16805 ( .A(n14843), .ZN(n22476) );
  NOR2_X1 U16806 ( .A1(n22457), .A2(n22476), .ZN(n22778) );
  AOI21_X1 U16807 ( .B1(n15213), .B2(n15038), .A(n22778), .ZN(n14842) );
  OAI211_X1 U16808 ( .C1(n14841), .C2(n22305), .A(n22434), .B(n14842), .ZN(
        n14840) );
  OAI211_X1 U16809 ( .C1(n22434), .C2(n14843), .A(n14840), .B(n15035), .ZN(
        n22780) );
  NAND2_X1 U16810 ( .A1(n22780), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n14847) );
  NOR2_X2 U16811 ( .A1(n14841), .A2(n15002), .ZN(n22787) );
  INV_X1 U16812 ( .A(n14842), .ZN(n14844) );
  AOI22_X1 U16813 ( .A1(n14844), .A2(n22434), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14843), .ZN(n22520) );
  INV_X1 U16814 ( .A(n22778), .ZN(n14851) );
  OAI22_X1 U16815 ( .A1(n22520), .A2(n22490), .B1(n22477), .B2(n14851), .ZN(
        n14845) );
  AOI21_X1 U16816 ( .B1(n22787), .B2(n22465), .A(n14845), .ZN(n14846) );
  OAI211_X1 U16817 ( .C1(n22407), .C2(n22783), .A(n14847), .B(n14846), .ZN(
        P1_U3137) );
  NAND2_X1 U16818 ( .A1(n22780), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n14850) );
  OAI22_X1 U16819 ( .A1(n22520), .A2(n22677), .B1(n22671), .B2(n14851), .ZN(
        n14848) );
  AOI21_X1 U16820 ( .B1(n22787), .B2(n22665), .A(n14848), .ZN(n14849) );
  OAI211_X1 U16821 ( .C1(n22655), .C2(n22783), .A(n14850), .B(n14849), .ZN(
        P1_U3143) );
  NAND2_X1 U16822 ( .A1(n22780), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n14854) );
  OAI22_X1 U16823 ( .A1(n22520), .A2(n22583), .B1(n22577), .B2(n14851), .ZN(
        n14852) );
  AOI21_X1 U16824 ( .B1(n22787), .B2(n22571), .A(n14852), .ZN(n14853) );
  OAI211_X1 U16825 ( .C1(n22564), .C2(n22783), .A(n14854), .B(n14853), .ZN(
        P1_U3140) );
  MUX2_X1 U16826 ( .A(n16297), .B(n16321), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n14855) );
  OAI21_X1 U16827 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16323), .A(
        n14855), .ZN(n14931) );
  INV_X1 U16828 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17077) );
  NAND2_X1 U16829 ( .A1(n14857), .A2(n17077), .ZN(n14858) );
  OAI211_X1 U16830 ( .C1(P1_EBX_REG_4__SCAN_IN), .C2(n11150), .A(n14858), .B(
        n16385), .ZN(n14859) );
  OAI21_X1 U16831 ( .B1(P1_EBX_REG_4__SCAN_IN), .B2(n16304), .A(n14859), .ZN(
        n14860) );
  OAI21_X1 U16832 ( .B1(n14861), .B2(n14860), .A(n15328), .ZN(n22105) );
  INV_X1 U16833 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n22104) );
  OAI222_X1 U16834 ( .A1(n22105), .A2(n16841), .B1(n22104), .B2(n20727), .C1(
        n20736), .C2(n20698), .ZN(P1_U2868) );
  XOR2_X1 U16835 ( .A(n14989), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n14866)
         );
  AOI21_X1 U16836 ( .B1(n14863), .B2(n14769), .A(n14862), .ZN(n17644) );
  INV_X1 U16837 ( .A(n17644), .ZN(n19144) );
  INV_X1 U16838 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n14864) );
  MUX2_X1 U16839 ( .A(n19144), .B(n14864), .S(n17423), .Z(n14865) );
  OAI21_X1 U16840 ( .B1(n14866), .B2(n17428), .A(n14865), .ZN(P2_U2880) );
  XNOR2_X1 U16841 ( .A(n14868), .B(n14867), .ZN(n22094) );
  INV_X1 U16842 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20612) );
  OAI222_X1 U16843 ( .A1(n22094), .A2(n16897), .B1(n16056), .B2(n14869), .C1(
        n16054), .C2(n20612), .ZN(P1_U2901) );
  NOR2_X1 U16844 ( .A1(n17330), .A2(n14874), .ZN(n14870) );
  NOR2_X1 U16845 ( .A1(n22441), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14876) );
  OAI21_X1 U16846 ( .B1(n14870), .B2(n14876), .A(n15035), .ZN(n22739) );
  INV_X1 U16847 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14887) );
  INV_X1 U16848 ( .A(DATAI_20_), .ZN(n14872) );
  INV_X1 U16849 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20805) );
  OR2_X1 U16850 ( .A1(n22686), .A2(n20805), .ZN(n14871) );
  OAI21_X1 U16851 ( .B1(n22688), .B2(n14872), .A(n14871), .ZN(n22616) );
  INV_X1 U16852 ( .A(DATAI_28_), .ZN(n14875) );
  INV_X1 U16853 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20822) );
  OAI22_X1 U16854 ( .A1(n14875), .A2(n22688), .B1(n20822), .B2(n22686), .ZN(
        n22608) );
  INV_X1 U16855 ( .A(n22608), .ZN(n22619) );
  NAND2_X1 U16856 ( .A1(n22438), .A2(n15022), .ZN(n14880) );
  INV_X1 U16857 ( .A(n14876), .ZN(n14877) );
  OAI22_X1 U16858 ( .A1(n22735), .A2(n22468), .B1(n14877), .B2(n22424), .ZN(
        n14878) );
  INV_X1 U16859 ( .A(n14878), .ZN(n14879) );
  NAND2_X1 U16860 ( .A1(n14880), .A2(n14879), .ZN(n22737) );
  NOR2_X1 U16861 ( .A1(n22678), .A2(n14881), .ZN(n22615) );
  NAND2_X1 U16862 ( .A1(n14882), .A2(n22682), .ZN(n22605) );
  NOR2_X1 U16863 ( .A1(n22605), .A2(n22735), .ZN(n14883) );
  AOI21_X1 U16864 ( .B1(n22737), .B2(n22615), .A(n14883), .ZN(n14884) );
  OAI21_X1 U16865 ( .B1(n22728), .B2(n22619), .A(n14884), .ZN(n14885) );
  AOI21_X1 U16866 ( .B1(n22746), .B2(n22616), .A(n14885), .ZN(n14886) );
  OAI21_X1 U16867 ( .B1(n14930), .B2(n14887), .A(n14886), .ZN(P1_U3093) );
  INV_X1 U16868 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14892) );
  NOR2_X1 U16869 ( .A1(n22671), .A2(n22735), .ZN(n14888) );
  AOI21_X1 U16870 ( .B1(n22737), .B2(n15248), .A(n14888), .ZN(n14889) );
  OAI21_X1 U16871 ( .B1(n22728), .B2(n22655), .A(n14889), .ZN(n14890) );
  AOI21_X1 U16872 ( .B1(n22746), .B2(n22665), .A(n14890), .ZN(n14891) );
  OAI21_X1 U16873 ( .B1(n14930), .B2(n14892), .A(n14891), .ZN(P1_U3095) );
  INV_X1 U16874 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14901) );
  INV_X1 U16875 ( .A(DATAI_26_), .ZN(n14893) );
  INV_X1 U16876 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20818) );
  OAI22_X1 U16877 ( .A1(n14893), .A2(n22688), .B1(n20818), .B2(n22686), .ZN(
        n22549) );
  NAND2_X1 U16878 ( .A1(n12886), .A2(n22682), .ZN(n22546) );
  NOR2_X1 U16879 ( .A1(n22678), .A2(n14894), .ZN(n22556) );
  NAND2_X1 U16880 ( .A1(n22737), .A2(n22556), .ZN(n14895) );
  OAI21_X1 U16881 ( .B1(n22546), .B2(n22735), .A(n14895), .ZN(n14899) );
  NAND2_X1 U16882 ( .A1(n14904), .A2(DATAI_18_), .ZN(n14897) );
  INV_X1 U16883 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20801) );
  OR2_X1 U16884 ( .A1(n22686), .A2(n20801), .ZN(n14896) );
  AND2_X1 U16885 ( .A1(n14897), .A2(n14896), .ZN(n22547) );
  NOR2_X1 U16886 ( .A1(n22742), .A2(n22547), .ZN(n14898) );
  AOI211_X1 U16887 ( .C1(n22738), .C2(n22549), .A(n14899), .B(n14898), .ZN(
        n14900) );
  OAI21_X1 U16888 ( .B1(n14930), .B2(n14901), .A(n14900), .ZN(P1_U3091) );
  INV_X1 U16889 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14910) );
  INV_X1 U16890 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20824) );
  INV_X1 U16891 ( .A(DATAI_29_), .ZN(n14902) );
  OAI22_X1 U16892 ( .A1(n20824), .A2(n22686), .B1(n14902), .B2(n22688), .ZN(
        n22643) );
  NAND2_X1 U16893 ( .A1(n11160), .A2(n22682), .ZN(n22640) );
  NOR2_X1 U16894 ( .A1(n22678), .A2(n14985), .ZN(n22650) );
  NAND2_X1 U16895 ( .A1(n22737), .A2(n22650), .ZN(n14903) );
  OAI21_X1 U16896 ( .B1(n22640), .B2(n22735), .A(n14903), .ZN(n14908) );
  NAND2_X1 U16897 ( .A1(n14904), .A2(DATAI_21_), .ZN(n14906) );
  INV_X1 U16898 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20807) );
  OR2_X1 U16899 ( .A1(n22686), .A2(n20807), .ZN(n14905) );
  AND2_X1 U16900 ( .A1(n14906), .A2(n14905), .ZN(n22641) );
  NOR2_X1 U16901 ( .A1(n22742), .A2(n22641), .ZN(n14907) );
  AOI211_X1 U16902 ( .C1(n22738), .C2(n22643), .A(n14908), .B(n14907), .ZN(
        n14909) );
  OAI21_X1 U16903 ( .B1(n14930), .B2(n14910), .A(n14909), .ZN(P1_U3094) );
  INV_X1 U16904 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14919) );
  INV_X1 U16905 ( .A(DATAI_17_), .ZN(n14912) );
  INV_X1 U16906 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20799) );
  OR2_X1 U16907 ( .A1(n22686), .A2(n20799), .ZN(n14911) );
  OAI21_X1 U16908 ( .B1(n22688), .B2(n14912), .A(n14911), .ZN(n22525) );
  INV_X1 U16909 ( .A(DATAI_25_), .ZN(n14913) );
  INV_X1 U16910 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20816) );
  OAI22_X1 U16911 ( .A1(n14913), .A2(n22688), .B1(n20816), .B2(n22686), .ZN(
        n22516) );
  INV_X1 U16912 ( .A(n22516), .ZN(n22528) );
  NOR2_X1 U16913 ( .A1(n22678), .A2(n14914), .ZN(n22524) );
  NAND2_X1 U16914 ( .A1(n12947), .A2(n22682), .ZN(n22513) );
  NOR2_X1 U16915 ( .A1(n22513), .A2(n22735), .ZN(n14915) );
  AOI21_X1 U16916 ( .B1(n22737), .B2(n22524), .A(n14915), .ZN(n14916) );
  OAI21_X1 U16917 ( .B1(n22728), .B2(n22528), .A(n14916), .ZN(n14917) );
  AOI21_X1 U16918 ( .B1(n22746), .B2(n22525), .A(n14917), .ZN(n14918) );
  OAI21_X1 U16919 ( .B1(n14930), .B2(n14919), .A(n14918), .ZN(P1_U3090) );
  INV_X1 U16920 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14924) );
  NOR2_X1 U16921 ( .A1(n22577), .A2(n22735), .ZN(n14920) );
  AOI21_X1 U16922 ( .B1(n22737), .B2(n15231), .A(n14920), .ZN(n14921) );
  OAI21_X1 U16923 ( .B1(n22728), .B2(n22564), .A(n14921), .ZN(n14922) );
  AOI21_X1 U16924 ( .B1(n22746), .B2(n22571), .A(n14922), .ZN(n14923) );
  OAI21_X1 U16925 ( .B1(n14930), .B2(n14924), .A(n14923), .ZN(P1_U3092) );
  INV_X1 U16926 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14929) );
  NOR2_X1 U16927 ( .A1(n22477), .A2(n22735), .ZN(n14925) );
  AOI21_X1 U16928 ( .B1(n22737), .B2(n15222), .A(n14925), .ZN(n14926) );
  OAI21_X1 U16929 ( .B1(n22728), .B2(n22407), .A(n14926), .ZN(n14927) );
  AOI21_X1 U16930 ( .B1(n22746), .B2(n22465), .A(n14927), .ZN(n14928) );
  OAI21_X1 U16931 ( .B1(n14930), .B2(n14929), .A(n14928), .ZN(P1_U3089) );
  XNOR2_X1 U16932 ( .A(n14856), .B(n14931), .ZN(n22103) );
  INV_X1 U16933 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n14932) );
  OAI222_X1 U16934 ( .A1(n22103), .A2(n16841), .B1(n20727), .B2(n14932), .C1(
        n22094), .C2(n20698), .ZN(P1_U2869) );
  INV_X1 U16935 ( .A(n15602), .ZN(n14938) );
  NAND2_X1 U16936 ( .A1(n14934), .A2(n14933), .ZN(n15290) );
  INV_X1 U16937 ( .A(n15289), .ZN(n14935) );
  XNOR2_X1 U16938 ( .A(n15290), .B(n14935), .ZN(n14936) );
  NAND2_X1 U16939 ( .A1(n14936), .A2(n15607), .ZN(n14937) );
  INV_X1 U16940 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n22011) );
  XNOR2_X1 U16941 ( .A(n15285), .B(n22011), .ZN(n14942) );
  NAND2_X1 U16942 ( .A1(n14940), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14941) );
  NAND2_X1 U16943 ( .A1(n21990), .A2(n14941), .ZN(n14943) );
  OR2_X1 U16944 ( .A1(n14942), .A2(n14943), .ZN(n14944) );
  NAND2_X1 U16945 ( .A1(n14943), .A2(n14942), .ZN(n15287) );
  AND2_X1 U16946 ( .A1(n14944), .A2(n15287), .ZN(n22008) );
  NAND2_X1 U16947 ( .A1(n20761), .A2(n22097), .ZN(n14945) );
  INV_X1 U16948 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n22090) );
  OR2_X1 U16949 ( .A1(n22066), .A2(n22090), .ZN(n22005) );
  OAI211_X1 U16950 ( .C1(n20728), .C2(n14946), .A(n14945), .B(n22005), .ZN(
        n14947) );
  AOI21_X1 U16951 ( .B1(n22008), .B2(n20756), .A(n14947), .ZN(n14948) );
  OAI21_X1 U16952 ( .B1(n17060), .B2(n22094), .A(n14948), .ZN(P1_U2996) );
  INV_X1 U16953 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14950) );
  AOI22_X1 U16954 ( .A1(n20633), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n14949) );
  OAI21_X1 U16955 ( .B1(n14950), .B2(n14974), .A(n14949), .ZN(P1_U2913) );
  AOI22_X1 U16956 ( .A1(n20633), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n14951) );
  OAI21_X1 U16957 ( .B1(n14952), .B2(n14974), .A(n14951), .ZN(P1_U2906) );
  AOI22_X1 U16958 ( .A1(n20633), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n14953) );
  OAI21_X1 U16959 ( .B1(n14954), .B2(n14974), .A(n14953), .ZN(P1_U2907) );
  AOI22_X1 U16960 ( .A1(n20633), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n14955) );
  OAI21_X1 U16961 ( .B1(n14956), .B2(n14974), .A(n14955), .ZN(P1_U2911) );
  AOI22_X1 U16962 ( .A1(n20633), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n14957) );
  OAI21_X1 U16963 ( .B1(n14958), .B2(n14974), .A(n14957), .ZN(P1_U2908) );
  INV_X1 U16964 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14960) );
  AOI22_X1 U16965 ( .A1(n20633), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n14959) );
  OAI21_X1 U16966 ( .B1(n14960), .B2(n14974), .A(n14959), .ZN(P1_U2912) );
  AOI22_X1 U16967 ( .A1(n20633), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n14961) );
  OAI21_X1 U16968 ( .B1(n14962), .B2(n14974), .A(n14961), .ZN(P1_U2909) );
  AOI22_X1 U16969 ( .A1(n20633), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n14963) );
  OAI21_X1 U16970 ( .B1(n14964), .B2(n14974), .A(n14963), .ZN(P1_U2914) );
  INV_X1 U16971 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14966) );
  AOI22_X1 U16972 ( .A1(n20633), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n14965) );
  OAI21_X1 U16973 ( .B1(n14966), .B2(n14974), .A(n14965), .ZN(P1_U2915) );
  INV_X1 U16974 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14968) );
  AOI22_X1 U16975 ( .A1(n20633), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n14967) );
  OAI21_X1 U16976 ( .B1(n14968), .B2(n14974), .A(n14967), .ZN(P1_U2916) );
  INV_X1 U16977 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14970) );
  AOI22_X1 U16978 ( .A1(n20633), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n14969) );
  OAI21_X1 U16979 ( .B1(n14970), .B2(n14974), .A(n14969), .ZN(P1_U2917) );
  AOI22_X1 U16980 ( .A1(n20633), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n14971) );
  OAI21_X1 U16981 ( .B1(n14972), .B2(n14974), .A(n14971), .ZN(P1_U2910) );
  INV_X1 U16982 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n14975) );
  AOI22_X1 U16983 ( .A1(n20633), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n20632), .ZN(n14973) );
  OAI21_X1 U16984 ( .B1(n14975), .B2(n14974), .A(n14973), .ZN(P1_U2920) );
  AOI21_X1 U16985 ( .B1(n19103), .B2(n18128), .A(n14976), .ZN(n15203) );
  XOR2_X1 U16986 ( .A(n18120), .B(n15203), .Z(n15202) );
  XNOR2_X1 U16987 ( .A(n15202), .B(n16017), .ZN(n14977) );
  NAND2_X1 U16988 ( .A1(n14977), .A2(n20322), .ZN(n14979) );
  AOI22_X1 U16989 ( .A1(n20321), .A2(n18120), .B1(n20319), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n14978) );
  OAI211_X1 U16990 ( .C1(n20328), .C2(n15324), .A(n14979), .B(n14978), .ZN(
        P2_U2917) );
  OR2_X1 U16991 ( .A1(n14814), .A2(n14982), .ZN(n14983) );
  AND2_X1 U16992 ( .A1(n14981), .A2(n14983), .ZN(n22126) );
  INV_X1 U16993 ( .A(n22126), .ZN(n14986) );
  INV_X1 U16994 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n14984) );
  OAI222_X1 U16995 ( .A1(n14986), .A2(n16897), .B1(n16056), .B2(n14985), .C1(
        n14984), .C2(n16054), .ZN(P1_U2899) );
  OR2_X1 U16996 ( .A1(n14987), .A2(n14862), .ZN(n14988) );
  AND2_X1 U16997 ( .A1(n15194), .A2(n14988), .ZN(n19397) );
  INV_X1 U16998 ( .A(n19397), .ZN(n14994) );
  INV_X1 U16999 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n20113) );
  INV_X1 U17000 ( .A(n15191), .ZN(n14990) );
  OAI211_X1 U17001 ( .C1(n11234), .C2(n14991), .A(n14990), .B(n17417), .ZN(
        n14993) );
  NAND2_X1 U17002 ( .A1(n17423), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14992) );
  OAI211_X1 U17003 ( .C1(n14994), .C2(n17420), .A(n14993), .B(n14992), .ZN(
        P2_U2879) );
  INV_X1 U17004 ( .A(n17431), .ZN(n14998) );
  AOI21_X1 U17005 ( .B1(n14996), .B2(n14820), .A(n14995), .ZN(n19383) );
  INV_X1 U17006 ( .A(n19383), .ZN(n14997) );
  INV_X1 U17007 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n18174) );
  OAI222_X1 U17008 ( .A1(n15324), .A2(n14998), .B1(n14997), .B2(n20171), .C1(
        n17475), .C2(n18174), .ZN(P2_U2907) );
  INV_X1 U17009 ( .A(n11195), .ZN(n14999) );
  INV_X1 U17010 ( .A(n15037), .ZN(n15000) );
  NOR3_X1 U17011 ( .A1(n15215), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15004) );
  INV_X1 U17012 ( .A(n15020), .ZN(n15017) );
  AND2_X1 U17013 ( .A1(n14427), .A2(n22418), .ZN(n22452) );
  INV_X1 U17014 ( .A(n15004), .ZN(n15253) );
  NOR2_X1 U17015 ( .A1(n22457), .A2(n15253), .ZN(n22750) );
  AOI21_X1 U17016 ( .B1(n22452), .B2(n15038), .A(n22750), .ZN(n15003) );
  OAI211_X1 U17017 ( .C1(n15017), .C2(n22305), .A(n22434), .B(n15003), .ZN(
        n15001) );
  OAI211_X1 U17018 ( .C1(n22434), .C2(n15004), .A(n15001), .B(n15035), .ZN(
        n22752) );
  NAND2_X1 U17019 ( .A1(n22752), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n15008) );
  INV_X1 U17020 ( .A(n15003), .ZN(n15005) );
  AOI22_X1 U17021 ( .A1(n15005), .A2(n22434), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15004), .ZN(n22504) );
  INV_X1 U17022 ( .A(n22750), .ZN(n15013) );
  OAI22_X1 U17023 ( .A1(n22504), .A2(n22583), .B1(n22577), .B2(n15013), .ZN(
        n15006) );
  AOI21_X1 U17024 ( .B1(n22758), .B2(n22571), .A(n15006), .ZN(n15007) );
  OAI211_X1 U17025 ( .C1(n22564), .C2(n22755), .A(n15008), .B(n15007), .ZN(
        P1_U3108) );
  INV_X1 U17026 ( .A(n22465), .ZN(n22478) );
  INV_X1 U17027 ( .A(n22758), .ZN(n15012) );
  NAND2_X1 U17028 ( .A1(n22752), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n15011) );
  INV_X1 U17029 ( .A(n22755), .ZN(n15254) );
  OAI22_X1 U17030 ( .A1(n22504), .A2(n22490), .B1(n22477), .B2(n15013), .ZN(
        n15009) );
  AOI21_X1 U17031 ( .B1(n15254), .B2(n22487), .A(n15009), .ZN(n15010) );
  OAI211_X1 U17032 ( .C1(n22478), .C2(n15012), .A(n15011), .B(n15010), .ZN(
        P1_U3105) );
  NAND2_X1 U17033 ( .A1(n22752), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n15016) );
  OAI22_X1 U17034 ( .A1(n22504), .A2(n22677), .B1(n22671), .B2(n15013), .ZN(
        n15014) );
  AOI21_X1 U17035 ( .B1(n22758), .B2(n22665), .A(n15014), .ZN(n15015) );
  OAI211_X1 U17036 ( .C1(n22655), .C2(n22755), .A(n15016), .B(n15015), .ZN(
        P1_U3111) );
  NOR2_X1 U17037 ( .A1(n15017), .A2(n17330), .ZN(n15018) );
  NOR3_X1 U17038 ( .A1(n15215), .A2(n22406), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22456) );
  OAI21_X1 U17039 ( .B1(n15018), .B2(n22456), .A(n15035), .ZN(n22765) );
  NAND2_X1 U17040 ( .A1(n22765), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n15025) );
  INV_X1 U17041 ( .A(n22456), .ZN(n15021) );
  NOR2_X1 U17042 ( .A1(n22457), .A2(n15021), .ZN(n22763) );
  AOI222_X1 U17043 ( .A1(n22456), .A2(P1_STATE2_REG_2__SCAN_IN), .B1(n22452), 
        .B2(n15022), .C1(n22434), .C2(n22763), .ZN(n22510) );
  INV_X1 U17044 ( .A(n22763), .ZN(n15029) );
  OAI22_X1 U17045 ( .A1(n22510), .A2(n22677), .B1(n22671), .B2(n15029), .ZN(
        n15023) );
  AOI21_X1 U17046 ( .B1(n22772), .B2(n22665), .A(n15023), .ZN(n15024) );
  OAI211_X1 U17047 ( .C1(n22655), .C2(n22768), .A(n15025), .B(n15024), .ZN(
        P1_U3127) );
  NAND2_X1 U17048 ( .A1(n22765), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n15028) );
  OAI22_X1 U17049 ( .A1(n22510), .A2(n22490), .B1(n22477), .B2(n15029), .ZN(
        n15026) );
  AOI21_X1 U17050 ( .B1(n22772), .B2(n22465), .A(n15026), .ZN(n15027) );
  OAI211_X1 U17051 ( .C1(n22407), .C2(n22768), .A(n15028), .B(n15027), .ZN(
        P1_U3121) );
  NAND2_X1 U17052 ( .A1(n22765), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n15032) );
  OAI22_X1 U17053 ( .A1(n22510), .A2(n22583), .B1(n22577), .B2(n15029), .ZN(
        n15030) );
  AOI21_X1 U17054 ( .B1(n22772), .B2(n22571), .A(n15030), .ZN(n15031) );
  OAI211_X1 U17055 ( .C1(n22564), .C2(n22768), .A(n15032), .B(n15031), .ZN(
        P1_U3124) );
  NOR3_X1 U17056 ( .A1(n22423), .A2(n22468), .A3(n22305), .ZN(n15036) );
  NOR3_X1 U17057 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22391) );
  NAND2_X1 U17058 ( .A1(n22698), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n15044) );
  NAND2_X1 U17059 ( .A1(n22418), .A2(n15038), .ZN(n15040) );
  INV_X1 U17060 ( .A(n22391), .ZN(n15039) );
  NOR2_X1 U17061 ( .A1(n22457), .A2(n15039), .ZN(n22695) );
  INV_X1 U17062 ( .A(n22695), .ZN(n15060) );
  OAI21_X1 U17063 ( .B1(n14427), .B2(n15040), .A(n15060), .ZN(n15041) );
  AOI22_X1 U17064 ( .A1(n15041), .A2(n22434), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n22391), .ZN(n22694) );
  OAI22_X1 U17065 ( .A1(n22694), .A2(n22583), .B1(n22577), .B2(n15060), .ZN(
        n15042) );
  AOI21_X1 U17066 ( .B1(n22697), .B2(n22580), .A(n15042), .ZN(n15043) );
  OAI211_X1 U17067 ( .C1(n22578), .C2(n22701), .A(n15044), .B(n15043), .ZN(
        P1_U3044) );
  NAND2_X1 U17068 ( .A1(n22698), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n15047) );
  OAI22_X1 U17069 ( .A1(n22694), .A2(n22677), .B1(n22671), .B2(n15060), .ZN(
        n15045) );
  AOI21_X1 U17070 ( .B1(n22697), .B2(n22674), .A(n15045), .ZN(n15046) );
  OAI211_X1 U17071 ( .C1(n22672), .C2(n22701), .A(n15047), .B(n15046), .ZN(
        P1_U3047) );
  NAND2_X1 U17072 ( .A1(n22698), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n15050) );
  OAI22_X1 U17073 ( .A1(n22694), .A2(n22490), .B1(n22477), .B2(n15060), .ZN(
        n15048) );
  AOI21_X1 U17074 ( .B1(n22697), .B2(n22487), .A(n15048), .ZN(n15049) );
  OAI211_X1 U17075 ( .C1(n22478), .C2(n22701), .A(n15050), .B(n15049), .ZN(
        P1_U3041) );
  NAND2_X1 U17076 ( .A1(n22698), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n15053) );
  INV_X1 U17077 ( .A(n22556), .ZN(n22552) );
  OAI22_X1 U17078 ( .A1(n22694), .A2(n22552), .B1(n22546), .B2(n15060), .ZN(
        n15051) );
  AOI21_X1 U17079 ( .B1(n22697), .B2(n22549), .A(n15051), .ZN(n15052) );
  OAI211_X1 U17080 ( .C1(n22547), .C2(n22701), .A(n15053), .B(n15052), .ZN(
        P1_U3043) );
  NAND2_X1 U17081 ( .A1(n22698), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n15056) );
  INV_X1 U17082 ( .A(n22650), .ZN(n22646) );
  OAI22_X1 U17083 ( .A1(n22694), .A2(n22646), .B1(n22640), .B2(n15060), .ZN(
        n15054) );
  AOI21_X1 U17084 ( .B1(n22697), .B2(n22643), .A(n15054), .ZN(n15055) );
  OAI211_X1 U17085 ( .C1(n22641), .C2(n22701), .A(n15056), .B(n15055), .ZN(
        P1_U3046) );
  INV_X1 U17086 ( .A(n22616), .ZN(n22606) );
  NAND2_X1 U17087 ( .A1(n22698), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n15059) );
  INV_X1 U17088 ( .A(n22615), .ZN(n22611) );
  OAI22_X1 U17089 ( .A1(n22694), .A2(n22611), .B1(n22605), .B2(n15060), .ZN(
        n15057) );
  AOI21_X1 U17090 ( .B1(n22697), .B2(n22608), .A(n15057), .ZN(n15058) );
  OAI211_X1 U17091 ( .C1(n22606), .C2(n22701), .A(n15059), .B(n15058), .ZN(
        P1_U3045) );
  INV_X1 U17092 ( .A(n22525), .ZN(n22514) );
  NAND2_X1 U17093 ( .A1(n22698), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n15063) );
  INV_X1 U17094 ( .A(n22524), .ZN(n22519) );
  OAI22_X1 U17095 ( .A1(n22694), .A2(n22519), .B1(n22513), .B2(n15060), .ZN(
        n15061) );
  AOI21_X1 U17096 ( .B1(n22697), .B2(n22516), .A(n15061), .ZN(n15062) );
  OAI211_X1 U17097 ( .C1(n22514), .C2(n22701), .A(n15063), .B(n15062), .ZN(
        P1_U3042) );
  OAI211_X1 U17098 ( .C1(P1_STATE2_REG_0__SCAN_IN), .C2(n22305), .A(
        P1_STATE2_REG_1__SCAN_IN), .B(n22424), .ZN(n18019) );
  NOR2_X1 U17099 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22297) );
  NAND2_X1 U17100 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n22297), .ZN(n18018) );
  OAI221_X1 U17101 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n18019), .C1(n22287), 
        .C2(n18018), .A(n21967), .ZN(n15066) );
  NAND2_X1 U17102 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15066), .ZN(n15071) );
  INV_X1 U17103 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16327) );
  INV_X1 U17104 ( .A(n15066), .ZN(n15067) );
  NAND2_X1 U17105 ( .A1(n22091), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15068) );
  OAI21_X1 U17106 ( .B1(n15071), .B2(n11359), .A(n22269), .ZN(n22125) );
  INV_X1 U17107 ( .A(n22125), .ZN(n22095) );
  INV_X1 U17108 ( .A(n15068), .ZN(n15069) );
  INV_X1 U17109 ( .A(n22091), .ZN(n16309) );
  NOR2_X1 U17110 ( .A1(n15070), .A2(n15071), .ZN(n22108) );
  INV_X1 U17111 ( .A(n22108), .ZN(n15182) );
  NAND2_X1 U17112 ( .A1(n22322), .A2(n22305), .ZN(n17981) );
  INV_X1 U17113 ( .A(n15071), .ZN(n15074) );
  AND3_X1 U17114 ( .A1(n17981), .A2(P1_EBX_REG_31__SCAN_IN), .A3(n15074), .ZN(
        n15072) );
  OR2_X1 U17115 ( .A1(n15073), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15079) );
  INV_X1 U17116 ( .A(n15079), .ZN(n15075) );
  AND2_X1 U17117 ( .A1(n16710), .A2(n15074), .ZN(n15077) );
  NAND2_X2 U17118 ( .A1(n15075), .A2(n15077), .ZN(n22245) );
  NAND2_X1 U17119 ( .A1(n12947), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n15076) );
  AND2_X1 U17120 ( .A1(n15077), .A2(n15076), .ZN(n15078) );
  OAI22_X1 U17121 ( .A1(n22245), .A2(P1_REIP_REG_1__SCAN_IN), .B1(n22262), 
        .B2(n15080), .ZN(n15081) );
  AOI21_X1 U17122 ( .B1(n15082), .B2(n22217), .A(n15081), .ZN(n15083) );
  OAI21_X1 U17123 ( .B1(n11193), .B2(n15182), .A(n15083), .ZN(n15084) );
  AOI21_X1 U17124 ( .B1(n16309), .B2(P1_REIP_REG_1__SCAN_IN), .A(n15084), .ZN(
        n15086) );
  NAND2_X1 U17125 ( .A1(n22264), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15085) );
  NAND2_X1 U17126 ( .A1(n15086), .A2(n15085), .ZN(n15087) );
  AOI21_X1 U17127 ( .B1(n22266), .B2(n15088), .A(n15087), .ZN(n15089) );
  OAI21_X1 U17128 ( .B1(n22095), .B2(n15090), .A(n15089), .ZN(P1_U2839) );
  NAND2_X1 U17129 ( .A1(n22099), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n15094) );
  NAND2_X1 U17130 ( .A1(n22236), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n15093) );
  OAI21_X1 U17131 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n22245), .A(n22091), .ZN(
        n15091) );
  NAND2_X1 U17132 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n15091), .ZN(n15092) );
  OAI211_X1 U17133 ( .C1(n22245), .C2(n15094), .A(n15093), .B(n15092), .ZN(
        n15095) );
  AOI21_X1 U17134 ( .B1(n21995), .B2(n22217), .A(n15095), .ZN(n15096) );
  OAI21_X1 U17135 ( .B1(n22418), .B2(n15182), .A(n15096), .ZN(n15097) );
  AOI21_X1 U17136 ( .B1(n22264), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n15097), .ZN(n15100) );
  NAND2_X1 U17137 ( .A1(n22125), .A2(n15098), .ZN(n15099) );
  OAI211_X1 U17138 ( .C1(n22257), .C2(n15101), .A(n15100), .B(n15099), .ZN(
        P1_U2838) );
  INV_X1 U17139 ( .A(n15102), .ZN(n15103) );
  NAND2_X1 U17140 ( .A1(n15103), .A2(n15164), .ZN(n15111) );
  INV_X1 U17141 ( .A(n15165), .ZN(n15105) );
  OAI21_X1 U17142 ( .B1(n15166), .B2(n15105), .A(n15104), .ZN(n15106) );
  INV_X1 U17143 ( .A(n15106), .ZN(n15107) );
  AND2_X1 U17144 ( .A1(n15108), .A2(n15107), .ZN(n15110) );
  INV_X1 U17145 ( .A(n15150), .ZN(n15132) );
  INV_X1 U17146 ( .A(n15112), .ZN(n15114) );
  NAND2_X1 U17147 ( .A1(n15114), .A2(n15113), .ZN(n15118) );
  INV_X1 U17148 ( .A(n15118), .ZN(n15116) );
  INV_X1 U17149 ( .A(n15115), .ZN(n15144) );
  MUX2_X1 U17150 ( .A(n15116), .B(n15144), .S(n19360), .Z(n15117) );
  OAI21_X1 U17151 ( .B1(n16344), .B2(n15132), .A(n15117), .ZN(n19355) );
  NAND2_X1 U17152 ( .A1(n19105), .A2(n15150), .ZN(n15120) );
  OAI21_X1 U17153 ( .B1(n11864), .B2(n11849), .A(n15118), .ZN(n15119) );
  OAI211_X1 U17154 ( .C1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n15144), .A(
        n15120), .B(n15119), .ZN(n16165) );
  OAI21_X1 U17155 ( .B1(n15121), .B2(n19355), .A(n16165), .ZN(n15123) );
  OAI21_X1 U17156 ( .B1(n19355), .B2(n20094), .A(n20092), .ZN(n15122) );
  AOI21_X1 U17157 ( .B1(n15123), .B2(n15122), .A(n16063), .ZN(n15137) );
  INV_X1 U17158 ( .A(n15137), .ZN(n15135) );
  INV_X1 U17159 ( .A(n15163), .ZN(n15124) );
  NAND2_X1 U17160 ( .A1(n15161), .A2(n15124), .ZN(n15141) );
  INV_X1 U17161 ( .A(n11850), .ZN(n15125) );
  NAND2_X1 U17162 ( .A1(n15125), .A2(n11830), .ZN(n15142) );
  NAND2_X1 U17163 ( .A1(n15126), .A2(n15142), .ZN(n15130) );
  XNOR2_X1 U17164 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15128) );
  NOR2_X1 U17165 ( .A1(n11164), .A2(n15127), .ZN(n15138) );
  OAI22_X1 U17166 ( .A1(n15144), .A2(n15128), .B1(n15138), .B2(n15130), .ZN(
        n15129) );
  AOI21_X1 U17167 ( .B1(n15141), .B2(n15130), .A(n15129), .ZN(n15131) );
  OAI21_X1 U17168 ( .B1(n15133), .B2(n15132), .A(n15131), .ZN(n16062) );
  NAND2_X1 U17169 ( .A1(n16063), .A2(n11830), .ZN(n15134) );
  OAI21_X1 U17170 ( .B1(n16062), .B2(n16063), .A(n15134), .ZN(n15172) );
  OAI21_X1 U17171 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15135), .A(
        n15172), .ZN(n15136) );
  OAI21_X1 U17172 ( .B1(n15137), .B2(n19998), .A(n15136), .ZN(n15152) );
  NAND2_X1 U17173 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15143) );
  INV_X1 U17174 ( .A(n15143), .ZN(n15140) );
  OR2_X1 U17175 ( .A1(n15138), .A2(n16676), .ZN(n15139) );
  OAI211_X1 U17176 ( .C1(n15144), .C2(n15140), .A(n15139), .B(n15142), .ZN(
        n15148) );
  INV_X1 U17177 ( .A(n15141), .ZN(n15146) );
  INV_X1 U17178 ( .A(n15142), .ZN(n15145) );
  OAI22_X1 U17179 ( .A1(n15146), .A2(n15145), .B1(n15144), .B2(n15143), .ZN(
        n15147) );
  MUX2_X1 U17180 ( .A(n15148), .B(n15147), .S(n11571), .Z(n15149) );
  AOI211_X1 U17181 ( .C1(n12303), .C2(n15150), .A(n16481), .B(n15149), .ZN(
        n17932) );
  MUX2_X1 U17182 ( .A(n17932), .B(n11571), .S(n16063), .Z(n15173) );
  OR2_X1 U17183 ( .A1(n15173), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15151) );
  AOI221_X1 U17184 ( .B1(n15152), .B2(n15151), .C1(n15173), .C2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15175) );
  INV_X1 U17185 ( .A(n17965), .ZN(n15154) );
  AOI22_X1 U17186 ( .A1(n15156), .A2(n15155), .B1(n15154), .B2(n15153), .ZN(
        n15160) );
  NAND2_X1 U17187 ( .A1(n15158), .A2(n15157), .ZN(n15159) );
  OAI211_X1 U17188 ( .C1(n16020), .C2(n15161), .A(n15160), .B(n15159), .ZN(
        n15162) );
  AOI21_X1 U17189 ( .B1(n15163), .B2(n16020), .A(n15162), .ZN(n19447) );
  NOR3_X1 U17190 ( .A1(n15166), .A2(n15165), .A3(n15164), .ZN(n19449) );
  OR2_X1 U17191 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n15170) );
  INV_X1 U17192 ( .A(n15167), .ZN(n15168) );
  NOR3_X1 U17193 ( .A1(n11846), .A2(n15168), .A3(n19079), .ZN(n19361) );
  AOI211_X1 U17194 ( .C1(n19449), .C2(n15170), .A(n19361), .B(n15169), .ZN(
        n15171) );
  OAI211_X1 U17195 ( .C1(n15173), .C2(n15172), .A(n19447), .B(n15171), .ZN(
        n15174) );
  AOI211_X1 U17196 ( .C1(n16063), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n15175), .B(n15174), .ZN(n19446) );
  NAND3_X1 U17197 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19446), .A3(n17963), 
        .ZN(n15179) );
  AND2_X1 U17198 ( .A1(n12601), .A2(n15176), .ZN(n15177) );
  AOI21_X1 U17199 ( .B1(n15179), .B2(n15178), .A(n15177), .ZN(n19443) );
  OAI21_X1 U17200 ( .B1(n19443), .B2(n19436), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n15180) );
  NOR2_X1 U17201 ( .A1(n19436), .A2(n18114), .ZN(n17962) );
  INV_X1 U17202 ( .A(n17962), .ZN(n17966) );
  NAND2_X1 U17203 ( .A1(n15180), .A2(n17966), .ZN(P2_U3593) );
  NAND2_X1 U17204 ( .A1(n22091), .A2(n22245), .ZN(n22210) );
  OAI22_X1 U17205 ( .A1(n22200), .A2(n20696), .B1(n22276), .B2(n15181), .ZN(
        n15185) );
  INV_X1 U17206 ( .A(n22417), .ZN(n15183) );
  NOR2_X1 U17207 ( .A1(n15183), .A2(n15182), .ZN(n15184) );
  AOI211_X1 U17208 ( .C1(n22236), .C2(P1_EBX_REG_0__SCAN_IN), .A(n15185), .B(
        n15184), .ZN(n15187) );
  OAI21_X1 U17209 ( .B1(n22266), .B2(n22264), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15186) );
  OAI211_X1 U17210 ( .C1(n22095), .C2(n20730), .A(n15187), .B(n15186), .ZN(
        P1_U2840) );
  INV_X1 U17211 ( .A(n16654), .ZN(n15189) );
  OAI21_X1 U17212 ( .B1(n14995), .B2(n15188), .A(n11231), .ZN(n19199) );
  INV_X1 U17213 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n18176) );
  OAI222_X1 U17214 ( .A1(n15324), .A2(n15189), .B1(n19199), .B2(n20171), .C1(
        n17475), .C2(n18176), .ZN(P2_U2906) );
  INV_X1 U17215 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n19150) );
  INV_X1 U17216 ( .A(n15190), .ZN(n15192) );
  OAI211_X1 U17217 ( .C1(n15191), .C2(n15192), .A(n17417), .B(n15368), .ZN(
        n15197) );
  AOI21_X1 U17218 ( .B1(n15195), .B2(n15194), .A(n15193), .ZN(n19157) );
  NAND2_X1 U17219 ( .A1(n14580), .A2(n19157), .ZN(n15196) );
  OAI211_X1 U17220 ( .C1(n14580), .C2(n19150), .A(n15197), .B(n15196), .ZN(
        P2_U2878) );
  OR2_X1 U17221 ( .A1(n15199), .A2(n15198), .ZN(n15201) );
  NAND2_X1 U17222 ( .A1(n15201), .A2(n15200), .ZN(n15389) );
  NAND2_X1 U17223 ( .A1(n15202), .A2(n18127), .ZN(n15206) );
  INV_X1 U17224 ( .A(n15389), .ZN(n19409) );
  XNOR2_X1 U17225 ( .A(n20058), .B(n19409), .ZN(n15204) );
  NAND2_X1 U17226 ( .A1(n15203), .A2(n18120), .ZN(n15205) );
  NAND3_X1 U17227 ( .A1(n15206), .A2(n15204), .A3(n15205), .ZN(n15377) );
  INV_X1 U17228 ( .A(n15377), .ZN(n15208) );
  AOI21_X1 U17229 ( .B1(n15206), .B2(n15205), .A(n15204), .ZN(n15207) );
  OAI21_X1 U17230 ( .B1(n15208), .B2(n15207), .A(n20322), .ZN(n15211) );
  INV_X1 U17231 ( .A(n16241), .ZN(n15209) );
  AOI22_X1 U17232 ( .A1(n20164), .A2(n15209), .B1(n20319), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n15210) );
  OAI211_X1 U17233 ( .C1(n15389), .C2(n17477), .A(n15211), .B(n15210), .ZN(
        P2_U2916) );
  OAI21_X1 U17234 ( .B1(n22787), .B2(n15212), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15214) );
  NAND2_X1 U17235 ( .A1(n15213), .A2(n22471), .ZN(n15221) );
  AOI21_X1 U17236 ( .B1(n15214), .B2(n15221), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n15217) );
  INV_X1 U17237 ( .A(n22404), .ZN(n15421) );
  NAND2_X1 U17238 ( .A1(n15421), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15218) );
  NAND2_X1 U17239 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15218), .ZN(n22459) );
  INV_X1 U17240 ( .A(n15219), .ZN(n15216) );
  NOR2_X1 U17241 ( .A1(n15216), .A2(n22424), .ZN(n22453) );
  NOR2_X1 U17242 ( .A1(n22453), .A2(n22678), .ZN(n22480) );
  OAI211_X1 U17243 ( .C1(n15217), .C2(n22784), .A(n22459), .B(n22480), .ZN(
        n22788) );
  NAND2_X1 U17244 ( .A1(n22787), .A2(n22487), .ZN(n15224) );
  INV_X1 U17245 ( .A(n15218), .ZN(n22454) );
  NOR2_X1 U17246 ( .A1(n15219), .A2(n22424), .ZN(n22474) );
  NAND2_X1 U17247 ( .A1(n22454), .A2(n22474), .ZN(n15220) );
  OAI21_X1 U17248 ( .B1(n15221), .B2(n22468), .A(n15220), .ZN(n22785) );
  INV_X1 U17249 ( .A(n22477), .ZN(n22458) );
  AOI22_X1 U17250 ( .A1(n22785), .A2(n15222), .B1(n22458), .B2(n22784), .ZN(
        n15223) );
  OAI211_X1 U17251 ( .C1(n22478), .C2(n22801), .A(n15224), .B(n15223), .ZN(
        n15225) );
  AOI21_X1 U17252 ( .B1(n22788), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n15225), .ZN(n15226) );
  INV_X1 U17253 ( .A(n15226), .ZN(P1_U3145) );
  NAND2_X1 U17254 ( .A1(n22787), .A2(n22643), .ZN(n15228) );
  AOI22_X1 U17255 ( .A1(n22785), .A2(n22650), .B1(n22784), .B2(n22649), .ZN(
        n15227) );
  OAI211_X1 U17256 ( .C1(n22641), .C2(n22801), .A(n15228), .B(n15227), .ZN(
        n15229) );
  AOI21_X1 U17257 ( .B1(n22788), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n15229), .ZN(n15230) );
  INV_X1 U17258 ( .A(n15230), .ZN(P1_U3150) );
  NAND2_X1 U17259 ( .A1(n22787), .A2(n22580), .ZN(n15233) );
  AOI22_X1 U17260 ( .A1(n22785), .A2(n15231), .B1(n22784), .B2(n22570), .ZN(
        n15232) );
  OAI211_X1 U17261 ( .C1(n22578), .C2(n22801), .A(n15233), .B(n15232), .ZN(
        n15234) );
  AOI21_X1 U17262 ( .B1(n22788), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n15234), .ZN(n15235) );
  INV_X1 U17263 ( .A(n15235), .ZN(P1_U3148) );
  NAND2_X1 U17264 ( .A1(n22787), .A2(n22608), .ZN(n15237) );
  INV_X1 U17265 ( .A(n22605), .ZN(n22614) );
  AOI22_X1 U17266 ( .A1(n22785), .A2(n22615), .B1(n22784), .B2(n22614), .ZN(
        n15236) );
  OAI211_X1 U17267 ( .C1(n22606), .C2(n22801), .A(n15237), .B(n15236), .ZN(
        n15238) );
  AOI21_X1 U17268 ( .B1(n22788), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n15238), .ZN(n15239) );
  INV_X1 U17269 ( .A(n15239), .ZN(P1_U3149) );
  NAND2_X1 U17270 ( .A1(n22787), .A2(n22516), .ZN(n15241) );
  AOI22_X1 U17271 ( .A1(n22785), .A2(n22524), .B1(n22784), .B2(n22523), .ZN(
        n15240) );
  OAI211_X1 U17272 ( .C1(n22514), .C2(n22801), .A(n15241), .B(n15240), .ZN(
        n15242) );
  AOI21_X1 U17273 ( .B1(n22788), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n15242), .ZN(n15243) );
  INV_X1 U17274 ( .A(n15243), .ZN(P1_U3146) );
  NAND2_X1 U17275 ( .A1(n22787), .A2(n22549), .ZN(n15245) );
  AOI22_X1 U17276 ( .A1(n22785), .A2(n22556), .B1(n22784), .B2(n22555), .ZN(
        n15244) );
  OAI211_X1 U17277 ( .C1(n22547), .C2(n22801), .A(n15245), .B(n15244), .ZN(
        n15246) );
  AOI21_X1 U17278 ( .B1(n22788), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n15246), .ZN(n15247) );
  INV_X1 U17279 ( .A(n15247), .ZN(P1_U3147) );
  NAND2_X1 U17280 ( .A1(n22787), .A2(n22674), .ZN(n15250) );
  INV_X1 U17281 ( .A(n22671), .ZN(n22663) );
  AOI22_X1 U17282 ( .A1(n22785), .A2(n15248), .B1(n22784), .B2(n22663), .ZN(
        n15249) );
  OAI211_X1 U17283 ( .C1(n22672), .C2(n22801), .A(n15250), .B(n15249), .ZN(
        n15251) );
  AOI21_X1 U17284 ( .B1(n22788), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n15251), .ZN(n15252) );
  INV_X1 U17285 ( .A(n15252), .ZN(P1_U3151) );
  NOR2_X1 U17286 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15253), .ZN(
        n22744) );
  OAI21_X1 U17287 ( .B1(n15254), .B2(n22746), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15255) );
  AOI21_X1 U17288 ( .B1(n22452), .B2(n11193), .A(n22744), .ZN(n15257) );
  NAND2_X1 U17289 ( .A1(n15255), .A2(n15257), .ZN(n15256) );
  NOR2_X1 U17290 ( .A1(n22474), .A2(n22678), .ZN(n22410) );
  NAND2_X1 U17291 ( .A1(n22747), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n15261) );
  INV_X1 U17292 ( .A(n15257), .ZN(n15258) );
  NAND2_X1 U17293 ( .A1(n15422), .A2(n22404), .ZN(n22483) );
  INV_X1 U17294 ( .A(n22483), .ZN(n22473) );
  AOI22_X1 U17295 ( .A1(n15258), .A2(n22434), .B1(n22473), .B2(n22453), .ZN(
        n22743) );
  INV_X1 U17296 ( .A(n22744), .ZN(n15277) );
  OAI22_X1 U17297 ( .A1(n22743), .A2(n22583), .B1(n22577), .B2(n15277), .ZN(
        n15259) );
  AOI21_X1 U17298 ( .B1(n22746), .B2(n22580), .A(n15259), .ZN(n15260) );
  OAI211_X1 U17299 ( .C1(n22578), .C2(n22755), .A(n15261), .B(n15260), .ZN(
        P1_U3100) );
  NAND2_X1 U17300 ( .A1(n22747), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n15264) );
  OAI22_X1 U17301 ( .A1(n22743), .A2(n22611), .B1(n22605), .B2(n15277), .ZN(
        n15262) );
  AOI21_X1 U17302 ( .B1(n22608), .B2(n22746), .A(n15262), .ZN(n15263) );
  OAI211_X1 U17303 ( .C1(n22606), .C2(n22755), .A(n15264), .B(n15263), .ZN(
        P1_U3101) );
  NAND2_X1 U17304 ( .A1(n22747), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n15267) );
  OAI22_X1 U17305 ( .A1(n22743), .A2(n22646), .B1(n22640), .B2(n15277), .ZN(
        n15265) );
  AOI21_X1 U17306 ( .B1(n22643), .B2(n22746), .A(n15265), .ZN(n15266) );
  OAI211_X1 U17307 ( .C1(n22641), .C2(n22755), .A(n15267), .B(n15266), .ZN(
        P1_U3102) );
  NAND2_X1 U17308 ( .A1(n22747), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n15270) );
  OAI22_X1 U17309 ( .A1(n22743), .A2(n22519), .B1(n22513), .B2(n15277), .ZN(
        n15268) );
  AOI21_X1 U17310 ( .B1(n22516), .B2(n22746), .A(n15268), .ZN(n15269) );
  OAI211_X1 U17311 ( .C1(n22514), .C2(n22755), .A(n15270), .B(n15269), .ZN(
        P1_U3098) );
  NAND2_X1 U17312 ( .A1(n22747), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n15273) );
  OAI22_X1 U17313 ( .A1(n22743), .A2(n22552), .B1(n22546), .B2(n15277), .ZN(
        n15271) );
  AOI21_X1 U17314 ( .B1(n22549), .B2(n22746), .A(n15271), .ZN(n15272) );
  OAI211_X1 U17315 ( .C1(n22547), .C2(n22755), .A(n15273), .B(n15272), .ZN(
        P1_U3099) );
  NAND2_X1 U17316 ( .A1(n22747), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n15276) );
  OAI22_X1 U17317 ( .A1(n22743), .A2(n22490), .B1(n22477), .B2(n15277), .ZN(
        n15274) );
  AOI21_X1 U17318 ( .B1(n22746), .B2(n22487), .A(n15274), .ZN(n15275) );
  OAI211_X1 U17319 ( .C1(n22478), .C2(n22755), .A(n15276), .B(n15275), .ZN(
        P1_U3097) );
  NAND2_X1 U17320 ( .A1(n22747), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n15280) );
  OAI22_X1 U17321 ( .A1(n22743), .A2(n22677), .B1(n22671), .B2(n15277), .ZN(
        n15278) );
  AOI21_X1 U17322 ( .B1(n22746), .B2(n22674), .A(n15278), .ZN(n15279) );
  OAI211_X1 U17323 ( .C1(n22672), .C2(n22755), .A(n15280), .B(n15279), .ZN(
        P1_U3103) );
  XOR2_X1 U17324 ( .A(n14981), .B(n15281), .Z(n22134) );
  INV_X1 U17325 ( .A(n22134), .ZN(n15282) );
  OAI222_X1 U17326 ( .A1(n16054), .A2(n15284), .B1(n16056), .B2(n15283), .C1(
        n16897), .C2(n15282), .ZN(P1_U2898) );
  NAND2_X1 U17327 ( .A1(n15285), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15286) );
  NAND2_X1 U17328 ( .A1(n15287), .A2(n15286), .ZN(n15573) );
  XNOR2_X1 U17329 ( .A(n15573), .B(n17077), .ZN(n15296) );
  NAND2_X1 U17330 ( .A1(n15288), .A2(n15602), .ZN(n15294) );
  NAND2_X1 U17331 ( .A1(n15290), .A2(n15289), .ZN(n15578) );
  INV_X1 U17332 ( .A(n15577), .ZN(n15291) );
  XNOR2_X1 U17333 ( .A(n15578), .B(n15291), .ZN(n15292) );
  NAND2_X1 U17334 ( .A1(n15292), .A2(n15607), .ZN(n15293) );
  NAND2_X1 U17335 ( .A1(n15294), .A2(n15293), .ZN(n15295) );
  OAI21_X1 U17336 ( .B1(n15296), .B2(n15295), .A(n15575), .ZN(n15297) );
  INV_X1 U17337 ( .A(n15297), .ZN(n20737) );
  AOI21_X1 U17338 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21989) );
  INV_X1 U17339 ( .A(n22053), .ZN(n21987) );
  NAND2_X1 U17340 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17078) );
  NOR2_X1 U17341 ( .A1(n15301), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n15299) );
  AOI21_X1 U17342 ( .B1(n21987), .B2(n17078), .A(n22030), .ZN(n15300) );
  INV_X1 U17343 ( .A(n15300), .ZN(n22028) );
  AOI21_X1 U17344 ( .B1(n22056), .B2(n21989), .A(n22028), .ZN(n22013) );
  INV_X1 U17345 ( .A(n15301), .ZN(n15302) );
  NAND2_X1 U17346 ( .A1(n15302), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n15304) );
  OAI22_X1 U17347 ( .A1(n21999), .A2(n21989), .B1(n17078), .B2(n21992), .ZN(
        n15305) );
  NAND2_X1 U17348 ( .A1(n22011), .A2(n15305), .ZN(n22009) );
  AOI21_X1 U17349 ( .B1(n22013), .B2(n22009), .A(n17077), .ZN(n15309) );
  INV_X1 U17350 ( .A(n15305), .ZN(n22033) );
  NOR3_X1 U17351 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n22033), .A3(
        n22011), .ZN(n15306) );
  AOI21_X1 U17352 ( .B1(n22021), .B2(P1_REIP_REG_4__SCAN_IN), .A(n15306), .ZN(
        n15307) );
  OAI21_X1 U17353 ( .B1(n22082), .B2(n22105), .A(n15307), .ZN(n15308) );
  AOI211_X1 U17354 ( .C1(n20737), .C2(n22075), .A(n15309), .B(n15308), .ZN(
        n15310) );
  INV_X1 U17355 ( .A(n15310), .ZN(P1_U3027) );
  OR2_X1 U17356 ( .A1(n15311), .A2(n15312), .ZN(n15352) );
  NAND2_X1 U17357 ( .A1(n15311), .A2(n15312), .ZN(n15313) );
  INV_X1 U17358 ( .A(n22152), .ZN(n15315) );
  INV_X1 U17359 ( .A(n16865), .ZN(n22679) );
  OAI222_X1 U17360 ( .A1(n15315), .A2(n16897), .B1(n16056), .B2(n22679), .C1(
        n15314), .C2(n16054), .ZN(P1_U2897) );
  XNOR2_X1 U17361 ( .A(n15316), .B(n15317), .ZN(n19223) );
  OAI222_X1 U17362 ( .A1(n15324), .A2(n15318), .B1(n17475), .B2(n18183), .C1(
        n20171), .C2(n19223), .ZN(P2_U2904) );
  INV_X1 U17363 ( .A(n16691), .ZN(n15323) );
  INV_X1 U17364 ( .A(n15319), .ZN(n15321) );
  INV_X1 U17365 ( .A(n15316), .ZN(n15320) );
  AOI21_X1 U17366 ( .B1(n15321), .B2(n11231), .A(n15320), .ZN(n19207) );
  INV_X1 U17367 ( .A(n19207), .ZN(n15322) );
  INV_X1 U17368 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n18178) );
  OAI222_X1 U17369 ( .A1(n15324), .A2(n15323), .B1(n15322), .B2(n20171), .C1(
        n17475), .C2(n18178), .ZN(P2_U2905) );
  OAI21_X1 U17370 ( .B1(n15325), .B2(n15327), .A(n15326), .ZN(n15407) );
  INV_X1 U17371 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15779) );
  INV_X1 U17372 ( .A(n15328), .ZN(n15332) );
  NAND2_X1 U17373 ( .A1(n16321), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15329) );
  OAI211_X1 U17374 ( .C1(P1_EBX_REG_5__SCAN_IN), .C2(n11150), .A(n14857), .B(
        n15329), .ZN(n15330) );
  OAI21_X1 U17375 ( .B1(n16297), .B2(P1_EBX_REG_5__SCAN_IN), .A(n15330), .ZN(
        n20722) );
  MUX2_X1 U17376 ( .A(n16297), .B(n16321), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n15334) );
  OR2_X1 U17377 ( .A1(n16323), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15333) );
  AND2_X1 U17378 ( .A1(n15334), .A2(n15333), .ZN(n20715) );
  INV_X1 U17379 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n22012) );
  NAND2_X1 U17380 ( .A1(n14857), .A2(n22012), .ZN(n15336) );
  INV_X1 U17381 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20701) );
  NAND2_X1 U17382 ( .A1(n11192), .A2(n20701), .ZN(n15335) );
  NAND3_X1 U17383 ( .A1(n15336), .A2(n16321), .A3(n15335), .ZN(n15337) );
  OAI21_X1 U17384 ( .B1(P1_EBX_REG_6__SCAN_IN), .B2(n16304), .A(n15337), .ZN(
        n20716) );
  NAND2_X1 U17385 ( .A1(n20715), .A2(n20716), .ZN(n15338) );
  INV_X1 U17386 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n22047) );
  NAND2_X1 U17387 ( .A1(n14857), .A2(n22047), .ZN(n15339) );
  OAI211_X1 U17388 ( .C1(P1_EBX_REG_8__SCAN_IN), .C2(n11150), .A(n15339), .B(
        n16385), .ZN(n15340) );
  OAI21_X1 U17389 ( .B1(P1_EBX_REG_8__SCAN_IN), .B2(n16304), .A(n15340), .ZN(
        n15356) );
  INV_X1 U17390 ( .A(n16297), .ZN(n15544) );
  INV_X1 U17391 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n15960) );
  NAND2_X1 U17392 ( .A1(n15544), .A2(n15960), .ZN(n15343) );
  NAND2_X1 U17393 ( .A1(n16385), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15341) );
  OAI211_X1 U17394 ( .C1(P1_EBX_REG_9__SCAN_IN), .C2(n11150), .A(n14857), .B(
        n15341), .ZN(n15342) );
  NAND2_X1 U17395 ( .A1(n16293), .A2(n15779), .ZN(n15346) );
  INV_X1 U17396 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n22073) );
  NAND2_X1 U17397 ( .A1(n14857), .A2(n22073), .ZN(n15344) );
  OAI211_X1 U17398 ( .C1(P1_EBX_REG_10__SCAN_IN), .C2(n11150), .A(n15344), .B(
        n16385), .ZN(n15345) );
  NAND2_X1 U17399 ( .A1(n15458), .A2(n15349), .ZN(n15350) );
  NAND2_X1 U17400 ( .A1(n17320), .A2(n15350), .ZN(n22068) );
  OAI222_X1 U17401 ( .A1(n15407), .A2(n20698), .B1(n15779), .B2(n20727), .C1(
        n22068), .C2(n16841), .ZN(P1_U2862) );
  OR2_X1 U17402 ( .A1(n15352), .A2(n15351), .ZN(n15453) );
  NAND2_X1 U17403 ( .A1(n15352), .A2(n15351), .ZN(n15353) );
  NAND2_X1 U17404 ( .A1(n15453), .A2(n15353), .ZN(n15612) );
  AOI22_X1 U17405 ( .A1(n16008), .A2(n16862), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n16890), .ZN(n15354) );
  OAI21_X1 U17406 ( .B1(n15612), .B2(n16897), .A(n15354), .ZN(P1_U2896) );
  INV_X1 U17407 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n15613) );
  INV_X1 U17408 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n22136) );
  NAND3_X1 U17409 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .ZN(n22113) );
  NOR2_X1 U17410 ( .A1(n22136), .A2(n22113), .ZN(n15355) );
  NAND4_X1 U17411 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_4__SCAN_IN), .A4(n15355), .ZN(n15360) );
  NOR2_X1 U17412 ( .A1(n15613), .A2(n15360), .ZN(n15455) );
  OAI21_X1 U17413 ( .B1(n15455), .B2(n22245), .A(n22091), .ZN(n15461) );
  NOR2_X1 U17414 ( .A1(n20718), .A2(n15356), .ZN(n15357) );
  OR2_X1 U17415 ( .A1(n15460), .A2(n15357), .ZN(n22038) );
  INV_X1 U17416 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n15373) );
  OAI22_X1 U17417 ( .A1(n22038), .A2(n22276), .B1(n22262), .B2(n15373), .ZN(
        n15358) );
  NAND2_X1 U17418 ( .A1(n22091), .A2(n22810), .ZN(n22193) );
  INV_X1 U17419 ( .A(n22193), .ZN(n22223) );
  AOI211_X1 U17420 ( .C1(n15461), .C2(P1_REIP_REG_8__SCAN_IN), .A(n15358), .B(
        n22223), .ZN(n15365) );
  INV_X1 U17421 ( .A(n15615), .ZN(n15363) );
  OR2_X1 U17422 ( .A1(n22245), .A2(n15455), .ZN(n15359) );
  OAI22_X1 U17423 ( .A1(n15361), .A2(n22213), .B1(n15360), .B2(n15359), .ZN(
        n15362) );
  AOI21_X1 U17424 ( .B1(n22266), .B2(n15363), .A(n15362), .ZN(n15364) );
  OAI211_X1 U17425 ( .C1(n15612), .C2(n22269), .A(n15365), .B(n15364), .ZN(
        P1_U2832) );
  OR2_X1 U17426 ( .A1(n15366), .A2(n15193), .ZN(n15367) );
  AND2_X1 U17427 ( .A1(n11202), .A2(n15367), .ZN(n19168) );
  INV_X1 U17428 ( .A(n19168), .ZN(n17869) );
  OAI211_X1 U17429 ( .C1(n11506), .C2(n15370), .A(n17417), .B(n15446), .ZN(
        n15372) );
  NAND2_X1 U17430 ( .A1(n17423), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n15371) );
  OAI211_X1 U17431 ( .C1(n17869), .C2(n17420), .A(n15372), .B(n15371), .ZN(
        P2_U2877) );
  OAI222_X1 U17432 ( .A1(n15612), .A2(n20698), .B1(n15373), .B2(n20727), .C1(
        n22038), .C2(n16841), .ZN(P1_U2864) );
  NAND2_X1 U17433 ( .A1(n20058), .A2(n15389), .ZN(n15376) );
  INV_X1 U17434 ( .A(n15200), .ZN(n15374) );
  XNOR2_X1 U17435 ( .A(n15375), .B(n15374), .ZN(n15500) );
  AOI21_X1 U17436 ( .B1(n15377), .B2(n15376), .A(n15500), .ZN(n20167) );
  XNOR2_X1 U17437 ( .A(n20167), .B(n20166), .ZN(n15382) );
  INV_X1 U17438 ( .A(n20230), .ZN(n15380) );
  INV_X1 U17439 ( .A(n15500), .ZN(n15378) );
  INV_X1 U17440 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n18156) );
  OAI22_X1 U17441 ( .A1(n17477), .A2(n15378), .B1(n17475), .B2(n18156), .ZN(
        n15379) );
  AOI21_X1 U17442 ( .B1(n20164), .B2(n15380), .A(n15379), .ZN(n15381) );
  OAI21_X1 U17443 ( .B1(n15382), .B2(n20165), .A(n15381), .ZN(P2_U2915) );
  INV_X1 U17444 ( .A(n19110), .ZN(n15518) );
  NAND2_X1 U17445 ( .A1(n19263), .A2(n15383), .ZN(n15384) );
  XNOR2_X1 U17446 ( .A(n15400), .B(n15384), .ZN(n15385) );
  NAND2_X1 U17447 ( .A1(n15385), .A2(n19316), .ZN(n15392) );
  AOI22_X1 U17448 ( .A1(n19323), .A2(n15397), .B1(P2_EBX_REG_3__SCAN_IN), .B2(
        n19328), .ZN(n15388) );
  OAI22_X1 U17449 ( .A1(n15402), .A2(n19237), .B1(n11736), .B2(n19338), .ZN(
        n15386) );
  INV_X1 U17450 ( .A(n15386), .ZN(n15387) );
  OAI211_X1 U17451 ( .C1(n15389), .C2(n19336), .A(n15388), .B(n15387), .ZN(
        n15390) );
  AOI21_X1 U17452 ( .B1(n12303), .B2(n19349), .A(n15390), .ZN(n15391) );
  OAI211_X1 U17453 ( .C1(n15518), .C2(n20058), .A(n15392), .B(n15391), .ZN(
        P2_U2852) );
  INV_X1 U17454 ( .A(n15393), .ZN(n15394) );
  AOI21_X1 U17455 ( .B1(n15396), .B2(n15395), .A(n15394), .ZN(n19421) );
  NAND2_X1 U17456 ( .A1(n19421), .A2(n18095), .ZN(n15406) );
  XNOR2_X1 U17457 ( .A(n15397), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15398) );
  XNOR2_X1 U17458 ( .A(n15399), .B(n15398), .ZN(n19418) );
  INV_X1 U17459 ( .A(n15400), .ZN(n15401) );
  NOR2_X1 U17460 ( .A1(n18112), .A2(n15401), .ZN(n15404) );
  INV_X1 U17461 ( .A(n19407), .ZN(n19258) );
  OAI22_X1 U17462 ( .A1(n15402), .A2(n18076), .B1(n11736), .B2(n19258), .ZN(
        n15403) );
  AOI211_X1 U17463 ( .C1(n18079), .C2(n19418), .A(n15404), .B(n15403), .ZN(
        n15405) );
  OAI211_X1 U17464 ( .C1(n18105), .C2(n12312), .A(n15406), .B(n15405), .ZN(
        P2_U3011) );
  INV_X1 U17465 ( .A(n15407), .ZN(n17073) );
  OAI22_X1 U17466 ( .A1(n22068), .A2(n22276), .B1(n22262), .B2(n15779), .ZN(
        n15408) );
  AOI211_X1 U17467 ( .C1(n22264), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15408), .B(n22223), .ZN(n15412) );
  INV_X1 U17468 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n22067) );
  NAND2_X1 U17469 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n15455), .ZN(n15409) );
  NOR2_X1 U17470 ( .A1(n22067), .A2(n15409), .ZN(n22161) );
  OAI21_X1 U17471 ( .B1(n22161), .B2(n22245), .A(n22091), .ZN(n22164) );
  OAI21_X1 U17472 ( .B1(n22245), .B2(n15409), .A(n22067), .ZN(n15410) );
  NAND2_X1 U17473 ( .A1(n22164), .A2(n15410), .ZN(n15411) );
  OAI211_X1 U17474 ( .C1(n22257), .C2(n17071), .A(n15412), .B(n15411), .ZN(
        n15413) );
  AOI21_X1 U17475 ( .B1(n17073), .B2(n22253), .A(n15413), .ZN(n15414) );
  INV_X1 U17476 ( .A(n15414), .ZN(P1_U2830) );
  INV_X1 U17477 ( .A(n22717), .ZN(n15416) );
  AOI21_X1 U17478 ( .B1(n15416), .B2(n22726), .A(n22305), .ZN(n15417) );
  AOI21_X1 U17479 ( .B1(n22438), .B2(n11193), .A(n15417), .ZN(n15418) );
  NOR2_X1 U17480 ( .A1(n15418), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15420) );
  NOR2_X1 U17481 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15419), .ZN(
        n22715) );
  NAND2_X1 U17482 ( .A1(n22718), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n15426) );
  NOR2_X1 U17483 ( .A1(n22471), .A2(n22468), .ZN(n15423) );
  NOR2_X1 U17484 ( .A1(n15422), .A2(n15421), .ZN(n22393) );
  AOI22_X1 U17485 ( .A1(n22438), .A2(n15423), .B1(n22474), .B2(n22393), .ZN(
        n22714) );
  INV_X1 U17486 ( .A(n22715), .ZN(n15442) );
  OAI22_X1 U17487 ( .A1(n22714), .A2(n22490), .B1(n22477), .B2(n15442), .ZN(
        n15424) );
  AOI21_X1 U17488 ( .B1(n22717), .B2(n22487), .A(n15424), .ZN(n15425) );
  OAI211_X1 U17489 ( .C1(n22478), .C2(n22726), .A(n15426), .B(n15425), .ZN(
        P1_U3065) );
  NAND2_X1 U17490 ( .A1(n22718), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n15429) );
  OAI22_X1 U17491 ( .A1(n22714), .A2(n22519), .B1(n22513), .B2(n15442), .ZN(
        n15427) );
  AOI21_X1 U17492 ( .B1(n22717), .B2(n22516), .A(n15427), .ZN(n15428) );
  OAI211_X1 U17493 ( .C1(n22514), .C2(n22726), .A(n15429), .B(n15428), .ZN(
        P1_U3066) );
  NAND2_X1 U17494 ( .A1(n22718), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n15432) );
  OAI22_X1 U17495 ( .A1(n22714), .A2(n22646), .B1(n22640), .B2(n15442), .ZN(
        n15430) );
  AOI21_X1 U17496 ( .B1(n22717), .B2(n22643), .A(n15430), .ZN(n15431) );
  OAI211_X1 U17497 ( .C1(n22641), .C2(n22726), .A(n15432), .B(n15431), .ZN(
        P1_U3070) );
  NAND2_X1 U17498 ( .A1(n22718), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n15435) );
  OAI22_X1 U17499 ( .A1(n22714), .A2(n22583), .B1(n22577), .B2(n15442), .ZN(
        n15433) );
  AOI21_X1 U17500 ( .B1(n22717), .B2(n22580), .A(n15433), .ZN(n15434) );
  OAI211_X1 U17501 ( .C1(n22578), .C2(n22726), .A(n15435), .B(n15434), .ZN(
        P1_U3068) );
  NAND2_X1 U17502 ( .A1(n22718), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n15438) );
  OAI22_X1 U17503 ( .A1(n22714), .A2(n22552), .B1(n22546), .B2(n15442), .ZN(
        n15436) );
  AOI21_X1 U17504 ( .B1(n22717), .B2(n22549), .A(n15436), .ZN(n15437) );
  OAI211_X1 U17505 ( .C1(n22547), .C2(n22726), .A(n15438), .B(n15437), .ZN(
        P1_U3067) );
  NAND2_X1 U17506 ( .A1(n22718), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n15441) );
  OAI22_X1 U17507 ( .A1(n22714), .A2(n22677), .B1(n22671), .B2(n15442), .ZN(
        n15439) );
  AOI21_X1 U17508 ( .B1(n22717), .B2(n22674), .A(n15439), .ZN(n15440) );
  OAI211_X1 U17509 ( .C1(n22672), .C2(n22726), .A(n15441), .B(n15440), .ZN(
        P1_U3071) );
  NAND2_X1 U17510 ( .A1(n22718), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n15445) );
  OAI22_X1 U17511 ( .A1(n22714), .A2(n22611), .B1(n22605), .B2(n15442), .ZN(
        n15443) );
  AOI21_X1 U17512 ( .B1(n22717), .B2(n22608), .A(n15443), .ZN(n15444) );
  OAI211_X1 U17513 ( .C1(n22606), .C2(n22726), .A(n15445), .B(n15444), .ZN(
        P1_U3069) );
  XNOR2_X1 U17514 ( .A(n15534), .B(n15536), .ZN(n15452) );
  NAND2_X1 U17515 ( .A1(n15489), .A2(n15448), .ZN(n15449) );
  AND2_X1 U17516 ( .A1(n15539), .A2(n15449), .ZN(n19385) );
  INV_X1 U17517 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n15524) );
  NOR2_X1 U17518 ( .A1(n14580), .A2(n15524), .ZN(n15450) );
  AOI21_X1 U17519 ( .B1(n19385), .B2(n14580), .A(n15450), .ZN(n15451) );
  OAI21_X1 U17520 ( .B1(n15452), .B2(n17428), .A(n15451), .ZN(P2_U2875) );
  AOI21_X1 U17521 ( .B1(n15454), .B2(n15453), .A(n15325), .ZN(n16096) );
  INV_X1 U17522 ( .A(n16096), .ZN(n15493) );
  INV_X1 U17523 ( .A(n22245), .ZN(n22235) );
  INV_X1 U17524 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n22059) );
  NAND3_X1 U17525 ( .A1(n22235), .A2(n15455), .A3(n22059), .ZN(n15456) );
  OAI211_X1 U17526 ( .C1(n22213), .C2(n15457), .A(n22193), .B(n15456), .ZN(
        n15465) );
  OAI21_X1 U17527 ( .B1(n15460), .B2(n15459), .A(n15458), .ZN(n22060) );
  NAND2_X1 U17528 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n15461), .ZN(n15463) );
  NAND2_X1 U17529 ( .A1(n22236), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n15462) );
  OAI211_X1 U17530 ( .C1(n22060), .C2(n22276), .A(n15463), .B(n15462), .ZN(
        n15464) );
  AOI211_X1 U17531 ( .C1(n22266), .C2(n15466), .A(n15465), .B(n15464), .ZN(
        n15467) );
  OAI21_X1 U17532 ( .B1(n15493), .B2(n22269), .A(n15467), .ZN(P1_U2831) );
  AOI22_X1 U17533 ( .A1(n16008), .A2(n16858), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n16890), .ZN(n15468) );
  OAI21_X1 U17534 ( .B1(n15493), .B2(n16897), .A(n15468), .ZN(P1_U2895) );
  XNOR2_X1 U17535 ( .A(n15469), .B(n16076), .ZN(n18042) );
  INV_X1 U17536 ( .A(n18042), .ZN(n15485) );
  NAND2_X1 U17537 ( .A1(n15471), .A2(n15470), .ZN(n15472) );
  AND2_X1 U17538 ( .A1(n15473), .A2(n15472), .ZN(n18041) );
  NOR2_X1 U17539 ( .A1(n18045), .A2(n19416), .ZN(n15483) );
  NAND3_X1 U17540 ( .A1(n19411), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n19410), .ZN(n16074) );
  INV_X1 U17541 ( .A(n17923), .ZN(n17786) );
  NAND2_X1 U17542 ( .A1(n17786), .A2(n15474), .ZN(n15475) );
  NAND2_X1 U17543 ( .A1(n15476), .A2(n15475), .ZN(n15478) );
  NOR2_X1 U17544 ( .A1(n15478), .A2(n15477), .ZN(n19412) );
  OAI21_X1 U17545 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17791), .A(
        n19412), .ZN(n16078) );
  NOR2_X1 U17546 ( .A1(n11748), .A2(n19258), .ZN(n15479) );
  AOI21_X1 U17547 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n16078), .A(
        n15479), .ZN(n15481) );
  NAND2_X1 U17548 ( .A1(n19408), .A2(n15500), .ZN(n15480) );
  OAI211_X1 U17549 ( .C1(n16074), .C2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n15481), .B(n15480), .ZN(n15482) );
  AOI211_X1 U17550 ( .C1(n18041), .C2(n19419), .A(n15483), .B(n15482), .ZN(
        n15484) );
  OAI21_X1 U17551 ( .B1(n15485), .B2(n19375), .A(n15484), .ZN(P2_U3042) );
  INV_X1 U17552 ( .A(n15446), .ZN(n15488) );
  INV_X1 U17553 ( .A(n15534), .ZN(n15487) );
  OAI211_X1 U17554 ( .C1(n15488), .C2(n11508), .A(n15487), .B(n17417), .ZN(
        n15492) );
  AOI21_X1 U17555 ( .B1(n15490), .B2(n11202), .A(n15447), .ZN(n19173) );
  NAND2_X1 U17556 ( .A1(n14580), .A2(n19173), .ZN(n15491) );
  OAI211_X1 U17557 ( .C1(n14580), .C2(n12199), .A(n15492), .B(n15491), .ZN(
        P2_U2876) );
  OAI222_X1 U17558 ( .A1(n15493), .A2(n20698), .B1(n15960), .B2(n20727), .C1(
        n22060), .C2(n16841), .ZN(P1_U2863) );
  INV_X1 U17559 ( .A(n18039), .ZN(n15497) );
  NOR2_X1 U17560 ( .A1(n11181), .A2(n15494), .ZN(n15496) );
  AOI21_X1 U17561 ( .B1(n15497), .B2(n15496), .A(n19432), .ZN(n15495) );
  OAI21_X1 U17562 ( .B1(n15497), .B2(n15496), .A(n15495), .ZN(n15506) );
  INV_X1 U17563 ( .A(n18045), .ZN(n15504) );
  AOI22_X1 U17564 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19346), .B1(
        P2_EBX_REG_4__SCAN_IN), .B2(n19328), .ZN(n15498) );
  OAI211_X1 U17565 ( .C1(n19338), .C2(n11748), .A(n15498), .B(n19380), .ZN(
        n15499) );
  AOI21_X1 U17566 ( .B1(n19348), .B2(n15500), .A(n15499), .ZN(n15501) );
  OAI21_X1 U17567 ( .B1(n15502), .B2(n19342), .A(n15501), .ZN(n15503) );
  AOI21_X1 U17568 ( .B1(n15504), .B2(n19349), .A(n15503), .ZN(n15505) );
  OAI211_X1 U17569 ( .C1(n20166), .C2(n15518), .A(n15506), .B(n15505), .ZN(
        P2_U2851) );
  NOR2_X1 U17570 ( .A1(n11181), .A2(n16058), .ZN(n15507) );
  XNOR2_X1 U17571 ( .A(n15507), .B(n18031), .ZN(n15508) );
  NAND2_X1 U17572 ( .A1(n15508), .A2(n19316), .ZN(n15517) );
  AOI22_X1 U17573 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19346), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n19307), .ZN(n15509) );
  INV_X1 U17574 ( .A(n15509), .ZN(n15515) );
  AND2_X1 U17575 ( .A1(n18033), .A2(n19349), .ZN(n15514) );
  NAND2_X1 U17576 ( .A1(n18120), .A2(n19348), .ZN(n15511) );
  NAND2_X1 U17577 ( .A1(n19328), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n15510) );
  OAI211_X1 U17578 ( .C1(n19342), .C2(n15512), .A(n15511), .B(n15510), .ZN(
        n15513) );
  NOR3_X1 U17579 ( .A1(n15515), .A2(n15514), .A3(n15513), .ZN(n15516) );
  OAI211_X1 U17580 ( .C1(n15518), .C2(n16017), .A(n15517), .B(n15516), .ZN(
        P2_U2853) );
  NOR2_X1 U17581 ( .A1(n11181), .A2(n15519), .ZN(n19182) );
  XNOR2_X1 U17582 ( .A(n19182), .B(n18101), .ZN(n15520) );
  NAND2_X1 U17583 ( .A1(n15520), .A2(n19316), .ZN(n15527) );
  INV_X1 U17584 ( .A(n19328), .ZN(n19188) );
  OAI21_X1 U17585 ( .B1(n11776), .B2(n19338), .A(n19258), .ZN(n15521) );
  AOI21_X1 U17586 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19346), .A(
        n15521), .ZN(n15523) );
  NAND2_X1 U17587 ( .A1(n19348), .A2(n19383), .ZN(n15522) );
  OAI211_X1 U17588 ( .C1(n19188), .C2(n15524), .A(n15523), .B(n15522), .ZN(
        n15525) );
  AOI21_X1 U17589 ( .B1(n19385), .B2(n19349), .A(n15525), .ZN(n15526) );
  OAI211_X1 U17590 ( .C1(n19342), .C2(n15528), .A(n15527), .B(n15526), .ZN(
        P2_U2843) );
  OAI21_X1 U17591 ( .B1(n15529), .B2(n15531), .A(n15530), .ZN(n17039) );
  AOI22_X1 U17592 ( .A1(n16008), .A2(n16843), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n16890), .ZN(n15532) );
  OAI21_X1 U17593 ( .B1(n17039), .B2(n16897), .A(n15532), .ZN(P1_U2890) );
  AND2_X1 U17594 ( .A1(n15536), .A2(n15535), .ZN(n15533) );
  AOI21_X1 U17595 ( .B1(n15534), .B2(n15536), .A(n15535), .ZN(n15537) );
  OR3_X1 U17596 ( .A1(n16115), .A2(n15537), .A3(n17428), .ZN(n15542) );
  AND2_X1 U17597 ( .A1(n15539), .A2(n15538), .ZN(n15540) );
  OR2_X1 U17598 ( .A1(n15540), .A2(n15569), .ZN(n17617) );
  INV_X1 U17599 ( .A(n17617), .ZN(n19195) );
  NAND2_X1 U17600 ( .A1(n19195), .A2(n14580), .ZN(n15541) );
  OAI211_X1 U17601 ( .C1(n14580), .C2(n12200), .A(n15542), .B(n15541), .ZN(
        P2_U2874) );
  INV_X1 U17602 ( .A(n17034), .ZN(n15561) );
  NAND2_X1 U17603 ( .A1(n22264), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15559) );
  MUX2_X1 U17604 ( .A(n16297), .B(n16321), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n15543) );
  OAI21_X1 U17605 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16323), .A(
        n15543), .ZN(n17319) );
  INV_X1 U17606 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15774) );
  NAND2_X1 U17607 ( .A1(n15544), .A2(n15774), .ZN(n15547) );
  NAND2_X1 U17608 ( .A1(n16385), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15545) );
  OAI211_X1 U17609 ( .C1(P1_EBX_REG_13__SCAN_IN), .C2(n11150), .A(n14857), .B(
        n15545), .ZN(n15546) );
  AND2_X1 U17610 ( .A1(n15547), .A2(n15546), .ZN(n16003) );
  NAND2_X1 U17611 ( .A1(n16385), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15548) );
  NAND2_X1 U17612 ( .A1(n14857), .A2(n15548), .ZN(n15550) );
  INV_X1 U17613 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n22171) );
  NAND2_X1 U17614 ( .A1(n11192), .A2(n22171), .ZN(n15549) );
  NAND2_X1 U17615 ( .A1(n15550), .A2(n15549), .ZN(n15551) );
  OAI21_X1 U17616 ( .B1(n16304), .B2(P1_EBX_REG_12__SCAN_IN), .A(n15551), .ZN(
        n17299) );
  NAND2_X1 U17617 ( .A1(n16003), .A2(n17299), .ZN(n15552) );
  INV_X1 U17618 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16348) );
  NAND2_X1 U17619 ( .A1(n14857), .A2(n16348), .ZN(n15553) );
  OAI211_X1 U17620 ( .C1(P1_EBX_REG_14__SCAN_IN), .C2(n11150), .A(n15553), .B(
        n16385), .ZN(n15554) );
  OAI21_X1 U17621 ( .B1(P1_EBX_REG_14__SCAN_IN), .B2(n16304), .A(n15554), .ZN(
        n15555) );
  OR2_X1 U17622 ( .A1(n16005), .A2(n15555), .ZN(n15556) );
  NAND2_X1 U17623 ( .A1(n16155), .A2(n15556), .ZN(n21980) );
  INV_X1 U17624 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15626) );
  OAI22_X1 U17625 ( .A1(n21980), .A2(n22276), .B1(n22262), .B2(n15626), .ZN(
        n15557) );
  INV_X1 U17626 ( .A(n15557), .ZN(n15558) );
  NAND3_X1 U17627 ( .A1(n15559), .A2(n15558), .A3(n22193), .ZN(n15560) );
  AOI21_X1 U17628 ( .B1(n22266), .B2(n15561), .A(n15560), .ZN(n15566) );
  INV_X1 U17629 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20651) );
  INV_X1 U17630 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n22177) );
  NAND2_X1 U17631 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n22161), .ZN(n22170) );
  NOR3_X1 U17632 ( .A1(n22177), .A2(n22245), .A3(n22170), .ZN(n16014) );
  NAND2_X1 U17633 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n16014), .ZN(n15562) );
  NOR2_X1 U17634 ( .A1(n20651), .A2(n15562), .ZN(n22182) );
  INV_X1 U17635 ( .A(n22182), .ZN(n15564) );
  OAI21_X1 U17636 ( .B1(n22200), .B2(n20651), .A(n15562), .ZN(n15563) );
  NAND2_X1 U17637 ( .A1(n15564), .A2(n15563), .ZN(n15565) );
  OAI211_X1 U17638 ( .C1(n17039), .C2(n22269), .A(n15566), .B(n15565), .ZN(
        P1_U2826) );
  OR2_X1 U17639 ( .A1(n15569), .A2(n15568), .ZN(n15570) );
  NAND2_X1 U17640 ( .A1(n15567), .A2(n15570), .ZN(n19206) );
  NAND2_X1 U17641 ( .A1(n16115), .A2(n16112), .ZN(n16046) );
  OAI211_X1 U17642 ( .C1(n16115), .C2(n16112), .A(n16046), .B(n17417), .ZN(
        n15572) );
  NAND2_X1 U17643 ( .A1(n17423), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15571) );
  OAI211_X1 U17644 ( .C1(n19206), .C2(n17420), .A(n15572), .B(n15571), .ZN(
        P2_U2873) );
  NAND2_X1 U17645 ( .A1(n15573), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n15574) );
  NAND2_X1 U17646 ( .A1(n15576), .A2(n15602), .ZN(n15581) );
  OR2_X1 U17647 ( .A1(n15578), .A2(n15577), .ZN(n15586) );
  XNOR2_X1 U17648 ( .A(n15586), .B(n15587), .ZN(n15579) );
  NAND2_X1 U17649 ( .A1(n15579), .A2(n15607), .ZN(n15580) );
  NAND2_X1 U17650 ( .A1(n15581), .A2(n15580), .ZN(n15582) );
  INV_X1 U17651 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n22020) );
  XNOR2_X1 U17652 ( .A(n15582), .B(n22020), .ZN(n20741) );
  NAND2_X1 U17653 ( .A1(n15582), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15583) );
  INV_X1 U17654 ( .A(n15586), .ZN(n15588) );
  NAND2_X1 U17655 ( .A1(n15588), .A2(n15587), .ZN(n15594) );
  INV_X1 U17656 ( .A(n15589), .ZN(n15595) );
  XNOR2_X1 U17657 ( .A(n15594), .B(n15595), .ZN(n15590) );
  NAND2_X1 U17658 ( .A1(n15590), .A2(n15607), .ZN(n15591) );
  NAND2_X1 U17659 ( .A1(n15593), .A2(n15602), .ZN(n15599) );
  INV_X1 U17660 ( .A(n15594), .ZN(n15596) );
  NAND2_X1 U17661 ( .A1(n15596), .A2(n15595), .ZN(n15605) );
  XNOR2_X1 U17662 ( .A(n15605), .B(n15606), .ZN(n15597) );
  NAND2_X1 U17663 ( .A1(n15597), .A2(n15607), .ZN(n15598) );
  NAND2_X1 U17664 ( .A1(n15599), .A2(n15598), .ZN(n15600) );
  INV_X1 U17665 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n22037) );
  XNOR2_X1 U17666 ( .A(n15600), .B(n22037), .ZN(n20753) );
  NAND2_X1 U17667 ( .A1(n15600), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15601) );
  NAND2_X1 U17668 ( .A1(n20752), .A2(n15601), .ZN(n15611) );
  NOR2_X1 U17669 ( .A1(n15603), .A2(n14938), .ZN(n15604) );
  INV_X1 U17670 ( .A(n15605), .ZN(n15608) );
  NAND3_X1 U17671 ( .A1(n15608), .A2(n15607), .A3(n15606), .ZN(n15609) );
  NAND2_X1 U17672 ( .A1(n17256), .A2(n15609), .ZN(n16088) );
  XNOR2_X1 U17673 ( .A(n16088), .B(n22047), .ZN(n15610) );
  NAND2_X1 U17674 ( .A1(n15611), .A2(n15610), .ZN(n16090) );
  OAI21_X1 U17675 ( .B1(n11168), .B2(n15610), .A(n16090), .ZN(n22039) );
  INV_X1 U17676 ( .A(n15612), .ZN(n15617) );
  NOR2_X1 U17677 ( .A1(n22066), .A2(n15613), .ZN(n22041) );
  AOI21_X1 U17678 ( .B1(n20760), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n22041), .ZN(n15614) );
  OAI21_X1 U17679 ( .B1(n15615), .B2(n20759), .A(n15614), .ZN(n15616) );
  AOI21_X1 U17680 ( .B1(n15617), .B2(n20762), .A(n15616), .ZN(n15618) );
  OAI21_X1 U17681 ( .B1(n22039), .B2(n22277), .A(n15618), .ZN(P1_U2991) );
  NAND2_X1 U17682 ( .A1(n15326), .A2(n15620), .ZN(n15621) );
  NAND2_X1 U17683 ( .A1(n15619), .A2(n15621), .ZN(n16039) );
  OAI21_X1 U17684 ( .B1(n16039), .B2(n16040), .A(n15619), .ZN(n15623) );
  NAND2_X1 U17685 ( .A1(n15623), .A2(n15622), .ZN(n16002) );
  OR2_X1 U17686 ( .A1(n15623), .A2(n15622), .ZN(n15624) );
  AOI22_X1 U17687 ( .A1(n16008), .A2(n16267), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n16890), .ZN(n15625) );
  OAI21_X1 U17688 ( .B1(n17059), .B2(n16897), .A(n15625), .ZN(P1_U2892) );
  OAI222_X1 U17689 ( .A1(n17039), .A2(n20698), .B1(n15626), .B2(n20727), .C1(
        n21980), .C2(n16841), .ZN(P1_U2858) );
  XOR2_X1 U17690 ( .A(DATAI_30_), .B(keyinput_130), .Z(n15630) );
  XNOR2_X1 U17691 ( .A(keyinput_128), .B(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(
        n15629) );
  XNOR2_X1 U17692 ( .A(DATAI_29_), .B(keyinput_131), .ZN(n15628) );
  XNOR2_X1 U17693 ( .A(DATAI_31_), .B(keyinput_129), .ZN(n15627) );
  NOR4_X1 U17694 ( .A1(n15630), .A2(n15629), .A3(n15628), .A4(n15627), .ZN(
        n15633) );
  XNOR2_X1 U17695 ( .A(DATAI_28_), .B(keyinput_132), .ZN(n15632) );
  XOR2_X1 U17696 ( .A(DATAI_27_), .B(keyinput_133), .Z(n15631) );
  OAI21_X1 U17697 ( .B1(n15633), .B2(n15632), .A(n15631), .ZN(n15636) );
  XOR2_X1 U17698 ( .A(DATAI_25_), .B(keyinput_135), .Z(n15635) );
  XOR2_X1 U17699 ( .A(DATAI_26_), .B(keyinput_134), .Z(n15634) );
  NAND3_X1 U17700 ( .A1(n15636), .A2(n15635), .A3(n15634), .ZN(n15639) );
  XOR2_X1 U17701 ( .A(DATAI_24_), .B(keyinput_136), .Z(n15638) );
  XOR2_X1 U17702 ( .A(DATAI_23_), .B(keyinput_137), .Z(n15637) );
  NAND3_X1 U17703 ( .A1(n15639), .A2(n15638), .A3(n15637), .ZN(n15643) );
  XNOR2_X1 U17704 ( .A(DATAI_22_), .B(keyinput_138), .ZN(n15642) );
  XOR2_X1 U17705 ( .A(DATAI_20_), .B(keyinput_140), .Z(n15641) );
  XOR2_X1 U17706 ( .A(DATAI_21_), .B(keyinput_139), .Z(n15640) );
  AOI211_X1 U17707 ( .C1(n15643), .C2(n15642), .A(n15641), .B(n15640), .ZN(
        n15646) );
  XOR2_X1 U17708 ( .A(DATAI_19_), .B(keyinput_141), .Z(n15645) );
  XOR2_X1 U17709 ( .A(DATAI_18_), .B(keyinput_142), .Z(n15644) );
  NOR3_X1 U17710 ( .A1(n15646), .A2(n15645), .A3(n15644), .ZN(n15649) );
  XOR2_X1 U17711 ( .A(DATAI_17_), .B(keyinput_143), .Z(n15648) );
  XNOR2_X1 U17712 ( .A(DATAI_16_), .B(keyinput_144), .ZN(n15647) );
  NOR3_X1 U17713 ( .A1(n15649), .A2(n15648), .A3(n15647), .ZN(n15653) );
  XOR2_X1 U17714 ( .A(DATAI_14_), .B(keyinput_146), .Z(n15652) );
  XNOR2_X1 U17715 ( .A(DATAI_13_), .B(keyinput_147), .ZN(n15651) );
  XNOR2_X1 U17716 ( .A(DATAI_15_), .B(keyinput_145), .ZN(n15650) );
  NOR4_X1 U17717 ( .A1(n15653), .A2(n15652), .A3(n15651), .A4(n15650), .ZN(
        n15657) );
  XOR2_X1 U17718 ( .A(DATAI_12_), .B(keyinput_148), .Z(n15656) );
  XOR2_X1 U17719 ( .A(DATAI_11_), .B(keyinput_149), .Z(n15655) );
  XNOR2_X1 U17720 ( .A(DATAI_10_), .B(keyinput_150), .ZN(n15654) );
  NOR4_X1 U17721 ( .A1(n15657), .A2(n15656), .A3(n15655), .A4(n15654), .ZN(
        n15670) );
  XOR2_X1 U17722 ( .A(DATAI_7_), .B(keyinput_153), .Z(n15661) );
  XOR2_X1 U17723 ( .A(DATAI_9_), .B(keyinput_151), .Z(n15660) );
  XOR2_X1 U17724 ( .A(DATAI_8_), .B(keyinput_152), .Z(n15659) );
  XOR2_X1 U17725 ( .A(DATAI_6_), .B(keyinput_154), .Z(n15658) );
  NAND4_X1 U17726 ( .A1(n15661), .A2(n15660), .A3(n15659), .A4(n15658), .ZN(
        n15669) );
  XOR2_X1 U17727 ( .A(DATAI_5_), .B(keyinput_155), .Z(n15667) );
  XOR2_X1 U17728 ( .A(DATAI_3_), .B(keyinput_157), .Z(n15666) );
  XNOR2_X1 U17729 ( .A(DATAI_1_), .B(keyinput_159), .ZN(n15664) );
  XNOR2_X1 U17730 ( .A(DATAI_4_), .B(keyinput_156), .ZN(n15663) );
  XNOR2_X1 U17731 ( .A(DATAI_2_), .B(keyinput_158), .ZN(n15662) );
  NAND3_X1 U17732 ( .A1(n15664), .A2(n15663), .A3(n15662), .ZN(n15665) );
  NOR3_X1 U17733 ( .A1(n15667), .A2(n15666), .A3(n15665), .ZN(n15668) );
  OAI21_X1 U17734 ( .B1(n15670), .B2(n15669), .A(n15668), .ZN(n15677) );
  INV_X1 U17735 ( .A(keyinput_162), .ZN(n15671) );
  XNOR2_X1 U17736 ( .A(n15671), .B(NA), .ZN(n15676) );
  INV_X1 U17737 ( .A(DATAI_0_), .ZN(n15673) );
  OAI22_X1 U17738 ( .A1(n15673), .A2(keyinput_160), .B1(keyinput_161), .B2(
        HOLD), .ZN(n15672) );
  AOI21_X1 U17739 ( .B1(n15673), .B2(keyinput_160), .A(n15672), .ZN(n15675) );
  NAND2_X1 U17740 ( .A1(HOLD), .A2(keyinput_161), .ZN(n15674) );
  NAND4_X1 U17741 ( .A1(n15677), .A2(n15676), .A3(n15675), .A4(n15674), .ZN(
        n15680) );
  INV_X1 U17742 ( .A(BS16), .ZN(n17944) );
  XNOR2_X1 U17743 ( .A(n17944), .B(keyinput_163), .ZN(n15679) );
  XNOR2_X1 U17744 ( .A(READY1), .B(keyinput_164), .ZN(n15678) );
  AOI21_X1 U17745 ( .B1(n15680), .B2(n15679), .A(n15678), .ZN(n15683) );
  XNOR2_X1 U17746 ( .A(keyinput_165), .B(READY2), .ZN(n15682) );
  XNOR2_X1 U17747 ( .A(keyinput_166), .B(P1_READREQUEST_REG_SCAN_IN), .ZN(
        n15681) );
  NOR3_X1 U17748 ( .A1(n15683), .A2(n15682), .A3(n15681), .ZN(n15690) );
  INV_X1 U17749 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n18025) );
  XNOR2_X1 U17750 ( .A(n18025), .B(keyinput_167), .ZN(n15686) );
  XOR2_X1 U17751 ( .A(keyinput_168), .B(P1_CODEFETCH_REG_SCAN_IN), .Z(n15685)
         );
  INV_X1 U17752 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n22804) );
  XNOR2_X1 U17753 ( .A(n22804), .B(keyinput_169), .ZN(n15684) );
  NAND3_X1 U17754 ( .A1(n15686), .A2(n15685), .A3(n15684), .ZN(n15689) );
  XOR2_X1 U17755 ( .A(keyinput_170), .B(P1_D_C_N_REG_SCAN_IN), .Z(n15688) );
  XNOR2_X1 U17756 ( .A(keyinput_171), .B(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15687) );
  OAI211_X1 U17757 ( .C1(n15690), .C2(n15689), .A(n15688), .B(n15687), .ZN(
        n15693) );
  XNOR2_X1 U17758 ( .A(n22305), .B(keyinput_172), .ZN(n15692) );
  INV_X1 U17759 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n17987) );
  XNOR2_X1 U17760 ( .A(n17987), .B(keyinput_173), .ZN(n15691) );
  AOI21_X1 U17761 ( .B1(n15693), .B2(n15692), .A(n15691), .ZN(n15700) );
  XOR2_X1 U17762 ( .A(keyinput_176), .B(P1_BYTEENABLE_REG_0__SCAN_IN), .Z(
        n15697) );
  XOR2_X1 U17763 ( .A(keyinput_174), .B(P1_FLUSH_REG_SCAN_IN), .Z(n15696) );
  XNOR2_X1 U17764 ( .A(keyinput_175), .B(P1_W_R_N_REG_SCAN_IN), .ZN(n15695) );
  XNOR2_X1 U17765 ( .A(keyinput_177), .B(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(
        n15694) );
  NAND4_X1 U17766 ( .A1(n15697), .A2(n15696), .A3(n15695), .A4(n15694), .ZN(
        n15699) );
  XNOR2_X1 U17767 ( .A(keyinput_178), .B(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(
        n15698) );
  OAI21_X1 U17768 ( .B1(n15700), .B2(n15699), .A(n15698), .ZN(n15707) );
  XOR2_X1 U17769 ( .A(P1_REIP_REG_29__SCAN_IN), .B(keyinput_182), .Z(n15704)
         );
  XNOR2_X1 U17770 ( .A(P1_REIP_REG_30__SCAN_IN), .B(keyinput_181), .ZN(n15703)
         );
  XNOR2_X1 U17771 ( .A(keyinput_179), .B(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(
        n15702) );
  XNOR2_X1 U17772 ( .A(P1_REIP_REG_31__SCAN_IN), .B(keyinput_180), .ZN(n15701)
         );
  NOR4_X1 U17773 ( .A1(n15704), .A2(n15703), .A3(n15702), .A4(n15701), .ZN(
        n15706) );
  XNOR2_X1 U17774 ( .A(P1_REIP_REG_28__SCAN_IN), .B(keyinput_183), .ZN(n15705)
         );
  AOI21_X1 U17775 ( .B1(n15707), .B2(n15706), .A(n15705), .ZN(n15710) );
  XNOR2_X1 U17776 ( .A(P1_REIP_REG_27__SCAN_IN), .B(keyinput_184), .ZN(n15709)
         );
  XOR2_X1 U17777 ( .A(P1_REIP_REG_26__SCAN_IN), .B(keyinput_185), .Z(n15708)
         );
  OAI21_X1 U17778 ( .B1(n15710), .B2(n15709), .A(n15708), .ZN(n15713) );
  XOR2_X1 U17779 ( .A(P1_REIP_REG_24__SCAN_IN), .B(keyinput_187), .Z(n15712)
         );
  XOR2_X1 U17780 ( .A(P1_REIP_REG_25__SCAN_IN), .B(keyinput_186), .Z(n15711)
         );
  NAND3_X1 U17781 ( .A1(n15713), .A2(n15712), .A3(n15711), .ZN(n15716) );
  XOR2_X1 U17782 ( .A(P1_REIP_REG_23__SCAN_IN), .B(keyinput_188), .Z(n15715)
         );
  XNOR2_X1 U17783 ( .A(P1_REIP_REG_22__SCAN_IN), .B(keyinput_189), .ZN(n15714)
         );
  AOI21_X1 U17784 ( .B1(n15716), .B2(n15715), .A(n15714), .ZN(n15722) );
  XNOR2_X1 U17785 ( .A(P1_REIP_REG_21__SCAN_IN), .B(keyinput_190), .ZN(n15721)
         );
  XOR2_X1 U17786 ( .A(P1_REIP_REG_19__SCAN_IN), .B(keyinput_192), .Z(n15719)
         );
  XNOR2_X1 U17787 ( .A(P1_REIP_REG_18__SCAN_IN), .B(keyinput_193), .ZN(n15718)
         );
  XNOR2_X1 U17788 ( .A(P1_REIP_REG_20__SCAN_IN), .B(keyinput_191), .ZN(n15717)
         );
  NOR3_X1 U17789 ( .A1(n15719), .A2(n15718), .A3(n15717), .ZN(n15720) );
  OAI21_X1 U17790 ( .B1(n15722), .B2(n15721), .A(n15720), .ZN(n15726) );
  XNOR2_X1 U17791 ( .A(P1_REIP_REG_17__SCAN_IN), .B(keyinput_194), .ZN(n15725)
         );
  XOR2_X1 U17792 ( .A(P1_REIP_REG_16__SCAN_IN), .B(keyinput_195), .Z(n15724)
         );
  XNOR2_X1 U17793 ( .A(P1_REIP_REG_15__SCAN_IN), .B(keyinput_196), .ZN(n15723)
         );
  AOI211_X1 U17794 ( .C1(n15726), .C2(n15725), .A(n15724), .B(n15723), .ZN(
        n15733) );
  XNOR2_X1 U17795 ( .A(P1_REIP_REG_14__SCAN_IN), .B(keyinput_197), .ZN(n15732)
         );
  XNOR2_X1 U17796 ( .A(P1_REIP_REG_11__SCAN_IN), .B(keyinput_200), .ZN(n15731)
         );
  XOR2_X1 U17797 ( .A(P1_REIP_REG_10__SCAN_IN), .B(keyinput_201), .Z(n15729)
         );
  XNOR2_X1 U17798 ( .A(P1_REIP_REG_13__SCAN_IN), .B(keyinput_198), .ZN(n15728)
         );
  XNOR2_X1 U17799 ( .A(P1_REIP_REG_12__SCAN_IN), .B(keyinput_199), .ZN(n15727)
         );
  NAND3_X1 U17800 ( .A1(n15729), .A2(n15728), .A3(n15727), .ZN(n15730) );
  NOR4_X1 U17801 ( .A1(n15733), .A2(n15732), .A3(n15731), .A4(n15730), .ZN(
        n15738) );
  XNOR2_X1 U17802 ( .A(P1_REIP_REG_9__SCAN_IN), .B(keyinput_202), .ZN(n15737)
         );
  XOR2_X1 U17803 ( .A(keyinput_206), .B(P1_REIP_REG_5__SCAN_IN), .Z(n15735) );
  XNOR2_X1 U17804 ( .A(keyinput_205), .B(P1_REIP_REG_6__SCAN_IN), .ZN(n15734)
         );
  NOR2_X1 U17805 ( .A1(n15735), .A2(n15734), .ZN(n15742) );
  XNOR2_X1 U17806 ( .A(P1_REIP_REG_8__SCAN_IN), .B(keyinput_203), .ZN(n15736)
         );
  OAI211_X1 U17807 ( .C1(n15738), .C2(n15737), .A(n15742), .B(n15736), .ZN(
        n15746) );
  XNOR2_X1 U17808 ( .A(keyinput_204), .B(P1_REIP_REG_7__SCAN_IN), .ZN(n15741)
         );
  XNOR2_X1 U17809 ( .A(keyinput_207), .B(P1_REIP_REG_4__SCAN_IN), .ZN(n15740)
         );
  XOR2_X1 U17810 ( .A(keyinput_208), .B(P1_REIP_REG_3__SCAN_IN), .Z(n15739) );
  AOI211_X1 U17811 ( .C1(n15742), .C2(n15741), .A(n15740), .B(n15739), .ZN(
        n15745) );
  XOR2_X1 U17812 ( .A(keyinput_210), .B(P1_REIP_REG_1__SCAN_IN), .Z(n15744) );
  XNOR2_X1 U17813 ( .A(keyinput_209), .B(P1_REIP_REG_2__SCAN_IN), .ZN(n15743)
         );
  AOI211_X1 U17814 ( .C1(n15746), .C2(n15745), .A(n15744), .B(n15743), .ZN(
        n15749) );
  XNOR2_X1 U17815 ( .A(keyinput_211), .B(P1_REIP_REG_0__SCAN_IN), .ZN(n15748)
         );
  XNOR2_X1 U17816 ( .A(P1_EBX_REG_31__SCAN_IN), .B(keyinput_212), .ZN(n15747)
         );
  NOR3_X1 U17817 ( .A1(n15749), .A2(n15748), .A3(n15747), .ZN(n15752) );
  XOR2_X1 U17818 ( .A(P1_EBX_REG_30__SCAN_IN), .B(keyinput_213), .Z(n15751) );
  INV_X1 U17819 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n16815) );
  XNOR2_X1 U17820 ( .A(n16815), .B(keyinput_214), .ZN(n15750) );
  OAI21_X1 U17821 ( .B1(n15752), .B2(n15751), .A(n15750), .ZN(n15757) );
  XOR2_X1 U17822 ( .A(P1_EBX_REG_28__SCAN_IN), .B(keyinput_215), .Z(n15756) );
  INV_X1 U17823 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n16817) );
  OAI22_X1 U17824 ( .A1(n16817), .A2(keyinput_216), .B1(P1_EBX_REG_26__SCAN_IN), .B2(keyinput_217), .ZN(n15753) );
  AOI21_X1 U17825 ( .B1(n16817), .B2(keyinput_216), .A(n15753), .ZN(n15755) );
  NAND2_X1 U17826 ( .A1(P1_EBX_REG_26__SCAN_IN), .A2(keyinput_217), .ZN(n15754) );
  NAND4_X1 U17827 ( .A1(n15757), .A2(n15756), .A3(n15755), .A4(n15754), .ZN(
        n15760) );
  XOR2_X1 U17828 ( .A(P1_EBX_REG_25__SCAN_IN), .B(keyinput_218), .Z(n15759) );
  XOR2_X1 U17829 ( .A(P1_EBX_REG_24__SCAN_IN), .B(keyinput_219), .Z(n15758) );
  AOI21_X1 U17830 ( .B1(n15760), .B2(n15759), .A(n15758), .ZN(n15773) );
  XOR2_X1 U17831 ( .A(P1_EBX_REG_21__SCAN_IN), .B(keyinput_222), .Z(n15764) );
  XOR2_X1 U17832 ( .A(P1_EBX_REG_23__SCAN_IN), .B(keyinput_220), .Z(n15763) );
  XOR2_X1 U17833 ( .A(P1_EBX_REG_19__SCAN_IN), .B(keyinput_224), .Z(n15762) );
  INV_X1 U17834 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n16842) );
  XNOR2_X1 U17835 ( .A(n16842), .B(keyinput_225), .ZN(n15761) );
  NOR4_X1 U17836 ( .A1(n15764), .A2(n15763), .A3(n15762), .A4(n15761), .ZN(
        n15767) );
  INV_X1 U17837 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n22261) );
  XNOR2_X1 U17838 ( .A(n22261), .B(keyinput_221), .ZN(n15766) );
  XOR2_X1 U17839 ( .A(P1_EBX_REG_20__SCAN_IN), .B(keyinput_223), .Z(n15765) );
  NAND3_X1 U17840 ( .A1(n15767), .A2(n15766), .A3(n15765), .ZN(n15772) );
  XOR2_X1 U17841 ( .A(P1_EBX_REG_17__SCAN_IN), .B(keyinput_226), .Z(n15771) );
  INV_X1 U17842 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n22195) );
  OAI22_X1 U17843 ( .A1(n22195), .A2(keyinput_227), .B1(P1_EBX_REG_15__SCAN_IN), .B2(keyinput_228), .ZN(n15769) );
  AND2_X1 U17844 ( .A1(P1_EBX_REG_15__SCAN_IN), .A2(keyinput_228), .ZN(n15768)
         );
  AOI211_X1 U17845 ( .C1(keyinput_227), .C2(n22195), .A(n15769), .B(n15768), 
        .ZN(n15770) );
  OAI211_X1 U17846 ( .C1(n15773), .C2(n15772), .A(n15771), .B(n15770), .ZN(
        n15778) );
  XNOR2_X1 U17847 ( .A(n15774), .B(keyinput_230), .ZN(n15777) );
  XNOR2_X1 U17848 ( .A(n22171), .B(keyinput_231), .ZN(n15776) );
  XNOR2_X1 U17849 ( .A(P1_EBX_REG_14__SCAN_IN), .B(keyinput_229), .ZN(n15775)
         );
  NAND4_X1 U17850 ( .A1(n15778), .A2(n15777), .A3(n15776), .A4(n15775), .ZN(
        n15783) );
  XOR2_X1 U17851 ( .A(P1_EBX_REG_11__SCAN_IN), .B(keyinput_232), .Z(n15782) );
  XNOR2_X1 U17852 ( .A(n15779), .B(keyinput_233), .ZN(n15781) );
  XNOR2_X1 U17853 ( .A(P1_EBX_REG_9__SCAN_IN), .B(keyinput_234), .ZN(n15780)
         );
  NAND4_X1 U17854 ( .A1(n15783), .A2(n15782), .A3(n15781), .A4(n15780), .ZN(
        n15786) );
  XNOR2_X1 U17855 ( .A(P1_EBX_REG_8__SCAN_IN), .B(keyinput_235), .ZN(n15785)
         );
  XNOR2_X1 U17856 ( .A(P1_EBX_REG_7__SCAN_IN), .B(keyinput_236), .ZN(n15784)
         );
  AOI21_X1 U17857 ( .B1(n15786), .B2(n15785), .A(n15784), .ZN(n15789) );
  XNOR2_X1 U17858 ( .A(n20701), .B(keyinput_237), .ZN(n15788) );
  XNOR2_X1 U17859 ( .A(P1_EBX_REG_5__SCAN_IN), .B(keyinput_238), .ZN(n15787)
         );
  OAI21_X1 U17860 ( .B1(n15789), .B2(n15788), .A(n15787), .ZN(n15793) );
  XOR2_X1 U17861 ( .A(P1_EBX_REG_4__SCAN_IN), .B(keyinput_239), .Z(n15792) );
  XNOR2_X1 U17862 ( .A(n15971), .B(keyinput_241), .ZN(n15791) );
  XNOR2_X1 U17863 ( .A(P1_EBX_REG_3__SCAN_IN), .B(keyinput_240), .ZN(n15790)
         );
  AOI211_X1 U17864 ( .C1(n15793), .C2(n15792), .A(n15791), .B(n15790), .ZN(
        n15800) );
  XOR2_X1 U17865 ( .A(P1_EAX_REG_31__SCAN_IN), .B(keyinput_244), .Z(n15796) );
  XNOR2_X1 U17866 ( .A(P1_EBX_REG_0__SCAN_IN), .B(keyinput_243), .ZN(n15795)
         );
  XNOR2_X1 U17867 ( .A(P1_EBX_REG_1__SCAN_IN), .B(keyinput_242), .ZN(n15794)
         );
  NAND3_X1 U17868 ( .A1(n15796), .A2(n15795), .A3(n15794), .ZN(n15799) );
  XOR2_X1 U17869 ( .A(P1_EAX_REG_29__SCAN_IN), .B(keyinput_246), .Z(n15798) );
  XOR2_X1 U17870 ( .A(P1_EAX_REG_30__SCAN_IN), .B(keyinput_245), .Z(n15797) );
  OAI211_X1 U17871 ( .C1(n15800), .C2(n15799), .A(n15798), .B(n15797), .ZN(
        n15804) );
  XNOR2_X1 U17872 ( .A(P1_EAX_REG_28__SCAN_IN), .B(keyinput_247), .ZN(n15803)
         );
  XOR2_X1 U17873 ( .A(P1_EAX_REG_27__SCAN_IN), .B(keyinput_248), .Z(n15802) );
  XNOR2_X1 U17874 ( .A(P1_EAX_REG_26__SCAN_IN), .B(keyinput_249), .ZN(n15801)
         );
  AOI211_X1 U17875 ( .C1(n15804), .C2(n15803), .A(n15802), .B(n15801), .ZN(
        n15808) );
  XOR2_X1 U17876 ( .A(P1_EAX_REG_25__SCAN_IN), .B(keyinput_250), .Z(n15807) );
  XOR2_X1 U17877 ( .A(P1_EAX_REG_24__SCAN_IN), .B(keyinput_251), .Z(n15806) );
  XNOR2_X1 U17878 ( .A(P1_EAX_REG_23__SCAN_IN), .B(keyinput_252), .ZN(n15805)
         );
  OAI211_X1 U17879 ( .C1(n15808), .C2(n15807), .A(n15806), .B(n15805), .ZN(
        n15812) );
  XOR2_X1 U17880 ( .A(P1_EAX_REG_22__SCAN_IN), .B(keyinput_253), .Z(n15811) );
  XNOR2_X1 U17881 ( .A(P1_EAX_REG_21__SCAN_IN), .B(keyinput_254), .ZN(n15810)
         );
  XNOR2_X1 U17882 ( .A(P1_EAX_REG_20__SCAN_IN), .B(keyinput_255), .ZN(n15809)
         );
  AOI211_X1 U17883 ( .C1(n15812), .C2(n15811), .A(n15810), .B(n15809), .ZN(
        n15996) );
  XOR2_X1 U17884 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(keyinput_0), .Z(n15816)
         );
  XOR2_X1 U17885 ( .A(DATAI_29_), .B(keyinput_3), .Z(n15815) );
  XOR2_X1 U17886 ( .A(DATAI_31_), .B(keyinput_1), .Z(n15814) );
  XOR2_X1 U17887 ( .A(DATAI_30_), .B(keyinput_2), .Z(n15813) );
  NAND4_X1 U17888 ( .A1(n15816), .A2(n15815), .A3(n15814), .A4(n15813), .ZN(
        n15819) );
  XOR2_X1 U17889 ( .A(DATAI_28_), .B(keyinput_4), .Z(n15818) );
  XNOR2_X1 U17890 ( .A(DATAI_27_), .B(keyinput_5), .ZN(n15817) );
  AOI21_X1 U17891 ( .B1(n15819), .B2(n15818), .A(n15817), .ZN(n15822) );
  XNOR2_X1 U17892 ( .A(DATAI_26_), .B(keyinput_6), .ZN(n15821) );
  XNOR2_X1 U17893 ( .A(DATAI_25_), .B(keyinput_7), .ZN(n15820) );
  NOR3_X1 U17894 ( .A1(n15822), .A2(n15821), .A3(n15820), .ZN(n15825) );
  XOR2_X1 U17895 ( .A(DATAI_24_), .B(keyinput_8), .Z(n15824) );
  XNOR2_X1 U17896 ( .A(DATAI_23_), .B(keyinput_9), .ZN(n15823) );
  NOR3_X1 U17897 ( .A1(n15825), .A2(n15824), .A3(n15823), .ZN(n15829) );
  XOR2_X1 U17898 ( .A(DATAI_22_), .B(keyinput_10), .Z(n15828) );
  XOR2_X1 U17899 ( .A(DATAI_20_), .B(keyinput_12), .Z(n15827) );
  XOR2_X1 U17900 ( .A(DATAI_21_), .B(keyinput_11), .Z(n15826) );
  OAI211_X1 U17901 ( .C1(n15829), .C2(n15828), .A(n15827), .B(n15826), .ZN(
        n15832) );
  XOR2_X1 U17902 ( .A(DATAI_18_), .B(keyinput_14), .Z(n15831) );
  XNOR2_X1 U17903 ( .A(DATAI_19_), .B(keyinput_13), .ZN(n15830) );
  NAND3_X1 U17904 ( .A1(n15832), .A2(n15831), .A3(n15830), .ZN(n15835) );
  XOR2_X1 U17905 ( .A(DATAI_17_), .B(keyinput_15), .Z(n15834) );
  XNOR2_X1 U17906 ( .A(DATAI_16_), .B(keyinput_16), .ZN(n15833) );
  NAND3_X1 U17907 ( .A1(n15835), .A2(n15834), .A3(n15833), .ZN(n15839) );
  XOR2_X1 U17908 ( .A(DATAI_14_), .B(keyinput_18), .Z(n15838) );
  XNOR2_X1 U17909 ( .A(DATAI_15_), .B(keyinput_17), .ZN(n15837) );
  XNOR2_X1 U17910 ( .A(DATAI_13_), .B(keyinput_19), .ZN(n15836) );
  NAND4_X1 U17911 ( .A1(n15839), .A2(n15838), .A3(n15837), .A4(n15836), .ZN(
        n15843) );
  XOR2_X1 U17912 ( .A(DATAI_10_), .B(keyinput_22), .Z(n15842) );
  XOR2_X1 U17913 ( .A(DATAI_11_), .B(keyinput_21), .Z(n15841) );
  XNOR2_X1 U17914 ( .A(DATAI_12_), .B(keyinput_20), .ZN(n15840) );
  NAND4_X1 U17915 ( .A1(n15843), .A2(n15842), .A3(n15841), .A4(n15840), .ZN(
        n15849) );
  XNOR2_X1 U17916 ( .A(DATAI_9_), .B(keyinput_23), .ZN(n15845) );
  XNOR2_X1 U17917 ( .A(DATAI_7_), .B(keyinput_25), .ZN(n15844) );
  NOR2_X1 U17918 ( .A1(n15845), .A2(n15844), .ZN(n15848) );
  XNOR2_X1 U17919 ( .A(DATAI_6_), .B(keyinput_26), .ZN(n15847) );
  XNOR2_X1 U17920 ( .A(DATAI_8_), .B(keyinput_24), .ZN(n15846) );
  NAND4_X1 U17921 ( .A1(n15849), .A2(n15848), .A3(n15847), .A4(n15846), .ZN(
        n15856) );
  XOR2_X1 U17922 ( .A(DATAI_1_), .B(keyinput_31), .Z(n15855) );
  XOR2_X1 U17923 ( .A(DATAI_5_), .B(keyinput_27), .Z(n15852) );
  XOR2_X1 U17924 ( .A(DATAI_2_), .B(keyinput_30), .Z(n15851) );
  XNOR2_X1 U17925 ( .A(DATAI_3_), .B(keyinput_29), .ZN(n15850) );
  NOR3_X1 U17926 ( .A1(n15852), .A2(n15851), .A3(n15850), .ZN(n15854) );
  XNOR2_X1 U17927 ( .A(DATAI_4_), .B(keyinput_28), .ZN(n15853) );
  NAND4_X1 U17928 ( .A1(n15856), .A2(n15855), .A3(n15854), .A4(n15853), .ZN(
        n15860) );
  XNOR2_X1 U17929 ( .A(NA), .B(keyinput_34), .ZN(n15859) );
  XNOR2_X1 U17930 ( .A(HOLD), .B(keyinput_33), .ZN(n15858) );
  XNOR2_X1 U17931 ( .A(DATAI_0_), .B(keyinput_32), .ZN(n15857) );
  NAND4_X1 U17932 ( .A1(n15860), .A2(n15859), .A3(n15858), .A4(n15857), .ZN(
        n15863) );
  XNOR2_X1 U17933 ( .A(BS16), .B(keyinput_35), .ZN(n15862) );
  XNOR2_X1 U17934 ( .A(READY1), .B(keyinput_36), .ZN(n15861) );
  AOI21_X1 U17935 ( .B1(n15863), .B2(n15862), .A(n15861), .ZN(n15866) );
  XNOR2_X1 U17936 ( .A(READY2), .B(keyinput_37), .ZN(n15865) );
  XNOR2_X1 U17937 ( .A(P1_READREQUEST_REG_SCAN_IN), .B(keyinput_38), .ZN(
        n15864) );
  NOR3_X1 U17938 ( .A1(n15866), .A2(n15865), .A3(n15864), .ZN(n15870) );
  XNOR2_X1 U17939 ( .A(n18025), .B(keyinput_39), .ZN(n15869) );
  XNOR2_X1 U17940 ( .A(n22804), .B(keyinput_41), .ZN(n15868) );
  XNOR2_X1 U17941 ( .A(P1_CODEFETCH_REG_SCAN_IN), .B(keyinput_40), .ZN(n15867)
         );
  NOR4_X1 U17942 ( .A1(n15870), .A2(n15869), .A3(n15868), .A4(n15867), .ZN(
        n15873) );
  XNOR2_X1 U17943 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .B(keyinput_43), .ZN(
        n15872) );
  XNOR2_X1 U17944 ( .A(P1_D_C_N_REG_SCAN_IN), .B(keyinput_42), .ZN(n15871) );
  NOR3_X1 U17945 ( .A1(n15873), .A2(n15872), .A3(n15871), .ZN(n15876) );
  XNOR2_X1 U17946 ( .A(n22305), .B(keyinput_44), .ZN(n15875) );
  XNOR2_X1 U17947 ( .A(n17987), .B(keyinput_45), .ZN(n15874) );
  OAI21_X1 U17948 ( .B1(n15876), .B2(n15875), .A(n15874), .ZN(n15883) );
  XOR2_X1 U17949 ( .A(P1_W_R_N_REG_SCAN_IN), .B(keyinput_47), .Z(n15880) );
  INV_X1 U17950 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20690) );
  XNOR2_X1 U17951 ( .A(n20690), .B(keyinput_49), .ZN(n15879) );
  XNOR2_X1 U17952 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .B(keyinput_48), .ZN(
        n15878) );
  XNOR2_X1 U17953 ( .A(P1_FLUSH_REG_SCAN_IN), .B(keyinput_46), .ZN(n15877) );
  NOR4_X1 U17954 ( .A1(n15880), .A2(n15879), .A3(n15878), .A4(n15877), .ZN(
        n15882) );
  XOR2_X1 U17955 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .B(keyinput_50), .Z(
        n15881) );
  AOI21_X1 U17956 ( .B1(n15883), .B2(n15882), .A(n15881), .ZN(n15890) );
  XOR2_X1 U17957 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(keyinput_51), .Z(
        n15887) );
  XNOR2_X1 U17958 ( .A(P1_REIP_REG_30__SCAN_IN), .B(keyinput_53), .ZN(n15886)
         );
  XNOR2_X1 U17959 ( .A(P1_REIP_REG_31__SCAN_IN), .B(keyinput_52), .ZN(n15885)
         );
  XNOR2_X1 U17960 ( .A(P1_REIP_REG_29__SCAN_IN), .B(keyinput_54), .ZN(n15884)
         );
  NAND4_X1 U17961 ( .A1(n15887), .A2(n15886), .A3(n15885), .A4(n15884), .ZN(
        n15889) );
  XOR2_X1 U17962 ( .A(P1_REIP_REG_28__SCAN_IN), .B(keyinput_55), .Z(n15888) );
  OAI21_X1 U17963 ( .B1(n15890), .B2(n15889), .A(n15888), .ZN(n15893) );
  XNOR2_X1 U17964 ( .A(P1_REIP_REG_27__SCAN_IN), .B(keyinput_56), .ZN(n15892)
         );
  XNOR2_X1 U17965 ( .A(P1_REIP_REG_26__SCAN_IN), .B(keyinput_57), .ZN(n15891)
         );
  AOI21_X1 U17966 ( .B1(n15893), .B2(n15892), .A(n15891), .ZN(n15896) );
  XNOR2_X1 U17967 ( .A(P1_REIP_REG_24__SCAN_IN), .B(keyinput_59), .ZN(n15895)
         );
  XNOR2_X1 U17968 ( .A(P1_REIP_REG_25__SCAN_IN), .B(keyinput_58), .ZN(n15894)
         );
  NOR3_X1 U17969 ( .A1(n15896), .A2(n15895), .A3(n15894), .ZN(n15899) );
  XNOR2_X1 U17970 ( .A(P1_REIP_REG_23__SCAN_IN), .B(keyinput_60), .ZN(n15898)
         );
  XNOR2_X1 U17971 ( .A(P1_REIP_REG_22__SCAN_IN), .B(keyinput_61), .ZN(n15897)
         );
  OAI21_X1 U17972 ( .B1(n15899), .B2(n15898), .A(n15897), .ZN(n15905) );
  XOR2_X1 U17973 ( .A(P1_REIP_REG_21__SCAN_IN), .B(keyinput_62), .Z(n15904) );
  XOR2_X1 U17974 ( .A(P1_REIP_REG_19__SCAN_IN), .B(keyinput_64), .Z(n15902) );
  XNOR2_X1 U17975 ( .A(P1_REIP_REG_18__SCAN_IN), .B(keyinput_65), .ZN(n15901)
         );
  XNOR2_X1 U17976 ( .A(P1_REIP_REG_20__SCAN_IN), .B(keyinput_63), .ZN(n15900)
         );
  NAND3_X1 U17977 ( .A1(n15902), .A2(n15901), .A3(n15900), .ZN(n15903) );
  AOI21_X1 U17978 ( .B1(n15905), .B2(n15904), .A(n15903), .ZN(n15909) );
  XNOR2_X1 U17979 ( .A(P1_REIP_REG_17__SCAN_IN), .B(keyinput_66), .ZN(n15908)
         );
  XOR2_X1 U17980 ( .A(P1_REIP_REG_16__SCAN_IN), .B(keyinput_67), .Z(n15907) );
  INV_X1 U17981 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n17024) );
  XNOR2_X1 U17982 ( .A(n17024), .B(keyinput_68), .ZN(n15906) );
  OAI211_X1 U17983 ( .C1(n15909), .C2(n15908), .A(n15907), .B(n15906), .ZN(
        n15916) );
  XOR2_X1 U17984 ( .A(P1_REIP_REG_10__SCAN_IN), .B(keyinput_73), .Z(n15915) );
  INV_X1 U17985 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n17064) );
  XNOR2_X1 U17986 ( .A(n17064), .B(keyinput_72), .ZN(n15914) );
  XOR2_X1 U17987 ( .A(P1_REIP_REG_14__SCAN_IN), .B(keyinput_69), .Z(n15912) );
  XOR2_X1 U17988 ( .A(P1_REIP_REG_12__SCAN_IN), .B(keyinput_71), .Z(n15911) );
  XNOR2_X1 U17989 ( .A(P1_REIP_REG_13__SCAN_IN), .B(keyinput_70), .ZN(n15910)
         );
  NOR3_X1 U17990 ( .A1(n15912), .A2(n15911), .A3(n15910), .ZN(n15913) );
  NAND4_X1 U17991 ( .A1(n15916), .A2(n15915), .A3(n15914), .A4(n15913), .ZN(
        n15922) );
  XOR2_X1 U17992 ( .A(P1_REIP_REG_9__SCAN_IN), .B(keyinput_74), .Z(n15921) );
  XNOR2_X1 U17993 ( .A(P1_REIP_REG_8__SCAN_IN), .B(keyinput_75), .ZN(n15920)
         );
  INV_X1 U17994 ( .A(keyinput_77), .ZN(n15917) );
  XNOR2_X1 U17995 ( .A(n15917), .B(P1_REIP_REG_6__SCAN_IN), .ZN(n15919) );
  XNOR2_X1 U17996 ( .A(P1_REIP_REG_5__SCAN_IN), .B(keyinput_78), .ZN(n15918)
         );
  NAND2_X1 U17997 ( .A1(n15919), .A2(n15918), .ZN(n15925) );
  AOI211_X1 U17998 ( .C1(n15922), .C2(n15921), .A(n15920), .B(n15925), .ZN(
        n15930) );
  XOR2_X1 U17999 ( .A(P1_REIP_REG_7__SCAN_IN), .B(keyinput_76), .Z(n15926) );
  XOR2_X1 U18000 ( .A(P1_REIP_REG_4__SCAN_IN), .B(keyinput_79), .Z(n15924) );
  XNOR2_X1 U18001 ( .A(P1_REIP_REG_3__SCAN_IN), .B(keyinput_80), .ZN(n15923)
         );
  OAI211_X1 U18002 ( .C1(n15926), .C2(n15925), .A(n15924), .B(n15923), .ZN(
        n15929) );
  XNOR2_X1 U18003 ( .A(P1_REIP_REG_1__SCAN_IN), .B(keyinput_82), .ZN(n15928)
         );
  XNOR2_X1 U18004 ( .A(P1_REIP_REG_2__SCAN_IN), .B(keyinput_81), .ZN(n15927)
         );
  OAI211_X1 U18005 ( .C1(n15930), .C2(n15929), .A(n15928), .B(n15927), .ZN(
        n15933) );
  XOR2_X1 U18006 ( .A(P1_REIP_REG_0__SCAN_IN), .B(keyinput_83), .Z(n15932) );
  XNOR2_X1 U18007 ( .A(P1_EBX_REG_31__SCAN_IN), .B(keyinput_84), .ZN(n15931)
         );
  NAND3_X1 U18008 ( .A1(n15933), .A2(n15932), .A3(n15931), .ZN(n15936) );
  XNOR2_X1 U18009 ( .A(P1_EBX_REG_30__SCAN_IN), .B(keyinput_85), .ZN(n15935)
         );
  XNOR2_X1 U18010 ( .A(P1_EBX_REG_29__SCAN_IN), .B(keyinput_86), .ZN(n15934)
         );
  AOI21_X1 U18011 ( .B1(n15936), .B2(n15935), .A(n15934), .ZN(n15940) );
  XOR2_X1 U18012 ( .A(P1_EBX_REG_27__SCAN_IN), .B(keyinput_88), .Z(n15939) );
  XNOR2_X1 U18013 ( .A(P1_EBX_REG_28__SCAN_IN), .B(keyinput_87), .ZN(n15938)
         );
  XNOR2_X1 U18014 ( .A(P1_EBX_REG_26__SCAN_IN), .B(keyinput_89), .ZN(n15937)
         );
  NOR4_X1 U18015 ( .A1(n15940), .A2(n15939), .A3(n15938), .A4(n15937), .ZN(
        n15943) );
  XOR2_X1 U18016 ( .A(P1_EBX_REG_25__SCAN_IN), .B(keyinput_90), .Z(n15942) );
  XOR2_X1 U18017 ( .A(P1_EBX_REG_24__SCAN_IN), .B(keyinput_91), .Z(n15941) );
  OAI21_X1 U18018 ( .B1(n15943), .B2(n15942), .A(n15941), .ZN(n15951) );
  XOR2_X1 U18019 ( .A(P1_EBX_REG_23__SCAN_IN), .B(keyinput_92), .Z(n15950) );
  XOR2_X1 U18020 ( .A(P1_EBX_REG_21__SCAN_IN), .B(keyinput_94), .Z(n15949) );
  XOR2_X1 U18021 ( .A(P1_EBX_REG_20__SCAN_IN), .B(keyinput_95), .Z(n15947) );
  XNOR2_X1 U18022 ( .A(n22261), .B(keyinput_93), .ZN(n15946) );
  XNOR2_X1 U18023 ( .A(n16842), .B(keyinput_97), .ZN(n15945) );
  XNOR2_X1 U18024 ( .A(P1_EBX_REG_19__SCAN_IN), .B(keyinput_96), .ZN(n15944)
         );
  NOR4_X1 U18025 ( .A1(n15947), .A2(n15946), .A3(n15945), .A4(n15944), .ZN(
        n15948) );
  NAND4_X1 U18026 ( .A1(n15951), .A2(n15950), .A3(n15949), .A4(n15948), .ZN(
        n15955) );
  XOR2_X1 U18027 ( .A(P1_EBX_REG_15__SCAN_IN), .B(keyinput_100), .Z(n15954) );
  XNOR2_X1 U18028 ( .A(P1_EBX_REG_16__SCAN_IN), .B(keyinput_99), .ZN(n15953)
         );
  XNOR2_X1 U18029 ( .A(P1_EBX_REG_17__SCAN_IN), .B(keyinput_98), .ZN(n15952)
         );
  NAND4_X1 U18030 ( .A1(n15955), .A2(n15954), .A3(n15953), .A4(n15952), .ZN(
        n15959) );
  XNOR2_X1 U18031 ( .A(n22171), .B(keyinput_103), .ZN(n15958) );
  XNOR2_X1 U18032 ( .A(P1_EBX_REG_13__SCAN_IN), .B(keyinput_102), .ZN(n15957)
         );
  XNOR2_X1 U18033 ( .A(P1_EBX_REG_14__SCAN_IN), .B(keyinput_101), .ZN(n15956)
         );
  NAND4_X1 U18034 ( .A1(n15959), .A2(n15958), .A3(n15957), .A4(n15956), .ZN(
        n15964) );
  XOR2_X1 U18035 ( .A(P1_EBX_REG_11__SCAN_IN), .B(keyinput_104), .Z(n15963) );
  XNOR2_X1 U18036 ( .A(n15960), .B(keyinput_106), .ZN(n15962) );
  XNOR2_X1 U18037 ( .A(P1_EBX_REG_10__SCAN_IN), .B(keyinput_105), .ZN(n15961)
         );
  NAND4_X1 U18038 ( .A1(n15964), .A2(n15963), .A3(n15962), .A4(n15961), .ZN(
        n15967) );
  XOR2_X1 U18039 ( .A(P1_EBX_REG_8__SCAN_IN), .B(keyinput_107), .Z(n15966) );
  XOR2_X1 U18040 ( .A(P1_EBX_REG_7__SCAN_IN), .B(keyinput_108), .Z(n15965) );
  AOI21_X1 U18041 ( .B1(n15967), .B2(n15966), .A(n15965), .ZN(n15970) );
  XNOR2_X1 U18042 ( .A(P1_EBX_REG_6__SCAN_IN), .B(keyinput_109), .ZN(n15969)
         );
  XOR2_X1 U18043 ( .A(P1_EBX_REG_5__SCAN_IN), .B(keyinput_110), .Z(n15968) );
  OAI21_X1 U18044 ( .B1(n15970), .B2(n15969), .A(n15968), .ZN(n15975) );
  XNOR2_X1 U18045 ( .A(P1_EBX_REG_4__SCAN_IN), .B(keyinput_111), .ZN(n15974)
         );
  XNOR2_X1 U18046 ( .A(n15971), .B(keyinput_113), .ZN(n15973) );
  XNOR2_X1 U18047 ( .A(P1_EBX_REG_3__SCAN_IN), .B(keyinput_112), .ZN(n15972)
         );
  AOI211_X1 U18048 ( .C1(n15975), .C2(n15974), .A(n15973), .B(n15972), .ZN(
        n15979) );
  XOR2_X1 U18049 ( .A(P1_EBX_REG_0__SCAN_IN), .B(keyinput_115), .Z(n15978) );
  XOR2_X1 U18050 ( .A(P1_EAX_REG_31__SCAN_IN), .B(keyinput_116), .Z(n15977) );
  XNOR2_X1 U18051 ( .A(P1_EBX_REG_1__SCAN_IN), .B(keyinput_114), .ZN(n15976)
         );
  NOR4_X1 U18052 ( .A1(n15979), .A2(n15978), .A3(n15977), .A4(n15976), .ZN(
        n15982) );
  XOR2_X1 U18053 ( .A(P1_EAX_REG_29__SCAN_IN), .B(keyinput_118), .Z(n15981) );
  XNOR2_X1 U18054 ( .A(P1_EAX_REG_30__SCAN_IN), .B(keyinput_117), .ZN(n15980)
         );
  NOR3_X1 U18055 ( .A1(n15982), .A2(n15981), .A3(n15980), .ZN(n15986) );
  XOR2_X1 U18056 ( .A(P1_EAX_REG_28__SCAN_IN), .B(keyinput_119), .Z(n15985) );
  XOR2_X1 U18057 ( .A(P1_EAX_REG_27__SCAN_IN), .B(keyinput_120), .Z(n15984) );
  XNOR2_X1 U18058 ( .A(P1_EAX_REG_26__SCAN_IN), .B(keyinput_121), .ZN(n15983)
         );
  OAI211_X1 U18059 ( .C1(n15986), .C2(n15985), .A(n15984), .B(n15983), .ZN(
        n15990) );
  XNOR2_X1 U18060 ( .A(P1_EAX_REG_25__SCAN_IN), .B(keyinput_122), .ZN(n15989)
         );
  XOR2_X1 U18061 ( .A(P1_EAX_REG_24__SCAN_IN), .B(keyinput_123), .Z(n15988) );
  XOR2_X1 U18062 ( .A(P1_EAX_REG_23__SCAN_IN), .B(keyinput_124), .Z(n15987) );
  AOI211_X1 U18063 ( .C1(n15990), .C2(n15989), .A(n15988), .B(n15987), .ZN(
        n15994) );
  XOR2_X1 U18064 ( .A(P1_EAX_REG_22__SCAN_IN), .B(keyinput_125), .Z(n15993) );
  XOR2_X1 U18065 ( .A(P1_EAX_REG_20__SCAN_IN), .B(keyinput_127), .Z(n15992) );
  XNOR2_X1 U18066 ( .A(P1_EAX_REG_21__SCAN_IN), .B(keyinput_126), .ZN(n15991)
         );
  OAI211_X1 U18067 ( .C1(n15994), .C2(n15993), .A(n15992), .B(n15991), .ZN(
        n15995) );
  NOR2_X1 U18068 ( .A1(n15996), .A2(n15995), .ZN(n15999) );
  AOI222_X1 U18069 ( .A1(n16855), .A2(n16008), .B1(n15997), .B2(n17073), .C1(
        P1_EAX_REG_10__SCAN_IN), .C2(n16890), .ZN(n15998) );
  XNOR2_X1 U18070 ( .A(n15999), .B(n15998), .ZN(P1_U2894) );
  INV_X1 U18071 ( .A(n16000), .ZN(n16001) );
  AOI21_X1 U18072 ( .B1(n16002), .B2(n16001), .A(n15529), .ZN(n17051) );
  INV_X1 U18073 ( .A(n17051), .ZN(n16010) );
  INV_X1 U18074 ( .A(n17322), .ZN(n16004) );
  AOI21_X1 U18075 ( .B1(n16004), .B2(n17299), .A(n16003), .ZN(n16006) );
  NOR2_X1 U18076 ( .A1(n16006), .A2(n16005), .ZN(n17296) );
  AOI22_X1 U18077 ( .A1(n17296), .A2(n20724), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n16821), .ZN(n16007) );
  OAI21_X1 U18078 ( .B1(n16010), .B2(n20698), .A(n16007), .ZN(P1_U2859) );
  AOI22_X1 U18079 ( .A1(n16008), .A2(n16847), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n16890), .ZN(n16009) );
  OAI21_X1 U18080 ( .B1(n16010), .B2(n16897), .A(n16009), .ZN(P1_U2891) );
  NAND2_X1 U18081 ( .A1(n17051), .A2(n22253), .ZN(n16016) );
  NOR2_X1 U18082 ( .A1(n22200), .A2(n16014), .ZN(n22179) );
  INV_X1 U18083 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n17047) );
  AOI22_X1 U18084 ( .A1(n17296), .A2(n22217), .B1(n22236), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n16011) );
  OAI211_X1 U18085 ( .C1(n22213), .C2(n16012), .A(n16011), .B(n22193), .ZN(
        n16013) );
  AOI221_X1 U18086 ( .B1(n22179), .B2(P1_REIP_REG_13__SCAN_IN), .C1(n16014), 
        .C2(n17047), .A(n16013), .ZN(n16015) );
  OAI211_X1 U18087 ( .C1(n22257), .C2(n17049), .A(n16016), .B(n16015), .ZN(
        P1_U2827) );
  OAI21_X1 U18088 ( .B1(n20545), .B2(n20274), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n16018) );
  NAND2_X1 U18089 ( .A1(n16018), .A2(n20100), .ZN(n16028) );
  INV_X1 U18090 ( .A(n16019), .ZN(n20430) );
  AOI21_X1 U18091 ( .B1(n17963), .B2(n19999), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19434) );
  NAND2_X1 U18092 ( .A1(n18114), .A2(n19434), .ZN(n16021) );
  NOR2_X1 U18093 ( .A1(n16021), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20101) );
  INV_X1 U18094 ( .A(n20101), .ZN(n20032) );
  OAI21_X1 U18095 ( .B1(n16023), .B2(n20032), .A(n19985), .ZN(n16024) );
  OAI21_X1 U18096 ( .B1(n16028), .B2(n20430), .A(n16024), .ZN(n16025) );
  NAND2_X1 U18097 ( .A1(n19998), .A2(n19952), .ZN(n20078) );
  INV_X1 U18098 ( .A(n20078), .ZN(n20093) );
  NAND2_X1 U18099 ( .A1(n20045), .A2(n20093), .ZN(n20538) );
  INV_X1 U18100 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16223) );
  INV_X1 U18101 ( .A(n20538), .ZN(n20268) );
  NOR2_X1 U18102 ( .A1(n20430), .A2(n20268), .ZN(n16027) );
  OAI21_X1 U18103 ( .B1(n12356), .B2(n20268), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16026) );
  AOI22_X1 U18104 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n11143), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20424), .ZN(n20310) );
  AOI22_X1 U18105 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n11143), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n20424), .ZN(n20315) );
  INV_X1 U18106 ( .A(n20315), .ZN(n20307) );
  NAND2_X1 U18107 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20086), .ZN(n20232) );
  AND2_X1 U18108 ( .A1(n16031), .A2(n20428), .ZN(n20311) );
  AOI22_X1 U18109 ( .A1(n20274), .A2(n20307), .B1(n20268), .B2(n20311), .ZN(
        n16032) );
  OAI21_X1 U18110 ( .B1(n20310), .B2(n20536), .A(n16032), .ZN(n16033) );
  AOI21_X1 U18111 ( .B1(n20543), .B2(n16029), .A(n16033), .ZN(n16034) );
  OAI21_X1 U18112 ( .B1(n20548), .B2(n16223), .A(n16034), .ZN(P2_U3051) );
  NOR2_X2 U18113 ( .A1(n16035), .A2(n20426), .ZN(n20419) );
  AOI22_X1 U18114 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n11143), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n20424), .ZN(n20423) );
  INV_X1 U18115 ( .A(n20423), .ZN(n20412) );
  AOI22_X1 U18116 ( .A1(n20274), .A2(n20412), .B1(n20268), .B2(n20418), .ZN(
        n16036) );
  OAI21_X1 U18117 ( .B1(n20415), .B2(n20536), .A(n16036), .ZN(n16037) );
  AOI21_X1 U18118 ( .B1(n20543), .B2(n20419), .A(n16037), .ZN(n16038) );
  OAI21_X1 U18119 ( .B1(n20548), .B2(n16516), .A(n16038), .ZN(P2_U3049) );
  XOR2_X1 U18120 ( .A(n16040), .B(n16039), .Z(n22163) );
  INV_X1 U18121 ( .A(n22163), .ZN(n16043) );
  INV_X1 U18122 ( .A(n16851), .ZN(n16042) );
  OAI222_X1 U18123 ( .A1(n16897), .A2(n16043), .B1(n16056), .B2(n16042), .C1(
        n16041), .C2(n16054), .ZN(P1_U2893) );
  INV_X1 U18124 ( .A(n16187), .ZN(n16044) );
  AOI21_X1 U18125 ( .B1(n16045), .B2(n15567), .A(n16044), .ZN(n17811) );
  INV_X1 U18126 ( .A(n17811), .ZN(n19215) );
  INV_X1 U18127 ( .A(n16046), .ZN(n16048) );
  INV_X1 U18128 ( .A(n16111), .ZN(n16047) );
  OR2_X1 U18129 ( .A1(n16046), .A2(n16111), .ZN(n16168) );
  OAI211_X1 U18130 ( .C1(n16048), .C2(n16047), .A(n17417), .B(n16168), .ZN(
        n16050) );
  NAND2_X1 U18131 ( .A1(n17423), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n16049) );
  OAI211_X1 U18132 ( .C1(n19215), .C2(n17420), .A(n16050), .B(n16049), .ZN(
        P2_U2872) );
  INV_X1 U18133 ( .A(n16051), .ZN(n16145) );
  NAND2_X1 U18134 ( .A1(n15530), .A2(n16052), .ZN(n16053) );
  NAND2_X1 U18135 ( .A1(n16145), .A2(n16053), .ZN(n20707) );
  OAI222_X1 U18136 ( .A1(n20707), .A2(n16897), .B1(n16056), .B2(n16055), .C1(
        n16054), .C2(n14214), .ZN(P1_U2889) );
  NOR2_X1 U18137 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19362) );
  AOI221_X1 U18138 ( .B1(n19100), .B2(n16057), .C1(n12397), .C2(n11181), .A(
        n17963), .ZN(n19357) );
  AOI211_X1 U18139 ( .C1(n16060), .C2(n16059), .A(n11181), .B(n16058), .ZN(
        n19111) );
  AOI21_X1 U18140 ( .B1(n11181), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n19111), .ZN(n16164) );
  INV_X1 U18141 ( .A(n16164), .ZN(n16061) );
  INV_X1 U18142 ( .A(n19435), .ZN(n16163) );
  AOI222_X1 U18143 ( .A1(n16062), .A2(n19362), .B1(n19357), .B2(n16061), .C1(
        n18127), .C2(n16163), .ZN(n16066) );
  OAI22_X1 U18144 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20083), .B1(n16063), 
        .B2(n19448), .ZN(n16064) );
  AOI21_X1 U18145 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n17962), .A(n16064), .ZN(
        n19358) );
  NAND2_X1 U18146 ( .A1(n19358), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16065) );
  OAI21_X1 U18147 ( .B1(n16066), .B2(n19358), .A(n16065), .ZN(P2_U3599) );
  AND2_X1 U18148 ( .A1(n16068), .A2(n16067), .ZN(n16070) );
  OAI21_X1 U18149 ( .B1(n16070), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n16069), .ZN(n18046) );
  OAI21_X1 U18150 ( .B1(n16073), .B2(n16072), .A(n16071), .ZN(n20170) );
  INV_X1 U18151 ( .A(n20170), .ZN(n16086) );
  AOI221_X1 U18152 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n16076), .C2(n16075), .A(
        n16074), .ZN(n16077) );
  AOI21_X1 U18153 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16078), .A(
        n16077), .ZN(n16080) );
  OR2_X1 U18154 ( .A1(n19258), .A2(n16079), .ZN(n18049) );
  OAI211_X1 U18155 ( .C1(n19416), .C2(n19122), .A(n16080), .B(n18049), .ZN(
        n16085) );
  OAI21_X1 U18156 ( .B1(n16081), .B2(n16083), .A(n16082), .ZN(n18048) );
  NOR2_X1 U18157 ( .A1(n18048), .A2(n19388), .ZN(n16084) );
  AOI211_X1 U18158 ( .C1(n19408), .C2(n16086), .A(n16085), .B(n16084), .ZN(
        n16087) );
  OAI21_X1 U18159 ( .B1(n19375), .B2(n18046), .A(n16087), .ZN(P2_U3041) );
  NAND2_X1 U18160 ( .A1(n16088), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16089) );
  NAND2_X1 U18161 ( .A1(n16090), .A2(n16089), .ZN(n16092) );
  XNOR2_X1 U18162 ( .A(n17256), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16091) );
  OAI21_X1 U18163 ( .B1(n16092), .B2(n16091), .A(n17061), .ZN(n22057) );
  AOI22_X1 U18164 ( .A1(n20760), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n22021), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n16093) );
  OAI21_X1 U18165 ( .B1(n20759), .B2(n16094), .A(n16093), .ZN(n16095) );
  AOI21_X1 U18166 ( .B1(n16096), .B2(n20762), .A(n16095), .ZN(n16097) );
  OAI21_X1 U18167 ( .B1(n22057), .B2(n22277), .A(n16097), .ZN(P1_U2990) );
  AOI22_X1 U18168 ( .A1(n16472), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n16416), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16104) );
  INV_X1 U18169 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n16099) );
  INV_X1 U18170 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16098) );
  OAI22_X1 U18171 ( .A1(n16474), .A2(n16099), .B1(n16473), .B2(n16098), .ZN(
        n16100) );
  AOI21_X1 U18172 ( .B1(n12024), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        n16100), .ZN(n16103) );
  AOI22_X1 U18173 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11944), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16102) );
  AOI22_X1 U18174 ( .A1(n16418), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11939), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16101) );
  NAND4_X1 U18175 ( .A1(n16104), .A2(n16103), .A3(n16102), .A4(n16101), .ZN(
        n16110) );
  AOI22_X1 U18176 ( .A1(n11978), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11905), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16108) );
  AOI22_X1 U18177 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n16481), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16107) );
  AOI22_X1 U18178 ( .A1(n16482), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n16424), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16106) );
  NAND2_X1 U18179 ( .A1(n16217), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n16105) );
  NAND4_X1 U18180 ( .A1(n16108), .A2(n16107), .A3(n16106), .A4(n16105), .ZN(
        n16109) );
  NOR2_X1 U18181 ( .A1(n16110), .A2(n16109), .ZN(n16169) );
  NOR2_X1 U18182 ( .A1(n16169), .A2(n16111), .ZN(n16113) );
  AND2_X1 U18183 ( .A1(n16113), .A2(n16112), .ZN(n16114) );
  AOI22_X1 U18184 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n16472), .B1(
        n16416), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n16122) );
  OAI22_X1 U18185 ( .A1(n16117), .A2(n16474), .B1(n16473), .B2(n16116), .ZN(
        n16118) );
  AOI21_X1 U18186 ( .B1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n12024), .A(
        n16118), .ZN(n16121) );
  AOI22_X1 U18187 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11944), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n16120) );
  AOI22_X1 U18188 ( .A1(n16418), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11939), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16119) );
  NAND4_X1 U18189 ( .A1(n16122), .A2(n16121), .A3(n16120), .A4(n16119), .ZN(
        n16128) );
  AOI22_X1 U18190 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11905), .B1(
        n11978), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16126) );
  AOI22_X1 U18191 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n16481), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16125) );
  AOI22_X1 U18192 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n16482), .B1(
        n16424), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16124) );
  NAND2_X1 U18193 ( .A1(n16217), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n16123) );
  NAND4_X1 U18194 ( .A1(n16126), .A2(n16125), .A3(n16124), .A4(n16123), .ZN(
        n16127) );
  OR2_X1 U18195 ( .A1(n16128), .A2(n16127), .ZN(n16131) );
  INV_X1 U18196 ( .A(n16210), .ZN(n16130) );
  OAI21_X1 U18197 ( .B1(n16129), .B2(n16131), .A(n16130), .ZN(n16185) );
  NOR2_X2 U18198 ( .A1(n16141), .A2(n20174), .ZN(n17479) );
  XNOR2_X1 U18199 ( .A(n16172), .B(n16132), .ZN(n19241) );
  OAI22_X1 U18200 ( .A1(n19241), .A2(n17477), .B1(n17475), .B2(n16133), .ZN(
        n16134) );
  AOI21_X1 U18201 ( .B1(n17479), .B2(n16135), .A(n16134), .ZN(n16143) );
  INV_X1 U18202 ( .A(n16141), .ZN(n16138) );
  NOR2_X1 U18203 ( .A1(n16136), .A2(n16139), .ZN(n16137) );
  NAND2_X1 U18204 ( .A1(n16138), .A2(n16137), .ZN(n20327) );
  NAND2_X1 U18205 ( .A1(n11649), .A2(n16139), .ZN(n16140) );
  NOR2_X2 U18206 ( .A1(n16141), .A2(n16140), .ZN(n19915) );
  AOI22_X1 U18207 ( .A1(n19914), .A2(BUF2_REG_17__SCAN_IN), .B1(n19915), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n16142) );
  OAI211_X1 U18208 ( .C1(n16185), .C2(n20165), .A(n16143), .B(n16142), .ZN(
        P2_U2902) );
  AND2_X1 U18209 ( .A1(n16145), .A2(n16144), .ZN(n16148) );
  INV_X1 U18210 ( .A(n16146), .ZN(n16147) );
  OR2_X1 U18211 ( .A1(n16148), .A2(n16147), .ZN(n22205) );
  AOI22_X1 U18212 ( .A1(n16891), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n16890), .ZN(n16154) );
  NOR3_X1 U18213 ( .A1(n16890), .A2(n16150), .A3(n11160), .ZN(n16151) );
  AOI22_X1 U18214 ( .A1(n16894), .A2(n16152), .B1(n16892), .B2(DATAI_16_), 
        .ZN(n16153) );
  OAI211_X1 U18215 ( .C1(n22205), .C2(n16897), .A(n16154), .B(n16153), .ZN(
        P1_U2888) );
  MUX2_X1 U18216 ( .A(n16297), .B(n16321), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n16156) );
  OAI21_X1 U18217 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16323), .A(
        n16156), .ZN(n17279) );
  INV_X1 U18218 ( .A(n17281), .ZN(n16162) );
  NAND2_X1 U18219 ( .A1(n16293), .A2(n22195), .ZN(n16159) );
  INV_X1 U18220 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17076) );
  NAND2_X1 U18221 ( .A1(n14857), .A2(n17076), .ZN(n16157) );
  OAI211_X1 U18222 ( .C1(P1_EBX_REG_16__SCAN_IN), .C2(n11150), .A(n16157), .B(
        n16385), .ZN(n16158) );
  INV_X1 U18223 ( .A(n16160), .ZN(n16161) );
  INV_X1 U18224 ( .A(n16275), .ZN(n17259) );
  OAI21_X1 U18225 ( .B1(n16162), .B2(n16161), .A(n17259), .ZN(n22208) );
  OAI222_X1 U18226 ( .A1(n22205), .A2(n20698), .B1(n22195), .B2(n20727), .C1(
        n22208), .C2(n16841), .ZN(P1_U2856) );
  AOI222_X1 U18227 ( .A1(n19362), .A2(n16165), .B1(n19357), .B2(n16164), .C1(
        n19944), .C2(n16163), .ZN(n16167) );
  NAND2_X1 U18228 ( .A1(n19358), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n16166) );
  OAI21_X1 U18229 ( .B1(n16167), .B2(n19358), .A(n16166), .ZN(P2_U3600) );
  AOI21_X1 U18230 ( .B1(n16169), .B2(n16168), .A(n16129), .ZN(n16190) );
  INV_X1 U18231 ( .A(n16190), .ZN(n16180) );
  AND2_X1 U18232 ( .A1(n16171), .A2(n16170), .ZN(n16173) );
  OR2_X1 U18233 ( .A1(n16173), .A2(n16172), .ZN(n19233) );
  OAI22_X1 U18234 ( .A1(n17477), .A2(n19233), .B1(n17475), .B2(n16174), .ZN(
        n16177) );
  INV_X1 U18235 ( .A(n19915), .ZN(n20317) );
  INV_X1 U18236 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n16175) );
  OAI22_X1 U18237 ( .A1(n20317), .A2(n20797), .B1(n20327), .B2(n16175), .ZN(
        n16176) );
  AOI211_X1 U18238 ( .C1(n17479), .C2(n16178), .A(n16177), .B(n16176), .ZN(
        n16179) );
  OAI21_X1 U18239 ( .B1(n16180), .B2(n20165), .A(n16179), .ZN(P2_U2903) );
  AND2_X1 U18240 ( .A1(n16189), .A2(n16181), .ZN(n16182) );
  OR2_X1 U18241 ( .A1(n16182), .A2(n16194), .ZN(n19242) );
  NOR2_X1 U18242 ( .A1(n19242), .A2(n17420), .ZN(n16183) );
  AOI21_X1 U18243 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n17420), .A(n16183), .ZN(
        n16184) );
  OAI21_X1 U18244 ( .B1(n16185), .B2(n17428), .A(n16184), .ZN(P2_U2870) );
  NAND2_X1 U18245 ( .A1(n16187), .A2(n16186), .ZN(n16188) );
  NAND2_X1 U18246 ( .A1(n16189), .A2(n16188), .ZN(n17799) );
  NAND2_X1 U18247 ( .A1(n16190), .A2(n17417), .ZN(n16192) );
  NAND2_X1 U18248 ( .A1(n17423), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n16191) );
  OAI211_X1 U18249 ( .C1(n17799), .C2(n17420), .A(n16192), .B(n16191), .ZN(
        P2_U2871) );
  OR2_X1 U18250 ( .A1(n16194), .A2(n16193), .ZN(n16196) );
  AND2_X1 U18251 ( .A1(n16196), .A2(n16195), .ZN(n19253) );
  INV_X1 U18252 ( .A(n19253), .ZN(n17773) );
  AOI22_X1 U18253 ( .A1(n16472), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16416), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16203) );
  INV_X1 U18254 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16197) );
  OAI22_X1 U18255 ( .A1(n16474), .A2(n16198), .B1(n16473), .B2(n16197), .ZN(
        n16199) );
  AOI21_X1 U18256 ( .B1(n12024), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n16199), .ZN(n16202) );
  AOI22_X1 U18257 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11944), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16201) );
  AOI22_X1 U18258 ( .A1(n16418), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11939), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16200) );
  NAND4_X1 U18259 ( .A1(n16203), .A2(n16202), .A3(n16201), .A4(n16200), .ZN(
        n16209) );
  AOI22_X1 U18260 ( .A1(n11978), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11905), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16207) );
  AOI22_X1 U18261 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16481), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n16206) );
  AOI22_X1 U18262 ( .A1(n16482), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16424), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16205) );
  NAND2_X1 U18263 ( .A1(n16217), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n16204) );
  NAND4_X1 U18264 ( .A1(n16207), .A2(n16206), .A3(n16205), .A4(n16204), .ZN(
        n16208) );
  OR2_X1 U18265 ( .A1(n16209), .A2(n16208), .ZN(n16211) );
  OR2_X1 U18266 ( .A1(n16210), .A2(n16211), .ZN(n16212) );
  AND2_X1 U18267 ( .A1(n16233), .A2(n16212), .ZN(n20323) );
  NAND2_X1 U18268 ( .A1(n20323), .A2(n17417), .ZN(n16214) );
  NAND2_X1 U18269 ( .A1(n17423), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n16213) );
  OAI211_X1 U18270 ( .C1(n17773), .C2(n17420), .A(n16214), .B(n16213), .ZN(
        P2_U2869) );
  AOI21_X1 U18271 ( .B1(n16216), .B2(n16195), .A(n11400), .ZN(n19266) );
  INV_X1 U18272 ( .A(n19266), .ZN(n16237) );
  INV_X1 U18273 ( .A(n16217), .ZN(n16436) );
  INV_X1 U18274 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16220) );
  AOI22_X1 U18275 ( .A1(n11978), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11905), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16219) );
  AOI22_X1 U18276 ( .A1(n16482), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16424), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16218) );
  OAI211_X1 U18277 ( .C1(n16436), .C2(n16220), .A(n16219), .B(n16218), .ZN(
        n16232) );
  AOI22_X1 U18278 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11944), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16222) );
  AOI22_X1 U18279 ( .A1(n16449), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16448), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16221) );
  OAI211_X1 U18280 ( .C1(n16452), .C2(n16223), .A(n16222), .B(n16221), .ZN(
        n16231) );
  AOI22_X1 U18281 ( .A1(n16472), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n16416), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16225) );
  AOI22_X1 U18282 ( .A1(n16418), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11939), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16224) );
  NAND2_X1 U18283 ( .A1(n16225), .A2(n16224), .ZN(n16230) );
  INV_X1 U18284 ( .A(n16226), .ZN(n16443) );
  INV_X1 U18285 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16228) );
  INV_X1 U18286 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16227) );
  OAI22_X1 U18287 ( .A1(n16443), .A2(n16228), .B1(n16441), .B2(n16227), .ZN(
        n16229) );
  NOR4_X1 U18288 ( .A1(n16232), .A2(n16231), .A3(n16230), .A4(n16229), .ZN(
        n16234) );
  AOI21_X1 U18289 ( .B1(n16234), .B2(n16233), .A(n16432), .ZN(n16243) );
  NAND2_X1 U18290 ( .A1(n16243), .A2(n17417), .ZN(n16236) );
  NAND2_X1 U18291 ( .A1(n17423), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n16235) );
  OAI211_X1 U18292 ( .C1(n16237), .C2(n17420), .A(n16236), .B(n16235), .ZN(
        P2_U2868) );
  INV_X1 U18293 ( .A(n17479), .ZN(n20316) );
  AOI22_X1 U18294 ( .A1(n19914), .A2(BUF2_REG_19__SCAN_IN), .B1(n19915), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n16240) );
  AOI21_X1 U18295 ( .B1(n16238), .B2(n17770), .A(n17743), .ZN(n17754) );
  AOI22_X1 U18296 ( .A1(n20321), .A2(n17754), .B1(n20319), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n16239) );
  OAI211_X1 U18297 ( .C1(n16241), .C2(n20316), .A(n16240), .B(n16239), .ZN(
        n16242) );
  AOI21_X1 U18298 ( .B1(n16243), .B2(n20322), .A(n16242), .ZN(n16244) );
  INV_X1 U18299 ( .A(n16244), .ZN(P2_U2900) );
  NAND4_X1 U18300 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .A3(P3_EBX_REG_13__SCAN_IN), .A4(P3_EBX_REG_12__SCAN_IN), .ZN(n18322)
         );
  NOR2_X1 U18301 ( .A1(n18322), .A2(n18291), .ZN(n18239) );
  AND3_X1 U18302 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_12__SCAN_IN), .ZN(n16245) );
  AOI21_X1 U18303 ( .B1(n16245), .B2(n18290), .A(P3_EBX_REG_15__SCAN_IN), .ZN(
        n16246) );
  NOR2_X1 U18304 ( .A1(n18239), .A2(n16246), .ZN(n16258) );
  AOI22_X1 U18305 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16250) );
  AOI22_X1 U18306 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18381), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16249) );
  AOI22_X1 U18307 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16248) );
  AOI22_X1 U18308 ( .A1(n18279), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16247) );
  NAND4_X1 U18309 ( .A1(n16250), .A2(n16249), .A3(n16248), .A4(n16247), .ZN(
        n16256) );
  AOI22_X1 U18310 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16254) );
  AOI22_X1 U18311 ( .A1(n18547), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11157), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16253) );
  AOI22_X1 U18312 ( .A1(n18393), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18480), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16252) );
  NAND4_X1 U18313 ( .A1(n16254), .A2(n16253), .A3(n16252), .A4(n16251), .ZN(
        n16255) );
  NOR2_X1 U18314 ( .A1(n16256), .A2(n16255), .ZN(n21508) );
  INV_X1 U18315 ( .A(n21508), .ZN(n16257) );
  MUX2_X1 U18316 ( .A(n16258), .B(n16257), .S(n18565), .Z(P3_U2688) );
  NOR2_X1 U18317 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21555) );
  INV_X1 U18318 ( .A(n21555), .ZN(n21545) );
  NOR2_X1 U18319 ( .A1(n16259), .A2(n21545), .ZN(n16262) );
  NAND2_X1 U18320 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18572), .ZN(n17935) );
  INV_X1 U18321 ( .A(n17935), .ZN(n21946) );
  NOR2_X1 U18322 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21949), .ZN(n21945) );
  NOR2_X1 U18323 ( .A1(n16260), .A2(n21961), .ZN(n16261) );
  AOI211_X2 U18324 ( .C1(n21946), .C2(P3_FLUSH_REG_SCAN_IN), .A(n21945), .B(
        n16261), .ZN(n21560) );
  MUX2_X1 U18325 ( .A(n16262), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n21560), .Z(P3_U3284) );
  NAND2_X2 U18326 ( .A1(n16266), .A2(n16265), .ZN(n16927) );
  AOI22_X1 U18327 ( .A1(n16891), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n16890), .ZN(n16269) );
  AOI22_X1 U18328 ( .A1(n16894), .A2(n16267), .B1(n16892), .B2(DATAI_28_), 
        .ZN(n16268) );
  OAI211_X1 U18329 ( .C1(n16927), .C2(n16897), .A(n16269), .B(n16268), .ZN(
        P1_U2876) );
  INV_X1 U18330 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n16306) );
  MUX2_X1 U18331 ( .A(n16297), .B(n16321), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n16273) );
  INV_X1 U18332 ( .A(n16323), .ZN(n16271) );
  INV_X1 U18333 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16270) );
  NAND2_X1 U18334 ( .A1(n16271), .A2(n16270), .ZN(n16272) );
  NAND2_X1 U18335 ( .A1(n16273), .A2(n16272), .ZN(n17260) );
  INV_X1 U18336 ( .A(n17260), .ZN(n16274) );
  NAND2_X1 U18337 ( .A1(n16275), .A2(n16274), .ZN(n16837) );
  NAND2_X1 U18338 ( .A1(n16293), .A2(n16842), .ZN(n16279) );
  NAND2_X1 U18339 ( .A1(n16385), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16276) );
  NAND2_X1 U18340 ( .A1(n14857), .A2(n16276), .ZN(n16277) );
  OAI21_X1 U18341 ( .B1(P1_EBX_REG_18__SCAN_IN), .B2(n11150), .A(n16277), .ZN(
        n16278) );
  AND2_X1 U18342 ( .A1(n16279), .A2(n16278), .ZN(n16838) );
  OR2_X2 U18343 ( .A1(n16837), .A2(n16838), .ZN(n16839) );
  MUX2_X1 U18344 ( .A(n16297), .B(n16321), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n16280) );
  OAI21_X1 U18345 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16323), .A(
        n16280), .ZN(n16805) );
  INV_X1 U18346 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17222) );
  NAND2_X1 U18347 ( .A1(n14857), .A2(n17222), .ZN(n16281) );
  OAI211_X1 U18348 ( .C1(P1_EBX_REG_20__SCAN_IN), .C2(n11150), .A(n16281), .B(
        n16385), .ZN(n16282) );
  OAI21_X1 U18349 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(n16304), .A(n16282), .ZN(
        n16829) );
  MUX2_X1 U18350 ( .A(n16297), .B(n16321), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n16283) );
  OAI21_X1 U18351 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n16323), .A(
        n16283), .ZN(n17209) );
  NAND2_X1 U18352 ( .A1(n16293), .A2(n22261), .ZN(n16287) );
  NAND2_X1 U18353 ( .A1(n16385), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16284) );
  NAND2_X1 U18354 ( .A1(n14857), .A2(n16284), .ZN(n16285) );
  OAI21_X1 U18355 ( .B1(P1_EBX_REG_22__SCAN_IN), .B2(n11150), .A(n16285), .ZN(
        n16286) );
  MUX2_X1 U18356 ( .A(n16297), .B(n16321), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n16288) );
  OAI21_X1 U18357 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16323), .A(
        n16288), .ZN(n16793) );
  INV_X1 U18358 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17172) );
  NAND2_X1 U18359 ( .A1(n14857), .A2(n17172), .ZN(n16289) );
  OAI211_X1 U18360 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n11150), .A(n16289), .B(
        n16385), .ZN(n16290) );
  OAI21_X1 U18361 ( .B1(P1_EBX_REG_24__SCAN_IN), .B2(n16304), .A(n16290), .ZN(
        n16783) );
  NAND2_X1 U18362 ( .A1(n16792), .A2(n16783), .ZN(n16770) );
  MUX2_X1 U18363 ( .A(n16297), .B(n16321), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n16291) );
  OAI21_X1 U18364 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n16323), .A(
        n16291), .ZN(n16771) );
  INV_X1 U18365 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n16292) );
  NAND2_X1 U18366 ( .A1(n16293), .A2(n16292), .ZN(n16296) );
  INV_X1 U18367 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17097) );
  NAND2_X1 U18368 ( .A1(n14857), .A2(n17097), .ZN(n16294) );
  OAI211_X1 U18369 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n11150), .A(n16294), .B(
        n16385), .ZN(n16295) );
  AND2_X1 U18370 ( .A1(n16296), .A2(n16295), .ZN(n16759) );
  MUX2_X1 U18371 ( .A(n16297), .B(n16321), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n16299) );
  OR2_X1 U18372 ( .A1(n16323), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16298) );
  NAND2_X1 U18373 ( .A1(n16299), .A2(n16298), .ZN(n16749) );
  INV_X1 U18374 ( .A(n16749), .ZN(n16300) );
  INV_X1 U18375 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16301) );
  NAND2_X1 U18376 ( .A1(n14857), .A2(n16301), .ZN(n16302) );
  OAI211_X1 U18377 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n11150), .A(n16302), .B(
        n16385), .ZN(n16303) );
  OAI21_X1 U18378 ( .B1(P1_EBX_REG_28__SCAN_IN), .B2(n16304), .A(n16303), .ZN(
        n16305) );
  OAI21_X1 U18379 ( .B1(n16747), .B2(n16305), .A(n16736), .ZN(n17136) );
  OAI222_X1 U18380 ( .A1(n20698), .A2(n16927), .B1(n16306), .B2(n20727), .C1(
        n17136), .C2(n16841), .ZN(P1_U2844) );
  NAND4_X1 U18381 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(P1_REIP_REG_16__SCAN_IN), .A4(P1_REIP_REG_14__SCAN_IN), .ZN(n16308) );
  NAND4_X1 U18382 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .A4(P1_REIP_REG_13__SCAN_IN), .ZN(n16307) );
  NOR3_X1 U18383 ( .A1(n22170), .A2(n16308), .A3(n16307), .ZN(n22234) );
  NAND2_X1 U18384 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n22234), .ZN(n22244) );
  OAI21_X1 U18385 ( .B1(n16309), .B2(n22244), .A(n22210), .ZN(n22248) );
  OAI21_X1 U18386 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n22245), .A(n22248), 
        .ZN(n22259) );
  NOR2_X1 U18387 ( .A1(n22245), .A2(n22259), .ZN(n22273) );
  NAND3_X1 U18388 ( .A1(n16797), .A2(P1_REIP_REG_23__SCAN_IN), .A3(
        P1_REIP_REG_24__SCAN_IN), .ZN(n16776) );
  INV_X1 U18389 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n16952) );
  NAND2_X1 U18390 ( .A1(n16774), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n16762) );
  INV_X1 U18391 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n16934) );
  NOR2_X1 U18392 ( .A1(n16762), .A2(n16934), .ZN(n16310) );
  NAND2_X1 U18393 ( .A1(n16310), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n16733) );
  INV_X1 U18394 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n16311) );
  INV_X1 U18395 ( .A(n16310), .ZN(n16754) );
  OAI21_X1 U18396 ( .B1(n22200), .B2(n16311), .A(n16754), .ZN(n16315) );
  AOI22_X1 U18397 ( .A1(n22264), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n22236), .B2(P1_EBX_REG_28__SCAN_IN), .ZN(n16313) );
  NAND2_X1 U18398 ( .A1(n22266), .A2(n16930), .ZN(n16312) );
  OAI211_X1 U18399 ( .C1(n17136), .C2(n22276), .A(n16313), .B(n16312), .ZN(
        n16314) );
  AOI21_X1 U18400 ( .B1(n16733), .B2(n16315), .A(n16314), .ZN(n16316) );
  OAI21_X1 U18401 ( .B1(n16927), .B2(n22269), .A(n16316), .ZN(P1_U2812) );
  INV_X1 U18402 ( .A(n16380), .ZN(n16333) );
  AND2_X1 U18403 ( .A1(n11150), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16317) );
  AOI21_X1 U18404 ( .B1(n16323), .B2(P1_EBX_REG_30__SCAN_IN), .A(n16317), .ZN(
        n16387) );
  OR2_X1 U18405 ( .A1(n16323), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16319) );
  NAND2_X1 U18406 ( .A1(n11192), .A2(n16815), .ZN(n16318) );
  NAND2_X1 U18407 ( .A1(n16319), .A2(n16318), .ZN(n16384) );
  MUX2_X1 U18408 ( .A(n16384), .B(P1_EBX_REG_29__SCAN_IN), .S(n16320), .Z(
        n16735) );
  NOR2_X2 U18409 ( .A1(n16736), .A2(n16735), .ZN(n16738) );
  MUX2_X1 U18410 ( .A(n16321), .B(n16387), .S(n16738), .Z(n16326) );
  AOI22_X1 U18411 ( .A1(n16323), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n11150), .ZN(n16324) );
  INV_X1 U18412 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n16813) );
  OAI22_X1 U18413 ( .A1(n22213), .A2(n16327), .B1(n16813), .B2(n22262), .ZN(
        n16328) );
  AOI21_X1 U18414 ( .B1(n17106), .B2(n22217), .A(n16328), .ZN(n16332) );
  INV_X1 U18415 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n16912) );
  NOR2_X1 U18416 ( .A1(n16733), .A2(n16912), .ZN(n16732) );
  NAND2_X1 U18417 ( .A1(n16732), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n16330) );
  NAND2_X1 U18418 ( .A1(n16330), .A2(n22210), .ZN(n16329) );
  MUX2_X1 U18419 ( .A(n16330), .B(n16329), .S(P1_REIP_REG_31__SCAN_IN), .Z(
        n16331) );
  OAI211_X1 U18420 ( .C1(n16333), .C2(n22269), .A(n16332), .B(n16331), .ZN(
        P1_U2809) );
  INV_X1 U18421 ( .A(n16334), .ZN(n16335) );
  OAI21_X1 U18422 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19091), .A(
        n16335), .ZN(n19371) );
  INV_X1 U18423 ( .A(n19371), .ZN(n16340) );
  OAI21_X1 U18424 ( .B1(n16337), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n16336), .ZN(n19376) );
  OR2_X1 U18425 ( .A1(n19258), .A2(n16338), .ZN(n19373) );
  OAI21_X1 U18426 ( .B1(n18103), .B2(n19376), .A(n19373), .ZN(n16339) );
  AOI21_X1 U18427 ( .B1(n18079), .B2(n16340), .A(n16339), .ZN(n16343) );
  OAI21_X1 U18428 ( .B1(n18102), .B2(n16341), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16342) );
  OAI211_X1 U18429 ( .C1(n18105), .C2(n16344), .A(n16343), .B(n16342), .ZN(
        P2_U3014) );
  NAND2_X1 U18430 ( .A1(n11541), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16345) );
  XNOR2_X1 U18431 ( .A(n17250), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17046) );
  INV_X1 U18432 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17311) );
  NAND2_X1 U18433 ( .A1(n17250), .A2(n17311), .ZN(n17044) );
  NAND2_X1 U18434 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16346) );
  NAND2_X1 U18435 ( .A1(n17250), .A2(n16346), .ZN(n17042) );
  AND2_X1 U18436 ( .A1(n17044), .A2(n17042), .ZN(n16347) );
  NAND2_X1 U18437 ( .A1(n17046), .A2(n16347), .ZN(n17028) );
  AND2_X1 U18438 ( .A1(n17256), .A2(n16348), .ZN(n16349) );
  NOR2_X1 U18439 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16350) );
  XNOR2_X1 U18440 ( .A(n17256), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17016) );
  INV_X1 U18441 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17284) );
  NAND2_X1 U18442 ( .A1(n17256), .A2(n17284), .ZN(n17014) );
  NAND2_X1 U18443 ( .A1(n17016), .A2(n17014), .ZN(n16351) );
  AOI21_X1 U18444 ( .B1(n17009), .B2(n16354), .A(n16351), .ZN(n17252) );
  NAND2_X1 U18445 ( .A1(n17256), .A2(n16270), .ZN(n16352) );
  OR2_X1 U18446 ( .A1(n17250), .A2(n17311), .ZN(n17043) );
  NOR2_X1 U18447 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16353) );
  NAND2_X1 U18448 ( .A1(n17029), .A2(n16354), .ZN(n17010) );
  NOR2_X1 U18449 ( .A1(n17256), .A2(n17284), .ZN(n17013) );
  OAI21_X1 U18450 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n11541), .ZN(n16355) );
  NAND2_X1 U18451 ( .A1(n17251), .A2(n16355), .ZN(n16356) );
  AND2_X1 U18452 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17192) );
  NAND2_X1 U18453 ( .A1(n17192), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n17198) );
  INV_X1 U18454 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17244) );
  INV_X1 U18455 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17080) );
  NOR4_X1 U18456 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16357) );
  AOI21_X1 U18457 ( .B1(n17004), .B2(n16357), .A(n17256), .ZN(n16975) );
  NOR2_X1 U18458 ( .A1(n16358), .A2(n16975), .ZN(n16918) );
  NOR3_X1 U18459 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16920) );
  INV_X1 U18460 ( .A(n16358), .ZN(n16948) );
  NAND2_X1 U18461 ( .A1(n16358), .A2(n17256), .ZN(n16359) );
  AND2_X1 U18462 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17163) );
  NAND2_X1 U18463 ( .A1(n17163), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17155) );
  NAND2_X1 U18464 ( .A1(n17256), .A2(n17155), .ZN(n16919) );
  NAND2_X1 U18465 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17122) );
  INV_X1 U18466 ( .A(n17122), .ZN(n16360) );
  NOR2_X1 U18467 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17132) );
  NAND2_X1 U18468 ( .A1(n16363), .A2(n16899), .ZN(n16910) );
  INV_X1 U18469 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17099) );
  XNOR2_X1 U18470 ( .A(n17256), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16367) );
  INV_X1 U18471 ( .A(n16367), .ZN(n16364) );
  OAI21_X1 U18472 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(n11541), .ZN(n16369) );
  NAND2_X1 U18473 ( .A1(n16364), .A2(n16369), .ZN(n16365) );
  OR2_X2 U18474 ( .A1(n16368), .A2(n16365), .ZN(n16376) );
  INV_X1 U18475 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16366) );
  NAND2_X1 U18476 ( .A1(n17256), .A2(n16366), .ZN(n16370) );
  NAND3_X1 U18477 ( .A1(n16368), .A2(n16367), .A3(n16370), .ZN(n16375) );
  INV_X1 U18478 ( .A(n16369), .ZN(n16372) );
  INV_X1 U18479 ( .A(n16370), .ZN(n16371) );
  NOR2_X1 U18480 ( .A1(n16372), .A2(n16371), .ZN(n16373) );
  OR2_X1 U18481 ( .A1(n16373), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16374) );
  NAND2_X1 U18482 ( .A1(n22021), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n17101) );
  NAND2_X1 U18483 ( .A1(n20760), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16377) );
  OAI211_X1 U18484 ( .C1(n16378), .C2(n20759), .A(n17101), .B(n16377), .ZN(
        n16379) );
  AOI21_X1 U18485 ( .B1(n16380), .B2(n20762), .A(n16379), .ZN(n16381) );
  OAI21_X1 U18486 ( .B1(n17108), .B2(n22277), .A(n16381), .ZN(P1_U2968) );
  AOI21_X1 U18487 ( .B1(n16383), .B2(n16729), .A(n16382), .ZN(n16908) );
  INV_X1 U18488 ( .A(n16908), .ZN(n16846) );
  OAI22_X1 U18489 ( .A1(n16738), .A2(n16385), .B1(n16384), .B2(n16736), .ZN(
        n16386) );
  XOR2_X1 U18490 ( .A(n16387), .B(n16386), .Z(n17109) );
  XOR2_X1 U18491 ( .A(P1_REIP_REG_30__SCAN_IN), .B(n16732), .Z(n16391) );
  NAND2_X1 U18492 ( .A1(n22266), .A2(n16904), .ZN(n16389) );
  AOI22_X1 U18493 ( .A1(n22264), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n22236), .ZN(n16388) );
  NAND2_X1 U18494 ( .A1(n16389), .A2(n16388), .ZN(n16390) );
  OAI21_X1 U18495 ( .B1(n16846), .B2(n22269), .A(n16394), .ZN(P1_U2810) );
  INV_X1 U18496 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n16395) );
  OAI222_X1 U18497 ( .A1(n20698), .A2(n16846), .B1(n16395), .B2(n20727), .C1(
        n17109), .C2(n16841), .ZN(P1_U2842) );
  NAND2_X1 U18498 ( .A1(n19350), .A2(n18091), .ZN(n16403) );
  INV_X1 U18499 ( .A(n16396), .ZN(n16401) );
  AOI21_X1 U18500 ( .B1(n18102), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n16397), .ZN(n16398) );
  OAI21_X1 U18501 ( .B1(n18112), .B2(n16399), .A(n16398), .ZN(n16400) );
  OAI21_X1 U18502 ( .B1(n16405), .B2(n18106), .A(n16404), .ZN(P2_U2983) );
  NOR2_X1 U18503 ( .A1(n18112), .A2(n16406), .ZN(n16407) );
  AOI211_X1 U18504 ( .C1(n18102), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n16408), .B(n16407), .ZN(n16409) );
  OAI21_X1 U18505 ( .B1(n16686), .B2(n18105), .A(n16409), .ZN(n16410) );
  OAI21_X1 U18506 ( .B1(n16413), .B2(n18106), .A(n16412), .ZN(P2_U2984) );
  INV_X1 U18507 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n20273) );
  AOI22_X1 U18508 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11944), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16415) );
  AOI22_X1 U18509 ( .A1(n16449), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16448), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16414) );
  OAI211_X1 U18510 ( .C1(n20273), .C2(n16452), .A(n16415), .B(n16414), .ZN(
        n16423) );
  INV_X1 U18511 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16417) );
  INV_X1 U18512 ( .A(n16416), .ZN(n16455) );
  INV_X1 U18513 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16587) );
  OAI22_X1 U18514 ( .A1(n16417), .A2(n16455), .B1(n16454), .B2(n16587), .ZN(
        n16422) );
  INV_X1 U18515 ( .A(n16418), .ZN(n16460) );
  INV_X1 U18516 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16420) );
  INV_X1 U18517 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16419) );
  OAI22_X1 U18518 ( .A1(n16460), .A2(n16420), .B1(n16458), .B2(n16419), .ZN(
        n16421) );
  NOR3_X1 U18519 ( .A1(n16423), .A2(n16422), .A3(n16421), .ZN(n16431) );
  AOI22_X1 U18520 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16481), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16430) );
  AOI22_X1 U18521 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11905), .B1(
        n11978), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16429) );
  INV_X1 U18522 ( .A(n16482), .ZN(n16465) );
  INV_X1 U18523 ( .A(n16424), .ZN(n16464) );
  INV_X1 U18524 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16425) );
  OAI22_X1 U18525 ( .A1(n16426), .A2(n16465), .B1(n16464), .B2(n16425), .ZN(
        n16427) );
  AOI21_X1 U18526 ( .B1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B2(n16217), .A(
        n16427), .ZN(n16428) );
  NAND4_X1 U18527 ( .A1(n16431), .A2(n16430), .A3(n16429), .A4(n16428), .ZN(
        n17422) );
  INV_X1 U18528 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16435) );
  AOI22_X1 U18529 ( .A1(n11978), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11905), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16434) );
  AOI22_X1 U18530 ( .A1(n16482), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16424), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16433) );
  OAI211_X1 U18531 ( .C1(n16436), .C2(n16435), .A(n16434), .B(n16433), .ZN(
        n16447) );
  AOI22_X1 U18532 ( .A1(n12062), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11944), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16438) );
  AOI22_X1 U18533 ( .A1(n16449), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16448), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16437) );
  OAI211_X1 U18534 ( .C1(n16601), .C2(n16452), .A(n16438), .B(n16437), .ZN(
        n16446) );
  AOI22_X1 U18535 ( .A1(n16472), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16416), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16440) );
  AOI22_X1 U18536 ( .A1(n16418), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11939), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16439) );
  NAND2_X1 U18537 ( .A1(n16440), .A2(n16439), .ZN(n16445) );
  INV_X1 U18538 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16442) );
  INV_X1 U18539 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16612) );
  OAI22_X1 U18540 ( .A1(n16443), .A2(n16442), .B1(n16441), .B2(n16612), .ZN(
        n16444) );
  NOR4_X1 U18541 ( .A1(n16447), .A2(n16446), .A3(n16445), .A4(n16444), .ZN(
        n17416) );
  AOI22_X1 U18542 ( .A1(n12062), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11944), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16451) );
  AOI22_X1 U18543 ( .A1(n16449), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16448), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16450) );
  OAI211_X1 U18544 ( .C1(n20162), .C2(n16452), .A(n16451), .B(n16450), .ZN(
        n16463) );
  OAI22_X1 U18545 ( .A1(n16456), .A2(n16455), .B1(n16454), .B2(n16453), .ZN(
        n16462) );
  OAI22_X1 U18546 ( .A1(n16460), .A2(n16459), .B1(n16458), .B2(n16457), .ZN(
        n16461) );
  NOR3_X1 U18547 ( .A1(n16463), .A2(n16462), .A3(n16461), .ZN(n16471) );
  AOI22_X1 U18548 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16481), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16470) );
  AOI22_X1 U18549 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n11978), .B1(
        n11905), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16469) );
  INV_X1 U18550 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16466) );
  OAI22_X1 U18551 ( .A1(n16466), .A2(n16465), .B1(n16464), .B2(n20150), .ZN(
        n16467) );
  AOI21_X1 U18552 ( .B1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B2(n16217), .A(
        n16467), .ZN(n16468) );
  NAND4_X1 U18553 ( .A1(n16471), .A2(n16470), .A3(n16469), .A4(n16468), .ZN(
        n17411) );
  AOI22_X1 U18554 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n16472), .B1(
        n16416), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16480) );
  OAI22_X1 U18555 ( .A1(n16475), .A2(n16474), .B1(n16473), .B2(n16671), .ZN(
        n16476) );
  AOI21_X1 U18556 ( .B1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n12024), .A(
        n16476), .ZN(n16479) );
  AOI22_X1 U18557 ( .A1(n11987), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11944), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16478) );
  AOI22_X1 U18558 ( .A1(n16418), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11939), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16477) );
  NAND4_X1 U18559 ( .A1(n16480), .A2(n16479), .A3(n16478), .A4(n16477), .ZN(
        n16488) );
  AOI22_X1 U18560 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n11978), .B1(
        n11905), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16486) );
  AOI22_X1 U18561 ( .A1(n16226), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n16481), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16485) );
  AOI22_X1 U18562 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n16482), .B1(
        n16424), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16484) );
  NAND2_X1 U18563 ( .A1(n16217), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n16483) );
  NAND4_X1 U18564 ( .A1(n16486), .A2(n16485), .A3(n16484), .A4(n16483), .ZN(
        n16487) );
  OR2_X1 U18565 ( .A1(n16488), .A2(n16487), .ZN(n16513) );
  INV_X1 U18566 ( .A(n16559), .ZN(n16665) );
  AOI22_X1 U18567 ( .A1(n11158), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n16665), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16501) );
  INV_X1 U18568 ( .A(n11848), .ZN(n16673) );
  INV_X1 U18569 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16494) );
  INV_X1 U18570 ( .A(n16489), .ZN(n16491) );
  NAND2_X1 U18571 ( .A1(n16491), .A2(n16490), .ZN(n16669) );
  INV_X1 U18572 ( .A(n11862), .ZN(n16627) );
  INV_X1 U18573 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16492) );
  OR2_X1 U18574 ( .A1(n16627), .A2(n16492), .ZN(n16493) );
  OAI211_X1 U18575 ( .C1(n16673), .C2(n16494), .A(n16669), .B(n16493), .ZN(
        n16495) );
  INV_X1 U18576 ( .A(n16495), .ZN(n16500) );
  AOI22_X1 U18577 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16676), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16499) );
  INV_X1 U18578 ( .A(n11855), .ZN(n16496) );
  AOI22_X1 U18579 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11857), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16498) );
  NAND4_X1 U18580 ( .A1(n16501), .A2(n16500), .A3(n16499), .A4(n16498), .ZN(
        n16511) );
  AOI22_X1 U18581 ( .A1(n11847), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n16665), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16509) );
  INV_X1 U18582 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16504) );
  INV_X1 U18583 ( .A(n16669), .ZN(n16611) );
  INV_X1 U18584 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16502) );
  OR2_X1 U18585 ( .A1(n16627), .A2(n16502), .ZN(n16503) );
  OAI211_X1 U18586 ( .C1(n16673), .C2(n16504), .A(n16611), .B(n16503), .ZN(
        n16505) );
  INV_X1 U18587 ( .A(n16505), .ZN(n16508) );
  AOI22_X1 U18588 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16676), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n16507) );
  AOI22_X1 U18589 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11857), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16506) );
  NAND4_X1 U18590 ( .A1(n16509), .A2(n16508), .A3(n16507), .A4(n16506), .ZN(
        n16510) );
  AND2_X1 U18591 ( .A1(n16511), .A2(n16510), .ZN(n16512) );
  XNOR2_X1 U18592 ( .A(n16513), .B(n16512), .ZN(n17407) );
  NAND2_X1 U18593 ( .A1(n16513), .A2(n16512), .ZN(n16532) );
  INV_X1 U18594 ( .A(n16532), .ZN(n16514) );
  NAND2_X1 U18595 ( .A1(n16597), .A2(n16514), .ZN(n16534) );
  AOI22_X1 U18596 ( .A1(n11184), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11183), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n16521) );
  AOI22_X1 U18597 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n16665), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n16520) );
  AOI22_X1 U18598 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n16676), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16519) );
  NAND2_X1 U18599 ( .A1(n11857), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n16515) );
  OAI211_X1 U18600 ( .C1(n16627), .C2(n16516), .A(n16515), .B(n16669), .ZN(
        n16517) );
  INV_X1 U18601 ( .A(n16517), .ZN(n16518) );
  NAND4_X1 U18602 ( .A1(n16521), .A2(n16520), .A3(n16519), .A4(n16518), .ZN(
        n16531) );
  AOI22_X1 U18603 ( .A1(n11158), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11183), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16529) );
  AOI22_X1 U18604 ( .A1(n16665), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n16676), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n16528) );
  AOI22_X1 U18605 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11857), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16527) );
  INV_X1 U18606 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16524) );
  INV_X1 U18607 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16522) );
  OR2_X1 U18608 ( .A1(n16627), .A2(n16522), .ZN(n16523) );
  OAI211_X1 U18609 ( .C1(n16673), .C2(n16524), .A(n16611), .B(n16523), .ZN(
        n16525) );
  INV_X1 U18610 ( .A(n16525), .ZN(n16526) );
  NAND4_X1 U18611 ( .A1(n16529), .A2(n16528), .A3(n16527), .A4(n16526), .ZN(
        n16530) );
  NAND2_X1 U18612 ( .A1(n16531), .A2(n16530), .ZN(n16533) );
  NOR2_X1 U18613 ( .A1(n16532), .A2(n16533), .ZN(n16552) );
  AOI22_X1 U18614 ( .A1(n16534), .A2(n16533), .B1(n16552), .B2(n19079), .ZN(
        n17399) );
  AOI22_X1 U18615 ( .A1(n11158), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16665), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16541) );
  INV_X1 U18616 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16536) );
  INV_X1 U18617 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20378) );
  OR2_X1 U18618 ( .A1(n16627), .A2(n20378), .ZN(n16535) );
  OAI211_X1 U18619 ( .C1(n16673), .C2(n16536), .A(n16669), .B(n16535), .ZN(
        n16537) );
  INV_X1 U18620 ( .A(n16537), .ZN(n16540) );
  AOI22_X1 U18621 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n16676), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16539) );
  AOI22_X1 U18622 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11857), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n16538) );
  NAND4_X1 U18623 ( .A1(n16541), .A2(n16540), .A3(n16539), .A4(n16538), .ZN(
        n16551) );
  AOI22_X1 U18624 ( .A1(n11158), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n16665), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n16549) );
  INV_X1 U18625 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n16544) );
  INV_X1 U18626 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16542) );
  OR2_X1 U18627 ( .A1(n16627), .A2(n16542), .ZN(n16543) );
  OAI211_X1 U18628 ( .C1(n16673), .C2(n16544), .A(n16611), .B(n16543), .ZN(
        n16545) );
  INV_X1 U18629 ( .A(n16545), .ZN(n16548) );
  AOI22_X1 U18630 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16676), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16547) );
  AOI22_X1 U18631 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11857), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16546) );
  NAND4_X1 U18632 ( .A1(n16549), .A2(n16548), .A3(n16547), .A4(n16546), .ZN(
        n16550) );
  AND2_X1 U18633 ( .A1(n16551), .A2(n16550), .ZN(n16554) );
  NAND2_X1 U18634 ( .A1(n16552), .A2(n16554), .ZN(n16579) );
  OAI211_X1 U18635 ( .C1(n16552), .C2(n16554), .A(n16579), .B(n16597), .ZN(
        n16556) );
  INV_X1 U18636 ( .A(n16556), .ZN(n16553) );
  INV_X1 U18637 ( .A(n16554), .ZN(n16555) );
  NOR2_X1 U18638 ( .A1(n19079), .A2(n16555), .ZN(n17395) );
  NAND2_X1 U18639 ( .A1(n17393), .A2(n17395), .ZN(n17394) );
  AOI22_X1 U18640 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11855), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16564) );
  AOI22_X1 U18641 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16563) );
  AOI22_X1 U18642 ( .A1(n11158), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n16676), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16562) );
  INV_X1 U18643 ( .A(n11639), .ZN(n16559) );
  NAND2_X1 U18644 ( .A1(n11857), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n16557) );
  OAI211_X1 U18645 ( .C1(n16559), .C2(n16558), .A(n16557), .B(n16669), .ZN(
        n16560) );
  INV_X1 U18646 ( .A(n16560), .ZN(n16561) );
  NAND4_X1 U18647 ( .A1(n16564), .A2(n16563), .A3(n16562), .A4(n16561), .ZN(
        n16573) );
  AOI22_X1 U18648 ( .A1(n11158), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16665), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16571) );
  INV_X1 U18649 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16565) );
  OR2_X1 U18650 ( .A1(n16627), .A2(n16565), .ZN(n16566) );
  OAI211_X1 U18651 ( .C1(n16673), .C2(n16227), .A(n16611), .B(n16566), .ZN(
        n16567) );
  INV_X1 U18652 ( .A(n16567), .ZN(n16570) );
  AOI22_X1 U18653 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n16676), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16569) );
  AOI22_X1 U18654 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11857), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16568) );
  NAND4_X1 U18655 ( .A1(n16571), .A2(n16570), .A3(n16569), .A4(n16568), .ZN(
        n16572) );
  AND2_X1 U18656 ( .A1(n16573), .A2(n16572), .ZN(n16577) );
  XNOR2_X1 U18657 ( .A(n16579), .B(n16577), .ZN(n16574) );
  NAND2_X1 U18658 ( .A1(n12188), .A2(n16577), .ZN(n17390) );
  INV_X1 U18659 ( .A(n16577), .ZN(n16578) );
  NOR2_X1 U18660 ( .A1(n16579), .A2(n16578), .ZN(n16598) );
  AOI22_X1 U18661 ( .A1(n11184), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16665), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16586) );
  INV_X1 U18662 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16581) );
  OR2_X1 U18663 ( .A1(n16627), .A2(n20273), .ZN(n16580) );
  OAI211_X1 U18664 ( .C1(n16673), .C2(n16581), .A(n16669), .B(n16580), .ZN(
        n16582) );
  INV_X1 U18665 ( .A(n16582), .ZN(n16585) );
  AOI22_X1 U18666 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16676), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16584) );
  AOI22_X1 U18667 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11857), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16583) );
  NAND4_X1 U18668 ( .A1(n16586), .A2(n16585), .A3(n16584), .A4(n16583), .ZN(
        n16596) );
  AOI22_X1 U18669 ( .A1(n11184), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16665), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16594) );
  INV_X1 U18670 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16589) );
  OR2_X1 U18671 ( .A1(n16627), .A2(n16587), .ZN(n16588) );
  OAI211_X1 U18672 ( .C1(n16673), .C2(n16589), .A(n16611), .B(n16588), .ZN(
        n16590) );
  INV_X1 U18673 ( .A(n16590), .ZN(n16593) );
  AOI22_X1 U18674 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16676), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16592) );
  AOI22_X1 U18675 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11857), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16591) );
  NAND4_X1 U18676 ( .A1(n16594), .A2(n16593), .A3(n16592), .A4(n16591), .ZN(
        n16595) );
  AND2_X1 U18677 ( .A1(n16596), .A2(n16595), .ZN(n16599) );
  NAND2_X1 U18678 ( .A1(n16598), .A2(n16599), .ZN(n17374) );
  INV_X1 U18679 ( .A(n16599), .ZN(n16600) );
  NOR2_X1 U18680 ( .A1(n19079), .A2(n16600), .ZN(n17382) );
  AOI22_X1 U18681 ( .A1(n11184), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n16665), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16608) );
  INV_X1 U18682 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16603) );
  OR2_X1 U18683 ( .A1(n16627), .A2(n16601), .ZN(n16602) );
  OAI211_X1 U18684 ( .C1(n16673), .C2(n16603), .A(n16669), .B(n16602), .ZN(
        n16604) );
  INV_X1 U18685 ( .A(n16604), .ZN(n16607) );
  AOI22_X1 U18686 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16676), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16606) );
  AOI22_X1 U18687 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11857), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16605) );
  NAND4_X1 U18688 ( .A1(n16608), .A2(n16607), .A3(n16606), .A4(n16605), .ZN(
        n16619) );
  AOI22_X1 U18689 ( .A1(n11184), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16665), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16617) );
  INV_X1 U18690 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16609) );
  OR2_X1 U18691 ( .A1(n16627), .A2(n16609), .ZN(n16610) );
  OAI211_X1 U18692 ( .C1(n16673), .C2(n16612), .A(n16611), .B(n16610), .ZN(
        n16613) );
  INV_X1 U18693 ( .A(n16613), .ZN(n16616) );
  AOI22_X1 U18694 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16676), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16615) );
  AOI22_X1 U18695 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11857), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16614) );
  NAND4_X1 U18696 ( .A1(n16617), .A2(n16616), .A3(n16615), .A4(n16614), .ZN(
        n16618) );
  AND2_X1 U18697 ( .A1(n16619), .A2(n16618), .ZN(n17375) );
  NAND2_X1 U18698 ( .A1(n16621), .A2(n16620), .ZN(n17379) );
  OAI211_X1 U18699 ( .C1(n17373), .C2(n17382), .A(n17375), .B(n17379), .ZN(
        n16639) );
  AOI22_X1 U18700 ( .A1(n11184), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11183), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16623) );
  AOI22_X1 U18701 ( .A1(n16665), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11857), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16622) );
  NAND2_X1 U18702 ( .A1(n16623), .A2(n16622), .ZN(n16637) );
  AOI22_X1 U18703 ( .A1(n11855), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n16676), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16625) );
  AOI21_X1 U18704 ( .B1(n11862), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n16669), .ZN(n16624) );
  OAI211_X1 U18705 ( .C1(n16673), .C2(n16626), .A(n16625), .B(n16624), .ZN(
        n16636) );
  OAI21_X1 U18706 ( .B1(n16627), .B2(n20162), .A(n16669), .ZN(n16631) );
  INV_X1 U18707 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16629) );
  INV_X1 U18708 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16628) );
  OAI22_X1 U18709 ( .A1(n16496), .A2(n16629), .B1(n16497), .B2(n16628), .ZN(
        n16630) );
  AOI211_X1 U18710 ( .C1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .C2(n16676), .A(
        n16631), .B(n16630), .ZN(n16634) );
  AOI22_X1 U18711 ( .A1(n11184), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16665), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16633) );
  AOI22_X1 U18712 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11848), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16632) );
  NAND3_X1 U18713 ( .A1(n16634), .A2(n16633), .A3(n16632), .ZN(n16635) );
  OAI21_X1 U18714 ( .B1(n16637), .B2(n16636), .A(n16635), .ZN(n16638) );
  NAND2_X1 U18715 ( .A1(n16639), .A2(n16638), .ZN(n16660) );
  INV_X1 U18716 ( .A(n16660), .ZN(n16640) );
  NOR2_X1 U18717 ( .A1(n16639), .A2(n16638), .ZN(n16658) );
  NOR2_X1 U18718 ( .A1(n16640), .A2(n16658), .ZN(n16642) );
  INV_X1 U18719 ( .A(n17375), .ZN(n16641) );
  XNOR2_X1 U18720 ( .A(n16642), .B(n16659), .ZN(n16657) );
  NAND2_X1 U18721 ( .A1(n17423), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16647) );
  NAND2_X1 U18722 ( .A1(n19331), .A2(n14580), .ZN(n16646) );
  OAI211_X1 U18723 ( .C1(n16657), .C2(n17428), .A(n16647), .B(n16646), .ZN(
        P2_U2858) );
  NOR2_X1 U18724 ( .A1(n16649), .A2(n16648), .ZN(n16650) );
  OAI22_X1 U18725 ( .A1(n17477), .A2(n19337), .B1(n17475), .B2(n16652), .ZN(
        n16653) );
  AOI21_X1 U18726 ( .B1(n17479), .B2(n16654), .A(n16653), .ZN(n16656) );
  AOI22_X1 U18727 ( .A1(n19914), .A2(BUF2_REG_29__SCAN_IN), .B1(n19915), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n16655) );
  OAI211_X1 U18728 ( .C1(n16657), .C2(n20165), .A(n16656), .B(n16655), .ZN(
        P2_U2890) );
  INV_X1 U18729 ( .A(n16658), .ZN(n16662) );
  NAND2_X1 U18730 ( .A1(n16662), .A2(n16661), .ZN(n16685) );
  AOI22_X1 U18731 ( .A1(n11848), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16664) );
  AOI22_X1 U18732 ( .A1(n11184), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16676), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16663) );
  NAND2_X1 U18733 ( .A1(n16664), .A2(n16663), .ZN(n16682) );
  INV_X1 U18734 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16668) );
  AOI22_X1 U18735 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11855), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16667) );
  AOI21_X1 U18736 ( .B1(n16665), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n16669), .ZN(n16666) );
  OAI211_X1 U18737 ( .C1(n16497), .C2(n16668), .A(n16667), .B(n16666), .ZN(
        n16681) );
  OAI21_X1 U18738 ( .B1(n16559), .B2(n16670), .A(n16669), .ZN(n16675) );
  INV_X1 U18739 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16672) );
  OAI22_X1 U18740 ( .A1(n16673), .A2(n16672), .B1(n16496), .B2(n16671), .ZN(
        n16674) );
  AOI211_X1 U18741 ( .C1(n16676), .C2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n16675), .B(n16674), .ZN(n16679) );
  AOI22_X1 U18742 ( .A1(n11183), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16678) );
  AOI22_X1 U18743 ( .A1(n11184), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11857), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16677) );
  NAND3_X1 U18744 ( .A1(n16679), .A2(n16678), .A3(n16677), .ZN(n16680) );
  OAI21_X1 U18745 ( .B1(n16682), .B2(n16681), .A(n16680), .ZN(n16683) );
  INV_X1 U18746 ( .A(n16683), .ZN(n16684) );
  XNOR2_X1 U18747 ( .A(n16685), .B(n16684), .ZN(n16694) );
  NOR2_X1 U18748 ( .A1(n16686), .A2(n17423), .ZN(n16687) );
  AOI21_X1 U18749 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n17420), .A(n16687), .ZN(
        n16688) );
  OAI21_X1 U18750 ( .B1(n16694), .B2(n17428), .A(n16688), .ZN(P2_U2857) );
  OAI22_X1 U18751 ( .A1(n12800), .A2(n17477), .B1(n17475), .B2(n16689), .ZN(
        n16690) );
  AOI21_X1 U18752 ( .B1(n17479), .B2(n16691), .A(n16690), .ZN(n16693) );
  AOI22_X1 U18753 ( .A1(n19914), .A2(BUF2_REG_30__SCAN_IN), .B1(n19915), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n16692) );
  NAND2_X1 U18754 ( .A1(n16696), .A2(n16695), .ZN(n16698) );
  XOR2_X1 U18755 ( .A(n16698), .B(n16697), .Z(n17659) );
  INV_X1 U18756 ( .A(n17493), .ZN(n16701) );
  OAI21_X1 U18757 ( .B1(n16701), .B2(n16700), .A(n16699), .ZN(n16703) );
  NAND2_X1 U18758 ( .A1(n18070), .A2(n19329), .ZN(n16704) );
  NAND2_X1 U18759 ( .A1(n19407), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n17647) );
  OAI211_X1 U18760 ( .C1(n18076), .C2(n16705), .A(n16704), .B(n17647), .ZN(
        n16706) );
  OAI21_X1 U18761 ( .B1(n17659), .B2(n18106), .A(n16708), .ZN(P2_U2985) );
  INV_X1 U18762 ( .A(n16709), .ZN(n16718) );
  NAND3_X1 U18763 ( .A1(n16711), .A2(n12933), .A3(n16710), .ZN(n16712) );
  NAND2_X1 U18764 ( .A1(n16713), .A2(n16712), .ZN(n16714) );
  NAND2_X1 U18765 ( .A1(n16719), .A2(n16714), .ZN(n16717) );
  NAND2_X1 U18766 ( .A1(n16722), .A2(n16715), .ZN(n16716) );
  OAI211_X1 U18767 ( .C1(n16719), .C2(n16718), .A(n16717), .B(n16716), .ZN(
        n16720) );
  NAND2_X1 U18768 ( .A1(n16720), .A2(n12941), .ZN(n18009) );
  INV_X1 U18769 ( .A(n18009), .ZN(n16728) );
  INV_X1 U18770 ( .A(n13689), .ZN(n16723) );
  AND2_X1 U18771 ( .A1(n16722), .A2(n16721), .ZN(n22808) );
  OAI22_X1 U18772 ( .A1(n16725), .A2(n16724), .B1(n16723), .B2(n22808), .ZN(
        n20766) );
  INV_X1 U18773 ( .A(n16726), .ZN(n16727) );
  AOI21_X1 U18774 ( .B1(n16727), .B2(n22331), .A(n22330), .ZN(n21970) );
  NOR2_X1 U18775 ( .A1(n20766), .A2(n21970), .ZN(n18016) );
  NOR2_X1 U18776 ( .A1(n18016), .A2(n22302), .ZN(n22279) );
  MUX2_X1 U18777 ( .A(P1_MORE_REG_SCAN_IN), .B(n16728), .S(n22279), .Z(
        P1_U3484) );
  INV_X1 U18778 ( .A(n16729), .ZN(n16730) );
  AOI21_X1 U18779 ( .B1(n16731), .B2(n16265), .A(n16730), .ZN(n16916) );
  INV_X1 U18780 ( .A(n16916), .ZN(n16850) );
  INV_X1 U18781 ( .A(n16732), .ZN(n16742) );
  OAI21_X1 U18782 ( .B1(n22200), .B2(n16912), .A(n16733), .ZN(n16741) );
  AOI22_X1 U18783 ( .A1(n22264), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B1(
        n22236), .B2(P1_EBX_REG_29__SCAN_IN), .ZN(n16734) );
  OAI21_X1 U18784 ( .B1(n22257), .B2(n16914), .A(n16734), .ZN(n16740) );
  AND2_X1 U18785 ( .A1(n16736), .A2(n16735), .ZN(n16737) );
  NOR2_X1 U18786 ( .A1(n17126), .A2(n22276), .ZN(n16739) );
  AOI211_X1 U18787 ( .C1(n16742), .C2(n16741), .A(n16740), .B(n16739), .ZN(
        n16743) );
  OAI21_X1 U18788 ( .B1(n16850), .B2(n22269), .A(n16743), .ZN(P1_U2811) );
  AOI21_X1 U18789 ( .B1(n16745), .B2(n16757), .A(n16263), .ZN(n16938) );
  INV_X1 U18790 ( .A(n16938), .ZN(n16854) );
  OAI21_X1 U18791 ( .B1(n22200), .B2(n16934), .A(n16762), .ZN(n16753) );
  INV_X1 U18792 ( .A(n16746), .ZN(n16748) );
  AOI21_X1 U18793 ( .B1(n16749), .B2(n16748), .A(n16747), .ZN(n17148) );
  NAND2_X1 U18794 ( .A1(n17148), .A2(n22217), .ZN(n16751) );
  AOI22_X1 U18795 ( .A1(n22264), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(
        n22236), .B2(P1_EBX_REG_27__SCAN_IN), .ZN(n16750) );
  OAI211_X1 U18796 ( .C1(n22257), .C2(n16936), .A(n16751), .B(n16750), .ZN(
        n16752) );
  AOI21_X1 U18797 ( .B1(n16754), .B2(n16753), .A(n16752), .ZN(n16755) );
  OAI21_X1 U18798 ( .B1(n16854), .B2(n22269), .A(n16755), .ZN(P1_U2813) );
  OAI21_X1 U18799 ( .B1(n16756), .B2(n16758), .A(n16757), .ZN(n16947) );
  AOI21_X1 U18800 ( .B1(n16759), .B2(n11200), .A(n16746), .ZN(n17151) );
  INV_X1 U18801 ( .A(n16944), .ZN(n16761) );
  AOI22_X1 U18802 ( .A1(n22264), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n22236), .B2(P1_EBX_REG_26__SCAN_IN), .ZN(n16760) );
  OAI21_X1 U18803 ( .B1(n22257), .B2(n16761), .A(n16760), .ZN(n16766) );
  AOI21_X1 U18804 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(n22210), .A(n16774), 
        .ZN(n16764) );
  INV_X1 U18805 ( .A(n16762), .ZN(n16763) );
  NOR2_X1 U18806 ( .A1(n16764), .A2(n16763), .ZN(n16765) );
  AOI211_X1 U18807 ( .C1(n17151), .C2(n22217), .A(n16766), .B(n16765), .ZN(
        n16767) );
  OAI21_X1 U18808 ( .B1(n16947), .B2(n22269), .A(n16767), .ZN(P1_U2814) );
  INV_X1 U18809 ( .A(n16768), .ZN(n16769) );
  AOI21_X1 U18810 ( .B1(n16769), .B2(n11198), .A(n16756), .ZN(n16956) );
  INV_X1 U18811 ( .A(n16956), .ZN(n16861) );
  NAND2_X1 U18812 ( .A1(n16770), .A2(n16771), .ZN(n16772) );
  AND2_X1 U18813 ( .A1(n11200), .A2(n16772), .ZN(n17168) );
  AOI22_X1 U18814 ( .A1(n22264), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n22236), .B2(P1_EBX_REG_25__SCAN_IN), .ZN(n16773) );
  OAI21_X1 U18815 ( .B1(n22257), .B2(n16954), .A(n16773), .ZN(n16778) );
  NAND2_X1 U18816 ( .A1(n22210), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n16775) );
  AOI21_X1 U18817 ( .B1(n16776), .B2(n16775), .A(n16774), .ZN(n16777) );
  AOI211_X1 U18818 ( .C1(n17168), .C2(n22217), .A(n16778), .B(n16777), .ZN(
        n16779) );
  OAI21_X1 U18819 ( .B1(n16861), .B2(n22269), .A(n16779), .ZN(P1_U2815) );
  NAND2_X1 U18820 ( .A1(n16797), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n16787) );
  INV_X1 U18821 ( .A(n16787), .ZN(n16781) );
  NOR2_X1 U18822 ( .A1(n16781), .A2(n22200), .ZN(n16796) );
  INV_X1 U18823 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n16820) );
  NAND2_X1 U18824 ( .A1(n22264), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16782) );
  OAI21_X1 U18825 ( .B1(n16820), .B2(n22262), .A(n16782), .ZN(n16785) );
  OAI21_X1 U18826 ( .B1(n16792), .B2(n16783), .A(n16770), .ZN(n17175) );
  NOR2_X1 U18827 ( .A1(n17175), .A2(n22276), .ZN(n16784) );
  AOI211_X1 U18828 ( .C1(n22266), .C2(n16966), .A(n16785), .B(n16784), .ZN(
        n16786) );
  OAI21_X1 U18829 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n16787), .A(n16786), 
        .ZN(n16788) );
  AOI21_X1 U18830 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n16796), .A(n16788), 
        .ZN(n16789) );
  OAI21_X1 U18831 ( .B1(n16963), .B2(n22269), .A(n16789), .ZN(P1_U2816) );
  AOI21_X1 U18832 ( .B1(n16791), .B2(n16790), .A(n16780), .ZN(n16973) );
  INV_X1 U18833 ( .A(n16973), .ZN(n16868) );
  AOI21_X1 U18834 ( .B1(n16793), .B2(n16825), .A(n16792), .ZN(n17187) );
  AOI22_X1 U18835 ( .A1(n22264), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n22236), .B2(P1_EBX_REG_23__SCAN_IN), .ZN(n16794) );
  OAI21_X1 U18836 ( .B1(n22257), .B2(n16971), .A(n16794), .ZN(n16795) );
  AOI21_X1 U18837 ( .B1(n17187), .B2(n22217), .A(n16795), .ZN(n16799) );
  OAI21_X1 U18838 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(n16797), .A(n16796), 
        .ZN(n16798) );
  OAI211_X1 U18839 ( .C1(n16868), .C2(n22269), .A(n16799), .B(n16798), .ZN(
        P1_U2817) );
  NAND2_X1 U18840 ( .A1(n16800), .A2(n16801), .ZN(n16802) );
  AND2_X1 U18841 ( .A1(n11211), .A2(n16802), .ZN(n20712) );
  INV_X1 U18842 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n22199) );
  NAND2_X1 U18843 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n22182), .ZN(n22198) );
  NOR2_X1 U18844 ( .A1(n22199), .A2(n22198), .ZN(n22209) );
  NAND2_X1 U18845 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n22209), .ZN(n22233) );
  INV_X1 U18846 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n22232) );
  NOR2_X1 U18847 ( .A1(n22233), .A2(n22232), .ZN(n16804) );
  AOI21_X1 U18848 ( .B1(n16804), .B2(P1_REIP_REG_19__SCAN_IN), .A(n22200), 
        .ZN(n16803) );
  OAI21_X1 U18849 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(n16804), .A(n16803), 
        .ZN(n16810) );
  AND2_X1 U18850 ( .A1(n16839), .A2(n16805), .ZN(n16806) );
  NOR2_X1 U18851 ( .A1(n16830), .A2(n16806), .ZN(n20711) );
  INV_X1 U18852 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n20714) );
  AOI21_X1 U18853 ( .B1(n22264), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n22223), .ZN(n16807) );
  OAI21_X1 U18854 ( .B1(n22262), .B2(n20714), .A(n16807), .ZN(n16808) );
  AOI21_X1 U18855 ( .B1(n20711), .B2(n22217), .A(n16808), .ZN(n16809) );
  OAI211_X1 U18856 ( .C1(n17000), .C2(n22257), .A(n16810), .B(n16809), .ZN(
        n16811) );
  AOI21_X1 U18857 ( .B1(n20712), .B2(n22253), .A(n16811), .ZN(n16812) );
  INV_X1 U18858 ( .A(n16812), .ZN(P1_U2821) );
  INV_X1 U18859 ( .A(n17106), .ZN(n16814) );
  OAI22_X1 U18860 ( .A1(n16814), .A2(n16841), .B1(n20727), .B2(n16813), .ZN(
        P1_U2841) );
  OAI222_X1 U18861 ( .A1(n20698), .A2(n16850), .B1(n16815), .B2(n20727), .C1(
        n17126), .C2(n16841), .ZN(P1_U2843) );
  INV_X1 U18862 ( .A(n17148), .ZN(n16816) );
  OAI222_X1 U18863 ( .A1(n20698), .A2(n16854), .B1(n16817), .B2(n20727), .C1(
        n16816), .C2(n16841), .ZN(P1_U2845) );
  AOI22_X1 U18864 ( .A1(n17151), .A2(n20724), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n16821), .ZN(n16818) );
  OAI21_X1 U18865 ( .B1(n16947), .B2(n20698), .A(n16818), .ZN(P1_U2846) );
  AOI22_X1 U18866 ( .A1(n17168), .A2(n20724), .B1(P1_EBX_REG_25__SCAN_IN), 
        .B2(n16821), .ZN(n16819) );
  OAI21_X1 U18867 ( .B1(n16861), .B2(n20698), .A(n16819), .ZN(P1_U2847) );
  OAI222_X1 U18868 ( .A1(n16963), .A2(n20698), .B1(n16820), .B2(n20727), .C1(
        n17175), .C2(n16841), .ZN(P1_U2848) );
  AOI22_X1 U18869 ( .A1(n17187), .A2(n20724), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n16821), .ZN(n16822) );
  OAI21_X1 U18870 ( .B1(n16868), .B2(n20698), .A(n16822), .ZN(P1_U2849) );
  OAI21_X1 U18871 ( .B1(n16823), .B2(n16824), .A(n16790), .ZN(n22270) );
  OAI21_X1 U18872 ( .B1(n11370), .B2(n11241), .A(n16825), .ZN(n22275) );
  OAI222_X1 U18873 ( .A1(n22270), .A2(n20698), .B1(n22261), .B2(n20727), .C1(
        n22275), .C2(n16841), .ZN(P1_U2850) );
  INV_X1 U18874 ( .A(n16826), .ZN(n16827) );
  AOI21_X1 U18875 ( .B1(n16828), .B2(n11211), .A(n16827), .ZN(n16995) );
  INV_X1 U18876 ( .A(n16995), .ZN(n22238) );
  INV_X1 U18877 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n16832) );
  OR2_X1 U18878 ( .A1(n16830), .A2(n16829), .ZN(n16831) );
  AND2_X1 U18879 ( .A1(n17210), .A2(n16831), .ZN(n17226) );
  INV_X1 U18880 ( .A(n17226), .ZN(n22237) );
  OAI222_X1 U18881 ( .A1(n20698), .A2(n22238), .B1(n16832), .B2(n20727), .C1(
        n22237), .C2(n16841), .ZN(P1_U2852) );
  OR2_X1 U18883 ( .A1(n16834), .A2(n16835), .ZN(n16836) );
  AND2_X1 U18884 ( .A1(n16800), .A2(n16836), .ZN(n22229) );
  INV_X1 U18885 ( .A(n22229), .ZN(n16888) );
  INV_X1 U18886 ( .A(n16837), .ZN(n17258) );
  INV_X1 U18887 ( .A(n16838), .ZN(n16840) );
  OAI21_X1 U18888 ( .B1(n17258), .B2(n16840), .A(n16839), .ZN(n22226) );
  OAI222_X1 U18889 ( .A1(n16888), .A2(n20698), .B1(n16842), .B2(n20727), .C1(
        n22226), .C2(n16841), .ZN(P1_U2854) );
  AOI22_X1 U18890 ( .A1(n16891), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n16890), .ZN(n16845) );
  AOI22_X1 U18891 ( .A1(n16894), .A2(n16843), .B1(n16892), .B2(DATAI_30_), 
        .ZN(n16844) );
  OAI211_X1 U18892 ( .C1(n16846), .C2(n16897), .A(n16845), .B(n16844), .ZN(
        P1_U2874) );
  AOI22_X1 U18893 ( .A1(n16891), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n16890), .ZN(n16849) );
  AOI22_X1 U18894 ( .A1(n16894), .A2(n16847), .B1(n16892), .B2(DATAI_29_), 
        .ZN(n16848) );
  OAI211_X1 U18895 ( .C1(n16850), .C2(n16897), .A(n16849), .B(n16848), .ZN(
        P1_U2875) );
  AOI22_X1 U18896 ( .A1(n16891), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n16890), .ZN(n16853) );
  AOI22_X1 U18897 ( .A1(n16894), .A2(n16851), .B1(n16892), .B2(DATAI_27_), 
        .ZN(n16852) );
  OAI211_X1 U18898 ( .C1(n16854), .C2(n16897), .A(n16853), .B(n16852), .ZN(
        P1_U2877) );
  AOI22_X1 U18899 ( .A1(n16891), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n16890), .ZN(n16857) );
  AOI22_X1 U18900 ( .A1(n16894), .A2(n16855), .B1(n16892), .B2(DATAI_26_), 
        .ZN(n16856) );
  OAI211_X1 U18901 ( .C1(n16947), .C2(n16897), .A(n16857), .B(n16856), .ZN(
        P1_U2878) );
  AOI22_X1 U18902 ( .A1(n16891), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n16890), .ZN(n16860) );
  AOI22_X1 U18903 ( .A1(n16894), .A2(n16858), .B1(n16892), .B2(DATAI_25_), 
        .ZN(n16859) );
  OAI211_X1 U18904 ( .C1(n16861), .C2(n16897), .A(n16860), .B(n16859), .ZN(
        P1_U2879) );
  AOI22_X1 U18905 ( .A1(n16891), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n16890), .ZN(n16864) );
  AOI22_X1 U18906 ( .A1(n16894), .A2(n16862), .B1(n16892), .B2(DATAI_24_), 
        .ZN(n16863) );
  OAI211_X1 U18907 ( .C1(n16963), .C2(n16897), .A(n16864), .B(n16863), .ZN(
        P1_U2880) );
  AOI22_X1 U18908 ( .A1(n16891), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n16890), .ZN(n16867) );
  AOI22_X1 U18909 ( .A1(n16894), .A2(n16865), .B1(n16892), .B2(DATAI_23_), 
        .ZN(n16866) );
  OAI211_X1 U18910 ( .C1(n16868), .C2(n16897), .A(n16867), .B(n16866), .ZN(
        P1_U2881) );
  AOI22_X1 U18911 ( .A1(n16891), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n16890), .ZN(n16871) );
  AOI22_X1 U18912 ( .A1(n16894), .A2(n16869), .B1(n16892), .B2(DATAI_22_), 
        .ZN(n16870) );
  OAI211_X1 U18913 ( .C1(n22270), .C2(n16897), .A(n16871), .B(n16870), .ZN(
        P1_U2882) );
  AND2_X1 U18914 ( .A1(n16826), .A2(n16872), .ZN(n16873) );
  NOR2_X1 U18915 ( .A1(n16823), .A2(n16873), .ZN(n22254) );
  INV_X1 U18916 ( .A(n22254), .ZN(n16877) );
  AOI22_X1 U18917 ( .A1(n16891), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n16890), .ZN(n16876) );
  AOI22_X1 U18918 ( .A1(n16894), .A2(n16874), .B1(n16892), .B2(DATAI_21_), 
        .ZN(n16875) );
  OAI211_X1 U18919 ( .C1(n16877), .C2(n16897), .A(n16876), .B(n16875), .ZN(
        P1_U2883) );
  AOI22_X1 U18920 ( .A1(n16891), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n16890), .ZN(n16880) );
  AOI22_X1 U18921 ( .A1(n16894), .A2(n16878), .B1(n16892), .B2(DATAI_20_), 
        .ZN(n16879) );
  OAI211_X1 U18922 ( .C1(n22238), .C2(n16897), .A(n16880), .B(n16879), .ZN(
        P1_U2884) );
  INV_X1 U18923 ( .A(n20712), .ZN(n16884) );
  AOI22_X1 U18924 ( .A1(n16891), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n16890), .ZN(n16883) );
  AOI22_X1 U18925 ( .A1(n16894), .A2(n16881), .B1(n16892), .B2(DATAI_19_), 
        .ZN(n16882) );
  OAI211_X1 U18926 ( .C1(n16884), .C2(n16897), .A(n16883), .B(n16882), .ZN(
        P1_U2885) );
  AOI22_X1 U18927 ( .A1(n16891), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n16890), .ZN(n16887) );
  AOI22_X1 U18928 ( .A1(n16894), .A2(n16885), .B1(n16892), .B2(DATAI_18_), 
        .ZN(n16886) );
  OAI211_X1 U18929 ( .C1(n16888), .C2(n16897), .A(n16887), .B(n16886), .ZN(
        P1_U2886) );
  AOI21_X1 U18930 ( .B1(n13339), .B2(n16146), .A(n16834), .ZN(n22218) );
  INV_X1 U18931 ( .A(n22218), .ZN(n16898) );
  AOI22_X1 U18932 ( .A1(n16891), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n16890), .ZN(n16896) );
  AOI22_X1 U18933 ( .A1(n16894), .A2(n16893), .B1(n16892), .B2(DATAI_17_), 
        .ZN(n16895) );
  OAI211_X1 U18934 ( .C1(n16898), .C2(n16897), .A(n16896), .B(n16895), .ZN(
        P1_U2887) );
  INV_X1 U18935 ( .A(n16900), .ZN(n16901) );
  XNOR2_X1 U18936 ( .A(n17256), .B(n17099), .ZN(n16911) );
  XNOR2_X1 U18937 ( .A(n11520), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17121) );
  NAND2_X1 U18938 ( .A1(n16904), .A2(n20761), .ZN(n16905) );
  NAND2_X1 U18939 ( .A1(n22021), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n17116) );
  OAI211_X1 U18940 ( .C1(n20728), .C2(n16906), .A(n16905), .B(n17116), .ZN(
        n16907) );
  AOI21_X1 U18941 ( .B1(n16908), .B2(n20762), .A(n16907), .ZN(n16909) );
  OAI21_X1 U18942 ( .B1(n17121), .B2(n22277), .A(n16909), .ZN(P1_U2969) );
  XNOR2_X1 U18943 ( .A(n16910), .B(n16911), .ZN(n17130) );
  NOR2_X1 U18944 ( .A1(n22066), .A2(n16912), .ZN(n17124) );
  AOI21_X1 U18945 ( .B1(n20760), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n17124), .ZN(n16913) );
  OAI21_X1 U18946 ( .B1(n16914), .B2(n20759), .A(n16913), .ZN(n16915) );
  AOI21_X1 U18947 ( .B1(n16916), .B2(n20762), .A(n16915), .ZN(n16917) );
  OAI21_X1 U18948 ( .B1(n22277), .B2(n17130), .A(n16917), .ZN(P1_U2970) );
  INV_X1 U18949 ( .A(n16918), .ZN(n16958) );
  NAND2_X1 U18950 ( .A1(n16958), .A2(n16919), .ZN(n16924) );
  INV_X1 U18951 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17145) );
  NAND2_X1 U18952 ( .A1(n16920), .A2(n17145), .ZN(n16921) );
  MUX2_X1 U18953 ( .A(n16921), .B(n17097), .S(n17256), .Z(n16923) );
  NOR2_X1 U18954 ( .A1(n16924), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16922) );
  AOI211_X1 U18955 ( .C1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n16924), .A(
        n16923), .B(n16922), .ZN(n16925) );
  XNOR2_X1 U18956 ( .A(n16925), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17140) );
  INV_X1 U18957 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16926) );
  NAND2_X1 U18958 ( .A1(n22021), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n17131) );
  OAI21_X1 U18959 ( .B1(n20728), .B2(n16926), .A(n17131), .ZN(n16929) );
  NOR2_X1 U18960 ( .A1(n16927), .A2(n17060), .ZN(n16928) );
  OAI21_X1 U18961 ( .B1(n22277), .B2(n17140), .A(n16931), .ZN(P1_U2971) );
  XNOR2_X1 U18962 ( .A(n17256), .B(n17145), .ZN(n16932) );
  XNOR2_X1 U18963 ( .A(n16933), .B(n16932), .ZN(n17150) );
  NOR2_X1 U18964 ( .A1(n22066), .A2(n16934), .ZN(n17142) );
  AOI21_X1 U18965 ( .B1(n20760), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n17142), .ZN(n16935) );
  OAI21_X1 U18966 ( .B1(n16936), .B2(n20759), .A(n16935), .ZN(n16937) );
  AOI21_X1 U18967 ( .B1(n16938), .B2(n20762), .A(n16937), .ZN(n16939) );
  OAI21_X1 U18968 ( .B1(n17150), .B2(n22277), .A(n16939), .ZN(P1_U2972) );
  INV_X1 U18969 ( .A(n16940), .ZN(n17153) );
  NAND2_X1 U18970 ( .A1(n16941), .A2(n17097), .ZN(n17152) );
  NAND3_X1 U18971 ( .A1(n17153), .A2(n20756), .A3(n17152), .ZN(n16946) );
  INV_X1 U18972 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16942) );
  NAND2_X1 U18973 ( .A1(n22021), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n17154) );
  OAI21_X1 U18974 ( .B1(n20728), .B2(n16942), .A(n17154), .ZN(n16943) );
  AOI21_X1 U18975 ( .B1(n16944), .B2(n20761), .A(n16943), .ZN(n16945) );
  OAI211_X1 U18976 ( .C1(n17060), .C2(n16947), .A(n16946), .B(n16945), .ZN(
        P1_U2973) );
  NOR2_X1 U18977 ( .A1(n17172), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16950) );
  MUX2_X1 U18978 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n16948), .S(
        n17256), .Z(n16949) );
  AOI211_X1 U18979 ( .C1(n17172), .C2(n16958), .A(n16950), .B(n16949), .ZN(
        n16951) );
  XNOR2_X1 U18980 ( .A(n16951), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17170) );
  NOR2_X1 U18981 ( .A1(n22066), .A2(n16952), .ZN(n17167) );
  AOI21_X1 U18982 ( .B1(n20760), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n17167), .ZN(n16953) );
  OAI21_X1 U18983 ( .B1(n16954), .B2(n20759), .A(n16953), .ZN(n16955) );
  AOI21_X1 U18984 ( .B1(n16956), .B2(n20762), .A(n16955), .ZN(n16957) );
  OAI21_X1 U18985 ( .B1(n17170), .B2(n22277), .A(n16957), .ZN(P1_U2974) );
  NAND3_X1 U18986 ( .A1(n16958), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n17256), .ZN(n16960) );
  INV_X1 U18987 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17184) );
  NAND3_X1 U18988 ( .A1(n16918), .A2(n11541), .A3(n17184), .ZN(n16959) );
  NAND2_X1 U18989 ( .A1(n16960), .A2(n16959), .ZN(n16961) );
  XNOR2_X1 U18990 ( .A(n16961), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17180) );
  NAND2_X1 U18991 ( .A1(n22021), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n17173) );
  OAI21_X1 U18992 ( .B1(n20728), .B2(n16962), .A(n17173), .ZN(n16965) );
  NOR2_X1 U18993 ( .A1(n16963), .A2(n17060), .ZN(n16964) );
  AOI211_X1 U18994 ( .C1(n20761), .C2(n16966), .A(n16965), .B(n16964), .ZN(
        n16967) );
  OAI21_X1 U18995 ( .B1(n17180), .B2(n22277), .A(n16967), .ZN(P1_U2975) );
  XNOR2_X1 U18996 ( .A(n17256), .B(n17184), .ZN(n16968) );
  XNOR2_X1 U18997 ( .A(n16918), .B(n16968), .ZN(n17189) );
  INV_X1 U18998 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n16969) );
  NOR2_X1 U18999 ( .A1(n22066), .A2(n16969), .ZN(n17181) );
  AOI21_X1 U19000 ( .B1(n20760), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n17181), .ZN(n16970) );
  OAI21_X1 U19001 ( .B1(n16971), .B2(n20759), .A(n16970), .ZN(n16972) );
  AOI21_X1 U19002 ( .B1(n16973), .B2(n20762), .A(n16972), .ZN(n16974) );
  OAI21_X1 U19003 ( .B1(n17189), .B2(n22277), .A(n16974), .ZN(P1_U2976) );
  NOR2_X1 U19004 ( .A1(n16976), .A2(n16975), .ZN(n16977) );
  XNOR2_X1 U19005 ( .A(n16977), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17205) );
  NAND2_X1 U19006 ( .A1(n22021), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n17200) );
  OAI21_X1 U19007 ( .B1(n20728), .B2(n16978), .A(n17200), .ZN(n16980) );
  NOR2_X1 U19008 ( .A1(n22270), .A2(n17060), .ZN(n16979) );
  AOI211_X1 U19009 ( .C1(n20761), .C2(n22265), .A(n16980), .B(n16979), .ZN(
        n16981) );
  OAI21_X1 U19010 ( .B1(n22277), .B2(n17205), .A(n16981), .ZN(P1_U2977) );
  XNOR2_X1 U19011 ( .A(n17256), .B(n17244), .ZN(n17003) );
  OR2_X1 U19012 ( .A1(n11165), .A2(n17003), .ZN(n16983) );
  OR2_X1 U19013 ( .A1(n17256), .A2(n17244), .ZN(n16982) );
  MUX2_X1 U19014 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n16998), .S(
        n11541), .Z(n16989) );
  INV_X1 U19015 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17220) );
  INV_X1 U19016 ( .A(n16998), .ZN(n16990) );
  MUX2_X1 U19017 ( .A(n17220), .B(n16990), .S(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(n16984) );
  NAND2_X1 U19018 ( .A1(n16989), .A2(n16984), .ZN(n16985) );
  XOR2_X1 U19019 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n16985), .Z(
        n17216) );
  INV_X1 U19020 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n22247) );
  NOR2_X1 U19021 ( .A1(n22066), .A2(n22247), .ZN(n17207) );
  AOI21_X1 U19022 ( .B1(n20760), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n17207), .ZN(n16986) );
  OAI21_X1 U19023 ( .B1(n22258), .B2(n20759), .A(n16986), .ZN(n16987) );
  AOI21_X1 U19024 ( .B1(n22254), .B2(n20762), .A(n16987), .ZN(n16988) );
  OAI21_X1 U19025 ( .B1(n17216), .B2(n22277), .A(n16988), .ZN(P1_U2978) );
  OAI21_X1 U19026 ( .B1(n17220), .B2(n16990), .A(n16989), .ZN(n16991) );
  XNOR2_X1 U19027 ( .A(n16991), .B(n17222), .ZN(n17228) );
  NAND2_X1 U19028 ( .A1(n22240), .A2(n20761), .ZN(n16992) );
  NAND2_X1 U19029 ( .A1(n22021), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n17221) );
  OAI211_X1 U19030 ( .C1(n20728), .C2(n16993), .A(n16992), .B(n17221), .ZN(
        n16994) );
  AOI21_X1 U19031 ( .B1(n16995), .B2(n20762), .A(n16994), .ZN(n16996) );
  OAI21_X1 U19032 ( .B1(n22277), .B2(n17228), .A(n16996), .ZN(P1_U2979) );
  XNOR2_X1 U19033 ( .A(n17256), .B(n17220), .ZN(n16997) );
  XNOR2_X1 U19034 ( .A(n16998), .B(n16997), .ZN(n17235) );
  NAND2_X1 U19035 ( .A1(n22021), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n17230) );
  NAND2_X1 U19036 ( .A1(n20760), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16999) );
  OAI211_X1 U19037 ( .C1(n17000), .C2(n20759), .A(n17230), .B(n16999), .ZN(
        n17001) );
  AOI21_X1 U19038 ( .B1(n20712), .B2(n20762), .A(n17001), .ZN(n17002) );
  OAI21_X1 U19039 ( .B1(n17235), .B2(n22277), .A(n17002), .ZN(P1_U2980) );
  XNOR2_X1 U19040 ( .A(n11165), .B(n17003), .ZN(n17249) );
  NOR2_X1 U19041 ( .A1(n22066), .A2(n22232), .ZN(n17242) );
  AOI21_X1 U19042 ( .B1(n20760), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n17242), .ZN(n17005) );
  OAI21_X1 U19043 ( .B1(n22222), .B2(n20759), .A(n17005), .ZN(n17006) );
  AOI21_X1 U19044 ( .B1(n22229), .B2(n20762), .A(n17006), .ZN(n17007) );
  OAI21_X1 U19045 ( .B1(n17249), .B2(n22277), .A(n17007), .ZN(P1_U2981) );
  INV_X1 U19046 ( .A(n17009), .ZN(n17011) );
  AOI21_X1 U19047 ( .B1(n17008), .B2(n17011), .A(n17010), .ZN(n17023) );
  INV_X1 U19048 ( .A(n17014), .ZN(n17012) );
  NOR2_X1 U19049 ( .A1(n17013), .A2(n17012), .ZN(n17022) );
  NAND2_X1 U19050 ( .A1(n17023), .A2(n17022), .ZN(n17021) );
  NAND2_X1 U19051 ( .A1(n17021), .A2(n17014), .ZN(n17015) );
  XOR2_X1 U19052 ( .A(n17016), .B(n17015), .Z(n17277) );
  NAND2_X1 U19053 ( .A1(n22021), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n17267) );
  OAI21_X1 U19054 ( .B1(n20728), .B2(n17017), .A(n17267), .ZN(n17019) );
  NOR2_X1 U19055 ( .A1(n22205), .A2(n17060), .ZN(n17018) );
  AOI211_X1 U19056 ( .C1(n20761), .C2(n22197), .A(n17019), .B(n17018), .ZN(
        n17020) );
  OAI21_X1 U19057 ( .B1(n17277), .B2(n22277), .A(n17020), .ZN(P1_U2983) );
  OAI21_X1 U19058 ( .B1(n17023), .B2(n17022), .A(n17021), .ZN(n17278) );
  NAND2_X1 U19059 ( .A1(n17278), .A2(n20756), .ZN(n17027) );
  OAI22_X1 U19060 ( .A1(n20728), .A2(n22184), .B1(n22066), .B2(n17024), .ZN(
        n17025) );
  AOI21_X1 U19061 ( .B1(n20761), .B2(n22187), .A(n17025), .ZN(n17026) );
  OAI211_X1 U19062 ( .C1(n17060), .C2(n20707), .A(n17027), .B(n17026), .ZN(
        P1_U2984) );
  INV_X1 U19063 ( .A(n17008), .ZN(n17030) );
  AOI21_X1 U19064 ( .B1(n17030), .B2(n17029), .A(n17028), .ZN(n17031) );
  AOI21_X1 U19065 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n11541), .A(
        n17031), .ZN(n17033) );
  MUX2_X1 U19066 ( .A(n16348), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .S(
        n17256), .Z(n17032) );
  XNOR2_X1 U19067 ( .A(n17033), .B(n17032), .ZN(n21982) );
  NAND2_X1 U19068 ( .A1(n21982), .A2(n20756), .ZN(n17038) );
  NAND2_X1 U19069 ( .A1(n22021), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n21979) );
  INV_X1 U19070 ( .A(n21979), .ZN(n17036) );
  NOR2_X1 U19071 ( .A1(n20759), .A2(n17034), .ZN(n17035) );
  AOI211_X1 U19072 ( .C1(n20760), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17036), .B(n17035), .ZN(n17037) );
  OAI211_X1 U19073 ( .C1(n17060), .C2(n17039), .A(n17038), .B(n17037), .ZN(
        P1_U2985) );
  INV_X1 U19074 ( .A(n17040), .ZN(n17041) );
  AOI21_X1 U19075 ( .B1(n17008), .B2(n17042), .A(n17041), .ZN(n17055) );
  AND2_X1 U19076 ( .A1(n17043), .A2(n17044), .ZN(n17054) );
  NAND2_X1 U19077 ( .A1(n17055), .A2(n17054), .ZN(n17053) );
  NAND2_X1 U19078 ( .A1(n17053), .A2(n17044), .ZN(n17045) );
  XOR2_X1 U19079 ( .A(n17046), .B(n17045), .Z(n17298) );
  NOR2_X1 U19080 ( .A1(n22066), .A2(n17047), .ZN(n17292) );
  AOI21_X1 U19081 ( .B1(n20760), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n17292), .ZN(n17048) );
  OAI21_X1 U19082 ( .B1(n17049), .B2(n20759), .A(n17048), .ZN(n17050) );
  AOI21_X1 U19083 ( .B1(n17051), .B2(n20762), .A(n17050), .ZN(n17052) );
  OAI21_X1 U19084 ( .B1(n17298), .B2(n22277), .A(n17052), .ZN(P1_U2986) );
  OAI21_X1 U19085 ( .B1(n17055), .B2(n17054), .A(n17053), .ZN(n17301) );
  NAND2_X1 U19086 ( .A1(n17301), .A2(n20756), .ZN(n17058) );
  NOR2_X1 U19087 ( .A1(n22066), .A2(n22177), .ZN(n17314) );
  NOR2_X1 U19088 ( .A1(n20728), .A2(n22175), .ZN(n17056) );
  AOI211_X1 U19089 ( .C1(n20761), .C2(n22169), .A(n17314), .B(n17056), .ZN(
        n17057) );
  OAI211_X1 U19090 ( .C1(n17060), .C2(n17059), .A(n17058), .B(n17057), .ZN(
        P1_U2987) );
  NOR2_X1 U19091 ( .A1(n17008), .A2(n17256), .ZN(n17062) );
  MUX2_X1 U19092 ( .A(n17061), .B(n17008), .S(n11541), .Z(n17069) );
  NOR2_X1 U19093 ( .A1(n17069), .A2(n22073), .ZN(n17068) );
  MUX2_X1 U19094 ( .A(n17062), .B(n17256), .S(n17068), .Z(n17063) );
  XNOR2_X1 U19095 ( .A(n17063), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17326) );
  NOR2_X1 U19096 ( .A1(n22066), .A2(n17064), .ZN(n17323) );
  AOI21_X1 U19097 ( .B1(n20760), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n17323), .ZN(n17065) );
  OAI21_X1 U19098 ( .B1(n22167), .B2(n20759), .A(n17065), .ZN(n17066) );
  AOI21_X1 U19099 ( .B1(n22163), .B2(n20762), .A(n17066), .ZN(n17067) );
  OAI21_X1 U19100 ( .B1(n17326), .B2(n22277), .A(n17067), .ZN(P1_U2988) );
  AOI21_X1 U19101 ( .B1(n22073), .B2(n17069), .A(n17068), .ZN(n22071) );
  INV_X1 U19102 ( .A(n22071), .ZN(n17075) );
  AOI22_X1 U19103 ( .A1(n20760), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n22021), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n17070) );
  OAI21_X1 U19104 ( .B1(n17071), .B2(n20759), .A(n17070), .ZN(n17072) );
  AOI21_X1 U19105 ( .B1(n17073), .B2(n20762), .A(n17072), .ZN(n17074) );
  OAI21_X1 U19106 ( .B1(n17075), .B2(n22277), .A(n17074), .ZN(P1_U2989) );
  NAND2_X1 U19107 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17272) );
  NOR3_X1 U19108 ( .A1(n17284), .A2(n17076), .A3(n17272), .ZN(n17261) );
  NAND2_X1 U19109 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17261), .ZN(
        n17241) );
  NOR2_X1 U19110 ( .A1(n17244), .A2(n17241), .ZN(n17083) );
  INV_X1 U19111 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17308) );
  INV_X1 U19112 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n22065) );
  NOR2_X1 U19113 ( .A1(n22065), .A2(n22073), .ZN(n22064) );
  NAND2_X1 U19114 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n22044) );
  NOR3_X1 U19115 ( .A1(n22020), .A2(n17077), .A3(n22011), .ZN(n22014) );
  NAND2_X1 U19116 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n22014), .ZN(
        n22032) );
  NOR3_X1 U19117 ( .A1(n22044), .A2(n22032), .A3(n17078), .ZN(n22052) );
  NAND2_X1 U19118 ( .A1(n22064), .A2(n22052), .ZN(n17303) );
  NOR3_X1 U19119 ( .A1(n17308), .A2(n17311), .A3(n17303), .ZN(n17238) );
  NAND2_X1 U19120 ( .A1(n17083), .A2(n17238), .ZN(n17091) );
  NAND2_X1 U19121 ( .A1(n21987), .A2(n17091), .ZN(n17079) );
  NAND2_X1 U19122 ( .A1(n22051), .A2(n17079), .ZN(n17194) );
  NOR2_X1 U19123 ( .A1(n17198), .A2(n17080), .ZN(n17092) );
  NOR2_X1 U19124 ( .A1(n22053), .A2(n17092), .ZN(n17081) );
  OR2_X1 U19125 ( .A1(n17194), .A2(n17081), .ZN(n17088) );
  INV_X1 U19126 ( .A(n22064), .ZN(n17082) );
  INV_X1 U19127 ( .A(n22044), .ZN(n22050) );
  NOR2_X1 U19128 ( .A1(n21989), .A2(n22032), .ZN(n22027) );
  NAND2_X1 U19129 ( .A1(n22050), .A2(n22027), .ZN(n22055) );
  NOR2_X1 U19130 ( .A1(n17082), .A2(n22055), .ZN(n17190) );
  NAND2_X1 U19131 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17190), .ZN(
        n17302) );
  NOR2_X1 U19132 ( .A1(n17311), .A2(n17302), .ZN(n17240) );
  NAND2_X1 U19133 ( .A1(n17083), .A2(n17240), .ZN(n17195) );
  INV_X1 U19134 ( .A(n17092), .ZN(n17084) );
  NOR2_X1 U19135 ( .A1(n17195), .A2(n17084), .ZN(n17095) );
  AND2_X1 U19136 ( .A1(n17095), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17085) );
  NOR2_X1 U19137 ( .A1(n21999), .A2(n17085), .ZN(n17086) );
  NOR2_X1 U19138 ( .A1(n17088), .A2(n17086), .ZN(n17185) );
  NAND2_X1 U19139 ( .A1(n22053), .A2(n21999), .ZN(n22078) );
  NAND2_X1 U19140 ( .A1(n22078), .A2(n17155), .ZN(n17087) );
  NAND2_X1 U19141 ( .A1(n17185), .A2(n17087), .ZN(n17162) );
  OR2_X1 U19142 ( .A1(n17162), .A2(n17097), .ZN(n17090) );
  INV_X1 U19143 ( .A(n17088), .ZN(n17089) );
  INV_X1 U19144 ( .A(n22078), .ZN(n22015) );
  NAND2_X1 U19145 ( .A1(n17089), .A2(n22015), .ZN(n17110) );
  NAND2_X1 U19146 ( .A1(n17090), .A2(n17110), .ZN(n17146) );
  NAND2_X1 U19147 ( .A1(n17146), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17114) );
  NOR2_X1 U19148 ( .A1(n22015), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17112) );
  NOR3_X1 U19149 ( .A1(n17114), .A2(n17112), .A3(n17122), .ZN(n17104) );
  NAND2_X1 U19150 ( .A1(n17110), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17103) );
  INV_X1 U19151 ( .A(n17091), .ZN(n17093) );
  NAND2_X1 U19152 ( .A1(n17093), .A2(n17092), .ZN(n17094) );
  OR2_X1 U19153 ( .A1(n21992), .A2(n17094), .ZN(n17171) );
  NAND2_X1 U19154 ( .A1(n22056), .A2(n17095), .ZN(n17096) );
  NAND2_X1 U19155 ( .A1(n17171), .A2(n17096), .ZN(n17182) );
  NOR2_X1 U19156 ( .A1(n17155), .A2(n17097), .ZN(n17098) );
  NAND2_X1 U19157 ( .A1(n17182), .A2(n17098), .ZN(n17141) );
  NOR3_X1 U19158 ( .A1(n17141), .A2(n17122), .A3(n17099), .ZN(n17113) );
  NAND3_X1 U19159 ( .A1(n17113), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n17100), .ZN(n17102) );
  OAI211_X1 U19160 ( .C1(n17104), .C2(n17103), .A(n17102), .B(n17101), .ZN(
        n17105) );
  AOI21_X1 U19161 ( .B1(n17106), .B2(n22043), .A(n17105), .ZN(n17107) );
  OAI21_X1 U19162 ( .B1(n17108), .B2(n22058), .A(n17107), .ZN(P1_U3000) );
  INV_X1 U19163 ( .A(n17109), .ZN(n17119) );
  INV_X1 U19164 ( .A(n17110), .ZN(n17111) );
  OAI21_X1 U19165 ( .B1(n16360), .B2(n17111), .A(n17146), .ZN(n17125) );
  OAI21_X1 U19166 ( .B1(n17125), .B2(n17112), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17117) );
  NAND2_X1 U19167 ( .A1(n17114), .A2(n17113), .ZN(n17115) );
  NAND3_X1 U19168 ( .A1(n17117), .A2(n17116), .A3(n17115), .ZN(n17118) );
  AOI21_X1 U19169 ( .B1(n17119), .B2(n22043), .A(n17118), .ZN(n17120) );
  OAI21_X1 U19170 ( .B1(n17121), .B2(n22058), .A(n17120), .ZN(P1_U3001) );
  NOR3_X1 U19171 ( .A1(n17141), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n17122), .ZN(n17123) );
  AOI211_X1 U19172 ( .C1(n17125), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n17124), .B(n17123), .ZN(n17129) );
  INV_X1 U19173 ( .A(n17126), .ZN(n17127) );
  NAND2_X1 U19174 ( .A1(n17127), .A2(n22043), .ZN(n17128) );
  OAI211_X1 U19175 ( .C1(n17130), .C2(n22058), .A(n17129), .B(n17128), .ZN(
        P1_U3002) );
  INV_X1 U19176 ( .A(n17146), .ZN(n17135) );
  INV_X1 U19177 ( .A(n17131), .ZN(n17134) );
  NOR3_X1 U19178 ( .A1(n17141), .A2(n16360), .A3(n17132), .ZN(n17133) );
  AOI211_X1 U19179 ( .C1(n17135), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n17134), .B(n17133), .ZN(n17139) );
  INV_X1 U19180 ( .A(n17136), .ZN(n17137) );
  NAND2_X1 U19181 ( .A1(n17137), .A2(n22043), .ZN(n17138) );
  OAI211_X1 U19182 ( .C1(n17140), .C2(n22058), .A(n17139), .B(n17138), .ZN(
        P1_U3003) );
  INV_X1 U19183 ( .A(n17141), .ZN(n17143) );
  AOI21_X1 U19184 ( .B1(n17143), .B2(n17145), .A(n17142), .ZN(n17144) );
  OAI21_X1 U19185 ( .B1(n17146), .B2(n17145), .A(n17144), .ZN(n17147) );
  AOI21_X1 U19186 ( .B1(n17148), .B2(n22043), .A(n17147), .ZN(n17149) );
  OAI21_X1 U19187 ( .B1(n17150), .B2(n22058), .A(n17149), .ZN(P1_U3004) );
  INV_X1 U19188 ( .A(n17151), .ZN(n17161) );
  NAND3_X1 U19189 ( .A1(n17153), .A2(n22075), .A3(n17152), .ZN(n17160) );
  INV_X1 U19190 ( .A(n17154), .ZN(n17158) );
  INV_X1 U19191 ( .A(n17182), .ZN(n17156) );
  NOR3_X1 U19192 ( .A1(n17156), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n17155), .ZN(n17157) );
  AOI211_X1 U19193 ( .C1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n17162), .A(
        n17158), .B(n17157), .ZN(n17159) );
  OAI211_X1 U19194 ( .C1(n22082), .C2(n17161), .A(n17160), .B(n17159), .ZN(
        P1_U3005) );
  INV_X1 U19195 ( .A(n17162), .ZN(n17165) );
  AOI21_X1 U19196 ( .B1(n17182), .B2(n17163), .A(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17164) );
  NOR2_X1 U19197 ( .A1(n17165), .A2(n17164), .ZN(n17166) );
  AOI211_X1 U19198 ( .C1(n17168), .C2(n22043), .A(n17167), .B(n17166), .ZN(
        n17169) );
  OAI21_X1 U19199 ( .B1(n17170), .B2(n22058), .A(n17169), .ZN(P1_U3006) );
  OAI21_X1 U19200 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17171), .A(
        n17185), .ZN(n17178) );
  NAND3_X1 U19201 ( .A1(n17182), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n17172), .ZN(n17174) );
  NAND2_X1 U19202 ( .A1(n17174), .A2(n17173), .ZN(n17177) );
  NOR2_X1 U19203 ( .A1(n17175), .A2(n22082), .ZN(n17176) );
  AOI211_X1 U19204 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n17178), .A(
        n17177), .B(n17176), .ZN(n17179) );
  OAI21_X1 U19205 ( .B1(n17180), .B2(n22058), .A(n17179), .ZN(P1_U3007) );
  AOI21_X1 U19206 ( .B1(n17182), .B2(n17184), .A(n17181), .ZN(n17183) );
  OAI21_X1 U19207 ( .B1(n17185), .B2(n17184), .A(n17183), .ZN(n17186) );
  AOI21_X1 U19208 ( .B1(n17187), .B2(n22043), .A(n17186), .ZN(n17188) );
  OAI21_X1 U19209 ( .B1(n17189), .B2(n22058), .A(n17188), .ZN(P1_U3008) );
  INV_X1 U19210 ( .A(n22275), .ZN(n17203) );
  OR2_X1 U19211 ( .A1(n21992), .A2(n17303), .ZN(n17191) );
  NAND2_X1 U19212 ( .A1(n22056), .A2(n17190), .ZN(n17217) );
  NAND2_X1 U19213 ( .A1(n17191), .A2(n17217), .ZN(n17315) );
  INV_X1 U19214 ( .A(n17195), .ZN(n17219) );
  NAND2_X1 U19215 ( .A1(n17315), .A2(n17219), .ZN(n17232) );
  INV_X1 U19216 ( .A(n17192), .ZN(n17193) );
  NOR3_X1 U19217 ( .A1(n17232), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n17193), .ZN(n17206) );
  INV_X1 U19218 ( .A(n17194), .ZN(n17218) );
  NOR3_X1 U19219 ( .A1(n17222), .A2(n17220), .A3(n17195), .ZN(n17197) );
  NOR2_X1 U19220 ( .A1(n22078), .A2(n22030), .ZN(n17196) );
  AOI21_X1 U19221 ( .B1(n17218), .B2(n17197), .A(n17196), .ZN(n17208) );
  OAI21_X1 U19222 ( .B1(n17206), .B2(n17208), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17201) );
  OR3_X1 U19223 ( .A1(n17232), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n17198), .ZN(n17199) );
  NAND3_X1 U19224 ( .A1(n17201), .A2(n17200), .A3(n17199), .ZN(n17202) );
  AOI21_X1 U19225 ( .B1(n17203), .B2(n22043), .A(n17202), .ZN(n17204) );
  OAI21_X1 U19226 ( .B1(n17205), .B2(n22058), .A(n17204), .ZN(P1_U3009) );
  AOI211_X1 U19227 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n17208), .A(
        n17207), .B(n17206), .ZN(n17215) );
  NAND2_X1 U19228 ( .A1(n17210), .A2(n17209), .ZN(n17211) );
  NAND2_X1 U19229 ( .A1(n17212), .A2(n17211), .ZN(n22251) );
  INV_X1 U19230 ( .A(n22251), .ZN(n17213) );
  NAND2_X1 U19231 ( .A1(n17213), .A2(n22043), .ZN(n17214) );
  OAI211_X1 U19232 ( .C1(n17216), .C2(n22058), .A(n17215), .B(n17214), .ZN(
        P1_U3010) );
  NOR3_X1 U19233 ( .A1(n17232), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n17220), .ZN(n17225) );
  NAND2_X1 U19234 ( .A1(n21992), .A2(n17217), .ZN(n17291) );
  OAI21_X1 U19235 ( .B1(n21999), .B2(n17219), .A(n17218), .ZN(n17229) );
  AOI21_X1 U19236 ( .B1(n17220), .B2(n17291), .A(n17229), .ZN(n17223) );
  OAI21_X1 U19237 ( .B1(n17223), .B2(n17222), .A(n17221), .ZN(n17224) );
  AOI211_X1 U19238 ( .C1(n17226), .C2(n22043), .A(n17225), .B(n17224), .ZN(
        n17227) );
  OAI21_X1 U19239 ( .B1(n17228), .B2(n22058), .A(n17227), .ZN(P1_U3011) );
  NAND2_X1 U19240 ( .A1(n17229), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17231) );
  OAI211_X1 U19241 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17232), .A(
        n17231), .B(n17230), .ZN(n17233) );
  AOI21_X1 U19242 ( .B1(n20711), .B2(n22043), .A(n17233), .ZN(n17234) );
  OAI21_X1 U19243 ( .B1(n17235), .B2(n22058), .A(n17234), .ZN(P1_U3012) );
  INV_X1 U19244 ( .A(n22226), .ZN(n17247) );
  AND2_X1 U19245 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17236) );
  INV_X1 U19246 ( .A(n21976), .ZN(n17237) );
  NOR3_X1 U19247 ( .A1(n17237), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17241), .ZN(n17246) );
  OR2_X1 U19248 ( .A1(n22053), .A2(n17238), .ZN(n17239) );
  OAI211_X1 U19249 ( .C1(n17240), .C2(n21999), .A(n22051), .B(n17239), .ZN(
        n21977) );
  AOI21_X1 U19250 ( .B1(n22078), .B2(n17241), .A(n21977), .ZN(n17263) );
  INV_X1 U19251 ( .A(n17242), .ZN(n17243) );
  OAI21_X1 U19252 ( .B1(n17263), .B2(n17244), .A(n17243), .ZN(n17245) );
  AOI211_X1 U19253 ( .C1(n17247), .C2(n22043), .A(n17246), .B(n17245), .ZN(
        n17248) );
  OAI21_X1 U19254 ( .B1(n17249), .B2(n22058), .A(n17248), .ZN(P1_U3013) );
  NOR2_X1 U19255 ( .A1(n17256), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17255) );
  INV_X1 U19256 ( .A(n17251), .ZN(n17253) );
  OAI21_X1 U19257 ( .B1(n17008), .B2(n17253), .A(n17252), .ZN(n17254) );
  MUX2_X1 U19258 ( .A(n17256), .B(n17255), .S(n17254), .Z(n17257) );
  XNOR2_X1 U19259 ( .A(n17257), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n20765) );
  AOI21_X1 U19260 ( .B1(n17260), .B2(n17259), .A(n17258), .ZN(n22216) );
  AOI21_X1 U19261 ( .B1(n21976), .B2(n17261), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17264) );
  INV_X1 U19262 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n17262) );
  OAI22_X1 U19263 ( .A1(n17264), .A2(n17263), .B1(n22066), .B2(n17262), .ZN(
        n17265) );
  AOI21_X1 U19264 ( .B1(n22216), .B2(n22043), .A(n17265), .ZN(n17266) );
  OAI21_X1 U19265 ( .B1(n20765), .B2(n22058), .A(n17266), .ZN(P1_U3014) );
  INV_X1 U19266 ( .A(n22208), .ZN(n17270) );
  INV_X1 U19267 ( .A(n17267), .ZN(n17269) );
  NAND3_X1 U19268 ( .A1(n21976), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17271) );
  NOR3_X1 U19269 ( .A1(n17271), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n17284), .ZN(n17268) );
  AOI211_X1 U19270 ( .C1(n17270), .C2(n22043), .A(n17269), .B(n17268), .ZN(
        n17276) );
  NOR2_X1 U19271 ( .A1(n17271), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17286) );
  INV_X1 U19272 ( .A(n17272), .ZN(n17274) );
  INV_X1 U19273 ( .A(n21977), .ZN(n17273) );
  OAI21_X1 U19274 ( .B1(n22015), .B2(n17274), .A(n17273), .ZN(n17282) );
  OAI21_X1 U19275 ( .B1(n17286), .B2(n17282), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17275) );
  OAI211_X1 U19276 ( .C1(n17277), .C2(n22058), .A(n17276), .B(n17275), .ZN(
        P1_U3015) );
  INV_X1 U19277 ( .A(n17278), .ZN(n17289) );
  NAND2_X1 U19278 ( .A1(n16155), .A2(n17279), .ZN(n17280) );
  AND2_X1 U19279 ( .A1(n17281), .A2(n17280), .ZN(n22186) );
  INV_X1 U19280 ( .A(n17282), .ZN(n17285) );
  NAND2_X1 U19281 ( .A1(n22021), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n17283) );
  OAI21_X1 U19282 ( .B1(n17285), .B2(n17284), .A(n17283), .ZN(n17287) );
  AOI211_X1 U19283 ( .C1(n22043), .C2(n22186), .A(n17287), .B(n17286), .ZN(
        n17288) );
  OAI21_X1 U19284 ( .B1(n17289), .B2(n22058), .A(n17288), .ZN(P1_U3016) );
  INV_X1 U19285 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17290) );
  AND2_X1 U19286 ( .A1(n17291), .A2(n17290), .ZN(n21978) );
  NAND2_X1 U19287 ( .A1(n21976), .A2(n21978), .ZN(n17294) );
  AOI21_X1 U19288 ( .B1(n21977), .B2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n17292), .ZN(n17293) );
  NAND2_X1 U19289 ( .A1(n17294), .A2(n17293), .ZN(n17295) );
  AOI21_X1 U19290 ( .B1(n17296), .B2(n22043), .A(n17295), .ZN(n17297) );
  OAI21_X1 U19291 ( .B1(n17298), .B2(n22058), .A(n17297), .ZN(P1_U3018) );
  INV_X1 U19292 ( .A(n17299), .ZN(n17300) );
  XNOR2_X1 U19293 ( .A(n17322), .B(n17300), .ZN(n22172) );
  NAND2_X1 U19294 ( .A1(n17301), .A2(n22075), .ZN(n17318) );
  NOR2_X1 U19295 ( .A1(n17308), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17316) );
  INV_X1 U19296 ( .A(n17302), .ZN(n17307) );
  INV_X1 U19297 ( .A(n17303), .ZN(n17304) );
  OAI21_X1 U19298 ( .B1(n22053), .B2(n17304), .A(n22051), .ZN(n17305) );
  INV_X1 U19299 ( .A(n17305), .ZN(n17306) );
  OAI21_X1 U19300 ( .B1(n21999), .B2(n17307), .A(n17306), .ZN(n17310) );
  OR2_X1 U19301 ( .A1(n17310), .A2(n17308), .ZN(n17309) );
  OAI21_X1 U19302 ( .B1(n17315), .B2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n17309), .ZN(n17324) );
  INV_X1 U19303 ( .A(n17310), .ZN(n17312) );
  AOI21_X1 U19304 ( .B1(n17324), .B2(n17312), .A(n17311), .ZN(n17313) );
  AOI211_X1 U19305 ( .C1(n17316), .C2(n17315), .A(n17314), .B(n17313), .ZN(
        n17317) );
  OAI211_X1 U19306 ( .C1(n22172), .C2(n22082), .A(n17318), .B(n17317), .ZN(
        P1_U3019) );
  NAND2_X1 U19307 ( .A1(n17320), .A2(n17319), .ZN(n17321) );
  AND2_X1 U19308 ( .A1(n17322), .A2(n17321), .ZN(n22157) );
  AOI21_X1 U19309 ( .B1(n22157), .B2(n22043), .A(n17323), .ZN(n17325) );
  OAI211_X1 U19310 ( .C1(n17326), .C2(n22058), .A(n17325), .B(n17324), .ZN(
        P1_U3020) );
  NAND2_X1 U19311 ( .A1(n22422), .A2(n22434), .ZN(n17329) );
  NOR2_X1 U19312 ( .A1(n11196), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n17327) );
  INV_X1 U19313 ( .A(n22281), .ZN(n17332) );
  OAI22_X1 U19314 ( .A1(n17329), .A2(n17327), .B1(n11193), .B2(n17332), .ZN(
        n17328) );
  MUX2_X1 U19315 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n17328), .S(
        n18023), .Z(P1_U3477) );
  MUX2_X1 U19316 ( .A(n17330), .B(n17329), .S(n11195), .Z(n17331) );
  OAI21_X1 U19317 ( .B1(n17332), .B2(n22418), .A(n17331), .ZN(n17333) );
  MUX2_X1 U19318 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n17333), .S(
        n18023), .Z(P1_U3476) );
  OAI21_X1 U19319 ( .B1(n17402), .B2(n17335), .A(n17334), .ZN(n17688) );
  OR2_X1 U19320 ( .A1(n17337), .A2(n17338), .ZN(n17339) );
  AND2_X1 U19321 ( .A1(n17336), .A2(n17339), .ZN(n17684) );
  AOI22_X1 U19322 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19346), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n19328), .ZN(n17340) );
  OAI21_X1 U19323 ( .B1(n19338), .B2(n18199), .A(n17340), .ZN(n17341) );
  AOI21_X1 U19324 ( .B1(n17684), .B2(n19348), .A(n17341), .ZN(n17342) );
  OAI21_X1 U19325 ( .B1(n17688), .B2(n19310), .A(n17342), .ZN(n17346) );
  AOI211_X1 U19326 ( .C1(n17344), .C2(n17515), .A(n19432), .B(n17343), .ZN(
        n17345) );
  AOI211_X1 U19327 ( .C1(n19323), .C2(n17347), .A(n17346), .B(n17345), .ZN(
        n17348) );
  INV_X1 U19328 ( .A(n17348), .ZN(P2_U2830) );
  OR2_X1 U19329 ( .A1(n17350), .A2(n17349), .ZN(n17351) );
  NAND2_X1 U19330 ( .A1(n14104), .A2(n17351), .ZN(n17719) );
  XNOR2_X1 U19331 ( .A(n17353), .B(n17352), .ZN(n17720) );
  AOI22_X1 U19332 ( .A1(n17354), .A2(n19323), .B1(P2_REIP_REG_22__SCAN_IN), 
        .B2(n19307), .ZN(n17356) );
  AOI22_X1 U19333 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19346), .B1(
        P2_EBX_REG_22__SCAN_IN), .B2(n19328), .ZN(n17355) );
  OAI211_X1 U19334 ( .C1(n17720), .C2(n19336), .A(n17356), .B(n17355), .ZN(
        n17361) );
  AOI211_X1 U19335 ( .C1(n17359), .C2(n17358), .A(n17357), .B(n19432), .ZN(
        n17360) );
  NOR2_X1 U19336 ( .A1(n17361), .A2(n17360), .ZN(n17362) );
  OAI21_X1 U19337 ( .B1(n17719), .B2(n19310), .A(n17362), .ZN(P2_U2833) );
  NOR2_X1 U19338 ( .A1(n11181), .A2(n17363), .ZN(n17364) );
  XNOR2_X1 U19339 ( .A(n17364), .B(n18069), .ZN(n17365) );
  NAND2_X1 U19340 ( .A1(n17365), .A2(n19316), .ZN(n17371) );
  AOI22_X1 U19341 ( .A1(n17366), .A2(n19323), .B1(P2_EBX_REG_8__SCAN_IN), .B2(
        n19328), .ZN(n17367) );
  OAI211_X1 U19342 ( .C1(n11761), .C2(n19338), .A(n17367), .B(n19258), .ZN(
        n17368) );
  AOI21_X1 U19343 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19346), .A(
        n17368), .ZN(n17370) );
  AOI22_X1 U19344 ( .A1(n19349), .A2(n19397), .B1(n19348), .B2(n19395), .ZN(
        n17369) );
  NAND3_X1 U19345 ( .A1(n17371), .A2(n17370), .A3(n17369), .ZN(P2_U2847) );
  NAND2_X1 U19346 ( .A1(n19350), .A2(n14580), .ZN(n17372) );
  OAI21_X1 U19347 ( .B1(n14580), .B2(n12219), .A(n17372), .ZN(P2_U2856) );
  INV_X1 U19348 ( .A(n17373), .ZN(n17380) );
  NAND2_X1 U19349 ( .A1(n17380), .A2(n17374), .ZN(n17376) );
  XNOR2_X1 U19350 ( .A(n17376), .B(n17375), .ZN(n17434) );
  NOR2_X1 U19351 ( .A1(n19311), .A2(n17420), .ZN(n17377) );
  AOI21_X1 U19352 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n17423), .A(n17377), .ZN(
        n17378) );
  OAI21_X1 U19353 ( .B1(n17434), .B2(n17428), .A(n17378), .ZN(P2_U2859) );
  NAND2_X1 U19354 ( .A1(n17380), .A2(n17379), .ZN(n17381) );
  XOR2_X1 U19355 ( .A(n17382), .B(n17381), .Z(n17440) );
  NAND2_X1 U19356 ( .A1(n17423), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n17384) );
  NAND2_X1 U19357 ( .A1(n17491), .A2(n14580), .ZN(n17383) );
  OAI211_X1 U19358 ( .C1(n17440), .C2(n17428), .A(n17384), .B(n17383), .ZN(
        P2_U2860) );
  INV_X1 U19359 ( .A(n17385), .ZN(n17386) );
  AOI21_X1 U19360 ( .B1(n17387), .B2(n17334), .A(n17386), .ZN(n19297) );
  INV_X1 U19361 ( .A(n19297), .ZN(n17677) );
  AOI21_X1 U19362 ( .B1(n17388), .B2(n17390), .A(n17389), .ZN(n17441) );
  NAND2_X1 U19363 ( .A1(n17441), .A2(n17417), .ZN(n17392) );
  NAND2_X1 U19364 ( .A1(n17423), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n17391) );
  OAI211_X1 U19365 ( .C1(n17677), .C2(n17420), .A(n17392), .B(n17391), .ZN(
        P2_U2861) );
  OAI21_X1 U19366 ( .B1(n17393), .B2(n17395), .A(n17394), .ZN(n17455) );
  MUX2_X1 U19367 ( .A(n12208), .B(n17688), .S(n14580), .Z(n17396) );
  OAI21_X1 U19368 ( .B1(n17455), .B2(n17428), .A(n17396), .ZN(P2_U2862) );
  OAI21_X1 U19369 ( .B1(n17397), .B2(n17399), .A(n17398), .ZN(n17462) );
  AND2_X1 U19370 ( .A1(n17401), .A2(n17400), .ZN(n17403) );
  OR2_X1 U19371 ( .A1(n17403), .A2(n17402), .ZN(n19285) );
  NOR2_X1 U19372 ( .A1(n19285), .A2(n17420), .ZN(n17404) );
  AOI21_X1 U19373 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n17420), .A(n17404), .ZN(
        n17405) );
  OAI21_X1 U19374 ( .B1(n17462), .B2(n17428), .A(n17405), .ZN(P2_U2863) );
  XNOR2_X1 U19375 ( .A(n17406), .B(n17407), .ZN(n17467) );
  NAND2_X1 U19376 ( .A1(n17423), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n17409) );
  NAND2_X1 U19377 ( .A1(n17715), .A2(n14580), .ZN(n17408) );
  OAI211_X1 U19378 ( .C1(n17467), .C2(n17428), .A(n17409), .B(n17408), .ZN(
        P2_U2864) );
  OAI21_X1 U19379 ( .B1(n17410), .B2(n17411), .A(n17406), .ZN(n17473) );
  NOR2_X1 U19380 ( .A1(n17719), .A2(n17420), .ZN(n17412) );
  AOI21_X1 U19381 ( .B1(P2_EBX_REG_22__SCAN_IN), .B2(n17420), .A(n17412), .ZN(
        n17413) );
  OAI21_X1 U19382 ( .B1(n17473), .B2(n17428), .A(n17413), .ZN(P2_U2865) );
  AOI21_X1 U19383 ( .B1(n17416), .B2(n17414), .A(n17410), .ZN(n17474) );
  NAND2_X1 U19384 ( .A1(n17474), .A2(n17417), .ZN(n17419) );
  NAND2_X1 U19385 ( .A1(n17423), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n17418) );
  OAI211_X1 U19386 ( .C1(n17421), .C2(n17420), .A(n17419), .B(n17418), .ZN(
        P2_U2866) );
  OAI21_X1 U19387 ( .B1(n16432), .B2(n17422), .A(n17414), .ZN(n20224) );
  NAND2_X1 U19388 ( .A1(n17423), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n17427) );
  AND2_X1 U19389 ( .A1(n16215), .A2(n17424), .ZN(n17425) );
  NOR2_X1 U19390 ( .A1(n12769), .A2(n17425), .ZN(n19273) );
  NAND2_X1 U19391 ( .A1(n19273), .A2(n14580), .ZN(n17426) );
  OAI211_X1 U19392 ( .C1(n20224), .C2(n17428), .A(n17427), .B(n17426), .ZN(
        P2_U2867) );
  OAI22_X1 U19393 ( .A1(n17477), .A2(n19309), .B1(n17475), .B2(n17429), .ZN(
        n17430) );
  AOI21_X1 U19394 ( .B1(n17479), .B2(n17431), .A(n17430), .ZN(n17433) );
  AOI22_X1 U19395 ( .A1(n19914), .A2(BUF2_REG_28__SCAN_IN), .B1(n19915), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n17432) );
  OAI211_X1 U19396 ( .C1(n17434), .C2(n20165), .A(n17433), .B(n17432), .ZN(
        P2_U2891) );
  OAI22_X1 U19397 ( .A1(n17477), .A2(n17661), .B1(n17475), .B2(n17435), .ZN(
        n17436) );
  AOI21_X1 U19398 ( .B1(n17479), .B2(n17437), .A(n17436), .ZN(n17439) );
  AOI22_X1 U19399 ( .A1(n19914), .A2(BUF2_REG_27__SCAN_IN), .B1(n19915), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n17438) );
  OAI211_X1 U19400 ( .C1(n17440), .C2(n20165), .A(n17439), .B(n17438), .ZN(
        P2_U2892) );
  NAND2_X1 U19401 ( .A1(n17441), .A2(n20322), .ZN(n17448) );
  NAND2_X1 U19402 ( .A1(n17336), .A2(n17442), .ZN(n17443) );
  AND2_X1 U19403 ( .A1(n14084), .A2(n17443), .ZN(n19296) );
  AOI22_X1 U19404 ( .A1(n20321), .A2(n19296), .B1(n20319), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n17447) );
  AOI22_X1 U19405 ( .A1(n19914), .A2(BUF2_REG_26__SCAN_IN), .B1(n19915), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n17446) );
  NAND2_X1 U19406 ( .A1(n17479), .A2(n17444), .ZN(n17445) );
  NAND4_X1 U19407 ( .A1(n17448), .A2(n17447), .A3(n17446), .A4(n17445), .ZN(
        P2_U2893) );
  INV_X1 U19408 ( .A(n17684), .ZN(n17450) );
  OAI22_X1 U19409 ( .A1(n17477), .A2(n17450), .B1(n17475), .B2(n17449), .ZN(
        n17451) );
  AOI21_X1 U19410 ( .B1(n17479), .B2(n17452), .A(n17451), .ZN(n17454) );
  AOI22_X1 U19411 ( .A1(n19914), .A2(BUF2_REG_25__SCAN_IN), .B1(n19915), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n17453) );
  OAI211_X1 U19412 ( .C1(n17455), .C2(n20165), .A(n17454), .B(n17453), .ZN(
        P2_U2894) );
  AND2_X1 U19413 ( .A1(n14107), .A2(n17456), .ZN(n17457) );
  OR2_X1 U19414 ( .A1(n17337), .A2(n17457), .ZN(n19284) );
  OAI22_X1 U19415 ( .A1(n17477), .A2(n19284), .B1(n17475), .B2(n14277), .ZN(
        n17458) );
  AOI21_X1 U19416 ( .B1(n17479), .B2(n17459), .A(n17458), .ZN(n17461) );
  AOI22_X1 U19417 ( .A1(n19914), .A2(BUF2_REG_24__SCAN_IN), .B1(n19915), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n17460) );
  OAI211_X1 U19418 ( .C1(n17462), .C2(n20165), .A(n17461), .B(n17460), .ZN(
        P2_U2895) );
  OAI22_X1 U19419 ( .A1(n17477), .A2(n17712), .B1(n17475), .B2(n14275), .ZN(
        n17463) );
  AOI21_X1 U19420 ( .B1(n17479), .B2(n17464), .A(n17463), .ZN(n17466) );
  AOI22_X1 U19421 ( .A1(n19914), .A2(BUF2_REG_23__SCAN_IN), .B1(n19915), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n17465) );
  OAI211_X1 U19422 ( .C1(n17467), .C2(n20165), .A(n17466), .B(n17465), .ZN(
        P2_U2896) );
  OAI22_X1 U19423 ( .A1(n17477), .A2(n17720), .B1(n17475), .B2(n14271), .ZN(
        n17470) );
  INV_X1 U19424 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n17468) );
  OAI22_X1 U19425 ( .A1(n20317), .A2(n20809), .B1(n20327), .B2(n17468), .ZN(
        n17469) );
  AOI211_X1 U19426 ( .C1(n17479), .C2(n17471), .A(n17470), .B(n17469), .ZN(
        n17472) );
  OAI21_X1 U19427 ( .B1(n17473), .B2(n20165), .A(n17472), .ZN(P2_U2897) );
  INV_X1 U19428 ( .A(n17474), .ZN(n17482) );
  OAI22_X1 U19429 ( .A1(n17477), .A2(n17476), .B1(n17475), .B2(n14269), .ZN(
        n17478) );
  AOI21_X1 U19430 ( .B1(n17479), .B2(n20163), .A(n17478), .ZN(n17481) );
  AOI22_X1 U19431 ( .A1(n19914), .A2(BUF2_REG_21__SCAN_IN), .B1(n19915), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n17480) );
  OAI211_X1 U19432 ( .C1(n17482), .C2(n20165), .A(n17481), .B(n17480), .ZN(
        P2_U2898) );
  INV_X1 U19433 ( .A(n17483), .ZN(n17485) );
  XNOR2_X1 U19434 ( .A(n17486), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17670) );
  NAND2_X1 U19435 ( .A1(n18070), .A2(n17487), .ZN(n17488) );
  NAND2_X1 U19436 ( .A1(n19407), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n17660) );
  OAI211_X1 U19437 ( .C1(n18076), .C2(n17489), .A(n17488), .B(n17660), .ZN(
        n17490) );
  AOI21_X1 U19438 ( .B1(n17491), .B2(n18091), .A(n17490), .ZN(n17496) );
  INV_X1 U19439 ( .A(n17492), .ZN(n17498) );
  AOI21_X1 U19440 ( .B1(n17494), .B2(n17498), .A(n17493), .ZN(n17668) );
  NAND2_X1 U19441 ( .A1(n17668), .A2(n18095), .ZN(n17495) );
  OAI211_X1 U19442 ( .C1(n17670), .C2(n18106), .A(n17496), .B(n17495), .ZN(
        P2_U2987) );
  NOR2_X1 U19443 ( .A1(n17518), .A2(n17691), .ZN(n17511) );
  OAI21_X1 U19444 ( .B1(n17511), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17498), .ZN(n17681) );
  AOI21_X1 U19445 ( .B1(n17499), .B2(n17508), .A(n17507), .ZN(n17501) );
  XNOR2_X1 U19446 ( .A(n17501), .B(n17500), .ZN(n17679) );
  NAND2_X1 U19447 ( .A1(n19297), .A2(n18091), .ZN(n17503) );
  NOR2_X1 U19448 ( .A1(n19380), .A2(n18200), .ZN(n17673) );
  AOI21_X1 U19449 ( .B1(n18102), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n17673), .ZN(n17502) );
  OAI211_X1 U19450 ( .C1(n18112), .C2(n17504), .A(n17503), .B(n17502), .ZN(
        n17505) );
  AOI21_X1 U19451 ( .B1(n17679), .B2(n18079), .A(n17505), .ZN(n17506) );
  OAI21_X1 U19452 ( .B1(n18103), .B2(n17681), .A(n17506), .ZN(P2_U2988) );
  INV_X1 U19453 ( .A(n17507), .ZN(n17509) );
  NAND2_X1 U19454 ( .A1(n17509), .A2(n17508), .ZN(n17510) );
  XNOR2_X1 U19455 ( .A(n17499), .B(n17510), .ZN(n17695) );
  INV_X1 U19456 ( .A(n17511), .ZN(n17683) );
  NAND2_X1 U19457 ( .A1(n17518), .A2(n17691), .ZN(n17682) );
  NAND3_X1 U19458 ( .A1(n17683), .A2(n18095), .A3(n17682), .ZN(n17517) );
  NAND2_X1 U19459 ( .A1(n19407), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n17685) );
  OAI21_X1 U19460 ( .B1(n18076), .B2(n17512), .A(n17685), .ZN(n17514) );
  NOR2_X1 U19461 ( .A1(n17688), .A2(n18105), .ZN(n17513) );
  AOI211_X1 U19462 ( .C1(n18070), .C2(n17515), .A(n17514), .B(n17513), .ZN(
        n17516) );
  OAI211_X1 U19463 ( .C1(n18106), .C2(n17695), .A(n17517), .B(n17516), .ZN(
        P2_U2989) );
  OAI21_X1 U19464 ( .B1(n11208), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n17518), .ZN(n17705) );
  XOR2_X1 U19465 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17520), .Z(
        n17521) );
  XNOR2_X1 U19466 ( .A(n17519), .B(n17521), .ZN(n17703) );
  NOR2_X1 U19467 ( .A1(n19380), .A2(n18198), .ZN(n17696) );
  NOR2_X1 U19468 ( .A1(n18112), .A2(n17522), .ZN(n17523) );
  AOI211_X1 U19469 ( .C1(n18102), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n17696), .B(n17523), .ZN(n17524) );
  OAI21_X1 U19470 ( .B1(n19285), .B2(n18105), .A(n17524), .ZN(n17525) );
  AOI21_X1 U19471 ( .B1(n17703), .B2(n18079), .A(n17525), .ZN(n17526) );
  OAI21_X1 U19472 ( .B1(n17705), .B2(n18103), .A(n17526), .ZN(P2_U2990) );
  INV_X1 U19473 ( .A(n17528), .ZN(n17530) );
  NAND2_X1 U19474 ( .A1(n17530), .A2(n17529), .ZN(n17531) );
  XNOR2_X1 U19475 ( .A(n17527), .B(n17531), .ZN(n17718) );
  OR2_X1 U19476 ( .A1(n17537), .A2(n17708), .ZN(n17538) );
  AOI21_X1 U19477 ( .B1(n17709), .B2(n17538), .A(n11208), .ZN(n17706) );
  NAND2_X1 U19478 ( .A1(n17706), .A2(n18095), .ZN(n17536) );
  NAND2_X1 U19479 ( .A1(n18070), .A2(n17532), .ZN(n17533) );
  NAND2_X1 U19480 ( .A1(n19407), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n17710) );
  OAI211_X1 U19481 ( .C1(n18076), .C2(n12232), .A(n17533), .B(n17710), .ZN(
        n17534) );
  AOI21_X1 U19482 ( .B1(n17715), .B2(n18091), .A(n17534), .ZN(n17535) );
  OAI211_X1 U19483 ( .C1(n18106), .C2(n17718), .A(n17536), .B(n17535), .ZN(
        P2_U2991) );
  INV_X1 U19484 ( .A(n17537), .ZN(n17539) );
  OAI21_X1 U19485 ( .B1(n17539), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n17538), .ZN(n17731) );
  OAI21_X1 U19486 ( .B1(n17540), .B2(n17542), .A(n17541), .ZN(n17729) );
  NOR2_X1 U19487 ( .A1(n19380), .A2(n18195), .ZN(n17722) );
  NOR2_X1 U19488 ( .A1(n18112), .A2(n17543), .ZN(n17544) );
  AOI211_X1 U19489 ( .C1(n18102), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n17722), .B(n17544), .ZN(n17545) );
  OAI21_X1 U19490 ( .B1(n17719), .B2(n18105), .A(n17545), .ZN(n17546) );
  AOI21_X1 U19491 ( .B1(n17729), .B2(n18079), .A(n17546), .ZN(n17547) );
  OAI21_X1 U19492 ( .B1(n17731), .B2(n18103), .A(n17547), .ZN(P2_U2992) );
  XNOR2_X1 U19493 ( .A(n17548), .B(n17550), .ZN(n17752) );
  AOI21_X1 U19494 ( .B1(n17550), .B2(n17556), .A(n17549), .ZN(n17750) );
  NAND2_X1 U19495 ( .A1(n19273), .A2(n18091), .ZN(n17553) );
  NOR2_X1 U19496 ( .A1(n19380), .A2(n17551), .ZN(n17745) );
  AOI21_X1 U19497 ( .B1(n18102), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n17745), .ZN(n17552) );
  OAI211_X1 U19498 ( .C1(n18112), .C2(n19281), .A(n17553), .B(n17552), .ZN(
        n17554) );
  AOI21_X1 U19499 ( .B1(n17750), .B2(n18095), .A(n17554), .ZN(n17555) );
  OAI21_X1 U19500 ( .B1(n17752), .B2(n18106), .A(n17555), .ZN(P2_U2994) );
  OAI21_X1 U19501 ( .B1(n17575), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n17556), .ZN(n17766) );
  NAND2_X1 U19502 ( .A1(n18070), .A2(n19264), .ZN(n17557) );
  NAND2_X1 U19503 ( .A1(n19407), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n17755) );
  OAI211_X1 U19504 ( .C1(n18076), .C2(n17558), .A(n17557), .B(n17755), .ZN(
        n17565) );
  NAND2_X1 U19505 ( .A1(n17559), .A2(n17569), .ZN(n17563) );
  NAND2_X1 U19506 ( .A1(n17561), .A2(n17560), .ZN(n17562) );
  XNOR2_X1 U19507 ( .A(n17563), .B(n17562), .ZN(n17753) );
  NOR2_X1 U19508 ( .A1(n17753), .A2(n18106), .ZN(n17564) );
  AOI211_X1 U19509 ( .C1(n18091), .C2(n19266), .A(n17565), .B(n17564), .ZN(
        n17566) );
  OAI21_X1 U19510 ( .B1(n18103), .B2(n17766), .A(n17566), .ZN(P2_U2995) );
  NAND2_X1 U19511 ( .A1(n17569), .A2(n17568), .ZN(n17570) );
  XNOR2_X1 U19512 ( .A(n17567), .B(n17570), .ZN(n17780) );
  NOR2_X1 U19513 ( .A1(n19380), .A2(n17571), .ZN(n17771) );
  AOI21_X1 U19514 ( .B1(n18102), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n17771), .ZN(n17572) );
  OAI21_X1 U19515 ( .B1(n18112), .B2(n19248), .A(n17572), .ZN(n17573) );
  AOI21_X1 U19516 ( .B1(n19253), .B2(n18091), .A(n17573), .ZN(n17578) );
  INV_X1 U19517 ( .A(n17593), .ZN(n17574) );
  AOI21_X1 U19518 ( .B1(n17574), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17576) );
  NOR2_X1 U19519 ( .A1(n17576), .A2(n17575), .ZN(n17777) );
  NAND2_X1 U19520 ( .A1(n17777), .A2(n18095), .ZN(n17577) );
  OAI211_X1 U19521 ( .C1(n17780), .C2(n18106), .A(n17578), .B(n17577), .ZN(
        P2_U2996) );
  XNOR2_X1 U19522 ( .A(n17593), .B(n17794), .ZN(n17590) );
  NAND2_X1 U19523 ( .A1(n17580), .A2(n17579), .ZN(n17584) );
  NOR2_X1 U19524 ( .A1(n17582), .A2(n17581), .ZN(n17583) );
  XOR2_X1 U19525 ( .A(n17584), .B(n17583), .Z(n17785) );
  NOR2_X1 U19526 ( .A1(n19380), .A2(n17585), .ZN(n17781) );
  AOI21_X1 U19527 ( .B1(n18102), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n17781), .ZN(n17587) );
  NAND2_X1 U19528 ( .A1(n18070), .A2(n19236), .ZN(n17586) );
  OAI211_X1 U19529 ( .C1(n19242), .C2(n18105), .A(n17587), .B(n17586), .ZN(
        n17588) );
  AOI21_X1 U19530 ( .B1(n17785), .B2(n18079), .A(n17588), .ZN(n17589) );
  OAI21_X1 U19531 ( .B1(n18103), .B2(n17590), .A(n17589), .ZN(P2_U2997) );
  XNOR2_X1 U19532 ( .A(n17592), .B(n17591), .ZN(n17802) );
  INV_X1 U19533 ( .A(n17802), .ZN(n17598) );
  OAI211_X1 U19534 ( .C1(n17605), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n18095), .B(n17593), .ZN(n17597) );
  INV_X1 U19535 ( .A(n17799), .ZN(n19229) );
  AOI22_X1 U19536 ( .A1(n18102), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n19407), .ZN(n17594) );
  OAI21_X1 U19537 ( .B1(n18112), .B2(n19227), .A(n17594), .ZN(n17595) );
  AOI21_X1 U19538 ( .B1(n19229), .B2(n18091), .A(n17595), .ZN(n17596) );
  OAI211_X1 U19539 ( .C1(n17598), .C2(n18106), .A(n17597), .B(n17596), .ZN(
        P2_U2998) );
  NAND2_X1 U19540 ( .A1(n17600), .A2(n17599), .ZN(n17604) );
  NAND2_X1 U19541 ( .A1(n17601), .A2(n17613), .ZN(n17825) );
  NAND2_X1 U19542 ( .A1(n17828), .A2(n17823), .ZN(n17603) );
  XOR2_X1 U19543 ( .A(n17604), .B(n17603), .Z(n17819) );
  AOI21_X1 U19544 ( .B1(n17815), .B2(n12764), .A(n17605), .ZN(n17808) );
  NAND2_X1 U19545 ( .A1(n17808), .A2(n18095), .ZN(n17610) );
  INV_X1 U19546 ( .A(n17606), .ZN(n19219) );
  NOR2_X1 U19547 ( .A1(n19380), .A2(n18193), .ZN(n17810) );
  AOI21_X1 U19548 ( .B1(n18102), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n17810), .ZN(n17607) );
  OAI21_X1 U19549 ( .B1(n18112), .B2(n19219), .A(n17607), .ZN(n17608) );
  AOI21_X1 U19550 ( .B1(n17811), .B2(n18091), .A(n17608), .ZN(n17609) );
  OAI211_X1 U19551 ( .C1(n17819), .C2(n18106), .A(n17610), .B(n17609), .ZN(
        P2_U2999) );
  NAND2_X1 U19552 ( .A1(n17613), .A2(n17612), .ZN(n17614) );
  XNOR2_X1 U19553 ( .A(n17611), .B(n17614), .ZN(n17849) );
  NAND2_X1 U19554 ( .A1(n17615), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17883) );
  NAND2_X1 U19555 ( .A1(n17623), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18094) );
  AND2_X1 U19556 ( .A1(n17615), .A2(n17830), .ZN(n17820) );
  AOI21_X1 U19557 ( .B1(n18094), .B2(n17842), .A(n17820), .ZN(n17839) );
  NAND2_X1 U19558 ( .A1(n17839), .A2(n18095), .ZN(n17621) );
  NAND2_X1 U19559 ( .A1(n19407), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n17840) );
  OAI21_X1 U19560 ( .B1(n18076), .B2(n17616), .A(n17840), .ZN(n17619) );
  NOR2_X1 U19561 ( .A1(n17617), .A2(n18105), .ZN(n17618) );
  AOI211_X1 U19562 ( .C1(n18070), .C2(n19193), .A(n17619), .B(n17618), .ZN(
        n17620) );
  OAI211_X1 U19563 ( .C1(n18106), .C2(n17849), .A(n17621), .B(n17620), .ZN(
        P2_U3001) );
  INV_X1 U19564 ( .A(n17622), .ZN(n17864) );
  INV_X1 U19565 ( .A(n17623), .ZN(n18092) );
  OAI21_X1 U19566 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n17864), .A(
        n18092), .ZN(n17863) );
  NOR2_X1 U19567 ( .A1(n19380), .A2(n17624), .ZN(n17854) );
  INV_X1 U19568 ( .A(n17625), .ZN(n19186) );
  OAI22_X1 U19569 ( .A1(n19177), .A2(n18076), .B1(n18112), .B2(n19186), .ZN(
        n17626) );
  AOI211_X1 U19570 ( .C1(n18091), .C2(n19173), .A(n17854), .B(n17626), .ZN(
        n17633) );
  NOR2_X1 U19571 ( .A1(n17628), .A2(n17627), .ZN(n18083) );
  INV_X1 U19572 ( .A(n17630), .ZN(n17631) );
  NAND2_X1 U19573 ( .A1(n17629), .A2(n17631), .ZN(n18084) );
  XOR2_X1 U19574 ( .A(n18083), .B(n18084), .Z(n17861) );
  NAND2_X1 U19575 ( .A1(n17861), .A2(n18079), .ZN(n17632) );
  OAI211_X1 U19576 ( .C1(n17863), .C2(n18103), .A(n17633), .B(n17632), .ZN(
        P2_U3003) );
  INV_X1 U19577 ( .A(n18063), .ZN(n17636) );
  NOR2_X1 U19578 ( .A1(n17636), .A2(n17635), .ZN(n17637) );
  XNOR2_X1 U19579 ( .A(n17634), .B(n17637), .ZN(n17910) );
  OR2_X1 U19580 ( .A1(n17639), .A2(n17638), .ZN(n17899) );
  NAND3_X1 U19581 ( .A1(n17899), .A2(n18095), .A3(n17898), .ZN(n17646) );
  INV_X1 U19582 ( .A(n19140), .ZN(n17640) );
  NOR2_X1 U19583 ( .A1(n18112), .A2(n17640), .ZN(n17643) );
  OAI22_X1 U19584 ( .A1(n17641), .A2(n18076), .B1(n11757), .B2(n19258), .ZN(
        n17642) );
  AOI211_X1 U19585 ( .C1(n18091), .C2(n17644), .A(n17643), .B(n17642), .ZN(
        n17645) );
  OAI211_X1 U19586 ( .C1(n17910), .C2(n18106), .A(n17646), .B(n17645), .ZN(
        P2_U3007) );
  INV_X1 U19587 ( .A(n19331), .ZN(n17656) );
  NOR2_X1 U19588 ( .A1(n17928), .A2(n19337), .ZN(n17654) );
  XNOR2_X1 U19589 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17648) );
  OAI21_X1 U19590 ( .B1(n17649), .B2(n17648), .A(n17647), .ZN(n17652) );
  OR2_X1 U19591 ( .A1(n17652), .A2(n17651), .ZN(n17653) );
  OAI21_X1 U19592 ( .B1(n17659), .B2(n19388), .A(n17658), .ZN(P2_U3017) );
  OAI21_X1 U19593 ( .B1(n17928), .B2(n17661), .A(n17660), .ZN(n17662) );
  AOI21_X1 U19594 ( .B1(n17663), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n17662), .ZN(n17665) );
  OAI211_X1 U19595 ( .C1(n17666), .C2(n19416), .A(n17665), .B(n17664), .ZN(
        n17667) );
  AOI21_X1 U19596 ( .B1(n17668), .B2(n19420), .A(n17667), .ZN(n17669) );
  OAI21_X1 U19597 ( .B1(n17670), .B2(n19388), .A(n17669), .ZN(P2_U3019) );
  NOR2_X1 U19598 ( .A1(n17671), .A2(n17687), .ZN(n17672) );
  AOI211_X1 U19599 ( .C1(n19408), .C2(n19296), .A(n17673), .B(n17672), .ZN(
        n17676) );
  OAI211_X1 U19600 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n17692), .B(n17674), .ZN(
        n17675) );
  OAI211_X1 U19601 ( .C1(n17677), .C2(n19416), .A(n17676), .B(n17675), .ZN(
        n17678) );
  AOI21_X1 U19602 ( .B1(n17679), .B2(n19419), .A(n17678), .ZN(n17680) );
  OAI21_X1 U19603 ( .B1(n19375), .B2(n17681), .A(n17680), .ZN(P2_U3020) );
  NAND3_X1 U19604 ( .A1(n17683), .A2(n19420), .A3(n17682), .ZN(n17694) );
  NAND2_X1 U19605 ( .A1(n19408), .A2(n17684), .ZN(n17686) );
  OAI211_X1 U19606 ( .C1(n17687), .C2(n17691), .A(n17686), .B(n17685), .ZN(
        n17690) );
  NOR2_X1 U19607 ( .A1(n17688), .A2(n19416), .ZN(n17689) );
  AOI211_X1 U19608 ( .C1(n17692), .C2(n17691), .A(n17690), .B(n17689), .ZN(
        n17693) );
  OAI211_X1 U19609 ( .C1(n17695), .C2(n19388), .A(n17694), .B(n17693), .ZN(
        P2_U3021) );
  INV_X1 U19610 ( .A(n19284), .ZN(n17697) );
  AOI21_X1 U19611 ( .B1(n19408), .B2(n17697), .A(n17696), .ZN(n17701) );
  NOR2_X1 U19612 ( .A1(n17727), .A2(n12694), .ZN(n17699) );
  OAI21_X1 U19613 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17699), .A(
        n17698), .ZN(n17700) );
  OAI211_X1 U19614 ( .C1(n19285), .C2(n19416), .A(n17701), .B(n17700), .ZN(
        n17702) );
  AOI21_X1 U19615 ( .B1(n17703), .B2(n19419), .A(n17702), .ZN(n17704) );
  OAI21_X1 U19616 ( .B1(n17705), .B2(n19375), .A(n17704), .ZN(P2_U3022) );
  NAND2_X1 U19617 ( .A1(n17706), .A2(n19420), .ZN(n17717) );
  AOI211_X1 U19618 ( .C1(n17709), .C2(n17708), .A(n17707), .B(n17727), .ZN(
        n17714) );
  NAND2_X1 U19619 ( .A1(n17724), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17711) );
  OAI211_X1 U19620 ( .C1(n17928), .C2(n17712), .A(n17711), .B(n17710), .ZN(
        n17713) );
  AOI211_X1 U19621 ( .C1(n17715), .C2(n19398), .A(n17714), .B(n17713), .ZN(
        n17716) );
  OAI211_X1 U19622 ( .C1(n17718), .C2(n19388), .A(n17717), .B(n17716), .ZN(
        P2_U3023) );
  INV_X1 U19623 ( .A(n17719), .ZN(n17723) );
  NOR2_X1 U19624 ( .A1(n17928), .A2(n17720), .ZN(n17721) );
  AOI211_X1 U19625 ( .C1(n17723), .C2(n19398), .A(n17722), .B(n17721), .ZN(
        n17726) );
  NAND2_X1 U19626 ( .A1(n17724), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17725) );
  OAI211_X1 U19627 ( .C1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17727), .A(
        n17726), .B(n17725), .ZN(n17728) );
  AOI21_X1 U19628 ( .B1(n17729), .B2(n19419), .A(n17728), .ZN(n17730) );
  OAI21_X1 U19629 ( .B1(n17731), .B2(n19375), .A(n17730), .ZN(P2_U3024) );
  NOR2_X1 U19630 ( .A1(n17757), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17775) );
  AND2_X1 U19631 ( .A1(n17732), .A2(n17734), .ZN(n17733) );
  OAI22_X1 U19632 ( .A1(n17734), .A2(n17923), .B1(n17787), .B2(n17733), .ZN(
        n17736) );
  OR2_X1 U19633 ( .A1(n17736), .A2(n17735), .ZN(n17789) );
  INV_X1 U19634 ( .A(n17789), .ZN(n17737) );
  OAI21_X1 U19635 ( .B1(n17738), .B2(n17791), .A(n17737), .ZN(n17776) );
  NOR2_X1 U19636 ( .A1(n17775), .A2(n17776), .ZN(n17762) );
  OAI21_X1 U19637 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17757), .A(
        n17762), .ZN(n17739) );
  NAND2_X1 U19638 ( .A1(n17739), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17747) );
  INV_X1 U19639 ( .A(n17740), .ZN(n17741) );
  OAI21_X1 U19640 ( .B1(n17743), .B2(n17742), .A(n17741), .ZN(n20225) );
  NOR2_X1 U19641 ( .A1(n20225), .A2(n17928), .ZN(n17744) );
  AOI211_X1 U19642 ( .C1(n19273), .C2(n19398), .A(n17745), .B(n17744), .ZN(
        n17746) );
  OAI211_X1 U19643 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n17748), .A(
        n17747), .B(n17746), .ZN(n17749) );
  AOI21_X1 U19644 ( .B1(n17750), .B2(n19420), .A(n17749), .ZN(n17751) );
  OAI21_X1 U19645 ( .B1(n17752), .B2(n19388), .A(n17751), .ZN(P2_U3026) );
  INV_X1 U19646 ( .A(n17753), .ZN(n17764) );
  INV_X1 U19647 ( .A(n17754), .ZN(n19270) );
  OAI21_X1 U19648 ( .B1(n19270), .B2(n17928), .A(n17755), .ZN(n17759) );
  NOR3_X1 U19649 ( .A1(n17757), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n17756), .ZN(n17758) );
  AOI211_X1 U19650 ( .C1(n19266), .C2(n19398), .A(n17759), .B(n17758), .ZN(
        n17760) );
  OAI21_X1 U19651 ( .B1(n17762), .B2(n17761), .A(n17760), .ZN(n17763) );
  AOI21_X1 U19652 ( .B1(n17764), .B2(n19419), .A(n17763), .ZN(n17765) );
  OAI21_X1 U19653 ( .B1(n19375), .B2(n17766), .A(n17765), .ZN(P2_U3027) );
  NAND2_X1 U19654 ( .A1(n17768), .A2(n17767), .ZN(n17769) );
  AND2_X1 U19655 ( .A1(n17770), .A2(n17769), .ZN(n20320) );
  AOI21_X1 U19656 ( .B1(n19408), .B2(n20320), .A(n17771), .ZN(n17772) );
  OAI21_X1 U19657 ( .B1(n17773), .B2(n19416), .A(n17772), .ZN(n17774) );
  AOI211_X1 U19658 ( .C1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n17776), .A(
        n17775), .B(n17774), .ZN(n17779) );
  NAND2_X1 U19659 ( .A1(n17777), .A2(n19420), .ZN(n17778) );
  OAI211_X1 U19660 ( .C1(n17780), .C2(n19388), .A(n17779), .B(n17778), .ZN(
        P2_U3028) );
  NOR2_X1 U19661 ( .A1(n17928), .A2(n19241), .ZN(n17784) );
  INV_X1 U19662 ( .A(n17781), .ZN(n17782) );
  OAI21_X1 U19663 ( .B1(n19242), .B2(n19416), .A(n17782), .ZN(n17783) );
  AOI211_X1 U19664 ( .C1(n17785), .C2(n19419), .A(n17784), .B(n17783), .ZN(
        n17797) );
  NOR2_X1 U19665 ( .A1(n17787), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17788) );
  NOR2_X1 U19666 ( .A1(n17789), .A2(n17788), .ZN(n17813) );
  NAND2_X1 U19667 ( .A1(n17790), .A2(n17813), .ZN(n17798) );
  AOI21_X1 U19668 ( .B1(n17791), .B2(n19375), .A(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17792) );
  OAI21_X1 U19669 ( .B1(n17798), .B2(n17792), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17796) );
  NAND3_X1 U19670 ( .A1(n17803), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n17794), .ZN(n17795) );
  NAND3_X1 U19671 ( .A1(n17797), .A2(n17796), .A3(n17795), .ZN(P2_U3029) );
  INV_X1 U19672 ( .A(n17798), .ZN(n17807) );
  NOR2_X1 U19673 ( .A1(n17928), .A2(n19233), .ZN(n17801) );
  OAI22_X1 U19674 ( .A1(n17799), .A2(n19416), .B1(n11789), .B2(n19380), .ZN(
        n17800) );
  AOI211_X1 U19675 ( .C1(n17802), .C2(n19419), .A(n17801), .B(n17800), .ZN(
        n17805) );
  NAND2_X1 U19676 ( .A1(n17803), .A2(n17806), .ZN(n17804) );
  OAI211_X1 U19677 ( .C1(n17807), .C2(n17806), .A(n17805), .B(n17804), .ZN(
        P2_U3030) );
  NAND2_X1 U19678 ( .A1(n17808), .A2(n19420), .ZN(n17818) );
  NOR2_X1 U19679 ( .A1(n17928), .A2(n19223), .ZN(n17809) );
  AOI211_X1 U19680 ( .C1(n17811), .C2(n19398), .A(n17810), .B(n17809), .ZN(
        n17812) );
  OAI21_X1 U19681 ( .B1(n17813), .B2(n17815), .A(n17812), .ZN(n17814) );
  AOI21_X1 U19682 ( .B1(n17816), .B2(n17815), .A(n17814), .ZN(n17817) );
  OAI211_X1 U19683 ( .C1(n17819), .C2(n19388), .A(n17818), .B(n17817), .ZN(
        P2_U3031) );
  OR2_X1 U19684 ( .A1(n17820), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17821) );
  NAND2_X1 U19685 ( .A1(n17821), .A2(n12764), .ZN(n18104) );
  INV_X1 U19686 ( .A(n17823), .ZN(n17827) );
  NAND2_X1 U19687 ( .A1(n17823), .A2(n17822), .ZN(n17824) );
  NAND2_X1 U19688 ( .A1(n17825), .A2(n17824), .ZN(n17826) );
  OAI21_X1 U19689 ( .B1(n17828), .B2(n17827), .A(n17826), .ZN(n18107) );
  NAND2_X1 U19690 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19407), .ZN(n17829) );
  OAI21_X1 U19691 ( .B1(n19206), .B2(n19416), .A(n17829), .ZN(n17833) );
  INV_X1 U19692 ( .A(n17896), .ZN(n17852) );
  INV_X1 U19693 ( .A(n17830), .ZN(n17831) );
  NOR3_X1 U19694 ( .A1(n17852), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n17831), .ZN(n17832) );
  AOI211_X1 U19695 ( .C1(n19408), .C2(n19207), .A(n17833), .B(n17832), .ZN(
        n17836) );
  NOR3_X1 U19696 ( .A1(n17852), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n19379), .ZN(n19381) );
  AOI211_X1 U19697 ( .C1(n19379), .C2(n19378), .A(n19377), .B(n19381), .ZN(
        n17843) );
  INV_X1 U19698 ( .A(n17843), .ZN(n17834) );
  NOR3_X1 U19699 ( .A1(n17852), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n19379), .ZN(n17846) );
  OAI21_X1 U19700 ( .B1(n17834), .B2(n17846), .A(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17835) );
  OAI211_X1 U19701 ( .C1(n18107), .C2(n19388), .A(n17836), .B(n17835), .ZN(
        n17837) );
  INV_X1 U19702 ( .A(n17837), .ZN(n17838) );
  OAI21_X1 U19703 ( .B1(n19375), .B2(n18104), .A(n17838), .ZN(P2_U3032) );
  NAND2_X1 U19704 ( .A1(n17839), .A2(n19420), .ZN(n17848) );
  NAND2_X1 U19705 ( .A1(n19398), .A2(n19195), .ZN(n17841) );
  OAI211_X1 U19706 ( .C1(n17928), .C2(n19199), .A(n17841), .B(n17840), .ZN(
        n17845) );
  NOR2_X1 U19707 ( .A1(n17843), .A2(n17842), .ZN(n17844) );
  AOI211_X1 U19708 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n17846), .A(
        n17845), .B(n17844), .ZN(n17847) );
  OAI211_X1 U19709 ( .C1(n17849), .C2(n19388), .A(n17848), .B(n17847), .ZN(
        P2_U3033) );
  NOR2_X1 U19710 ( .A1(n17895), .A2(n19377), .ZN(n17850) );
  NOR2_X1 U19711 ( .A1(n17851), .A2(n17850), .ZN(n17868) );
  NOR3_X1 U19712 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17895), .A3(
        n17852), .ZN(n17867) );
  OAI21_X1 U19713 ( .B1(n17868), .B2(n17867), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17859) );
  NAND4_X1 U19714 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n17896), .A4(n17853), .ZN(
        n17856) );
  INV_X1 U19715 ( .A(n17854), .ZN(n17855) );
  OAI211_X1 U19716 ( .C1(n17928), .C2(n19176), .A(n17856), .B(n17855), .ZN(
        n17857) );
  AOI21_X1 U19717 ( .B1(n19398), .B2(n19173), .A(n17857), .ZN(n17858) );
  NAND2_X1 U19718 ( .A1(n17859), .A2(n17858), .ZN(n17860) );
  AOI21_X1 U19719 ( .B1(n17861), .B2(n19419), .A(n17860), .ZN(n17862) );
  OAI21_X1 U19720 ( .B1(n17863), .B2(n19375), .A(n17862), .ZN(P2_U3035) );
  AOI21_X1 U19721 ( .B1(n17865), .B2(n17883), .A(n17864), .ZN(n18078) );
  NAND2_X1 U19722 ( .A1(n18078), .A2(n19420), .ZN(n17882) );
  NOR2_X1 U19723 ( .A1(n11767), .A2(n19380), .ZN(n17866) );
  AOI211_X1 U19724 ( .C1(n17868), .C2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17867), .B(n17866), .ZN(n17881) );
  OAI22_X1 U19725 ( .A1(n19416), .A2(n17869), .B1(n17928), .B2(n19172), .ZN(
        n17870) );
  INV_X1 U19726 ( .A(n17870), .ZN(n17880) );
  NAND2_X1 U19727 ( .A1(n17871), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17872) );
  NAND2_X1 U19728 ( .A1(n17872), .A2(n18064), .ZN(n17874) );
  OR2_X1 U19729 ( .A1(n17871), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17873) );
  NAND2_X1 U19730 ( .A1(n17890), .A2(n17887), .ZN(n17892) );
  NAND2_X1 U19731 ( .A1(n17892), .A2(n17888), .ZN(n17878) );
  NAND2_X1 U19732 ( .A1(n17876), .A2(n17875), .ZN(n17877) );
  XNOR2_X1 U19733 ( .A(n17878), .B(n17877), .ZN(n18080) );
  NAND2_X1 U19734 ( .A1(n18080), .A2(n19419), .ZN(n17879) );
  NAND4_X1 U19735 ( .A1(n17882), .A2(n17881), .A3(n17880), .A4(n17879), .ZN(
        P2_U3036) );
  OAI21_X1 U19736 ( .B1(n17615), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17883), .ZN(n18072) );
  NAND2_X1 U19737 ( .A1(n19377), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17886) );
  NOR2_X1 U19738 ( .A1(n11763), .A2(n19380), .ZN(n17884) );
  AOI21_X1 U19739 ( .B1(n19398), .B2(n19157), .A(n17884), .ZN(n17885) );
  OAI211_X1 U19740 ( .C1(n17928), .C2(n19161), .A(n17886), .B(n17885), .ZN(
        n17894) );
  INV_X1 U19741 ( .A(n17888), .ZN(n17891) );
  AND2_X1 U19742 ( .A1(n17888), .A2(n17887), .ZN(n17889) );
  OAI22_X1 U19743 ( .A1(n17892), .A2(n17891), .B1(n17890), .B2(n17889), .ZN(
        n18071) );
  NOR2_X1 U19744 ( .A1(n18071), .A2(n19388), .ZN(n17893) );
  AOI211_X1 U19745 ( .C1(n17896), .C2(n17895), .A(n17894), .B(n17893), .ZN(
        n17897) );
  OAI21_X1 U19746 ( .B1(n19375), .B2(n18072), .A(n17897), .ZN(P2_U3037) );
  NAND3_X1 U19747 ( .A1(n17899), .A2(n19420), .A3(n17898), .ZN(n17909) );
  INV_X1 U19748 ( .A(n17900), .ZN(n17903) );
  AOI21_X1 U19749 ( .B1(n17902), .B2(n17901), .A(n19367), .ZN(n17922) );
  OAI21_X1 U19750 ( .B1(n17903), .B2(n17923), .A(n17922), .ZN(n19396) );
  AND2_X1 U19751 ( .A1(n17903), .A2(n19411), .ZN(n19402) );
  AOI22_X1 U19752 ( .A1(n19407), .A2(P2_REIP_REG_7__SCAN_IN), .B1(n19402), 
        .B2(n17904), .ZN(n17905) );
  OAI21_X1 U19753 ( .B1(n19416), .B2(n19144), .A(n17905), .ZN(n17907) );
  NOR2_X1 U19754 ( .A1(n19145), .A2(n17928), .ZN(n17906) );
  AOI211_X1 U19755 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n19396), .A(
        n17907), .B(n17906), .ZN(n17908) );
  OAI211_X1 U19756 ( .C1(n17910), .C2(n19388), .A(n17909), .B(n17908), .ZN(
        P2_U3039) );
  OAI21_X1 U19757 ( .B1(n17912), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n17911), .ZN(n18055) );
  OR2_X1 U19758 ( .A1(n17915), .A2(n17914), .ZN(n17916) );
  NAND2_X1 U19759 ( .A1(n17913), .A2(n17916), .ZN(n18054) );
  INV_X1 U19760 ( .A(n18054), .ZN(n17930) );
  NOR2_X1 U19761 ( .A1(n11754), .A2(n19380), .ZN(n17920) );
  INV_X1 U19762 ( .A(n19411), .ZN(n17918) );
  INV_X1 U19763 ( .A(n17924), .ZN(n17917) );
  NOR3_X1 U19764 ( .A1(n17918), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n17917), .ZN(n17919) );
  AOI211_X1 U19765 ( .C1(n19398), .C2(n17921), .A(n17920), .B(n17919), .ZN(
        n17927) );
  OAI21_X1 U19766 ( .B1(n17924), .B2(n17923), .A(n17922), .ZN(n17925) );
  NAND2_X1 U19767 ( .A1(n17925), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17926) );
  OAI211_X1 U19768 ( .C1(n19134), .C2(n17928), .A(n17927), .B(n17926), .ZN(
        n17929) );
  AOI21_X1 U19769 ( .B1(n17930), .B2(n19419), .A(n17929), .ZN(n17931) );
  OAI21_X1 U19770 ( .B1(n18055), .B2(n19375), .A(n17931), .ZN(P2_U3040) );
  INV_X1 U19771 ( .A(n19362), .ZN(n19425) );
  OAI22_X1 U19772 ( .A1(n20058), .A2(n19435), .B1(n17932), .B2(n19425), .ZN(
        n17933) );
  MUX2_X1 U19773 ( .A(n17933), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n19358), .Z(P2_U3596) );
  NAND2_X1 U19774 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19503) );
  NAND2_X1 U19775 ( .A1(n18933), .A2(n20833), .ZN(n17937) );
  INV_X1 U19776 ( .A(n17937), .ZN(n17936) );
  NAND2_X1 U19777 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19530), .ZN(n19497) );
  NOR2_X1 U19778 ( .A1(n18538), .A2(n17934), .ZN(n18573) );
  INV_X1 U19779 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n21965) );
  OAI221_X1 U19780 ( .B1(n17935), .B2(n18573), .C1(n17935), .C2(n21965), .A(
        n19686), .ZN(n18979) );
  NAND2_X1 U19781 ( .A1(n19497), .A2(n18979), .ZN(n18981) );
  AOI221_X1 U19782 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19503), .C1(n17936), 
        .C2(n19503), .A(n18981), .ZN(n18977) );
  INV_X1 U19783 ( .A(n19526), .ZN(n18980) );
  OAI21_X1 U19784 ( .B1(n19530), .B2(n21949), .A(n17937), .ZN(n18978) );
  OAI221_X1 U19785 ( .B1(n18980), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18980), .C2(n18978), .A(n18979), .ZN(n18975) );
  AOI22_X1 U19786 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18977), .B1(
        n18975), .B2(n19523), .ZN(P3_U2865) );
  NAND4_X1 U19787 ( .A1(n22107), .A2(n17940), .A3(n17939), .A4(n17938), .ZN(
        n17941) );
  OAI21_X1 U19788 ( .B1(n17943), .B2(n17942), .A(n17941), .ZN(P1_U3468) );
  INV_X1 U19789 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17945) );
  INV_X1 U19790 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n22364) );
  OAI21_X1 U19791 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n22364), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n19048) );
  NAND2_X1 U19792 ( .A1(n19068), .A2(n19048), .ZN(n17947) );
  INV_X1 U19793 ( .A(n17947), .ZN(n22318) );
  INV_X1 U19794 ( .A(n22318), .ZN(n17946) );
  NAND2_X1 U19795 ( .A1(n22356), .A2(n22364), .ZN(n22319) );
  AOI21_X1 U19796 ( .B1(n17944), .B2(n22319), .A(n17946), .ZN(n22314) );
  AOI21_X1 U19797 ( .B1(n17945), .B2(n17946), .A(n22314), .ZN(P3_U3280) );
  AND2_X1 U19798 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n17946), .ZN(P3_U3028) );
  AND2_X1 U19799 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n17946), .ZN(P3_U3027) );
  AND2_X1 U19800 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n17946), .ZN(P3_U3026) );
  AND2_X1 U19801 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n17946), .ZN(P3_U3025) );
  AND2_X1 U19802 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n17946), .ZN(P3_U3024) );
  AND2_X1 U19803 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n17946), .ZN(P3_U3023) );
  AND2_X1 U19804 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n17946), .ZN(P3_U3022) );
  AND2_X1 U19805 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n17946), .ZN(P3_U3021) );
  AND2_X1 U19806 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n17946), .ZN(
        P3_U3020) );
  AND2_X1 U19807 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n17946), .ZN(
        P3_U3019) );
  AND2_X1 U19808 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n17946), .ZN(
        P3_U3018) );
  AND2_X1 U19809 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n17946), .ZN(
        P3_U3017) );
  AND2_X1 U19810 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n17946), .ZN(
        P3_U3016) );
  AND2_X1 U19811 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n17947), .ZN(
        P3_U3015) );
  AND2_X1 U19812 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n17947), .ZN(
        P3_U3014) );
  AND2_X1 U19813 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n17947), .ZN(
        P3_U3013) );
  AND2_X1 U19814 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n17947), .ZN(
        P3_U3012) );
  AND2_X1 U19815 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n17947), .ZN(
        P3_U3011) );
  AND2_X1 U19816 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n17947), .ZN(
        P3_U3010) );
  AND2_X1 U19817 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n17947), .ZN(
        P3_U3009) );
  AND2_X1 U19818 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n17947), .ZN(
        P3_U3008) );
  AND2_X1 U19819 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n17946), .ZN(
        P3_U3007) );
  AND2_X1 U19820 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n17946), .ZN(
        P3_U3006) );
  AND2_X1 U19821 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n17946), .ZN(
        P3_U3005) );
  AND2_X1 U19822 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n17946), .ZN(
        P3_U3004) );
  AND2_X1 U19823 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n17946), .ZN(
        P3_U3003) );
  AND2_X1 U19824 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n17946), .ZN(
        P3_U3002) );
  AND2_X1 U19825 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n17946), .ZN(
        P3_U3001) );
  AND2_X1 U19826 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n17946), .ZN(
        P3_U3000) );
  AND2_X1 U19827 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n17947), .ZN(
        P3_U2999) );
  AOI21_X1 U19828 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n17949)
         );
  AOI211_X1 U19829 ( .C1(n18933), .C2(n17949), .A(n21946), .B(n17948), .ZN(
        P3_U2998) );
  NOR2_X1 U19830 ( .A1(n17950), .A2(n18979), .ZN(P3_U2867) );
  INV_X1 U19832 ( .A(n20842), .ZN(n18568) );
  AND2_X1 U19833 ( .A1(n19037), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U19834 ( .A1(n18571), .A2(n20899), .ZN(n17955) );
  OAI22_X1 U19835 ( .A1(P3_READREQUEST_REG_SCAN_IN), .A2(n17955), .B1(n20835), 
        .B2(n20899), .ZN(n17954) );
  INV_X1 U19836 ( .A(n17954), .ZN(P3_U3298) );
  NOR2_X1 U19837 ( .A1(n19027), .A2(n20899), .ZN(n21327) );
  NOR2_X1 U19838 ( .A1(P3_MEMORYFETCH_REG_SCAN_IN), .A2(n17955), .ZN(n17956)
         );
  NOR2_X1 U19839 ( .A1(n21327), .A2(n17956), .ZN(P3_U3299) );
  AND2_X1 U19840 ( .A1(n22354), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n22344) );
  AOI21_X1 U19841 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n22344), .A(n17957), 
        .ZN(n17959) );
  INV_X1 U19842 ( .A(n17959), .ZN(n22313) );
  NOR2_X1 U19843 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n22339) );
  OAI21_X1 U19844 ( .B1(BS16), .B2(n22339), .A(n22313), .ZN(n22311) );
  OAI21_X1 U19845 ( .B1(n22313), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n22311), 
        .ZN(n17958) );
  INV_X1 U19846 ( .A(n17958), .ZN(P2_U3591) );
  AND2_X1 U19847 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n17959), .ZN(P2_U3208) );
  AND2_X1 U19848 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n17959), .ZN(P2_U3207) );
  INV_X1 U19849 ( .A(n22313), .ZN(n17960) );
  AND2_X1 U19850 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n17960), .ZN(P2_U3206) );
  AND2_X1 U19851 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n17959), .ZN(P2_U3205) );
  AND2_X1 U19852 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n17960), .ZN(P2_U3204) );
  AND2_X1 U19853 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n17959), .ZN(P2_U3203) );
  AND2_X1 U19854 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n17960), .ZN(P2_U3202) );
  AND2_X1 U19855 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n17960), .ZN(P2_U3201) );
  AND2_X1 U19856 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n17960), .ZN(
        P2_U3200) );
  AND2_X1 U19857 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n17960), .ZN(
        P2_U3199) );
  AND2_X1 U19858 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n17960), .ZN(
        P2_U3198) );
  AND2_X1 U19859 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n17960), .ZN(
        P2_U3197) );
  AND2_X1 U19860 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n17959), .ZN(
        P2_U3196) );
  AND2_X1 U19861 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n17959), .ZN(
        P2_U3195) );
  AND2_X1 U19862 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n17959), .ZN(
        P2_U3194) );
  AND2_X1 U19863 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n17959), .ZN(
        P2_U3193) );
  AND2_X1 U19864 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n17959), .ZN(
        P2_U3192) );
  AND2_X1 U19865 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n17959), .ZN(
        P2_U3191) );
  AND2_X1 U19866 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n17959), .ZN(
        P2_U3190) );
  AND2_X1 U19867 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n17959), .ZN(
        P2_U3189) );
  AND2_X1 U19868 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n17959), .ZN(
        P2_U3188) );
  AND2_X1 U19869 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n17959), .ZN(
        P2_U3187) );
  AND2_X1 U19870 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n17960), .ZN(
        P2_U3186) );
  AND2_X1 U19871 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n17960), .ZN(
        P2_U3185) );
  AND2_X1 U19872 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n17960), .ZN(
        P2_U3184) );
  AND2_X1 U19873 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n17960), .ZN(
        P2_U3183) );
  AND2_X1 U19874 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n17960), .ZN(
        P2_U3182) );
  AND2_X1 U19875 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n17960), .ZN(
        P2_U3181) );
  AND2_X1 U19876 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n17960), .ZN(
        P2_U3180) );
  AND2_X1 U19877 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n17960), .ZN(
        P2_U3179) );
  NAND2_X1 U19878 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19073), .ZN(n19426) );
  AOI21_X1 U19879 ( .B1(n17961), .B2(n19436), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17964) );
  AOI221_X1 U19880 ( .B1(n19426), .B2(n17964), .C1(n17963), .C2(n17964), .A(
        n17962), .ZN(P2_U3178) );
  OAI221_X1 U19881 ( .B1(n12618), .B2(n17966), .C1(n17965), .C2(n17966), .A(
        n20426), .ZN(n18133) );
  NOR2_X1 U19882 ( .A1(n17967), .A2(n18133), .ZN(P2_U3047) );
  AND2_X1 U19883 ( .A1(n18159), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U19884 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17971) );
  NOR4_X1 U19885 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17970) );
  NOR4_X1 U19886 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17969) );
  NOR4_X1 U19887 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17968) );
  NAND4_X1 U19888 ( .A1(n17971), .A2(n17970), .A3(n17969), .A4(n17968), .ZN(
        n17977) );
  NOR4_X1 U19889 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n17975) );
  AOI211_X1 U19890 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17974) );
  NOR4_X1 U19891 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17973) );
  NOR4_X1 U19892 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17972) );
  NAND4_X1 U19893 ( .A1(n17975), .A2(n17974), .A3(n17973), .A4(n17972), .ZN(
        n17976) );
  NOR2_X1 U19894 ( .A1(n17977), .A2(n17976), .ZN(n18143) );
  INV_X1 U19895 ( .A(n18143), .ZN(n18141) );
  NOR2_X1 U19896 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18141), .ZN(n18136) );
  OR3_X1 U19897 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18140) );
  INV_X1 U19898 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17978) );
  AOI22_X1 U19899 ( .A1(n18136), .A2(n18140), .B1(n18141), .B2(n17978), .ZN(
        P2_U2821) );
  INV_X1 U19900 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n17979) );
  AOI22_X1 U19901 ( .A1(n18136), .A2(n16338), .B1(n18141), .B2(n17979), .ZN(
        P2_U2820) );
  INV_X1 U19902 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17980) );
  NOR2_X1 U19903 ( .A1(n12943), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n22805) );
  AND2_X1 U19904 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n22323), .ZN(n18026) );
  NOR2_X1 U19905 ( .A1(n22805), .A2(n18026), .ZN(n22306) );
  INV_X1 U19906 ( .A(n22306), .ZN(n22308) );
  OAI221_X1 U19907 ( .B1(n12943), .B2(BS16), .C1(n22329), .C2(BS16), .A(n22306), .ZN(n22304) );
  INV_X1 U19908 ( .A(n22304), .ZN(n22307) );
  AOI21_X1 U19909 ( .B1(n17980), .B2(n22308), .A(n22307), .ZN(P1_U3464) );
  AND2_X1 U19910 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n22308), .ZN(P1_U3193) );
  AND2_X1 U19911 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n22308), .ZN(P1_U3192) );
  AND2_X1 U19912 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n22308), .ZN(P1_U3191) );
  AND2_X1 U19913 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n22308), .ZN(P1_U3190) );
  AND2_X1 U19914 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n22308), .ZN(P1_U3189) );
  AND2_X1 U19915 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n22308), .ZN(P1_U3188) );
  AND2_X1 U19916 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n22308), .ZN(P1_U3187) );
  AND2_X1 U19917 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n22308), .ZN(P1_U3186) );
  AND2_X1 U19918 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n22308), .ZN(
        P1_U3185) );
  AND2_X1 U19919 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n22308), .ZN(
        P1_U3184) );
  AND2_X1 U19920 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n22308), .ZN(
        P1_U3183) );
  AND2_X1 U19921 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n22308), .ZN(
        P1_U3182) );
  AND2_X1 U19922 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n22308), .ZN(
        P1_U3181) );
  AND2_X1 U19923 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n22308), .ZN(
        P1_U3180) );
  AND2_X1 U19924 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n22308), .ZN(
        P1_U3179) );
  AND2_X1 U19925 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n22308), .ZN(
        P1_U3178) );
  AND2_X1 U19926 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n22308), .ZN(
        P1_U3177) );
  AND2_X1 U19927 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n22308), .ZN(
        P1_U3176) );
  AND2_X1 U19928 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n22308), .ZN(
        P1_U3175) );
  AND2_X1 U19929 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n22308), .ZN(
        P1_U3174) );
  AND2_X1 U19930 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n22308), .ZN(
        P1_U3173) );
  AND2_X1 U19931 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n22308), .ZN(
        P1_U3172) );
  AND2_X1 U19932 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n22308), .ZN(
        P1_U3171) );
  AND2_X1 U19933 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n22308), .ZN(
        P1_U3170) );
  AND2_X1 U19934 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n22308), .ZN(
        P1_U3169) );
  AND2_X1 U19935 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n22308), .ZN(
        P1_U3168) );
  AND2_X1 U19936 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n22308), .ZN(
        P1_U3167) );
  AND2_X1 U19937 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n22308), .ZN(
        P1_U3166) );
  AND2_X1 U19938 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n22308), .ZN(
        P1_U3165) );
  AND2_X1 U19939 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n22308), .ZN(
        P1_U3164) );
  NOR2_X1 U19940 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n22424), .ZN(n17984) );
  NOR3_X1 U19941 ( .A1(n21971), .A2(n22331), .A3(n17981), .ZN(n17982) );
  NAND2_X1 U19942 ( .A1(n17982), .A2(n14280), .ZN(n17983) );
  OAI221_X1 U19943 ( .B1(n17985), .B2(n17984), .C1(n17985), .C2(n22330), .A(
        n17983), .ZN(n17986) );
  INV_X1 U19944 ( .A(n17986), .ZN(n18021) );
  NAND2_X1 U19945 ( .A1(n22278), .A2(n17987), .ZN(n18015) );
  MUX2_X1 U19946 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n17988), .S(
        n17994), .Z(n18006) );
  MUX2_X1 U19947 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n17989), .S(
        n17994), .Z(n18007) );
  NAND2_X1 U19948 ( .A1(n17990), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n17991) );
  OR2_X1 U19949 ( .A1(n17992), .A2(n17991), .ZN(n17993) );
  INV_X1 U19950 ( .A(n17993), .ZN(n17998) );
  AOI22_X1 U19951 ( .A1(n17995), .A2(n17994), .B1(n22406), .B2(n17993), .ZN(
        n17997) );
  NOR2_X1 U19952 ( .A1(n18007), .A2(n18000), .ZN(n17996) );
  AOI211_X1 U19953 ( .C1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n17998), .A(
        n17997), .B(n17996), .ZN(n17999) );
  AOI21_X1 U19954 ( .B1(n18007), .B2(n18000), .A(n17999), .ZN(n18002) );
  INV_X1 U19955 ( .A(n18002), .ZN(n18004) );
  INV_X1 U19956 ( .A(n18006), .ZN(n18001) );
  AOI21_X1 U19957 ( .B1(n18002), .B2(n18001), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18003) );
  AOI21_X1 U19958 ( .B1(n18006), .B2(n18004), .A(n18003), .ZN(n18012) );
  INV_X1 U19959 ( .A(n18005), .ZN(n18010) );
  NAND2_X1 U19960 ( .A1(n18007), .A2(n18006), .ZN(n18008) );
  AND3_X1 U19961 ( .A1(n18010), .A2(n18009), .A3(n18008), .ZN(n18011) );
  OAI21_X1 U19962 ( .B1(n18012), .B2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n18011), .ZN(n18013) );
  AOI211_X1 U19963 ( .C1(n18016), .C2(n18015), .A(n18014), .B(n18013), .ZN(
        n22303) );
  NAND2_X1 U19964 ( .A1(n18021), .A2(n22303), .ZN(n18017) );
  OAI211_X1 U19965 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n22322), .A(n22293), 
        .B(n18018), .ZN(n22294) );
  AOI21_X1 U19966 ( .B1(n22322), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n18019), 
        .ZN(n18020) );
  INV_X1 U19967 ( .A(n18020), .ZN(n18022) );
  NAND2_X1 U19968 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n18021), .ZN(n22299) );
  OAI211_X1 U19969 ( .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n22294), .A(n18022), 
        .B(n22299), .ZN(P1_U3162) );
  NOR2_X1 U19970 ( .A1(n18024), .A2(n18023), .ZN(P1_U3032) );
  AND2_X1 U19971 ( .A1(n20620), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  AOI21_X1 U19972 ( .B1(n18026), .B2(n18025), .A(n22805), .ZN(P1_U2802) );
  INV_X1 U19973 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18028) );
  OAI22_X1 U19974 ( .A1(n19074), .A2(n18028), .B1(n19436), .B2(n18027), .ZN(
        P2_U2816) );
  AOI22_X1 U19975 ( .A1(n18029), .A2(n18095), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18102), .ZN(n18038) );
  NAND2_X1 U19976 ( .A1(n18030), .A2(n18079), .ZN(n18036) );
  INV_X1 U19977 ( .A(n18031), .ZN(n18032) );
  AOI22_X1 U19978 ( .A1(n18070), .A2(n18032), .B1(n19407), .B2(
        P2_REIP_REG_2__SCAN_IN), .ZN(n18035) );
  NAND2_X1 U19979 ( .A1(n18033), .A2(n18091), .ZN(n18034) );
  AND3_X1 U19980 ( .A1(n18036), .A2(n18035), .A3(n18034), .ZN(n18037) );
  NAND2_X1 U19981 ( .A1(n18038), .A2(n18037), .ZN(P2_U3012) );
  OAI22_X1 U19982 ( .A1(n11748), .A2(n19258), .B1(n18112), .B2(n18039), .ZN(
        n18040) );
  AOI21_X1 U19983 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18102), .A(
        n18040), .ZN(n18044) );
  AOI22_X1 U19984 ( .A1(n18042), .A2(n18095), .B1(n18079), .B2(n18041), .ZN(
        n18043) );
  OAI211_X1 U19985 ( .C1(n18105), .C2(n18045), .A(n18044), .B(n18043), .ZN(
        P2_U3010) );
  AOI22_X1 U19986 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n18102), .B1(
        n18070), .B2(n19121), .ZN(n18052) );
  OAI22_X1 U19987 ( .A1(n18046), .A2(n18103), .B1(n18105), .B2(n19122), .ZN(
        n18047) );
  INV_X1 U19988 ( .A(n18047), .ZN(n18051) );
  OR2_X1 U19989 ( .A1(n18048), .A2(n18106), .ZN(n18050) );
  NAND4_X1 U19990 ( .A1(n18052), .A2(n18051), .A3(n18050), .A4(n18049), .ZN(
        P2_U3009) );
  OAI22_X1 U19991 ( .A1(n11754), .A2(n19258), .B1(n18112), .B2(n19129), .ZN(
        n18053) );
  AOI21_X1 U19992 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18102), .A(
        n18053), .ZN(n18058) );
  OAI22_X1 U19993 ( .A1(n18055), .A2(n18103), .B1(n18106), .B2(n18054), .ZN(
        n18056) );
  INV_X1 U19994 ( .A(n18056), .ZN(n18057) );
  OAI211_X1 U19995 ( .C1(n18105), .C2(n19133), .A(n18058), .B(n18057), .ZN(
        P2_U3008) );
  AOI22_X1 U19996 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18102), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19407), .ZN(n18068) );
  OAI21_X1 U19997 ( .B1(n18061), .B2(n18060), .A(n18059), .ZN(n18062) );
  INV_X1 U19998 ( .A(n18062), .ZN(n19400) );
  NAND2_X1 U19999 ( .A1(n17871), .A2(n18063), .ZN(n18066) );
  XNOR2_X1 U20000 ( .A(n18064), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18065) );
  XNOR2_X1 U20001 ( .A(n18066), .B(n18065), .ZN(n19399) );
  AOI222_X1 U20002 ( .A1(n19400), .A2(n18095), .B1(n18079), .B2(n19399), .C1(
        n18091), .C2(n19397), .ZN(n18067) );
  OAI211_X1 U20003 ( .C1(n18112), .C2(n18069), .A(n18068), .B(n18067), .ZN(
        P2_U3006) );
  AOI22_X1 U20004 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19407), .B1(n18070), 
        .B2(n19156), .ZN(n18075) );
  OAI22_X1 U20005 ( .A1(n18072), .A2(n18103), .B1(n18106), .B2(n18071), .ZN(
        n18073) );
  AOI21_X1 U20006 ( .B1(n18091), .B2(n19157), .A(n18073), .ZN(n18074) );
  OAI211_X1 U20007 ( .C1(n18077), .C2(n18076), .A(n18075), .B(n18074), .ZN(
        P2_U3005) );
  AOI22_X1 U20008 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18102), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19407), .ZN(n18082) );
  AOI222_X1 U20009 ( .A1(n18080), .A2(n18079), .B1(n18091), .B2(n19168), .C1(
        n18095), .C2(n18078), .ZN(n18081) );
  OAI211_X1 U20010 ( .C1(n18112), .C2(n19166), .A(n18082), .B(n18081), .ZN(
        P2_U3004) );
  AOI22_X1 U20011 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18102), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19407), .ZN(n18100) );
  AND2_X1 U20012 ( .A1(n18084), .A2(n18083), .ZN(n18086) );
  NOR2_X1 U20013 ( .A1(n18086), .A2(n18085), .ZN(n18090) );
  NAND2_X1 U20014 ( .A1(n18088), .A2(n18087), .ZN(n18089) );
  XNOR2_X1 U20015 ( .A(n18090), .B(n18089), .ZN(n19389) );
  NAND2_X1 U20016 ( .A1(n19385), .A2(n18091), .ZN(n18097) );
  NAND2_X1 U20017 ( .A1(n18092), .A2(n19393), .ZN(n18093) );
  NAND2_X1 U20018 ( .A1(n19384), .A2(n18095), .ZN(n18096) );
  OAI211_X1 U20019 ( .C1(n19389), .C2(n18106), .A(n18097), .B(n18096), .ZN(
        n18098) );
  INV_X1 U20020 ( .A(n18098), .ZN(n18099) );
  OAI211_X1 U20021 ( .C1(n18112), .C2(n18101), .A(n18100), .B(n18099), .ZN(
        P2_U3002) );
  AOI22_X1 U20022 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18102), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19407), .ZN(n18111) );
  NOR2_X1 U20023 ( .A1(n18104), .A2(n18103), .ZN(n18109) );
  OAI22_X1 U20024 ( .A1(n18107), .A2(n18106), .B1(n18105), .B2(n19206), .ZN(
        n18108) );
  NOR2_X1 U20025 ( .A1(n18109), .A2(n18108), .ZN(n18110) );
  OAI211_X1 U20026 ( .C1(n18112), .C2(n19201), .A(n18111), .B(n18110), .ZN(
        P2_U3000) );
  INV_X1 U20027 ( .A(n18133), .ZN(n18135) );
  INV_X1 U20028 ( .A(n19077), .ZN(n18117) );
  INV_X1 U20029 ( .A(n18113), .ZN(n18115) );
  NOR2_X1 U20030 ( .A1(n18115), .A2(n18114), .ZN(n19442) );
  NOR2_X1 U20031 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20083), .ZN(
        n18116) );
  AOI211_X1 U20032 ( .C1(n20081), .C2(n18117), .A(n19442), .B(n18116), .ZN(
        n18118) );
  AOI22_X1 U20033 ( .A1(n18135), .A2(n20094), .B1(n18118), .B2(n18133), .ZN(
        P2_U3605) );
  NAND2_X1 U20034 ( .A1(n19944), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20008) );
  OR2_X1 U20035 ( .A1(n18127), .A2(n20008), .ZN(n20057) );
  NAND2_X1 U20036 ( .A1(n20008), .A2(n20100), .ZN(n18119) );
  NAND2_X1 U20037 ( .A1(n18119), .A2(n19425), .ZN(n18132) );
  AOI22_X1 U20038 ( .A1(n18127), .A2(n18132), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n18120), .ZN(n18121) );
  OAI21_X1 U20039 ( .B1(n20057), .B2(n20096), .A(n18121), .ZN(n18122) );
  INV_X1 U20040 ( .A(n18122), .ZN(n18123) );
  AOI22_X1 U20041 ( .A1(n18135), .A2(n19998), .B1(n18123), .B2(n18133), .ZN(
        P2_U3603) );
  NAND2_X1 U20042 ( .A1(n20100), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20082) );
  NAND2_X1 U20043 ( .A1(n18128), .A2(n20082), .ZN(n18124) );
  AOI22_X1 U20044 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n18125), .B1(n18132), 
        .B2(n18124), .ZN(n18126) );
  AOI22_X1 U20045 ( .A1(n18135), .A2(n20092), .B1(n18126), .B2(n18133), .ZN(
        P2_U3604) );
  INV_X1 U20046 ( .A(n20058), .ZN(n18131) );
  INV_X1 U20047 ( .A(n19982), .ZN(n19984) );
  OAI21_X1 U20048 ( .B1(n20030), .B2(n18128), .A(n19984), .ZN(n18130) );
  INV_X1 U20049 ( .A(n20082), .ZN(n18129) );
  AOI222_X1 U20050 ( .A1(n18132), .A2(n18131), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19409), .C1(n18130), .C2(n18129), .ZN(n18134) );
  AOI22_X1 U20051 ( .A1(n18135), .A2(n19952), .B1(n18134), .B2(n18133), .ZN(
        P2_U3602) );
  INV_X1 U20052 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22312) );
  NAND2_X1 U20053 ( .A1(n18136), .A2(n22312), .ZN(n18139) );
  OAI21_X1 U20054 ( .B1(n11689), .B2(n16338), .A(n18143), .ZN(n18137) );
  OAI21_X1 U20055 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18143), .A(n18137), 
        .ZN(n18138) );
  OAI221_X1 U20056 ( .B1(n18139), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18139), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18138), .ZN(P2_U2822) );
  INV_X1 U20057 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18142) );
  OAI221_X1 U20058 ( .B1(n18143), .B2(n18142), .C1(n18141), .C2(n18140), .A(
        n18139), .ZN(P2_U2823) );
  OAI22_X1 U20059 ( .A1(n22341), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n18205), .ZN(n18144) );
  INV_X1 U20060 ( .A(n18144), .ZN(P2_U3611) );
  INV_X1 U20061 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n18145) );
  AOI22_X1 U20062 ( .A1(n18205), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n18145), 
        .B2(n22341), .ZN(P2_U3608) );
  AOI21_X1 U20063 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n22313), .ZN(n18146) );
  INV_X1 U20064 ( .A(n18146), .ZN(P2_U2815) );
  AOI22_X1 U20065 ( .A1(n18180), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n18148) );
  OAI21_X1 U20066 ( .B1(n14417), .B2(n18182), .A(n18148), .ZN(P2_U2951) );
  INV_X1 U20067 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n18150) );
  AOI22_X1 U20068 ( .A1(n18180), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n18149) );
  OAI21_X1 U20069 ( .B1(n18150), .B2(n18182), .A(n18149), .ZN(P2_U2950) );
  INV_X1 U20070 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n18152) );
  AOI22_X1 U20071 ( .A1(n18180), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n18159), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n18151) );
  OAI21_X1 U20072 ( .B1(n18152), .B2(n18182), .A(n18151), .ZN(P2_U2949) );
  INV_X1 U20073 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n18154) );
  AOI22_X1 U20074 ( .A1(n18168), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n18159), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n18153) );
  OAI21_X1 U20075 ( .B1(n18154), .B2(n18182), .A(n18153), .ZN(P2_U2948) );
  AOI22_X1 U20076 ( .A1(n18180), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n18159), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n18155) );
  OAI21_X1 U20077 ( .B1(n18156), .B2(n18182), .A(n18155), .ZN(P2_U2947) );
  INV_X1 U20078 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n18158) );
  AOI22_X1 U20079 ( .A1(n18168), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n18159), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n18157) );
  OAI21_X1 U20080 ( .B1(n18158), .B2(n18182), .A(n18157), .ZN(P2_U2946) );
  AOI22_X1 U20081 ( .A1(n18168), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n18159), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n18160) );
  OAI21_X1 U20082 ( .B1(n18161), .B2(n18182), .A(n18160), .ZN(P2_U2945) );
  AOI22_X1 U20083 ( .A1(n18168), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n18162) );
  OAI21_X1 U20084 ( .B1(n18163), .B2(n18182), .A(n18162), .ZN(P2_U2944) );
  AOI22_X1 U20085 ( .A1(n18168), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n18164) );
  OAI21_X1 U20086 ( .B1(n18165), .B2(n18182), .A(n18164), .ZN(P2_U2943) );
  AOI22_X1 U20087 ( .A1(n18180), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n18166) );
  OAI21_X1 U20088 ( .B1(n18167), .B2(n18182), .A(n18166), .ZN(P2_U2942) );
  AOI22_X1 U20089 ( .A1(n18168), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n18169) );
  OAI21_X1 U20090 ( .B1(n18170), .B2(n18182), .A(n18169), .ZN(P2_U2941) );
  AOI22_X1 U20091 ( .A1(n18180), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n18171) );
  OAI21_X1 U20092 ( .B1(n18172), .B2(n18182), .A(n18171), .ZN(P2_U2940) );
  AOI22_X1 U20093 ( .A1(n18180), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n18173) );
  OAI21_X1 U20094 ( .B1(n18174), .B2(n18182), .A(n18173), .ZN(P2_U2939) );
  AOI22_X1 U20095 ( .A1(n18180), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n18175) );
  OAI21_X1 U20096 ( .B1(n18176), .B2(n18182), .A(n18175), .ZN(P2_U2938) );
  AOI22_X1 U20097 ( .A1(n18180), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n18177) );
  OAI21_X1 U20098 ( .B1(n18178), .B2(n18182), .A(n18177), .ZN(P2_U2937) );
  AOI22_X1 U20099 ( .A1(n18180), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n18179), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n18181) );
  OAI21_X1 U20100 ( .B1(n18183), .B2(n18182), .A(n18181), .ZN(P2_U2936) );
  AOI21_X1 U20101 ( .B1(n18185), .B2(n18184), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18186) );
  AOI21_X1 U20102 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n18205), .A(n18186), 
        .ZN(P2_U2817) );
  NOR2_X1 U20103 ( .A1(n22354), .A2(n22341), .ZN(n22343) );
  OAI222_X1 U20104 ( .A1(n18207), .A2(n14569), .B1(n20551), .B2(n18205), .C1(
        n11689), .C2(n22352), .ZN(P2_U3212) );
  INV_X1 U20105 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n18187) );
  OAI222_X1 U20106 ( .A1(n18202), .A2(n11736), .B1(n18187), .B2(n18205), .C1(
        n14569), .C2(n22352), .ZN(P2_U3213) );
  INV_X1 U20107 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n18188) );
  OAI222_X1 U20108 ( .A1(n18202), .A2(n11748), .B1(n18188), .B2(n18205), .C1(
        n11736), .C2(n22352), .ZN(P2_U3214) );
  INV_X1 U20109 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n18189) );
  OAI222_X1 U20110 ( .A1(n18202), .A2(n16079), .B1(n18189), .B2(n18205), .C1(
        n11748), .C2(n22352), .ZN(P2_U3215) );
  INV_X1 U20111 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n18190) );
  OAI222_X1 U20112 ( .A1(n18202), .A2(n11754), .B1(n18190), .B2(n18205), .C1(
        n16079), .C2(n22352), .ZN(P2_U3216) );
  INV_X1 U20113 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20557) );
  OAI222_X1 U20114 ( .A1(n18202), .A2(n11757), .B1(n20557), .B2(n18205), .C1(
        n11754), .C2(n22352), .ZN(P2_U3217) );
  INV_X1 U20115 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20559) );
  OAI222_X1 U20116 ( .A1(n18207), .A2(n11761), .B1(n20559), .B2(n18205), .C1(
        n11757), .C2(n22352), .ZN(P2_U3218) );
  INV_X1 U20117 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20561) );
  OAI222_X1 U20118 ( .A1(n18207), .A2(n11763), .B1(n20561), .B2(n18205), .C1(
        n11761), .C2(n22352), .ZN(P2_U3219) );
  INV_X1 U20119 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20563) );
  OAI222_X1 U20120 ( .A1(n22352), .A2(n11763), .B1(n20563), .B2(n18205), .C1(
        n11767), .C2(n18202), .ZN(P2_U3220) );
  INV_X1 U20121 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20565) );
  OAI222_X1 U20122 ( .A1(n22352), .A2(n11767), .B1(n20565), .B2(n18205), .C1(
        n17624), .C2(n18202), .ZN(P2_U3221) );
  INV_X1 U20123 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20567) );
  OAI222_X1 U20124 ( .A1(n22352), .A2(n17624), .B1(n20567), .B2(n18205), .C1(
        n11776), .C2(n18202), .ZN(P2_U3222) );
  INV_X1 U20125 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20569) );
  OAI222_X1 U20126 ( .A1(n22352), .A2(n11776), .B1(n20569), .B2(n18205), .C1(
        n19187), .C2(n18202), .ZN(P2_U3223) );
  INV_X1 U20127 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20571) );
  OAI222_X1 U20128 ( .A1(n22352), .A2(n19187), .B1(n20571), .B2(n18205), .C1(
        n11783), .C2(n18202), .ZN(P2_U3224) );
  INV_X1 U20129 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n18191) );
  OAI222_X1 U20130 ( .A1(n22352), .A2(n11783), .B1(n18191), .B2(n18205), .C1(
        n18193), .C2(n18202), .ZN(P2_U3225) );
  INV_X1 U20131 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n18192) );
  OAI222_X1 U20132 ( .A1(n22352), .A2(n18193), .B1(n18192), .B2(n18205), .C1(
        n11789), .C2(n18202), .ZN(P2_U3226) );
  INV_X1 U20133 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20575) );
  OAI222_X1 U20134 ( .A1(n22352), .A2(n11789), .B1(n20575), .B2(n18205), .C1(
        n17585), .C2(n18202), .ZN(P2_U3227) );
  INV_X1 U20135 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20577) );
  OAI222_X1 U20136 ( .A1(n22352), .A2(n17585), .B1(n20577), .B2(n18205), .C1(
        n17571), .C2(n18202), .ZN(P2_U3228) );
  INV_X1 U20137 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20579) );
  OAI222_X1 U20138 ( .A1(n18207), .A2(n19260), .B1(n20579), .B2(n18205), .C1(
        n17571), .C2(n22352), .ZN(P2_U3229) );
  INV_X1 U20139 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20581) );
  OAI222_X1 U20140 ( .A1(n22352), .A2(n19260), .B1(n20581), .B2(n18205), .C1(
        n17551), .C2(n18202), .ZN(P2_U3230) );
  INV_X1 U20141 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20583) );
  OAI222_X1 U20142 ( .A1(n18207), .A2(n11805), .B1(n20583), .B2(n18205), .C1(
        n17551), .C2(n22352), .ZN(P2_U3231) );
  INV_X1 U20143 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n18194) );
  OAI222_X1 U20144 ( .A1(n18207), .A2(n18195), .B1(n18194), .B2(n18205), .C1(
        n11805), .C2(n22352), .ZN(P2_U3232) );
  INV_X1 U20145 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n18196) );
  OAI222_X1 U20146 ( .A1(n18207), .A2(n18197), .B1(n18196), .B2(n18205), .C1(
        n18195), .C2(n22352), .ZN(P2_U3233) );
  INV_X1 U20147 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20587) );
  OAI222_X1 U20148 ( .A1(n18207), .A2(n18198), .B1(n20587), .B2(n18205), .C1(
        n18197), .C2(n22352), .ZN(P2_U3234) );
  INV_X1 U20149 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20589) );
  OAI222_X1 U20150 ( .A1(n18207), .A2(n18199), .B1(n20589), .B2(n18205), .C1(
        n18198), .C2(n22352), .ZN(P2_U3235) );
  INV_X1 U20151 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20591) );
  OAI222_X1 U20152 ( .A1(n22352), .A2(n18199), .B1(n20591), .B2(n18205), .C1(
        n18200), .C2(n18202), .ZN(P2_U3236) );
  INV_X1 U20153 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20593) );
  OAI222_X1 U20154 ( .A1(n18207), .A2(n18201), .B1(n20593), .B2(n18205), .C1(
        n18200), .C2(n22352), .ZN(P2_U3237) );
  INV_X1 U20155 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20595) );
  OAI222_X1 U20156 ( .A1(n22352), .A2(n18201), .B1(n20595), .B2(n18205), .C1(
        n14043), .C2(n18202), .ZN(P2_U3238) );
  INV_X1 U20157 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20597) );
  OAI222_X1 U20158 ( .A1(n22352), .A2(n14043), .B1(n20597), .B2(n18205), .C1(
        n19326), .C2(n18202), .ZN(P2_U3239) );
  INV_X1 U20159 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n18203) );
  OAI222_X1 U20160 ( .A1(n22352), .A2(n19326), .B1(n18203), .B2(n18205), .C1(
        n18204), .C2(n18202), .ZN(P2_U3240) );
  INV_X1 U20161 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n18206) );
  OAI222_X1 U20162 ( .A1(n18207), .A2(n19339), .B1(n18206), .B2(n18205), .C1(
        n18204), .C2(n22352), .ZN(P2_U3241) );
  OAI22_X1 U20163 ( .A1(n22341), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n18205), .ZN(n18208) );
  INV_X1 U20164 ( .A(n18208), .ZN(P2_U3588) );
  OAI22_X1 U20165 ( .A1(n22341), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n18205), .ZN(n18209) );
  INV_X1 U20166 ( .A(n18209), .ZN(P2_U3587) );
  MUX2_X1 U20167 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n22341), .Z(P2_U3586) );
  OAI22_X1 U20168 ( .A1(n22341), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n18205), .ZN(n18210) );
  INV_X1 U20169 ( .A(n18210), .ZN(P2_U3585) );
  NOR2_X1 U20170 ( .A1(n21443), .A2(n18564), .ZN(n18560) );
  AND2_X1 U20171 ( .A1(n18211), .A2(n18560), .ZN(n18217) );
  AND2_X1 U20172 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n18217), .ZN(n18215) );
  AOI21_X1 U20173 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n18562), .A(n18215), .ZN(
        n18212) );
  OAI22_X1 U20174 ( .A1(n18237), .A2(n18212), .B1(n11271), .B2(n18562), .ZN(
        P3_U2699) );
  AOI21_X1 U20175 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n18562), .A(n18217), .ZN(
        n18214) );
  OAI22_X1 U20176 ( .A1(n18215), .A2(n18214), .B1(n18213), .B2(n18562), .ZN(
        P3_U2700) );
  INV_X1 U20177 ( .A(n18216), .ZN(n18559) );
  INV_X1 U20178 ( .A(n18564), .ZN(n18324) );
  AOI221_X1 U20179 ( .B1(n18559), .B2(n18324), .C1(n21443), .C2(n18324), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n18218) );
  AOI211_X1 U20180 ( .C1(n18565), .C2(n11287), .A(n18218), .B(n18217), .ZN(
        P3_U2701) );
  AOI22_X1 U20181 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18222) );
  AOI22_X1 U20182 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18221) );
  AOI22_X1 U20183 ( .A1(n18523), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18220) );
  NAND4_X1 U20184 ( .A1(n18222), .A2(n18221), .A3(n18220), .A4(n18219), .ZN(
        n18228) );
  AOI22_X1 U20185 ( .A1(n18393), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18480), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18226) );
  AOI22_X1 U20186 ( .A1(n18540), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11157), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18225) );
  AOI22_X1 U20187 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18498), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18224) );
  AOI22_X1 U20188 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11156), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18223) );
  NAND4_X1 U20189 ( .A1(n18226), .A2(n18225), .A3(n18224), .A4(n18223), .ZN(
        n18227) );
  NOR2_X1 U20190 ( .A1(n18228), .A2(n18227), .ZN(n21515) );
  INV_X1 U20191 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n21012) );
  OAI33_X1 U20192 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n21443), .A3(n18316), .B1(
        n21012), .B2(n18565), .B3(n18229), .ZN(n18230) );
  INV_X1 U20193 ( .A(n18230), .ZN(n18231) );
  OAI21_X1 U20194 ( .B1(n21515), .B2(n18562), .A(n18231), .ZN(P3_U2695) );
  INV_X1 U20195 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18380) );
  INV_X1 U20196 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n20977) );
  NAND3_X1 U20197 ( .A1(n21524), .A2(P3_EBX_REG_5__SCAN_IN), .A3(n18237), .ZN(
        n18236) );
  NOR2_X1 U20198 ( .A1(n20977), .A2(n18236), .ZN(n18235) );
  OAI211_X1 U20199 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n18235), .A(n18316), .B(
        n18562), .ZN(n18232) );
  OAI21_X1 U20200 ( .B1(n18562), .B2(n18380), .A(n18232), .ZN(P3_U2696) );
  INV_X1 U20201 ( .A(n18236), .ZN(n18233) );
  AOI21_X1 U20202 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n18562), .A(n18233), .ZN(
        n18234) );
  OAI22_X1 U20203 ( .A1(n18235), .A2(n18234), .B1(n11261), .B2(n18562), .ZN(
        P3_U2697) );
  OAI21_X1 U20204 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n18237), .A(n18236), .ZN(
        n18238) );
  AOI22_X1 U20205 ( .A1(n18565), .A2(n11267), .B1(n18238), .B2(n18562), .ZN(
        P3_U2698) );
  NAND2_X1 U20206 ( .A1(n21524), .A2(n18239), .ZN(n18251) );
  AOI22_X1 U20207 ( .A1(n18547), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18243) );
  AOI22_X1 U20208 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18381), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18242) );
  AOI22_X1 U20209 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n20948), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18241) );
  AOI22_X1 U20210 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18240) );
  NAND4_X1 U20211 ( .A1(n18243), .A2(n18242), .A3(n18241), .A4(n18240), .ZN(
        n18249) );
  AOI22_X1 U20212 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18247) );
  AOI22_X1 U20213 ( .A1(n18393), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11157), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18246) );
  AOI22_X1 U20214 ( .A1(n18480), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18245) );
  NAND4_X1 U20215 ( .A1(n18247), .A2(n18246), .A3(n18245), .A4(n18244), .ZN(
        n18248) );
  NOR2_X1 U20216 ( .A1(n18249), .A2(n18248), .ZN(n21496) );
  NAND3_X1 U20217 ( .A1(n18251), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n18562), 
        .ZN(n18250) );
  OAI221_X1 U20218 ( .B1(n18251), .B2(P3_EBX_REG_16__SCAN_IN), .C1(n18562), 
        .C2(n21496), .A(n18250), .ZN(P3_U2687) );
  AOI22_X1 U20219 ( .A1(n18547), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n18263) );
  AOI22_X1 U20220 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11157), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18262) );
  INV_X1 U20221 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18253) );
  AOI22_X1 U20222 ( .A1(n18523), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n18252) );
  OAI21_X1 U20223 ( .B1(n18254), .B2(n18253), .A(n18252), .ZN(n18260) );
  AOI22_X1 U20224 ( .A1(n18540), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18480), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18258) );
  AOI22_X1 U20225 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18257) );
  AOI22_X1 U20226 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13798), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18256) );
  AOI22_X1 U20227 ( .A1(n18279), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18255) );
  NAND4_X1 U20228 ( .A1(n18258), .A2(n18257), .A3(n18256), .A4(n18255), .ZN(
        n18259) );
  AOI211_X1 U20229 ( .C1(n18393), .C2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n18260), .B(n18259), .ZN(n18261) );
  NAND3_X1 U20230 ( .A1(n18263), .A2(n18262), .A3(n18261), .ZN(n21346) );
  INV_X1 U20231 ( .A(n21346), .ZN(n18265) );
  AOI21_X1 U20232 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n18290), .A(
        P3_EBX_REG_13__SCAN_IN), .ZN(n18264) );
  NAND4_X1 U20233 ( .A1(n21524), .A2(P3_EBX_REG_13__SCAN_IN), .A3(
        P3_EBX_REG_12__SCAN_IN), .A4(n18290), .ZN(n18278) );
  NAND2_X1 U20234 ( .A1(n18562), .A2(n18278), .ZN(n18277) );
  OAI22_X1 U20235 ( .A1(n18265), .A2(n18562), .B1(n18264), .B2(n18277), .ZN(
        P3_U2690) );
  INV_X1 U20236 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n21087) );
  AOI22_X1 U20237 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18275) );
  AOI22_X1 U20238 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18498), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18274) );
  AOI22_X1 U20239 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18381), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18266) );
  OAI21_X1 U20240 ( .B1(n11206), .B2(n11261), .A(n18266), .ZN(n18272) );
  AOI22_X1 U20241 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18270) );
  AOI22_X1 U20242 ( .A1(n13798), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18269) );
  AOI22_X1 U20243 ( .A1(n18279), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18267) );
  NAND4_X1 U20244 ( .A1(n18270), .A2(n18269), .A3(n18268), .A4(n18267), .ZN(
        n18271) );
  AOI211_X1 U20245 ( .C1(n18388), .C2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n18272), .B(n18271), .ZN(n18273) );
  NAND3_X1 U20246 ( .A1(n18275), .A2(n18274), .A3(n18273), .ZN(n21498) );
  NAND2_X1 U20247 ( .A1(n18565), .A2(n21498), .ZN(n18276) );
  OAI221_X1 U20248 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n18278), .C1(n21087), 
        .C2(n18277), .A(n18276), .ZN(P3_U2689) );
  AOI22_X1 U20249 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18545), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18283) );
  AOI22_X1 U20250 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18281) );
  AOI22_X1 U20251 ( .A1(n18279), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18280) );
  NAND4_X1 U20252 ( .A1(n18283), .A2(n18282), .A3(n18281), .A4(n18280), .ZN(
        n18289) );
  AOI22_X1 U20253 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18287) );
  AOI22_X1 U20254 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18498), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18286) );
  AOI22_X1 U20255 ( .A1(n18480), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18285) );
  AOI22_X1 U20256 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18381), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18284) );
  NAND4_X1 U20257 ( .A1(n18287), .A2(n18286), .A3(n18285), .A4(n18284), .ZN(
        n18288) );
  NOR2_X1 U20258 ( .A1(n18289), .A2(n18288), .ZN(n21353) );
  INV_X1 U20259 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n21058) );
  AOI22_X1 U20260 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n18291), .B1(n18290), 
        .B2(n21058), .ZN(n18292) );
  AOI22_X1 U20261 ( .A1(n18565), .A2(n21353), .B1(n18292), .B2(n18562), .ZN(
        P3_U2691) );
  NOR2_X1 U20262 ( .A1(n18565), .A2(n18293), .ZN(n18317) );
  AOI22_X1 U20263 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18303) );
  AOI22_X1 U20264 ( .A1(n18547), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11157), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18302) );
  AOI22_X1 U20265 ( .A1(n20948), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18294) );
  OAI21_X1 U20266 ( .B1(n11206), .B2(n11287), .A(n18294), .ZN(n18300) );
  AOI22_X1 U20267 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18297) );
  AOI22_X1 U20268 ( .A1(n18480), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18296) );
  AOI22_X1 U20269 ( .A1(n13798), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18381), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18295) );
  NAND4_X1 U20270 ( .A1(n18298), .A2(n18297), .A3(n18296), .A4(n18295), .ZN(
        n18299) );
  AOI211_X1 U20271 ( .C1(n18388), .C2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A(
        n18300), .B(n18299), .ZN(n18301) );
  NAND3_X1 U20272 ( .A1(n18303), .A2(n18302), .A3(n18301), .ZN(n21359) );
  AOI22_X1 U20273 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18317), .B1(n18565), 
        .B2(n21359), .ZN(n18304) );
  OAI21_X1 U20274 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n18305), .A(n18304), .ZN(
        P3_U2693) );
  AOI22_X1 U20275 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18547), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n13899), .ZN(n18309) );
  AOI22_X1 U20276 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18545), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18308) );
  AOI22_X1 U20277 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20948), .B1(
        n18381), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18307) );
  AOI22_X1 U20278 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18548), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n11151), .ZN(n18306) );
  NAND4_X1 U20279 ( .A1(n18309), .A2(n18308), .A3(n18307), .A4(n18306), .ZN(
        n18315) );
  AOI22_X1 U20280 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18546), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n11157), .ZN(n18313) );
  AOI22_X1 U20281 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n18539), .ZN(n18312) );
  AOI22_X1 U20282 ( .A1(n18523), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18480), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18311) );
  AOI22_X1 U20283 ( .A1(n13798), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n11156), .ZN(n18310) );
  NAND4_X1 U20284 ( .A1(n18313), .A2(n18312), .A3(n18311), .A4(n18310), .ZN(
        n18314) );
  NOR2_X1 U20285 ( .A1(n18315), .A2(n18314), .ZN(n21364) );
  NOR2_X1 U20286 ( .A1(n21012), .A2(n18316), .ZN(n18318) );
  OAI21_X1 U20287 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n18318), .A(n18317), .ZN(
        n18319) );
  OAI21_X1 U20288 ( .B1(n21364), .B2(n18562), .A(n18319), .ZN(P3_U2694) );
  INV_X1 U20289 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n21172) );
  INV_X1 U20290 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n21145) );
  INV_X1 U20291 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n21129) );
  INV_X1 U20292 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n21108) );
  NOR4_X1 U20293 ( .A1(n21108), .A2(n18322), .A3(n18321), .A4(n18320), .ZN(
        n18323) );
  NAND4_X1 U20294 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .A4(n18323), .ZN(n18556) );
  NOR2_X1 U20295 ( .A1(n21129), .A2(n18556), .ZN(n18555) );
  NAND2_X1 U20296 ( .A1(n18324), .A2(n18555), .ZN(n18508) );
  NOR2_X1 U20297 ( .A1(n21145), .A2(n18508), .ZN(n18536) );
  NAND2_X1 U20298 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n18536), .ZN(n18535) );
  NOR2_X1 U20299 ( .A1(n21172), .A2(n18535), .ZN(n18439) );
  INV_X1 U20300 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n21254) );
  INV_X1 U20301 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n21238) );
  NAND4_X1 U20302 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n18442)
         );
  NAND2_X1 U20303 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n18446) );
  NOR4_X1 U20304 ( .A1(n21254), .A2(n21238), .A3(n18442), .A4(n18446), .ZN(
        n18449) );
  NAND4_X1 U20305 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(P3_EBX_REG_29__SCAN_IN), 
        .A3(n18439), .A4(n18449), .ZN(n18425) );
  INV_X1 U20306 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n18326) );
  INV_X1 U20307 ( .A(n18425), .ZN(n18325) );
  OAI33_X1 U20308 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n21443), .A3(n18425), 
        .B1(n18326), .B2(n18565), .B3(n18325), .ZN(P3_U2672) );
  AOI22_X1 U20309 ( .A1(n18523), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18330) );
  AOI22_X1 U20310 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11157), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18329) );
  AOI22_X1 U20311 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18480), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18328) );
  NAND4_X1 U20312 ( .A1(n18330), .A2(n18329), .A3(n18328), .A4(n18327), .ZN(
        n18337) );
  AOI22_X1 U20313 ( .A1(n18393), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18498), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18335) );
  AOI22_X1 U20314 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11156), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18334) );
  AOI22_X1 U20315 ( .A1(n18540), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18333) );
  AOI22_X1 U20316 ( .A1(n20948), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18332) );
  NAND4_X1 U20317 ( .A1(n18335), .A2(n18334), .A3(n18333), .A4(n18332), .ZN(
        n18336) );
  NOR2_X1 U20318 ( .A1(n18337), .A2(n18336), .ZN(n18424) );
  AOI22_X1 U20319 ( .A1(n18540), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18341) );
  AOI22_X1 U20320 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18340) );
  AOI22_X1 U20321 ( .A1(n18547), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n18339) );
  AOI22_X1 U20322 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n20948), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18338) );
  NAND4_X1 U20323 ( .A1(n18341), .A2(n18340), .A3(n18339), .A4(n18338), .ZN(
        n18347) );
  AOI22_X1 U20324 ( .A1(n18393), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18480), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18345) );
  AOI22_X1 U20325 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11157), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18344) );
  AOI22_X1 U20326 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n18342) );
  NAND4_X1 U20327 ( .A1(n18345), .A2(n18344), .A3(n18343), .A4(n18342), .ZN(
        n18346) );
  NOR2_X1 U20328 ( .A1(n18347), .A2(n18346), .ZN(n18453) );
  AOI22_X1 U20329 ( .A1(n18393), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18480), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18351) );
  AOI22_X1 U20330 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18381), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18350) );
  AOI22_X1 U20331 ( .A1(n18523), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18348) );
  NAND4_X1 U20332 ( .A1(n18351), .A2(n18350), .A3(n18349), .A4(n18348), .ZN(
        n18357) );
  AOI22_X1 U20333 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18498), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18355) );
  AOI22_X1 U20334 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18354) );
  AOI22_X1 U20335 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18353) );
  AOI22_X1 U20336 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11156), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18352) );
  NAND4_X1 U20337 ( .A1(n18355), .A2(n18354), .A3(n18353), .A4(n18352), .ZN(
        n18356) );
  NOR2_X1 U20338 ( .A1(n18357), .A2(n18356), .ZN(n18459) );
  AOI22_X1 U20339 ( .A1(n18547), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18361) );
  AOI22_X1 U20340 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18545), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n18538), .ZN(n18360) );
  AOI22_X1 U20341 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n20948), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18359) );
  AOI22_X1 U20342 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18546), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n11151), .ZN(n18358) );
  NAND4_X1 U20343 ( .A1(n18361), .A2(n18360), .A3(n18359), .A4(n18358), .ZN(
        n18367) );
  AOI22_X1 U20344 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n18514), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n18365) );
  AOI22_X1 U20345 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18364) );
  AOI22_X1 U20346 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n11157), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18363) );
  AOI22_X1 U20347 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18381), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18362) );
  NAND4_X1 U20348 ( .A1(n18365), .A2(n18364), .A3(n18363), .A4(n18362), .ZN(
        n18366) );
  NOR2_X1 U20349 ( .A1(n18367), .A2(n18366), .ZN(n18470) );
  AOI22_X1 U20350 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11156), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18378) );
  AOI22_X1 U20351 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18545), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18377) );
  INV_X1 U20352 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18369) );
  AOI22_X1 U20353 ( .A1(n18497), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18368) );
  OAI21_X1 U20354 ( .B1(n18414), .B2(n18369), .A(n18368), .ZN(n18375) );
  AOI22_X1 U20355 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18480), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18373) );
  AOI22_X1 U20356 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18372) );
  AOI22_X1 U20357 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n18371) );
  NAND4_X1 U20358 ( .A1(n18373), .A2(n18372), .A3(n18371), .A4(n18370), .ZN(
        n18374) );
  AOI211_X1 U20359 ( .C1(n18540), .C2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n18375), .B(n18374), .ZN(n18376) );
  NAND3_X1 U20360 ( .A1(n18378), .A2(n18377), .A3(n18376), .ZN(n18475) );
  AOI22_X1 U20361 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18391) );
  AOI22_X1 U20362 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11156), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18379) );
  OAI21_X1 U20363 ( .B1(n11514), .B2(n18380), .A(n18379), .ZN(n18387) );
  AOI22_X1 U20364 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18385) );
  AOI22_X1 U20365 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18381), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18384) );
  AOI22_X1 U20366 ( .A1(n18393), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18498), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18383) );
  AOI22_X1 U20367 ( .A1(n20948), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18382) );
  NAND4_X1 U20368 ( .A1(n18385), .A2(n18384), .A3(n18383), .A4(n18382), .ZN(
        n18386) );
  AOI211_X1 U20369 ( .C1(n18388), .C2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n18387), .B(n18386), .ZN(n18389) );
  NAND3_X1 U20370 ( .A1(n18391), .A2(n18390), .A3(n18389), .ZN(n18476) );
  NAND2_X1 U20371 ( .A1(n18475), .A2(n18476), .ZN(n18474) );
  NOR2_X1 U20372 ( .A1(n18470), .A2(n18474), .ZN(n18469) );
  AOI22_X1 U20373 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18402) );
  AOI22_X1 U20374 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18540), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18401) );
  AOI22_X1 U20375 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18392) );
  OAI21_X1 U20376 ( .B1(n18414), .B2(n11287), .A(n18392), .ZN(n18399) );
  AOI22_X1 U20377 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18480), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18396) );
  AOI22_X1 U20378 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18395) );
  AOI22_X1 U20379 ( .A1(n20948), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18394) );
  NAND4_X1 U20380 ( .A1(n18397), .A2(n18396), .A3(n18395), .A4(n18394), .ZN(
        n18398) );
  AOI211_X1 U20381 ( .C1(n13798), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n18399), .B(n18398), .ZN(n18400) );
  NAND3_X1 U20382 ( .A1(n18402), .A2(n18401), .A3(n18400), .ZN(n18464) );
  NAND2_X1 U20383 ( .A1(n18469), .A2(n18464), .ZN(n18463) );
  NOR2_X1 U20384 ( .A1(n18459), .A2(n18463), .ZN(n18458) );
  AOI22_X1 U20385 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18412) );
  AOI22_X1 U20386 ( .A1(n18523), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18480), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18411) );
  AOI22_X1 U20387 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18403) );
  OAI21_X1 U20388 ( .B1(n18414), .B2(n11271), .A(n18403), .ZN(n18409) );
  AOI22_X1 U20389 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18514), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n18407) );
  AOI22_X1 U20390 ( .A1(n18393), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11156), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18405) );
  AOI22_X1 U20391 ( .A1(n20948), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18404) );
  NAND4_X1 U20392 ( .A1(n18407), .A2(n18406), .A3(n18405), .A4(n18404), .ZN(
        n18408) );
  AOI211_X1 U20393 ( .C1(n11159), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n18409), .B(n18408), .ZN(n18410) );
  NAND3_X1 U20394 ( .A1(n18412), .A2(n18411), .A3(n18410), .ZN(n18441) );
  NAND2_X1 U20395 ( .A1(n18458), .A2(n18441), .ZN(n18452) );
  NOR2_X1 U20396 ( .A1(n18453), .A2(n18452), .ZN(n18451) );
  AOI22_X1 U20397 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18514), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18423) );
  AOI22_X1 U20398 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18540), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18422) );
  OAI21_X1 U20399 ( .B1(n18414), .B2(n11261), .A(n18413), .ZN(n18420) );
  AOI22_X1 U20400 ( .A1(n18497), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18538), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18418) );
  AOI22_X1 U20401 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18417) );
  AOI22_X1 U20402 ( .A1(n18393), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18416) );
  AOI22_X1 U20403 ( .A1(n20948), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18415) );
  NAND4_X1 U20404 ( .A1(n18418), .A2(n18417), .A3(n18416), .A4(n18415), .ZN(
        n18419) );
  AOI211_X1 U20405 ( .C1(n18388), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n18420), .B(n18419), .ZN(n18421) );
  NAND3_X1 U20406 ( .A1(n18423), .A2(n18422), .A3(n18421), .ZN(n18445) );
  NAND2_X1 U20407 ( .A1(n18451), .A2(n18445), .ZN(n18444) );
  XNOR2_X1 U20408 ( .A(n18424), .B(n18444), .ZN(n21460) );
  AND3_X1 U20409 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n18439), .A3(n18449), .ZN(
        n18426) );
  OAI211_X1 U20410 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n18426), .A(n18425), .B(
        n18562), .ZN(n18427) );
  OAI21_X1 U20411 ( .B1(n21460), .B2(n18562), .A(n18427), .ZN(P3_U2673) );
  AOI22_X1 U20412 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18431) );
  AOI22_X1 U20413 ( .A1(n18480), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18430) );
  AOI22_X1 U20414 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11157), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n18429) );
  AOI22_X1 U20415 ( .A1(n20948), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18428) );
  NAND4_X1 U20416 ( .A1(n18431), .A2(n18430), .A3(n18429), .A4(n18428), .ZN(
        n18438) );
  AOI22_X1 U20417 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18498), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18436) );
  AOI22_X1 U20418 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18540), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18435) );
  AOI22_X1 U20419 ( .A1(n18545), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18433) );
  NAND4_X1 U20420 ( .A1(n18436), .A2(n18435), .A3(n18434), .A4(n18433), .ZN(
        n18437) );
  NOR2_X1 U20421 ( .A1(n18438), .A2(n18437), .ZN(n21407) );
  NOR2_X1 U20422 ( .A1(n18565), .A2(n18439), .ZN(n18505) );
  NAND2_X1 U20423 ( .A1(n21524), .A2(n18439), .ZN(n18467) );
  INV_X1 U20424 ( .A(n18467), .ZN(n18479) );
  INV_X1 U20425 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n18468) );
  AOI22_X1 U20426 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n18505), .B1(n18479), 
        .B2(n18468), .ZN(n18440) );
  OAI21_X1 U20427 ( .B1(n21407), .B2(n18562), .A(n18440), .ZN(P3_U2682) );
  OAI21_X1 U20428 ( .B1(n18458), .B2(n18441), .A(n18452), .ZN(n21478) );
  NOR2_X1 U20429 ( .A1(n18467), .A2(n18442), .ZN(n18473) );
  NAND2_X1 U20430 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n18473), .ZN(n18457) );
  NOR2_X1 U20431 ( .A1(n21254), .A2(n18457), .ZN(n18462) );
  NAND2_X1 U20432 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n18462), .ZN(n18456) );
  OAI211_X1 U20433 ( .C1(n18462), .C2(P3_EBX_REG_27__SCAN_IN), .A(n18562), .B(
        n18456), .ZN(n18443) );
  OAI21_X1 U20434 ( .B1(n18562), .B2(n21478), .A(n18443), .ZN(P3_U2676) );
  OAI21_X1 U20435 ( .B1(n18451), .B2(n18445), .A(n18444), .ZN(n21467) );
  INV_X1 U20436 ( .A(n18446), .ZN(n18447) );
  INV_X1 U20437 ( .A(n18560), .ZN(n18567) );
  OAI22_X1 U20438 ( .A1(n18565), .A2(n18462), .B1(n18447), .B2(n18567), .ZN(
        n18454) );
  NOR2_X1 U20439 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n18467), .ZN(n18448) );
  AOI22_X1 U20440 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n18454), .B1(n18449), 
        .B2(n18448), .ZN(n18450) );
  OAI21_X1 U20441 ( .B1(n21467), .B2(n18562), .A(n18450), .ZN(P3_U2674) );
  AOI21_X1 U20442 ( .B1(n18453), .B2(n18452), .A(n18451), .ZN(n21468) );
  AOI22_X1 U20443 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18454), .B1(n21468), 
        .B2(n18565), .ZN(n18455) );
  OAI21_X1 U20444 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n18456), .A(n18455), .ZN(
        P3_U2675) );
  INV_X1 U20445 ( .A(n18457), .ZN(n18466) );
  AOI21_X1 U20446 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n18562), .A(n18466), .ZN(
        n18461) );
  AOI21_X1 U20447 ( .B1(n18459), .B2(n18463), .A(n18458), .ZN(n21448) );
  INV_X1 U20448 ( .A(n21448), .ZN(n18460) );
  OAI22_X1 U20449 ( .A1(n18462), .A2(n18461), .B1(n18460), .B2(n18562), .ZN(
        P3_U2677) );
  AOI21_X1 U20450 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18562), .A(n18473), .ZN(
        n18465) );
  OAI21_X1 U20451 ( .B1(n18469), .B2(n18464), .A(n18463), .ZN(n21447) );
  OAI22_X1 U20452 ( .A1(n18466), .A2(n18465), .B1(n21447), .B2(n18562), .ZN(
        P3_U2678) );
  INV_X1 U20453 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n21198) );
  NOR3_X1 U20454 ( .A1(n21198), .A2(n18468), .A3(n18467), .ZN(n18492) );
  AND2_X1 U20455 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n18492), .ZN(n18478) );
  AOI21_X1 U20456 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18562), .A(n18478), .ZN(
        n18472) );
  AOI21_X1 U20457 ( .B1(n18470), .B2(n18474), .A(n18469), .ZN(n21479) );
  INV_X1 U20458 ( .A(n21479), .ZN(n18471) );
  OAI22_X1 U20459 ( .A1(n18473), .A2(n18472), .B1(n18471), .B2(n18562), .ZN(
        P3_U2679) );
  AOI21_X1 U20460 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18562), .A(n18492), .ZN(
        n18477) );
  OAI21_X1 U20461 ( .B1(n18476), .B2(n18475), .A(n18474), .ZN(n21490) );
  OAI22_X1 U20462 ( .A1(n18478), .A2(n18477), .B1(n21490), .B2(n18562), .ZN(
        P3_U2680) );
  AOI22_X1 U20463 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n18562), .B1(
        P3_EBX_REG_21__SCAN_IN), .B2(n18479), .ZN(n18491) );
  AOI22_X1 U20464 ( .A1(n18393), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18484) );
  AOI22_X1 U20465 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11157), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18483) );
  AOI22_X1 U20466 ( .A1(n20948), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18481) );
  NAND4_X1 U20467 ( .A1(n18484), .A2(n18483), .A3(n18482), .A4(n18481), .ZN(
        n18490) );
  AOI22_X1 U20468 ( .A1(n18547), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18488) );
  AOI22_X1 U20469 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18540), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18487) );
  AOI22_X1 U20470 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18486) );
  AOI22_X1 U20471 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11159), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18485) );
  NAND4_X1 U20472 ( .A1(n18488), .A2(n18487), .A3(n18486), .A4(n18485), .ZN(
        n18489) );
  NOR2_X1 U20473 ( .A1(n18490), .A2(n18489), .ZN(n21419) );
  OAI22_X1 U20474 ( .A1(n18492), .A2(n18491), .B1(n21419), .B2(n18562), .ZN(
        P3_U2681) );
  AOI22_X1 U20475 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18496) );
  AOI22_X1 U20476 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18540), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18495) );
  AOI22_X1 U20477 ( .A1(n18545), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18494) );
  NAND4_X1 U20478 ( .A1(n18496), .A2(n18495), .A3(n18494), .A4(n18493), .ZN(
        n18504) );
  AOI22_X1 U20479 ( .A1(n13916), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n18502) );
  AOI22_X1 U20480 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18498), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18501) );
  AOI22_X1 U20481 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18500) );
  AOI22_X1 U20482 ( .A1(n11157), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18538), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18499) );
  NAND4_X1 U20483 ( .A1(n18502), .A2(n18501), .A3(n18500), .A4(n18499), .ZN(
        n18503) );
  NOR2_X1 U20484 ( .A1(n18504), .A2(n18503), .ZN(n21414) );
  INV_X1 U20485 ( .A(n18535), .ZN(n18506) );
  OAI21_X1 U20486 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n18506), .A(n18505), .ZN(
        n18507) );
  OAI21_X1 U20487 ( .B1(n21414), .B2(n18562), .A(n18507), .ZN(P3_U2683) );
  AOI21_X1 U20488 ( .B1(n21145), .B2(n18508), .A(n18565), .ZN(n18509) );
  INV_X1 U20489 ( .A(n18509), .ZN(n18521) );
  AOI22_X1 U20490 ( .A1(n18545), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18513) );
  AOI22_X1 U20491 ( .A1(n18547), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18497), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18512) );
  AOI22_X1 U20492 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n20948), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18511) );
  AOI22_X1 U20493 ( .A1(n18540), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18510) );
  NAND4_X1 U20494 ( .A1(n18513), .A2(n18512), .A3(n18511), .A4(n18510), .ZN(
        n18520) );
  AOI22_X1 U20495 ( .A1(n18514), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18538), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18518) );
  AOI22_X1 U20496 ( .A1(n13916), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11157), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18517) );
  AOI22_X1 U20497 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18539), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18515) );
  NAND4_X1 U20498 ( .A1(n18518), .A2(n18517), .A3(n18516), .A4(n18515), .ZN(
        n18519) );
  NOR2_X1 U20499 ( .A1(n18520), .A2(n18519), .ZN(n21434) );
  OAI22_X1 U20500 ( .A1(n18536), .A2(n18521), .B1(n21434), .B2(n18562), .ZN(
        P3_U2685) );
  AOI22_X1 U20501 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18522), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18527) );
  AOI22_X1 U20502 ( .A1(n18393), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11157), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18526) );
  AOI22_X1 U20503 ( .A1(n18540), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11151), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18525) );
  AOI22_X1 U20504 ( .A1(n18523), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n20948), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18524) );
  NAND4_X1 U20505 ( .A1(n18527), .A2(n18526), .A3(n18525), .A4(n18524), .ZN(
        n18534) );
  AOI22_X1 U20506 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18546), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18532) );
  AOI22_X1 U20507 ( .A1(n13798), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18547), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18531) );
  AOI22_X1 U20508 ( .A1(n11159), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18528), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18530) );
  AOI22_X1 U20509 ( .A1(n13916), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18538), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18529) );
  NAND4_X1 U20510 ( .A1(n18532), .A2(n18531), .A3(n18530), .A4(n18529), .ZN(
        n18533) );
  NOR2_X1 U20511 ( .A1(n18534), .A2(n18533), .ZN(n21429) );
  OAI21_X1 U20512 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n18536), .A(n18535), .ZN(
        n18537) );
  AOI22_X1 U20513 ( .A1(n18565), .A2(n21429), .B1(n18537), .B2(n18562), .ZN(
        P3_U2684) );
  AOI22_X1 U20514 ( .A1(n13798), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11157), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18544) );
  AOI22_X1 U20515 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18539), .B1(
        n18538), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18543) );
  AOI22_X1 U20516 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20948), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n18540), .ZN(n18542) );
  AOI22_X1 U20517 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n11151), .ZN(n18541) );
  NAND4_X1 U20518 ( .A1(n18544), .A2(n18543), .A3(n18542), .A4(n18541), .ZN(
        n18554) );
  AOI22_X1 U20519 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18545), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n13899), .ZN(n18552) );
  AOI22_X1 U20520 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18497), .B1(
        n18546), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18551) );
  AOI22_X1 U20521 ( .A1(n18548), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18547), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18550) );
  AOI22_X1 U20522 ( .A1(n13916), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n11159), .ZN(n18549) );
  NAND4_X1 U20523 ( .A1(n18552), .A2(n18551), .A3(n18550), .A4(n18549), .ZN(
        n18553) );
  NOR2_X1 U20524 ( .A1(n18554), .A2(n18553), .ZN(n21439) );
  AOI211_X1 U20525 ( .C1(n21129), .C2(n18556), .A(n18555), .B(n18567), .ZN(
        n18557) );
  AOI21_X1 U20526 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n18564), .A(n18557), .ZN(
        n18558) );
  OAI21_X1 U20527 ( .B1(n21439), .B2(n18562), .A(n18558), .ZN(P3_U2686) );
  NOR2_X1 U20528 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n20927) );
  NOR2_X1 U20529 ( .A1(n20927), .A2(n18559), .ZN(n20907) );
  AOI22_X1 U20530 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(n18564), .B1(n18560), .B2(
        n20907), .ZN(n18561) );
  OAI21_X1 U20531 ( .B1(n18563), .B2(n18562), .A(n18561), .ZN(P3_U2702) );
  AOI22_X1 U20532 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18565), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n18564), .ZN(n18566) );
  OAI21_X1 U20533 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n18567), .A(n18566), .ZN(
        P3_U2703) );
  OAI21_X1 U20534 ( .B1(n18569), .B2(n18568), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n18570) );
  OAI21_X1 U20535 ( .B1(n18571), .B2(n21960), .A(n18570), .ZN(P3_U2634) );
  INV_X1 U20536 ( .A(n18979), .ZN(n18575) );
  OAI21_X1 U20537 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n18573), .A(n18572), .ZN(
        n21958) );
  OAI21_X1 U20538 ( .B1(n20833), .B2(n18575), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18574) );
  OAI221_X1 U20539 ( .B1(n18575), .B2(n21958), .C1(n18575), .C2(n19497), .A(
        n18574), .ZN(P3_U2863) );
  AOI22_X1 U20540 ( .A1(n21869), .A2(n18962), .B1(n21720), .B2(n18883), .ZN(
        n18576) );
  INV_X1 U20541 ( .A(n18576), .ZN(n18617) );
  AOI21_X1 U20542 ( .B1(n18826), .B2(n21877), .A(n18617), .ZN(n18829) );
  NAND2_X1 U20543 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18609) );
  NOR2_X4 U20544 ( .A1(n18600), .A2(n18609), .ZN(n21122) );
  NAND2_X2 U20545 ( .A1(n21122), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n21134) );
  NOR2_X1 U20546 ( .A1(n21134), .A2(n20902), .ZN(n18817) );
  INV_X2 U20547 ( .A(n19813), .ZN(n19814) );
  OR2_X1 U20548 ( .A1(n18726), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18578) );
  AOI21_X1 U20549 ( .B1(n18728), .B2(n21134), .A(n18957), .ZN(n18820) );
  OAI211_X1 U20550 ( .C1(n18817), .C2(n18969), .A(n18578), .B(n18820), .ZN(
        n18592) );
  NOR2_X1 U20551 ( .A1(n18726), .A2(n21134), .ZN(n18581) );
  INV_X1 U20552 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n21888) );
  INV_X1 U20553 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18579) );
  NAND2_X1 U20554 ( .A1(n18594), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n21147) );
  OAI21_X1 U20555 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18817), .A(
        n21147), .ZN(n21138) );
  OAI22_X1 U20556 ( .A1(n14030), .A2(n21888), .B1(n18734), .B2(n21138), .ZN(
        n18580) );
  AOI221_X1 U20557 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18592), .C1(
        n18581), .C2(n18592), .A(n18580), .ZN(n18584) );
  AOI21_X1 U20558 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18755), .A(
        n18670), .ZN(n18582) );
  XNOR2_X1 U20559 ( .A(n18582), .B(n18587), .ZN(n21886) );
  NOR2_X1 U20560 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n21877), .ZN(
        n21885) );
  AOI22_X1 U20561 ( .A1(n18870), .A2(n21886), .B1(n18826), .B2(n21885), .ZN(
        n18583) );
  OAI211_X1 U20562 ( .C1(n18829), .C2(n18585), .A(n18584), .B(n18583), .ZN(
        P3_U2812) );
  NOR2_X1 U20563 ( .A1(n18845), .A2(n18586), .ZN(n18669) );
  NOR2_X1 U20564 ( .A1(n18588), .A2(n18587), .ZN(n18661) );
  NOR2_X1 U20565 ( .A1(n18669), .A2(n18661), .ZN(n18589) );
  XNOR2_X1 U20566 ( .A(n21854), .B(n18589), .ZN(n21857) );
  NAND2_X1 U20567 ( .A1(n18591), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n21562) );
  NOR2_X1 U20568 ( .A1(n21720), .A2(n21562), .ZN(n21849) );
  NOR2_X1 U20569 ( .A1(n21869), .A2(n21562), .ZN(n21848) );
  OAI22_X1 U20570 ( .A1(n21849), .A2(n18839), .B1(n21848), .B2(n18974), .ZN(
        n18678) );
  INV_X1 U20571 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18593) );
  CLKBUF_X1 U20572 ( .A(n18648), .Z(n21165) );
  AOI21_X1 U20573 ( .B1(n18593), .B2(n21147), .A(n21165), .ZN(n21149) );
  INV_X1 U20574 ( .A(n21149), .ZN(n18597) );
  AOI22_X1 U20575 ( .A1(n11153), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18592), .ZN(n18596) );
  INV_X1 U20576 ( .A(n18726), .ZN(n18775) );
  NAND3_X1 U20577 ( .A1(n18594), .A2(n18593), .A3(n18775), .ZN(n18595) );
  OAI211_X1 U20578 ( .C1(n18597), .C2(n18734), .A(n18596), .B(n18595), .ZN(
        n18598) );
  AOI221_X1 U20579 ( .B1(n18740), .B2(n21854), .C1(n18678), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n18598), .ZN(n18599) );
  OAI21_X1 U20580 ( .B1(n21857), .B2(n18881), .A(n18599), .ZN(P3_U2811) );
  NOR2_X1 U20581 ( .A1(n18600), .A2(n20902), .ZN(n21094) );
  NAND2_X1 U20582 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n21094), .ZN(
        n18607) );
  OAI21_X1 U20583 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n21094), .A(
        n18607), .ZN(n21099) );
  AOI21_X1 U20584 ( .B1(n18728), .B2(n18600), .A(n18957), .ZN(n18843) );
  OAI21_X1 U20585 ( .B1(n21094), .B2(n18969), .A(n18843), .ZN(n18614) );
  AOI22_X1 U20586 ( .A1(n11153), .A2(P3_REIP_REG_15__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18614), .ZN(n18606) );
  NOR2_X1 U20587 ( .A1(n18643), .A2(n21718), .ZN(n18604) );
  NAND4_X1 U20588 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n21074), .A3(
        n18624), .A4(n18775), .ZN(n18611) );
  INV_X1 U20589 ( .A(n18848), .ZN(n18866) );
  NOR3_X1 U20590 ( .A1(n21684), .A2(n21697), .A3(n18866), .ZN(n18835) );
  NAND2_X1 U20591 ( .A1(n18601), .A2(n18622), .ZN(n18638) );
  NOR3_X1 U20592 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n18638), .ZN(n18836) );
  AOI22_X1 U20593 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18835), .B1(
        n18836), .B2(n21693), .ZN(n18602) );
  XOR2_X1 U20594 ( .A(n18602), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Z(
        n21728) );
  OAI22_X1 U20595 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18611), .B1(
        n21728), .B2(n18881), .ZN(n18603) );
  AOI221_X1 U20596 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18617), 
        .C1(n18604), .C2(n18617), .A(n18603), .ZN(n18605) );
  OAI211_X1 U20597 ( .C1(n18734), .C2(n21099), .A(n18606), .B(n18605), .ZN(
        P3_U2815) );
  INV_X1 U20598 ( .A(n18826), .ZN(n18620) );
  INV_X1 U20599 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n21906) );
  NOR2_X1 U20600 ( .A1(n14030), .A2(n21906), .ZN(n18613) );
  INV_X1 U20601 ( .A(n18607), .ZN(n18608) );
  NAND2_X1 U20602 ( .A1(n21122), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18818) );
  OAI21_X1 U20603 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18608), .A(
        n18818), .ZN(n21106) );
  OAI21_X1 U20604 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18609), .ZN(n18610) );
  OAI22_X1 U20605 ( .A1(n18734), .A2(n21106), .B1(n18611), .B2(n18610), .ZN(
        n18612) );
  AOI211_X1 U20606 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n18614), .A(
        n18613), .B(n18612), .ZN(n18619) );
  AOI22_X1 U20607 ( .A1(n18755), .A2(n21902), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18845), .ZN(n18615) );
  XNOR2_X1 U20608 ( .A(n18616), .B(n18615), .ZN(n21904) );
  AOI22_X1 U20609 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18617), .B1(
        n18870), .B2(n21904), .ZN(n18618) );
  OAI211_X1 U20610 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n18620), .A(
        n18619), .B(n18618), .ZN(P3_U2814) );
  NAND2_X1 U20611 ( .A1(n21671), .A2(n18848), .ZN(n18621) );
  OAI21_X1 U20612 ( .B1(n18622), .B2(n18621), .A(n18638), .ZN(n18623) );
  XOR2_X1 U20613 ( .A(n18623), .B(n21688), .Z(n21692) );
  NAND2_X1 U20614 ( .A1(n18624), .A2(n18775), .ZN(n18632) );
  NAND2_X1 U20615 ( .A1(n11153), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n21690) );
  OAI21_X1 U20616 ( .B1(n18624), .B2(n18933), .A(n18969), .ZN(n18625) );
  AOI21_X1 U20617 ( .B1(n18626), .B2(n18625), .A(n18957), .ZN(n18635) );
  INV_X1 U20618 ( .A(n18635), .ZN(n18627) );
  NOR2_X1 U20619 ( .A1(n18633), .A2(n18626), .ZN(n18831) );
  AOI21_X1 U20620 ( .B1(n18633), .B2(n18626), .A(n18831), .ZN(n21056) );
  AOI22_X1 U20621 ( .A1(n18627), .A2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n18808), .B2(n21056), .ZN(n18628) );
  OAI211_X1 U20622 ( .C1(n18632), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n21690), .B(n18628), .ZN(n18629) );
  INV_X1 U20623 ( .A(n18629), .ZN(n18631) );
  OAI21_X1 U20624 ( .B1(n21681), .B2(n18643), .A(n18873), .ZN(n18640) );
  OAI221_X1 U20625 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n21685), 
        .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18869), .A(n18640), .ZN(
        n18630) );
  OAI211_X1 U20626 ( .C1(n21692), .C2(n18881), .A(n18631), .B(n18630), .ZN(
        P3_U2818) );
  NAND2_X1 U20627 ( .A1(n21681), .A2(n21697), .ZN(n21915) );
  AOI211_X1 U20628 ( .C1(n18633), .C2(n18634), .A(n21074), .B(n18632), .ZN(
        n18637) );
  INV_X1 U20629 ( .A(n18831), .ZN(n21067) );
  AOI22_X1 U20630 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n21067), .B1(
        n18831), .B2(n18634), .ZN(n21075) );
  OAI22_X1 U20631 ( .A1(n18635), .A2(n18634), .B1(n18734), .B2(n21075), .ZN(
        n18636) );
  AOI211_X1 U20632 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n11153), .A(n18637), 
        .B(n18636), .ZN(n18642) );
  OAI22_X1 U20633 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18638), .B1(
        n18866), .B2(n21684), .ZN(n18639) );
  XOR2_X1 U20634 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18639), .Z(
        n21908) );
  AOI22_X1 U20635 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18640), .B1(
        n18870), .B2(n21908), .ZN(n18641) );
  OAI211_X1 U20636 ( .C1(n18643), .C2(n21915), .A(n18642), .B(n18641), .ZN(
        P3_U2817) );
  NAND2_X1 U20637 ( .A1(n18741), .A2(n18740), .ZN(n18654) );
  INV_X1 U20638 ( .A(n21566), .ZN(n18692) );
  INV_X1 U20639 ( .A(n21567), .ZN(n18706) );
  AOI22_X1 U20640 ( .A1(n18962), .A2(n18692), .B1(n18883), .B2(n18706), .ZN(
        n18667) );
  NOR2_X1 U20641 ( .A1(n18645), .A2(n18644), .ZN(n18647) );
  OAI21_X1 U20642 ( .B1(n18647), .B2(n18646), .A(n18668), .ZN(n18694) );
  XOR2_X1 U20643 ( .A(n21737), .B(n18694), .Z(n21729) );
  INV_X1 U20644 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18659) );
  NOR2_X1 U20645 ( .A1(n18672), .A2(n18659), .ZN(n18655) );
  NAND2_X1 U20646 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18684) );
  NOR2_X2 U20647 ( .A1(n18672), .A2(n18684), .ZN(n18685) );
  INV_X1 U20648 ( .A(n18685), .ZN(n18681) );
  OAI21_X1 U20649 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18655), .A(
        n18681), .ZN(n21190) );
  INV_X1 U20650 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n21169) );
  OR2_X1 U20651 ( .A1(n18675), .A2(n21169), .ZN(n18683) );
  OAI21_X1 U20652 ( .B1(n21165), .B2(n18969), .A(n18970), .ZN(n18649) );
  AOI21_X1 U20653 ( .B1(n18728), .B2(n18683), .A(n18649), .ZN(n18674) );
  OAI21_X1 U20654 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18776), .A(
        n18674), .ZN(n18658) );
  AOI22_X1 U20655 ( .A1(n11153), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18658), .ZN(n18651) );
  NOR2_X1 U20656 ( .A1(n18726), .A2(n18683), .ZN(n18660) );
  OAI211_X1 U20657 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n18660), .B(n18684), .ZN(n18650) );
  OAI211_X1 U20658 ( .C1(n21190), .C2(n18734), .A(n18651), .B(n18650), .ZN(
        n18652) );
  AOI21_X1 U20659 ( .B1(n18870), .B2(n21729), .A(n18652), .ZN(n18653) );
  OAI221_X1 U20660 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18654), 
        .C1(n21737), .C2(n18667), .A(n18653), .ZN(P3_U2808) );
  INV_X1 U20661 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18666) );
  AOI21_X1 U20662 ( .B1(n18672), .B2(n18659), .A(n18655), .ZN(n21184) );
  AOI22_X1 U20663 ( .A1(n11153), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18808), 
        .B2(n21184), .ZN(n18656) );
  INV_X1 U20664 ( .A(n18656), .ZN(n18657) );
  AOI221_X1 U20665 ( .B1(n18660), .B2(n18659), .C1(n18658), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n18657), .ZN(n18665) );
  NOR2_X1 U20666 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18662) );
  AOI22_X1 U20667 ( .A1(n21570), .A2(n18669), .B1(n18662), .B2(n18661), .ZN(
        n18663) );
  XOR2_X1 U20668 ( .A(n18666), .B(n18663), .Z(n21574) );
  INV_X1 U20669 ( .A(n21570), .ZN(n21569) );
  NOR2_X1 U20670 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n21569), .ZN(
        n21573) );
  AOI22_X1 U20671 ( .A1(n18870), .A2(n21574), .B1(n18740), .B2(n21573), .ZN(
        n18664) );
  OAI211_X1 U20672 ( .C1(n18667), .C2(n18666), .A(n18665), .B(n18664), .ZN(
        P3_U2809) );
  OAI221_X1 U20673 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18670), 
        .C1(n21854), .C2(n18669), .A(n18668), .ZN(n18671) );
  XNOR2_X1 U20674 ( .A(n21863), .B(n18671), .ZN(n21867) );
  OAI21_X1 U20675 ( .B1(n21165), .B2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n18672), .ZN(n18673) );
  INV_X1 U20676 ( .A(n18673), .ZN(n21168) );
  INV_X1 U20677 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n21163) );
  NOR2_X1 U20678 ( .A1(n14030), .A2(n21163), .ZN(n21860) );
  AOI221_X1 U20679 ( .B1(n18675), .B2(n21169), .C1(n19813), .C2(n21169), .A(
        n18674), .ZN(n18676) );
  AOI211_X1 U20680 ( .C1(n21168), .C2(n18963), .A(n21860), .B(n18676), .ZN(
        n18680) );
  NOR2_X1 U20681 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21562), .ZN(
        n18677) );
  AOI22_X1 U20682 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18678), .B1(
        n18826), .B2(n18677), .ZN(n18679) );
  OAI211_X1 U20683 ( .C1(n18881), .C2(n21867), .A(n18680), .B(n18679), .ZN(
        P3_U2810) );
  AOI22_X1 U20684 ( .A1(n18962), .A2(n21825), .B1(n18883), .B2(n21827), .ZN(
        n18720) );
  INV_X1 U20685 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n21218) );
  NOR2_X4 U20686 ( .A1(n18681), .A2(n21218), .ZN(n18712) );
  AOI21_X1 U20687 ( .B1(n18681), .B2(n21218), .A(n18712), .ZN(n21213) );
  NAND2_X1 U20688 ( .A1(n21218), .A2(n18682), .ZN(n18700) );
  INV_X1 U20689 ( .A(n18700), .ZN(n18690) );
  NOR2_X1 U20690 ( .A1(n18684), .A2(n18683), .ZN(n18687) );
  NAND2_X1 U20691 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18687), .ZN(
        n18724) );
  OAI21_X1 U20692 ( .B1(n18685), .B2(n18969), .A(n18970), .ZN(n18686) );
  AOI21_X1 U20693 ( .B1(n19814), .B2(n18724), .A(n18686), .ZN(n18701) );
  AOI21_X1 U20694 ( .B1(n19814), .B2(n18687), .A(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18688) );
  INV_X1 U20695 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n21839) );
  OAI22_X1 U20696 ( .A1(n18701), .A2(n18688), .B1(n14030), .B2(n21839), .ZN(
        n18689) );
  AOI221_X1 U20697 ( .B1(n18808), .B2(n21213), .C1(n18690), .C2(n21213), .A(
        n18689), .ZN(n18699) );
  NAND2_X1 U20698 ( .A1(n18883), .A2(n21827), .ZN(n18693) );
  NAND2_X1 U20699 ( .A1(n18962), .A2(n21825), .ZN(n18691) );
  OAI22_X1 U20700 ( .A1(n18706), .A2(n18693), .B1(n18692), .B2(n18691), .ZN(
        n18697) );
  AOI221_X1 U20701 ( .B1(n21737), .B2(n18695), .C1(n18845), .C2(n18695), .A(
        n18694), .ZN(n18696) );
  XOR2_X1 U20702 ( .A(n18696), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(
        n21837) );
  AOI22_X1 U20703 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18697), .B1(
        n18870), .B2(n21837), .ZN(n18698) );
  OAI211_X1 U20704 ( .C1(n18720), .C2(n21833), .A(n18699), .B(n18698), .ZN(
        P3_U2807) );
  NAND2_X1 U20705 ( .A1(n18701), .A2(n18700), .ZN(n18715) );
  INV_X1 U20706 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n21239) );
  NAND2_X1 U20707 ( .A1(n18712), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18703) );
  NAND2_X1 U20708 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18725) );
  INV_X1 U20709 ( .A(n18725), .ZN(n18702) );
  AOI21_X1 U20710 ( .B1(n21239), .B2(n18703), .A(n18765), .ZN(n21236) );
  AOI22_X1 U20711 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18715), .B1(
        n18808), .B2(n21236), .ZN(n18711) );
  INV_X1 U20712 ( .A(n18736), .ZN(n18704) );
  AOI22_X1 U20713 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18736), .B1(
        n18704), .B2(n21762), .ZN(n21753) );
  NAND3_X1 U20714 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n18705), .ZN(n18739) );
  OAI22_X1 U20715 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18737), .B1(
        n18739), .B2(n18706), .ZN(n21748) );
  OAI21_X1 U20716 ( .B1(n18845), .B2(n18761), .A(n11515), .ZN(n18707) );
  XOR2_X1 U20717 ( .A(n18707), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n21750) );
  OAI22_X1 U20718 ( .A1(n18839), .A2(n21748), .B1(n18881), .B2(n21750), .ZN(
        n18708) );
  AOI21_X1 U20719 ( .B1(n18962), .B2(n21753), .A(n18708), .ZN(n18710) );
  NAND2_X1 U20720 ( .A1(n11153), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n21754) );
  NOR2_X1 U20721 ( .A1(n18726), .A2(n18724), .ZN(n18717) );
  OAI211_X1 U20722 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18717), .B(n18725), .ZN(n18709) );
  NAND4_X1 U20723 ( .A1(n18711), .A2(n18710), .A3(n21754), .A4(n18709), .ZN(
        P3_U2805) );
  INV_X1 U20724 ( .A(n18712), .ZN(n18713) );
  INV_X1 U20725 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18716) );
  OAI22_X1 U20726 ( .A1(n18713), .A2(n18716), .B1(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18712), .ZN(n21220) );
  INV_X1 U20727 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n21225) );
  NOR2_X1 U20728 ( .A1(n14030), .A2(n21225), .ZN(n18714) );
  AOI221_X1 U20729 ( .B1(n18717), .B2(n18716), .C1(n18715), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n18714), .ZN(n18723) );
  NOR2_X1 U20730 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21739), .ZN(
        n21840) );
  AOI21_X1 U20731 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18719), .A(
        n18718), .ZN(n21846) );
  OAI22_X1 U20732 ( .A1(n18720), .A2(n21740), .B1(n21846), .B2(n18881), .ZN(
        n18721) );
  AOI21_X1 U20733 ( .B1(n18740), .B2(n21840), .A(n18721), .ZN(n18722) );
  OAI211_X1 U20734 ( .C1(n18734), .C2(n21220), .A(n18723), .B(n18722), .ZN(
        P3_U2806) );
  NOR2_X1 U20735 ( .A1(n18725), .A2(n18724), .ZN(n18763) );
  NAND2_X1 U20736 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18763), .ZN(
        n18730) );
  NOR3_X1 U20737 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18726), .A3(
        n18730), .ZN(n18756) );
  OAI21_X1 U20738 ( .B1(n18765), .B2(n18969), .A(n18970), .ZN(n18727) );
  AOI21_X1 U20739 ( .B1(n18728), .B2(n18730), .A(n18727), .ZN(n18767) );
  OAI21_X1 U20740 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18776), .A(
        n18767), .ZN(n18752) );
  NAND2_X2 U20741 ( .A1(n11522), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n18764) );
  INV_X1 U20742 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18751) );
  NOR2_X4 U20743 ( .A1(n18764), .A2(n18751), .ZN(n18750) );
  NAND2_X2 U20744 ( .A1(n18750), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n18807) );
  OAI21_X1 U20745 ( .B1(n18750), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n18807), .ZN(n21271) );
  INV_X1 U20746 ( .A(n18729), .ZN(n18733) );
  NOR2_X1 U20747 ( .A1(n18751), .A2(n18730), .ZN(n18774) );
  INV_X1 U20748 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n18731) );
  NAND3_X1 U20749 ( .A1(n18774), .A2(n18731), .A3(n18775), .ZN(n18732) );
  OAI211_X1 U20750 ( .C1(n18734), .C2(n21271), .A(n18733), .B(n18732), .ZN(
        n18735) );
  AOI221_X1 U20751 ( .B1(n18756), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C1(
        n18752), .C2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n18735), .ZN(
        n18749) );
  NAND2_X1 U20752 ( .A1(n18738), .A2(n18736), .ZN(n21758) );
  NAND2_X1 U20753 ( .A1(n18738), .A2(n18737), .ZN(n21777) );
  AOI22_X1 U20754 ( .A1(n18962), .A2(n21758), .B1(n18883), .B2(n21777), .ZN(
        n18770) );
  NAND2_X1 U20755 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18770), .ZN(
        n18757) );
  OAI211_X1 U20756 ( .C1(n18962), .C2(n18883), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18757), .ZN(n18748) );
  INV_X1 U20757 ( .A(n18739), .ZN(n21756) );
  NAND3_X1 U20758 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18793), .A3(
        n18742), .ZN(n18747) );
  OAI211_X1 U20759 ( .C1(n18745), .C2(n18744), .A(n18870), .B(n18743), .ZN(
        n18746) );
  NAND4_X1 U20760 ( .A1(n18749), .A2(n18748), .A3(n18747), .A4(n18746), .ZN(
        P3_U2802) );
  AOI21_X1 U20761 ( .B1(n18764), .B2(n18751), .A(n18750), .ZN(n21264) );
  AOI22_X1 U20762 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n18752), .B1(
        n18808), .B2(n21264), .ZN(n18760) );
  OAI21_X1 U20763 ( .B1(n18755), .B2(n18754), .A(n18753), .ZN(n21771) );
  AOI21_X1 U20764 ( .B1(n18870), .B2(n21771), .A(n18756), .ZN(n18759) );
  OAI21_X1 U20765 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18793), .A(
        n18757), .ZN(n18758) );
  NAND2_X1 U20766 ( .A1(n11153), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n21784) );
  NAND4_X1 U20767 ( .A1(n18760), .A2(n18759), .A3(n18758), .A4(n21784), .ZN(
        P3_U2803) );
  OAI221_X1 U20768 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18845), 
        .C1(n21762), .C2(n18761), .A(n11515), .ZN(n18762) );
  XOR2_X1 U20769 ( .A(n21760), .B(n18762), .Z(n21767) );
  INV_X1 U20770 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n21260) );
  NOR2_X1 U20771 ( .A1(n14030), .A2(n21260), .ZN(n21766) );
  AOI21_X1 U20772 ( .B1(n19814), .B2(n18763), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n18766) );
  OAI21_X1 U20773 ( .B1(n18765), .B2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n18764), .ZN(n21247) );
  OAI22_X1 U20774 ( .A1(n18767), .A2(n18766), .B1(n18955), .B2(n21247), .ZN(
        n18768) );
  AOI211_X1 U20775 ( .C1(n21767), .C2(n18870), .A(n21766), .B(n18768), .ZN(
        n18769) );
  OAI221_X1 U20776 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n18771), 
        .C1(n21760), .C2(n18770), .A(n18769), .ZN(P3_U2804) );
  NAND2_X1 U20777 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21814) );
  NOR2_X1 U20778 ( .A1(n21814), .A2(n18796), .ZN(n18772) );
  INV_X1 U20779 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n21812) );
  XOR2_X1 U20780 ( .A(n18772), .B(n21812), .Z(n21817) );
  INV_X1 U20781 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n21299) );
  NAND2_X1 U20782 ( .A1(n18806), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n18773) );
  INV_X1 U20783 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n21319) );
  NAND2_X1 U20784 ( .A1(n11153), .A2(P3_REIP_REG_31__SCAN_IN), .ZN(n21822) );
  INV_X1 U20785 ( .A(n21822), .ZN(n18782) );
  NAND2_X1 U20786 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18774), .ZN(
        n18803) );
  NOR2_X1 U20787 ( .A1(n21299), .A2(n18803), .ZN(n18777) );
  NAND2_X1 U20788 ( .A1(n18777), .A2(n18775), .ZN(n18792) );
  XNOR2_X1 U20789 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n18780) );
  NOR2_X1 U20790 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18776), .ZN(
        n18809) );
  INV_X1 U20791 ( .A(n18807), .ZN(n18778) );
  OAI22_X1 U20792 ( .A1(n18969), .A2(n18778), .B1(n19813), .B2(n18777), .ZN(
        n18779) );
  OR2_X1 U20793 ( .A1(n18779), .A2(n18957), .ZN(n18805) );
  NOR2_X1 U20794 ( .A1(n18809), .A2(n18805), .ZN(n18790) );
  OAI22_X1 U20795 ( .A1(n18792), .A2(n18780), .B1(n18790), .B2(n21319), .ZN(
        n18781) );
  AOI211_X1 U20796 ( .C1(n21146), .C2(n18808), .A(n18782), .B(n18781), .ZN(
        n18786) );
  INV_X1 U20797 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21798) );
  NAND3_X1 U20798 ( .A1(n18801), .A2(n18800), .A3(n21798), .ZN(n18787) );
  OAI22_X1 U20799 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18787), .B1(
        n18788), .B2(n21814), .ZN(n18783) );
  XNOR2_X1 U20800 ( .A(n21812), .B(n18783), .ZN(n21821) );
  NOR2_X1 U20801 ( .A1(n18795), .A2(n21814), .ZN(n18784) );
  XNOR2_X1 U20802 ( .A(n21812), .B(n18784), .ZN(n21820) );
  AOI22_X1 U20803 ( .A1(n18870), .A2(n21821), .B1(n18962), .B2(n21820), .ZN(
        n18785) );
  OAI211_X1 U20804 ( .C1(n21817), .C2(n18839), .A(n18786), .B(n18785), .ZN(
        P3_U2799) );
  OAI21_X1 U20805 ( .B1(n18788), .B2(n21798), .A(n18787), .ZN(n18789) );
  INV_X1 U20806 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21803) );
  XOR2_X1 U20807 ( .A(n18789), .B(n21803), .Z(n21811) );
  INV_X1 U20808 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n18791) );
  XNOR2_X1 U20809 ( .A(n18791), .B(n18806), .ZN(n21314) );
  NAND2_X1 U20810 ( .A1(n11153), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n21809) );
  OAI221_X1 U20811 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n18792), .C1(
        n18791), .C2(n18790), .A(n21809), .ZN(n18798) );
  NAND3_X1 U20812 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21804) );
  NOR2_X1 U20813 ( .A1(n21804), .A2(n18794), .ZN(n18797) );
  INV_X1 U20814 ( .A(n18795), .ZN(n21793) );
  NAND2_X1 U20815 ( .A1(n21793), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n21789) );
  AOI21_X1 U20816 ( .B1(n21794), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n18839), .ZN(n18813) );
  AOI21_X1 U20817 ( .B1(n18962), .B2(n21789), .A(n18813), .ZN(n18816) );
  AOI21_X1 U20818 ( .B1(n21793), .B2(n18962), .A(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n18815) );
  AOI21_X1 U20819 ( .B1(n18801), .B2(n18800), .A(n18799), .ZN(n18802) );
  XOR2_X1 U20820 ( .A(n18802), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n21801) );
  OAI21_X1 U20821 ( .B1(n19813), .B2(n18803), .A(n21299), .ZN(n18804) );
  AOI22_X1 U20822 ( .A1(n11153), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n18805), 
        .B2(n18804), .ZN(n18811) );
  AOI21_X1 U20823 ( .B1(n18807), .B2(n21299), .A(n18806), .ZN(n21293) );
  OAI21_X1 U20824 ( .B1(n18809), .B2(n18808), .A(n21293), .ZN(n18810) );
  OAI211_X1 U20825 ( .C1(n21801), .C2(n18881), .A(n18811), .B(n18810), .ZN(
        n18812) );
  AOI21_X1 U20826 ( .B1(n21794), .B2(n18813), .A(n18812), .ZN(n18814) );
  OAI21_X1 U20827 ( .B1(n18816), .B2(n18815), .A(n18814), .ZN(P3_U2801) );
  INV_X1 U20828 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18819) );
  AOI21_X1 U20829 ( .B1(n18819), .B2(n18818), .A(n18817), .ZN(n21123) );
  INV_X1 U20830 ( .A(n21123), .ZN(n18822) );
  AOI21_X1 U20831 ( .B1(n21122), .B2(n19814), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18821) );
  OAI22_X1 U20832 ( .A1(n18955), .A2(n18822), .B1(n18821), .B2(n18820), .ZN(
        n18823) );
  AOI21_X1 U20833 ( .B1(n11153), .B2(P3_REIP_REG_17__SCAN_IN), .A(n18823), 
        .ZN(n18828) );
  OAI21_X1 U20834 ( .B1(n18825), .B2(n21882), .A(n18824), .ZN(n21892) );
  NOR2_X1 U20835 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21902), .ZN(
        n21891) );
  AOI22_X1 U20836 ( .A1(n18870), .A2(n21892), .B1(n18826), .B2(n21891), .ZN(
        n18827) );
  OAI211_X1 U20837 ( .C1(n18829), .C2(n21882), .A(n18828), .B(n18827), .ZN(
        P3_U2813) );
  AOI21_X1 U20838 ( .B1(n21074), .B2(n18830), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18844) );
  INV_X1 U20839 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18833) );
  NAND2_X1 U20840 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n18831), .ZN(
        n18832) );
  AOI21_X1 U20841 ( .B1(n18833), .B2(n18832), .A(n21094), .ZN(n21080) );
  AOI22_X1 U20842 ( .A1(n11153), .A2(P3_REIP_REG_14__SCAN_IN), .B1(n21080), 
        .B2(n18963), .ZN(n18842) );
  AOI21_X1 U20843 ( .B1(n21693), .B2(n18834), .A(n21724), .ZN(n21706) );
  NOR2_X1 U20844 ( .A1(n18836), .A2(n18835), .ZN(n18837) );
  XOR2_X1 U20845 ( .A(n18837), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n21710) );
  AND2_X1 U20846 ( .A1(n21928), .A2(n21700), .ZN(n18838) );
  NAND3_X1 U20847 ( .A1(n21928), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n21700), .ZN(n21714) );
  OAI21_X1 U20848 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18838), .A(
        n21714), .ZN(n21705) );
  OAI22_X1 U20849 ( .A1(n21710), .A2(n18881), .B1(n18839), .B2(n21705), .ZN(
        n18840) );
  AOI21_X1 U20850 ( .B1(n18962), .B2(n21706), .A(n18840), .ZN(n18841) );
  OAI211_X1 U20851 ( .C1(n18844), .C2(n18843), .A(n18842), .B(n18841), .ZN(
        P3_U2816) );
  INV_X1 U20852 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21916) );
  INV_X1 U20853 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21942) );
  AOI21_X1 U20854 ( .B1(n18845), .B2(n21942), .A(n18848), .ZN(n18846) );
  AOI211_X1 U20855 ( .C1(n21942), .C2(n18847), .A(n18846), .B(n21916), .ZN(
        n18850) );
  NOR3_X1 U20856 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18848), .A3(
        n21942), .ZN(n18849) );
  AOI211_X1 U20857 ( .C1(n18851), .C2(n18867), .A(n18850), .B(n18849), .ZN(
        n21917) );
  INV_X1 U20858 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n21033) );
  NOR2_X1 U20859 ( .A1(n14030), .A2(n21033), .ZN(n18857) );
  NOR2_X1 U20860 ( .A1(n18886), .A2(n19813), .ZN(n18889) );
  NAND3_X1 U20861 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(n18889), .ZN(n18863) );
  NOR2_X1 U20862 ( .A1(n18862), .A2(n18863), .ZN(n18861) );
  AOI21_X1 U20863 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18964), .A(
        n18861), .ZN(n18854) );
  NOR2_X1 U20864 ( .A1(n18862), .A2(n18874), .ZN(n21014) );
  INV_X1 U20865 ( .A(n18852), .ZN(n18853) );
  OAI21_X1 U20866 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n21014), .A(
        n18853), .ZN(n21028) );
  OAI22_X1 U20867 ( .A1(n18855), .A2(n18854), .B1(n18955), .B2(n21028), .ZN(
        n18856) );
  AOI211_X1 U20868 ( .C1(n21917), .C2(n18870), .A(n18857), .B(n18856), .ZN(
        n18860) );
  NAND3_X1 U20869 ( .A1(n21675), .A2(n18858), .A3(n18869), .ZN(n18859) );
  OAI211_X1 U20870 ( .C1(n18873), .C2(n21916), .A(n18860), .B(n18859), .ZN(
        P3_U2820) );
  AOI21_X1 U20871 ( .B1(n18862), .B2(n18874), .A(n21014), .ZN(n21018) );
  AOI211_X1 U20872 ( .C1(n18863), .C2(n18862), .A(n18908), .B(n18861), .ZN(
        n18865) );
  INV_X1 U20873 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n21025) );
  NOR2_X1 U20874 ( .A1(n14030), .A2(n21025), .ZN(n18864) );
  AOI211_X1 U20875 ( .C1(n21018), .C2(n18963), .A(n18865), .B(n18864), .ZN(
        n18872) );
  NAND2_X1 U20876 ( .A1(n18867), .A2(n18866), .ZN(n18868) );
  XOR2_X1 U20877 ( .A(n18868), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n21938) );
  AOI22_X1 U20878 ( .A1(n18870), .A2(n21938), .B1(n21942), .B2(n18869), .ZN(
        n18871) );
  OAI211_X1 U20879 ( .C1(n18873), .C2(n21942), .A(n18872), .B(n18871), .ZN(
        P3_U2821) );
  OAI21_X1 U20880 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18887), .A(
        n18874), .ZN(n21003) );
  OAI21_X1 U20881 ( .B1(n20970), .B2(n18933), .A(n18970), .ZN(n18897) );
  INV_X1 U20882 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20998) );
  NOR2_X1 U20883 ( .A1(n14030), .A2(n20998), .ZN(n21663) );
  AOI221_X1 U20884 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C1(n21000), .C2(n21007), .A(n19813), .ZN(n18875) );
  AOI211_X1 U20885 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18897), .A(
        n21663), .B(n18875), .ZN(n18885) );
  OAI21_X1 U20886 ( .B1(n18878), .B2(n18877), .A(n18876), .ZN(n21660) );
  OAI21_X1 U20887 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18880), .A(
        n18879), .ZN(n21665) );
  OAI22_X1 U20888 ( .A1(n18974), .A2(n21665), .B1(n18881), .B2(n21660), .ZN(
        n18882) );
  AOI21_X1 U20889 ( .B1(n18883), .B2(n21660), .A(n18882), .ZN(n18884) );
  OAI211_X1 U20890 ( .C1(n18955), .C2(n21003), .A(n18885), .B(n18884), .ZN(
        P3_U2822) );
  NOR2_X1 U20891 ( .A1(n18886), .A2(n20902), .ZN(n18910) );
  INV_X1 U20892 ( .A(n18887), .ZN(n18888) );
  OAI21_X1 U20893 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18910), .A(
        n18888), .ZN(n20981) );
  AOI22_X1 U20894 ( .A1(n11153), .A2(P3_REIP_REG_7__SCAN_IN), .B1(n18889), 
        .B2(n20984), .ZN(n18899) );
  OAI21_X1 U20895 ( .B1(n18892), .B2(n18891), .A(n18890), .ZN(n18893) );
  XOR2_X1 U20896 ( .A(n18893), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n21643) );
  OAI21_X1 U20897 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18895), .A(
        n18894), .ZN(n21654) );
  OAI22_X1 U20898 ( .A1(n18974), .A2(n21643), .B1(n18973), .B2(n21654), .ZN(
        n18896) );
  AOI21_X1 U20899 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18897), .A(
        n18896), .ZN(n18898) );
  OAI211_X1 U20900 ( .C1(n18955), .C2(n20981), .A(n18899), .B(n18898), .ZN(
        P3_U2823) );
  OAI21_X1 U20901 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18901), .A(
        n18900), .ZN(n21635) );
  CLKBUF_X1 U20902 ( .A(n18902), .Z(n18909) );
  NAND2_X1 U20903 ( .A1(n18909), .A2(n19814), .ZN(n18906) );
  OAI21_X1 U20904 ( .B1(n18905), .B2(n18904), .A(n18903), .ZN(n21636) );
  OAI22_X1 U20905 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18906), .B1(
        n18973), .B2(n21636), .ZN(n18907) );
  AOI21_X1 U20906 ( .B1(n11153), .B2(P3_REIP_REG_6__SCAN_IN), .A(n18907), .ZN(
        n18913) );
  AOI21_X1 U20907 ( .B1(n19814), .B2(n18909), .A(n18908), .ZN(n18923) );
  INV_X1 U20908 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18911) );
  NAND2_X1 U20909 ( .A1(n18909), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18917) );
  AOI21_X1 U20910 ( .B1(n18911), .B2(n18917), .A(n18910), .ZN(n20973) );
  AOI22_X1 U20911 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18923), .B1(
        n20973), .B2(n18963), .ZN(n18912) );
  OAI211_X1 U20912 ( .C1(n18974), .C2(n21635), .A(n18913), .B(n18912), .ZN(
        P3_U2824) );
  OAI21_X1 U20913 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18915), .A(
        n18914), .ZN(n21628) );
  OAI21_X1 U20914 ( .B1(n18957), .B2(n20943), .A(n18916), .ZN(n18922) );
  NOR2_X1 U20915 ( .A1(n20943), .A2(n20902), .ZN(n18935) );
  OAI21_X1 U20916 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18935), .A(
        n18917), .ZN(n20963) );
  OAI21_X1 U20917 ( .B1(n18920), .B2(n18919), .A(n18918), .ZN(n21627) );
  OAI22_X1 U20918 ( .A1(n18955), .A2(n20963), .B1(n18974), .B2(n21627), .ZN(
        n18921) );
  AOI21_X1 U20919 ( .B1(n18923), .B2(n18922), .A(n18921), .ZN(n18924) );
  NAND2_X1 U20920 ( .A1(n11153), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n21631) );
  OAI211_X1 U20921 ( .C1(n18973), .C2(n21628), .A(n18924), .B(n21631), .ZN(
        P3_U2825) );
  OAI21_X1 U20922 ( .B1(n18927), .B2(n18926), .A(n18925), .ZN(n21612) );
  NOR2_X1 U20923 ( .A1(n19813), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18932) );
  INV_X1 U20924 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20960) );
  OAI21_X1 U20925 ( .B1(n18930), .B2(n18929), .A(n18928), .ZN(n21613) );
  OAI22_X1 U20926 ( .A1(n14030), .A2(n20960), .B1(n18973), .B2(n21613), .ZN(
        n18931) );
  AOI21_X1 U20927 ( .B1(n18932), .B2(n18934), .A(n18931), .ZN(n18937) );
  OAI21_X1 U20928 ( .B1(n18934), .B2(n18933), .A(n18970), .ZN(n18947) );
  INV_X1 U20929 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20951) );
  NAND2_X1 U20930 ( .A1(n18934), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18941) );
  AOI21_X1 U20931 ( .B1(n20951), .B2(n18941), .A(n18935), .ZN(n20947) );
  AOI22_X1 U20932 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18947), .B1(
        n20947), .B2(n18963), .ZN(n18936) );
  OAI211_X1 U20933 ( .C1(n18974), .C2(n21612), .A(n18937), .B(n18936), .ZN(
        P3_U2826) );
  OAI21_X1 U20934 ( .B1(n18940), .B2(n18939), .A(n18938), .ZN(n21607) );
  INV_X1 U20935 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20920) );
  NOR2_X1 U20936 ( .A1(n18957), .A2(n20920), .ZN(n18946) );
  NOR2_X1 U20937 ( .A1(n20920), .A2(n20902), .ZN(n20916) );
  OAI21_X1 U20938 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n20916), .A(
        n18941), .ZN(n20937) );
  OAI21_X1 U20939 ( .B1(n18944), .B2(n18943), .A(n18942), .ZN(n21606) );
  OAI22_X1 U20940 ( .A1(n18955), .A2(n20937), .B1(n18974), .B2(n21606), .ZN(
        n18945) );
  AOI221_X1 U20941 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18947), .C1(
        n18946), .C2(n18947), .A(n18945), .ZN(n18948) );
  NAND2_X1 U20942 ( .A1(n11153), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n21610) );
  OAI211_X1 U20943 ( .C1(n18973), .C2(n21607), .A(n18948), .B(n21610), .ZN(
        P3_U2827) );
  OAI21_X1 U20944 ( .B1(n18951), .B2(n18950), .A(n18949), .ZN(n21599) );
  AOI21_X1 U20945 ( .B1(n20920), .B2(n20902), .A(n20916), .ZN(n20918) );
  INV_X1 U20946 ( .A(n20918), .ZN(n20919) );
  OAI21_X1 U20947 ( .B1(n18954), .B2(n18953), .A(n18952), .ZN(n21595) );
  OAI22_X1 U20948 ( .A1(n18955), .A2(n20919), .B1(n18973), .B2(n21595), .ZN(
        n18956) );
  AOI221_X1 U20949 ( .B1(n18957), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n19814), .C2(n20920), .A(n18956), .ZN(n18958) );
  NAND2_X1 U20950 ( .A1(n11153), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n21597) );
  OAI211_X1 U20951 ( .C1(n18974), .C2(n21599), .A(n18958), .B(n21597), .ZN(
        P3_U2828) );
  OAI21_X1 U20952 ( .B1(n18967), .B2(n18960), .A(n18959), .ZN(n21590) );
  NAND2_X1 U20953 ( .A1(n21732), .A2(n18968), .ZN(n18961) );
  XNOR2_X1 U20954 ( .A(n18961), .B(n18960), .ZN(n21586) );
  AOI22_X1 U20955 ( .A1(n11153), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18962), 
        .B2(n21586), .ZN(n18966) );
  AOI22_X1 U20956 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18964), .B1(
        n18963), .B2(n20902), .ZN(n18965) );
  OAI211_X1 U20957 ( .C1(n18973), .C2(n21590), .A(n18966), .B(n18965), .ZN(
        P3_U2829) );
  AOI21_X1 U20958 ( .B1(n18968), .B2(n21732), .A(n18967), .ZN(n21582) );
  INV_X1 U20959 ( .A(n21582), .ZN(n21581) );
  NAND3_X1 U20960 ( .A1(n21537), .A2(n18970), .A3(n18969), .ZN(n18971) );
  AOI22_X1 U20961 ( .A1(n11153), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18971), .ZN(n18972) );
  OAI221_X1 U20962 ( .B1(n21582), .B2(n18974), .C1(n21581), .C2(n18973), .A(
        n18972), .ZN(P3_U2830) );
  NAND2_X1 U20963 ( .A1(n19523), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19508) );
  INV_X1 U20964 ( .A(n19508), .ZN(n19510) );
  NAND2_X1 U20965 ( .A1(n19522), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19531) );
  INV_X1 U20966 ( .A(n19531), .ZN(n19532) );
  NOR2_X1 U20967 ( .A1(n19510), .A2(n19532), .ZN(n18976) );
  OAI22_X1 U20968 ( .A1(n18977), .A2(n19522), .B1(n18976), .B2(n18975), .ZN(
        P3_U2866) );
  NAND2_X1 U20969 ( .A1(n18979), .A2(n18978), .ZN(n18983) );
  OAI21_X1 U20970 ( .B1(n18981), .B2(n18980), .A(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18982) );
  OAI21_X1 U20971 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18983), .A(
        n18982), .ZN(P3_U2864) );
  NOR4_X1 U20972 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18987) );
  NOR4_X1 U20973 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18986) );
  NOR4_X1 U20974 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18985) );
  NOR4_X1 U20975 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18984) );
  NAND4_X1 U20976 ( .A1(n18987), .A2(n18986), .A3(n18985), .A4(n18984), .ZN(
        n18993) );
  NOR4_X1 U20977 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18991) );
  AOI211_X1 U20978 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18990) );
  NOR4_X1 U20979 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18989) );
  NOR4_X1 U20980 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18988) );
  NAND4_X1 U20981 ( .A1(n18991), .A2(n18990), .A3(n18989), .A4(n18988), .ZN(
        n18992) );
  NOR2_X1 U20982 ( .A1(n18993), .A2(n18992), .ZN(n19005) );
  INV_X1 U20983 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18995) );
  OAI21_X1 U20984 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n19005), .ZN(n18994) );
  OAI21_X1 U20985 ( .B1(n19005), .B2(n18995), .A(n18994), .ZN(P3_U3293) );
  INV_X1 U20986 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18998) );
  AOI21_X1 U20987 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18996) );
  INV_X1 U20988 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n20923) );
  OAI221_X1 U20989 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18996), .C1(n20923), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n19005), .ZN(n18997) );
  OAI21_X1 U20990 ( .B1(n19005), .B2(n18998), .A(n18997), .ZN(P3_U3292) );
  INV_X1 U20991 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19000) );
  NOR3_X1 U20992 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19001) );
  OAI21_X1 U20993 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n19001), .A(n19005), .ZN(
        n18999) );
  OAI21_X1 U20994 ( .B1(n19005), .B2(n19000), .A(n18999), .ZN(P3_U2638) );
  INV_X1 U20995 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22317) );
  AOI21_X1 U20996 ( .B1(n20923), .B2(n22317), .A(n19001), .ZN(n19004) );
  INV_X1 U20997 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19003) );
  INV_X1 U20998 ( .A(n19005), .ZN(n19002) );
  AOI22_X1 U20999 ( .A1(n19005), .A2(n19004), .B1(n19003), .B2(n19002), .ZN(
        P3_U2639) );
  OAI22_X1 U21000 ( .A1(n19068), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n22321), .ZN(n19006) );
  INV_X1 U21001 ( .A(n19006), .ZN(P3_U3297) );
  INV_X1 U21002 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19007) );
  AOI22_X1 U21003 ( .A1(n22321), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19007), 
        .B2(n19068), .ZN(P3_U3294) );
  AOI21_X1 U21004 ( .B1(n22356), .B2(n22361), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n19008) );
  AOI22_X1 U21005 ( .A1(n22321), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n19008), 
        .B2(n19068), .ZN(P3_U2635) );
  INV_X1 U21006 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n21530) );
  AOI22_X1 U21007 ( .A1(n19015), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n19009) );
  OAI21_X1 U21008 ( .B1(n21530), .B2(n19026), .A(n19009), .ZN(P3_U2767) );
  INV_X1 U21009 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n21518) );
  AOI22_X1 U21010 ( .A1(n19015), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n19010) );
  OAI21_X1 U21011 ( .B1(n21518), .B2(n19026), .A(n19010), .ZN(P3_U2766) );
  INV_X1 U21012 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n20872) );
  AOI22_X1 U21013 ( .A1(n19015), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n19011) );
  OAI21_X1 U21014 ( .B1(n20872), .B2(n19026), .A(n19011), .ZN(P3_U2765) );
  INV_X1 U21015 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n20874) );
  AOI22_X1 U21016 ( .A1(n19015), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n19037), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n19012) );
  OAI21_X1 U21017 ( .B1(n20874), .B2(n19026), .A(n19012), .ZN(P3_U2764) );
  INV_X1 U21018 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n21370) );
  AOI22_X1 U21019 ( .A1(n19015), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n19037), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n19013) );
  OAI21_X1 U21020 ( .B1(n21370), .B2(n19026), .A(n19013), .ZN(P3_U2763) );
  INV_X1 U21021 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n21343) );
  AOI22_X1 U21022 ( .A1(n19015), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n19037), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n19014) );
  OAI21_X1 U21023 ( .B1(n21343), .B2(n19026), .A(n19014), .ZN(P3_U2762) );
  INV_X1 U21024 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n21371) );
  AOI22_X1 U21025 ( .A1(n19015), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n19037), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n19016) );
  OAI21_X1 U21026 ( .B1(n21371), .B2(n19026), .A(n19016), .ZN(P3_U2761) );
  INV_X1 U21027 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n21342) );
  AOI22_X1 U21029 ( .A1(n19015), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n19017) );
  OAI21_X1 U21030 ( .B1(n21342), .B2(n19026), .A(n19017), .ZN(P3_U2760) );
  INV_X1 U21031 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n21509) );
  AOI22_X1 U21032 ( .A1(n19015), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n19018) );
  OAI21_X1 U21033 ( .B1(n21509), .B2(n19026), .A(n19018), .ZN(P3_U2759) );
  INV_X1 U21034 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n21400) );
  AOI22_X1 U21035 ( .A1(n19015), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n19019) );
  OAI21_X1 U21036 ( .B1(n21400), .B2(n19026), .A(n19019), .ZN(P3_U2758) );
  INV_X1 U21037 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n20883) );
  AOI22_X1 U21038 ( .A1(n19015), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n19020) );
  OAI21_X1 U21039 ( .B1(n20883), .B2(n19026), .A(n19020), .ZN(P3_U2757) );
  INV_X1 U21040 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n21351) );
  AOI22_X1 U21041 ( .A1(n19015), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n19021) );
  OAI21_X1 U21042 ( .B1(n21351), .B2(n19026), .A(n19021), .ZN(P3_U2756) );
  INV_X1 U21043 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n21350) );
  AOI22_X1 U21044 ( .A1(n19015), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n19022) );
  OAI21_X1 U21045 ( .B1(n21350), .B2(n19026), .A(n19022), .ZN(P3_U2755) );
  INV_X1 U21046 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n20887) );
  AOI22_X1 U21047 ( .A1(n19015), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n19023) );
  OAI21_X1 U21048 ( .B1(n20887), .B2(n19026), .A(n19023), .ZN(P3_U2754) );
  INV_X1 U21049 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n21501) );
  AOI22_X1 U21050 ( .A1(n19015), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n19024) );
  OAI21_X1 U21051 ( .B1(n21501), .B2(n19026), .A(n19024), .ZN(P3_U2753) );
  INV_X1 U21052 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n21504) );
  AOI22_X1 U21053 ( .A1(n19015), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n19025) );
  OAI21_X1 U21054 ( .B1(n21504), .B2(n19026), .A(n19025), .ZN(P3_U2752) );
  INV_X1 U21055 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n20845) );
  NAND2_X1 U21056 ( .A1(n19028), .A2(n19027), .ZN(n19047) );
  AOI22_X1 U21057 ( .A1(n19015), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n19029) );
  OAI21_X1 U21058 ( .B1(n20845), .B2(n19047), .A(n19029), .ZN(P3_U2751) );
  INV_X1 U21059 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n21416) );
  AOI22_X1 U21060 ( .A1(n19015), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n19030) );
  OAI21_X1 U21061 ( .B1(n21416), .B2(n19047), .A(n19030), .ZN(P3_U2750) );
  INV_X1 U21062 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n20848) );
  AOI22_X1 U21063 ( .A1(n19015), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n19031) );
  OAI21_X1 U21064 ( .B1(n20848), .B2(n19047), .A(n19031), .ZN(P3_U2749) );
  INV_X1 U21065 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n21425) );
  AOI22_X1 U21066 ( .A1(n19015), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n19037), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n19032) );
  OAI21_X1 U21067 ( .B1(n21425), .B2(n19047), .A(n19032), .ZN(P3_U2748) );
  INV_X1 U21068 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n21417) );
  AOI22_X1 U21069 ( .A1(n19015), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n19037), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n19033) );
  OAI21_X1 U21070 ( .B1(n21417), .B2(n19047), .A(n19033), .ZN(P3_U2747) );
  INV_X1 U21071 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n21415) );
  AOI22_X1 U21072 ( .A1(n19015), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n19037), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n19034) );
  OAI21_X1 U21073 ( .B1(n21415), .B2(n19047), .A(n19034), .ZN(P3_U2746) );
  INV_X1 U21074 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n21441) );
  AOI22_X1 U21075 ( .A1(n19015), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n19037), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n19035) );
  OAI21_X1 U21076 ( .B1(n21441), .B2(n19047), .A(n19035), .ZN(P3_U2745) );
  INV_X1 U21077 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n20855) );
  AOI22_X1 U21078 ( .A1(n19015), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n19037), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n19036) );
  OAI21_X1 U21079 ( .B1(n20855), .B2(n19047), .A(n19036), .ZN(P3_U2744) );
  INV_X1 U21080 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n20857) );
  AOI22_X1 U21081 ( .A1(n19015), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n19037), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n19038) );
  OAI21_X1 U21082 ( .B1(n20857), .B2(n19047), .A(n19038), .ZN(P3_U2743) );
  INV_X1 U21083 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20859) );
  AOI22_X1 U21084 ( .A1(n19015), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n19039) );
  OAI21_X1 U21085 ( .B1(n20859), .B2(n19047), .A(n19039), .ZN(P3_U2742) );
  INV_X1 U21086 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n21450) );
  AOI22_X1 U21087 ( .A1(n19015), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n19040) );
  OAI21_X1 U21088 ( .B1(n21450), .B2(n19047), .A(n19040), .ZN(P3_U2741) );
  INV_X1 U21089 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n20863) );
  AOI22_X1 U21090 ( .A1(n19015), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n19041) );
  OAI21_X1 U21091 ( .B1(n20863), .B2(n19047), .A(n19041), .ZN(P3_U2740) );
  INV_X1 U21092 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n20865) );
  AOI22_X1 U21093 ( .A1(n19015), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n19042) );
  OAI21_X1 U21094 ( .B1(n20865), .B2(n19047), .A(n19042), .ZN(P3_U2739) );
  INV_X1 U21095 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n21463) );
  AOI22_X1 U21096 ( .A1(n19015), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n19043) );
  OAI21_X1 U21097 ( .B1(n21463), .B2(n19047), .A(n19043), .ZN(P3_U2738) );
  INV_X1 U21098 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n20868) );
  AOI22_X1 U21099 ( .A1(n19015), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n19044), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n19046) );
  OAI21_X1 U21100 ( .B1(n20868), .B2(n19047), .A(n19046), .ZN(P3_U2737) );
  NOR2_X1 U21101 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(n19048), .ZN(n19049) );
  NOR2_X1 U21102 ( .A1(n22321), .A2(n19049), .ZN(P3_U2633) );
  NOR2_X1 U21103 ( .A1(n19068), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19060) );
  INV_X1 U21104 ( .A(n19060), .ZN(n19064) );
  INV_X1 U21105 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n20924) );
  INV_X1 U21106 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n20552) );
  OAI222_X1 U21107 ( .A1(n19064), .A2(n20924), .B1(n20552), .B2(n22321), .C1(
        n20923), .C2(n19059), .ZN(P3_U3032) );
  AOI22_X1 U21108 ( .A1(n19060), .A2(P3_REIP_REG_3__SCAN_IN), .B1(
        P3_ADDRESS_REG_1__SCAN_IN), .B2(n19068), .ZN(n19050) );
  OAI21_X1 U21109 ( .B1(n22359), .B2(n20924), .A(n19050), .ZN(P3_U3033) );
  AOI22_X1 U21110 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n19062), .B1(
        P3_ADDRESS_REG_2__SCAN_IN), .B2(n19068), .ZN(n19051) );
  OAI21_X1 U21111 ( .B1(n20960), .B2(n19064), .A(n19051), .ZN(P3_U3034) );
  AOI22_X1 U21112 ( .A1(n19060), .A2(P3_REIP_REG_5__SCAN_IN), .B1(
        P3_ADDRESS_REG_3__SCAN_IN), .B2(n19068), .ZN(n19052) );
  OAI21_X1 U21113 ( .B1(n22359), .B2(n20960), .A(n19052), .ZN(P3_U3035) );
  INV_X1 U21114 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20992) );
  AOI22_X1 U21115 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n19062), .B1(
        P3_ADDRESS_REG_4__SCAN_IN), .B2(n19068), .ZN(n19053) );
  OAI21_X1 U21116 ( .B1(n20992), .B2(n19064), .A(n19053), .ZN(P3_U3036) );
  INV_X1 U21117 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n20993) );
  INV_X1 U21118 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n20558) );
  OAI222_X1 U21119 ( .A1(n19064), .A2(n20993), .B1(n20558), .B2(n22321), .C1(
        n20992), .C2(n19059), .ZN(P3_U3037) );
  INV_X1 U21120 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n20560) );
  OAI222_X1 U21121 ( .A1(n19064), .A2(n20998), .B1(n20560), .B2(n22321), .C1(
        n20993), .C2(n19059), .ZN(P3_U3038) );
  INV_X1 U21122 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n20562) );
  OAI222_X1 U21123 ( .A1(n19064), .A2(n21025), .B1(n20562), .B2(n22321), .C1(
        n20998), .C2(n19059), .ZN(P3_U3039) );
  INV_X1 U21124 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n20564) );
  OAI222_X1 U21125 ( .A1(n21025), .A2(n22359), .B1(n20564), .B2(n22321), .C1(
        n21033), .C2(n19064), .ZN(P3_U3040) );
  INV_X1 U21126 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n20566) );
  OAI222_X1 U21127 ( .A1(n21033), .A2(n22359), .B1(n20566), .B2(n22321), .C1(
        n19054), .C2(n19064), .ZN(P3_U3041) );
  INV_X1 U21128 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n20568) );
  INV_X1 U21129 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n21062) );
  OAI222_X1 U21130 ( .A1(n19054), .A2(n22359), .B1(n20568), .B2(n22321), .C1(
        n21062), .C2(n19064), .ZN(P3_U3042) );
  INV_X1 U21131 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n21068) );
  INV_X1 U21132 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n20570) );
  OAI222_X1 U21133 ( .A1(n19064), .A2(n21068), .B1(n20570), .B2(n22321), .C1(
        n21062), .C2(n22359), .ZN(P3_U3043) );
  INV_X1 U21134 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n21082) );
  INV_X1 U21135 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n20572) );
  OAI222_X1 U21136 ( .A1(n19064), .A2(n21082), .B1(n20572), .B2(n22321), .C1(
        n21068), .C2(n22359), .ZN(P3_U3044) );
  AOI22_X1 U21137 ( .A1(n19060), .A2(P3_REIP_REG_15__SCAN_IN), .B1(
        P3_ADDRESS_REG_13__SCAN_IN), .B2(n19068), .ZN(n19055) );
  OAI21_X1 U21138 ( .B1(n22359), .B2(n21082), .A(n19055), .ZN(P3_U3045) );
  AOI22_X1 U21139 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n19062), .B1(
        P3_ADDRESS_REG_14__SCAN_IN), .B2(n19068), .ZN(n19056) );
  OAI21_X1 U21140 ( .B1(n21906), .B2(n19064), .A(n19056), .ZN(P3_U3046) );
  INV_X1 U21141 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n21894) );
  INV_X1 U21142 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n20576) );
  OAI222_X1 U21143 ( .A1(n19064), .A2(n21894), .B1(n20576), .B2(n22321), .C1(
        n21906), .C2(n22359), .ZN(P3_U3047) );
  INV_X1 U21144 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n20578) );
  OAI222_X1 U21145 ( .A1(n19064), .A2(n21888), .B1(n20578), .B2(n22321), .C1(
        n21894), .C2(n22359), .ZN(P3_U3048) );
  INV_X1 U21146 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n21156) );
  INV_X1 U21147 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n20580) );
  OAI222_X1 U21148 ( .A1(n19064), .A2(n21156), .B1(n20580), .B2(n22321), .C1(
        n21888), .C2(n22359), .ZN(P3_U3049) );
  INV_X1 U21149 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n20582) );
  OAI222_X1 U21150 ( .A1(n19064), .A2(n21163), .B1(n20582), .B2(n22321), .C1(
        n21156), .C2(n22359), .ZN(P3_U3050) );
  INV_X1 U21151 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n21576) );
  INV_X1 U21152 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n20584) );
  OAI222_X1 U21153 ( .A1(n19064), .A2(n21576), .B1(n20584), .B2(n22321), .C1(
        n21163), .C2(n19059), .ZN(P3_U3051) );
  AOI22_X1 U21154 ( .A1(n19060), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_ADDRESS_REG_20__SCAN_IN), .B2(n19068), .ZN(n19057) );
  OAI21_X1 U21155 ( .B1(n19059), .B2(n21576), .A(n19057), .ZN(P3_U3052) );
  AOI22_X1 U21156 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n19062), .B1(
        P3_ADDRESS_REG_21__SCAN_IN), .B2(n19068), .ZN(n19058) );
  OAI21_X1 U21157 ( .B1(n21839), .B2(n19064), .A(n19058), .ZN(P3_U3053) );
  INV_X1 U21158 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n20588) );
  OAI222_X1 U21159 ( .A1(n21839), .A2(n22359), .B1(n20588), .B2(n22321), .C1(
        n21225), .C2(n19064), .ZN(P3_U3054) );
  INV_X1 U21160 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n21261) );
  INV_X1 U21161 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n20590) );
  OAI222_X1 U21162 ( .A1(n19064), .A2(n21261), .B1(n20590), .B2(n22321), .C1(
        n21225), .C2(n19059), .ZN(P3_U3055) );
  INV_X1 U21163 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n20592) );
  OAI222_X1 U21164 ( .A1(n21261), .A2(n22359), .B1(n20592), .B2(n22321), .C1(
        n21260), .C2(n19064), .ZN(P3_U3056) );
  INV_X1 U21165 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n21270) );
  INV_X1 U21166 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n20594) );
  OAI222_X1 U21167 ( .A1(n19064), .A2(n21270), .B1(n20594), .B2(n22321), .C1(
        n21260), .C2(n19059), .ZN(P3_U3057) );
  INV_X1 U21168 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n20596) );
  OAI222_X1 U21169 ( .A1(n19064), .A2(n21275), .B1(n20596), .B2(n22321), .C1(
        n21270), .C2(n19059), .ZN(P3_U3058) );
  INV_X1 U21170 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n20598) );
  INV_X1 U21171 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n21283) );
  OAI222_X1 U21172 ( .A1(n21275), .A2(n22359), .B1(n20598), .B2(n22321), .C1(
        n21283), .C2(n19064), .ZN(P3_U3059) );
  AOI22_X1 U21173 ( .A1(n19060), .A2(P3_REIP_REG_30__SCAN_IN), .B1(
        P3_ADDRESS_REG_28__SCAN_IN), .B2(n19068), .ZN(n19061) );
  OAI21_X1 U21174 ( .B1(n22359), .B2(n21283), .A(n19061), .ZN(P3_U3060) );
  INV_X1 U21175 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n21315) );
  AOI22_X1 U21176 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n19062), .B1(
        P3_ADDRESS_REG_29__SCAN_IN), .B2(n19068), .ZN(n19063) );
  OAI21_X1 U21177 ( .B1(n21315), .B2(n19064), .A(n19063), .ZN(P3_U3061) );
  OAI22_X1 U21178 ( .A1(n19068), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n22321), .ZN(n19065) );
  INV_X1 U21179 ( .A(n19065), .ZN(P3_U3277) );
  OAI22_X1 U21180 ( .A1(n19068), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n22321), .ZN(n19066) );
  INV_X1 U21181 ( .A(n19066), .ZN(P3_U3276) );
  OAI22_X1 U21182 ( .A1(n19068), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n22321), .ZN(n19067) );
  INV_X1 U21183 ( .A(n19067), .ZN(P3_U3275) );
  OAI22_X1 U21184 ( .A1(n19068), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n22321), .ZN(n19069) );
  INV_X1 U21185 ( .A(n19069), .ZN(P3_U3274) );
  NOR4_X1 U21186 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n19072)
         );
  INV_X1 U21187 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n19070) );
  NOR4_X1 U21188 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n19070), .ZN(n19071) );
  NAND3_X1 U21189 ( .A1(n19072), .A2(n19071), .A3(U215), .ZN(U213) );
  NAND4_X1 U21190 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .A3(n19436), .A4(n19073), .ZN(n19076) );
  INV_X1 U21191 ( .A(n19074), .ZN(n19075) );
  OAI211_X1 U21192 ( .C1(n19078), .C2(n19077), .A(n19076), .B(n19075), .ZN(
        n19089) );
  INV_X1 U21193 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19088) );
  NOR2_X1 U21194 ( .A1(n22338), .A2(n19999), .ZN(n19082) );
  NAND4_X1 U21195 ( .A1(n19080), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n22347), 
        .A4(n19079), .ZN(n19081) );
  OAI21_X1 U21196 ( .B1(n19082), .B2(n19434), .A(n19081), .ZN(n19086) );
  AOI211_X1 U21197 ( .C1(P2_STATEBS16_REG_SCAN_IN), .C2(n19084), .A(n19436), 
        .B(n19083), .ZN(n19085) );
  OAI21_X1 U21198 ( .B1(n19086), .B2(n19085), .A(n19089), .ZN(n19087) );
  OAI21_X1 U21199 ( .B1(n19089), .B2(n19088), .A(n19087), .ZN(P2_U3610) );
  NAND2_X1 U21200 ( .A1(n19316), .A2(n16057), .ZN(n19353) );
  OAI22_X1 U21201 ( .A1(n16338), .A2(n19338), .B1(n19336), .B2(n19366), .ZN(
        n19090) );
  INV_X1 U21202 ( .A(n19090), .ZN(n19095) );
  NAND2_X1 U21203 ( .A1(n12300), .A2(n19349), .ZN(n19094) );
  NAND2_X1 U21204 ( .A1(n19328), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n19093) );
  NAND2_X1 U21205 ( .A1(n19323), .A2(n19091), .ZN(n19092) );
  AND4_X1 U21206 ( .A1(n19095), .A2(n19094), .A3(n19093), .A4(n19092), .ZN(
        n19099) );
  NAND2_X1 U21207 ( .A1(n11181), .A2(n19316), .ZN(n19282) );
  INV_X1 U21208 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19096) );
  AOI21_X1 U21209 ( .B1(n19237), .B2(n19282), .A(n19096), .ZN(n19097) );
  AOI21_X1 U21210 ( .B1(n19110), .B2(n20081), .A(n19097), .ZN(n19098) );
  OAI211_X1 U21211 ( .C1(n19100), .C2(n19353), .A(n19099), .B(n19098), .ZN(
        P2_U2855) );
  AOI22_X1 U21212 ( .A1(n19323), .A2(n19101), .B1(P2_EBX_REG_1__SCAN_IN), .B2(
        n19328), .ZN(n19109) );
  INV_X1 U21213 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19102) );
  OAI22_X1 U21214 ( .A1(n19336), .A2(n19103), .B1(n19237), .B2(n19102), .ZN(
        n19104) );
  INV_X1 U21215 ( .A(n19104), .ZN(n19108) );
  NAND2_X1 U21216 ( .A1(n19105), .A2(n19349), .ZN(n19107) );
  NAND2_X1 U21217 ( .A1(n19307), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n19106) );
  AND4_X1 U21218 ( .A1(n19109), .A2(n19108), .A3(n19107), .A4(n19106), .ZN(
        n19113) );
  AOI22_X1 U21219 ( .A1(n19111), .A2(n19316), .B1(n19944), .B2(n19110), .ZN(
        n19112) );
  OAI211_X1 U21220 ( .C1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19282), .A(
        n19113), .B(n19112), .ZN(P2_U2854) );
  INV_X1 U21221 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n19117) );
  OAI22_X1 U21222 ( .A1(n19342), .A2(n19114), .B1(n19237), .B2(n12256), .ZN(
        n19115) );
  INV_X1 U21223 ( .A(n19115), .ZN(n19116) );
  OAI21_X1 U21224 ( .B1(n19188), .B2(n19117), .A(n19116), .ZN(n19118) );
  AOI211_X1 U21225 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19307), .A(n19407), .B(
        n19118), .ZN(n19126) );
  NAND2_X1 U21226 ( .A1(n19263), .A2(n19119), .ZN(n19120) );
  XNOR2_X1 U21227 ( .A(n19121), .B(n19120), .ZN(n19124) );
  INV_X1 U21228 ( .A(n19122), .ZN(n19123) );
  AOI22_X1 U21229 ( .A1(n19124), .A2(n19316), .B1(n19349), .B2(n19123), .ZN(
        n19125) );
  OAI211_X1 U21230 ( .C1(n19336), .C2(n20170), .A(n19126), .B(n19125), .ZN(
        P2_U2850) );
  NOR2_X1 U21231 ( .A1(n11181), .A2(n19127), .ZN(n19128) );
  XOR2_X1 U21232 ( .A(n19129), .B(n19128), .Z(n19138) );
  INV_X1 U21233 ( .A(n19130), .ZN(n19131) );
  AOI22_X1 U21234 ( .A1(n19323), .A2(n19131), .B1(P2_EBX_REG_6__SCAN_IN), .B2(
        n19328), .ZN(n19132) );
  OAI211_X1 U21235 ( .C1(n11754), .C2(n19338), .A(n19132), .B(n19258), .ZN(
        n19136) );
  OAI22_X1 U21236 ( .A1(n19134), .A2(n19336), .B1(n19310), .B2(n19133), .ZN(
        n19135) );
  AOI211_X1 U21237 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19346), .A(
        n19136), .B(n19135), .ZN(n19137) );
  OAI21_X1 U21238 ( .B1(n19432), .B2(n19138), .A(n19137), .ZN(P2_U2849) );
  NAND2_X1 U21239 ( .A1(n19263), .A2(n19139), .ZN(n19141) );
  XOR2_X1 U21240 ( .A(n19141), .B(n19140), .Z(n19149) );
  AOI22_X1 U21241 ( .A1(n19142), .A2(n19323), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n19328), .ZN(n19143) );
  OAI211_X1 U21242 ( .C1(n11757), .C2(n19338), .A(n19143), .B(n19258), .ZN(
        n19147) );
  OAI22_X1 U21243 ( .A1(n19145), .A2(n19336), .B1(n19310), .B2(n19144), .ZN(
        n19146) );
  AOI211_X1 U21244 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19346), .A(
        n19147), .B(n19146), .ZN(n19148) );
  OAI21_X1 U21245 ( .B1(n19149), .B2(n19432), .A(n19148), .ZN(P2_U2848) );
  OAI21_X1 U21246 ( .B1(n11763), .B2(n19338), .A(n19258), .ZN(n19153) );
  OAI22_X1 U21247 ( .A1(n19151), .A2(n19342), .B1(n19188), .B2(n19150), .ZN(
        n19152) );
  AOI211_X1 U21248 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19346), .A(
        n19153), .B(n19152), .ZN(n19160) );
  NAND2_X1 U21249 ( .A1(n19263), .A2(n19154), .ZN(n19155) );
  XNOR2_X1 U21250 ( .A(n19156), .B(n19155), .ZN(n19158) );
  AOI22_X1 U21251 ( .A1(n19158), .A2(n19316), .B1(n19157), .B2(n19349), .ZN(
        n19159) );
  OAI211_X1 U21252 ( .C1(n19161), .C2(n19336), .A(n19160), .B(n19159), .ZN(
        P2_U2846) );
  AOI22_X1 U21253 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19346), .B1(
        P2_EBX_REG_10__SCAN_IN), .B2(n19328), .ZN(n19162) );
  OAI21_X1 U21254 ( .B1(n19163), .B2(n19342), .A(n19162), .ZN(n19164) );
  AOI211_X1 U21255 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n19307), .A(n19407), 
        .B(n19164), .ZN(n19171) );
  NOR2_X1 U21256 ( .A1(n11181), .A2(n19165), .ZN(n19167) );
  XNOR2_X1 U21257 ( .A(n19167), .B(n19166), .ZN(n19169) );
  AOI22_X1 U21258 ( .A1(n19169), .A2(n19316), .B1(n19168), .B2(n19349), .ZN(
        n19170) );
  OAI211_X1 U21259 ( .C1(n19172), .C2(n19336), .A(n19171), .B(n19170), .ZN(
        P2_U2845) );
  NAND2_X1 U21260 ( .A1(n19173), .A2(n19349), .ZN(n19175) );
  AOI21_X1 U21261 ( .B1(n19307), .B2(P2_REIP_REG_11__SCAN_IN), .A(n19407), 
        .ZN(n19174) );
  OAI211_X1 U21262 ( .C1(n19336), .C2(n19176), .A(n19175), .B(n19174), .ZN(
        n19179) );
  OAI22_X1 U21263 ( .A1(n19188), .A2(n12199), .B1(n19177), .B2(n19237), .ZN(
        n19178) );
  AOI211_X1 U21264 ( .C1(n19323), .C2(n19180), .A(n19179), .B(n19178), .ZN(
        n19185) );
  INV_X1 U21265 ( .A(n19181), .ZN(n19183) );
  OAI211_X1 U21266 ( .C1(n19183), .C2(n19186), .A(n19316), .B(n19182), .ZN(
        n19184) );
  OAI211_X1 U21267 ( .C1(n19282), .C2(n19186), .A(n19185), .B(n19184), .ZN(
        P2_U2844) );
  OAI21_X1 U21268 ( .B1(n19187), .B2(n19338), .A(n19258), .ZN(n19191) );
  OAI22_X1 U21269 ( .A1(n19189), .A2(n19342), .B1(n12200), .B2(n19188), .ZN(
        n19190) );
  AOI211_X1 U21270 ( .C1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n19346), .A(
        n19191), .B(n19190), .ZN(n19198) );
  NAND2_X1 U21271 ( .A1(n19263), .A2(n19192), .ZN(n19194) );
  XNOR2_X1 U21272 ( .A(n19194), .B(n19193), .ZN(n19196) );
  AOI22_X1 U21273 ( .A1(n19196), .A2(n19316), .B1(n19195), .B2(n19349), .ZN(
        n19197) );
  OAI211_X1 U21274 ( .C1(n19199), .C2(n19336), .A(n19198), .B(n19197), .ZN(
        P2_U2842) );
  NOR2_X1 U21275 ( .A1(n11181), .A2(n19200), .ZN(n19202) );
  XOR2_X1 U21276 ( .A(n19202), .B(n19201), .Z(n19211) );
  AOI22_X1 U21277 ( .A1(P2_EBX_REG_14__SCAN_IN), .A2(n19328), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19346), .ZN(n19203) );
  OAI21_X1 U21278 ( .B1(n19204), .B2(n19342), .A(n19203), .ZN(n19205) );
  AOI211_X1 U21279 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19307), .A(n19407), 
        .B(n19205), .ZN(n19210) );
  INV_X1 U21280 ( .A(n19206), .ZN(n19208) );
  AOI22_X1 U21281 ( .A1(n19208), .A2(n19349), .B1(n19207), .B2(n19348), .ZN(
        n19209) );
  OAI211_X1 U21282 ( .C1(n19432), .C2(n19211), .A(n19210), .B(n19209), .ZN(
        P2_U2841) );
  AOI22_X1 U21283 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(n19328), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n19346), .ZN(n19212) );
  OAI211_X1 U21284 ( .C1(n19219), .C2(n19282), .A(n19212), .B(n19380), .ZN(
        n19213) );
  AOI21_X1 U21285 ( .B1(n19307), .B2(P2_REIP_REG_15__SCAN_IN), .A(n19213), 
        .ZN(n19214) );
  OAI21_X1 U21286 ( .B1(n19215), .B2(n19310), .A(n19214), .ZN(n19216) );
  AOI21_X1 U21287 ( .B1(n11210), .B2(n19323), .A(n19216), .ZN(n19222) );
  INV_X1 U21288 ( .A(n19217), .ZN(n19220) );
  NOR2_X1 U21289 ( .A1(n11181), .A2(n19218), .ZN(n19228) );
  OAI211_X1 U21290 ( .C1(n19220), .C2(n19219), .A(n19316), .B(n19228), .ZN(
        n19221) );
  OAI211_X1 U21291 ( .C1(n19336), .C2(n19223), .A(n19222), .B(n19221), .ZN(
        P2_U2840) );
  AOI22_X1 U21292 ( .A1(P2_EBX_REG_16__SCAN_IN), .A2(n19328), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19346), .ZN(n19224) );
  OAI21_X1 U21293 ( .B1(n19225), .B2(n19342), .A(n19224), .ZN(n19226) );
  AOI211_X1 U21294 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n19307), .A(n19407), 
        .B(n19226), .ZN(n19232) );
  XNOR2_X1 U21295 ( .A(n19228), .B(n19227), .ZN(n19230) );
  AOI22_X1 U21296 ( .A1(n19230), .A2(n19316), .B1(n19229), .B2(n19349), .ZN(
        n19231) );
  OAI211_X1 U21297 ( .C1(n19233), .C2(n19336), .A(n19232), .B(n19231), .ZN(
        P2_U2839) );
  NAND2_X1 U21298 ( .A1(n16057), .A2(n19234), .ZN(n19235) );
  XOR2_X1 U21299 ( .A(n19236), .B(n19235), .Z(n19246) );
  OAI21_X1 U21300 ( .B1(n17585), .B2(n19338), .A(n19258), .ZN(n19240) );
  OAI22_X1 U21301 ( .A1(n19238), .A2(n19342), .B1(n19237), .B2(n12231), .ZN(
        n19239) );
  AOI211_X1 U21302 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19328), .A(n19240), .B(
        n19239), .ZN(n19245) );
  OAI22_X1 U21303 ( .A1(n19242), .A2(n19310), .B1(n19241), .B2(n19336), .ZN(
        n19243) );
  INV_X1 U21304 ( .A(n19243), .ZN(n19244) );
  OAI211_X1 U21305 ( .C1(n19432), .C2(n19246), .A(n19245), .B(n19244), .ZN(
        P2_U2838) );
  NOR2_X1 U21306 ( .A1(n11181), .A2(n19247), .ZN(n19249) );
  XOR2_X1 U21307 ( .A(n19249), .B(n19248), .Z(n19256) );
  AOI22_X1 U21308 ( .A1(n19250), .A2(n19323), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n19328), .ZN(n19251) );
  OAI211_X1 U21309 ( .C1(n17571), .C2(n19338), .A(n19251), .B(n19258), .ZN(
        n19252) );
  AOI21_X1 U21310 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19346), .A(
        n19252), .ZN(n19255) );
  AOI22_X1 U21311 ( .A1(n19253), .A2(n19349), .B1(n20320), .B2(n19348), .ZN(
        n19254) );
  OAI211_X1 U21312 ( .C1(n19432), .C2(n19256), .A(n19255), .B(n19254), .ZN(
        P2_U2837) );
  AOI22_X1 U21313 ( .A1(n19257), .A2(n19323), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n19328), .ZN(n19259) );
  OAI211_X1 U21314 ( .C1(n19260), .C2(n19338), .A(n19259), .B(n19258), .ZN(
        n19261) );
  AOI21_X1 U21315 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19346), .A(
        n19261), .ZN(n19269) );
  NAND2_X1 U21316 ( .A1(n19263), .A2(n19262), .ZN(n19265) );
  XNOR2_X1 U21317 ( .A(n19265), .B(n19264), .ZN(n19267) );
  AOI22_X1 U21318 ( .A1(n19267), .A2(n19316), .B1(n19266), .B2(n19349), .ZN(
        n19268) );
  OAI211_X1 U21319 ( .C1(n19270), .C2(n19336), .A(n19269), .B(n19268), .ZN(
        P2_U2836) );
  AOI22_X1 U21320 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19346), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19307), .ZN(n19271) );
  OAI21_X1 U21321 ( .B1(n19272), .B2(n19342), .A(n19271), .ZN(n19276) );
  INV_X1 U21322 ( .A(n19273), .ZN(n19274) );
  OAI22_X1 U21323 ( .A1(n19274), .A2(n19310), .B1(n20225), .B2(n19336), .ZN(
        n19275) );
  AOI211_X1 U21324 ( .C1(P2_EBX_REG_20__SCAN_IN), .C2(n19328), .A(n19276), .B(
        n19275), .ZN(n19280) );
  OAI211_X1 U21325 ( .C1(n19278), .C2(n19281), .A(n19277), .B(n19316), .ZN(
        n19279) );
  OAI211_X1 U21326 ( .C1(n19282), .C2(n19281), .A(n19280), .B(n19279), .ZN(
        P2_U2835) );
  AOI22_X1 U21327 ( .A1(n19283), .A2(n19323), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19346), .ZN(n19294) );
  AOI22_X1 U21328 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n19328), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19307), .ZN(n19293) );
  OAI22_X1 U21329 ( .A1(n19285), .A2(n19310), .B1(n19284), .B2(n19336), .ZN(
        n19286) );
  INV_X1 U21330 ( .A(n19286), .ZN(n19292) );
  AOI21_X1 U21331 ( .B1(n19289), .B2(n19288), .A(n19287), .ZN(n19290) );
  NAND2_X1 U21332 ( .A1(n19316), .A2(n19290), .ZN(n19291) );
  NAND4_X1 U21333 ( .A1(n19294), .A2(n19293), .A3(n19292), .A4(n19291), .ZN(
        P2_U2831) );
  AOI22_X1 U21334 ( .A1(n19295), .A2(n19323), .B1(P2_REIP_REG_26__SCAN_IN), 
        .B2(n19307), .ZN(n19305) );
  AOI22_X1 U21335 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n19328), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19346), .ZN(n19304) );
  AOI22_X1 U21336 ( .A1(n19297), .A2(n19349), .B1(n19296), .B2(n19348), .ZN(
        n19303) );
  AOI21_X1 U21337 ( .B1(n19300), .B2(n19299), .A(n19298), .ZN(n19301) );
  NAND2_X1 U21338 ( .A1(n19316), .A2(n19301), .ZN(n19302) );
  NAND4_X1 U21339 ( .A1(n19305), .A2(n19304), .A3(n19303), .A4(n19302), .ZN(
        P2_U2829) );
  INV_X1 U21340 ( .A(n19306), .ZN(n19308) );
  AOI22_X1 U21341 ( .A1(n19308), .A2(n19323), .B1(P2_REIP_REG_28__SCAN_IN), 
        .B2(n19307), .ZN(n19322) );
  AOI22_X1 U21342 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19346), .B1(
        P2_EBX_REG_28__SCAN_IN), .B2(n19328), .ZN(n19321) );
  OAI22_X1 U21343 ( .A1(n19311), .A2(n19310), .B1(n19309), .B2(n19336), .ZN(
        n19312) );
  INV_X1 U21344 ( .A(n19312), .ZN(n19320) );
  OR2_X1 U21345 ( .A1(n19313), .A2(n11181), .ZN(n19317) );
  OAI21_X1 U21346 ( .B1(n11181), .B2(n19318), .A(n19313), .ZN(n19315) );
  OAI211_X1 U21347 ( .C1(n19318), .C2(n19317), .A(n19316), .B(n19315), .ZN(
        n19319) );
  NAND4_X1 U21348 ( .A1(n19322), .A2(n19321), .A3(n19320), .A4(n19319), .ZN(
        P2_U2827) );
  AOI22_X1 U21349 ( .A1(n19324), .A2(n19323), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19346), .ZN(n19325) );
  OAI21_X1 U21350 ( .B1(n19326), .B2(n19338), .A(n19325), .ZN(n19327) );
  AOI21_X1 U21351 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n19328), .A(n19327), .ZN(
        n19335) );
  AOI21_X1 U21352 ( .B1(n19330), .B2(n19329), .A(n19432), .ZN(n19333) );
  AOI22_X1 U21353 ( .A1(n19333), .A2(n19332), .B1(n19331), .B2(n19349), .ZN(
        n19334) );
  OAI211_X1 U21354 ( .C1(n19337), .C2(n19336), .A(n19335), .B(n19334), .ZN(
        P2_U2826) );
  NOR2_X1 U21355 ( .A1(n19339), .A2(n19338), .ZN(n19345) );
  INV_X1 U21356 ( .A(n19340), .ZN(n19343) );
  OAI22_X1 U21357 ( .A1(n19343), .A2(n19342), .B1(n12219), .B2(n19341), .ZN(
        n19344) );
  AOI211_X1 U21358 ( .C1(n19346), .C2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n19345), .B(n19344), .ZN(n19352) );
  AOI22_X1 U21359 ( .A1(n19350), .A2(n19349), .B1(n19348), .B2(n19347), .ZN(
        n19351) );
  OAI211_X1 U21360 ( .C1(n19354), .C2(n19353), .A(n19352), .B(n19351), .ZN(
        P2_U2824) );
  AOI21_X1 U21361 ( .B1(n19355), .B2(n20083), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n19356) );
  OAI22_X1 U21362 ( .A1(n19357), .A2(n19356), .B1(n19929), .B2(n19435), .ZN(
        n19359) );
  INV_X1 U21363 ( .A(n19358), .ZN(n19365) );
  MUX2_X1 U21364 ( .A(n19360), .B(n19359), .S(n19365), .Z(P2_U3601) );
  NAND3_X1 U21365 ( .A1(n19365), .A2(n19362), .A3(n19361), .ZN(n19363) );
  OAI21_X1 U21366 ( .B1(n19365), .B2(n19364), .A(n19363), .ZN(P2_U3595) );
  INV_X1 U21367 ( .A(n19366), .ZN(n19368) );
  AOI22_X1 U21368 ( .A1(n19408), .A2(n19368), .B1(n19367), .B2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19370) );
  NAND2_X1 U21369 ( .A1(n19398), .A2(n12300), .ZN(n19369) );
  OAI211_X1 U21370 ( .C1(n19388), .C2(n19371), .A(n19370), .B(n19369), .ZN(
        n19372) );
  AOI21_X1 U21371 ( .B1(n12397), .B2(n19378), .A(n19372), .ZN(n19374) );
  OAI211_X1 U21372 ( .C1(n19376), .C2(n19375), .A(n19374), .B(n19373), .ZN(
        P2_U3046) );
  AOI21_X1 U21373 ( .B1(n19379), .B2(n19378), .A(n19377), .ZN(n19394) );
  NOR2_X1 U21374 ( .A1(n19380), .A2(n11776), .ZN(n19382) );
  AOI211_X1 U21375 ( .C1(n19408), .C2(n19383), .A(n19382), .B(n19381), .ZN(
        n19392) );
  NAND2_X1 U21376 ( .A1(n19384), .A2(n19420), .ZN(n19387) );
  NAND2_X1 U21377 ( .A1(n19398), .A2(n19385), .ZN(n19386) );
  OAI211_X1 U21378 ( .C1(n19389), .C2(n19388), .A(n19387), .B(n19386), .ZN(
        n19390) );
  INV_X1 U21379 ( .A(n19390), .ZN(n19391) );
  OAI211_X1 U21380 ( .C1(n19394), .C2(n19393), .A(n19392), .B(n19391), .ZN(
        P2_U3034) );
  AOI22_X1 U21381 ( .A1(n19396), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19408), .B2(n19395), .ZN(n19406) );
  AOI222_X1 U21382 ( .A1(n19400), .A2(n19420), .B1(n19419), .B2(n19399), .C1(
        n19398), .C2(n19397), .ZN(n19405) );
  NAND2_X1 U21383 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19407), .ZN(n19404) );
  OAI211_X1 U21384 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n19402), .B(n19401), .ZN(n19403) );
  NAND4_X1 U21385 ( .A1(n19406), .A2(n19405), .A3(n19404), .A4(n19403), .ZN(
        P2_U3038) );
  AOI22_X1 U21386 ( .A1(n19409), .A2(n19408), .B1(P2_REIP_REG_3__SCAN_IN), 
        .B2(n19407), .ZN(n19415) );
  NAND2_X1 U21387 ( .A1(n19411), .A2(n19410), .ZN(n19413) );
  MUX2_X1 U21388 ( .A(n19413), .B(n19412), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n19414) );
  OAI211_X1 U21389 ( .C1(n19416), .C2(n12312), .A(n19415), .B(n19414), .ZN(
        n19417) );
  INV_X1 U21390 ( .A(n19417), .ZN(n19423) );
  AOI22_X1 U21391 ( .A1(n19421), .A2(n19420), .B1(n19419), .B2(n19418), .ZN(
        n19422) );
  NAND2_X1 U21392 ( .A1(n19423), .A2(n19422), .ZN(P2_U3043) );
  AND2_X1 U21393 ( .A1(n19443), .A2(n19424), .ZN(n19438) );
  INV_X1 U21394 ( .A(n19438), .ZN(n19431) );
  OAI21_X1 U21395 ( .B1(n19426), .B2(n19425), .A(n19448), .ZN(n19430) );
  NAND2_X1 U21396 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n22338), .ZN(n19427) );
  AOI21_X1 U21397 ( .B1(n19428), .B2(n19431), .A(n19427), .ZN(n19429) );
  AOI21_X1 U21398 ( .B1(n19431), .B2(n19430), .A(n19429), .ZN(n19433) );
  NAND2_X1 U21399 ( .A1(n19433), .A2(n19432), .ZN(P2_U3177) );
  AOI21_X1 U21400 ( .B1(n19436), .B2(n19435), .A(n19434), .ZN(n19437) );
  AOI21_X1 U21401 ( .B1(n19438), .B2(n22338), .A(n19437), .ZN(n19439) );
  AOI211_X1 U21402 ( .C1(n19441), .C2(n22338), .A(n19440), .B(n19439), .ZN(
        n19445) );
  OAI21_X1 U21403 ( .B1(n19443), .B2(n19442), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19444) );
  OAI211_X1 U21404 ( .C1(n19446), .C2(n19448), .A(n19445), .B(n19444), .ZN(
        P2_U3176) );
  INV_X1 U21405 ( .A(n19447), .ZN(n19450) );
  NOR2_X1 U21406 ( .A1(n19449), .A2(n19448), .ZN(n19452) );
  MUX2_X1 U21407 ( .A(P2_MORE_REG_SCAN_IN), .B(n19450), .S(n19452), .Z(
        P2_U3609) );
  OAI21_X1 U21408 ( .B1(n19452), .B2(n12618), .A(n19451), .ZN(P2_U2819) );
  INV_X1 U21409 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20828) );
  INV_X1 U21410 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19922) );
  AOI22_X1 U21411 ( .A1(n19811), .A2(n20828), .B1(n19922), .B2(U215), .ZN(U282) );
  OAI22_X1 U21412 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19811), .ZN(n19453) );
  INV_X1 U21413 ( .A(n19453), .ZN(U281) );
  OAI22_X1 U21414 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19811), .ZN(n19454) );
  INV_X1 U21415 ( .A(n19454), .ZN(U280) );
  OAI22_X1 U21416 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19811), .ZN(n19455) );
  INV_X1 U21417 ( .A(n19455), .ZN(U279) );
  OAI22_X1 U21418 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19811), .ZN(n19456) );
  INV_X1 U21419 ( .A(n19456), .ZN(U278) );
  OAI22_X1 U21420 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19811), .ZN(n19457) );
  INV_X1 U21421 ( .A(n19457), .ZN(U277) );
  OAI22_X1 U21422 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19811), .ZN(n19458) );
  INV_X1 U21423 ( .A(n19458), .ZN(U276) );
  OAI22_X1 U21424 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19811), .ZN(n19459) );
  INV_X1 U21425 ( .A(n19459), .ZN(U275) );
  OAI22_X1 U21426 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19811), .ZN(n19460) );
  INV_X1 U21427 ( .A(n19460), .ZN(U274) );
  OAI22_X1 U21428 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19811), .ZN(n19461) );
  INV_X1 U21429 ( .A(n19461), .ZN(U273) );
  OAI22_X1 U21430 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19811), .ZN(n19462) );
  INV_X1 U21431 ( .A(n19462), .ZN(U272) );
  OAI22_X1 U21432 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19811), .ZN(n19463) );
  INV_X1 U21433 ( .A(n19463), .ZN(U271) );
  OAI22_X1 U21434 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19476), .ZN(n19464) );
  INV_X1 U21435 ( .A(n19464), .ZN(U270) );
  OAI22_X1 U21436 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19811), .ZN(n19465) );
  INV_X1 U21437 ( .A(n19465), .ZN(U269) );
  OAI22_X1 U21438 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19476), .ZN(n19466) );
  INV_X1 U21439 ( .A(n19466), .ZN(U268) );
  OAI22_X1 U21440 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19811), .ZN(n19467) );
  INV_X1 U21441 ( .A(n19467), .ZN(U267) );
  OAI22_X1 U21442 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19476), .ZN(n19468) );
  INV_X1 U21443 ( .A(n19468), .ZN(U266) );
  OAI22_X1 U21444 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n19811), .ZN(n19469) );
  INV_X1 U21445 ( .A(n19469), .ZN(U265) );
  OAI22_X1 U21446 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n19476), .ZN(n19470) );
  INV_X1 U21447 ( .A(n19470), .ZN(U264) );
  OAI22_X1 U21448 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n19476), .ZN(n19471) );
  INV_X1 U21449 ( .A(n19471), .ZN(U263) );
  OAI22_X1 U21450 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n19476), .ZN(n19472) );
  INV_X1 U21451 ( .A(n19472), .ZN(U262) );
  OAI22_X1 U21452 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n19476), .ZN(n19473) );
  INV_X1 U21453 ( .A(n19473), .ZN(U261) );
  OAI22_X1 U21454 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n19476), .ZN(n19474) );
  INV_X1 U21455 ( .A(n19474), .ZN(U260) );
  OAI22_X1 U21456 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n19476), .ZN(n19475) );
  INV_X1 U21457 ( .A(n19475), .ZN(U259) );
  OAI22_X1 U21458 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19476), .ZN(n19477) );
  INV_X1 U21459 ( .A(n19477), .ZN(U258) );
  NOR2_X1 U21460 ( .A1(n19522), .A2(n19503), .ZN(n19552) );
  NAND2_X1 U21461 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19552), .ZN(
        n19803) );
  NAND2_X1 U21462 ( .A1(n19478), .A2(n21945), .ZN(n19817) );
  OR2_X1 U21463 ( .A1(n19817), .A2(n21524), .ZN(n19564) );
  NAND2_X1 U21464 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19486) );
  NOR2_X2 U21465 ( .A1(n19542), .A2(n19486), .ZN(n19833) );
  NOR2_X2 U21466 ( .A1(n19922), .A2(n19813), .ZN(n19557) );
  AND2_X1 U21467 ( .A1(n19555), .A2(n19552), .ZN(n19816) );
  INV_X1 U21468 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n21374) );
  NOR2_X2 U21469 ( .A1(n21374), .A2(n19686), .ZN(n19556) );
  AOI22_X1 U21470 ( .A1(n19833), .A2(n19557), .B1(n19816), .B2(n19556), .ZN(
        n19481) );
  NOR2_X1 U21471 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19486), .ZN(
        n19487) );
  INV_X1 U21472 ( .A(n19686), .ZN(n19815) );
  NAND2_X1 U21473 ( .A1(n19497), .A2(n19815), .ZN(n19509) );
  INV_X1 U21474 ( .A(n19509), .ZN(n19488) );
  AOI22_X1 U21475 ( .A1(n19814), .A2(n19487), .B1(n19552), .B2(n19488), .ZN(
        n19818) );
  NOR2_X1 U21476 ( .A1(n19530), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19491) );
  INV_X1 U21477 ( .A(n19491), .ZN(n19536) );
  NOR2_X2 U21478 ( .A1(n19486), .A2(n19536), .ZN(n19906) );
  INV_X1 U21479 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n19479) );
  NOR2_X2 U21480 ( .A1(n19479), .A2(n19813), .ZN(n19561) );
  AOI22_X1 U21481 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19818), .B1(
        n19906), .B2(n19561), .ZN(n19480) );
  OAI211_X1 U21482 ( .C1(n19803), .C2(n19564), .A(n19481), .B(n19480), .ZN(
        P3_U2995) );
  NAND2_X1 U21483 ( .A1(n19552), .A2(n19530), .ZN(n19913) );
  INV_X1 U21484 ( .A(n19906), .ZN(n19810) );
  NAND2_X1 U21485 ( .A1(n19810), .A2(n19913), .ZN(n19560) );
  INV_X1 U21486 ( .A(n19560), .ZN(n19482) );
  NOR2_X1 U21487 ( .A1(n20894), .A2(n19482), .ZN(n19821) );
  AOI22_X1 U21488 ( .A1(n19561), .A2(n19833), .B1(n19556), .B2(n19821), .ZN(
        n19485) );
  INV_X1 U21489 ( .A(n19913), .ZN(n19822) );
  INV_X1 U21490 ( .A(n19833), .ZN(n19826) );
  NOR2_X1 U21491 ( .A1(n19524), .A2(n19508), .ZN(n19499) );
  NAND2_X1 U21492 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19499), .ZN(
        n19732) );
  NAND2_X1 U21493 ( .A1(n19826), .A2(n19732), .ZN(n19493) );
  INV_X1 U21494 ( .A(n19493), .ZN(n19492) );
  OAI21_X1 U21495 ( .B1(n19492), .B2(n19526), .A(n19482), .ZN(n19483) );
  OAI211_X1 U21496 ( .C1(n19822), .C2(n21949), .A(n19815), .B(n19483), .ZN(
        n19823) );
  INV_X1 U21497 ( .A(n19732), .ZN(n19840) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19823), .B1(
        n19557), .B2(n19840), .ZN(n19484) );
  OAI211_X1 U21499 ( .C1(n19564), .C2(n19913), .A(n19485), .B(n19484), .ZN(
        P3_U2987) );
  NAND2_X1 U21500 ( .A1(n19530), .A2(n19499), .ZN(n19831) );
  INV_X1 U21501 ( .A(n19831), .ZN(n19845) );
  NAND2_X1 U21502 ( .A1(n19524), .A2(n19555), .ZN(n19549) );
  NOR2_X1 U21503 ( .A1(n19486), .A2(n19549), .ZN(n19827) );
  AOI22_X1 U21504 ( .A1(n19557), .A2(n19845), .B1(n19556), .B2(n19827), .ZN(
        n19490) );
  AOI22_X1 U21505 ( .A1(n19814), .A2(n19499), .B1(n19488), .B2(n19487), .ZN(
        n19828) );
  AOI22_X1 U21506 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19828), .B1(
        n19561), .B2(n19840), .ZN(n19489) );
  OAI211_X1 U21507 ( .C1(n19810), .C2(n19564), .A(n19490), .B(n19489), .ZN(
        P3_U2979) );
  NAND2_X1 U21508 ( .A1(n19510), .A2(n19491), .ZN(n19837) );
  INV_X1 U21509 ( .A(n19837), .ZN(n19850) );
  NOR2_X1 U21510 ( .A1(n20894), .A2(n19492), .ZN(n19832) );
  AOI22_X1 U21511 ( .A1(n19557), .A2(n19850), .B1(n19556), .B2(n19832), .ZN(
        n19496) );
  NOR2_X1 U21512 ( .A1(n19845), .A2(n19850), .ZN(n19504) );
  INV_X1 U21513 ( .A(n19504), .ZN(n19494) );
  AOI21_X1 U21514 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n19686), .ZN(n19559) );
  AOI22_X1 U21515 ( .A1(n19814), .A2(n19494), .B1(n19559), .B2(n19493), .ZN(
        n19834) );
  AOI22_X1 U21516 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19834), .B1(
        n19561), .B2(n19845), .ZN(n19495) );
  OAI211_X1 U21517 ( .C1(n19564), .C2(n19826), .A(n19496), .B(n19495), .ZN(
        P3_U2971) );
  NOR2_X1 U21518 ( .A1(n19526), .A2(n19508), .ZN(n19498) );
  OAI211_X1 U21519 ( .C1(n19498), .C2(n19499), .A(n19497), .B(n19815), .ZN(
        n19839) );
  INV_X1 U21520 ( .A(n19499), .ZN(n19500) );
  NOR2_X1 U21521 ( .A1(n20894), .A2(n19500), .ZN(n19838) );
  AOI22_X1 U21522 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19839), .B1(
        n19556), .B2(n19838), .ZN(n19502) );
  NOR2_X2 U21523 ( .A1(n19542), .A2(n19508), .ZN(n19856) );
  AOI22_X1 U21524 ( .A1(n19561), .A2(n19850), .B1(n19557), .B2(n19856), .ZN(
        n19501) );
  OAI211_X1 U21525 ( .C1(n19564), .C2(n19732), .A(n19502), .B(n19501), .ZN(
        P3_U2963) );
  NOR2_X1 U21526 ( .A1(n19503), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19518) );
  NAND2_X1 U21527 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19518), .ZN(
        n19854) );
  INV_X1 U21528 ( .A(n19854), .ZN(n19862) );
  NOR2_X1 U21529 ( .A1(n20894), .A2(n19504), .ZN(n19844) );
  AOI22_X1 U21530 ( .A1(n19557), .A2(n19862), .B1(n19556), .B2(n19844), .ZN(
        n19507) );
  INV_X1 U21531 ( .A(n19856), .ZN(n19843) );
  NAND2_X1 U21532 ( .A1(n19843), .A2(n19854), .ZN(n19514) );
  INV_X1 U21533 ( .A(n19514), .ZN(n19513) );
  OAI21_X1 U21534 ( .B1(n19513), .B2(n19526), .A(n19504), .ZN(n19505) );
  OAI211_X1 U21535 ( .C1(n19845), .C2(n21949), .A(n19815), .B(n19505), .ZN(
        n19846) );
  AOI22_X1 U21536 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19846), .B1(
        n19561), .B2(n19856), .ZN(n19506) );
  OAI211_X1 U21537 ( .C1(n19564), .C2(n19831), .A(n19507), .B(n19506), .ZN(
        P3_U2955) );
  NOR2_X1 U21538 ( .A1(n19508), .A2(n19549), .ZN(n19849) );
  AOI22_X1 U21539 ( .A1(n19561), .A2(n19862), .B1(n19556), .B2(n19849), .ZN(
        n19512) );
  NOR2_X1 U21540 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19509), .ZN(
        n19551) );
  AOI22_X1 U21541 ( .A1(n19814), .A2(n19518), .B1(n19510), .B2(n19551), .ZN(
        n19851) );
  NAND2_X1 U21542 ( .A1(n19530), .A2(n19518), .ZN(n19785) );
  INV_X1 U21543 ( .A(n19785), .ZN(n19868) );
  AOI22_X1 U21544 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19851), .B1(
        n19557), .B2(n19868), .ZN(n19511) );
  OAI211_X1 U21545 ( .C1(n19564), .C2(n19837), .A(n19512), .B(n19511), .ZN(
        P3_U2947) );
  NOR2_X1 U21546 ( .A1(n20894), .A2(n19513), .ZN(n19855) );
  AOI22_X1 U21547 ( .A1(n19561), .A2(n19868), .B1(n19556), .B2(n19855), .ZN(
        n19517) );
  NOR2_X2 U21548 ( .A1(n19531), .A2(n19536), .ZN(n19873) );
  NOR2_X1 U21549 ( .A1(n19868), .A2(n19873), .ZN(n19525) );
  INV_X1 U21550 ( .A(n19525), .ZN(n19515) );
  AOI22_X1 U21551 ( .A1(n19814), .A2(n19515), .B1(n19559), .B2(n19514), .ZN(
        n19857) );
  AOI22_X1 U21552 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19857), .B1(
        n19557), .B2(n19873), .ZN(n19516) );
  OAI211_X1 U21553 ( .C1(n19564), .C2(n19843), .A(n19517), .B(n19516), .ZN(
        P3_U2939) );
  INV_X1 U21554 ( .A(n19518), .ZN(n19519) );
  NOR2_X1 U21555 ( .A1(n20894), .A2(n19519), .ZN(n19861) );
  AOI22_X1 U21556 ( .A1(n19561), .A2(n19873), .B1(n19556), .B2(n19861), .ZN(
        n19521) );
  AOI21_X1 U21557 ( .B1(n19524), .B2(n19526), .A(n19686), .ZN(n19541) );
  OAI211_X1 U21558 ( .C1(n19862), .C2(n21949), .A(n19532), .B(n19541), .ZN(
        n19863) );
  NOR2_X2 U21559 ( .A1(n19542), .A2(n19531), .ZN(n19879) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19863), .B1(
        n19557), .B2(n19879), .ZN(n19520) );
  OAI211_X1 U21561 ( .C1(n19564), .C2(n19854), .A(n19521), .B(n19520), .ZN(
        P3_U2931) );
  NAND2_X1 U21562 ( .A1(n19523), .A2(n19522), .ZN(n19548) );
  NOR2_X1 U21563 ( .A1(n19524), .A2(n19548), .ZN(n19540) );
  NAND2_X1 U21564 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19540), .ZN(
        n19877) );
  INV_X1 U21565 ( .A(n19877), .ZN(n19886) );
  NOR2_X1 U21566 ( .A1(n20894), .A2(n19525), .ZN(n19867) );
  AOI22_X1 U21567 ( .A1(n19557), .A2(n19886), .B1(n19556), .B2(n19867), .ZN(
        n19529) );
  INV_X1 U21568 ( .A(n19879), .ZN(n19866) );
  NAND2_X1 U21569 ( .A1(n19866), .A2(n19877), .ZN(n19537) );
  INV_X1 U21570 ( .A(n19537), .ZN(n19535) );
  OAI21_X1 U21571 ( .B1(n19535), .B2(n19526), .A(n19525), .ZN(n19527) );
  OAI211_X1 U21572 ( .C1(n19868), .C2(n21949), .A(n19815), .B(n19527), .ZN(
        n19869) );
  AOI22_X1 U21573 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19869), .B1(
        n19561), .B2(n19879), .ZN(n19528) );
  OAI211_X1 U21574 ( .C1(n19564), .C2(n19785), .A(n19529), .B(n19528), .ZN(
        P3_U2923) );
  INV_X1 U21575 ( .A(n19873), .ZN(n19860) );
  NAND2_X1 U21576 ( .A1(n19530), .A2(n19540), .ZN(n19794) );
  INV_X1 U21577 ( .A(n19794), .ZN(n19890) );
  NOR2_X1 U21578 ( .A1(n19531), .A2(n19549), .ZN(n19872) );
  AOI22_X1 U21579 ( .A1(n19557), .A2(n19890), .B1(n19556), .B2(n19872), .ZN(
        n19534) );
  AOI22_X1 U21580 ( .A1(n19814), .A2(n19540), .B1(n19532), .B2(n19551), .ZN(
        n19874) );
  AOI22_X1 U21581 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19874), .B1(
        n19561), .B2(n19886), .ZN(n19533) );
  OAI211_X1 U21582 ( .C1(n19564), .C2(n19860), .A(n19534), .B(n19533), .ZN(
        P3_U2915) );
  NOR2_X1 U21583 ( .A1(n20894), .A2(n19535), .ZN(n19878) );
  AOI22_X1 U21584 ( .A1(n19561), .A2(n19890), .B1(n19556), .B2(n19878), .ZN(
        n19539) );
  NOR2_X2 U21585 ( .A1(n19536), .A2(n19548), .ZN(n19898) );
  INV_X1 U21586 ( .A(n19898), .ZN(n19883) );
  NAND2_X1 U21587 ( .A1(n19794), .A2(n19883), .ZN(n19545) );
  AOI22_X1 U21588 ( .A1(n19814), .A2(n19545), .B1(n19559), .B2(n19537), .ZN(
        n19880) );
  AOI22_X1 U21589 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19880), .B1(
        n19557), .B2(n19898), .ZN(n19538) );
  OAI211_X1 U21590 ( .C1(n19564), .C2(n19866), .A(n19539), .B(n19538), .ZN(
        P3_U2907) );
  AND2_X1 U21591 ( .A1(n19555), .A2(n19540), .ZN(n19884) );
  AOI22_X1 U21592 ( .A1(n19561), .A2(n19898), .B1(n19556), .B2(n19884), .ZN(
        n19544) );
  INV_X1 U21593 ( .A(n19548), .ZN(n19550) );
  OAI211_X1 U21594 ( .C1(n19886), .C2(n21949), .A(n19550), .B(n19541), .ZN(
        n19885) );
  NOR2_X2 U21595 ( .A1(n19542), .A2(n19548), .ZN(n19908) );
  AOI22_X1 U21596 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19885), .B1(
        n19557), .B2(n19908), .ZN(n19543) );
  OAI211_X1 U21597 ( .C1(n19564), .C2(n19877), .A(n19544), .B(n19543), .ZN(
        P3_U2899) );
  AND2_X1 U21598 ( .A1(n19555), .A2(n19545), .ZN(n19889) );
  AOI22_X1 U21599 ( .A1(n19561), .A2(n19908), .B1(n19556), .B2(n19889), .ZN(
        n19547) );
  INV_X1 U21600 ( .A(n19908), .ZN(n19894) );
  NAND2_X1 U21601 ( .A1(n19803), .A2(n19894), .ZN(n19558) );
  AOI22_X1 U21602 ( .A1(n19814), .A2(n19558), .B1(n19559), .B2(n19545), .ZN(
        n19891) );
  INV_X1 U21603 ( .A(n19803), .ZN(n19897) );
  AOI22_X1 U21604 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19891), .B1(
        n19897), .B2(n19557), .ZN(n19546) );
  OAI211_X1 U21605 ( .C1(n19564), .C2(n19794), .A(n19547), .B(n19546), .ZN(
        P3_U2891) );
  NOR2_X1 U21606 ( .A1(n19549), .A2(n19548), .ZN(n19895) );
  AOI22_X1 U21607 ( .A1(n19557), .A2(n19822), .B1(n19556), .B2(n19895), .ZN(
        n19554) );
  AOI22_X1 U21608 ( .A1(n19814), .A2(n19552), .B1(n19551), .B2(n19550), .ZN(
        n19899) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19899), .B1(
        n19561), .B2(n19897), .ZN(n19553) );
  OAI211_X1 U21610 ( .C1(n19564), .C2(n19883), .A(n19554), .B(n19553), .ZN(
        P3_U2883) );
  AND2_X1 U21611 ( .A1(n19555), .A2(n19558), .ZN(n19904) );
  AOI22_X1 U21612 ( .A1(n19906), .A2(n19557), .B1(n19556), .B2(n19904), .ZN(
        n19563) );
  AOI22_X1 U21613 ( .A1(n19814), .A2(n19560), .B1(n19559), .B2(n19558), .ZN(
        n19909) );
  AOI22_X1 U21614 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19909), .B1(
        n19561), .B2(n19822), .ZN(n19562) );
  OAI211_X1 U21615 ( .C1(n19564), .C2(n19894), .A(n19563), .B(n19562), .ZN(
        P3_U2875) );
  OAI22_X1 U21616 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19811), .ZN(n19565) );
  INV_X1 U21617 ( .A(n19565), .ZN(U257) );
  INV_X1 U21618 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n20116) );
  NOR2_X1 U21619 ( .A1(n20116), .A2(n19813), .ZN(n19599) );
  INV_X1 U21620 ( .A(n19599), .ZN(n19597) );
  NAND2_X1 U21621 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n19814), .ZN(n19603) );
  INV_X1 U21622 ( .A(n19603), .ZN(n19594) );
  INV_X1 U21623 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n21380) );
  NOR2_X2 U21624 ( .A1(n21380), .A2(n19686), .ZN(n19598) );
  AOI22_X1 U21625 ( .A1(n19906), .A2(n19594), .B1(n19816), .B2(n19598), .ZN(
        n19567) );
  NOR2_X2 U21626 ( .A1(n21405), .A2(n19817), .ZN(n19600) );
  AOI22_X1 U21627 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19818), .B1(
        n19897), .B2(n19600), .ZN(n19566) );
  OAI211_X1 U21628 ( .C1(n19826), .C2(n19597), .A(n19567), .B(n19566), .ZN(
        P3_U2994) );
  AOI22_X1 U21629 ( .A1(n19833), .A2(n19594), .B1(n19821), .B2(n19598), .ZN(
        n19569) );
  AOI22_X1 U21630 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19823), .B1(
        n19822), .B2(n19600), .ZN(n19568) );
  OAI211_X1 U21631 ( .C1(n19732), .C2(n19597), .A(n19569), .B(n19568), .ZN(
        P3_U2986) );
  AOI22_X1 U21632 ( .A1(n19845), .A2(n19599), .B1(n19827), .B2(n19598), .ZN(
        n19571) );
  AOI22_X1 U21633 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19828), .B1(
        n19906), .B2(n19600), .ZN(n19570) );
  OAI211_X1 U21634 ( .C1(n19732), .C2(n19603), .A(n19571), .B(n19570), .ZN(
        P3_U2978) );
  AOI22_X1 U21635 ( .A1(n19845), .A2(n19594), .B1(n19832), .B2(n19598), .ZN(
        n19573) );
  AOI22_X1 U21636 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19834), .B1(
        n19833), .B2(n19600), .ZN(n19572) );
  OAI211_X1 U21637 ( .C1(n19837), .C2(n19597), .A(n19573), .B(n19572), .ZN(
        P3_U2970) );
  AOI22_X1 U21638 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19839), .B1(
        n19838), .B2(n19598), .ZN(n19575) );
  AOI22_X1 U21639 ( .A1(n19840), .A2(n19600), .B1(n19850), .B2(n19594), .ZN(
        n19574) );
  OAI211_X1 U21640 ( .C1(n19843), .C2(n19597), .A(n19575), .B(n19574), .ZN(
        P3_U2962) );
  AOI22_X1 U21641 ( .A1(n19862), .A2(n19599), .B1(n19844), .B2(n19598), .ZN(
        n19577) );
  AOI22_X1 U21642 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19846), .B1(
        n19845), .B2(n19600), .ZN(n19576) );
  OAI211_X1 U21643 ( .C1(n19843), .C2(n19603), .A(n19577), .B(n19576), .ZN(
        P3_U2954) );
  AOI22_X1 U21644 ( .A1(n19868), .A2(n19599), .B1(n19849), .B2(n19598), .ZN(
        n19579) );
  AOI22_X1 U21645 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n19600), .ZN(n19578) );
  OAI211_X1 U21646 ( .C1(n19854), .C2(n19603), .A(n19579), .B(n19578), .ZN(
        P3_U2946) );
  AOI22_X1 U21647 ( .A1(n19868), .A2(n19594), .B1(n19855), .B2(n19598), .ZN(
        n19581) );
  AOI22_X1 U21648 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19857), .B1(
        n19856), .B2(n19600), .ZN(n19580) );
  OAI211_X1 U21649 ( .C1(n19860), .C2(n19597), .A(n19581), .B(n19580), .ZN(
        P3_U2938) );
  AOI22_X1 U21650 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19863), .B1(
        n19861), .B2(n19598), .ZN(n19583) );
  AOI22_X1 U21651 ( .A1(n19862), .A2(n19600), .B1(n19879), .B2(n19599), .ZN(
        n19582) );
  OAI211_X1 U21652 ( .C1(n19860), .C2(n19603), .A(n19583), .B(n19582), .ZN(
        P3_U2930) );
  AOI22_X1 U21653 ( .A1(n19886), .A2(n19599), .B1(n19867), .B2(n19598), .ZN(
        n19585) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19869), .B1(
        n19868), .B2(n19600), .ZN(n19584) );
  OAI211_X1 U21655 ( .C1(n19866), .C2(n19603), .A(n19585), .B(n19584), .ZN(
        P3_U2922) );
  AOI22_X1 U21656 ( .A1(n19890), .A2(n19599), .B1(n19872), .B2(n19598), .ZN(
        n19587) );
  AOI22_X1 U21657 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19874), .B1(
        n19873), .B2(n19600), .ZN(n19586) );
  OAI211_X1 U21658 ( .C1(n19877), .C2(n19603), .A(n19587), .B(n19586), .ZN(
        P3_U2914) );
  AOI22_X1 U21659 ( .A1(n19890), .A2(n19594), .B1(n19878), .B2(n19598), .ZN(
        n19589) );
  AOI22_X1 U21660 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19880), .B1(
        n19879), .B2(n19600), .ZN(n19588) );
  OAI211_X1 U21661 ( .C1(n19883), .C2(n19597), .A(n19589), .B(n19588), .ZN(
        P3_U2906) );
  AOI22_X1 U21662 ( .A1(n19898), .A2(n19594), .B1(n19884), .B2(n19598), .ZN(
        n19591) );
  AOI22_X1 U21663 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19885), .B1(
        n19886), .B2(n19600), .ZN(n19590) );
  OAI211_X1 U21664 ( .C1(n19894), .C2(n19597), .A(n19591), .B(n19590), .ZN(
        P3_U2898) );
  AOI22_X1 U21665 ( .A1(n19908), .A2(n19594), .B1(n19889), .B2(n19598), .ZN(
        n19593) );
  AOI22_X1 U21666 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19891), .B1(
        n19890), .B2(n19600), .ZN(n19592) );
  OAI211_X1 U21667 ( .C1(n19803), .C2(n19597), .A(n19593), .B(n19592), .ZN(
        P3_U2890) );
  AOI22_X1 U21668 ( .A1(n19897), .A2(n19594), .B1(n19895), .B2(n19598), .ZN(
        n19596) );
  AOI22_X1 U21669 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19899), .B1(
        n19898), .B2(n19600), .ZN(n19595) );
  OAI211_X1 U21670 ( .C1(n19913), .C2(n19597), .A(n19596), .B(n19595), .ZN(
        P3_U2882) );
  AOI22_X1 U21671 ( .A1(n19906), .A2(n19599), .B1(n19904), .B2(n19598), .ZN(
        n19602) );
  AOI22_X1 U21672 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19909), .B1(
        n19908), .B2(n19600), .ZN(n19601) );
  OAI211_X1 U21673 ( .C1(n19913), .C2(n19603), .A(n19602), .B(n19601), .ZN(
        P3_U2874) );
  OAI22_X1 U21674 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19811), .ZN(n19604) );
  INV_X1 U21675 ( .A(n19604), .ZN(U256) );
  INV_X1 U21676 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n21406) );
  NOR2_X1 U21677 ( .A1(n21406), .A2(n19813), .ZN(n19634) );
  INV_X1 U21678 ( .A(n19634), .ZN(n19643) );
  NAND2_X1 U21679 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19814), .ZN(n19637) );
  INV_X1 U21680 ( .A(n19637), .ZN(n19639) );
  INV_X1 U21681 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n21384) );
  NOR2_X2 U21682 ( .A1(n21384), .A2(n19686), .ZN(n19638) );
  AOI22_X1 U21683 ( .A1(n19833), .A2(n19639), .B1(n19816), .B2(n19638), .ZN(
        n19607) );
  NOR2_X2 U21684 ( .A1(n19605), .A2(n19817), .ZN(n19640) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19818), .B1(
        n19897), .B2(n19640), .ZN(n19606) );
  OAI211_X1 U21686 ( .C1(n19810), .C2(n19643), .A(n19607), .B(n19606), .ZN(
        P3_U2993) );
  AOI22_X1 U21687 ( .A1(n19833), .A2(n19634), .B1(n19821), .B2(n19638), .ZN(
        n19609) );
  AOI22_X1 U21688 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19823), .B1(
        n19822), .B2(n19640), .ZN(n19608) );
  OAI211_X1 U21689 ( .C1(n19732), .C2(n19637), .A(n19609), .B(n19608), .ZN(
        P3_U2985) );
  AOI22_X1 U21690 ( .A1(n19840), .A2(n19634), .B1(n19827), .B2(n19638), .ZN(
        n19611) );
  AOI22_X1 U21691 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19828), .B1(
        n19906), .B2(n19640), .ZN(n19610) );
  OAI211_X1 U21692 ( .C1(n19831), .C2(n19637), .A(n19611), .B(n19610), .ZN(
        P3_U2977) );
  AOI22_X1 U21693 ( .A1(n19845), .A2(n19634), .B1(n19832), .B2(n19638), .ZN(
        n19613) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19834), .B1(
        n19833), .B2(n19640), .ZN(n19612) );
  OAI211_X1 U21695 ( .C1(n19837), .C2(n19637), .A(n19613), .B(n19612), .ZN(
        P3_U2969) );
  AOI22_X1 U21696 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19839), .B1(
        n19838), .B2(n19638), .ZN(n19615) );
  AOI22_X1 U21697 ( .A1(n19840), .A2(n19640), .B1(n19850), .B2(n19634), .ZN(
        n19614) );
  OAI211_X1 U21698 ( .C1(n19843), .C2(n19637), .A(n19615), .B(n19614), .ZN(
        P3_U2961) );
  AOI22_X1 U21699 ( .A1(n19856), .A2(n19634), .B1(n19844), .B2(n19638), .ZN(
        n19617) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19846), .B1(
        n19845), .B2(n19640), .ZN(n19616) );
  OAI211_X1 U21701 ( .C1(n19854), .C2(n19637), .A(n19617), .B(n19616), .ZN(
        P3_U2953) );
  AOI22_X1 U21702 ( .A1(n19862), .A2(n19634), .B1(n19849), .B2(n19638), .ZN(
        n19619) );
  AOI22_X1 U21703 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n19640), .ZN(n19618) );
  OAI211_X1 U21704 ( .C1(n19785), .C2(n19637), .A(n19619), .B(n19618), .ZN(
        P3_U2945) );
  AOI22_X1 U21705 ( .A1(n19873), .A2(n19639), .B1(n19855), .B2(n19638), .ZN(
        n19621) );
  AOI22_X1 U21706 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19857), .B1(
        n19856), .B2(n19640), .ZN(n19620) );
  OAI211_X1 U21707 ( .C1(n19785), .C2(n19643), .A(n19621), .B(n19620), .ZN(
        P3_U2937) );
  AOI22_X1 U21708 ( .A1(n19879), .A2(n19639), .B1(n19861), .B2(n19638), .ZN(
        n19623) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19863), .B1(
        n19862), .B2(n19640), .ZN(n19622) );
  OAI211_X1 U21710 ( .C1(n19860), .C2(n19643), .A(n19623), .B(n19622), .ZN(
        P3_U2929) );
  AOI22_X1 U21711 ( .A1(n19886), .A2(n19639), .B1(n19867), .B2(n19638), .ZN(
        n19625) );
  AOI22_X1 U21712 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19869), .B1(
        n19868), .B2(n19640), .ZN(n19624) );
  OAI211_X1 U21713 ( .C1(n19866), .C2(n19643), .A(n19625), .B(n19624), .ZN(
        P3_U2921) );
  AOI22_X1 U21714 ( .A1(n19890), .A2(n19639), .B1(n19872), .B2(n19638), .ZN(
        n19627) );
  AOI22_X1 U21715 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19874), .B1(
        n19873), .B2(n19640), .ZN(n19626) );
  OAI211_X1 U21716 ( .C1(n19877), .C2(n19643), .A(n19627), .B(n19626), .ZN(
        P3_U2913) );
  AOI22_X1 U21717 ( .A1(n19898), .A2(n19639), .B1(n19878), .B2(n19638), .ZN(
        n19629) );
  AOI22_X1 U21718 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19880), .B1(
        n19879), .B2(n19640), .ZN(n19628) );
  OAI211_X1 U21719 ( .C1(n19794), .C2(n19643), .A(n19629), .B(n19628), .ZN(
        P3_U2905) );
  AOI22_X1 U21720 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19885), .B1(
        n19884), .B2(n19638), .ZN(n19631) );
  AOI22_X1 U21721 ( .A1(n19886), .A2(n19640), .B1(n19898), .B2(n19634), .ZN(
        n19630) );
  OAI211_X1 U21722 ( .C1(n19894), .C2(n19637), .A(n19631), .B(n19630), .ZN(
        P3_U2897) );
  AOI22_X1 U21723 ( .A1(n19908), .A2(n19634), .B1(n19889), .B2(n19638), .ZN(
        n19633) );
  AOI22_X1 U21724 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19891), .B1(
        n19890), .B2(n19640), .ZN(n19632) );
  OAI211_X1 U21725 ( .C1(n19803), .C2(n19637), .A(n19633), .B(n19632), .ZN(
        P3_U2889) );
  AOI22_X1 U21726 ( .A1(n19897), .A2(n19634), .B1(n19895), .B2(n19638), .ZN(
        n19636) );
  AOI22_X1 U21727 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19899), .B1(
        n19898), .B2(n19640), .ZN(n19635) );
  OAI211_X1 U21728 ( .C1(n19913), .C2(n19637), .A(n19636), .B(n19635), .ZN(
        P3_U2881) );
  AOI22_X1 U21729 ( .A1(n19906), .A2(n19639), .B1(n19904), .B2(n19638), .ZN(
        n19642) );
  AOI22_X1 U21730 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19909), .B1(
        n19908), .B2(n19640), .ZN(n19641) );
  OAI211_X1 U21731 ( .C1(n19913), .C2(n19643), .A(n19642), .B(n19641), .ZN(
        P3_U2873) );
  OAI22_X1 U21732 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19811), .ZN(n19644) );
  INV_X1 U21733 ( .A(n19644), .ZN(U255) );
  INV_X1 U21734 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n20222) );
  NOR2_X1 U21735 ( .A1(n20222), .A2(n19813), .ZN(n19672) );
  INV_X1 U21736 ( .A(n19672), .ZN(n19683) );
  NAND2_X1 U21737 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19814), .ZN(n19675) );
  INV_X1 U21738 ( .A(n19675), .ZN(n19679) );
  INV_X1 U21739 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n21390) );
  NOR2_X2 U21740 ( .A1(n21390), .A2(n19686), .ZN(n19678) );
  AOI22_X1 U21741 ( .A1(n19833), .A2(n19679), .B1(n19816), .B2(n19678), .ZN(
        n19647) );
  NOR2_X2 U21742 ( .A1(n19645), .A2(n19817), .ZN(n19680) );
  AOI22_X1 U21743 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19818), .B1(
        n19897), .B2(n19680), .ZN(n19646) );
  OAI211_X1 U21744 ( .C1(n19810), .C2(n19683), .A(n19647), .B(n19646), .ZN(
        P3_U2992) );
  AOI22_X1 U21745 ( .A1(n19840), .A2(n19679), .B1(n19821), .B2(n19678), .ZN(
        n19649) );
  AOI22_X1 U21746 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19823), .B1(
        n19822), .B2(n19680), .ZN(n19648) );
  OAI211_X1 U21747 ( .C1(n19826), .C2(n19683), .A(n19649), .B(n19648), .ZN(
        P3_U2984) );
  AOI22_X1 U21748 ( .A1(n19845), .A2(n19679), .B1(n19827), .B2(n19678), .ZN(
        n19651) );
  AOI22_X1 U21749 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19828), .B1(
        n19906), .B2(n19680), .ZN(n19650) );
  OAI211_X1 U21750 ( .C1(n19732), .C2(n19683), .A(n19651), .B(n19650), .ZN(
        P3_U2976) );
  AOI22_X1 U21751 ( .A1(n19850), .A2(n19679), .B1(n19832), .B2(n19678), .ZN(
        n19653) );
  AOI22_X1 U21752 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19834), .B1(
        n19833), .B2(n19680), .ZN(n19652) );
  OAI211_X1 U21753 ( .C1(n19831), .C2(n19683), .A(n19653), .B(n19652), .ZN(
        P3_U2968) );
  AOI22_X1 U21754 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19839), .B1(
        n19838), .B2(n19678), .ZN(n19655) );
  AOI22_X1 U21755 ( .A1(n19840), .A2(n19680), .B1(n19856), .B2(n19679), .ZN(
        n19654) );
  OAI211_X1 U21756 ( .C1(n19837), .C2(n19683), .A(n19655), .B(n19654), .ZN(
        P3_U2960) );
  AOI22_X1 U21757 ( .A1(n19862), .A2(n19679), .B1(n19844), .B2(n19678), .ZN(
        n19657) );
  AOI22_X1 U21758 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19846), .B1(
        n19845), .B2(n19680), .ZN(n19656) );
  OAI211_X1 U21759 ( .C1(n19843), .C2(n19683), .A(n19657), .B(n19656), .ZN(
        P3_U2952) );
  AOI22_X1 U21760 ( .A1(n19862), .A2(n19672), .B1(n19849), .B2(n19678), .ZN(
        n19659) );
  AOI22_X1 U21761 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n19680), .ZN(n19658) );
  OAI211_X1 U21762 ( .C1(n19785), .C2(n19675), .A(n19659), .B(n19658), .ZN(
        P3_U2944) );
  AOI22_X1 U21763 ( .A1(n19873), .A2(n19679), .B1(n19855), .B2(n19678), .ZN(
        n19661) );
  AOI22_X1 U21764 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19857), .B1(
        n19856), .B2(n19680), .ZN(n19660) );
  OAI211_X1 U21765 ( .C1(n19785), .C2(n19683), .A(n19661), .B(n19660), .ZN(
        P3_U2936) );
  AOI22_X1 U21766 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19863), .B1(
        n19861), .B2(n19678), .ZN(n19663) );
  AOI22_X1 U21767 ( .A1(n19862), .A2(n19680), .B1(n19879), .B2(n19679), .ZN(
        n19662) );
  OAI211_X1 U21768 ( .C1(n19860), .C2(n19683), .A(n19663), .B(n19662), .ZN(
        P3_U2928) );
  AOI22_X1 U21769 ( .A1(n19879), .A2(n19672), .B1(n19867), .B2(n19678), .ZN(
        n19665) );
  AOI22_X1 U21770 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19869), .B1(
        n19868), .B2(n19680), .ZN(n19664) );
  OAI211_X1 U21771 ( .C1(n19877), .C2(n19675), .A(n19665), .B(n19664), .ZN(
        P3_U2920) );
  AOI22_X1 U21772 ( .A1(n19886), .A2(n19672), .B1(n19872), .B2(n19678), .ZN(
        n19667) );
  AOI22_X1 U21773 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19874), .B1(
        n19873), .B2(n19680), .ZN(n19666) );
  OAI211_X1 U21774 ( .C1(n19794), .C2(n19675), .A(n19667), .B(n19666), .ZN(
        P3_U2912) );
  AOI22_X1 U21775 ( .A1(n19898), .A2(n19679), .B1(n19878), .B2(n19678), .ZN(
        n19669) );
  AOI22_X1 U21776 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19880), .B1(
        n19879), .B2(n19680), .ZN(n19668) );
  OAI211_X1 U21777 ( .C1(n19794), .C2(n19683), .A(n19669), .B(n19668), .ZN(
        P3_U2904) );
  AOI22_X1 U21778 ( .A1(n19898), .A2(n19672), .B1(n19884), .B2(n19678), .ZN(
        n19671) );
  AOI22_X1 U21779 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19885), .B1(
        n19886), .B2(n19680), .ZN(n19670) );
  OAI211_X1 U21780 ( .C1(n19894), .C2(n19675), .A(n19671), .B(n19670), .ZN(
        P3_U2896) );
  AOI22_X1 U21781 ( .A1(n19908), .A2(n19672), .B1(n19889), .B2(n19678), .ZN(
        n19674) );
  AOI22_X1 U21782 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19891), .B1(
        n19890), .B2(n19680), .ZN(n19673) );
  OAI211_X1 U21783 ( .C1(n19803), .C2(n19675), .A(n19674), .B(n19673), .ZN(
        P3_U2888) );
  AOI22_X1 U21784 ( .A1(n19822), .A2(n19679), .B1(n19895), .B2(n19678), .ZN(
        n19677) );
  AOI22_X1 U21785 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19899), .B1(
        n19898), .B2(n19680), .ZN(n19676) );
  OAI211_X1 U21786 ( .C1(n19803), .C2(n19683), .A(n19677), .B(n19676), .ZN(
        P3_U2880) );
  AOI22_X1 U21787 ( .A1(n19906), .A2(n19679), .B1(n19904), .B2(n19678), .ZN(
        n19682) );
  AOI22_X1 U21788 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19909), .B1(
        n19908), .B2(n19680), .ZN(n19681) );
  OAI211_X1 U21789 ( .C1(n19913), .C2(n19683), .A(n19682), .B(n19681), .ZN(
        P3_U2872) );
  OAI22_X1 U21790 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19811), .ZN(n19684) );
  INV_X1 U21791 ( .A(n19684), .ZN(U254) );
  INV_X1 U21792 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n19685) );
  NOR2_X1 U21793 ( .A1(n19685), .A2(n19813), .ZN(n19721) );
  INV_X1 U21794 ( .A(n19721), .ZN(n19717) );
  NAND2_X1 U21795 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19814), .ZN(n19725) );
  INV_X1 U21796 ( .A(n19725), .ZN(n19714) );
  INV_X1 U21797 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n21395) );
  NOR2_X2 U21798 ( .A1(n21395), .A2(n19686), .ZN(n19720) );
  AOI22_X1 U21799 ( .A1(n19833), .A2(n19714), .B1(n19816), .B2(n19720), .ZN(
        n19689) );
  NOR2_X2 U21800 ( .A1(n19687), .A2(n19817), .ZN(n19722) );
  AOI22_X1 U21801 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19818), .B1(
        n19897), .B2(n19722), .ZN(n19688) );
  OAI211_X1 U21802 ( .C1(n19810), .C2(n19717), .A(n19689), .B(n19688), .ZN(
        P3_U2991) );
  AOI22_X1 U21803 ( .A1(n19833), .A2(n19721), .B1(n19821), .B2(n19720), .ZN(
        n19691) );
  AOI22_X1 U21804 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19823), .B1(
        n19822), .B2(n19722), .ZN(n19690) );
  OAI211_X1 U21805 ( .C1(n19732), .C2(n19725), .A(n19691), .B(n19690), .ZN(
        P3_U2983) );
  AOI22_X1 U21806 ( .A1(n19845), .A2(n19714), .B1(n19827), .B2(n19720), .ZN(
        n19693) );
  AOI22_X1 U21807 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19828), .B1(
        n19906), .B2(n19722), .ZN(n19692) );
  OAI211_X1 U21808 ( .C1(n19732), .C2(n19717), .A(n19693), .B(n19692), .ZN(
        P3_U2975) );
  AOI22_X1 U21809 ( .A1(n19845), .A2(n19721), .B1(n19832), .B2(n19720), .ZN(
        n19695) );
  AOI22_X1 U21810 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19834), .B1(
        n19833), .B2(n19722), .ZN(n19694) );
  OAI211_X1 U21811 ( .C1(n19837), .C2(n19725), .A(n19695), .B(n19694), .ZN(
        P3_U2967) );
  AOI22_X1 U21812 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19839), .B1(
        n19838), .B2(n19720), .ZN(n19697) );
  AOI22_X1 U21813 ( .A1(n19840), .A2(n19722), .B1(n19850), .B2(n19721), .ZN(
        n19696) );
  OAI211_X1 U21814 ( .C1(n19843), .C2(n19725), .A(n19697), .B(n19696), .ZN(
        P3_U2959) );
  AOI22_X1 U21815 ( .A1(n19862), .A2(n19714), .B1(n19844), .B2(n19720), .ZN(
        n19699) );
  AOI22_X1 U21816 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19846), .B1(
        n19845), .B2(n19722), .ZN(n19698) );
  OAI211_X1 U21817 ( .C1(n19843), .C2(n19717), .A(n19699), .B(n19698), .ZN(
        P3_U2951) );
  AOI22_X1 U21818 ( .A1(n19862), .A2(n19721), .B1(n19849), .B2(n19720), .ZN(
        n19701) );
  AOI22_X1 U21819 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n19722), .ZN(n19700) );
  OAI211_X1 U21820 ( .C1(n19785), .C2(n19725), .A(n19701), .B(n19700), .ZN(
        P3_U2943) );
  AOI22_X1 U21821 ( .A1(n19868), .A2(n19721), .B1(n19855), .B2(n19720), .ZN(
        n19703) );
  AOI22_X1 U21822 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19857), .B1(
        n19856), .B2(n19722), .ZN(n19702) );
  OAI211_X1 U21823 ( .C1(n19860), .C2(n19725), .A(n19703), .B(n19702), .ZN(
        P3_U2935) );
  AOI22_X1 U21824 ( .A1(n19879), .A2(n19714), .B1(n19861), .B2(n19720), .ZN(
        n19705) );
  AOI22_X1 U21825 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19863), .B1(
        n19862), .B2(n19722), .ZN(n19704) );
  OAI211_X1 U21826 ( .C1(n19860), .C2(n19717), .A(n19705), .B(n19704), .ZN(
        P3_U2927) );
  AOI22_X1 U21827 ( .A1(n19879), .A2(n19721), .B1(n19867), .B2(n19720), .ZN(
        n19707) );
  AOI22_X1 U21828 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19869), .B1(
        n19868), .B2(n19722), .ZN(n19706) );
  OAI211_X1 U21829 ( .C1(n19877), .C2(n19725), .A(n19707), .B(n19706), .ZN(
        P3_U2919) );
  AOI22_X1 U21830 ( .A1(n19886), .A2(n19721), .B1(n19872), .B2(n19720), .ZN(
        n19709) );
  AOI22_X1 U21831 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19874), .B1(
        n19873), .B2(n19722), .ZN(n19708) );
  OAI211_X1 U21832 ( .C1(n19794), .C2(n19725), .A(n19709), .B(n19708), .ZN(
        P3_U2911) );
  AOI22_X1 U21833 ( .A1(n19898), .A2(n19714), .B1(n19878), .B2(n19720), .ZN(
        n19711) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19880), .B1(
        n19879), .B2(n19722), .ZN(n19710) );
  OAI211_X1 U21835 ( .C1(n19794), .C2(n19717), .A(n19711), .B(n19710), .ZN(
        P3_U2903) );
  AOI22_X1 U21836 ( .A1(n19908), .A2(n19714), .B1(n19884), .B2(n19720), .ZN(
        n19713) );
  AOI22_X1 U21837 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19885), .B1(
        n19886), .B2(n19722), .ZN(n19712) );
  OAI211_X1 U21838 ( .C1(n19883), .C2(n19717), .A(n19713), .B(n19712), .ZN(
        P3_U2895) );
  AOI22_X1 U21839 ( .A1(n19897), .A2(n19714), .B1(n19889), .B2(n19720), .ZN(
        n19716) );
  AOI22_X1 U21840 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19891), .B1(
        n19890), .B2(n19722), .ZN(n19715) );
  OAI211_X1 U21841 ( .C1(n19894), .C2(n19717), .A(n19716), .B(n19715), .ZN(
        P3_U2887) );
  AOI22_X1 U21842 ( .A1(n19897), .A2(n19721), .B1(n19895), .B2(n19720), .ZN(
        n19719) );
  AOI22_X1 U21843 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19899), .B1(
        n19898), .B2(n19722), .ZN(n19718) );
  OAI211_X1 U21844 ( .C1(n19913), .C2(n19725), .A(n19719), .B(n19718), .ZN(
        P3_U2879) );
  AOI22_X1 U21845 ( .A1(n19822), .A2(n19721), .B1(n19904), .B2(n19720), .ZN(
        n19724) );
  AOI22_X1 U21846 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19909), .B1(
        n19908), .B2(n19722), .ZN(n19723) );
  OAI211_X1 U21847 ( .C1(n19810), .C2(n19725), .A(n19724), .B(n19723), .ZN(
        P3_U2871) );
  OAI22_X1 U21848 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19811), .ZN(n19726) );
  INV_X1 U21849 ( .A(n19726), .ZN(U253) );
  INV_X1 U21850 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n20326) );
  NOR2_X1 U21851 ( .A1(n19813), .A2(n20326), .ZN(n19757) );
  INV_X1 U21852 ( .A(n19757), .ZN(n19766) );
  NAND2_X1 U21853 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19814), .ZN(n19760) );
  INV_X1 U21854 ( .A(n19760), .ZN(n19762) );
  AND2_X1 U21855 ( .A1(n19815), .A2(BUF2_REG_2__SCAN_IN), .ZN(n19761) );
  AOI22_X1 U21856 ( .A1(n19833), .A2(n19762), .B1(n19816), .B2(n19761), .ZN(
        n19729) );
  NOR2_X2 U21857 ( .A1(n19727), .A2(n19817), .ZN(n19763) );
  AOI22_X1 U21858 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19818), .B1(
        n19897), .B2(n19763), .ZN(n19728) );
  OAI211_X1 U21859 ( .C1(n19810), .C2(n19766), .A(n19729), .B(n19728), .ZN(
        P3_U2990) );
  AOI22_X1 U21860 ( .A1(n19833), .A2(n19757), .B1(n19821), .B2(n19761), .ZN(
        n19731) );
  AOI22_X1 U21861 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19823), .B1(
        n19822), .B2(n19763), .ZN(n19730) );
  OAI211_X1 U21862 ( .C1(n19732), .C2(n19760), .A(n19731), .B(n19730), .ZN(
        P3_U2982) );
  AOI22_X1 U21863 ( .A1(n19840), .A2(n19757), .B1(n19827), .B2(n19761), .ZN(
        n19734) );
  AOI22_X1 U21864 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19828), .B1(
        n19906), .B2(n19763), .ZN(n19733) );
  OAI211_X1 U21865 ( .C1(n19831), .C2(n19760), .A(n19734), .B(n19733), .ZN(
        P3_U2974) );
  AOI22_X1 U21866 ( .A1(n19850), .A2(n19762), .B1(n19832), .B2(n19761), .ZN(
        n19736) );
  AOI22_X1 U21867 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19834), .B1(
        n19833), .B2(n19763), .ZN(n19735) );
  OAI211_X1 U21868 ( .C1(n19831), .C2(n19766), .A(n19736), .B(n19735), .ZN(
        P3_U2966) );
  AOI22_X1 U21869 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19839), .B1(
        n19838), .B2(n19761), .ZN(n19738) );
  AOI22_X1 U21870 ( .A1(n19840), .A2(n19763), .B1(n19856), .B2(n19762), .ZN(
        n19737) );
  OAI211_X1 U21871 ( .C1(n19837), .C2(n19766), .A(n19738), .B(n19737), .ZN(
        P3_U2958) );
  AOI22_X1 U21872 ( .A1(n19856), .A2(n19757), .B1(n19844), .B2(n19761), .ZN(
        n19740) );
  AOI22_X1 U21873 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19846), .B1(
        n19845), .B2(n19763), .ZN(n19739) );
  OAI211_X1 U21874 ( .C1(n19854), .C2(n19760), .A(n19740), .B(n19739), .ZN(
        P3_U2950) );
  AOI22_X1 U21875 ( .A1(n19868), .A2(n19762), .B1(n19849), .B2(n19761), .ZN(
        n19742) );
  AOI22_X1 U21876 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n19763), .ZN(n19741) );
  OAI211_X1 U21877 ( .C1(n19854), .C2(n19766), .A(n19742), .B(n19741), .ZN(
        P3_U2942) );
  AOI22_X1 U21878 ( .A1(n19873), .A2(n19762), .B1(n19855), .B2(n19761), .ZN(
        n19744) );
  AOI22_X1 U21879 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19857), .B1(
        n19856), .B2(n19763), .ZN(n19743) );
  OAI211_X1 U21880 ( .C1(n19785), .C2(n19766), .A(n19744), .B(n19743), .ZN(
        P3_U2934) );
  AOI22_X1 U21881 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19863), .B1(
        n19861), .B2(n19761), .ZN(n19746) );
  AOI22_X1 U21882 ( .A1(n19862), .A2(n19763), .B1(n19879), .B2(n19762), .ZN(
        n19745) );
  OAI211_X1 U21883 ( .C1(n19860), .C2(n19766), .A(n19746), .B(n19745), .ZN(
        P3_U2926) );
  AOI22_X1 U21884 ( .A1(n19879), .A2(n19757), .B1(n19867), .B2(n19761), .ZN(
        n19748) );
  AOI22_X1 U21885 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19869), .B1(
        n19868), .B2(n19763), .ZN(n19747) );
  OAI211_X1 U21886 ( .C1(n19877), .C2(n19760), .A(n19748), .B(n19747), .ZN(
        P3_U2918) );
  AOI22_X1 U21887 ( .A1(n19890), .A2(n19762), .B1(n19872), .B2(n19761), .ZN(
        n19750) );
  AOI22_X1 U21888 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19874), .B1(
        n19873), .B2(n19763), .ZN(n19749) );
  OAI211_X1 U21889 ( .C1(n19877), .C2(n19766), .A(n19750), .B(n19749), .ZN(
        P3_U2910) );
  AOI22_X1 U21890 ( .A1(n19890), .A2(n19757), .B1(n19878), .B2(n19761), .ZN(
        n19752) );
  AOI22_X1 U21891 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19880), .B1(
        n19879), .B2(n19763), .ZN(n19751) );
  OAI211_X1 U21892 ( .C1(n19883), .C2(n19760), .A(n19752), .B(n19751), .ZN(
        P3_U2902) );
  AOI22_X1 U21893 ( .A1(n19898), .A2(n19757), .B1(n19884), .B2(n19761), .ZN(
        n19754) );
  AOI22_X1 U21894 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19885), .B1(
        n19886), .B2(n19763), .ZN(n19753) );
  OAI211_X1 U21895 ( .C1(n19894), .C2(n19760), .A(n19754), .B(n19753), .ZN(
        P3_U2894) );
  AOI22_X1 U21896 ( .A1(n19897), .A2(n19762), .B1(n19889), .B2(n19761), .ZN(
        n19756) );
  AOI22_X1 U21897 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19891), .B1(
        n19890), .B2(n19763), .ZN(n19755) );
  OAI211_X1 U21898 ( .C1(n19894), .C2(n19766), .A(n19756), .B(n19755), .ZN(
        P3_U2886) );
  AOI22_X1 U21899 ( .A1(n19897), .A2(n19757), .B1(n19895), .B2(n19761), .ZN(
        n19759) );
  AOI22_X1 U21900 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19899), .B1(
        n19898), .B2(n19763), .ZN(n19758) );
  OAI211_X1 U21901 ( .C1(n19913), .C2(n19760), .A(n19759), .B(n19758), .ZN(
        P3_U2878) );
  AOI22_X1 U21902 ( .A1(n19906), .A2(n19762), .B1(n19904), .B2(n19761), .ZN(
        n19765) );
  AOI22_X1 U21903 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19909), .B1(
        n19908), .B2(n19763), .ZN(n19764) );
  OAI211_X1 U21904 ( .C1(n19913), .C2(n19766), .A(n19765), .B(n19764), .ZN(
        P3_U2870) );
  OAI22_X1 U21905 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19811), .ZN(n19767) );
  INV_X1 U21906 ( .A(n19767), .ZN(U252) );
  INV_X1 U21907 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n19768) );
  NOR2_X1 U21908 ( .A1(n19813), .A2(n19768), .ZN(n19805) );
  INV_X1 U21909 ( .A(n19805), .ZN(n19802) );
  NAND2_X1 U21910 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19814), .ZN(n19809) );
  INV_X1 U21911 ( .A(n19809), .ZN(n19799) );
  AND2_X1 U21912 ( .A1(n19815), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19804) );
  AOI22_X1 U21913 ( .A1(n19833), .A2(n19799), .B1(n19816), .B2(n19804), .ZN(
        n19770) );
  NOR2_X2 U21914 ( .A1(n21337), .A2(n19817), .ZN(n19806) );
  AOI22_X1 U21915 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19818), .B1(
        n19897), .B2(n19806), .ZN(n19769) );
  OAI211_X1 U21916 ( .C1(n19810), .C2(n19802), .A(n19770), .B(n19769), .ZN(
        P3_U2989) );
  AOI22_X1 U21917 ( .A1(n19840), .A2(n19799), .B1(n19821), .B2(n19804), .ZN(
        n19772) );
  AOI22_X1 U21918 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19823), .B1(
        n19822), .B2(n19806), .ZN(n19771) );
  OAI211_X1 U21919 ( .C1(n19826), .C2(n19802), .A(n19772), .B(n19771), .ZN(
        P3_U2981) );
  AOI22_X1 U21920 ( .A1(n19840), .A2(n19805), .B1(n19827), .B2(n19804), .ZN(
        n19774) );
  AOI22_X1 U21921 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19828), .B1(
        n19906), .B2(n19806), .ZN(n19773) );
  OAI211_X1 U21922 ( .C1(n19831), .C2(n19809), .A(n19774), .B(n19773), .ZN(
        P3_U2973) );
  AOI22_X1 U21923 ( .A1(n19845), .A2(n19805), .B1(n19832), .B2(n19804), .ZN(
        n19776) );
  AOI22_X1 U21924 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19834), .B1(
        n19833), .B2(n19806), .ZN(n19775) );
  OAI211_X1 U21925 ( .C1(n19837), .C2(n19809), .A(n19776), .B(n19775), .ZN(
        P3_U2965) );
  AOI22_X1 U21926 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19839), .B1(
        n19838), .B2(n19804), .ZN(n19778) );
  AOI22_X1 U21927 ( .A1(n19840), .A2(n19806), .B1(n19850), .B2(n19805), .ZN(
        n19777) );
  OAI211_X1 U21928 ( .C1(n19843), .C2(n19809), .A(n19778), .B(n19777), .ZN(
        P3_U2957) );
  AOI22_X1 U21929 ( .A1(n19862), .A2(n19799), .B1(n19844), .B2(n19804), .ZN(
        n19780) );
  AOI22_X1 U21930 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19846), .B1(
        n19845), .B2(n19806), .ZN(n19779) );
  OAI211_X1 U21931 ( .C1(n19843), .C2(n19802), .A(n19780), .B(n19779), .ZN(
        P3_U2949) );
  AOI22_X1 U21932 ( .A1(n19862), .A2(n19805), .B1(n19849), .B2(n19804), .ZN(
        n19782) );
  AOI22_X1 U21933 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n19806), .ZN(n19781) );
  OAI211_X1 U21934 ( .C1(n19785), .C2(n19809), .A(n19782), .B(n19781), .ZN(
        P3_U2941) );
  AOI22_X1 U21935 ( .A1(n19873), .A2(n19799), .B1(n19855), .B2(n19804), .ZN(
        n19784) );
  AOI22_X1 U21936 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19857), .B1(
        n19856), .B2(n19806), .ZN(n19783) );
  OAI211_X1 U21937 ( .C1(n19785), .C2(n19802), .A(n19784), .B(n19783), .ZN(
        P3_U2933) );
  AOI22_X1 U21938 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19863), .B1(
        n19861), .B2(n19804), .ZN(n19787) );
  AOI22_X1 U21939 ( .A1(n19862), .A2(n19806), .B1(n19873), .B2(n19805), .ZN(
        n19786) );
  OAI211_X1 U21940 ( .C1(n19866), .C2(n19809), .A(n19787), .B(n19786), .ZN(
        P3_U2925) );
  AOI22_X1 U21941 ( .A1(n19886), .A2(n19799), .B1(n19867), .B2(n19804), .ZN(
        n19789) );
  AOI22_X1 U21942 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19869), .B1(
        n19868), .B2(n19806), .ZN(n19788) );
  OAI211_X1 U21943 ( .C1(n19866), .C2(n19802), .A(n19789), .B(n19788), .ZN(
        P3_U2917) );
  AOI22_X1 U21944 ( .A1(n19886), .A2(n19805), .B1(n19872), .B2(n19804), .ZN(
        n19791) );
  AOI22_X1 U21945 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19874), .B1(
        n19873), .B2(n19806), .ZN(n19790) );
  OAI211_X1 U21946 ( .C1(n19794), .C2(n19809), .A(n19791), .B(n19790), .ZN(
        P3_U2909) );
  AOI22_X1 U21947 ( .A1(n19898), .A2(n19799), .B1(n19878), .B2(n19804), .ZN(
        n19793) );
  AOI22_X1 U21948 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19880), .B1(
        n19879), .B2(n19806), .ZN(n19792) );
  OAI211_X1 U21949 ( .C1(n19794), .C2(n19802), .A(n19793), .B(n19792), .ZN(
        P3_U2901) );
  AOI22_X1 U21950 ( .A1(n19908), .A2(n19799), .B1(n19884), .B2(n19804), .ZN(
        n19796) );
  AOI22_X1 U21951 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19885), .B1(
        n19886), .B2(n19806), .ZN(n19795) );
  OAI211_X1 U21952 ( .C1(n19883), .C2(n19802), .A(n19796), .B(n19795), .ZN(
        P3_U2893) );
  AOI22_X1 U21953 ( .A1(n19908), .A2(n19805), .B1(n19889), .B2(n19804), .ZN(
        n19798) );
  AOI22_X1 U21954 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19891), .B1(
        n19890), .B2(n19806), .ZN(n19797) );
  OAI211_X1 U21955 ( .C1(n19803), .C2(n19809), .A(n19798), .B(n19797), .ZN(
        P3_U2885) );
  AOI22_X1 U21956 ( .A1(n19822), .A2(n19799), .B1(n19895), .B2(n19804), .ZN(
        n19801) );
  AOI22_X1 U21957 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19899), .B1(
        n19898), .B2(n19806), .ZN(n19800) );
  OAI211_X1 U21958 ( .C1(n19803), .C2(n19802), .A(n19801), .B(n19800), .ZN(
        P3_U2877) );
  AOI22_X1 U21959 ( .A1(n19822), .A2(n19805), .B1(n19904), .B2(n19804), .ZN(
        n19808) );
  AOI22_X1 U21960 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19909), .B1(
        n19908), .B2(n19806), .ZN(n19807) );
  OAI211_X1 U21961 ( .C1(n19810), .C2(n19809), .A(n19808), .B(n19807), .ZN(
        P3_U2869) );
  OAI22_X1 U21962 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19811), .ZN(n19812) );
  INV_X1 U21963 ( .A(n19812), .ZN(U251) );
  INV_X1 U21964 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n21484) );
  NOR2_X1 U21965 ( .A1(n21484), .A2(n19813), .ZN(n19905) );
  INV_X1 U21966 ( .A(n19905), .ZN(n19902) );
  NAND2_X1 U21967 ( .A1(n19814), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19912) );
  INV_X1 U21968 ( .A(n19912), .ZN(n19896) );
  AND2_X1 U21969 ( .A1(n19815), .A2(BUF2_REG_0__SCAN_IN), .ZN(n19903) );
  AOI22_X1 U21970 ( .A1(n19906), .A2(n19896), .B1(n19816), .B2(n19903), .ZN(
        n19820) );
  NOR2_X2 U21971 ( .A1(n21336), .A2(n19817), .ZN(n19907) );
  AOI22_X1 U21972 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19818), .B1(
        n19897), .B2(n19907), .ZN(n19819) );
  OAI211_X1 U21973 ( .C1(n19826), .C2(n19902), .A(n19820), .B(n19819), .ZN(
        P3_U2988) );
  AOI22_X1 U21974 ( .A1(n19840), .A2(n19905), .B1(n19821), .B2(n19903), .ZN(
        n19825) );
  AOI22_X1 U21975 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19823), .B1(
        n19822), .B2(n19907), .ZN(n19824) );
  OAI211_X1 U21976 ( .C1(n19826), .C2(n19912), .A(n19825), .B(n19824), .ZN(
        P3_U2980) );
  AOI22_X1 U21977 ( .A1(n19840), .A2(n19896), .B1(n19827), .B2(n19903), .ZN(
        n19830) );
  AOI22_X1 U21978 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19828), .B1(
        n19906), .B2(n19907), .ZN(n19829) );
  OAI211_X1 U21979 ( .C1(n19831), .C2(n19902), .A(n19830), .B(n19829), .ZN(
        P3_U2972) );
  AOI22_X1 U21980 ( .A1(n19845), .A2(n19896), .B1(n19832), .B2(n19903), .ZN(
        n19836) );
  AOI22_X1 U21981 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19834), .B1(
        n19833), .B2(n19907), .ZN(n19835) );
  OAI211_X1 U21982 ( .C1(n19837), .C2(n19902), .A(n19836), .B(n19835), .ZN(
        P3_U2964) );
  AOI22_X1 U21983 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19839), .B1(
        n19838), .B2(n19903), .ZN(n19842) );
  AOI22_X1 U21984 ( .A1(n19840), .A2(n19907), .B1(n19850), .B2(n19896), .ZN(
        n19841) );
  OAI211_X1 U21985 ( .C1(n19843), .C2(n19902), .A(n19842), .B(n19841), .ZN(
        P3_U2956) );
  AOI22_X1 U21986 ( .A1(n19856), .A2(n19896), .B1(n19844), .B2(n19903), .ZN(
        n19848) );
  AOI22_X1 U21987 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19846), .B1(
        n19845), .B2(n19907), .ZN(n19847) );
  OAI211_X1 U21988 ( .C1(n19854), .C2(n19902), .A(n19848), .B(n19847), .ZN(
        P3_U2948) );
  AOI22_X1 U21989 ( .A1(n19868), .A2(n19905), .B1(n19849), .B2(n19903), .ZN(
        n19853) );
  AOI22_X1 U21990 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19851), .B1(
        n19850), .B2(n19907), .ZN(n19852) );
  OAI211_X1 U21991 ( .C1(n19854), .C2(n19912), .A(n19853), .B(n19852), .ZN(
        P3_U2940) );
  AOI22_X1 U21992 ( .A1(n19868), .A2(n19896), .B1(n19855), .B2(n19903), .ZN(
        n19859) );
  AOI22_X1 U21993 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19857), .B1(
        n19856), .B2(n19907), .ZN(n19858) );
  OAI211_X1 U21994 ( .C1(n19860), .C2(n19902), .A(n19859), .B(n19858), .ZN(
        P3_U2932) );
  AOI22_X1 U21995 ( .A1(n19873), .A2(n19896), .B1(n19861), .B2(n19903), .ZN(
        n19865) );
  AOI22_X1 U21996 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19863), .B1(
        n19862), .B2(n19907), .ZN(n19864) );
  OAI211_X1 U21997 ( .C1(n19866), .C2(n19902), .A(n19865), .B(n19864), .ZN(
        P3_U2924) );
  AOI22_X1 U21998 ( .A1(n19879), .A2(n19896), .B1(n19867), .B2(n19903), .ZN(
        n19871) );
  AOI22_X1 U21999 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19869), .B1(
        n19868), .B2(n19907), .ZN(n19870) );
  OAI211_X1 U22000 ( .C1(n19877), .C2(n19902), .A(n19871), .B(n19870), .ZN(
        P3_U2916) );
  AOI22_X1 U22001 ( .A1(n19890), .A2(n19905), .B1(n19872), .B2(n19903), .ZN(
        n19876) );
  AOI22_X1 U22002 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19874), .B1(
        n19873), .B2(n19907), .ZN(n19875) );
  OAI211_X1 U22003 ( .C1(n19877), .C2(n19912), .A(n19876), .B(n19875), .ZN(
        P3_U2908) );
  AOI22_X1 U22004 ( .A1(n19890), .A2(n19896), .B1(n19878), .B2(n19903), .ZN(
        n19882) );
  AOI22_X1 U22005 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19880), .B1(
        n19879), .B2(n19907), .ZN(n19881) );
  OAI211_X1 U22006 ( .C1(n19883), .C2(n19902), .A(n19882), .B(n19881), .ZN(
        P3_U2900) );
  AOI22_X1 U22007 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19885), .B1(
        n19884), .B2(n19903), .ZN(n19888) );
  AOI22_X1 U22008 ( .A1(n19886), .A2(n19907), .B1(n19898), .B2(n19896), .ZN(
        n19887) );
  OAI211_X1 U22009 ( .C1(n19894), .C2(n19902), .A(n19888), .B(n19887), .ZN(
        P3_U2892) );
  AOI22_X1 U22010 ( .A1(n19897), .A2(n19905), .B1(n19889), .B2(n19903), .ZN(
        n19893) );
  AOI22_X1 U22011 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19891), .B1(
        n19890), .B2(n19907), .ZN(n19892) );
  OAI211_X1 U22012 ( .C1(n19894), .C2(n19912), .A(n19893), .B(n19892), .ZN(
        P3_U2884) );
  AOI22_X1 U22013 ( .A1(n19897), .A2(n19896), .B1(n19895), .B2(n19903), .ZN(
        n19901) );
  AOI22_X1 U22014 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19899), .B1(
        n19898), .B2(n19907), .ZN(n19900) );
  OAI211_X1 U22015 ( .C1(n19913), .C2(n19902), .A(n19901), .B(n19900), .ZN(
        P3_U2876) );
  AOI22_X1 U22016 ( .A1(n19906), .A2(n19905), .B1(n19904), .B2(n19903), .ZN(
        n19911) );
  AOI22_X1 U22017 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19909), .B1(
        n19908), .B2(n19907), .ZN(n19910) );
  OAI211_X1 U22018 ( .C1(n19913), .C2(n19912), .A(n19911), .B(n19910), .ZN(
        P3_U2868) );
  AOI22_X1 U22019 ( .A1(n19914), .A2(BUF2_REG_31__SCAN_IN), .B1(n20321), .B2(
        n19347), .ZN(n19917) );
  AOI22_X1 U22020 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n20319), .B1(n19915), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19916) );
  NAND2_X1 U22021 ( .A1(n19917), .A2(n19916), .ZN(P2_U2888) );
  AOI22_X1 U22022 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n11143), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n20424), .ZN(n20091) );
  NAND3_X1 U22023 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19930) );
  OAI21_X1 U22024 ( .B1(n19923), .B2(n20430), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19918) );
  OAI21_X1 U22025 ( .B1(n19930), .B2(n20096), .A(n19918), .ZN(n20431) );
  AND2_X1 U22026 ( .A1(n19921), .A2(n20428), .ZN(n20108) );
  AOI22_X1 U22027 ( .A1(n20431), .A2(n19920), .B1(n20430), .B2(n20108), .ZN(
        n19928) );
  NAND2_X1 U22028 ( .A1(n19944), .A2(n19929), .ZN(n20073) );
  INV_X1 U22029 ( .A(n20073), .ZN(n19964) );
  INV_X1 U22030 ( .A(n20439), .ZN(n20434) );
  INV_X1 U22031 ( .A(n19941), .ZN(n19945) );
  OAI21_X1 U22032 ( .B1(n19945), .B2(n20008), .A(n19930), .ZN(n19926) );
  AOI211_X1 U22033 ( .C1(n19923), .C2(n20101), .A(n20100), .B(n20430), .ZN(
        n19924) );
  NOR2_X1 U22034 ( .A1(n20426), .A2(n19924), .ZN(n19925) );
  NAND2_X1 U22035 ( .A1(n19926), .A2(n19925), .ZN(n20435) );
  AOI22_X1 U22036 ( .A1(n20109), .A2(n20434), .B1(
        P2_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n20435), .ZN(n19927) );
  OAI211_X1 U22037 ( .C1(n20091), .C2(n20540), .A(n19928), .B(n19927), .ZN(
        P2_U3175) );
  INV_X1 U22038 ( .A(n20108), .ZN(n20066) );
  NOR2_X1 U22039 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19930), .ZN(
        n20236) );
  INV_X1 U22040 ( .A(n20236), .ZN(n20438) );
  OAI22_X1 U22041 ( .A1(n20439), .A2(n20091), .B1(n20066), .B2(n20438), .ZN(
        n19931) );
  INV_X1 U22042 ( .A(n19931), .ZN(n19940) );
  NAND2_X1 U22043 ( .A1(n20445), .A2(n20439), .ZN(n19932) );
  AOI21_X1 U22044 ( .B1(n19932), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20096), 
        .ZN(n19935) );
  NAND3_X1 U22045 ( .A1(n20092), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19953) );
  NOR2_X1 U22046 ( .A1(n20094), .A2(n19953), .ZN(n20446) );
  INV_X1 U22047 ( .A(n20446), .ZN(n19946) );
  NAND2_X1 U22048 ( .A1(n19936), .A2(n20101), .ZN(n19933) );
  AOI22_X1 U22049 ( .A1(n19935), .A2(n19946), .B1(n19985), .B2(n19933), .ZN(
        n19934) );
  OAI21_X1 U22050 ( .B1(n20236), .B2(n20446), .A(n19935), .ZN(n19938) );
  OAI21_X1 U22051 ( .B1(n19936), .B2(n20236), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19937) );
  NAND2_X1 U22052 ( .A1(n19938), .A2(n19937), .ZN(n20441) );
  AOI22_X1 U22053 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20442), .B1(
        n19920), .B2(n20441), .ZN(n19939) );
  OAI211_X1 U22054 ( .C1(n20107), .C2(n20445), .A(n19940), .B(n19939), .ZN(
        P2_U3167) );
  OAI21_X1 U22055 ( .B1(n19942), .B2(n20446), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19943) );
  OAI21_X1 U22056 ( .B1(n19953), .B2(n20096), .A(n19943), .ZN(n20447) );
  AOI22_X1 U22057 ( .A1(n20447), .A2(n19920), .B1(n20108), .B2(n20446), .ZN(
        n19950) );
  OR2_X1 U22058 ( .A1(n19944), .A2(n22310), .ZN(n20029) );
  OAI21_X1 U22059 ( .B1(n19945), .B2(n20029), .A(n19953), .ZN(n19948) );
  OAI211_X1 U22060 ( .C1(n12371), .C2(n20032), .A(n19946), .B(n20096), .ZN(
        n19947) );
  NAND3_X1 U22061 ( .A1(n19948), .A2(n20086), .A3(n19947), .ZN(n20449) );
  INV_X1 U22062 ( .A(n20445), .ZN(n20448) );
  INV_X1 U22063 ( .A(n20091), .ZN(n20110) );
  AOI22_X1 U22064 ( .A1(n20449), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n20448), .B2(n20110), .ZN(n19949) );
  OAI211_X1 U22065 ( .C1(n20107), .C2(n20452), .A(n19950), .B(n19949), .ZN(
        P2_U3159) );
  NAND2_X1 U22066 ( .A1(n19951), .A2(n20017), .ZN(n20048) );
  NOR2_X1 U22067 ( .A1(n19952), .A2(n20048), .ZN(n19959) );
  INV_X1 U22068 ( .A(n19959), .ZN(n19956) );
  NOR2_X1 U22069 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19953), .ZN(
        n20453) );
  OAI21_X1 U22070 ( .B1(n19954), .B2(n20453), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19955) );
  OAI21_X1 U22071 ( .B1(n19956), .B2(n20096), .A(n19955), .ZN(n20454) );
  AOI22_X1 U22072 ( .A1(n20454), .A2(n19920), .B1(n20108), .B2(n20453), .ZN(
        n19962) );
  AOI21_X1 U22073 ( .B1(n20464), .B2(n20452), .A(n22310), .ZN(n19960) );
  INV_X1 U22074 ( .A(n20453), .ZN(n19957) );
  OAI211_X1 U22075 ( .C1(n12367), .C2(n20032), .A(n19957), .B(n20096), .ZN(
        n19958) );
  OAI211_X1 U22076 ( .C1(n19960), .C2(n19959), .A(n20086), .B(n19958), .ZN(
        n20456) );
  AOI22_X1 U22077 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20110), .ZN(n19961) );
  OAI211_X1 U22078 ( .C1(n20107), .C2(n20464), .A(n19962), .B(n19961), .ZN(
        P2_U3151) );
  NAND3_X1 U22079 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19998), .ZN(n19972) );
  NOR2_X1 U22080 ( .A1(n20094), .A2(n19972), .ZN(n20459) );
  OAI21_X1 U22081 ( .B1(n12358), .B2(n20459), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19963) );
  OAI21_X1 U22082 ( .B1(n19972), .B2(n20096), .A(n19963), .ZN(n20460) );
  AOI22_X1 U22083 ( .A1(n20460), .A2(n19920), .B1(n20108), .B2(n20459), .ZN(
        n19969) );
  AND2_X1 U22084 ( .A1(n12358), .A2(n20101), .ZN(n19967) );
  OR2_X1 U22085 ( .A1(n20100), .A2(n20459), .ZN(n19966) );
  OAI21_X1 U22086 ( .B1(n20058), .B2(n20057), .A(n19972), .ZN(n19965) );
  OAI211_X1 U22087 ( .C1(n19967), .C2(n19966), .A(n19965), .B(n20086), .ZN(
        n20461) );
  AOI22_X1 U22088 ( .A1(n20109), .A2(n20466), .B1(
        P2_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n20461), .ZN(n19968) );
  OAI211_X1 U22089 ( .C1(n20091), .C2(n20464), .A(n19969), .B(n19968), .ZN(
        P2_U3143) );
  INV_X1 U22090 ( .A(n20466), .ZN(n19970) );
  AOI21_X1 U22091 ( .B1(n19970), .B2(n20478), .A(n22310), .ZN(n19971) );
  NOR2_X1 U22092 ( .A1(n19971), .A2(n20096), .ZN(n19974) );
  NOR2_X1 U22093 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19972), .ZN(
        n20465) );
  NAND3_X1 U22094 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20092), .A3(
        n19998), .ZN(n19995) );
  NOR2_X1 U22095 ( .A1(n20094), .A2(n19995), .ZN(n20344) );
  NOR2_X1 U22096 ( .A1(n20465), .A2(n20344), .ZN(n19977) );
  AOI211_X1 U22097 ( .C1(n19975), .C2(n20083), .A(n20465), .B(n20100), .ZN(
        n19973) );
  INV_X1 U22098 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n19981) );
  AOI22_X1 U22099 ( .A1(n20466), .A2(n20110), .B1(n20108), .B2(n20465), .ZN(
        n19980) );
  INV_X1 U22100 ( .A(n19974), .ZN(n19978) );
  OAI21_X1 U22101 ( .B1(n19975), .B2(n20465), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19976) );
  AOI22_X1 U22102 ( .A1(n19920), .A2(n20468), .B1(n20467), .B2(n20109), .ZN(
        n19979) );
  OAI211_X1 U22103 ( .C1(n20471), .C2(n19981), .A(n19980), .B(n19979), .ZN(
        P2_U3135) );
  INV_X1 U22104 ( .A(n20344), .ZN(n20472) );
  OAI22_X1 U22105 ( .A1(n20478), .A2(n20091), .B1(n20472), .B2(n20066), .ZN(
        n19983) );
  INV_X1 U22106 ( .A(n19983), .ZN(n19994) );
  OAI21_X1 U22107 ( .B1(n19984), .B2(n20029), .A(n20100), .ZN(n19992) );
  INV_X1 U22108 ( .A(n19995), .ZN(n19989) );
  INV_X1 U22109 ( .A(n19985), .ZN(n19988) );
  NOR2_X1 U22110 ( .A1(n20344), .A2(n19990), .ZN(n19986) );
  AOI211_X1 U22111 ( .C1(n20032), .C2(n20472), .A(n20426), .B(n19986), .ZN(
        n19987) );
  OAI22_X1 U22112 ( .A1(n19992), .A2(n19989), .B1(n19988), .B2(n19987), .ZN(
        n20475) );
  OAI21_X1 U22113 ( .B1(n19990), .B2(n20344), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19991) );
  OAI21_X1 U22114 ( .B1(n19992), .B2(n19995), .A(n19991), .ZN(n20474) );
  AOI22_X1 U22115 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20475), .B1(
        n19920), .B2(n20474), .ZN(n19993) );
  OAI211_X1 U22116 ( .C1(n20107), .C2(n20480), .A(n19994), .B(n19993), .ZN(
        P2_U3127) );
  NOR2_X1 U22117 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19995), .ZN(
        n20347) );
  INV_X1 U22118 ( .A(n20347), .ZN(n20479) );
  OAI22_X1 U22119 ( .A1(n20480), .A2(n20091), .B1(n20066), .B2(n20479), .ZN(
        n19996) );
  INV_X1 U22120 ( .A(n19996), .ZN(n20006) );
  NAND2_X1 U22121 ( .A1(n20480), .A2(n20492), .ZN(n19997) );
  AOI21_X1 U22122 ( .B1(n19997), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20096), 
        .ZN(n20002) );
  NOR2_X1 U22123 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19998), .ZN(
        n20044) );
  NAND2_X1 U22124 ( .A1(n20061), .A2(n20044), .ZN(n20009) );
  OAI21_X1 U22125 ( .B1(n12317), .B2(n19999), .A(n20083), .ZN(n20000) );
  AOI21_X1 U22126 ( .B1(n20002), .B2(n20009), .A(n20000), .ZN(n20001) );
  INV_X1 U22127 ( .A(n20009), .ZN(n20486) );
  OAI21_X1 U22128 ( .B1(n20486), .B2(n20347), .A(n20002), .ZN(n20004) );
  OAI21_X1 U22129 ( .B1(n12317), .B2(n20347), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20003) );
  NAND2_X1 U22130 ( .A1(n20004), .A2(n20003), .ZN(n20482) );
  AOI22_X1 U22131 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20483), .B1(
        n20482), .B2(n19920), .ZN(n20005) );
  OAI211_X1 U22132 ( .C1(n20107), .C2(n20492), .A(n20006), .B(n20005), .ZN(
        P2_U3119) );
  NAND2_X1 U22133 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20044), .ZN(
        n20018) );
  OAI21_X1 U22134 ( .B1(n12365), .B2(n20486), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20007) );
  OAI21_X1 U22135 ( .B1(n20018), .B2(n20096), .A(n20007), .ZN(n20487) );
  AOI22_X1 U22136 ( .A1(n20487), .A2(n19920), .B1(n20486), .B2(n20108), .ZN(
        n20014) );
  OAI21_X1 U22137 ( .B1(n20030), .B2(n20008), .A(n20018), .ZN(n20012) );
  INV_X1 U22138 ( .A(n12365), .ZN(n20010) );
  OAI211_X1 U22139 ( .C1(n20010), .C2(n20032), .A(n20096), .B(n20009), .ZN(
        n20011) );
  NAND3_X1 U22140 ( .A1(n20012), .A2(n20086), .A3(n20011), .ZN(n20489) );
  AOI22_X1 U22141 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20489), .B1(
        n20495), .B2(n20109), .ZN(n20013) );
  OAI211_X1 U22142 ( .C1(n20091), .C2(n20492), .A(n20014), .B(n20013), .ZN(
        P2_U3111) );
  INV_X1 U22143 ( .A(n20044), .ZN(n20016) );
  OR2_X1 U22144 ( .A1(n20017), .A2(n20016), .ZN(n20022) );
  NOR2_X1 U22145 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20018), .ZN(
        n20493) );
  OAI21_X1 U22146 ( .B1(n12364), .B2(n20493), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20019) );
  OAI21_X1 U22147 ( .B1(n20096), .B2(n20022), .A(n20019), .ZN(n20494) );
  AOI22_X1 U22148 ( .A1(n20494), .A2(n19920), .B1(n20108), .B2(n20493), .ZN(
        n20026) );
  INV_X1 U22149 ( .A(n20493), .ZN(n20020) );
  OAI211_X1 U22150 ( .C1(n20021), .C2(n20032), .A(n20096), .B(n20020), .ZN(
        n20024) );
  OAI221_X1 U22151 ( .B1(n22310), .B2(n20402), .C1(n22310), .C2(n20505), .A(
        n20022), .ZN(n20023) );
  NAND3_X1 U22152 ( .A1(n20024), .A2(n20023), .A3(n20086), .ZN(n20496) );
  AOI22_X1 U22153 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20496), .B1(
        n20495), .B2(n20110), .ZN(n20025) );
  OAI211_X1 U22154 ( .C1(n20107), .C2(n20505), .A(n20026), .B(n20025), .ZN(
        P2_U3103) );
  NAND2_X1 U22155 ( .A1(n20044), .A2(n20092), .ZN(n20038) );
  NOR2_X1 U22156 ( .A1(n20094), .A2(n20038), .ZN(n20403) );
  AOI22_X1 U22157 ( .A1(n20109), .A2(n20359), .B1(n20108), .B2(n20403), .ZN(
        n20041) );
  OAI21_X1 U22158 ( .B1(n20030), .B2(n20029), .A(n20100), .ZN(n20039) );
  INV_X1 U22159 ( .A(n20038), .ZN(n20035) );
  OAI21_X1 U22160 ( .B1(n20100), .B2(n20403), .A(n20086), .ZN(n20031) );
  OAI21_X1 U22161 ( .B1(n20033), .B2(n20032), .A(n20031), .ZN(n20034) );
  OAI21_X1 U22162 ( .B1(n20039), .B2(n20035), .A(n20034), .ZN(n20502) );
  OAI21_X1 U22163 ( .B1(n20036), .B2(n20403), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20037) );
  OAI21_X1 U22164 ( .B1(n20039), .B2(n20038), .A(n20037), .ZN(n20501) );
  AOI22_X1 U22165 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20502), .B1(
        n19920), .B2(n20501), .ZN(n20040) );
  OAI211_X1 U22166 ( .C1(n20091), .C2(n20505), .A(n20041), .B(n20040), .ZN(
        P2_U3095) );
  INV_X1 U22167 ( .A(n20074), .ZN(n20043) );
  NAND2_X1 U22168 ( .A1(n20045), .A2(n20044), .ZN(n20506) );
  OAI22_X1 U22169 ( .A1(n20507), .A2(n20091), .B1(n20066), .B2(n20506), .ZN(
        n20046) );
  INV_X1 U22170 ( .A(n20046), .ZN(n20056) );
  OAI21_X1 U22171 ( .B1(n20362), .B2(n20359), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20047) );
  NAND2_X1 U22172 ( .A1(n20047), .A2(n20100), .ZN(n20054) );
  NOR2_X1 U22173 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20048), .ZN(
        n20051) );
  NAND2_X1 U22174 ( .A1(n12366), .A2(n20101), .ZN(n20049) );
  NAND3_X1 U22175 ( .A1(n20049), .A2(n20506), .A3(n20096), .ZN(n20050) );
  OAI211_X1 U22176 ( .C1(n20054), .C2(n20051), .A(n20086), .B(n20050), .ZN(
        n20510) );
  INV_X1 U22177 ( .A(n20051), .ZN(n20053) );
  INV_X1 U22178 ( .A(n20506), .ZN(n20358) );
  OAI21_X1 U22179 ( .B1(n12366), .B2(n20358), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20052) );
  AOI22_X1 U22180 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20510), .B1(
        n19920), .B2(n20509), .ZN(n20055) );
  OAI211_X1 U22181 ( .C1(n20107), .C2(n20515), .A(n20056), .B(n20055), .ZN(
        P2_U3087) );
  INV_X1 U22182 ( .A(n20057), .ZN(n20059) );
  NAND2_X1 U22183 ( .A1(n20059), .A2(n20058), .ZN(n20060) );
  NAND2_X1 U22184 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20093), .ZN(
        n20068) );
  NAND2_X1 U22185 ( .A1(n20060), .A2(n20068), .ZN(n20065) );
  NAND2_X1 U22186 ( .A1(n20070), .A2(n20101), .ZN(n20063) );
  AND2_X1 U22187 ( .A1(n20061), .A2(n20093), .ZN(n20411) );
  OAI21_X1 U22188 ( .B1(n20100), .B2(n20411), .A(n20086), .ZN(n20062) );
  NAND2_X1 U22189 ( .A1(n20063), .A2(n20062), .ZN(n20064) );
  AND2_X1 U22190 ( .A1(n20065), .A2(n20064), .ZN(n20206) );
  INV_X1 U22191 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n20077) );
  INV_X1 U22192 ( .A(n20411), .ZN(n20513) );
  OAI22_X1 U22193 ( .A1(n20515), .A2(n20091), .B1(n20513), .B2(n20066), .ZN(
        n20067) );
  INV_X1 U22194 ( .A(n20067), .ZN(n20076) );
  INV_X1 U22195 ( .A(n20068), .ZN(n20069) );
  NAND2_X1 U22196 ( .A1(n20069), .A2(n20100), .ZN(n20072) );
  OAI21_X1 U22197 ( .B1(n20070), .B2(n20411), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20071) );
  NAND2_X1 U22198 ( .A1(n20072), .A2(n20071), .ZN(n20517) );
  AOI22_X1 U22199 ( .A1(n19920), .A2(n20517), .B1(n20524), .B2(n20109), .ZN(
        n20075) );
  OAI211_X1 U22200 ( .C1(n20206), .C2(n20077), .A(n20076), .B(n20075), .ZN(
        P2_U3079) );
  NOR3_X2 U22201 ( .A1(n20092), .A2(n20078), .A3(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20522) );
  OAI21_X1 U22202 ( .B1(n12355), .B2(n20522), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20080) );
  OR2_X1 U22203 ( .A1(n20079), .A2(n20078), .ZN(n20084) );
  NAND2_X1 U22204 ( .A1(n20080), .A2(n20084), .ZN(n20523) );
  AOI22_X1 U22205 ( .A1(n20523), .A2(n19920), .B1(n20108), .B2(n20522), .ZN(
        n20090) );
  AOI21_X1 U22206 ( .B1(n20521), .B2(n20528), .A(n20082), .ZN(n20088) );
  AOI21_X1 U22207 ( .B1(n12355), .B2(n20083), .A(n20522), .ZN(n20085) );
  OAI21_X1 U22208 ( .B1(n20085), .B2(n20100), .A(n20084), .ZN(n20087) );
  OAI21_X1 U22209 ( .B1(n20088), .B2(n20087), .A(n20086), .ZN(n20525) );
  AOI22_X1 U22210 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20525), .B1(
        n20532), .B2(n20109), .ZN(n20089) );
  OAI211_X1 U22211 ( .C1(n20091), .C2(n20521), .A(n20090), .B(n20089), .ZN(
        P2_U3071) );
  NAND2_X1 U22212 ( .A1(n20093), .A2(n20092), .ZN(n20098) );
  NOR2_X1 U22213 ( .A1(n20094), .A2(n20098), .ZN(n20529) );
  OAI21_X1 U22214 ( .B1(n12357), .B2(n20529), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20095) );
  OAI21_X1 U22215 ( .B1(n20098), .B2(n20096), .A(n20095), .ZN(n20531) );
  AOI22_X1 U22216 ( .A1(n20531), .A2(n19920), .B1(n20108), .B2(n20529), .ZN(
        n20106) );
  INV_X1 U22217 ( .A(n20097), .ZN(n20099) );
  OAI21_X1 U22218 ( .B1(n20099), .B2(n22310), .A(n20098), .ZN(n20104) );
  AOI211_X1 U22219 ( .C1(n12357), .C2(n20101), .A(n20100), .B(n20529), .ZN(
        n20102) );
  NOR2_X1 U22220 ( .A1(n20426), .A2(n20102), .ZN(n20103) );
  NAND2_X1 U22221 ( .A1(n20104), .A2(n20103), .ZN(n20533) );
  AOI22_X1 U22222 ( .A1(n20533), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n20532), .B2(n20110), .ZN(n20105) );
  OAI211_X1 U22223 ( .C1(n20107), .C2(n20536), .A(n20106), .B(n20105), .ZN(
        P2_U3063) );
  AOI22_X1 U22224 ( .A1(n20109), .A2(n20274), .B1(n20268), .B2(n20108), .ZN(
        n20112) );
  AOI22_X1 U22225 ( .A1(n19920), .A2(n20543), .B1(n20545), .B2(n20110), .ZN(
        n20111) );
  OAI211_X1 U22226 ( .C1(n20548), .C2(n20113), .A(n20112), .B(n20111), .ZN(
        P2_U3055) );
  AOI22_X1 U22227 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n11143), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n20424), .ZN(n20145) );
  NAND2_X1 U22228 ( .A1(n11649), .A2(n20428), .ZN(n20156) );
  AOI22_X1 U22229 ( .A1(n20431), .A2(n20115), .B1(n20430), .B2(n20153), .ZN(
        n20118) );
  OAI22_X1 U22230 ( .A1(n20827), .A2(n20433), .B1(n20116), .B2(n20432), .ZN(
        n20147) );
  AOI22_X1 U22231 ( .A1(n20435), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n20434), .B2(n20147), .ZN(n20117) );
  OAI211_X1 U22232 ( .C1(n20145), .C2(n20540), .A(n20118), .B(n20117), .ZN(
        P2_U3174) );
  OAI22_X1 U22233 ( .A1(n20439), .A2(n20145), .B1(n20156), .B2(n20438), .ZN(
        n20119) );
  INV_X1 U22234 ( .A(n20119), .ZN(n20121) );
  AOI22_X1 U22235 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20442), .B1(
        n20115), .B2(n20441), .ZN(n20120) );
  OAI211_X1 U22236 ( .C1(n20157), .C2(n20445), .A(n20121), .B(n20120), .ZN(
        P2_U3166) );
  AOI22_X1 U22237 ( .A1(n20447), .A2(n20115), .B1(n20153), .B2(n20446), .ZN(
        n20123) );
  AOI22_X1 U22238 ( .A1(n20449), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n20147), .B2(n20455), .ZN(n20122) );
  OAI211_X1 U22239 ( .C1(n20145), .C2(n20445), .A(n20123), .B(n20122), .ZN(
        P2_U3158) );
  AOI22_X1 U22240 ( .A1(n20454), .A2(n20115), .B1(n20153), .B2(n20453), .ZN(
        n20125) );
  INV_X1 U22241 ( .A(n20145), .ZN(n20159) );
  AOI22_X1 U22242 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20159), .ZN(n20124) );
  OAI211_X1 U22243 ( .C1(n20157), .C2(n20464), .A(n20125), .B(n20124), .ZN(
        P2_U3150) );
  AOI22_X1 U22244 ( .A1(n20460), .A2(n20115), .B1(n20153), .B2(n20459), .ZN(
        n20127) );
  AOI22_X1 U22245 ( .A1(n20466), .A2(n20147), .B1(n20461), .B2(
        P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n20126) );
  OAI211_X1 U22246 ( .C1(n20145), .C2(n20464), .A(n20127), .B(n20126), .ZN(
        P2_U3142) );
  AOI22_X1 U22247 ( .A1(n20466), .A2(n20159), .B1(n20153), .B2(n20465), .ZN(
        n20129) );
  AOI22_X1 U22248 ( .A1(n20115), .A2(n20468), .B1(n20467), .B2(n20147), .ZN(
        n20128) );
  OAI211_X1 U22249 ( .C1(n20471), .C2(n16626), .A(n20129), .B(n20128), .ZN(
        P2_U3134) );
  OAI22_X1 U22250 ( .A1(n20480), .A2(n20157), .B1(n20472), .B2(n20156), .ZN(
        n20130) );
  INV_X1 U22251 ( .A(n20130), .ZN(n20132) );
  AOI22_X1 U22252 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20475), .B1(
        n20115), .B2(n20474), .ZN(n20131) );
  OAI211_X1 U22253 ( .C1(n20145), .C2(n20478), .A(n20132), .B(n20131), .ZN(
        P2_U3126) );
  OAI22_X1 U22254 ( .A1(n20480), .A2(n20145), .B1(n20156), .B2(n20479), .ZN(
        n20133) );
  INV_X1 U22255 ( .A(n20133), .ZN(n20135) );
  AOI22_X1 U22256 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20483), .B1(
        n20482), .B2(n20115), .ZN(n20134) );
  OAI211_X1 U22257 ( .C1(n20157), .C2(n20492), .A(n20135), .B(n20134), .ZN(
        P2_U3118) );
  AOI22_X1 U22258 ( .A1(n20487), .A2(n20115), .B1(n20486), .B2(n20153), .ZN(
        n20137) );
  AOI22_X1 U22259 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20489), .B1(
        n20495), .B2(n20147), .ZN(n20136) );
  OAI211_X1 U22260 ( .C1(n20145), .C2(n20492), .A(n20137), .B(n20136), .ZN(
        P2_U3110) );
  AOI22_X1 U22261 ( .A1(n20494), .A2(n20115), .B1(n20153), .B2(n20493), .ZN(
        n20139) );
  AOI22_X1 U22262 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20496), .B1(
        n20495), .B2(n20159), .ZN(n20138) );
  OAI211_X1 U22263 ( .C1(n20157), .C2(n20505), .A(n20139), .B(n20138), .ZN(
        P2_U3102) );
  AOI22_X1 U22264 ( .A1(n20404), .A2(n20159), .B1(n20153), .B2(n20403), .ZN(
        n20141) );
  AOI22_X1 U22265 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20502), .B1(
        n20115), .B2(n20501), .ZN(n20140) );
  OAI211_X1 U22266 ( .C1(n20157), .C2(n20507), .A(n20141), .B(n20140), .ZN(
        P2_U3094) );
  OAI22_X1 U22267 ( .A1(n20507), .A2(n20145), .B1(n20506), .B2(n20156), .ZN(
        n20142) );
  INV_X1 U22268 ( .A(n20142), .ZN(n20144) );
  AOI22_X1 U22269 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20510), .B1(
        n20115), .B2(n20509), .ZN(n20143) );
  OAI211_X1 U22270 ( .C1(n20157), .C2(n20515), .A(n20144), .B(n20143), .ZN(
        P2_U3086) );
  OAI22_X1 U22271 ( .A1(n20515), .A2(n20145), .B1(n20513), .B2(n20156), .ZN(
        n20146) );
  INV_X1 U22272 ( .A(n20146), .ZN(n20149) );
  AOI22_X1 U22273 ( .A1(n20115), .A2(n20517), .B1(n20524), .B2(n20147), .ZN(
        n20148) );
  OAI211_X1 U22274 ( .C1(n20206), .C2(n20150), .A(n20149), .B(n20148), .ZN(
        P2_U3078) );
  AOI22_X1 U22275 ( .A1(n20523), .A2(n20115), .B1(n20153), .B2(n20522), .ZN(
        n20152) );
  AOI22_X1 U22276 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20525), .B1(
        n20524), .B2(n20159), .ZN(n20151) );
  OAI211_X1 U22277 ( .C1(n20157), .C2(n20528), .A(n20152), .B(n20151), .ZN(
        P2_U3070) );
  AOI22_X1 U22278 ( .A1(n20531), .A2(n20115), .B1(n20153), .B2(n20529), .ZN(
        n20155) );
  AOI22_X1 U22279 ( .A1(n20533), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n20532), .B2(n20159), .ZN(n20154) );
  OAI211_X1 U22280 ( .C1(n20157), .C2(n20536), .A(n20155), .B(n20154), .ZN(
        P2_U3062) );
  OAI22_X1 U22281 ( .A1(n20540), .A2(n20157), .B1(n20538), .B2(n20156), .ZN(
        n20158) );
  INV_X1 U22282 ( .A(n20158), .ZN(n20161) );
  AOI22_X1 U22283 ( .A1(n20545), .A2(n20159), .B1(n20543), .B2(n20115), .ZN(
        n20160) );
  OAI211_X1 U22284 ( .C1(n20548), .C2(n20162), .A(n20161), .B(n20160), .ZN(
        P2_U3054) );
  AOI22_X1 U22285 ( .A1(n20164), .A2(n20163), .B1(n20319), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n20169) );
  OR3_X1 U22286 ( .A1(n20167), .A2(n20166), .A3(n20165), .ZN(n20168) );
  OAI211_X1 U22287 ( .C1(n20171), .C2(n20170), .A(n20169), .B(n20168), .ZN(
        P2_U2914) );
  AOI22_X2 U22288 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n20424), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n11143), .ZN(n20217) );
  NAND2_X1 U22289 ( .A1(n20174), .A2(n20428), .ZN(n20216) );
  AOI22_X1 U22290 ( .A1(n20431), .A2(n20173), .B1(n20430), .B2(n20211), .ZN(
        n20176) );
  AOI22_X1 U22291 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n11143), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n20424), .ZN(n20215) );
  INV_X1 U22292 ( .A(n20215), .ZN(n20219) );
  AOI22_X1 U22293 ( .A1(n20435), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n20274), .B2(n20219), .ZN(n20175) );
  OAI211_X1 U22294 ( .C1(n20217), .C2(n20439), .A(n20176), .B(n20175), .ZN(
        P2_U3173) );
  OAI22_X1 U22295 ( .A1(n20445), .A2(n20217), .B1(n20216), .B2(n20438), .ZN(
        n20177) );
  INV_X1 U22296 ( .A(n20177), .ZN(n20179) );
  AOI22_X1 U22297 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20442), .B1(
        n20173), .B2(n20441), .ZN(n20178) );
  OAI211_X1 U22298 ( .C1(n20215), .C2(n20439), .A(n20179), .B(n20178), .ZN(
        P2_U3165) );
  AOI22_X1 U22299 ( .A1(n20447), .A2(n20173), .B1(n20211), .B2(n20446), .ZN(
        n20181) );
  INV_X1 U22300 ( .A(n20217), .ZN(n20212) );
  AOI22_X1 U22301 ( .A1(n20449), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n20455), .B2(n20212), .ZN(n20180) );
  OAI211_X1 U22302 ( .C1(n20215), .C2(n20445), .A(n20181), .B(n20180), .ZN(
        P2_U3157) );
  AOI22_X1 U22303 ( .A1(n20454), .A2(n20173), .B1(n20211), .B2(n20453), .ZN(
        n20183) );
  AOI22_X1 U22304 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20219), .ZN(n20182) );
  OAI211_X1 U22305 ( .C1(n20217), .C2(n20464), .A(n20183), .B(n20182), .ZN(
        P2_U3149) );
  AOI22_X1 U22306 ( .A1(n20460), .A2(n20173), .B1(n20211), .B2(n20459), .ZN(
        n20185) );
  AOI22_X1 U22307 ( .A1(n20466), .A2(n20212), .B1(n20461), .B2(
        P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n20184) );
  OAI211_X1 U22308 ( .C1(n20215), .C2(n20464), .A(n20185), .B(n20184), .ZN(
        P2_U3141) );
  INV_X1 U22309 ( .A(n20465), .ZN(n20186) );
  OAI22_X1 U22310 ( .A1(n20478), .A2(n20217), .B1(n20216), .B2(n20186), .ZN(
        n20187) );
  INV_X1 U22311 ( .A(n20187), .ZN(n20189) );
  AOI22_X1 U22312 ( .A1(n20173), .A2(n20468), .B1(n20466), .B2(n20219), .ZN(
        n20188) );
  OAI211_X1 U22313 ( .C1(n20471), .C2(n16612), .A(n20189), .B(n20188), .ZN(
        P2_U3133) );
  OAI22_X1 U22314 ( .A1(n20480), .A2(n20217), .B1(n20472), .B2(n20216), .ZN(
        n20190) );
  INV_X1 U22315 ( .A(n20190), .ZN(n20192) );
  AOI22_X1 U22316 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20475), .B1(
        n20173), .B2(n20474), .ZN(n20191) );
  OAI211_X1 U22317 ( .C1(n20215), .C2(n20478), .A(n20192), .B(n20191), .ZN(
        P2_U3125) );
  OAI22_X1 U22318 ( .A1(n20480), .A2(n20215), .B1(n20216), .B2(n20479), .ZN(
        n20193) );
  INV_X1 U22319 ( .A(n20193), .ZN(n20195) );
  AOI22_X1 U22320 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20483), .B1(
        n20482), .B2(n20173), .ZN(n20194) );
  OAI211_X1 U22321 ( .C1(n20217), .C2(n20492), .A(n20195), .B(n20194), .ZN(
        P2_U3117) );
  AOI22_X1 U22322 ( .A1(n20487), .A2(n20173), .B1(n20486), .B2(n20211), .ZN(
        n20197) );
  INV_X1 U22323 ( .A(n20492), .ZN(n20351) );
  AOI22_X1 U22324 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20489), .B1(
        n20351), .B2(n20219), .ZN(n20196) );
  OAI211_X1 U22325 ( .C1(n20217), .C2(n20402), .A(n20197), .B(n20196), .ZN(
        P2_U3109) );
  AOI22_X1 U22326 ( .A1(n20494), .A2(n20173), .B1(n20211), .B2(n20493), .ZN(
        n20199) );
  AOI22_X1 U22327 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20496), .B1(
        n20495), .B2(n20219), .ZN(n20198) );
  OAI211_X1 U22328 ( .C1(n20217), .C2(n20505), .A(n20199), .B(n20198), .ZN(
        P2_U3101) );
  AOI22_X1 U22329 ( .A1(n20404), .A2(n20219), .B1(n20211), .B2(n20403), .ZN(
        n20201) );
  AOI22_X1 U22330 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20502), .B1(
        n20173), .B2(n20501), .ZN(n20200) );
  OAI211_X1 U22331 ( .C1(n20217), .C2(n20507), .A(n20201), .B(n20200), .ZN(
        P2_U3093) );
  OAI22_X1 U22332 ( .A1(n20507), .A2(n20215), .B1(n20506), .B2(n20216), .ZN(
        n20202) );
  INV_X1 U22333 ( .A(n20202), .ZN(n20204) );
  AOI22_X1 U22334 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20510), .B1(
        n20173), .B2(n20509), .ZN(n20203) );
  OAI211_X1 U22335 ( .C1(n20217), .C2(n20515), .A(n20204), .B(n20203), .ZN(
        P2_U3085) );
  OAI22_X1 U22336 ( .A1(n20515), .A2(n20215), .B1(n20513), .B2(n20216), .ZN(
        n20205) );
  INV_X1 U22337 ( .A(n20205), .ZN(n20208) );
  INV_X1 U22338 ( .A(n20206), .ZN(n20518) );
  AOI22_X1 U22339 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20518), .B1(
        n20173), .B2(n20517), .ZN(n20207) );
  OAI211_X1 U22340 ( .C1(n20217), .C2(n20521), .A(n20208), .B(n20207), .ZN(
        P2_U3077) );
  AOI22_X1 U22341 ( .A1(n20523), .A2(n20173), .B1(n20211), .B2(n20522), .ZN(
        n20210) );
  AOI22_X1 U22342 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20525), .B1(
        n20532), .B2(n20212), .ZN(n20209) );
  OAI211_X1 U22343 ( .C1(n20215), .C2(n20521), .A(n20210), .B(n20209), .ZN(
        P2_U3069) );
  AOI22_X1 U22344 ( .A1(n20531), .A2(n20173), .B1(n20211), .B2(n20529), .ZN(
        n20214) );
  AOI22_X1 U22345 ( .A1(n20533), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n20545), .B2(n20212), .ZN(n20213) );
  OAI211_X1 U22346 ( .C1(n20215), .C2(n20528), .A(n20214), .B(n20213), .ZN(
        P2_U3061) );
  OAI22_X1 U22347 ( .A1(n20540), .A2(n20217), .B1(n20538), .B2(n20216), .ZN(
        n20218) );
  INV_X1 U22348 ( .A(n20218), .ZN(n20221) );
  AOI22_X1 U22349 ( .A1(n20545), .A2(n20219), .B1(n20543), .B2(n20173), .ZN(
        n20220) );
  OAI211_X1 U22350 ( .C1(n20548), .C2(n16601), .A(n20221), .B(n20220), .ZN(
        P2_U3053) );
  OAI22_X1 U22351 ( .A1(n20316), .A2(n20230), .B1(n20222), .B2(n20327), .ZN(
        n20223) );
  AOI21_X1 U22352 ( .B1(P2_EAX_REG_20__SCAN_IN), .B2(n20319), .A(n20223), .ZN(
        n20229) );
  INV_X1 U22353 ( .A(n20224), .ZN(n20227) );
  INV_X1 U22354 ( .A(n20225), .ZN(n20226) );
  AOI22_X1 U22355 ( .A1(n20227), .A2(n20322), .B1(n20321), .B2(n20226), .ZN(
        n20228) );
  OAI211_X1 U22356 ( .C1(n20317), .C2(n20805), .A(n20229), .B(n20228), .ZN(
        P2_U2899) );
  INV_X1 U22357 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n21473) );
  OAI22_X1 U22358 ( .A1(n21473), .A2(n20432), .B1(n20822), .B2(n20433), .ZN(
        n20269) );
  NOR2_X2 U22359 ( .A1(n20233), .A2(n20232), .ZN(n20267) );
  AOI22_X1 U22360 ( .A1(n20431), .A2(n20231), .B1(n20430), .B2(n20267), .ZN(
        n20235) );
  AOI22_X1 U22361 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n11143), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n20424), .ZN(n20249) );
  AOI22_X1 U22362 ( .A1(n20270), .A2(n20274), .B1(
        P2_INSTQUEUE_REG_15__4__SCAN_IN), .B2(n20435), .ZN(n20234) );
  OAI211_X1 U22363 ( .C1(n20266), .C2(n20439), .A(n20235), .B(n20234), .ZN(
        P2_U3172) );
  AOI22_X1 U22364 ( .A1(n20270), .A2(n20434), .B1(n20267), .B2(n20236), .ZN(
        n20238) );
  AOI22_X1 U22365 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20442), .B1(
        n20231), .B2(n20441), .ZN(n20237) );
  OAI211_X1 U22366 ( .C1(n20266), .C2(n20445), .A(n20238), .B(n20237), .ZN(
        P2_U3164) );
  AOI22_X1 U22367 ( .A1(n20447), .A2(n20231), .B1(n20267), .B2(n20446), .ZN(
        n20240) );
  AOI22_X1 U22368 ( .A1(n20269), .A2(n20455), .B1(n20449), .B2(
        P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n20239) );
  OAI211_X1 U22369 ( .C1(n20249), .C2(n20445), .A(n20240), .B(n20239), .ZN(
        P2_U3156) );
  AOI22_X1 U22370 ( .A1(n20454), .A2(n20231), .B1(n20267), .B2(n20453), .ZN(
        n20242) );
  AOI22_X1 U22371 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20270), .ZN(n20241) );
  OAI211_X1 U22372 ( .C1(n20266), .C2(n20464), .A(n20242), .B(n20241), .ZN(
        P2_U3148) );
  AOI22_X1 U22373 ( .A1(n20460), .A2(n20231), .B1(n20267), .B2(n20459), .ZN(
        n20244) );
  AOI22_X1 U22374 ( .A1(n20269), .A2(n20466), .B1(
        P2_INSTQUEUE_REG_11__4__SCAN_IN), .B2(n20461), .ZN(n20243) );
  OAI211_X1 U22375 ( .C1(n20249), .C2(n20464), .A(n20244), .B(n20243), .ZN(
        P2_U3140) );
  AOI22_X1 U22376 ( .A1(n20269), .A2(n20467), .B1(n20267), .B2(n20465), .ZN(
        n20246) );
  AOI22_X1 U22377 ( .A1(n20231), .A2(n20468), .B1(n20466), .B2(n20270), .ZN(
        n20245) );
  OAI211_X1 U22378 ( .C1(n20471), .C2(n16589), .A(n20246), .B(n20245), .ZN(
        P2_U3132) );
  INV_X1 U22379 ( .A(n20480), .ZN(n20348) );
  AOI22_X1 U22380 ( .A1(n20269), .A2(n20348), .B1(n20344), .B2(n20267), .ZN(
        n20248) );
  AOI22_X1 U22381 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20475), .B1(
        n20231), .B2(n20474), .ZN(n20247) );
  OAI211_X1 U22382 ( .C1(n20249), .C2(n20478), .A(n20248), .B(n20247), .ZN(
        P2_U3124) );
  AOI22_X1 U22383 ( .A1(n20270), .A2(n20348), .B1(n20267), .B2(n20347), .ZN(
        n20251) );
  AOI22_X1 U22384 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20483), .B1(
        n20482), .B2(n20231), .ZN(n20250) );
  OAI211_X1 U22385 ( .C1(n20266), .C2(n20492), .A(n20251), .B(n20250), .ZN(
        P2_U3116) );
  AOI22_X1 U22386 ( .A1(n20487), .A2(n20231), .B1(n20486), .B2(n20267), .ZN(
        n20253) );
  AOI22_X1 U22387 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20489), .B1(
        n20351), .B2(n20270), .ZN(n20252) );
  OAI211_X1 U22388 ( .C1(n20266), .C2(n20402), .A(n20253), .B(n20252), .ZN(
        P2_U3108) );
  AOI22_X1 U22389 ( .A1(n20494), .A2(n20231), .B1(n20267), .B2(n20493), .ZN(
        n20255) );
  AOI22_X1 U22390 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20496), .B1(
        n20495), .B2(n20270), .ZN(n20254) );
  OAI211_X1 U22391 ( .C1(n20266), .C2(n20505), .A(n20255), .B(n20254), .ZN(
        P2_U3100) );
  AOI22_X1 U22392 ( .A1(n20270), .A2(n20404), .B1(n20267), .B2(n20403), .ZN(
        n20257) );
  AOI22_X1 U22393 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20502), .B1(
        n20231), .B2(n20501), .ZN(n20256) );
  OAI211_X1 U22394 ( .C1(n20266), .C2(n20507), .A(n20257), .B(n20256), .ZN(
        P2_U3092) );
  AOI22_X1 U22395 ( .A1(n20270), .A2(n20359), .B1(n20358), .B2(n20267), .ZN(
        n20259) );
  AOI22_X1 U22396 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20510), .B1(
        n20231), .B2(n20509), .ZN(n20258) );
  OAI211_X1 U22397 ( .C1(n20266), .C2(n20515), .A(n20259), .B(n20258), .ZN(
        P2_U3084) );
  AOI22_X1 U22398 ( .A1(n20270), .A2(n20362), .B1(n20411), .B2(n20267), .ZN(
        n20261) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20518), .B1(
        n20231), .B2(n20517), .ZN(n20260) );
  OAI211_X1 U22400 ( .C1(n20266), .C2(n20521), .A(n20261), .B(n20260), .ZN(
        P2_U3076) );
  AOI22_X1 U22401 ( .A1(n20523), .A2(n20231), .B1(n20267), .B2(n20522), .ZN(
        n20263) );
  AOI22_X1 U22402 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20525), .B1(
        n20524), .B2(n20270), .ZN(n20262) );
  OAI211_X1 U22403 ( .C1(n20266), .C2(n20528), .A(n20263), .B(n20262), .ZN(
        P2_U3068) );
  AOI22_X1 U22404 ( .A1(n20531), .A2(n20231), .B1(n20267), .B2(n20529), .ZN(
        n20265) );
  AOI22_X1 U22405 ( .A1(n20270), .A2(n20532), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n20533), .ZN(n20264) );
  OAI211_X1 U22406 ( .C1(n20266), .C2(n20536), .A(n20265), .B(n20264), .ZN(
        P2_U3060) );
  AOI22_X1 U22407 ( .A1(n20269), .A2(n20274), .B1(n20268), .B2(n20267), .ZN(
        n20272) );
  AOI22_X1 U22408 ( .A1(n20545), .A2(n20270), .B1(n20543), .B2(n20231), .ZN(
        n20271) );
  OAI211_X1 U22409 ( .C1(n20548), .C2(n20273), .A(n20272), .B(n20271), .ZN(
        P2_U3052) );
  AOI22_X1 U22410 ( .A1(n20431), .A2(n16029), .B1(n20430), .B2(n20311), .ZN(
        n20276) );
  INV_X1 U22411 ( .A(n20310), .ZN(n20312) );
  AOI22_X1 U22412 ( .A1(n20435), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n20274), .B2(n20312), .ZN(n20275) );
  OAI211_X1 U22413 ( .C1(n20315), .C2(n20439), .A(n20276), .B(n20275), .ZN(
        P2_U3171) );
  INV_X1 U22414 ( .A(n20311), .ZN(n20301) );
  OAI22_X1 U22415 ( .A1(n20445), .A2(n20315), .B1(n20301), .B2(n20438), .ZN(
        n20277) );
  INV_X1 U22416 ( .A(n20277), .ZN(n20279) );
  AOI22_X1 U22417 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20442), .B1(
        n16029), .B2(n20441), .ZN(n20278) );
  OAI211_X1 U22418 ( .C1(n20310), .C2(n20439), .A(n20279), .B(n20278), .ZN(
        P2_U3163) );
  AOI22_X1 U22419 ( .A1(n20447), .A2(n16029), .B1(n20311), .B2(n20446), .ZN(
        n20281) );
  AOI22_X1 U22420 ( .A1(n20449), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n20455), .B2(n20307), .ZN(n20280) );
  OAI211_X1 U22421 ( .C1(n20310), .C2(n20445), .A(n20281), .B(n20280), .ZN(
        P2_U3155) );
  AOI22_X1 U22422 ( .A1(n20454), .A2(n16029), .B1(n20311), .B2(n20453), .ZN(
        n20283) );
  AOI22_X1 U22423 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20312), .ZN(n20282) );
  OAI211_X1 U22424 ( .C1(n20315), .C2(n20464), .A(n20283), .B(n20282), .ZN(
        P2_U3147) );
  AOI22_X1 U22425 ( .A1(n20460), .A2(n16029), .B1(n20311), .B2(n20459), .ZN(
        n20285) );
  AOI22_X1 U22426 ( .A1(n20466), .A2(n20307), .B1(n20461), .B2(
        P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n20284) );
  OAI211_X1 U22427 ( .C1(n20310), .C2(n20464), .A(n20285), .B(n20284), .ZN(
        P2_U3139) );
  AOI22_X1 U22428 ( .A1(n20466), .A2(n20312), .B1(n20465), .B2(n20311), .ZN(
        n20287) );
  AOI22_X1 U22429 ( .A1(n16029), .A2(n20468), .B1(n20467), .B2(n20307), .ZN(
        n20286) );
  OAI211_X1 U22430 ( .C1(n20471), .C2(n16227), .A(n20287), .B(n20286), .ZN(
        P2_U3131) );
  OAI22_X1 U22431 ( .A1(n20478), .A2(n20310), .B1(n20472), .B2(n20301), .ZN(
        n20288) );
  INV_X1 U22432 ( .A(n20288), .ZN(n20290) );
  AOI22_X1 U22433 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20475), .B1(
        n16029), .B2(n20474), .ZN(n20289) );
  OAI211_X1 U22434 ( .C1(n20315), .C2(n20480), .A(n20290), .B(n20289), .ZN(
        P2_U3123) );
  OAI22_X1 U22435 ( .A1(n20480), .A2(n20310), .B1(n20479), .B2(n20301), .ZN(
        n20291) );
  INV_X1 U22436 ( .A(n20291), .ZN(n20293) );
  AOI22_X1 U22437 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20483), .B1(
        n20482), .B2(n16029), .ZN(n20292) );
  OAI211_X1 U22438 ( .C1(n20315), .C2(n20492), .A(n20293), .B(n20292), .ZN(
        P2_U3115) );
  AOI22_X1 U22439 ( .A1(n20487), .A2(n16029), .B1(n20311), .B2(n20486), .ZN(
        n20295) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20489), .B1(
        n20351), .B2(n20312), .ZN(n20294) );
  OAI211_X1 U22441 ( .C1(n20315), .C2(n20402), .A(n20295), .B(n20294), .ZN(
        P2_U3107) );
  AOI22_X1 U22442 ( .A1(n20494), .A2(n16029), .B1(n20311), .B2(n20493), .ZN(
        n20297) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20496), .B1(
        n20495), .B2(n20312), .ZN(n20296) );
  OAI211_X1 U22444 ( .C1(n20315), .C2(n20505), .A(n20297), .B(n20296), .ZN(
        P2_U3099) );
  INV_X1 U22445 ( .A(n20403), .ZN(n20499) );
  OAI22_X1 U22446 ( .A1(n20507), .A2(n20315), .B1(n20301), .B2(n20499), .ZN(
        n20298) );
  INV_X1 U22447 ( .A(n20298), .ZN(n20300) );
  AOI22_X1 U22448 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20502), .B1(
        n16029), .B2(n20501), .ZN(n20299) );
  OAI211_X1 U22449 ( .C1(n20310), .C2(n20505), .A(n20300), .B(n20299), .ZN(
        P2_U3091) );
  OAI22_X1 U22450 ( .A1(n20507), .A2(n20310), .B1(n20506), .B2(n20301), .ZN(
        n20302) );
  INV_X1 U22451 ( .A(n20302), .ZN(n20304) );
  AOI22_X1 U22452 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20510), .B1(
        n16029), .B2(n20509), .ZN(n20303) );
  OAI211_X1 U22453 ( .C1(n20315), .C2(n20515), .A(n20304), .B(n20303), .ZN(
        P2_U3083) );
  AOI22_X1 U22454 ( .A1(n20524), .A2(n20307), .B1(n20311), .B2(n20411), .ZN(
        n20306) );
  AOI22_X1 U22455 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20518), .B1(
        n16029), .B2(n20517), .ZN(n20305) );
  OAI211_X1 U22456 ( .C1(n20310), .C2(n20515), .A(n20306), .B(n20305), .ZN(
        P2_U3075) );
  AOI22_X1 U22457 ( .A1(n20523), .A2(n16029), .B1(n20311), .B2(n20522), .ZN(
        n20309) );
  AOI22_X1 U22458 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20525), .B1(
        n20532), .B2(n20307), .ZN(n20308) );
  OAI211_X1 U22459 ( .C1(n20310), .C2(n20521), .A(n20309), .B(n20308), .ZN(
        P2_U3067) );
  AOI22_X1 U22460 ( .A1(n20531), .A2(n16029), .B1(n20311), .B2(n20529), .ZN(
        n20314) );
  AOI22_X1 U22461 ( .A1(n20533), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n20532), .B2(n20312), .ZN(n20313) );
  OAI211_X1 U22462 ( .C1(n20315), .C2(n20536), .A(n20314), .B(n20313), .ZN(
        P2_U3059) );
  OAI22_X1 U22463 ( .A1(n20317), .A2(n20801), .B1(n20316), .B2(n20328), .ZN(
        n20318) );
  AOI21_X1 U22464 ( .B1(P2_EAX_REG_18__SCAN_IN), .B2(n20319), .A(n20318), .ZN(
        n20325) );
  AOI22_X1 U22465 ( .A1(n20323), .A2(n20322), .B1(n20321), .B2(n20320), .ZN(
        n20324) );
  OAI211_X1 U22466 ( .C1(n20327), .C2(n20326), .A(n20325), .B(n20324), .ZN(
        P2_U2901) );
  AOI22_X1 U22467 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n11143), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20424), .ZN(n20371) );
  AND2_X1 U22468 ( .A1(n20330), .A2(n20428), .ZN(n20367) );
  AOI22_X1 U22469 ( .A1(n20431), .A2(n20329), .B1(n20430), .B2(n20367), .ZN(
        n20332) );
  INV_X1 U22470 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n21454) );
  OAI22_X1 U22471 ( .A1(n20818), .A2(n20433), .B1(n21454), .B2(n20432), .ZN(
        n20368) );
  AOI22_X1 U22472 ( .A1(n20435), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n20434), .B2(n20368), .ZN(n20331) );
  OAI211_X1 U22473 ( .C1(n20371), .C2(n20540), .A(n20332), .B(n20331), .ZN(
        P2_U3170) );
  INV_X1 U22474 ( .A(n20367), .ZN(n20372) );
  OAI22_X1 U22475 ( .A1(n20445), .A2(n20373), .B1(n20372), .B2(n20438), .ZN(
        n20333) );
  INV_X1 U22476 ( .A(n20333), .ZN(n20335) );
  AOI22_X1 U22477 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20442), .B1(
        n20329), .B2(n20441), .ZN(n20334) );
  OAI211_X1 U22478 ( .C1(n20371), .C2(n20439), .A(n20335), .B(n20334), .ZN(
        P2_U3162) );
  AOI22_X1 U22479 ( .A1(n20447), .A2(n20329), .B1(n20367), .B2(n20446), .ZN(
        n20337) );
  AOI22_X1 U22480 ( .A1(n20375), .A2(n20448), .B1(
        P2_INSTQUEUE_REG_13__2__SCAN_IN), .B2(n20449), .ZN(n20336) );
  OAI211_X1 U22481 ( .C1(n20373), .C2(n20452), .A(n20337), .B(n20336), .ZN(
        P2_U3154) );
  AOI22_X1 U22482 ( .A1(n20454), .A2(n20329), .B1(n20367), .B2(n20453), .ZN(
        n20339) );
  AOI22_X1 U22483 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20375), .ZN(n20338) );
  OAI211_X1 U22484 ( .C1(n20373), .C2(n20464), .A(n20339), .B(n20338), .ZN(
        P2_U3146) );
  AOI22_X1 U22485 ( .A1(n20460), .A2(n20329), .B1(n20367), .B2(n20459), .ZN(
        n20341) );
  AOI22_X1 U22486 ( .A1(n20466), .A2(n20368), .B1(n20461), .B2(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n20340) );
  OAI211_X1 U22487 ( .C1(n20371), .C2(n20464), .A(n20341), .B(n20340), .ZN(
        P2_U3138) );
  AOI22_X1 U22488 ( .A1(n20375), .A2(n20466), .B1(n20367), .B2(n20465), .ZN(
        n20343) );
  AOI22_X1 U22489 ( .A1(n20329), .A2(n20468), .B1(n20467), .B2(n20368), .ZN(
        n20342) );
  OAI211_X1 U22490 ( .C1(n20471), .C2(n16544), .A(n20343), .B(n20342), .ZN(
        P2_U3130) );
  AOI22_X1 U22491 ( .A1(n20375), .A2(n20467), .B1(n20344), .B2(n20367), .ZN(
        n20346) );
  AOI22_X1 U22492 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20475), .B1(
        n20329), .B2(n20474), .ZN(n20345) );
  OAI211_X1 U22493 ( .C1(n20373), .C2(n20480), .A(n20346), .B(n20345), .ZN(
        P2_U3122) );
  AOI22_X1 U22494 ( .A1(n20375), .A2(n20348), .B1(n20367), .B2(n20347), .ZN(
        n20350) );
  AOI22_X1 U22495 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20483), .B1(
        n20482), .B2(n20329), .ZN(n20349) );
  OAI211_X1 U22496 ( .C1(n20373), .C2(n20492), .A(n20350), .B(n20349), .ZN(
        P2_U3114) );
  AOI22_X1 U22497 ( .A1(n20487), .A2(n20329), .B1(n20486), .B2(n20367), .ZN(
        n20353) );
  AOI22_X1 U22498 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20489), .B1(
        n20351), .B2(n20375), .ZN(n20352) );
  OAI211_X1 U22499 ( .C1(n20373), .C2(n20402), .A(n20353), .B(n20352), .ZN(
        P2_U3106) );
  AOI22_X1 U22500 ( .A1(n20494), .A2(n20329), .B1(n20367), .B2(n20493), .ZN(
        n20355) );
  AOI22_X1 U22501 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20496), .B1(
        n20404), .B2(n20368), .ZN(n20354) );
  OAI211_X1 U22502 ( .C1(n20371), .C2(n20402), .A(n20355), .B(n20354), .ZN(
        P2_U3098) );
  AOI22_X1 U22503 ( .A1(n20375), .A2(n20404), .B1(n20367), .B2(n20403), .ZN(
        n20357) );
  AOI22_X1 U22504 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20502), .B1(
        n20329), .B2(n20501), .ZN(n20356) );
  OAI211_X1 U22505 ( .C1(n20373), .C2(n20507), .A(n20357), .B(n20356), .ZN(
        P2_U3090) );
  AOI22_X1 U22506 ( .A1(n20375), .A2(n20359), .B1(n20358), .B2(n20367), .ZN(
        n20361) );
  AOI22_X1 U22507 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20510), .B1(
        n20329), .B2(n20509), .ZN(n20360) );
  OAI211_X1 U22508 ( .C1(n20373), .C2(n20515), .A(n20361), .B(n20360), .ZN(
        P2_U3082) );
  AOI22_X1 U22509 ( .A1(n20375), .A2(n20362), .B1(n20411), .B2(n20367), .ZN(
        n20364) );
  AOI22_X1 U22510 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20518), .B1(
        n20329), .B2(n20517), .ZN(n20363) );
  OAI211_X1 U22511 ( .C1(n20373), .C2(n20521), .A(n20364), .B(n20363), .ZN(
        P2_U3074) );
  AOI22_X1 U22512 ( .A1(n20523), .A2(n20329), .B1(n20367), .B2(n20522), .ZN(
        n20366) );
  AOI22_X1 U22513 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20525), .B1(
        n20524), .B2(n20375), .ZN(n20365) );
  OAI211_X1 U22514 ( .C1(n20373), .C2(n20528), .A(n20366), .B(n20365), .ZN(
        P2_U3066) );
  AOI22_X1 U22515 ( .A1(n20531), .A2(n20329), .B1(n20367), .B2(n20529), .ZN(
        n20370) );
  AOI22_X1 U22516 ( .A1(n20533), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n20545), .B2(n20368), .ZN(n20369) );
  OAI211_X1 U22517 ( .C1(n20371), .C2(n20528), .A(n20370), .B(n20369), .ZN(
        P2_U3058) );
  OAI22_X1 U22518 ( .A1(n20540), .A2(n20373), .B1(n20538), .B2(n20372), .ZN(
        n20374) );
  INV_X1 U22519 ( .A(n20374), .ZN(n20377) );
  AOI22_X1 U22520 ( .A1(n20545), .A2(n20375), .B1(n20543), .B2(n20329), .ZN(
        n20376) );
  OAI211_X1 U22521 ( .C1(n20548), .C2(n20378), .A(n20377), .B(n20376), .ZN(
        P2_U3050) );
  AOI22_X1 U22522 ( .A1(n20431), .A2(n20419), .B1(n20430), .B2(n20418), .ZN(
        n20380) );
  AOI22_X1 U22523 ( .A1(n20435), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n20434), .B2(n20412), .ZN(n20379) );
  OAI211_X1 U22524 ( .C1(n20415), .C2(n20540), .A(n20380), .B(n20379), .ZN(
        P2_U3169) );
  INV_X1 U22525 ( .A(n20418), .ZN(n20407) );
  OAI22_X1 U22526 ( .A1(n20445), .A2(n20423), .B1(n20407), .B2(n20438), .ZN(
        n20381) );
  INV_X1 U22527 ( .A(n20381), .ZN(n20383) );
  AOI22_X1 U22528 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20442), .B1(
        n20419), .B2(n20441), .ZN(n20382) );
  OAI211_X1 U22529 ( .C1(n20415), .C2(n20439), .A(n20383), .B(n20382), .ZN(
        P2_U3161) );
  AOI22_X1 U22530 ( .A1(n20447), .A2(n20419), .B1(n20418), .B2(n20446), .ZN(
        n20385) );
  AOI22_X1 U22531 ( .A1(n20449), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n20455), .B2(n20412), .ZN(n20384) );
  OAI211_X1 U22532 ( .C1(n20415), .C2(n20445), .A(n20385), .B(n20384), .ZN(
        P2_U3153) );
  AOI22_X1 U22533 ( .A1(n20454), .A2(n20419), .B1(n20418), .B2(n20453), .ZN(
        n20387) );
  INV_X1 U22534 ( .A(n20415), .ZN(n20420) );
  AOI22_X1 U22535 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20420), .ZN(n20386) );
  OAI211_X1 U22536 ( .C1(n20423), .C2(n20464), .A(n20387), .B(n20386), .ZN(
        P2_U3145) );
  AOI22_X1 U22537 ( .A1(n20460), .A2(n20419), .B1(n20418), .B2(n20459), .ZN(
        n20389) );
  AOI22_X1 U22538 ( .A1(n20466), .A2(n20412), .B1(n20461), .B2(
        P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n20388) );
  OAI211_X1 U22539 ( .C1(n20415), .C2(n20464), .A(n20389), .B(n20388), .ZN(
        P2_U3137) );
  AOI22_X1 U22540 ( .A1(n20466), .A2(n20420), .B1(n20465), .B2(n20418), .ZN(
        n20391) );
  AOI22_X1 U22541 ( .A1(n20419), .A2(n20468), .B1(n20467), .B2(n20412), .ZN(
        n20390) );
  OAI211_X1 U22542 ( .C1(n20471), .C2(n16524), .A(n20391), .B(n20390), .ZN(
        P2_U3129) );
  OAI22_X1 U22543 ( .A1(n20478), .A2(n20415), .B1(n20472), .B2(n20407), .ZN(
        n20392) );
  INV_X1 U22544 ( .A(n20392), .ZN(n20394) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20475), .B1(
        n20419), .B2(n20474), .ZN(n20393) );
  OAI211_X1 U22546 ( .C1(n20423), .C2(n20480), .A(n20394), .B(n20393), .ZN(
        P2_U3121) );
  OAI22_X1 U22547 ( .A1(n20480), .A2(n20415), .B1(n20479), .B2(n20407), .ZN(
        n20395) );
  INV_X1 U22548 ( .A(n20395), .ZN(n20397) );
  AOI22_X1 U22549 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20483), .B1(
        n20482), .B2(n20419), .ZN(n20396) );
  OAI211_X1 U22550 ( .C1(n20423), .C2(n20492), .A(n20397), .B(n20396), .ZN(
        P2_U3113) );
  AOI22_X1 U22551 ( .A1(n20487), .A2(n20419), .B1(n20418), .B2(n20486), .ZN(
        n20399) );
  AOI22_X1 U22552 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20489), .B1(
        n20495), .B2(n20412), .ZN(n20398) );
  OAI211_X1 U22553 ( .C1(n20415), .C2(n20492), .A(n20399), .B(n20398), .ZN(
        P2_U3105) );
  AOI22_X1 U22554 ( .A1(n20494), .A2(n20419), .B1(n20418), .B2(n20493), .ZN(
        n20401) );
  AOI22_X1 U22555 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20496), .B1(
        n20404), .B2(n20412), .ZN(n20400) );
  OAI211_X1 U22556 ( .C1(n20415), .C2(n20402), .A(n20401), .B(n20400), .ZN(
        P2_U3097) );
  AOI22_X1 U22557 ( .A1(n20404), .A2(n20420), .B1(n20403), .B2(n20418), .ZN(
        n20406) );
  AOI22_X1 U22558 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20502), .B1(
        n20419), .B2(n20501), .ZN(n20405) );
  OAI211_X1 U22559 ( .C1(n20423), .C2(n20507), .A(n20406), .B(n20405), .ZN(
        P2_U3089) );
  OAI22_X1 U22560 ( .A1(n20507), .A2(n20415), .B1(n20506), .B2(n20407), .ZN(
        n20408) );
  INV_X1 U22561 ( .A(n20408), .ZN(n20410) );
  AOI22_X1 U22562 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20510), .B1(
        n20419), .B2(n20509), .ZN(n20409) );
  OAI211_X1 U22563 ( .C1(n20423), .C2(n20515), .A(n20410), .B(n20409), .ZN(
        P2_U3081) );
  AOI22_X1 U22564 ( .A1(n20524), .A2(n20412), .B1(n20418), .B2(n20411), .ZN(
        n20414) );
  AOI22_X1 U22565 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20518), .B1(
        n20419), .B2(n20517), .ZN(n20413) );
  OAI211_X1 U22566 ( .C1(n20415), .C2(n20515), .A(n20414), .B(n20413), .ZN(
        P2_U3073) );
  AOI22_X1 U22567 ( .A1(n20523), .A2(n20419), .B1(n20418), .B2(n20522), .ZN(
        n20417) );
  AOI22_X1 U22568 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20525), .B1(
        n20524), .B2(n20420), .ZN(n20416) );
  OAI211_X1 U22569 ( .C1(n20423), .C2(n20528), .A(n20417), .B(n20416), .ZN(
        P2_U3065) );
  AOI22_X1 U22570 ( .A1(n20531), .A2(n20419), .B1(n20418), .B2(n20529), .ZN(
        n20422) );
  AOI22_X1 U22571 ( .A1(n20533), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n20532), .B2(n20420), .ZN(n20421) );
  OAI211_X1 U22572 ( .C1(n20423), .C2(n20536), .A(n20422), .B(n20421), .ZN(
        P2_U3057) );
  AOI22_X1 U22573 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n11143), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20424), .ZN(n20514) );
  NOR2_X2 U22574 ( .A1(n20427), .A2(n20426), .ZN(n20542) );
  NAND2_X1 U22575 ( .A1(n20429), .A2(n20428), .ZN(n20537) );
  AOI22_X1 U22576 ( .A1(n20431), .A2(n20542), .B1(n20430), .B2(n20530), .ZN(
        n20437) );
  OAI22_X1 U22577 ( .A1(n20814), .A2(n20433), .B1(n21484), .B2(n20432), .ZN(
        n20488) );
  AOI22_X1 U22578 ( .A1(n20435), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n20434), .B2(n20488), .ZN(n20436) );
  OAI211_X1 U22579 ( .C1(n20514), .C2(n20540), .A(n20437), .B(n20436), .ZN(
        P2_U3168) );
  OAI22_X1 U22580 ( .A1(n20439), .A2(n20514), .B1(n20537), .B2(n20438), .ZN(
        n20440) );
  INV_X1 U22581 ( .A(n20440), .ZN(n20444) );
  AOI22_X1 U22582 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20442), .B1(
        n20542), .B2(n20441), .ZN(n20443) );
  OAI211_X1 U22583 ( .C1(n20539), .C2(n20445), .A(n20444), .B(n20443), .ZN(
        P2_U3160) );
  AOI22_X1 U22584 ( .A1(n20447), .A2(n20542), .B1(n20530), .B2(n20446), .ZN(
        n20451) );
  INV_X1 U22585 ( .A(n20514), .ZN(n20544) );
  AOI22_X1 U22586 ( .A1(n20449), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n20448), .B2(n20544), .ZN(n20450) );
  OAI211_X1 U22587 ( .C1(n20539), .C2(n20452), .A(n20451), .B(n20450), .ZN(
        P2_U3152) );
  AOI22_X1 U22588 ( .A1(n20454), .A2(n20542), .B1(n20530), .B2(n20453), .ZN(
        n20458) );
  AOI22_X1 U22589 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20456), .B1(
        n20455), .B2(n20544), .ZN(n20457) );
  OAI211_X1 U22590 ( .C1(n20539), .C2(n20464), .A(n20458), .B(n20457), .ZN(
        P2_U3144) );
  AOI22_X1 U22591 ( .A1(n20460), .A2(n20542), .B1(n20530), .B2(n20459), .ZN(
        n20463) );
  AOI22_X1 U22592 ( .A1(n20466), .A2(n20488), .B1(n20461), .B2(
        P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n20462) );
  OAI211_X1 U22593 ( .C1(n20514), .C2(n20464), .A(n20463), .B(n20462), .ZN(
        P2_U3136) );
  AOI22_X1 U22594 ( .A1(n20466), .A2(n20544), .B1(n20530), .B2(n20465), .ZN(
        n20470) );
  AOI22_X1 U22595 ( .A1(n20542), .A2(n20468), .B1(n20467), .B2(n20488), .ZN(
        n20469) );
  OAI211_X1 U22596 ( .C1(n20471), .C2(n16504), .A(n20470), .B(n20469), .ZN(
        P2_U3128) );
  OAI22_X1 U22597 ( .A1(n20480), .A2(n20539), .B1(n20472), .B2(n20537), .ZN(
        n20473) );
  INV_X1 U22598 ( .A(n20473), .ZN(n20477) );
  AOI22_X1 U22599 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20475), .B1(
        n20542), .B2(n20474), .ZN(n20476) );
  OAI211_X1 U22600 ( .C1(n20514), .C2(n20478), .A(n20477), .B(n20476), .ZN(
        P2_U3120) );
  OAI22_X1 U22601 ( .A1(n20480), .A2(n20514), .B1(n20537), .B2(n20479), .ZN(
        n20481) );
  INV_X1 U22602 ( .A(n20481), .ZN(n20485) );
  AOI22_X1 U22603 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20483), .B1(
        n20482), .B2(n20542), .ZN(n20484) );
  OAI211_X1 U22604 ( .C1(n20539), .C2(n20492), .A(n20485), .B(n20484), .ZN(
        P2_U3112) );
  AOI22_X1 U22605 ( .A1(n20487), .A2(n20542), .B1(n20486), .B2(n20530), .ZN(
        n20491) );
  AOI22_X1 U22606 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20489), .B1(
        n20495), .B2(n20488), .ZN(n20490) );
  OAI211_X1 U22607 ( .C1(n20514), .C2(n20492), .A(n20491), .B(n20490), .ZN(
        P2_U3104) );
  AOI22_X1 U22608 ( .A1(n20494), .A2(n20542), .B1(n20530), .B2(n20493), .ZN(
        n20498) );
  AOI22_X1 U22609 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20496), .B1(
        n20495), .B2(n20544), .ZN(n20497) );
  OAI211_X1 U22610 ( .C1(n20539), .C2(n20505), .A(n20498), .B(n20497), .ZN(
        P2_U3096) );
  OAI22_X1 U22611 ( .A1(n20507), .A2(n20539), .B1(n20499), .B2(n20537), .ZN(
        n20500) );
  INV_X1 U22612 ( .A(n20500), .ZN(n20504) );
  AOI22_X1 U22613 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20502), .B1(
        n20542), .B2(n20501), .ZN(n20503) );
  OAI211_X1 U22614 ( .C1(n20514), .C2(n20505), .A(n20504), .B(n20503), .ZN(
        P2_U3088) );
  OAI22_X1 U22615 ( .A1(n20507), .A2(n20514), .B1(n20506), .B2(n20537), .ZN(
        n20508) );
  INV_X1 U22616 ( .A(n20508), .ZN(n20512) );
  AOI22_X1 U22617 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20510), .B1(
        n20542), .B2(n20509), .ZN(n20511) );
  OAI211_X1 U22618 ( .C1(n20539), .C2(n20515), .A(n20512), .B(n20511), .ZN(
        P2_U3080) );
  OAI22_X1 U22619 ( .A1(n20515), .A2(n20514), .B1(n20513), .B2(n20537), .ZN(
        n20516) );
  INV_X1 U22620 ( .A(n20516), .ZN(n20520) );
  AOI22_X1 U22621 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20518), .B1(
        n20542), .B2(n20517), .ZN(n20519) );
  OAI211_X1 U22622 ( .C1(n20539), .C2(n20521), .A(n20520), .B(n20519), .ZN(
        P2_U3072) );
  AOI22_X1 U22623 ( .A1(n20523), .A2(n20542), .B1(n20530), .B2(n20522), .ZN(
        n20527) );
  AOI22_X1 U22624 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20525), .B1(
        n20524), .B2(n20544), .ZN(n20526) );
  OAI211_X1 U22625 ( .C1(n20539), .C2(n20528), .A(n20527), .B(n20526), .ZN(
        P2_U3064) );
  AOI22_X1 U22626 ( .A1(n20531), .A2(n20542), .B1(n20530), .B2(n20529), .ZN(
        n20535) );
  AOI22_X1 U22627 ( .A1(n20533), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n20532), .B2(n20544), .ZN(n20534) );
  OAI211_X1 U22628 ( .C1(n20539), .C2(n20536), .A(n20535), .B(n20534), .ZN(
        P2_U3056) );
  OAI22_X1 U22629 ( .A1(n20540), .A2(n20539), .B1(n20538), .B2(n20537), .ZN(
        n20541) );
  INV_X1 U22630 ( .A(n20541), .ZN(n20547) );
  AOI22_X1 U22631 ( .A1(n20545), .A2(n20544), .B1(n20543), .B2(n20542), .ZN(
        n20546) );
  OAI211_X1 U22632 ( .C1(n20548), .C2(n16492), .A(n20547), .B(n20546), .ZN(
        P2_U3048) );
  INV_X1 U22633 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20829) );
  INV_X1 U22634 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n20549) );
  AOI222_X1 U22635 ( .A1(n20828), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n20829), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n20549), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n20550) );
  INV_X1 U22636 ( .A(n20600), .ZN(n20602) );
  AOI22_X1 U22637 ( .A1(n20602), .A2(n20552), .B1(n20551), .B2(n20600), .ZN(
        U376) );
  OAI22_X1 U22638 ( .A1(n20600), .A2(P3_ADDRESS_REG_1__SCAN_IN), .B1(
        P2_ADDRESS_REG_1__SCAN_IN), .B2(n20602), .ZN(n20553) );
  INV_X1 U22639 ( .A(n20553), .ZN(U365) );
  OAI22_X1 U22640 ( .A1(n20600), .A2(P3_ADDRESS_REG_2__SCAN_IN), .B1(
        P2_ADDRESS_REG_2__SCAN_IN), .B2(n20602), .ZN(n20554) );
  INV_X1 U22641 ( .A(n20554), .ZN(U354) );
  OAI22_X1 U22642 ( .A1(n20600), .A2(P3_ADDRESS_REG_3__SCAN_IN), .B1(
        P2_ADDRESS_REG_3__SCAN_IN), .B2(n20602), .ZN(n20555) );
  INV_X1 U22643 ( .A(n20555), .ZN(U353) );
  OAI22_X1 U22644 ( .A1(n20600), .A2(P3_ADDRESS_REG_4__SCAN_IN), .B1(
        P2_ADDRESS_REG_4__SCAN_IN), .B2(n20602), .ZN(n20556) );
  INV_X1 U22645 ( .A(n20556), .ZN(U352) );
  INV_X1 U22646 ( .A(n20600), .ZN(n20599) );
  AOI22_X1 U22647 ( .A1(n20599), .A2(n20558), .B1(n20557), .B2(n20600), .ZN(
        U351) );
  AOI22_X1 U22648 ( .A1(n20599), .A2(n20560), .B1(n20559), .B2(n20600), .ZN(
        U350) );
  AOI22_X1 U22649 ( .A1(n20599), .A2(n20562), .B1(n20561), .B2(n20600), .ZN(
        U349) );
  AOI22_X1 U22650 ( .A1(n20599), .A2(n20564), .B1(n20563), .B2(n20600), .ZN(
        U348) );
  AOI22_X1 U22651 ( .A1(n20599), .A2(n20566), .B1(n20565), .B2(n20600), .ZN(
        U347) );
  AOI22_X1 U22652 ( .A1(n20599), .A2(n20568), .B1(n20567), .B2(n20600), .ZN(
        U375) );
  AOI22_X1 U22653 ( .A1(n20599), .A2(n20570), .B1(n20569), .B2(n20600), .ZN(
        U374) );
  AOI22_X1 U22654 ( .A1(n20599), .A2(n20572), .B1(n20571), .B2(n20600), .ZN(
        U373) );
  OAI22_X1 U22655 ( .A1(n20600), .A2(P3_ADDRESS_REG_13__SCAN_IN), .B1(
        P2_ADDRESS_REG_13__SCAN_IN), .B2(n20599), .ZN(n20573) );
  INV_X1 U22656 ( .A(n20573), .ZN(U372) );
  OAI22_X1 U22657 ( .A1(n20600), .A2(P3_ADDRESS_REG_14__SCAN_IN), .B1(
        P2_ADDRESS_REG_14__SCAN_IN), .B2(n20599), .ZN(n20574) );
  INV_X1 U22658 ( .A(n20574), .ZN(U371) );
  AOI22_X1 U22659 ( .A1(n20599), .A2(n20576), .B1(n20575), .B2(n20600), .ZN(
        U370) );
  AOI22_X1 U22660 ( .A1(n20599), .A2(n20578), .B1(n20577), .B2(n20600), .ZN(
        U369) );
  AOI22_X1 U22661 ( .A1(n20599), .A2(n20580), .B1(n20579), .B2(n20600), .ZN(
        U368) );
  AOI22_X1 U22662 ( .A1(n20599), .A2(n20582), .B1(n20581), .B2(n20600), .ZN(
        U367) );
  AOI22_X1 U22663 ( .A1(n20599), .A2(n20584), .B1(n20583), .B2(n20600), .ZN(
        U366) );
  OAI22_X1 U22664 ( .A1(n20600), .A2(P3_ADDRESS_REG_20__SCAN_IN), .B1(
        P2_ADDRESS_REG_20__SCAN_IN), .B2(n20599), .ZN(n20585) );
  INV_X1 U22665 ( .A(n20585), .ZN(U364) );
  OAI22_X1 U22666 ( .A1(n20600), .A2(P3_ADDRESS_REG_21__SCAN_IN), .B1(
        P2_ADDRESS_REG_21__SCAN_IN), .B2(n20599), .ZN(n20586) );
  INV_X1 U22667 ( .A(n20586), .ZN(U363) );
  AOI22_X1 U22668 ( .A1(n20599), .A2(n20588), .B1(n20587), .B2(n20600), .ZN(
        U362) );
  AOI22_X1 U22669 ( .A1(n20599), .A2(n20590), .B1(n20589), .B2(n20600), .ZN(
        U361) );
  AOI22_X1 U22670 ( .A1(n20602), .A2(n20592), .B1(n20591), .B2(n20600), .ZN(
        U360) );
  AOI22_X1 U22671 ( .A1(n20599), .A2(n20594), .B1(n20593), .B2(n20600), .ZN(
        U359) );
  AOI22_X1 U22672 ( .A1(n20599), .A2(n20596), .B1(n20595), .B2(n20600), .ZN(
        U358) );
  AOI22_X1 U22673 ( .A1(n20599), .A2(n20598), .B1(n20597), .B2(n20600), .ZN(
        U357) );
  OAI22_X1 U22674 ( .A1(n20600), .A2(P3_ADDRESS_REG_28__SCAN_IN), .B1(
        P2_ADDRESS_REG_28__SCAN_IN), .B2(n20602), .ZN(n20601) );
  INV_X1 U22675 ( .A(n20601), .ZN(U356) );
  OAI22_X1 U22676 ( .A1(n20600), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n20602), .ZN(n20603) );
  INV_X1 U22677 ( .A(n20603), .ZN(U355) );
  AOI22_X1 U22678 ( .A1(n20633), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20620), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20605) );
  OAI21_X1 U22679 ( .B1(n20606), .B2(n20635), .A(n20605), .ZN(P1_U2936) );
  AOI22_X1 U22680 ( .A1(n20633), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20620), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20607) );
  OAI21_X1 U22681 ( .B1(n20608), .B2(n20635), .A(n20607), .ZN(P1_U2935) );
  AOI22_X1 U22682 ( .A1(n20633), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20620), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20609) );
  OAI21_X1 U22683 ( .B1(n20610), .B2(n20635), .A(n20609), .ZN(P1_U2934) );
  AOI22_X1 U22684 ( .A1(n20633), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20611) );
  OAI21_X1 U22685 ( .B1(n20612), .B2(n20635), .A(n20611), .ZN(P1_U2933) );
  AOI22_X1 U22686 ( .A1(n20633), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20620), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20613) );
  OAI21_X1 U22687 ( .B1(n20614), .B2(n20635), .A(n20613), .ZN(P1_U2932) );
  AOI22_X1 U22688 ( .A1(n20633), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20615) );
  OAI21_X1 U22689 ( .B1(n14984), .B2(n20635), .A(n20615), .ZN(P1_U2931) );
  AOI22_X1 U22690 ( .A1(n20633), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20620), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20616) );
  OAI21_X1 U22691 ( .B1(n15284), .B2(n20635), .A(n20616), .ZN(P1_U2930) );
  AOI22_X1 U22692 ( .A1(n20633), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20620), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20617) );
  OAI21_X1 U22693 ( .B1(n15314), .B2(n20635), .A(n20617), .ZN(P1_U2929) );
  AOI22_X1 U22694 ( .A1(n20633), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20620), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20618) );
  OAI21_X1 U22695 ( .B1(n20619), .B2(n20635), .A(n20618), .ZN(P1_U2928) );
  INV_X1 U22696 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20622) );
  AOI22_X1 U22697 ( .A1(n20633), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20620), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20621) );
  OAI21_X1 U22698 ( .B1(n20622), .B2(n20635), .A(n20621), .ZN(P1_U2927) );
  INV_X1 U22699 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20624) );
  AOI22_X1 U22700 ( .A1(n20633), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20623) );
  OAI21_X1 U22701 ( .B1(n20624), .B2(n20635), .A(n20623), .ZN(P1_U2926) );
  AOI22_X1 U22702 ( .A1(n20633), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20625) );
  OAI21_X1 U22703 ( .B1(n16041), .B2(n20635), .A(n20625), .ZN(P1_U2925) );
  INV_X1 U22704 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20627) );
  AOI22_X1 U22705 ( .A1(n20633), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20626) );
  OAI21_X1 U22706 ( .B1(n20627), .B2(n20635), .A(n20626), .ZN(P1_U2924) );
  INV_X1 U22707 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20629) );
  AOI22_X1 U22708 ( .A1(n20633), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20628) );
  OAI21_X1 U22709 ( .B1(n20629), .B2(n20635), .A(n20628), .ZN(P1_U2923) );
  INV_X1 U22710 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20631) );
  AOI22_X1 U22711 ( .A1(n20633), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20630) );
  OAI21_X1 U22712 ( .B1(n20631), .B2(n20635), .A(n20630), .ZN(P1_U2922) );
  AOI22_X1 U22713 ( .A1(n20633), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20632), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20634) );
  OAI21_X1 U22714 ( .B1(n14214), .B2(n20635), .A(n20634), .ZN(P1_U2921) );
  CLKBUF_X1 U22715 ( .A(n22803), .Z(n20692) );
  OR2_X1 U22716 ( .A1(n22329), .A2(n20692), .ZN(n20650) );
  INV_X1 U22717 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n22098) );
  OR2_X1 U22718 ( .A1(n22803), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20653) );
  OAI222_X1 U22719 ( .A1(n20650), .A2(n22098), .B1(n20636), .B2(n22805), .C1(
        n22099), .C2(n20653), .ZN(P1_U3197) );
  INV_X1 U22720 ( .A(n20650), .ZN(n20669) );
  INV_X1 U22721 ( .A(n20653), .ZN(n20668) );
  AOI222_X1 U22722 ( .A1(n20669), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n22803), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20668), .ZN(n20637) );
  INV_X1 U22723 ( .A(n20637), .ZN(P1_U3198) );
  AOI22_X1 U22724 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(n20692), .B1(
        P1_REIP_REG_4__SCAN_IN), .B2(n20668), .ZN(n20638) );
  OAI21_X1 U22725 ( .B1(n22090), .B2(n20650), .A(n20638), .ZN(P1_U3199) );
  AOI22_X1 U22726 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(n20692), .B1(
        P1_REIP_REG_4__SCAN_IN), .B2(n20669), .ZN(n20639) );
  OAI21_X1 U22727 ( .B1(n22136), .B2(n20653), .A(n20639), .ZN(P1_U3200) );
  AOI22_X1 U22728 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(n20692), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n20668), .ZN(n20640) );
  OAI21_X1 U22729 ( .B1(n22136), .B2(n20650), .A(n20640), .ZN(P1_U3201) );
  INV_X1 U22730 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n22155) );
  AOI22_X1 U22731 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20692), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(n20669), .ZN(n20641) );
  OAI21_X1 U22732 ( .B1(n22155), .B2(n20653), .A(n20641), .ZN(P1_U3202) );
  AOI222_X1 U22733 ( .A1(n20669), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n22803), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20668), .ZN(n20642) );
  INV_X1 U22734 ( .A(n20642), .ZN(P1_U3203) );
  AOI222_X1 U22735 ( .A1(n20669), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20692), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n20668), .ZN(n20643) );
  INV_X1 U22736 ( .A(n20643), .ZN(P1_U3204) );
  AOI222_X1 U22737 ( .A1(n20669), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n22803), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20668), .ZN(n20644) );
  INV_X1 U22738 ( .A(n20644), .ZN(P1_U3205) );
  AOI22_X1 U22739 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n20692), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n20668), .ZN(n20645) );
  OAI21_X1 U22740 ( .B1(n22067), .B2(n20650), .A(n20645), .ZN(P1_U3206) );
  AOI22_X1 U22741 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20692), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n20669), .ZN(n20646) );
  OAI21_X1 U22742 ( .B1(n22177), .B2(n20653), .A(n20646), .ZN(P1_U3207) );
  AOI222_X1 U22743 ( .A1(n20668), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20692), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20669), .ZN(n20647) );
  INV_X1 U22744 ( .A(n20647), .ZN(P1_U3208) );
  AOI222_X1 U22745 ( .A1(n20669), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n22803), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20668), .ZN(n20648) );
  INV_X1 U22746 ( .A(n20648), .ZN(P1_U3209) );
  AOI22_X1 U22747 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20692), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(n20668), .ZN(n20649) );
  OAI21_X1 U22748 ( .B1(n20651), .B2(n20650), .A(n20649), .ZN(P1_U3210) );
  AOI22_X1 U22749 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n20692), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(n20669), .ZN(n20652) );
  OAI21_X1 U22750 ( .B1(n22199), .B2(n20653), .A(n20652), .ZN(P1_U3211) );
  AOI222_X1 U22751 ( .A1(n20669), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n22803), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20668), .ZN(n20654) );
  INV_X1 U22752 ( .A(n20654), .ZN(P1_U3212) );
  AOI222_X1 U22753 ( .A1(n20669), .A2(P1_REIP_REG_17__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n22803), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n20668), .ZN(n20655) );
  INV_X1 U22754 ( .A(n20655), .ZN(P1_U3213) );
  AOI222_X1 U22755 ( .A1(n20668), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n22803), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n20669), .ZN(n20656) );
  INV_X1 U22756 ( .A(n20656), .ZN(P1_U3214) );
  AOI222_X1 U22757 ( .A1(n20669), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n22803), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n20668), .ZN(n20657) );
  INV_X1 U22758 ( .A(n20657), .ZN(P1_U3215) );
  AOI222_X1 U22759 ( .A1(n20668), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n22803), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n20669), .ZN(n20658) );
  INV_X1 U22760 ( .A(n20658), .ZN(P1_U3216) );
  AOI222_X1 U22761 ( .A1(n20669), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n22803), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20668), .ZN(n20659) );
  INV_X1 U22762 ( .A(n20659), .ZN(P1_U3217) );
  AOI222_X1 U22763 ( .A1(n20669), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n22803), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20668), .ZN(n20660) );
  INV_X1 U22764 ( .A(n20660), .ZN(P1_U3218) );
  AOI222_X1 U22765 ( .A1(n20669), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n22803), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20668), .ZN(n20661) );
  INV_X1 U22766 ( .A(n20661), .ZN(P1_U3219) );
  AOI222_X1 U22767 ( .A1(n20669), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n22803), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20668), .ZN(n20662) );
  INV_X1 U22768 ( .A(n20662), .ZN(P1_U3220) );
  AOI222_X1 U22769 ( .A1(n20669), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n22803), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20668), .ZN(n20663) );
  INV_X1 U22770 ( .A(n20663), .ZN(P1_U3221) );
  AOI222_X1 U22771 ( .A1(n20669), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n22803), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20668), .ZN(n20664) );
  INV_X1 U22772 ( .A(n20664), .ZN(P1_U3222) );
  AOI222_X1 U22773 ( .A1(n20669), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n22803), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20668), .ZN(n20665) );
  INV_X1 U22774 ( .A(n20665), .ZN(P1_U3223) );
  AOI222_X1 U22775 ( .A1(n20669), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n22803), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20668), .ZN(n20666) );
  INV_X1 U22776 ( .A(n20666), .ZN(P1_U3224) );
  AOI222_X1 U22777 ( .A1(n20669), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n22803), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n20668), .ZN(n20667) );
  INV_X1 U22778 ( .A(n20667), .ZN(P1_U3225) );
  AOI222_X1 U22779 ( .A1(n20669), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n22803), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20668), .ZN(n20670) );
  INV_X1 U22780 ( .A(n20670), .ZN(P1_U3226) );
  OAI22_X1 U22781 ( .A1(n22803), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n22805), .ZN(n20671) );
  INV_X1 U22782 ( .A(n20671), .ZN(P1_U3458) );
  NOR2_X1 U22783 ( .A1(P1_DATAWIDTH_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20672) );
  NAND2_X1 U22784 ( .A1(n20672), .A2(n20696), .ZN(n20691) );
  OAI21_X1 U22785 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(n20691), .ZN(n20683) );
  NOR4_X1 U22786 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20676) );
  NOR4_X1 U22787 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20675) );
  NOR4_X1 U22788 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20674) );
  NOR4_X1 U22789 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20673) );
  NAND4_X1 U22790 ( .A1(n20676), .A2(n20675), .A3(n20674), .A4(n20673), .ZN(
        n20682) );
  NOR4_X1 U22791 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20680) );
  AOI211_X1 U22792 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20679) );
  NOR4_X1 U22793 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20678) );
  NOR4_X1 U22794 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20677) );
  NAND4_X1 U22795 ( .A1(n20680), .A2(n20679), .A3(n20678), .A4(n20677), .ZN(
        n20681) );
  OR2_X1 U22796 ( .A1(n20682), .A2(n20681), .ZN(n20694) );
  MUX2_X1 U22797 ( .A(n20683), .B(P1_BYTEENABLE_REG_3__SCAN_IN), .S(n20694), 
        .Z(P1_U2808) );
  OAI22_X1 U22798 ( .A1(n20692), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n22805), .ZN(n20684) );
  INV_X1 U22799 ( .A(n20684), .ZN(P1_U3459) );
  NAND2_X1 U22800 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20688) );
  NOR2_X1 U22801 ( .A1(n20694), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20697) );
  INV_X1 U22802 ( .A(n20697), .ZN(n20685) );
  AOI211_X1 U22803 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(n20685), .B(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20686) );
  AOI21_X1 U22804 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(n20694), .A(n20686), 
        .ZN(n20687) );
  OAI21_X1 U22805 ( .B1(n20688), .B2(n20694), .A(n20687), .ZN(P1_U3481) );
  OAI22_X1 U22806 ( .A1(n20692), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n22805), .ZN(n20689) );
  INV_X1 U22807 ( .A(n20689), .ZN(P1_U3460) );
  AOI22_X1 U22808 ( .A1(n20697), .A2(n20691), .B1(n20690), .B2(n20694), .ZN(
        P1_U2807) );
  OAI22_X1 U22809 ( .A1(n20692), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n22805), .ZN(n20693) );
  INV_X1 U22810 ( .A(n20693), .ZN(P1_U3461) );
  INV_X1 U22811 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20695) );
  AOI22_X1 U22812 ( .A1(n20697), .A2(n20696), .B1(n20695), .B2(n20694), .ZN(
        P1_U3482) );
  XNOR2_X1 U22813 ( .A(n20699), .B(n20716), .ZN(n22130) );
  AOI22_X1 U22814 ( .A1(n22134), .A2(n20725), .B1(n20724), .B2(n22130), .ZN(
        n20700) );
  OAI21_X1 U22815 ( .B1(n20727), .B2(n20701), .A(n20700), .ZN(P1_U2866) );
  INV_X1 U22816 ( .A(n22172), .ZN(n20702) );
  AOI22_X1 U22817 ( .A1(n22168), .A2(n20725), .B1(n20724), .B2(n20702), .ZN(
        n20703) );
  OAI21_X1 U22818 ( .B1(n20727), .B2(n22171), .A(n20703), .ZN(P1_U2860) );
  INV_X1 U22819 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n20705) );
  AOI22_X1 U22820 ( .A1(n22163), .A2(n20725), .B1(n22157), .B2(n20724), .ZN(
        n20704) );
  OAI21_X1 U22821 ( .B1(n20727), .B2(n20705), .A(n20704), .ZN(P1_U2861) );
  INV_X1 U22822 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n22211) );
  AOI22_X1 U22823 ( .A1(n22218), .A2(n20725), .B1(n20724), .B2(n22216), .ZN(
        n20706) );
  OAI21_X1 U22824 ( .B1(n20727), .B2(n22211), .A(n20706), .ZN(P1_U2855) );
  INV_X1 U22825 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n22183) );
  INV_X1 U22826 ( .A(n20707), .ZN(n22188) );
  AOI22_X1 U22827 ( .A1(n22188), .A2(n20725), .B1(n20724), .B2(n22186), .ZN(
        n20708) );
  OAI21_X1 U22828 ( .B1(n20727), .B2(n22183), .A(n20708), .ZN(P1_U2857) );
  INV_X1 U22829 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n22246) );
  NOR2_X1 U22830 ( .A1(n22251), .A2(n16841), .ZN(n20709) );
  AOI21_X1 U22831 ( .B1(n22254), .B2(n20725), .A(n20709), .ZN(n20710) );
  OAI21_X1 U22832 ( .B1(n20727), .B2(n22246), .A(n20710), .ZN(P1_U2851) );
  AOI22_X1 U22833 ( .A1(n20712), .A2(n20725), .B1(n20724), .B2(n20711), .ZN(
        n20713) );
  OAI21_X1 U22834 ( .B1(n20727), .B2(n20714), .A(n20713), .ZN(P1_U2853) );
  INV_X1 U22835 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n22146) );
  INV_X1 U22836 ( .A(n20699), .ZN(n20717) );
  AOI21_X1 U22837 ( .B1(n20717), .B2(n20716), .A(n20715), .ZN(n20719) );
  OR2_X1 U22838 ( .A1(n20719), .A2(n20718), .ZN(n22144) );
  NOR2_X1 U22839 ( .A1(n22144), .A2(n16841), .ZN(n20720) );
  AOI21_X1 U22840 ( .B1(n22152), .B2(n20725), .A(n20720), .ZN(n20721) );
  OAI21_X1 U22841 ( .B1(n20727), .B2(n22146), .A(n20721), .ZN(P1_U2865) );
  INV_X1 U22842 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n22120) );
  NAND2_X1 U22843 ( .A1(n15328), .A2(n20722), .ZN(n20723) );
  AND2_X1 U22844 ( .A1(n20699), .A2(n20723), .ZN(n22123) );
  AOI22_X1 U22845 ( .A1(n22126), .A2(n20725), .B1(n20724), .B2(n22123), .ZN(
        n20726) );
  OAI21_X1 U22846 ( .B1(n20727), .B2(n22120), .A(n20726), .ZN(P1_U2867) );
  NAND2_X1 U22847 ( .A1(n20729), .A2(n20728), .ZN(n20732) );
  INV_X1 U22848 ( .A(n20730), .ZN(n20731) );
  AOI22_X1 U22849 ( .A1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20732), .B1(
        n20762), .B2(n20731), .ZN(n20734) );
  NAND2_X1 U22850 ( .A1(n22021), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20733) );
  OAI211_X1 U22851 ( .C1(n22277), .C2(n20735), .A(n20734), .B(n20733), .ZN(
        P1_U2999) );
  AOI22_X1 U22852 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n20760), .B1(
        n22021), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20739) );
  INV_X1 U22853 ( .A(n20736), .ZN(n22112) );
  AOI22_X1 U22854 ( .A1(n20737), .A2(n20756), .B1(n20762), .B2(n22112), .ZN(
        n20738) );
  OAI211_X1 U22855 ( .C1(n20759), .C2(n22118), .A(n20739), .B(n20738), .ZN(
        P1_U2995) );
  AOI22_X1 U22856 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20760), .B1(
        n22021), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n20745) );
  OAI21_X1 U22857 ( .B1(n20742), .B2(n20741), .A(n20740), .ZN(n20743) );
  INV_X1 U22858 ( .A(n20743), .ZN(n22023) );
  AOI22_X1 U22859 ( .A1(n22023), .A2(n20756), .B1(n20762), .B2(n22126), .ZN(
        n20744) );
  OAI211_X1 U22860 ( .C1(n20759), .C2(n22129), .A(n20745), .B(n20744), .ZN(
        P1_U2994) );
  AOI22_X1 U22861 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20760), .B1(
        n22021), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n20751) );
  OAI21_X1 U22862 ( .B1(n20748), .B2(n20747), .A(n20746), .ZN(n20749) );
  INV_X1 U22863 ( .A(n20749), .ZN(n22016) );
  AOI22_X1 U22864 ( .A1(n22016), .A2(n20756), .B1(n20762), .B2(n22134), .ZN(
        n20750) );
  OAI211_X1 U22865 ( .C1(n20759), .C2(n22141), .A(n20751), .B(n20750), .ZN(
        P1_U2993) );
  AOI22_X1 U22866 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n20760), .B1(
        n22021), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n20758) );
  OAI21_X1 U22867 ( .B1(n20754), .B2(n20753), .A(n20752), .ZN(n20755) );
  INV_X1 U22868 ( .A(n20755), .ZN(n22034) );
  AOI22_X1 U22869 ( .A1(n22034), .A2(n20756), .B1(n20762), .B2(n22152), .ZN(
        n20757) );
  OAI211_X1 U22870 ( .C1(n20759), .C2(n22142), .A(n20758), .B(n20757), .ZN(
        P1_U2992) );
  AOI22_X1 U22871 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n20760), .B1(
        n22021), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n20764) );
  AOI22_X1 U22872 ( .A1(n22218), .A2(n20762), .B1(n22215), .B2(n20761), .ZN(
        n20763) );
  OAI211_X1 U22873 ( .C1(n22277), .C2(n20765), .A(n20764), .B(n20763), .ZN(
        P1_U2982) );
  OAI21_X1 U22874 ( .B1(n20766), .B2(n22302), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20767) );
  OAI21_X1 U22875 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20768), .A(n20767), 
        .ZN(P1_U2803) );
  INV_X1 U22876 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n20770) );
  OAI21_X1 U22877 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n22329), .A(n22335), 
        .ZN(n20769) );
  AOI22_X1 U22878 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(n22805), .B1(n20770), 
        .B2(n20769), .ZN(P1_U2804) );
  AOI22_X1 U22879 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n20825), .ZN(n20772) );
  OAI21_X1 U22880 ( .B1(n14388), .B2(n20811), .A(n20772), .ZN(U247) );
  AOI22_X1 U22881 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n20825), .ZN(n20773) );
  OAI21_X1 U22882 ( .B1(n14533), .B2(n20811), .A(n20773), .ZN(U246) );
  AOI22_X1 U22883 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n20825), .ZN(n20774) );
  OAI21_X1 U22884 ( .B1(n14523), .B2(n20811), .A(n20774), .ZN(U245) );
  AOI22_X1 U22885 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n20825), .ZN(n20775) );
  OAI21_X1 U22886 ( .B1(n14528), .B2(n20811), .A(n20775), .ZN(U244) );
  AOI22_X1 U22887 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n20825), .ZN(n20776) );
  OAI21_X1 U22888 ( .B1(n14202), .B2(n20811), .A(n20776), .ZN(U243) );
  AOI22_X1 U22889 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n20825), .ZN(n20777) );
  OAI21_X1 U22890 ( .B1(n14220), .B2(n20811), .A(n20777), .ZN(U242) );
  AOI22_X1 U22891 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n20825), .ZN(n20778) );
  OAI21_X1 U22892 ( .B1(n14215), .B2(n20811), .A(n20778), .ZN(U241) );
  AOI22_X1 U22893 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n20825), .ZN(n20779) );
  OAI21_X1 U22894 ( .B1(n14235), .B2(n20811), .A(n20779), .ZN(U240) );
  INV_X1 U22895 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n20781) );
  AOI22_X1 U22896 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n20825), .ZN(n20780) );
  OAI21_X1 U22897 ( .B1(n20781), .B2(n20811), .A(n20780), .ZN(U239) );
  INV_X1 U22898 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n20783) );
  AOI22_X1 U22899 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n20825), .ZN(n20782) );
  OAI21_X1 U22900 ( .B1(n20783), .B2(n20811), .A(n20782), .ZN(U238) );
  INV_X1 U22901 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n20785) );
  AOI22_X1 U22902 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n20825), .ZN(n20784) );
  OAI21_X1 U22903 ( .B1(n20785), .B2(n20811), .A(n20784), .ZN(U237) );
  INV_X1 U22904 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n20787) );
  AOI22_X1 U22905 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n20825), .ZN(n20786) );
  OAI21_X1 U22906 ( .B1(n20787), .B2(n20811), .A(n20786), .ZN(U236) );
  INV_X1 U22907 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20789) );
  AOI22_X1 U22908 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n20825), .ZN(n20788) );
  OAI21_X1 U22909 ( .B1(n20789), .B2(n20811), .A(n20788), .ZN(U235) );
  INV_X1 U22910 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n20791) );
  AOI22_X1 U22911 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n20825), .ZN(n20790) );
  OAI21_X1 U22912 ( .B1(n20791), .B2(n20811), .A(n20790), .ZN(U234) );
  INV_X1 U22913 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n20793) );
  AOI22_X1 U22914 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n20825), .ZN(n20792) );
  OAI21_X1 U22915 ( .B1(n20793), .B2(n20811), .A(n20792), .ZN(U233) );
  INV_X1 U22916 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n20795) );
  AOI22_X1 U22917 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n20825), .ZN(n20794) );
  OAI21_X1 U22918 ( .B1(n20795), .B2(n20811), .A(n20794), .ZN(U232) );
  AOI22_X1 U22919 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n20825), .ZN(n20796) );
  OAI21_X1 U22920 ( .B1(n20797), .B2(n20811), .A(n20796), .ZN(U231) );
  AOI22_X1 U22921 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n20825), .ZN(n20798) );
  OAI21_X1 U22922 ( .B1(n20799), .B2(n20811), .A(n20798), .ZN(U230) );
  AOI22_X1 U22923 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n20825), .ZN(n20800) );
  OAI21_X1 U22924 ( .B1(n20801), .B2(n20811), .A(n20800), .ZN(U229) );
  AOI22_X1 U22925 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n20825), .ZN(n20802) );
  OAI21_X1 U22926 ( .B1(n20803), .B2(n20811), .A(n20802), .ZN(U228) );
  AOI22_X1 U22927 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n20825), .ZN(n20804) );
  OAI21_X1 U22928 ( .B1(n20805), .B2(n20811), .A(n20804), .ZN(U227) );
  AOI22_X1 U22929 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n20825), .ZN(n20806) );
  OAI21_X1 U22930 ( .B1(n20807), .B2(n20811), .A(n20806), .ZN(U226) );
  AOI22_X1 U22931 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n20825), .ZN(n20808) );
  OAI21_X1 U22932 ( .B1(n20809), .B2(n20811), .A(n20808), .ZN(U225) );
  INV_X1 U22933 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n22687) );
  AOI22_X1 U22934 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n20825), .ZN(n20810) );
  OAI21_X1 U22935 ( .B1(n22687), .B2(n20811), .A(n20810), .ZN(U224) );
  AOI22_X1 U22936 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n20825), .ZN(n20813) );
  OAI21_X1 U22937 ( .B1(n20814), .B2(n20811), .A(n20813), .ZN(U223) );
  AOI22_X1 U22938 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n20825), .ZN(n20815) );
  OAI21_X1 U22939 ( .B1(n20816), .B2(n20811), .A(n20815), .ZN(U222) );
  AOI22_X1 U22940 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n20825), .ZN(n20817) );
  OAI21_X1 U22941 ( .B1(n20818), .B2(n20811), .A(n20817), .ZN(U221) );
  AOI22_X1 U22942 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n20825), .ZN(n20819) );
  OAI21_X1 U22943 ( .B1(n20820), .B2(n20811), .A(n20819), .ZN(U220) );
  AOI22_X1 U22944 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n20825), .ZN(n20821) );
  OAI21_X1 U22945 ( .B1(n20822), .B2(n20811), .A(n20821), .ZN(U219) );
  AOI22_X1 U22946 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n20825), .ZN(n20823) );
  OAI21_X1 U22947 ( .B1(n20824), .B2(n20811), .A(n20823), .ZN(U218) );
  AOI22_X1 U22948 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n20812), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n20825), .ZN(n20826) );
  OAI21_X1 U22949 ( .B1(n20827), .B2(n20811), .A(n20826), .ZN(U217) );
  OAI222_X1 U22950 ( .A1(U214), .A2(n20829), .B1(n20811), .B2(n22680), .C1(
        U212), .C2(n20828), .ZN(U216) );
  AOI22_X1 U22951 ( .A1(n22805), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20830), 
        .B2(n22803), .ZN(P1_U3483) );
  OAI21_X1 U22952 ( .B1(n22367), .B2(n20831), .A(n20899), .ZN(n20832) );
  AOI21_X1 U22953 ( .B1(n20833), .B2(n21961), .A(n20832), .ZN(n20840) );
  AOI21_X1 U22954 ( .B1(n21337), .B2(n22315), .A(n20834), .ZN(n20836) );
  OAI211_X1 U22955 ( .C1(n20836), .C2(n20835), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n22363), .ZN(n20837) );
  AOI21_X1 U22956 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n20837), .A(n21952), 
        .ZN(n20839) );
  NAND2_X1 U22957 ( .A1(n20840), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20838) );
  OAI21_X1 U22958 ( .B1(n20840), .B2(n20839), .A(n20838), .ZN(P3_U3296) );
  NAND2_X1 U22959 ( .A1(n20841), .A2(n20842), .ZN(n20893) );
  NAND2_X1 U22960 ( .A1(n20842), .A2(n22363), .ZN(n21339) );
  AOI22_X1 U22961 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20891), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20860), .ZN(n20844) );
  OAI21_X1 U22962 ( .B1(n20845), .B2(n20893), .A(n20844), .ZN(P3_U2768) );
  AOI22_X1 U22963 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20891), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20860), .ZN(n20846) );
  OAI21_X1 U22964 ( .B1(n21416), .B2(n20893), .A(n20846), .ZN(P3_U2769) );
  AOI22_X1 U22965 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20891), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20860), .ZN(n20847) );
  OAI21_X1 U22966 ( .B1(n20848), .B2(n20893), .A(n20847), .ZN(P3_U2770) );
  AOI22_X1 U22967 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20891), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20860), .ZN(n20850) );
  OAI21_X1 U22968 ( .B1(n21425), .B2(n20889), .A(n20850), .ZN(P3_U2771) );
  AOI22_X1 U22969 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20891), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20860), .ZN(n20851) );
  OAI21_X1 U22970 ( .B1(n21417), .B2(n20889), .A(n20851), .ZN(P3_U2772) );
  AOI22_X1 U22971 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20891), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20860), .ZN(n20852) );
  OAI21_X1 U22972 ( .B1(n21415), .B2(n20889), .A(n20852), .ZN(P3_U2773) );
  AOI22_X1 U22973 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20891), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20860), .ZN(n20853) );
  OAI21_X1 U22974 ( .B1(n21441), .B2(n20889), .A(n20853), .ZN(P3_U2774) );
  AOI22_X1 U22975 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20891), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20860), .ZN(n20854) );
  OAI21_X1 U22976 ( .B1(n20855), .B2(n20889), .A(n20854), .ZN(P3_U2775) );
  AOI22_X1 U22977 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20891), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20860), .ZN(n20856) );
  OAI21_X1 U22978 ( .B1(n20857), .B2(n20889), .A(n20856), .ZN(P3_U2776) );
  AOI22_X1 U22979 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20891), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20860), .ZN(n20858) );
  OAI21_X1 U22980 ( .B1(n20859), .B2(n20889), .A(n20858), .ZN(P3_U2777) );
  AOI22_X1 U22981 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20891), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n20890), .ZN(n20861) );
  OAI21_X1 U22982 ( .B1(n21450), .B2(n20889), .A(n20861), .ZN(P3_U2778) );
  AOI22_X1 U22983 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20891), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n20890), .ZN(n20862) );
  OAI21_X1 U22984 ( .B1(n20863), .B2(n20889), .A(n20862), .ZN(P3_U2779) );
  AOI22_X1 U22985 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20891), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20890), .ZN(n20864) );
  OAI21_X1 U22986 ( .B1(n20865), .B2(n20889), .A(n20864), .ZN(P3_U2780) );
  AOI22_X1 U22987 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20878), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n20890), .ZN(n20866) );
  OAI21_X1 U22988 ( .B1(n21463), .B2(n20889), .A(n20866), .ZN(P3_U2781) );
  AOI22_X1 U22989 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20878), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n20890), .ZN(n20867) );
  OAI21_X1 U22990 ( .B1(n20868), .B2(n20889), .A(n20867), .ZN(P3_U2782) );
  AOI22_X1 U22991 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20878), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n20890), .ZN(n20869) );
  OAI21_X1 U22992 ( .B1(n21530), .B2(n20889), .A(n20869), .ZN(P3_U2783) );
  AOI22_X1 U22993 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20878), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20890), .ZN(n20870) );
  OAI21_X1 U22994 ( .B1(n21518), .B2(n20889), .A(n20870), .ZN(P3_U2784) );
  AOI22_X1 U22995 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20878), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n20890), .ZN(n20871) );
  OAI21_X1 U22996 ( .B1(n20872), .B2(n20889), .A(n20871), .ZN(P3_U2785) );
  AOI22_X1 U22997 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20878), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n20890), .ZN(n20873) );
  OAI21_X1 U22998 ( .B1(n20874), .B2(n20889), .A(n20873), .ZN(P3_U2786) );
  AOI22_X1 U22999 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20878), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n20890), .ZN(n20875) );
  OAI21_X1 U23000 ( .B1(n21370), .B2(n20889), .A(n20875), .ZN(P3_U2787) );
  AOI22_X1 U23001 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20878), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n20890), .ZN(n20876) );
  OAI21_X1 U23002 ( .B1(n21343), .B2(n20889), .A(n20876), .ZN(P3_U2788) );
  AOI22_X1 U23003 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20878), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n20890), .ZN(n20877) );
  OAI21_X1 U23004 ( .B1(n21371), .B2(n20889), .A(n20877), .ZN(P3_U2789) );
  AOI22_X1 U23005 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20878), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n20890), .ZN(n20879) );
  OAI21_X1 U23006 ( .B1(n21342), .B2(n20889), .A(n20879), .ZN(P3_U2790) );
  AOI22_X1 U23007 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20891), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n20890), .ZN(n20880) );
  OAI21_X1 U23008 ( .B1(n21509), .B2(n20889), .A(n20880), .ZN(P3_U2791) );
  AOI22_X1 U23009 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20891), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n20890), .ZN(n20881) );
  OAI21_X1 U23010 ( .B1(n21400), .B2(n20893), .A(n20881), .ZN(P3_U2792) );
  AOI22_X1 U23011 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20891), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n20890), .ZN(n20882) );
  OAI21_X1 U23012 ( .B1(n20883), .B2(n20889), .A(n20882), .ZN(P3_U2793) );
  AOI22_X1 U23013 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20891), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n20890), .ZN(n20884) );
  OAI21_X1 U23014 ( .B1(n21351), .B2(n20893), .A(n20884), .ZN(P3_U2794) );
  AOI22_X1 U23015 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20891), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n20890), .ZN(n20885) );
  OAI21_X1 U23016 ( .B1(n21350), .B2(n20889), .A(n20885), .ZN(P3_U2795) );
  AOI22_X1 U23017 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20891), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n20890), .ZN(n20886) );
  OAI21_X1 U23018 ( .B1(n20887), .B2(n20893), .A(n20886), .ZN(P3_U2796) );
  AOI22_X1 U23019 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20891), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n20890), .ZN(n20888) );
  OAI21_X1 U23020 ( .B1(n21501), .B2(n20889), .A(n20888), .ZN(P3_U2797) );
  AOI22_X1 U23021 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20891), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n20890), .ZN(n20892) );
  OAI21_X1 U23022 ( .B1(n21504), .B2(n20893), .A(n20892), .ZN(P3_U2798) );
  AND2_X1 U23023 ( .A1(n20895), .A2(n20894), .ZN(n21954) );
  NAND2_X1 U23024 ( .A1(n14030), .A2(n21311), .ZN(n20896) );
  INV_X1 U23025 ( .A(n20898), .ZN(n21538) );
  AOI22_X1 U23026 ( .A1(n21119), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n21538), 
        .B2(n21327), .ZN(n20913) );
  INV_X1 U23027 ( .A(n20906), .ZN(n20901) );
  NAND2_X1 U23028 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n20904), .ZN(n20900) );
  NAND3_X1 U23029 ( .A1(n20905), .A2(n20901), .A3(n20900), .ZN(n21303) );
  AOI21_X1 U23030 ( .B1(n21146), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n21311), .ZN(n21065) );
  AOI22_X1 U23031 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(n21331), .B1(n20902), .B2(
        n21065), .ZN(n20912) );
  NAND2_X1 U23032 ( .A1(n22363), .A2(n22315), .ZN(n20903) );
  NAND4_X1 U23033 ( .A1(n20905), .A2(P3_EBX_REG_31__SCAN_IN), .A3(n20904), 
        .A4(n20903), .ZN(n21287) );
  AOI22_X1 U23034 ( .A1(n21330), .A2(n20907), .B1(n21179), .B2(n20923), .ZN(
        n20911) );
  INV_X4 U23035 ( .A(n20908), .ZN(n21312) );
  NOR2_X1 U23036 ( .A1(n21312), .A2(n21311), .ZN(n20909) );
  OAI221_X1 U23037 ( .B1(n21301), .B2(n20909), .C1(n21301), .C2(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20910) );
  NAND4_X1 U23038 ( .A1(n20913), .A2(n20912), .A3(n20911), .A4(n20910), .ZN(
        P3_U2670) );
  INV_X1 U23039 ( .A(n20914), .ZN(n20915) );
  AOI22_X1 U23040 ( .A1(n21119), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n20915), 
        .B2(n21327), .ZN(n20931) );
  INV_X1 U23041 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n21164) );
  NAND2_X1 U23042 ( .A1(n21164), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n21133) );
  AOI21_X1 U23043 ( .B1(n21164), .B2(n20916), .A(n21312), .ZN(n20917) );
  INV_X1 U23044 ( .A(n20917), .ZN(n20936) );
  AOI211_X1 U23045 ( .C1(n20918), .C2(n21133), .A(n21311), .B(n20936), .ZN(
        n20922) );
  NAND2_X1 U23046 ( .A1(n21135), .A2(n21312), .ZN(n21097) );
  OAI22_X1 U23047 ( .A1(n20920), .A2(n21318), .B1(n20919), .B2(n21097), .ZN(
        n20921) );
  AOI211_X1 U23048 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n21331), .A(n20922), .B(
        n20921), .ZN(n20930) );
  NOR2_X1 U23049 ( .A1(n20924), .A2(n20923), .ZN(n20932) );
  AOI211_X1 U23050 ( .C1(n20924), .C2(n20923), .A(n21162), .B(n20932), .ZN(
        n20925) );
  INV_X1 U23051 ( .A(n20925), .ZN(n20929) );
  NAND2_X1 U23052 ( .A1(n20927), .A2(n20926), .ZN(n20934) );
  OAI211_X1 U23053 ( .C1(n20927), .C2(n20926), .A(n21330), .B(n20934), .ZN(
        n20928) );
  NAND4_X1 U23054 ( .A1(n20931), .A2(n20930), .A3(n20929), .A4(n20928), .ZN(
        P3_U2669) );
  NAND3_X1 U23055 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .A3(P3_REIP_REG_1__SCAN_IN), .ZN(n20959) );
  AOI21_X1 U23056 ( .B1(n21179), .B2(n20959), .A(n21119), .ZN(n20957) );
  AOI21_X1 U23057 ( .B1(n21179), .B2(n20932), .A(P3_REIP_REG_3__SCAN_IN), .ZN(
        n20942) );
  AOI22_X1 U23058 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n21301), .B1(
        n21331), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n20941) );
  OR2_X1 U23059 ( .A1(n11151), .A2(n20933), .ZN(n21556) );
  NOR2_X1 U23060 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n20934), .ZN(n20945) );
  AOI211_X1 U23061 ( .C1(P3_EBX_REG_3__SCAN_IN), .C2(n20934), .A(n20945), .B(
        n21287), .ZN(n20939) );
  OAI21_X1 U23062 ( .B1(n20937), .B2(n20936), .A(n21135), .ZN(n20935) );
  AOI21_X1 U23063 ( .B1(n20937), .B2(n20936), .A(n20935), .ZN(n20938) );
  AOI211_X1 U23064 ( .C1(n21327), .C2(n21556), .A(n20939), .B(n20938), .ZN(
        n20940) );
  OAI211_X1 U23065 ( .C1(n20957), .C2(n20942), .A(n20941), .B(n20940), .ZN(
        P3_U2668) );
  OAI21_X1 U23066 ( .B1(n20943), .B2(n21133), .A(n21146), .ZN(n20962) );
  NOR3_X1 U23067 ( .A1(n20947), .A2(n21311), .A3(n20962), .ZN(n20944) );
  AOI211_X1 U23068 ( .C1(n21331), .C2(P3_EBX_REG_4__SCAN_IN), .A(n11153), .B(
        n20944), .ZN(n20956) );
  INV_X1 U23069 ( .A(n20945), .ZN(n20946) );
  AOI21_X1 U23070 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n20946), .A(n21287), .ZN(
        n20954) );
  NOR3_X1 U23071 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n21162), .A3(n20959), .ZN(
        n20953) );
  OAI211_X1 U23072 ( .C1(n21312), .C2(n20951), .A(n20947), .B(n21065), .ZN(
        n20950) );
  OAI21_X1 U23073 ( .B1(n20948), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n21327), .ZN(n20949) );
  OAI211_X1 U23074 ( .C1(n21318), .C2(n20951), .A(n20950), .B(n20949), .ZN(
        n20952) );
  AOI211_X1 U23075 ( .C1(n20954), .C2(n20958), .A(n20953), .B(n20952), .ZN(
        n20955) );
  OAI211_X1 U23076 ( .C1(n20957), .C2(n20960), .A(n20956), .B(n20955), .ZN(
        P3_U2667) );
  INV_X1 U23077 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n20969) );
  AOI211_X1 U23078 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n20958), .A(n20974), .B(
        n21287), .ZN(n20967) );
  NOR2_X1 U23079 ( .A1(n20960), .A2(n20959), .ZN(n20961) );
  NAND2_X1 U23080 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n20961), .ZN(n20991) );
  AOI21_X1 U23081 ( .B1(n21179), .B2(n20991), .A(n21119), .ZN(n20988) );
  AOI21_X1 U23082 ( .B1(n21179), .B2(n20961), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n20965) );
  XNOR2_X1 U23083 ( .A(n20963), .B(n20962), .ZN(n20964) );
  OAI22_X1 U23084 ( .A1(n20988), .A2(n20965), .B1(n21311), .B2(n20964), .ZN(
        n20966) );
  AOI211_X1 U23085 ( .C1(n21301), .C2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n20967), .B(n20966), .ZN(n20968) );
  OAI211_X1 U23086 ( .C1(n21303), .C2(n20969), .A(n20968), .B(n14030), .ZN(
        P3_U2666) );
  NOR3_X1 U23087 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n21162), .A3(n20991), .ZN(
        n20990) );
  NAND2_X1 U23088 ( .A1(n21135), .A2(n21164), .ZN(n21013) );
  OAI21_X1 U23089 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n21013), .A(
        n21097), .ZN(n20972) );
  INV_X1 U23090 ( .A(n21133), .ZN(n21121) );
  NAND2_X1 U23091 ( .A1(n20970), .A2(n21121), .ZN(n21040) );
  NAND2_X1 U23092 ( .A1(n21146), .A2(n21040), .ZN(n20980) );
  NOR3_X1 U23093 ( .A1(n20973), .A2(n21311), .A3(n20980), .ZN(n20971) );
  AOI211_X1 U23094 ( .C1(n20973), .C2(n20972), .A(n11153), .B(n20971), .ZN(
        n20976) );
  NAND2_X1 U23095 ( .A1(n20974), .A2(n20977), .ZN(n20982) );
  OAI211_X1 U23096 ( .C1(n20974), .C2(n20977), .A(n21330), .B(n20982), .ZN(
        n20975) );
  OAI211_X1 U23097 ( .C1(n20977), .C2(n21303), .A(n20976), .B(n20975), .ZN(
        n20978) );
  AOI211_X1 U23098 ( .C1(n21301), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n20990), .B(n20978), .ZN(n20979) );
  OAI21_X1 U23099 ( .B1(n20988), .B2(n20992), .A(n20979), .ZN(P3_U2665) );
  XOR2_X1 U23100 ( .A(n20981), .B(n20980), .Z(n20987) );
  AOI211_X1 U23101 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n20982), .A(n21004), .B(
        n21287), .ZN(n20986) );
  INV_X1 U23102 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n20983) );
  OAI22_X1 U23103 ( .A1(n20984), .A2(n21318), .B1(n21303), .B2(n20983), .ZN(
        n20985) );
  AOI211_X1 U23104 ( .C1(n21135), .C2(n20987), .A(n20986), .B(n20985), .ZN(
        n20996) );
  INV_X1 U23105 ( .A(n20988), .ZN(n20989) );
  OAI21_X1 U23106 ( .B1(n20990), .B2(n20989), .A(P3_REIP_REG_7__SCAN_IN), .ZN(
        n20995) );
  NOR2_X1 U23107 ( .A1(n20992), .A2(n20991), .ZN(n20997) );
  NAND3_X1 U23108 ( .A1(n21179), .A2(n20997), .A3(n20993), .ZN(n20994) );
  NAND4_X1 U23109 ( .A1(n20996), .A2(n14030), .A3(n20995), .A4(n20994), .ZN(
        P3_U2664) );
  NAND2_X1 U23110 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n20997), .ZN(n20999) );
  NOR2_X1 U23111 ( .A1(n20998), .A2(n20999), .ZN(n21038) );
  OAI21_X1 U23112 ( .B1(n21038), .B2(n21162), .A(n21329), .ZN(n21010) );
  OAI21_X1 U23113 ( .B1(n21162), .B2(n20999), .A(n20998), .ZN(n21009) );
  OAI21_X1 U23114 ( .B1(n21000), .B2(n21133), .A(n21146), .ZN(n21002) );
  AOI21_X1 U23115 ( .B1(n21003), .B2(n21002), .A(n21311), .ZN(n21001) );
  OAI21_X1 U23116 ( .B1(n21003), .B2(n21002), .A(n21001), .ZN(n21006) );
  NAND2_X1 U23117 ( .A1(n21004), .A2(n21012), .ZN(n21019) );
  OAI211_X1 U23118 ( .C1(n21004), .C2(n21012), .A(n21330), .B(n21019), .ZN(
        n21005) );
  OAI211_X1 U23119 ( .C1(n21318), .C2(n21007), .A(n21006), .B(n21005), .ZN(
        n21008) );
  AOI21_X1 U23120 ( .B1(n21010), .B2(n21009), .A(n21008), .ZN(n21011) );
  OAI211_X1 U23121 ( .C1(n21303), .C2(n21012), .A(n21011), .B(n14030), .ZN(
        P3_U2663) );
  AOI22_X1 U23122 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n21301), .B1(
        n21331), .B2(P3_EBX_REG_9__SCAN_IN), .ZN(n21023) );
  OAI21_X1 U23123 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n21013), .A(
        n21097), .ZN(n21017) );
  AOI21_X1 U23124 ( .B1(n21164), .B2(n21014), .A(n21312), .ZN(n21015) );
  INV_X1 U23125 ( .A(n21015), .ZN(n21027) );
  NOR3_X1 U23126 ( .A1(n21018), .A2(n21311), .A3(n21027), .ZN(n21016) );
  AOI211_X1 U23127 ( .C1(n21018), .C2(n21017), .A(n11153), .B(n21016), .ZN(
        n21022) );
  OAI221_X1 U23128 ( .B1(n21162), .B2(P3_REIP_REG_9__SCAN_IN), .C1(n21162), 
        .C2(n21038), .A(n21329), .ZN(n21032) );
  NAND2_X1 U23129 ( .A1(n21179), .A2(n21038), .ZN(n21024) );
  INV_X1 U23130 ( .A(n21024), .ZN(n21050) );
  AOI211_X1 U23131 ( .C1(P3_EBX_REG_9__SCAN_IN), .C2(n21019), .A(n21034), .B(
        n21287), .ZN(n21020) );
  AOI221_X1 U23132 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n21032), .C1(n21050), 
        .C2(n21032), .A(n21020), .ZN(n21021) );
  NAND3_X1 U23133 ( .A1(n21023), .A2(n21022), .A3(n21021), .ZN(P3_U2662) );
  INV_X1 U23134 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n21037) );
  NOR2_X1 U23135 ( .A1(n21025), .A2(n21024), .ZN(n21039) );
  AOI21_X1 U23136 ( .B1(n21028), .B2(n21027), .A(n21311), .ZN(n21026) );
  OAI21_X1 U23137 ( .B1(n21028), .B2(n21027), .A(n21026), .ZN(n21029) );
  OAI211_X1 U23138 ( .C1(n21030), .C2(n21318), .A(n14030), .B(n21029), .ZN(
        n21031) );
  AOI221_X1 U23139 ( .B1(n21039), .B2(n21033), .C1(n21032), .C2(
        P3_REIP_REG_10__SCAN_IN), .A(n21031), .ZN(n21036) );
  NAND2_X1 U23140 ( .A1(n21034), .A2(n21037), .ZN(n21044) );
  OAI211_X1 U23141 ( .C1(n21034), .C2(n21037), .A(n21330), .B(n21044), .ZN(
        n21035) );
  OAI211_X1 U23142 ( .C1(n21037), .C2(n21303), .A(n21036), .B(n21035), .ZN(
        P3_U2661) );
  NAND4_X1 U23143 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(P3_REIP_REG_10__SCAN_IN), 
        .A3(P3_REIP_REG_11__SCAN_IN), .A4(n21038), .ZN(n21081) );
  AOI21_X1 U23144 ( .B1(n21179), .B2(n21081), .A(n21119), .ZN(n21069) );
  AOI21_X1 U23145 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n21039), .A(
        P3_REIP_REG_11__SCAN_IN), .ZN(n21049) );
  AOI22_X1 U23146 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n21301), .B1(
        n21331), .B2(P3_EBX_REG_11__SCAN_IN), .ZN(n21048) );
  OAI21_X1 U23147 ( .B1(n21041), .B2(n21040), .A(n21146), .ZN(n21042) );
  XOR2_X1 U23148 ( .A(n21043), .B(n21042), .Z(n21046) );
  AOI211_X1 U23149 ( .C1(P3_EBX_REG_11__SCAN_IN), .C2(n21044), .A(n21051), .B(
        n21287), .ZN(n21045) );
  AOI211_X1 U23150 ( .C1(n21135), .C2(n21046), .A(n11153), .B(n21045), .ZN(
        n21047) );
  OAI211_X1 U23151 ( .C1(n21069), .C2(n21049), .A(n21048), .B(n21047), .ZN(
        P3_U2660) );
  NAND4_X1 U23152 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(P3_REIP_REG_10__SCAN_IN), 
        .A3(P3_REIP_REG_11__SCAN_IN), .A4(n21050), .ZN(n21083) );
  NAND2_X1 U23153 ( .A1(n21051), .A2(n21058), .ZN(n21063) );
  OAI211_X1 U23154 ( .C1(n21058), .C2(n21051), .A(n21063), .B(n21330), .ZN(
        n21052) );
  INV_X1 U23155 ( .A(n21052), .ZN(n21060) );
  AOI21_X1 U23156 ( .B1(n21164), .B2(n21053), .A(n21312), .ZN(n21055) );
  INV_X1 U23157 ( .A(n21056), .ZN(n21054) );
  INV_X1 U23158 ( .A(n21055), .ZN(n21073) );
  OAI221_X1 U23159 ( .B1(n21056), .B2(n21055), .C1(n21054), .C2(n21073), .A(
        n21135), .ZN(n21057) );
  OAI211_X1 U23160 ( .C1(n21303), .C2(n21058), .A(n14030), .B(n21057), .ZN(
        n21059) );
  AOI211_X1 U23161 ( .C1(n21301), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n21060), .B(n21059), .ZN(n21061) );
  OAI221_X1 U23162 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n21083), .C1(n21062), 
        .C2(n21069), .A(n21061), .ZN(P3_U2659) );
  AOI211_X1 U23163 ( .C1(P3_EBX_REG_13__SCAN_IN), .C2(n21063), .A(n21088), .B(
        n21287), .ZN(n21064) );
  AOI211_X1 U23164 ( .C1(n21331), .C2(P3_EBX_REG_13__SCAN_IN), .A(n11153), .B(
        n21064), .ZN(n21078) );
  INV_X1 U23165 ( .A(n21065), .ZN(n21066) );
  AOI211_X1 U23166 ( .C1(n21067), .C2(n21097), .A(n21066), .B(n21075), .ZN(
        n21072) );
  XNOR2_X1 U23167 ( .A(P3_REIP_REG_13__SCAN_IN), .B(P3_REIP_REG_12__SCAN_IN), 
        .ZN(n21070) );
  OAI22_X1 U23168 ( .A1(n21083), .A2(n21070), .B1(n21069), .B2(n21068), .ZN(
        n21071) );
  AOI211_X1 U23169 ( .C1(n21301), .C2(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n21072), .B(n21071), .ZN(n21077) );
  OAI21_X1 U23170 ( .B1(n21074), .B2(n21312), .A(n21073), .ZN(n21079) );
  NAND3_X1 U23171 ( .A1(n21135), .A2(n21075), .A3(n21079), .ZN(n21076) );
  NAND3_X1 U23172 ( .A1(n21078), .A2(n21077), .A3(n21076), .ZN(P3_U2658) );
  AOI22_X1 U23173 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n21301), .B1(
        n21331), .B2(P3_EBX_REG_14__SCAN_IN), .ZN(n21091) );
  XOR2_X1 U23174 ( .A(n21080), .B(n21079), .Z(n21086) );
  NAND2_X1 U23175 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(P3_REIP_REG_12__SCAN_IN), 
        .ZN(n21084) );
  NOR3_X1 U23176 ( .A1(n21082), .A2(n21081), .A3(n21084), .ZN(n21107) );
  OAI21_X1 U23177 ( .B1(n21107), .B2(n21162), .A(n21329), .ZN(n21115) );
  OAI21_X1 U23178 ( .B1(n21084), .B2(n21083), .A(n21082), .ZN(n21085) );
  AOI22_X1 U23179 ( .A1(n21135), .A2(n21086), .B1(n21115), .B2(n21085), .ZN(
        n21090) );
  NAND2_X1 U23180 ( .A1(n21088), .A2(n21087), .ZN(n21092) );
  OAI211_X1 U23181 ( .C1(n21088), .C2(n21087), .A(n21330), .B(n21092), .ZN(
        n21089) );
  NAND4_X1 U23182 ( .A1(n21091), .A2(n21090), .A3(n14030), .A4(n21089), .ZN(
        P3_U2657) );
  NOR2_X1 U23183 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n21092), .ZN(n21109) );
  AOI211_X1 U23184 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n21092), .A(n21109), .B(
        n21287), .ZN(n21093) );
  AOI21_X1 U23185 ( .B1(n21301), .B2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n21093), .ZN(n21104) );
  AND2_X1 U23186 ( .A1(n21094), .A2(n21164), .ZN(n21095) );
  AOI21_X1 U23187 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n21095), .A(
        n21312), .ZN(n21105) );
  INV_X1 U23188 ( .A(n21105), .ZN(n21098) );
  OAI21_X1 U23189 ( .B1(n21095), .B2(n21099), .A(n21135), .ZN(n21096) );
  AOI22_X1 U23190 ( .A1(n21099), .A2(n21098), .B1(n21097), .B2(n21096), .ZN(
        n21100) );
  AOI211_X1 U23191 ( .C1(n21331), .C2(P3_EBX_REG_15__SCAN_IN), .A(n11153), .B(
        n21100), .ZN(n21103) );
  INV_X1 U23192 ( .A(n21107), .ZN(n21101) );
  NOR3_X1 U23193 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n21162), .A3(n21101), 
        .ZN(n21114) );
  AOI21_X1 U23194 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n21115), .A(n21114), 
        .ZN(n21102) );
  NAND3_X1 U23195 ( .A1(n21104), .A2(n21103), .A3(n21102), .ZN(P3_U2656) );
  XOR2_X1 U23196 ( .A(n21106), .B(n21105), .Z(n21117) );
  NAND2_X1 U23197 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n21107), .ZN(n21118) );
  NAND2_X1 U23198 ( .A1(n21179), .A2(n21906), .ZN(n21112) );
  AOI22_X1 U23199 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n21301), .B1(
        n21331), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n21111) );
  NAND2_X1 U23200 ( .A1(n21109), .A2(n21108), .ZN(n21120) );
  OAI211_X1 U23201 ( .C1(n21109), .C2(n21108), .A(n21330), .B(n21120), .ZN(
        n21110) );
  OAI211_X1 U23202 ( .C1(n21118), .C2(n21112), .A(n21111), .B(n21110), .ZN(
        n21113) );
  AOI221_X1 U23203 ( .B1(n21115), .B2(P3_REIP_REG_16__SCAN_IN), .C1(n21114), 
        .C2(P3_REIP_REG_16__SCAN_IN), .A(n21113), .ZN(n21116) );
  OAI211_X1 U23204 ( .C1(n21117), .C2(n21311), .A(n21116), .B(n14030), .ZN(
        P3_U2655) );
  NOR2_X1 U23205 ( .A1(n21906), .A2(n21118), .ZN(n21126) );
  NAND2_X1 U23206 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n21126), .ZN(n21151) );
  AOI21_X1 U23207 ( .B1(n21179), .B2(n21151), .A(n21119), .ZN(n21155) );
  NOR2_X1 U23208 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n21120), .ZN(n21142) );
  AOI211_X1 U23209 ( .C1(P3_EBX_REG_17__SCAN_IN), .C2(n21120), .A(n21142), .B(
        n21287), .ZN(n21131) );
  AOI21_X1 U23210 ( .B1(n21122), .B2(n21121), .A(n21312), .ZN(n21124) );
  XOR2_X1 U23211 ( .A(n21124), .B(n21123), .Z(n21127) );
  INV_X1 U23212 ( .A(n21151), .ZN(n21139) );
  NOR2_X1 U23213 ( .A1(n21139), .A2(n21162), .ZN(n21125) );
  AOI22_X1 U23214 ( .A1(n21135), .A2(n21127), .B1(n21126), .B2(n21125), .ZN(
        n21128) );
  OAI211_X1 U23215 ( .C1(n21303), .C2(n21129), .A(n21128), .B(n14030), .ZN(
        n21130) );
  AOI211_X1 U23216 ( .C1(n21301), .C2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n21131), .B(n21130), .ZN(n21132) );
  OAI21_X1 U23217 ( .B1(n21155), .B2(n21894), .A(n21132), .ZN(P3_U2654) );
  OAI21_X1 U23218 ( .B1(n21134), .B2(n21133), .A(n21146), .ZN(n21137) );
  OAI21_X1 U23219 ( .B1(n21138), .B2(n21137), .A(n21135), .ZN(n21136) );
  AOI21_X1 U23220 ( .B1(n21138), .B2(n21137), .A(n21136), .ZN(n21141) );
  NAND3_X1 U23221 ( .A1(n21179), .A2(n21139), .A3(n21888), .ZN(n21154) );
  OAI211_X1 U23222 ( .C1(n21155), .C2(n21888), .A(n14030), .B(n21154), .ZN(
        n21140) );
  AOI211_X1 U23223 ( .C1(n21301), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n21141), .B(n21140), .ZN(n21144) );
  NAND2_X1 U23224 ( .A1(n21142), .A2(n21145), .ZN(n21150) );
  OAI211_X1 U23225 ( .C1(n21142), .C2(n21145), .A(n21330), .B(n21150), .ZN(
        n21143) );
  OAI211_X1 U23226 ( .C1(n21145), .C2(n21303), .A(n21144), .B(n21143), .ZN(
        P3_U2653) );
  OAI21_X1 U23227 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n21147), .A(
        n21146), .ZN(n21148) );
  XOR2_X1 U23228 ( .A(n21149), .B(n21148), .Z(n21160) );
  NOR2_X1 U23229 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n21150), .ZN(n21173) );
  AOI211_X1 U23230 ( .C1(P3_EBX_REG_19__SCAN_IN), .C2(n21150), .A(n21173), .B(
        n21287), .ZN(n21158) );
  NOR2_X1 U23231 ( .A1(n21888), .A2(n21151), .ZN(n21161) );
  NOR2_X1 U23232 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n21162), .ZN(n21152) );
  AOI22_X1 U23233 ( .A1(n21331), .A2(P3_EBX_REG_19__SCAN_IN), .B1(n21161), 
        .B2(n21152), .ZN(n21153) );
  OAI221_X1 U23234 ( .B1(n21156), .B2(n21155), .C1(n21156), .C2(n21154), .A(
        n21153), .ZN(n21157) );
  AOI211_X1 U23235 ( .C1(n21301), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n21158), .B(n21157), .ZN(n21159) );
  OAI211_X1 U23236 ( .C1(n21160), .C2(n21311), .A(n21159), .B(n14030), .ZN(
        P3_U2652) );
  NAND2_X1 U23237 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n21161), .ZN(n21177) );
  NAND2_X1 U23238 ( .A1(n21179), .A2(n21163), .ZN(n21176) );
  NAND2_X1 U23239 ( .A1(n21329), .A2(n21162), .ZN(n21328) );
  NOR2_X1 U23240 ( .A1(n21163), .A2(n21177), .ZN(n21178) );
  NAND2_X1 U23241 ( .A1(n21178), .A2(n21329), .ZN(n21205) );
  NAND2_X1 U23242 ( .A1(n21328), .A2(n21205), .ZN(n21189) );
  INV_X1 U23243 ( .A(n21189), .ZN(n21197) );
  AND2_X1 U23244 ( .A1(n21165), .A2(n21164), .ZN(n21166) );
  AOI211_X1 U23245 ( .C1(n21168), .C2(n21167), .A(n21181), .B(n21311), .ZN(
        n21171) );
  OAI22_X1 U23246 ( .A1(n21169), .A2(n21318), .B1(n21303), .B2(n21172), .ZN(
        n21170) );
  AOI211_X1 U23247 ( .C1(n21197), .C2(P3_REIP_REG_20__SCAN_IN), .A(n21171), 
        .B(n21170), .ZN(n21175) );
  NAND2_X1 U23248 ( .A1(n21173), .A2(n21172), .ZN(n21180) );
  OAI211_X1 U23249 ( .C1(n21173), .C2(n21172), .A(n21330), .B(n21180), .ZN(
        n21174) );
  OAI211_X1 U23250 ( .C1(n21177), .C2(n21176), .A(n21175), .B(n21174), .ZN(
        P3_U2651) );
  AOI22_X1 U23251 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n21301), .B1(
        n21331), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n21188) );
  NOR2_X1 U23252 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n21180), .ZN(n21199) );
  AOI211_X1 U23253 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n21180), .A(n21199), .B(
        n21287), .ZN(n21186) );
  NOR2_X1 U23254 ( .A1(n21181), .A2(n21312), .ZN(n21183) );
  OR2_X2 U23255 ( .A1(n21183), .A2(n21184), .ZN(n21191) );
  INV_X1 U23256 ( .A(n21191), .ZN(n21182) );
  AOI211_X1 U23257 ( .C1(n21184), .C2(n21183), .A(n21182), .B(n21311), .ZN(
        n21185) );
  AOI211_X1 U23258 ( .C1(n21207), .C2(n21576), .A(n21186), .B(n21185), .ZN(
        n21187) );
  OAI211_X1 U23259 ( .C1(n21576), .C2(n21189), .A(n21188), .B(n21187), .ZN(
        P3_U2650) );
  INV_X1 U23260 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n21202) );
  INV_X1 U23261 ( .A(n21190), .ZN(n21193) );
  AND2_X2 U23262 ( .A1(n21191), .A2(n21146), .ZN(n21192) );
  AOI211_X1 U23263 ( .C1(n21193), .C2(n21192), .A(n21208), .B(n21311), .ZN(
        n21196) );
  NAND2_X1 U23264 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n21206) );
  OAI211_X1 U23265 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(P3_REIP_REG_21__SCAN_IN), .A(n21207), .B(n21206), .ZN(n21194) );
  OAI21_X1 U23266 ( .B1(n21198), .B2(n21303), .A(n21194), .ZN(n21195) );
  AOI211_X1 U23267 ( .C1(n21197), .C2(P3_REIP_REG_22__SCAN_IN), .A(n21196), 
        .B(n21195), .ZN(n21201) );
  NAND2_X1 U23268 ( .A1(n21199), .A2(n21198), .ZN(n21203) );
  OAI211_X1 U23269 ( .C1(n21199), .C2(n21198), .A(n21330), .B(n21203), .ZN(
        n21200) );
  OAI211_X1 U23270 ( .C1(n21318), .C2(n21202), .A(n21201), .B(n21200), .ZN(
        P3_U2649) );
  NOR2_X1 U23271 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n21203), .ZN(n21228) );
  AOI211_X1 U23272 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n21203), .A(n21228), .B(
        n21287), .ZN(n21204) );
  AOI21_X1 U23273 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n21331), .A(n21204), .ZN(
        n21217) );
  INV_X1 U23274 ( .A(n21328), .ZN(n21286) );
  NOR3_X1 U23275 ( .A1(n21839), .A2(n21206), .A3(n21205), .ZN(n21233) );
  NOR2_X1 U23276 ( .A1(n21286), .A2(n21233), .ZN(n21226) );
  NAND3_X1 U23277 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .A3(n21207), .ZN(n21219) );
  INV_X1 U23278 ( .A(n21219), .ZN(n21215) );
  NOR2_X1 U23279 ( .A1(n21208), .A2(n21312), .ZN(n21212) );
  INV_X1 U23280 ( .A(n21212), .ZN(n21210) );
  INV_X1 U23281 ( .A(n21213), .ZN(n21209) );
  NAND2_X1 U23282 ( .A1(n21210), .A2(n21209), .ZN(n21221) );
  INV_X1 U23283 ( .A(n21221), .ZN(n21211) );
  AOI211_X1 U23284 ( .C1(n21213), .C2(n21212), .A(n21211), .B(n21311), .ZN(
        n21214) );
  AOI221_X1 U23285 ( .B1(n21226), .B2(P3_REIP_REG_23__SCAN_IN), .C1(n21215), 
        .C2(n21839), .A(n21214), .ZN(n21216) );
  OAI211_X1 U23286 ( .C1(n21218), .C2(n21318), .A(n21217), .B(n21216), .ZN(
        P3_U2648) );
  AOI22_X1 U23287 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n21301), .B1(
        n21331), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n21231) );
  NOR2_X1 U23288 ( .A1(n21839), .A2(n21219), .ZN(n21232) );
  INV_X1 U23289 ( .A(n21220), .ZN(n21223) );
  NOR2_X1 U23290 ( .A1(n21223), .A2(n21222), .ZN(n21234) );
  AOI211_X1 U23291 ( .C1(n21223), .C2(n21222), .A(n21234), .B(n21311), .ZN(
        n21224) );
  AOI221_X1 U23292 ( .B1(n21226), .B2(P3_REIP_REG_24__SCAN_IN), .C1(n21232), 
        .C2(n21225), .A(n21224), .ZN(n21230) );
  INV_X1 U23293 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n21227) );
  NAND2_X1 U23294 ( .A1(n21228), .A2(n21227), .ZN(n21237) );
  OAI211_X1 U23295 ( .C1(n21228), .C2(n21227), .A(n21330), .B(n21237), .ZN(
        n21229) );
  NAND3_X1 U23296 ( .A1(n21231), .A2(n21230), .A3(n21229), .ZN(P3_U2647) );
  NAND2_X1 U23297 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n21232), .ZN(n21259) );
  NAND2_X1 U23298 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n21233), .ZN(n21245) );
  NAND2_X1 U23299 ( .A1(n21328), .A2(n21245), .ZN(n21244) );
  NOR2_X1 U23300 ( .A1(n21234), .A2(n21312), .ZN(n21235) );
  NOR2_X1 U23301 ( .A1(n21236), .A2(n21235), .ZN(n21248) );
  AOI211_X1 U23302 ( .C1(n21236), .C2(n21235), .A(n21248), .B(n21311), .ZN(
        n21242) );
  NOR2_X1 U23303 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n21237), .ZN(n21255) );
  AOI211_X1 U23304 ( .C1(P3_EBX_REG_25__SCAN_IN), .C2(n21237), .A(n21255), .B(
        n21287), .ZN(n21241) );
  OAI22_X1 U23305 ( .A1(n21239), .A2(n21318), .B1(n21303), .B2(n21238), .ZN(
        n21240) );
  NOR3_X1 U23306 ( .A1(n21242), .A2(n21241), .A3(n21240), .ZN(n21243) );
  OAI221_X1 U23307 ( .B1(P3_REIP_REG_25__SCAN_IN), .B2(n21259), .C1(n21261), 
        .C2(n21244), .A(n21243), .ZN(P3_U2646) );
  AOI22_X1 U23308 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n21301), .B1(
        n21331), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n21258) );
  NAND2_X1 U23309 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(P3_REIP_REG_26__SCAN_IN), 
        .ZN(n21246) );
  OAI21_X1 U23310 ( .B1(n21246), .B2(n21245), .A(n21328), .ZN(n21284) );
  INV_X1 U23311 ( .A(n21284), .ZN(n21253) );
  NOR2_X1 U23312 ( .A1(n21261), .A2(n21259), .ZN(n21252) );
  INV_X1 U23313 ( .A(n21247), .ZN(n21250) );
  NOR2_X1 U23314 ( .A1(n21248), .A2(n21312), .ZN(n21249) );
  NOR2_X1 U23315 ( .A1(n21250), .A2(n21249), .ZN(n21262) );
  AOI211_X1 U23316 ( .C1(n21250), .C2(n21249), .A(n21262), .B(n21311), .ZN(
        n21251) );
  AOI221_X1 U23317 ( .B1(n21253), .B2(P3_REIP_REG_26__SCAN_IN), .C1(n21252), 
        .C2(n21260), .A(n21251), .ZN(n21257) );
  NAND2_X1 U23318 ( .A1(n21255), .A2(n21254), .ZN(n21265) );
  OAI211_X1 U23319 ( .C1(n21255), .C2(n21254), .A(n21330), .B(n21265), .ZN(
        n21256) );
  NAND3_X1 U23320 ( .A1(n21258), .A2(n21257), .A3(n21256), .ZN(P3_U2645) );
  AOI22_X1 U23321 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n21301), .B1(
        n21331), .B2(P3_EBX_REG_27__SCAN_IN), .ZN(n21269) );
  NOR3_X1 U23322 ( .A1(n21261), .A2(n21260), .A3(n21259), .ZN(n21304) );
  NOR2_X1 U23323 ( .A1(n21262), .A2(n21312), .ZN(n21263) );
  NOR2_X1 U23324 ( .A1(n21264), .A2(n21263), .ZN(n21272) );
  AOI211_X1 U23325 ( .C1(n21264), .C2(n21263), .A(n21272), .B(n21311), .ZN(
        n21267) );
  NOR2_X1 U23326 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n21265), .ZN(n21279) );
  AOI211_X1 U23327 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n21265), .A(n21279), .B(
        n21287), .ZN(n21266) );
  AOI211_X1 U23328 ( .C1(n21304), .C2(n21270), .A(n21267), .B(n21266), .ZN(
        n21268) );
  OAI211_X1 U23329 ( .C1(n21270), .C2(n21284), .A(n21269), .B(n21268), .ZN(
        P3_U2644) );
  INV_X1 U23330 ( .A(n21271), .ZN(n21274) );
  NOR2_X1 U23331 ( .A1(n21272), .A2(n21312), .ZN(n21273) );
  NOR2_X1 U23332 ( .A1(n21274), .A2(n21273), .ZN(n21291) );
  AOI211_X1 U23333 ( .C1(n21274), .C2(n21273), .A(n21291), .B(n21311), .ZN(
        n21277) );
  INV_X1 U23334 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n21278) );
  OAI22_X1 U23335 ( .A1(n21275), .A2(n21284), .B1(n21303), .B2(n21278), .ZN(
        n21276) );
  AOI211_X1 U23336 ( .C1(n21301), .C2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n21277), .B(n21276), .ZN(n21282) );
  NAND2_X1 U23337 ( .A1(n21279), .A2(n21278), .ZN(n21288) );
  OAI211_X1 U23338 ( .C1(n21279), .C2(n21278), .A(n21330), .B(n21288), .ZN(
        n21281) );
  NAND2_X1 U23339 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n21290) );
  OAI211_X1 U23340 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n21304), .B(n21290), .ZN(n21280) );
  NAND3_X1 U23341 ( .A1(n21282), .A2(n21281), .A3(n21280), .ZN(P3_U2643) );
  NOR2_X1 U23342 ( .A1(n21283), .A2(n21290), .ZN(n21285) );
  OAI21_X1 U23343 ( .B1(n21286), .B2(n21285), .A(n21284), .ZN(n21322) );
  AOI22_X1 U23344 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n21322), .B1(n21331), 
        .B2(P3_EBX_REG_29__SCAN_IN), .ZN(n21298) );
  NOR2_X1 U23345 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n21288), .ZN(n21302) );
  NOR2_X1 U23346 ( .A1(n21302), .A2(n21287), .ZN(n21307) );
  NAND2_X1 U23347 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n21288), .ZN(n21296) );
  INV_X1 U23348 ( .A(n21304), .ZN(n21289) );
  NOR3_X1 U23349 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n21290), .A3(n21289), 
        .ZN(n21295) );
  NOR2_X1 U23350 ( .A1(n21291), .A2(n21312), .ZN(n21292) );
  NOR2_X1 U23351 ( .A1(n21293), .A2(n21292), .ZN(n21300) );
  AOI211_X1 U23352 ( .C1(n21293), .C2(n21292), .A(n21300), .B(n21311), .ZN(
        n21294) );
  AOI211_X1 U23353 ( .C1(n21307), .C2(n21296), .A(n21295), .B(n21294), .ZN(
        n21297) );
  OAI211_X1 U23354 ( .C1(n21299), .C2(n21318), .A(n21298), .B(n21297), .ZN(
        P3_U2642) );
  NOR2_X1 U23355 ( .A1(n21300), .A2(n21312), .ZN(n21313) );
  XNOR2_X1 U23356 ( .A(n21314), .B(n21313), .ZN(n21310) );
  AOI22_X1 U23357 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n21301), .B1(
        P3_REIP_REG_30__SCAN_IN), .B2(n21322), .ZN(n21309) );
  INV_X1 U23358 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n21306) );
  NAND2_X1 U23359 ( .A1(n21330), .A2(n21302), .ZN(n21326) );
  NAND2_X1 U23360 ( .A1(n21303), .A2(n21326), .ZN(n21305) );
  NAND4_X1 U23361 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n21304), .ZN(n21317) );
  NOR2_X1 U23362 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n21317), .ZN(n21323) );
  AOI221_X1 U23363 ( .B1(n21307), .B2(n21306), .C1(n21305), .C2(
        P3_EBX_REG_30__SCAN_IN), .A(n21323), .ZN(n21308) );
  OAI211_X1 U23364 ( .C1(n21311), .C2(n21310), .A(n21309), .B(n21308), .ZN(
        P3_U2641) );
  NOR4_X1 U23365 ( .A1(n21314), .A2(n21313), .A3(n21312), .A4(n21311), .ZN(
        n21321) );
  NAND2_X1 U23366 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n21315), .ZN(n21316) );
  OAI22_X1 U23367 ( .A1(n21319), .A2(n21318), .B1(n21317), .B2(n21316), .ZN(
        n21320) );
  OAI21_X1 U23368 ( .B1(n21323), .B2(n21322), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n21324) );
  OAI211_X1 U23369 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n21326), .A(n21325), .B(
        n21324), .ZN(P3_U2640) );
  AOI22_X1 U23370 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n21328), .B1(n21327), 
        .B2(n21535), .ZN(n21334) );
  NAND3_X1 U23371 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n21329), .A3(
        n21545), .ZN(n21333) );
  OAI21_X1 U23372 ( .B1(n21331), .B2(n21330), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n21332) );
  NAND3_X1 U23373 ( .A1(n21334), .A2(n21333), .A3(n21332), .ZN(P3_U2671) );
  NAND2_X1 U23374 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .ZN(n21401) );
  NAND3_X1 U23375 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .A3(P3_EAX_REG_2__SCAN_IN), .ZN(n21368) );
  NAND3_X1 U23376 ( .A1(n21337), .A2(n21336), .A3(n21335), .ZN(n21338) );
  NAND4_X1 U23377 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_4__SCAN_IN), .A4(n21529), .ZN(n21341) );
  INV_X1 U23378 ( .A(n21403), .ZN(n21511) );
  NOR3_X1 U23379 ( .A1(n21443), .A2(n21511), .A3(n21509), .ZN(n21363) );
  NAND2_X1 U23380 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n21366), .ZN(n21360) );
  NOR2_X1 U23381 ( .A1(n21401), .A2(n21360), .ZN(n21497) );
  INV_X1 U23382 ( .A(n21497), .ZN(n21349) );
  NAND3_X1 U23383 ( .A1(n21512), .A2(P3_EAX_REG_13__SCAN_IN), .A3(n21349), 
        .ZN(n21348) );
  INV_X1 U23384 ( .A(n21529), .ZN(n21369) );
  NOR2_X1 U23385 ( .A1(n21345), .A2(n21369), .ZN(n21526) );
  AOI22_X1 U23386 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21527), .B1(n21526), .B2(
        n21346), .ZN(n21347) );
  OAI211_X1 U23387 ( .C1(P3_EAX_REG_13__SCAN_IN), .C2(n21349), .A(n21348), .B(
        n21347), .ZN(P3_U2722) );
  INV_X1 U23388 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n21355) );
  OAI22_X1 U23389 ( .A1(n21360), .A2(n21351), .B1(n21350), .B2(n21461), .ZN(
        n21352) );
  INV_X1 U23390 ( .A(n21352), .ZN(n21354) );
  OAI222_X1 U23391 ( .A1(n21394), .A2(n21355), .B1(n21497), .B2(n21354), .C1(
        n21522), .C2(n21353), .ZN(P3_U2723) );
  NAND3_X1 U23392 ( .A1(n21512), .A2(P3_EAX_REG_11__SCAN_IN), .A3(n21360), 
        .ZN(n21358) );
  AOI22_X1 U23393 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n21527), .B1(n21526), .B2(
        n21356), .ZN(n21357) );
  OAI211_X1 U23394 ( .C1(P3_EAX_REG_11__SCAN_IN), .C2(n21360), .A(n21358), .B(
        n21357), .ZN(P3_U2724) );
  AOI22_X1 U23395 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n21527), .B1(n21526), .B2(
        n21359), .ZN(n21362) );
  OAI211_X1 U23396 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n21366), .A(n21512), .B(
        n21360), .ZN(n21361) );
  NAND2_X1 U23397 ( .A1(n21362), .A2(n21361), .ZN(P3_U2725) );
  INV_X1 U23398 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n21367) );
  AOI21_X1 U23399 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n21519), .A(n21363), .ZN(
        n21365) );
  OAI222_X1 U23400 ( .A1(n21394), .A2(n21367), .B1(n21366), .B2(n21365), .C1(
        n21522), .C2(n21364), .ZN(P3_U2726) );
  NOR2_X1 U23401 ( .A1(n21443), .A2(n21511), .ZN(n21510) );
  NOR3_X1 U23402 ( .A1(n21369), .A2(n21443), .A3(n21368), .ZN(n21399) );
  NAND2_X1 U23403 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n21399), .ZN(n21385) );
  NOR2_X1 U23404 ( .A1(n21370), .A2(n21385), .ZN(n21389) );
  NAND2_X1 U23405 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n21389), .ZN(n21375) );
  NOR2_X1 U23406 ( .A1(n21371), .A2(n21375), .ZN(n21379) );
  AOI21_X1 U23407 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n21512), .A(n21379), .ZN(
        n21373) );
  OAI222_X1 U23408 ( .A1(n21394), .A2(n21374), .B1(n21510), .B2(n21373), .C1(
        n21522), .C2(n11148), .ZN(P3_U2728) );
  INV_X1 U23409 ( .A(n21375), .ZN(n21383) );
  AOI21_X1 U23410 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n21512), .A(n21383), .ZN(
        n21378) );
  INV_X1 U23411 ( .A(n21376), .ZN(n21377) );
  OAI222_X1 U23412 ( .A1(n21380), .A2(n21394), .B1(n21379), .B2(n21378), .C1(
        n21522), .C2(n21377), .ZN(P3_U2729) );
  AOI21_X1 U23413 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n21512), .A(n21389), .ZN(
        n21382) );
  OAI222_X1 U23414 ( .A1(n21384), .A2(n21394), .B1(n21383), .B2(n21382), .C1(
        n21522), .C2(n21381), .ZN(P3_U2730) );
  INV_X1 U23415 ( .A(n21385), .ZN(n21393) );
  AOI21_X1 U23416 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n21512), .A(n21393), .ZN(
        n21388) );
  INV_X1 U23417 ( .A(n21386), .ZN(n21387) );
  OAI222_X1 U23418 ( .A1(n21390), .A2(n21394), .B1(n21389), .B2(n21388), .C1(
        n21522), .C2(n21387), .ZN(P3_U2731) );
  AOI21_X1 U23419 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n21519), .A(n21399), .ZN(
        n21392) );
  OAI222_X1 U23420 ( .A1(n21395), .A2(n21394), .B1(n21393), .B2(n21392), .C1(
        n21522), .C2(n21391), .ZN(P3_U2732) );
  NAND2_X1 U23421 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n21529), .ZN(n21517) );
  NOR2_X1 U23422 ( .A1(n21518), .A2(n21517), .ZN(n21516) );
  OAI21_X1 U23423 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n21516), .A(n21519), .ZN(
        n21398) );
  AOI22_X1 U23424 ( .A1(n21527), .A2(BUF2_REG_2__SCAN_IN), .B1(n21526), .B2(
        n21396), .ZN(n21397) );
  OAI21_X1 U23425 ( .B1(n21399), .B2(n21398), .A(n21397), .ZN(P3_U2733) );
  NAND2_X1 U23426 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .ZN(n21418) );
  NOR4_X1 U23427 ( .A1(n21509), .A2(n21501), .A3(n21401), .A4(n21400), .ZN(
        n21402) );
  NAND4_X1 U23428 ( .A1(n21403), .A2(P3_EAX_REG_10__SCAN_IN), .A3(
        P3_EAX_REG_13__SCAN_IN), .A4(n21402), .ZN(n21505) );
  NOR2_X1 U23429 ( .A1(n21443), .A2(n21493), .ZN(n21436) );
  NAND2_X1 U23430 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n21436), .ZN(n21435) );
  NOR2_X1 U23431 ( .A1(n21418), .A2(n21435), .ZN(n21424) );
  NAND2_X1 U23432 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n21424), .ZN(n21411) );
  NAND3_X1 U23433 ( .A1(n21512), .A2(P3_EAX_REG_21__SCAN_IN), .A3(n21411), 
        .ZN(n21410) );
  NOR2_X2 U23434 ( .A1(n21404), .A2(n21519), .ZN(n21491) );
  INV_X1 U23435 ( .A(n21492), .ZN(n21485) );
  OAI22_X1 U23436 ( .A1(n21407), .A2(n21522), .B1(n21406), .B2(n21485), .ZN(
        n21408) );
  AOI21_X1 U23437 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n21491), .A(n21408), .ZN(
        n21409) );
  OAI211_X1 U23438 ( .C1(P3_EAX_REG_21__SCAN_IN), .C2(n21411), .A(n21410), .B(
        n21409), .ZN(P3_U2714) );
  AOI22_X1 U23439 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n21492), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n21491), .ZN(n21413) );
  OAI211_X1 U23440 ( .C1(n21424), .C2(P3_EAX_REG_20__SCAN_IN), .A(n21519), .B(
        n21411), .ZN(n21412) );
  OAI211_X1 U23441 ( .C1(n21414), .C2(n21522), .A(n21413), .B(n21412), .ZN(
        P3_U2715) );
  NOR4_X1 U23442 ( .A1(n21418), .A2(n21417), .A3(n21416), .A4(n21415), .ZN(
        n21440) );
  NAND2_X1 U23443 ( .A1(n21440), .A2(n21436), .ZN(n21423) );
  NAND3_X1 U23444 ( .A1(n21512), .A2(P3_EAX_REG_22__SCAN_IN), .A3(n21423), 
        .ZN(n21422) );
  OAI22_X1 U23445 ( .A1(n21419), .A2(n21522), .B1(n17468), .B2(n21485), .ZN(
        n21420) );
  AOI21_X1 U23446 ( .B1(BUF2_REG_6__SCAN_IN), .B2(n21491), .A(n21420), .ZN(
        n21421) );
  OAI211_X1 U23447 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n21423), .A(n21422), .B(
        n21421), .ZN(P3_U2713) );
  AOI22_X1 U23448 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n21492), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n21491), .ZN(n21428) );
  INV_X1 U23449 ( .A(n21435), .ZN(n21431) );
  NAND2_X1 U23450 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n21431), .ZN(n21430) );
  AOI211_X1 U23451 ( .C1(n21425), .C2(n21430), .A(n21424), .B(n21461), .ZN(
        n21426) );
  INV_X1 U23452 ( .A(n21426), .ZN(n21427) );
  OAI211_X1 U23453 ( .C1(n21429), .C2(n21522), .A(n21428), .B(n21427), .ZN(
        P3_U2716) );
  AOI22_X1 U23454 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n21492), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n21491), .ZN(n21433) );
  OAI211_X1 U23455 ( .C1(n21431), .C2(P3_EAX_REG_18__SCAN_IN), .A(n21519), .B(
        n21430), .ZN(n21432) );
  OAI211_X1 U23456 ( .C1(n21434), .C2(n21522), .A(n21433), .B(n21432), .ZN(
        P3_U2717) );
  AOI22_X1 U23457 ( .A1(BUF2_REG_17__SCAN_IN), .A2(n21492), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n21491), .ZN(n21438) );
  OAI211_X1 U23458 ( .C1(n21436), .C2(P3_EAX_REG_17__SCAN_IN), .A(n21519), .B(
        n21435), .ZN(n21437) );
  OAI211_X1 U23459 ( .C1(n21439), .C2(n21522), .A(n21438), .B(n21437), .ZN(
        P3_U2718) );
  AOI22_X1 U23460 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n21492), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n21491), .ZN(n21446) );
  INV_X1 U23461 ( .A(n21440), .ZN(n21442) );
  NAND2_X1 U23462 ( .A1(n21487), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n21486) );
  NAND2_X1 U23463 ( .A1(n21481), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n21480) );
  OAI211_X1 U23464 ( .C1(n21444), .C2(P3_EAX_REG_25__SCAN_IN), .A(n21519), .B(
        n21449), .ZN(n21445) );
  OAI211_X1 U23465 ( .C1(n21447), .C2(n21522), .A(n21446), .B(n21445), .ZN(
        P3_U2710) );
  AOI22_X1 U23466 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n21491), .B1(n21526), .B2(
        n21448), .ZN(n21453) );
  AOI211_X1 U23467 ( .C1(n21450), .C2(n21449), .A(n21475), .B(n21461), .ZN(
        n21451) );
  INV_X1 U23468 ( .A(n21451), .ZN(n21452) );
  OAI211_X1 U23469 ( .C1(n21485), .C2(n21454), .A(n21453), .B(n21452), .ZN(
        P3_U2709) );
  NAND2_X1 U23470 ( .A1(n21475), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n21474) );
  NAND2_X1 U23471 ( .A1(n21462), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n21457) );
  NAND3_X1 U23472 ( .A1(n21512), .A2(P3_EAX_REG_31__SCAN_IN), .A3(n21457), 
        .ZN(n21456) );
  NAND2_X1 U23473 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n21492), .ZN(n21455) );
  OAI211_X1 U23474 ( .C1(P3_EAX_REG_31__SCAN_IN), .C2(n21457), .A(n21456), .B(
        n21455), .ZN(P3_U2704) );
  AOI22_X1 U23475 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n21492), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n21491), .ZN(n21459) );
  OAI211_X1 U23476 ( .C1(n21462), .C2(P3_EAX_REG_30__SCAN_IN), .A(n21519), .B(
        n21457), .ZN(n21458) );
  OAI211_X1 U23477 ( .C1(n21460), .C2(n21522), .A(n21459), .B(n21458), .ZN(
        P3_U2705) );
  AOI22_X1 U23478 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n21492), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n21491), .ZN(n21466) );
  AOI211_X1 U23479 ( .C1(n21463), .C2(n21469), .A(n21462), .B(n21461), .ZN(
        n21464) );
  INV_X1 U23480 ( .A(n21464), .ZN(n21465) );
  OAI211_X1 U23481 ( .C1(n21467), .C2(n21522), .A(n21466), .B(n21465), .ZN(
        P3_U2706) );
  AOI22_X1 U23482 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n21491), .B1(n21526), .B2(
        n21468), .ZN(n21472) );
  OAI211_X1 U23483 ( .C1(n21470), .C2(P3_EAX_REG_28__SCAN_IN), .A(n21519), .B(
        n21469), .ZN(n21471) );
  OAI211_X1 U23484 ( .C1(n21485), .C2(n21473), .A(n21472), .B(n21471), .ZN(
        P3_U2707) );
  AOI22_X1 U23485 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n21492), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n21491), .ZN(n21477) );
  OAI211_X1 U23486 ( .C1(n21475), .C2(P3_EAX_REG_27__SCAN_IN), .A(n21519), .B(
        n21474), .ZN(n21476) );
  OAI211_X1 U23487 ( .C1(n21478), .C2(n21522), .A(n21477), .B(n21476), .ZN(
        P3_U2708) );
  AOI22_X1 U23488 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n21491), .B1(n21526), .B2(
        n21479), .ZN(n21483) );
  OAI211_X1 U23489 ( .C1(n21481), .C2(P3_EAX_REG_24__SCAN_IN), .A(n21519), .B(
        n21480), .ZN(n21482) );
  OAI211_X1 U23490 ( .C1(n21485), .C2(n21484), .A(n21483), .B(n21482), .ZN(
        P3_U2711) );
  AOI22_X1 U23491 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n21492), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n21491), .ZN(n21489) );
  OAI211_X1 U23492 ( .C1(n21487), .C2(P3_EAX_REG_23__SCAN_IN), .A(n21512), .B(
        n21486), .ZN(n21488) );
  OAI211_X1 U23493 ( .C1(n21490), .C2(n21522), .A(n21489), .B(n21488), .ZN(
        P3_U2712) );
  AOI22_X1 U23494 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n21492), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n21491), .ZN(n21495) );
  OAI211_X1 U23495 ( .C1(n21503), .C2(P3_EAX_REG_16__SCAN_IN), .A(n21512), .B(
        n21493), .ZN(n21494) );
  OAI211_X1 U23496 ( .C1(n21496), .C2(n21522), .A(n21495), .B(n21494), .ZN(
        P3_U2719) );
  NAND2_X1 U23497 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n21497), .ZN(n21502) );
  NAND2_X1 U23498 ( .A1(n21512), .A2(n21505), .ZN(n21500) );
  AOI22_X1 U23499 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21527), .B1(n21526), .B2(
        n21498), .ZN(n21499) );
  OAI221_X1 U23500 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n21502), .C1(n21501), 
        .C2(n21500), .A(n21499), .ZN(P3_U2721) );
  AOI21_X1 U23501 ( .B1(n21505), .B2(n21504), .A(n21503), .ZN(n21506) );
  AOI22_X1 U23502 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n21527), .B1(n21506), .B2(
        n21519), .ZN(n21507) );
  OAI21_X1 U23503 ( .B1(n21508), .B2(n21522), .A(n21507), .ZN(P3_U2720) );
  AOI22_X1 U23504 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n21527), .B1(n21510), .B2(
        n21509), .ZN(n21514) );
  NAND3_X1 U23505 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n21512), .A3(n21511), .ZN(
        n21513) );
  OAI211_X1 U23506 ( .C1(n21515), .C2(n21522), .A(n21514), .B(n21513), .ZN(
        P3_U2727) );
  AOI21_X1 U23507 ( .B1(n21518), .B2(n21517), .A(n21516), .ZN(n21520) );
  AOI22_X1 U23508 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n21527), .B1(n21520), .B2(
        n21519), .ZN(n21521) );
  OAI21_X1 U23509 ( .B1(n21523), .B2(n21522), .A(n21521), .ZN(P3_U2734) );
  NAND2_X1 U23510 ( .A1(n21524), .A2(n21529), .ZN(n21531) );
  AOI22_X1 U23511 ( .A1(n21527), .A2(BUF2_REG_0__SCAN_IN), .B1(n21526), .B2(
        n21525), .ZN(n21528) );
  OAI221_X1 U23512 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n21531), .C1(n21530), 
        .C2(n21529), .A(n21528), .ZN(P3_U2735) );
  INV_X1 U23513 ( .A(n21532), .ZN(n21951) );
  AOI222_X1 U23514 ( .A1(n21732), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n21533), 
        .B2(n21555), .C1(n21535), .C2(n21951), .ZN(n21534) );
  INV_X1 U23515 ( .A(n21560), .ZN(n21557) );
  AOI22_X1 U23516 ( .A1(n21560), .A2(n21535), .B1(n21534), .B2(n21557), .ZN(
        P3_U3290) );
  AOI22_X1 U23517 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21812), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n21536), .ZN(n21543) );
  NOR2_X1 U23518 ( .A1(n21537), .A2(n21732), .ZN(n21542) );
  AOI222_X1 U23519 ( .A1(n21539), .A2(n21555), .B1(n21538), .B2(n21951), .C1(
        n21543), .C2(n21542), .ZN(n21540) );
  AOI22_X1 U23520 ( .A1(n21560), .A2(n21541), .B1(n21540), .B2(n21557), .ZN(
        P3_U3289) );
  NOR2_X1 U23521 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21549), .ZN(
        n21548) );
  INV_X1 U23522 ( .A(n21542), .ZN(n21544) );
  OAI22_X1 U23523 ( .A1(n21546), .A2(n21545), .B1(n21544), .B2(n21543), .ZN(
        n21547) );
  AOI21_X1 U23524 ( .B1(n21548), .B2(n21951), .A(n21547), .ZN(n21552) );
  AOI21_X1 U23525 ( .B1(n21951), .B2(n21549), .A(n21560), .ZN(n21551) );
  OAI22_X1 U23526 ( .A1(n21560), .A2(n21552), .B1(n21551), .B2(n21550), .ZN(
        P3_U3288) );
  INV_X1 U23527 ( .A(n21553), .ZN(n21554) );
  AOI22_X1 U23528 ( .A1(n21951), .A2(n21556), .B1(n21555), .B2(n21554), .ZN(
        n21558) );
  AOI22_X1 U23529 ( .A1(n21560), .A2(n21559), .B1(n21558), .B2(n21557), .ZN(
        P3_U3285) );
  OAI21_X1 U23530 ( .B1(n21925), .B2(n21561), .A(n21897), .ZN(n21850) );
  NAND2_X1 U23531 ( .A1(n21911), .A2(n21936), .ZN(n21730) );
  OAI21_X1 U23532 ( .B1(n21563), .B2(n21562), .A(n21746), .ZN(n21564) );
  OAI21_X1 U23533 ( .B1(n21565), .B2(n21911), .A(n21564), .ZN(n21851) );
  OAI22_X1 U23534 ( .A1(n21567), .A2(n21927), .B1(n21566), .B2(n21847), .ZN(
        n21568) );
  AOI211_X1 U23535 ( .C1(n21569), .C2(n21730), .A(n21851), .B(n21568), .ZN(
        n21733) );
  OAI21_X1 U23536 ( .B1(n21925), .B2(n21570), .A(n21733), .ZN(n21571) );
  OAI21_X1 U23537 ( .B1(n21850), .B2(n21571), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n21577) );
  NOR2_X1 U23538 ( .A1(n21572), .A2(n21930), .ZN(n21864) );
  AOI22_X1 U23539 ( .A1(n21939), .A2(n21574), .B1(n21573), .B2(n21864), .ZN(
        n21575) );
  OAI221_X1 U23540 ( .B1(n11153), .B2(n21577), .C1(n14030), .C2(n21576), .A(
        n21575), .ZN(P3_U2841) );
  NAND2_X1 U23541 ( .A1(n21897), .A2(n21826), .ZN(n21666) );
  AND2_X1 U23542 ( .A1(n11153), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n21579) );
  NAND2_X1 U23543 ( .A1(n21911), .A2(n21925), .ZN(n21696) );
  INV_X1 U23544 ( .A(n21696), .ZN(n21859) );
  AOI221_X1 U23545 ( .B1(n21936), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C1(
        n21859), .C2(n21732), .A(n21930), .ZN(n21578) );
  AOI211_X1 U23546 ( .C1(n21835), .C2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n21579), .B(n21578), .ZN(n21580) );
  OAI221_X1 U23547 ( .B1(n21582), .B2(n21666), .C1(n21581), .C2(n21653), .A(
        n21580), .ZN(P3_U2862) );
  AOI22_X1 U23548 ( .A1(n11153), .A2(P3_REIP_REG_1__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21835), .ZN(n21589) );
  NOR2_X1 U23549 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21746), .ZN(
        n21583) );
  NOR2_X1 U23550 ( .A1(n21899), .A2(n21583), .ZN(n21585) );
  AND2_X1 U23551 ( .A1(n21732), .A2(n21696), .ZN(n21584) );
  MUX2_X1 U23552 ( .A(n21585), .B(n21584), .S(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n21587) );
  OAI221_X1 U23553 ( .B1(n21587), .B2(n21826), .C1(n21587), .C2(n21586), .A(
        n21897), .ZN(n21588) );
  OAI211_X1 U23554 ( .C1(n21590), .C2(n21653), .A(n21589), .B(n21588), .ZN(
        P3_U2861) );
  NAND2_X1 U23555 ( .A1(n21732), .A2(n21731), .ZN(n21872) );
  AOI211_X1 U23556 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n21872), .A(
        n11304), .B(n13796), .ZN(n21592) );
  NAND2_X1 U23557 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21601), .ZN(
        n21602) );
  AOI21_X1 U23558 ( .B1(n21602), .B2(n21605), .A(n21911), .ZN(n21591) );
  NOR2_X1 U23559 ( .A1(n21592), .A2(n21591), .ZN(n21594) );
  AOI21_X1 U23560 ( .B1(n21936), .B2(n21732), .A(n11304), .ZN(n21600) );
  NAND3_X1 U23561 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21600), .A3(
        n13796), .ZN(n21593) );
  OAI211_X1 U23562 ( .C1(n21595), .C2(n21614), .A(n21594), .B(n21593), .ZN(
        n21596) );
  AOI22_X1 U23563 ( .A1(n21897), .A2(n21596), .B1(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n21835), .ZN(n21598) );
  OAI211_X1 U23564 ( .C1(n21666), .C2(n21599), .A(n21598), .B(n21597), .ZN(
        P3_U2860) );
  AOI22_X1 U23565 ( .A1(n21875), .A2(n21605), .B1(n21601), .B2(n21600), .ZN(
        n21634) );
  AOI21_X1 U23566 ( .B1(n21634), .B2(n21626), .A(n21930), .ZN(n21609) );
  AOI22_X1 U23567 ( .A1(n21746), .A2(n21603), .B1(n21731), .B2(n21602), .ZN(
        n21604) );
  OAI211_X1 U23568 ( .C1(n21911), .C2(n21605), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n21604), .ZN(n21615) );
  OAI22_X1 U23569 ( .A1(n21653), .A2(n21607), .B1(n21666), .B2(n21606), .ZN(
        n21608) );
  AOI21_X1 U23570 ( .B1(n21609), .B2(n21615), .A(n21608), .ZN(n21611) );
  OAI211_X1 U23571 ( .C1(n21828), .C2(n21626), .A(n21611), .B(n21610), .ZN(
        P3_U2859) );
  NAND2_X1 U23572 ( .A1(n11153), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n21621) );
  OAI22_X1 U23573 ( .A1(n21614), .A2(n21613), .B1(n21847), .B2(n21612), .ZN(
        n21619) );
  NOR2_X1 U23574 ( .A1(n21634), .A2(n21626), .ZN(n21617) );
  AND2_X1 U23575 ( .A1(n21843), .A2(n21615), .ZN(n21616) );
  MUX2_X1 U23576 ( .A(n21617), .B(n21616), .S(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(n21618) );
  OAI21_X1 U23577 ( .B1(n21619), .B2(n21618), .A(n21897), .ZN(n21620) );
  OAI211_X1 U23578 ( .C1(n21828), .C2(n21625), .A(n21621), .B(n21620), .ZN(
        P3_U2858) );
  OAI211_X1 U23579 ( .C1(n11304), .C2(n21622), .A(n21897), .B(n21872), .ZN(
        n21624) );
  OAI221_X1 U23580 ( .B1(n21624), .B2(n21875), .C1(n21624), .C2(n21623), .A(
        n14030), .ZN(n21641) );
  NOR4_X1 U23581 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21634), .A3(
        n21626), .A4(n21625), .ZN(n21630) );
  OAI22_X1 U23582 ( .A1(n21653), .A2(n21628), .B1(n21666), .B2(n21627), .ZN(
        n21629) );
  AOI21_X1 U23583 ( .B1(n21897), .B2(n21630), .A(n21629), .ZN(n21632) );
  OAI211_X1 U23584 ( .C1(n11439), .C2(n21641), .A(n21632), .B(n21631), .ZN(
        P3_U2857) );
  NOR2_X1 U23585 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21930), .ZN(
        n21638) );
  NOR2_X1 U23586 ( .A1(n21634), .A2(n21633), .ZN(n21644) );
  OAI22_X1 U23587 ( .A1(n21653), .A2(n21636), .B1(n21666), .B2(n21635), .ZN(
        n21637) );
  AOI21_X1 U23588 ( .B1(n21638), .B2(n21644), .A(n21637), .ZN(n21640) );
  NAND2_X1 U23589 ( .A1(n11153), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n21639) );
  OAI211_X1 U23590 ( .C1(n21642), .C2(n21641), .A(n21640), .B(n21639), .ZN(
        P3_U2856) );
  INV_X1 U23591 ( .A(n21666), .ZN(n21759) );
  INV_X1 U23592 ( .A(n21643), .ZN(n21650) );
  NAND2_X1 U23593 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21644), .ZN(
        n21667) );
  NAND2_X1 U23594 ( .A1(n21655), .A2(n21667), .ZN(n21649) );
  OAI211_X1 U23595 ( .C1(n21645), .C2(n21911), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n21872), .ZN(n21646) );
  AOI21_X1 U23596 ( .B1(n21883), .B2(n21647), .A(n21646), .ZN(n21657) );
  OAI22_X1 U23597 ( .A1(n21657), .A2(n21930), .B1(n21655), .B2(n21828), .ZN(
        n21648) );
  AOI22_X1 U23598 ( .A1(n21759), .A2(n21650), .B1(n21649), .B2(n21648), .ZN(
        n21652) );
  NAND2_X1 U23599 ( .A1(n11153), .A2(P3_REIP_REG_7__SCAN_IN), .ZN(n21651) );
  OAI211_X1 U23600 ( .C1(n21654), .C2(n21653), .A(n21652), .B(n21651), .ZN(
        P3_U2855) );
  NOR3_X1 U23601 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21655), .A3(
        n21667), .ZN(n21659) );
  NOR3_X1 U23602 ( .A1(n21899), .A2(n21657), .A3(n21656), .ZN(n21658) );
  AOI211_X1 U23603 ( .C1(n21871), .C2(n21660), .A(n21659), .B(n21658), .ZN(
        n21661) );
  OAI22_X1 U23604 ( .A1(n21661), .A2(n21930), .B1(n21868), .B2(n21660), .ZN(
        n21662) );
  AOI211_X1 U23605 ( .C1(n21835), .C2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n21663), .B(n21662), .ZN(n21664) );
  OAI21_X1 U23606 ( .B1(n21666), .B2(n21665), .A(n21664), .ZN(P3_U2854) );
  NOR2_X1 U23607 ( .A1(n21668), .A2(n21667), .ZN(n21713) );
  OAI21_X1 U23608 ( .B1(n21713), .B2(n21686), .A(n21897), .ZN(n21943) );
  NOR2_X1 U23609 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n21943), .ZN(
        n21669) );
  AOI22_X1 U23610 ( .A1(n11153), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n21671), 
        .B2(n21669), .ZN(n21678) );
  NOR2_X1 U23611 ( .A1(n21871), .A2(n21826), .ZN(n21881) );
  NAND2_X1 U23612 ( .A1(n21826), .A2(n21670), .ZN(n21933) );
  OAI211_X1 U23613 ( .C1(n21671), .C2(n21881), .A(n21897), .B(n21933), .ZN(
        n21672) );
  AOI221_X1 U23614 ( .B1(n21942), .B2(n21731), .C1(n21931), .C2(n21731), .A(
        n21672), .ZN(n21918) );
  NOR2_X1 U23615 ( .A1(n21685), .A2(n21911), .ZN(n21695) );
  NAND2_X1 U23616 ( .A1(n21875), .A2(n21673), .ZN(n21926) );
  NAND2_X1 U23617 ( .A1(n21746), .A2(n21674), .ZN(n21712) );
  OAI211_X1 U23618 ( .C1(n21928), .C2(n21927), .A(n21926), .B(n21712), .ZN(
        n21921) );
  AOI211_X1 U23619 ( .C1(n21675), .C2(n21746), .A(n21695), .B(n21921), .ZN(
        n21680) );
  OAI211_X1 U23620 ( .C1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n21925), .A(
        n21918), .B(n21680), .ZN(n21676) );
  NAND3_X1 U23621 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14030), .A3(
        n21676), .ZN(n21677) );
  OAI211_X1 U23622 ( .C1(n21679), .C2(n21868), .A(n21678), .B(n21677), .ZN(
        P3_U2851) );
  NAND2_X1 U23623 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21683) );
  OAI211_X1 U23624 ( .C1(n21681), .C2(n21881), .A(n21680), .B(n21933), .ZN(
        n21682) );
  AOI21_X1 U23625 ( .B1(n21683), .B2(n21746), .A(n21682), .ZN(n21910) );
  OAI21_X1 U23626 ( .B1(n21684), .B2(n21931), .A(n21731), .ZN(n21909) );
  OAI21_X1 U23627 ( .B1(n21713), .B2(n21686), .A(n21685), .ZN(n21687) );
  OAI222_X1 U23628 ( .A1(n21688), .A2(n21910), .B1(n21688), .B2(n21909), .C1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n21687), .ZN(n21689) );
  AOI22_X1 U23629 ( .A1(n21897), .A2(n21689), .B1(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n21835), .ZN(n21691) );
  OAI211_X1 U23630 ( .C1(n21692), .C2(n21868), .A(n21691), .B(n21690), .ZN(
        P3_U2850) );
  AOI22_X1 U23631 ( .A1(n11153), .A2(P3_REIP_REG_14__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n21835), .ZN(n21709) );
  NAND3_X1 U23632 ( .A1(n21700), .A2(n21713), .A3(n21693), .ZN(n21704) );
  OAI21_X1 U23633 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n21911), .A(
        n21909), .ZN(n21702) );
  INV_X1 U23634 ( .A(n21926), .ZN(n21694) );
  AOI211_X1 U23635 ( .C1(n21697), .C2(n21696), .A(n21695), .B(n21694), .ZN(
        n21698) );
  OAI221_X1 U23636 ( .B1(n21936), .B2(n21700), .C1(n21936), .C2(n21699), .A(
        n21698), .ZN(n21701) );
  OAI21_X1 U23637 ( .B1(n21702), .B2(n21701), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21703) );
  OAI211_X1 U23638 ( .C1(n21927), .C2(n21705), .A(n21704), .B(n21703), .ZN(
        n21707) );
  AOI22_X1 U23639 ( .A1(n21897), .A2(n21707), .B1(n21759), .B2(n21706), .ZN(
        n21708) );
  OAI211_X1 U23640 ( .C1(n21710), .C2(n21868), .A(n21709), .B(n21708), .ZN(
        P3_U2848) );
  OAI21_X1 U23641 ( .B1(n21718), .B2(n21931), .A(n21731), .ZN(n21711) );
  NAND4_X1 U23642 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21712), .A3(
        n21926), .A4(n21711), .ZN(n21717) );
  NAND2_X1 U23643 ( .A1(n21713), .A2(n21717), .ZN(n21715) );
  NAND2_X1 U23644 ( .A1(n21871), .A2(n21720), .ZN(n21896) );
  OAI22_X1 U23645 ( .A1(n21718), .A2(n21715), .B1(n21896), .B2(n21714), .ZN(
        n21716) );
  AOI22_X1 U23646 ( .A1(n11153), .A2(P3_REIP_REG_15__SCAN_IN), .B1(n21897), 
        .B2(n21716), .ZN(n21727) );
  INV_X1 U23647 ( .A(n21869), .ZN(n21719) );
  NOR3_X1 U23648 ( .A1(n21719), .A2(n21847), .A3(n21930), .ZN(n21725) );
  AOI21_X1 U23649 ( .B1(n21718), .B2(n21730), .A(n21717), .ZN(n21898) );
  NOR2_X1 U23650 ( .A1(n21719), .A2(n21847), .ZN(n21901) );
  AOI211_X1 U23651 ( .C1(n21871), .C2(n21720), .A(n21901), .B(n21930), .ZN(
        n21722) );
  AOI211_X1 U23652 ( .C1(n21898), .C2(n21722), .A(n11153), .B(n21721), .ZN(
        n21723) );
  AOI21_X1 U23653 ( .B1(n21725), .B2(n21724), .A(n21723), .ZN(n21726) );
  OAI211_X1 U23654 ( .C1(n21728), .C2(n21868), .A(n21727), .B(n21726), .ZN(
        P3_U2847) );
  AOI22_X1 U23655 ( .A1(n11153), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n21939), 
        .B2(n21729), .ZN(n21736) );
  INV_X1 U23656 ( .A(n21730), .ZN(n21919) );
  OAI21_X1 U23657 ( .B1(n21732), .B2(n21745), .A(n21731), .ZN(n21743) );
  OAI211_X1 U23658 ( .C1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n21919), .A(
        n21743), .B(n21733), .ZN(n21734) );
  OAI221_X1 U23659 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n21757), 
        .C1(n21737), .C2(n21734), .A(n21897), .ZN(n21735) );
  OAI211_X1 U23660 ( .C1(n21828), .C2(n21737), .A(n21736), .B(n21735), .ZN(
        P3_U2840) );
  INV_X1 U23661 ( .A(n21738), .ZN(n21741) );
  NOR3_X1 U23662 ( .A1(n21741), .A2(n21740), .A3(n21739), .ZN(n21795) );
  NAND2_X1 U23663 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21747) );
  AND2_X1 U23664 ( .A1(n21875), .A2(n21742), .ZN(n21831) );
  INV_X1 U23665 ( .A(n21743), .ZN(n21744) );
  AOI21_X1 U23666 ( .B1(n21746), .B2(n21745), .A(n21744), .ZN(n21830) );
  INV_X1 U23667 ( .A(n21830), .ZN(n21776) );
  AOI211_X1 U23668 ( .C1(n21843), .C2(n21747), .A(n21831), .B(n21776), .ZN(
        n21764) );
  OAI22_X1 U23669 ( .A1(n21764), .A2(n21762), .B1(n21927), .B2(n21748), .ZN(
        n21749) );
  AOI21_X1 U23670 ( .B1(n21795), .B2(n21762), .A(n21749), .ZN(n21751) );
  OAI22_X1 U23671 ( .A1(n21751), .A2(n21930), .B1(n21868), .B2(n21750), .ZN(
        n21752) );
  AOI21_X1 U23672 ( .B1(n21759), .B2(n21753), .A(n21752), .ZN(n21755) );
  OAI211_X1 U23673 ( .C1(n21828), .C2(n21762), .A(n21755), .B(n21754), .ZN(
        P3_U2837) );
  AOI21_X1 U23674 ( .B1(n21757), .B2(n21756), .A(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21770) );
  AND2_X1 U23675 ( .A1(n21759), .A2(n21758), .ZN(n21782) );
  AND2_X1 U23676 ( .A1(n21871), .A2(n21777), .ZN(n21761) );
  AOI211_X1 U23677 ( .C1(n21843), .C2(n21762), .A(n21761), .B(n21760), .ZN(
        n21763) );
  AOI21_X1 U23678 ( .B1(n21764), .B2(n21763), .A(n21930), .ZN(n21765) );
  AOI211_X1 U23679 ( .C1(n21835), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n21782), .B(n21765), .ZN(n21769) );
  AOI21_X1 U23680 ( .B1(n21767), .B2(n21939), .A(n21766), .ZN(n21768) );
  OAI21_X1 U23681 ( .B1(n21770), .B2(n21769), .A(n21768), .ZN(P3_U2836) );
  INV_X1 U23682 ( .A(n21771), .ZN(n21785) );
  INV_X1 U23683 ( .A(n21772), .ZN(n21774) );
  OAI211_X1 U23684 ( .C1(n11304), .C2(n21774), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n21773), .ZN(n21775) );
  AOI211_X1 U23685 ( .C1(n21871), .C2(n21777), .A(n21776), .B(n21775), .ZN(
        n21779) );
  OAI22_X1 U23686 ( .A1(n21779), .A2(n21930), .B1(n21778), .B2(n21828), .ZN(
        n21781) );
  OAI22_X1 U23687 ( .A1(n21782), .A2(n21781), .B1(n21780), .B2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21783) );
  OAI211_X1 U23688 ( .C1(n21785), .C2(n21868), .A(n21784), .B(n21783), .ZN(
        P3_U2835) );
  OAI21_X1 U23689 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n21936), .A(
        n21786), .ZN(n21802) );
  OAI211_X1 U23690 ( .C1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n21859), .A(
        n21897), .B(n21787), .ZN(n21788) );
  NOR2_X1 U23691 ( .A1(n21802), .A2(n21788), .ZN(n21791) );
  NAND2_X1 U23692 ( .A1(n21794), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n21790) );
  AOI22_X1 U23693 ( .A1(n21871), .A2(n21790), .B1(n21826), .B2(n21789), .ZN(
        n21807) );
  AOI21_X1 U23694 ( .B1(n21791), .B2(n21807), .A(n21798), .ZN(n21792) );
  AOI22_X1 U23695 ( .A1(n11153), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n21792), 
        .B2(n14030), .ZN(n21800) );
  AOI22_X1 U23696 ( .A1(n21871), .A2(n21794), .B1(n21826), .B2(n21793), .ZN(
        n21797) );
  NAND2_X1 U23697 ( .A1(n21796), .A2(n21795), .ZN(n21815) );
  NAND2_X1 U23698 ( .A1(n21797), .A2(n21815), .ZN(n21805) );
  NAND3_X1 U23699 ( .A1(n21897), .A2(n21798), .A3(n21805), .ZN(n21799) );
  OAI211_X1 U23700 ( .C1(n21801), .C2(n21868), .A(n21800), .B(n21799), .ZN(
        P3_U2833) );
  AOI211_X1 U23701 ( .C1(n21843), .C2(n21804), .A(n21803), .B(n21802), .ZN(
        n21813) );
  AOI21_X1 U23702 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n21805), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21806) );
  AOI211_X1 U23703 ( .C1(n21813), .C2(n21807), .A(n21806), .B(n21930), .ZN(
        n21808) );
  AOI21_X1 U23704 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n21835), .A(
        n21808), .ZN(n21810) );
  OAI211_X1 U23705 ( .C1(n21811), .C2(n21868), .A(n21810), .B(n21809), .ZN(
        P3_U2832) );
  NOR3_X1 U23706 ( .A1(n21899), .A2(n21813), .A3(n21812), .ZN(n21819) );
  OR2_X1 U23707 ( .A1(n21814), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n21816) );
  OAI22_X1 U23708 ( .A1(n21817), .A2(n21927), .B1(n21816), .B2(n21815), .ZN(
        n21818) );
  AOI211_X1 U23709 ( .C1(n21826), .C2(n21820), .A(n21819), .B(n21818), .ZN(
        n21824) );
  AOI22_X1 U23710 ( .A1(n21835), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n21939), .B2(n21821), .ZN(n21823) );
  OAI211_X1 U23711 ( .C1(n21824), .C2(n21930), .A(n21823), .B(n21822), .ZN(
        P3_U2831) );
  AOI22_X1 U23712 ( .A1(n21871), .A2(n21827), .B1(n21826), .B2(n21825), .ZN(
        n21829) );
  NAND3_X1 U23713 ( .A1(n21830), .A2(n21829), .A3(n21828), .ZN(n21842) );
  NOR3_X1 U23714 ( .A1(n21831), .A2(n21833), .A3(n21842), .ZN(n21832) );
  NOR2_X1 U23715 ( .A1(n11153), .A2(n21832), .ZN(n21841) );
  OAI21_X1 U23716 ( .B1(n21835), .B2(n21834), .A(n21833), .ZN(n21836) );
  AOI22_X1 U23717 ( .A1(n21939), .A2(n21837), .B1(n21841), .B2(n21836), .ZN(
        n21838) );
  OAI21_X1 U23718 ( .B1(n14030), .B2(n21839), .A(n21838), .ZN(P3_U2839) );
  AOI22_X1 U23719 ( .A1(n11153), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n21864), 
        .B2(n21840), .ZN(n21845) );
  OAI211_X1 U23720 ( .C1(n21843), .C2(n21842), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n21841), .ZN(n21844) );
  OAI211_X1 U23721 ( .C1(n21846), .C2(n21868), .A(n21845), .B(n21844), .ZN(
        P3_U2838) );
  OAI22_X1 U23722 ( .A1(n21849), .A2(n21927), .B1(n21848), .B2(n21847), .ZN(
        n21852) );
  NOR3_X1 U23723 ( .A1(n21852), .A2(n21851), .A3(n21850), .ZN(n21853) );
  NOR2_X1 U23724 ( .A1(n21853), .A2(n11153), .ZN(n21862) );
  AOI22_X1 U23725 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21862), .B1(
        n21864), .B2(n21854), .ZN(n21856) );
  NAND2_X1 U23726 ( .A1(n11153), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n21855) );
  OAI211_X1 U23727 ( .C1(n21857), .C2(n21868), .A(n21856), .B(n21855), .ZN(
        P3_U2843) );
  NOR3_X1 U23728 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21859), .A3(
        n21858), .ZN(n21861) );
  AOI221_X1 U23729 ( .B1(n21862), .B2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), 
        .C1(n21861), .C2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A(n21860), .ZN(
        n21866) );
  NAND3_X1 U23730 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21864), .A3(
        n21863), .ZN(n21865) );
  OAI211_X1 U23731 ( .C1(n21868), .C2(n21867), .A(n21866), .B(n21865), .ZN(
        P3_U2842) );
  AOI211_X1 U23732 ( .C1(n21871), .C2(n21870), .A(n21877), .B(n21869), .ZN(
        n21880) );
  NAND3_X1 U23733 ( .A1(n21873), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n21872), .ZN(n21874) );
  AOI21_X1 U23734 ( .B1(n21883), .B2(n21874), .A(n21930), .ZN(n21879) );
  OAI21_X1 U23735 ( .B1(n21877), .B2(n21876), .A(n21875), .ZN(n21878) );
  OAI211_X1 U23736 ( .C1(n21881), .C2(n21880), .A(n21879), .B(n21878), .ZN(
        n21890) );
  OAI221_X1 U23737 ( .B1(n21890), .B2(n21883), .C1(n21890), .C2(n21882), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21889) );
  NOR2_X1 U23738 ( .A1(n21884), .A2(n21943), .ZN(n21903) );
  AOI22_X1 U23739 ( .A1(n21939), .A2(n21886), .B1(n21903), .B2(n21885), .ZN(
        n21887) );
  OAI221_X1 U23740 ( .B1(n11153), .B2(n21889), .C1(n14030), .C2(n21888), .A(
        n21887), .ZN(P3_U2844) );
  NAND2_X1 U23741 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21890), .ZN(
        n21895) );
  AOI22_X1 U23742 ( .A1(n21939), .A2(n21892), .B1(n21903), .B2(n21891), .ZN(
        n21893) );
  OAI221_X1 U23743 ( .B1(n11153), .B2(n21895), .C1(n14030), .C2(n21894), .A(
        n21893), .ZN(P3_U2845) );
  OAI211_X1 U23744 ( .C1(n21899), .C2(n21898), .A(n21897), .B(n21896), .ZN(
        n21900) );
  OAI21_X1 U23745 ( .B1(n21901), .B2(n21900), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21907) );
  AOI22_X1 U23746 ( .A1(n21904), .A2(n21939), .B1(n21903), .B2(n21902), .ZN(
        n21905) );
  OAI221_X1 U23747 ( .B1(n11153), .B2(n21907), .C1(n14030), .C2(n21906), .A(
        n21905), .ZN(P3_U2846) );
  AOI22_X1 U23748 ( .A1(n11153), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n21939), 
        .B2(n21908), .ZN(n21914) );
  OAI211_X1 U23749 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n21911), .A(
        n21910), .B(n21909), .ZN(n21912) );
  OAI211_X1 U23750 ( .C1(n21930), .C2(n21912), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n14030), .ZN(n21913) );
  OAI211_X1 U23751 ( .C1(n21943), .C2(n21915), .A(n21914), .B(n21913), .ZN(
        P3_U2849) );
  NAND2_X1 U23752 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n21916), .ZN(
        n21924) );
  AOI22_X1 U23753 ( .A1(n11153), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n21939), 
        .B2(n21917), .ZN(n21923) );
  OAI21_X1 U23754 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21919), .A(
        n21918), .ZN(n21920) );
  OAI211_X1 U23755 ( .C1(n21921), .C2(n21920), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n14030), .ZN(n21922) );
  OAI211_X1 U23756 ( .C1(n21924), .C2(n21943), .A(n21923), .B(n21922), .ZN(
        P3_U2852) );
  AOI21_X1 U23757 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n21925), .A(
        n11304), .ZN(n21932) );
  OAI21_X1 U23758 ( .B1(n21928), .B2(n21927), .A(n21926), .ZN(n21929) );
  AOI211_X1 U23759 ( .C1(n21932), .C2(n21931), .A(n21930), .B(n21929), .ZN(
        n21934) );
  OAI211_X1 U23760 ( .C1(n21936), .C2(n21935), .A(n21934), .B(n21933), .ZN(
        n21937) );
  NAND2_X1 U23761 ( .A1(n14030), .A2(n21937), .ZN(n21941) );
  AOI22_X1 U23762 ( .A1(n11153), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n21939), 
        .B2(n21938), .ZN(n21940) );
  OAI221_X1 U23763 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21943), .C1(
        n21942), .C2(n21941), .A(n21940), .ZN(P3_U2853) );
  INV_X1 U23764 ( .A(n21944), .ZN(n21948) );
  NOR2_X1 U23765 ( .A1(n21946), .A2(n21945), .ZN(n21947) );
  OAI21_X1 U23766 ( .B1(n21949), .B2(n21948), .A(n21947), .ZN(P3_U3282) );
  AOI211_X1 U23767 ( .C1(n21952), .C2(n21951), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n21950), .ZN(n21953) );
  AOI211_X1 U23768 ( .C1(n21956), .C2(n21955), .A(n21954), .B(n21953), .ZN(
        n21957) );
  OAI221_X1 U23769 ( .B1(n21960), .B2(n21959), .C1(n21960), .C2(n21958), .A(
        n21957), .ZN(P3_U2996) );
  NOR2_X1 U23770 ( .A1(n21962), .A2(n21961), .ZN(n21966) );
  MUX2_X1 U23771 ( .A(P3_MORE_REG_SCAN_IN), .B(n21963), .S(n21966), .Z(
        P3_U3295) );
  OAI21_X1 U23772 ( .B1(n21966), .B2(n21965), .A(n21964), .ZN(P3_U2637) );
  INV_X1 U23773 ( .A(n21967), .ZN(n21968) );
  AOI211_X1 U23774 ( .C1(n20633), .C2(n22322), .A(n21969), .B(n21968), .ZN(
        n21975) );
  OAI211_X1 U23775 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21971), .A(n21970), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21972) );
  AOI21_X1 U23776 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n21972), .A(n22297), 
        .ZN(n21974) );
  NAND2_X1 U23777 ( .A1(n21975), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21973) );
  OAI21_X1 U23778 ( .B1(n21975), .B2(n21974), .A(n21973), .ZN(P1_U3485) );
  NAND2_X1 U23779 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21976), .ZN(
        n21985) );
  NOR2_X1 U23780 ( .A1(n21978), .A2(n21977), .ZN(n21984) );
  OAI21_X1 U23781 ( .B1(n21980), .B2(n22082), .A(n21979), .ZN(n21981) );
  AOI21_X1 U23782 ( .B1(n21982), .B2(n22075), .A(n21981), .ZN(n21983) );
  OAI221_X1 U23783 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n21985), 
        .C1(n16348), .C2(n21984), .A(n21983), .ZN(P1_U3017) );
  NOR2_X1 U23784 ( .A1(n21986), .A2(n22087), .ZN(n21988) );
  AOI22_X1 U23785 ( .A1(n21988), .A2(n22056), .B1(n22087), .B2(n21987), .ZN(
        n22002) );
  INV_X1 U23786 ( .A(n21989), .ZN(n21998) );
  NAND3_X1 U23787 ( .A1(n21991), .A2(n21990), .A3(n22075), .ZN(n21997) );
  NOR3_X1 U23788 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n21992), .A3(
        n22087), .ZN(n21993) );
  AOI211_X1 U23789 ( .C1(n22043), .C2(n21995), .A(n21994), .B(n21993), .ZN(
        n21996) );
  OAI211_X1 U23790 ( .C1(n21999), .C2(n21998), .A(n21997), .B(n21996), .ZN(
        n22000) );
  INV_X1 U23791 ( .A(n22000), .ZN(n22001) );
  OAI221_X1 U23792 ( .B1(n22003), .B2(n22051), .C1(n22003), .C2(n22002), .A(
        n22001), .ZN(P1_U3029) );
  INV_X1 U23793 ( .A(n22103), .ZN(n22004) );
  NAND2_X1 U23794 ( .A1(n22043), .A2(n22004), .ZN(n22006) );
  NAND2_X1 U23795 ( .A1(n22006), .A2(n22005), .ZN(n22007) );
  AOI21_X1 U23796 ( .B1(n22008), .B2(n22075), .A(n22007), .ZN(n22010) );
  OAI211_X1 U23797 ( .C1(n22013), .C2(n22011), .A(n22010), .B(n22009), .ZN(
        P1_U3028) );
  NAND2_X1 U23798 ( .A1(n22014), .A2(n22012), .ZN(n22019) );
  AOI22_X1 U23799 ( .A1(n22130), .A2(n22043), .B1(n22021), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n22018) );
  OAI21_X1 U23800 ( .B1(n22015), .B2(n22014), .A(n22013), .ZN(n22022) );
  AOI22_X1 U23801 ( .A1(n22016), .A2(n22075), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n22022), .ZN(n22017) );
  OAI211_X1 U23802 ( .C1(n22033), .C2(n22019), .A(n22018), .B(n22017), .ZN(
        P1_U3025) );
  NAND3_X1 U23803 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n22020), .ZN(n22026) );
  AOI22_X1 U23804 ( .A1(n22043), .A2(n22123), .B1(n22021), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n22025) );
  AOI22_X1 U23805 ( .A1(n22023), .A2(n22075), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n22022), .ZN(n22024) );
  OAI211_X1 U23806 ( .C1(n22033), .C2(n22026), .A(n22025), .B(n22024), .ZN(
        P1_U3026) );
  INV_X1 U23807 ( .A(n22027), .ZN(n22029) );
  OAI22_X1 U23808 ( .A1(n22078), .A2(n22030), .B1(n22029), .B2(n22028), .ZN(
        n22048) );
  OAI22_X1 U23809 ( .A1(n22144), .A2(n22082), .B1(n22066), .B2(n22155), .ZN(
        n22031) );
  INV_X1 U23810 ( .A(n22031), .ZN(n22036) );
  NOR2_X1 U23811 ( .A1(n22033), .A2(n22032), .ZN(n22049) );
  AOI22_X1 U23812 ( .A1(n22034), .A2(n22075), .B1(n22049), .B2(n22037), .ZN(
        n22035) );
  OAI211_X1 U23813 ( .C1(n22037), .C2(n22048), .A(n22036), .B(n22035), .ZN(
        P1_U3024) );
  INV_X1 U23814 ( .A(n22038), .ZN(n22042) );
  NOR2_X1 U23815 ( .A1(n22039), .A2(n22058), .ZN(n22040) );
  AOI211_X1 U23816 ( .C1(n22043), .C2(n22042), .A(n22041), .B(n22040), .ZN(
        n22046) );
  OAI211_X1 U23817 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n22049), .B(n22044), .ZN(n22045) );
  OAI211_X1 U23818 ( .C1(n22048), .C2(n22047), .A(n22046), .B(n22045), .ZN(
        P1_U3023) );
  NAND2_X1 U23819 ( .A1(n22050), .A2(n22049), .ZN(n22063) );
  OAI21_X1 U23820 ( .B1(n22053), .B2(n22052), .A(n22051), .ZN(n22054) );
  AOI21_X1 U23821 ( .B1(n22056), .B2(n22055), .A(n22054), .ZN(n22074) );
  OAI222_X1 U23822 ( .A1(n22060), .A2(n22082), .B1(n22066), .B2(n22059), .C1(
        n22058), .C2(n22057), .ZN(n22061) );
  INV_X1 U23823 ( .A(n22061), .ZN(n22062) );
  OAI221_X1 U23824 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n22063), .C1(
        n22065), .C2(n22074), .A(n22062), .ZN(P1_U3022) );
  AOI211_X1 U23825 ( .C1(n22065), .C2(n22073), .A(n22064), .B(n22063), .ZN(
        n22070) );
  OAI22_X1 U23826 ( .A1(n22068), .A2(n22082), .B1(n22067), .B2(n22066), .ZN(
        n22069) );
  AOI211_X1 U23827 ( .C1(n22071), .C2(n22075), .A(n22070), .B(n22069), .ZN(
        n22072) );
  OAI21_X1 U23828 ( .B1(n22074), .B2(n22073), .A(n22072), .ZN(P1_U3021) );
  AND3_X1 U23829 ( .A1(n22077), .A2(n22076), .A3(n22075), .ZN(n22085) );
  OAI211_X1 U23830 ( .C1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n22079), .A(
        n22078), .B(n22087), .ZN(n22081) );
  OAI211_X1 U23831 ( .C1(n22083), .C2(n22082), .A(n22081), .B(n22080), .ZN(
        n22084) );
  NOR2_X1 U23832 ( .A1(n22085), .A2(n22084), .ZN(n22086) );
  OAI21_X1 U23833 ( .B1(n22088), .B2(n22087), .A(n22086), .ZN(P1_U3030) );
  AOI22_X1 U23834 ( .A1(n14427), .A2(n22108), .B1(n22236), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n22089) );
  OAI21_X1 U23835 ( .B1(n22091), .B2(n22090), .A(n22089), .ZN(n22092) );
  AOI21_X1 U23836 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n22264), .A(
        n22092), .ZN(n22093) );
  OAI21_X1 U23837 ( .B1(n22095), .B2(n22094), .A(n22093), .ZN(n22096) );
  AOI21_X1 U23838 ( .B1(n22097), .B2(n22266), .A(n22096), .ZN(n22102) );
  NOR2_X1 U23839 ( .A1(n22099), .A2(n22098), .ZN(n22100) );
  OAI211_X1 U23840 ( .C1(P1_REIP_REG_3__SCAN_IN), .C2(n22100), .A(n22235), .B(
        n22113), .ZN(n22101) );
  OAI211_X1 U23841 ( .C1(n22103), .C2(n22276), .A(n22102), .B(n22101), .ZN(
        P1_U2837) );
  OAI22_X1 U23842 ( .A1(n22105), .A2(n22276), .B1(n22262), .B2(n22104), .ZN(
        n22106) );
  AOI211_X1 U23843 ( .C1(n22108), .C2(n22107), .A(n22106), .B(n22223), .ZN(
        n22109) );
  OAI21_X1 U23844 ( .B1(n22110), .B2(n22213), .A(n22109), .ZN(n22111) );
  AOI21_X1 U23845 ( .B1(n22112), .B2(n22125), .A(n22111), .ZN(n22117) );
  NOR2_X1 U23846 ( .A1(n22245), .A2(n22113), .ZN(n22115) );
  NAND2_X1 U23847 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n22115), .ZN(n22135) );
  INV_X1 U23848 ( .A(n22135), .ZN(n22114) );
  NOR2_X1 U23849 ( .A1(n22114), .A2(n22200), .ZN(n22124) );
  OAI21_X1 U23850 ( .B1(P1_REIP_REG_4__SCAN_IN), .B2(n22115), .A(n22124), .ZN(
        n22116) );
  OAI211_X1 U23851 ( .C1(n22257), .C2(n22118), .A(n22117), .B(n22116), .ZN(
        P1_U2836) );
  OAI21_X1 U23852 ( .B1(n22213), .B2(n22119), .A(n22193), .ZN(n22122) );
  OAI22_X1 U23853 ( .A1(n22135), .A2(P1_REIP_REG_5__SCAN_IN), .B1(n22262), 
        .B2(n22120), .ZN(n22121) );
  AOI211_X1 U23854 ( .C1(n22217), .C2(n22123), .A(n22122), .B(n22121), .ZN(
        n22128) );
  AOI22_X1 U23855 ( .A1(n22126), .A2(n22125), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n22124), .ZN(n22127) );
  OAI211_X1 U23856 ( .C1(n22129), .C2(n22257), .A(n22128), .B(n22127), .ZN(
        P1_U2835) );
  INV_X1 U23857 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n22132) );
  AOI22_X1 U23858 ( .A1(n22130), .A2(n22217), .B1(n22236), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n22131) );
  OAI211_X1 U23859 ( .C1(n22213), .C2(n22132), .A(n22131), .B(n22193), .ZN(
        n22133) );
  AOI21_X1 U23860 ( .B1(n22134), .B2(n22253), .A(n22133), .ZN(n22140) );
  NOR2_X1 U23861 ( .A1(n22136), .A2(n22135), .ZN(n22138) );
  NAND2_X1 U23862 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n22138), .ZN(n22156) );
  NAND2_X1 U23863 ( .A1(n22210), .A2(n22156), .ZN(n22154) );
  INV_X1 U23864 ( .A(n22154), .ZN(n22137) );
  OAI21_X1 U23865 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n22138), .A(n22137), .ZN(
        n22139) );
  OAI211_X1 U23866 ( .C1(n22257), .C2(n22141), .A(n22140), .B(n22139), .ZN(
        P1_U2834) );
  INV_X1 U23867 ( .A(n22142), .ZN(n22143) );
  NAND2_X1 U23868 ( .A1(n22266), .A2(n22143), .ZN(n22150) );
  INV_X1 U23869 ( .A(n22144), .ZN(n22148) );
  AOI21_X1 U23870 ( .B1(n22264), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n22223), .ZN(n22145) );
  OAI21_X1 U23871 ( .B1(n22262), .B2(n22146), .A(n22145), .ZN(n22147) );
  AOI21_X1 U23872 ( .B1(n22148), .B2(n22217), .A(n22147), .ZN(n22149) );
  NAND2_X1 U23873 ( .A1(n22150), .A2(n22149), .ZN(n22151) );
  AOI21_X1 U23874 ( .B1(n22152), .B2(n22253), .A(n22151), .ZN(n22153) );
  OAI221_X1 U23875 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(n22156), .C1(n22155), 
        .C2(n22154), .A(n22153), .ZN(P1_U2833) );
  NOR2_X1 U23876 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n22245), .ZN(n22162) );
  AOI22_X1 U23877 ( .A1(n22157), .A2(n22217), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n22236), .ZN(n22158) );
  OAI211_X1 U23878 ( .C1(n22213), .C2(n22159), .A(n22158), .B(n22193), .ZN(
        n22160) );
  AOI21_X1 U23879 ( .B1(n22162), .B2(n22161), .A(n22160), .ZN(n22166) );
  AOI22_X1 U23880 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n22164), .B1(n22253), 
        .B2(n22163), .ZN(n22165) );
  OAI211_X1 U23881 ( .C1(n22167), .C2(n22257), .A(n22166), .B(n22165), .ZN(
        P1_U2829) );
  AOI22_X1 U23882 ( .A1(n22169), .A2(n22266), .B1(n22253), .B2(n22168), .ZN(
        n22181) );
  NOR2_X1 U23883 ( .A1(n22245), .A2(n22170), .ZN(n22178) );
  OAI22_X1 U23884 ( .A1(n22172), .A2(n22276), .B1(n22171), .B2(n22262), .ZN(
        n22173) );
  INV_X1 U23885 ( .A(n22173), .ZN(n22174) );
  OAI211_X1 U23886 ( .C1(n22213), .C2(n22175), .A(n22174), .B(n22193), .ZN(
        n22176) );
  AOI221_X1 U23887 ( .B1(n22179), .B2(P1_REIP_REG_12__SCAN_IN), .C1(n22178), 
        .C2(n22177), .A(n22176), .ZN(n22180) );
  NAND2_X1 U23888 ( .A1(n22181), .A2(n22180), .ZN(P1_U2828) );
  INV_X1 U23889 ( .A(n22198), .ZN(n22192) );
  AOI21_X1 U23890 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n22210), .A(n22182), 
        .ZN(n22191) );
  OAI22_X1 U23891 ( .A1(n22213), .A2(n22184), .B1(n22183), .B2(n22262), .ZN(
        n22185) );
  AOI211_X1 U23892 ( .C1(n22186), .C2(n22217), .A(n22223), .B(n22185), .ZN(
        n22190) );
  AOI22_X1 U23893 ( .A1(n22188), .A2(n22253), .B1(n22266), .B2(n22187), .ZN(
        n22189) );
  OAI211_X1 U23894 ( .C1(n22192), .C2(n22191), .A(n22190), .B(n22189), .ZN(
        P1_U2825) );
  NAND2_X1 U23895 ( .A1(n22264), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n22194) );
  OAI211_X1 U23896 ( .C1(n22262), .C2(n22195), .A(n22194), .B(n22193), .ZN(
        n22196) );
  AOI21_X1 U23897 ( .B1(n22266), .B2(n22197), .A(n22196), .ZN(n22204) );
  OAI21_X1 U23898 ( .B1(n22200), .B2(n22199), .A(n22198), .ZN(n22202) );
  INV_X1 U23899 ( .A(n22209), .ZN(n22201) );
  NAND2_X1 U23900 ( .A1(n22202), .A2(n22201), .ZN(n22203) );
  OAI211_X1 U23901 ( .C1(n22205), .C2(n22269), .A(n22204), .B(n22203), .ZN(
        n22206) );
  INV_X1 U23902 ( .A(n22206), .ZN(n22207) );
  OAI21_X1 U23903 ( .B1(n22276), .B2(n22208), .A(n22207), .ZN(P1_U2824) );
  NOR2_X1 U23904 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n22209), .ZN(n22221) );
  NAND2_X1 U23905 ( .A1(n22210), .A2(n22233), .ZN(n22231) );
  OAI22_X1 U23906 ( .A1(n22213), .A2(n22212), .B1(n22262), .B2(n22211), .ZN(
        n22214) );
  AOI211_X1 U23907 ( .C1(n22266), .C2(n22215), .A(n22223), .B(n22214), .ZN(
        n22220) );
  AOI22_X1 U23908 ( .A1(n22218), .A2(n22253), .B1(n22217), .B2(n22216), .ZN(
        n22219) );
  OAI211_X1 U23909 ( .C1(n22221), .C2(n22231), .A(n22220), .B(n22219), .ZN(
        P1_U2823) );
  NOR2_X1 U23910 ( .A1(n22257), .A2(n22222), .ZN(n22228) );
  AOI21_X1 U23911 ( .B1(n22264), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n22223), .ZN(n22225) );
  NAND2_X1 U23912 ( .A1(n22236), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n22224) );
  OAI211_X1 U23913 ( .C1(n22226), .C2(n22276), .A(n22225), .B(n22224), .ZN(
        n22227) );
  AOI211_X1 U23914 ( .C1(n22229), .C2(n22253), .A(n22228), .B(n22227), .ZN(
        n22230) );
  OAI221_X1 U23915 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n22233), .C1(n22232), 
        .C2(n22231), .A(n22230), .ZN(P1_U2822) );
  AOI21_X1 U23916 ( .B1(n22235), .B2(n22234), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n22243) );
  AOI22_X1 U23917 ( .A1(n22264), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n22236), .B2(P1_EBX_REG_20__SCAN_IN), .ZN(n22242) );
  OAI22_X1 U23918 ( .A1(n22238), .A2(n22269), .B1(n22276), .B2(n22237), .ZN(
        n22239) );
  AOI21_X1 U23919 ( .B1(n22240), .B2(n22266), .A(n22239), .ZN(n22241) );
  OAI211_X1 U23920 ( .C1(n22248), .C2(n22243), .A(n22242), .B(n22241), .ZN(
        P1_U2820) );
  NOR3_X1 U23921 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n22245), .A3(n22244), 
        .ZN(n22250) );
  OAI22_X1 U23922 ( .A1(n22248), .A2(n22247), .B1(n22262), .B2(n22246), .ZN(
        n22249) );
  AOI211_X1 U23923 ( .C1(n22264), .C2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n22250), .B(n22249), .ZN(n22256) );
  NOR2_X1 U23924 ( .A1(n22251), .A2(n22276), .ZN(n22252) );
  AOI21_X1 U23925 ( .B1(n22254), .B2(n22253), .A(n22252), .ZN(n22255) );
  OAI211_X1 U23926 ( .C1(n22258), .C2(n22257), .A(n22256), .B(n22255), .ZN(
        P1_U2819) );
  INV_X1 U23927 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n22272) );
  INV_X1 U23928 ( .A(n22259), .ZN(n22260) );
  OAI22_X1 U23929 ( .A1(n22262), .A2(n22261), .B1(n22272), .B2(n22260), .ZN(
        n22263) );
  AOI21_X1 U23930 ( .B1(n22264), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n22263), .ZN(n22268) );
  NAND2_X1 U23931 ( .A1(n22266), .A2(n22265), .ZN(n22267) );
  OAI211_X1 U23932 ( .C1(n22270), .C2(n22269), .A(n22268), .B(n22267), .ZN(
        n22271) );
  AOI21_X1 U23933 ( .B1(n22273), .B2(n22272), .A(n22271), .ZN(n22274) );
  OAI21_X1 U23934 ( .B1(n22276), .B2(n22275), .A(n22274), .ZN(P1_U2818) );
  OAI21_X1 U23935 ( .B1(n22279), .B2(n22278), .A(n22277), .ZN(P1_U2806) );
  AOI22_X1 U23936 ( .A1(n22417), .A2(n22281), .B1(n22280), .B2(n22434), .ZN(
        n22285) );
  INV_X1 U23937 ( .A(n22290), .ZN(n22282) );
  NOR2_X1 U23938 ( .A1(n22283), .A2(n22282), .ZN(n22295) );
  NOR2_X1 U23939 ( .A1(n22286), .A2(n22295), .ZN(n22284) );
  AOI22_X1 U23940 ( .A1(n22457), .A2(n22286), .B1(n22285), .B2(n22284), .ZN(
        P1_U3478) );
  NOR2_X1 U23941 ( .A1(n22330), .A2(n22287), .ZN(n22288) );
  AOI21_X1 U23942 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(n22288), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n22291) );
  OAI221_X1 U23943 ( .B1(n22291), .B2(n22290), .C1(n22291), .C2(n22293), .A(
        n22289), .ZN(P1_U3163) );
  OAI21_X1 U23944 ( .B1(n22293), .B2(n14188), .A(n22292), .ZN(P1_U3466) );
  NOR2_X1 U23945 ( .A1(n22295), .A2(n22294), .ZN(n22301) );
  NAND2_X1 U23946 ( .A1(n22297), .A2(n22296), .ZN(n22298) );
  AOI21_X1 U23947 ( .B1(n22299), .B2(n22298), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n22300) );
  OAI22_X1 U23948 ( .A1(n22303), .A2(n22302), .B1(n22301), .B2(n22300), .ZN(
        P1_U3161) );
  OAI21_X1 U23949 ( .B1(n22306), .B2(n22305), .A(n22304), .ZN(P1_U2805) );
  AOI21_X1 U23950 ( .B1(n22308), .B2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n22307), 
        .ZN(n22309) );
  INV_X1 U23951 ( .A(n22309), .ZN(P1_U3465) );
  OAI21_X1 U23952 ( .B1(n22313), .B2(n22310), .A(n22311), .ZN(P2_U2818) );
  OAI21_X1 U23953 ( .B1(n22313), .B2(n22312), .A(n22311), .ZN(P2_U3592) );
  INV_X1 U23954 ( .A(n22314), .ZN(n22316) );
  OAI21_X1 U23955 ( .B1(n22318), .B2(n22315), .A(n22316), .ZN(P3_U2636) );
  OAI21_X1 U23956 ( .B1(n22318), .B2(n22317), .A(n22316), .ZN(P3_U3281) );
  INV_X1 U23957 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22357) );
  AOI21_X1 U23958 ( .B1(HOLD), .B2(n22319), .A(n22357), .ZN(n22320) );
  AOI21_X1 U23959 ( .B1(n22367), .B2(P3_STATE_REG_1__SCAN_IN), .A(n22361), 
        .ZN(n22374) );
  AOI21_X1 U23960 ( .B1(n22364), .B2(NA), .A(n22356), .ZN(n22366) );
  OAI22_X1 U23961 ( .A1(n22321), .A2(n22320), .B1(n22374), .B2(n22366), .ZN(
        P3_U3029) );
  INV_X1 U23962 ( .A(NA), .ZN(n22348) );
  NAND4_X1 U23963 ( .A1(n22330), .A2(P1_STATE_REG_1__SCAN_IN), .A3(
        P1_REQUESTPENDING_REG_SCAN_IN), .A4(n22348), .ZN(n22328) );
  NOR2_X1 U23964 ( .A1(NA), .A2(n22322), .ZN(n22324) );
  INV_X1 U23965 ( .A(HOLD), .ZN(n22358) );
  OAI21_X1 U23966 ( .B1(n22329), .B2(n22358), .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n22333) );
  OAI211_X1 U23967 ( .C1(n22324), .C2(n22323), .A(HOLD), .B(n22333), .ZN(
        n22327) );
  AOI21_X1 U23968 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n22330), .A(n22335), 
        .ZN(n22337) );
  INV_X1 U23969 ( .A(n22337), .ZN(n22325) );
  OAI211_X1 U23970 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n22348), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n22325), .ZN(n22326) );
  OAI221_X1 U23971 ( .B1(n22335), .B2(n22328), .C1(n22335), .C2(n22327), .A(
        n22326), .ZN(P1_U3196) );
  OAI221_X1 U23972 ( .B1(n22330), .B2(HOLD), .C1(n22330), .C2(n22329), .A(
        P1_STATE_REG_1__SCAN_IN), .ZN(n22332) );
  OAI211_X1 U23973 ( .C1(n22335), .C2(n22333), .A(n22332), .B(n22331), .ZN(
        P1_U3195) );
  NOR2_X1 U23974 ( .A1(n12943), .A2(n22358), .ZN(n22334) );
  AOI211_X1 U23975 ( .C1(NA), .C2(n22335), .A(n22334), .B(n22333), .ZN(n22336)
         );
  OAI22_X1 U23976 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n22337), .B1(n22805), 
        .B2(n22336), .ZN(P1_U3194) );
  NAND2_X1 U23977 ( .A1(n22338), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n22350) );
  NAND2_X1 U23978 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n22350), .ZN(n22349) );
  OAI22_X1 U23979 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n22348), .B1(n22339), 
        .B2(n22358), .ZN(n22340) );
  AOI22_X1 U23980 ( .A1(n22354), .A2(n22349), .B1(n22341), .B2(n22340), .ZN(
        n22342) );
  OAI21_X1 U23981 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(n22343), .A(n22342), .ZN(P2_U3209) );
  NAND2_X1 U23982 ( .A1(n22344), .A2(HOLD), .ZN(n22346) );
  OAI211_X1 U23983 ( .C1(n22354), .C2(n22358), .A(P2_STATE_REG_0__SCAN_IN), 
        .B(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22345) );
  NAND4_X1 U23984 ( .A1(n22347), .A2(n22346), .A3(n22350), .A4(n22345), .ZN(
        P2_U3210) );
  OAI22_X1 U23985 ( .A1(HOLD), .A2(n22349), .B1(P2_STATE_REG_0__SCAN_IN), .B2(
        n22348), .ZN(n22355) );
  OAI22_X1 U23986 ( .A1(NA), .A2(n22350), .B1(P2_STATE_REG_1__SCAN_IN), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22351) );
  OAI211_X1 U23987 ( .C1(HOLD), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n22351), .ZN(n22353) );
  OAI211_X1 U23988 ( .C1(n22355), .C2(n22354), .A(n22353), .B(n22352), .ZN(
        P2_U3211) );
  NOR2_X1 U23989 ( .A1(n22358), .A2(n22356), .ZN(n22371) );
  INV_X1 U23990 ( .A(n22371), .ZN(n22360) );
  OAI222_X1 U23991 ( .A1(n22361), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .B1(
        n22361), .B2(n22360), .C1(P3_STATE_REG_2__SCAN_IN), .C2(
        P3_STATE_REG_0__SCAN_IN), .ZN(n22365) );
  NAND2_X1 U23992 ( .A1(n22358), .A2(n22357), .ZN(n22369) );
  OAI221_X1 U23993 ( .B1(n22361), .B2(n22360), .C1(n22361), .C2(n22369), .A(
        n22359), .ZN(n22362) );
  AOI22_X1 U23994 ( .A1(n22365), .A2(n22364), .B1(n22363), .B2(n22362), .ZN(
        P3_U3030) );
  INV_X1 U23995 ( .A(n22366), .ZN(n22373) );
  NAND2_X1 U23996 ( .A1(n22367), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n22368) );
  OAI22_X1 U23997 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n22368), .ZN(n22370) );
  OAI211_X1 U23998 ( .C1(n22371), .C2(n22370), .A(P3_STATE_REG_0__SCAN_IN), 
        .B(n22369), .ZN(n22372) );
  OAI21_X1 U23999 ( .B1(n22374), .B2(n22373), .A(n22372), .ZN(P3_U3031) );
  AOI22_X1 U24000 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n22381), .B1(n22384), 
        .B2(P1_EAX_REG_9__SCAN_IN), .ZN(n22376) );
  NAND2_X1 U24001 ( .A1(n22376), .A2(n22375), .ZN(P1_U2961) );
  AOI22_X1 U24002 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n22385), .B1(n22384), 
        .B2(P1_EAX_REG_11__SCAN_IN), .ZN(n22378) );
  NAND2_X1 U24003 ( .A1(n22378), .A2(n22377), .ZN(P1_U2963) );
  AOI22_X1 U24004 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n22385), .B1(n22384), 
        .B2(P1_EAX_REG_12__SCAN_IN), .ZN(n22380) );
  NAND2_X1 U24005 ( .A1(n22380), .A2(n22379), .ZN(P1_U2964) );
  AOI22_X1 U24006 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n22381), .B1(n22384), 
        .B2(P1_EAX_REG_13__SCAN_IN), .ZN(n22383) );
  NAND2_X1 U24007 ( .A1(n22383), .A2(n22382), .ZN(P1_U2965) );
  AOI22_X1 U24008 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n22385), .B1(n22384), 
        .B2(P1_EAX_REG_14__SCAN_IN), .ZN(n22387) );
  NAND2_X1 U24009 ( .A1(n22387), .A2(n22386), .ZN(P1_U2966) );
  NOR3_X1 U24010 ( .A1(n22697), .A2(n22797), .A3(n22468), .ZN(n22388) );
  NOR2_X1 U24011 ( .A1(n22468), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22469) );
  NOR2_X1 U24012 ( .A1(n22388), .A2(n22469), .ZN(n22397) );
  INV_X1 U24013 ( .A(n22397), .ZN(n22390) );
  NAND2_X1 U24014 ( .A1(n22418), .A2(n11193), .ZN(n22389) );
  NOR2_X1 U24015 ( .A1(n14427), .A2(n22389), .ZN(n22396) );
  NAND2_X1 U24016 ( .A1(n22457), .A2(n22391), .ZN(n22683) );
  OAI22_X1 U24017 ( .A1(n22684), .A2(n22407), .B1(n22683), .B2(n22477), .ZN(
        n22392) );
  INV_X1 U24018 ( .A(n22392), .ZN(n22399) );
  INV_X1 U24019 ( .A(n22410), .ZN(n22460) );
  NOR2_X1 U24020 ( .A1(n22393), .A2(n22424), .ZN(n22394) );
  AOI211_X1 U24021 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n22683), .A(n22460), 
        .B(n22394), .ZN(n22395) );
  OAI21_X1 U24022 ( .B1(n22397), .B2(n22396), .A(n22395), .ZN(n22690) );
  AOI22_X1 U24023 ( .A1(n22690), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n22697), .B2(n22465), .ZN(n22398) );
  OAI211_X1 U24024 ( .C1(n22693), .C2(n22490), .A(n22399), .B(n22398), .ZN(
        P1_U3033) );
  NOR3_X1 U24025 ( .A1(n22703), .A2(n22709), .A3(n22468), .ZN(n22402) );
  NOR2_X1 U24026 ( .A1(n22402), .A2(n22469), .ZN(n22412) );
  INV_X1 U24027 ( .A(n22412), .ZN(n22405) );
  NAND2_X1 U24028 ( .A1(n22418), .A2(n22471), .ZN(n22403) );
  NOR2_X1 U24029 ( .A1(n14427), .A2(n22403), .ZN(n22411) );
  NOR2_X1 U24030 ( .A1(n22404), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22439) );
  NOR3_X1 U24031 ( .A1(n22406), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22415) );
  NAND2_X1 U24032 ( .A1(n22457), .A2(n22415), .ZN(n22587) );
  OAI22_X1 U24033 ( .A1(n22701), .A2(n22407), .B1(n22587), .B2(n22477), .ZN(
        n22408) );
  INV_X1 U24034 ( .A(n22408), .ZN(n22414) );
  NOR2_X1 U24035 ( .A1(n22439), .A2(n22424), .ZN(n22445) );
  AOI21_X1 U24036 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22587), .A(n22445), 
        .ZN(n22409) );
  OAI211_X1 U24037 ( .C1(n22412), .C2(n22411), .A(n22410), .B(n22409), .ZN(
        n22704) );
  AOI22_X1 U24038 ( .A1(n22704), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n22709), .B2(n22465), .ZN(n22413) );
  OAI211_X1 U24039 ( .C1(n22707), .C2(n22490), .A(n22414), .B(n22413), .ZN(
        P1_U3049) );
  INV_X1 U24040 ( .A(n22415), .ZN(n22428) );
  NAND3_X1 U24041 ( .A1(n22418), .A2(n22417), .A3(n22416), .ZN(n22419) );
  OR2_X1 U24042 ( .A1(n22419), .A2(n14427), .ZN(n22421) );
  NOR2_X1 U24043 ( .A1(n22457), .A2(n22428), .ZN(n22708) );
  INV_X1 U24044 ( .A(n22708), .ZN(n22420) );
  AND2_X1 U24045 ( .A1(n22421), .A2(n22420), .ZN(n22426) );
  OAI21_X1 U24046 ( .B1(n22423), .B2(n22422), .A(n22434), .ZN(n22431) );
  OAI22_X1 U24047 ( .A1(n22424), .A2(n22428), .B1(n22426), .B2(n22431), .ZN(
        n22425) );
  AOI22_X1 U24048 ( .A1(n22717), .A2(n22465), .B1(n22708), .B2(n22458), .ZN(
        n22433) );
  INV_X1 U24049 ( .A(n22426), .ZN(n22430) );
  AOI21_X1 U24050 ( .B1(n22468), .B2(n22428), .A(n22427), .ZN(n22429) );
  OAI21_X1 U24051 ( .B1(n22431), .B2(n22430), .A(n22429), .ZN(n22710) );
  AOI22_X1 U24052 ( .A1(n22710), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n22709), .B2(n22487), .ZN(n22432) );
  OAI211_X1 U24053 ( .C1(n22713), .C2(n22490), .A(n22433), .B(n22432), .ZN(
        P1_U3057) );
  INV_X1 U24054 ( .A(n22730), .ZN(n22435) );
  NAND3_X1 U24055 ( .A1(n22435), .A2(n22434), .A3(n22728), .ZN(n22437) );
  INV_X1 U24056 ( .A(n22469), .ZN(n22436) );
  NAND2_X1 U24057 ( .A1(n22437), .A2(n22436), .ZN(n22444) );
  NAND2_X1 U24058 ( .A1(n22438), .A2(n22471), .ZN(n22443) );
  INV_X1 U24059 ( .A(n22443), .ZN(n22440) );
  NOR3_X1 U24060 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n22441), .ZN(n22664) );
  INV_X1 U24061 ( .A(n22664), .ZN(n22727) );
  OAI22_X1 U24062 ( .A1(n22728), .A2(n22478), .B1(n22727), .B2(n22477), .ZN(
        n22442) );
  INV_X1 U24063 ( .A(n22442), .ZN(n22450) );
  NAND2_X1 U24064 ( .A1(n22444), .A2(n22443), .ZN(n22448) );
  INV_X1 U24065 ( .A(n22480), .ZN(n22446) );
  NOR2_X1 U24066 ( .A1(n22446), .A2(n22445), .ZN(n22447) );
  OAI211_X1 U24067 ( .C1(n14188), .C2(n22664), .A(n22448), .B(n22447), .ZN(
        n22731) );
  AOI22_X1 U24068 ( .A1(n22731), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n22730), .B2(n22487), .ZN(n22449) );
  OAI211_X1 U24069 ( .C1(n22734), .C2(n22490), .A(n22450), .B(n22449), .ZN(
        P1_U3081) );
  NOR2_X1 U24070 ( .A1(n22758), .A2(n22468), .ZN(n22451) );
  AOI21_X1 U24071 ( .B1(n22451), .B2(n22768), .A(n22469), .ZN(n22464) );
  INV_X1 U24072 ( .A(n22464), .ZN(n22455) );
  AND2_X1 U24073 ( .A1(n22452), .A2(n22471), .ZN(n22463) );
  NAND2_X1 U24074 ( .A1(n22457), .A2(n22456), .ZN(n22756) );
  INV_X1 U24075 ( .A(n22756), .ZN(n22634) );
  AOI22_X1 U24076 ( .A1(n22758), .A2(n22487), .B1(n22634), .B2(n22458), .ZN(
        n22467) );
  INV_X1 U24077 ( .A(n22459), .ZN(n22461) );
  AOI211_X1 U24078 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n22756), .A(n22461), 
        .B(n22460), .ZN(n22462) );
  OAI21_X1 U24079 ( .B1(n22464), .B2(n22463), .A(n22462), .ZN(n22759) );
  INV_X1 U24080 ( .A(n22768), .ZN(n22635) );
  AOI22_X1 U24081 ( .A1(n22759), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n22635), .B2(n22465), .ZN(n22466) );
  OAI211_X1 U24082 ( .C1(n22762), .C2(n22490), .A(n22467), .B(n22466), .ZN(
        P1_U3113) );
  NOR2_X1 U24083 ( .A1(n22772), .A2(n22468), .ZN(n22470) );
  AOI21_X1 U24084 ( .B1(n22470), .B2(n22783), .A(n22469), .ZN(n22486) );
  INV_X1 U24085 ( .A(n22486), .ZN(n22475) );
  NOR2_X1 U24086 ( .A1(n22472), .A2(n22471), .ZN(n22485) );
  NOR2_X1 U24087 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22476), .ZN(
        n22481) );
  INV_X1 U24088 ( .A(n22481), .ZN(n22770) );
  OAI22_X1 U24089 ( .A1(n22783), .A2(n22478), .B1(n22770), .B2(n22477), .ZN(
        n22479) );
  INV_X1 U24090 ( .A(n22479), .ZN(n22489) );
  OAI21_X1 U24091 ( .B1(n14188), .B2(n22481), .A(n22480), .ZN(n22482) );
  AOI21_X1 U24092 ( .B1(n22483), .B2(P1_STATE2_REG_2__SCAN_IN), .A(n22482), 
        .ZN(n22484) );
  OAI21_X1 U24093 ( .B1(n22486), .B2(n22485), .A(n22484), .ZN(n22773) );
  AOI22_X1 U24094 ( .A1(n22773), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n22772), .B2(n22487), .ZN(n22488) );
  OAI211_X1 U24095 ( .C1(n22777), .C2(n22490), .A(n22489), .B(n22488), .ZN(
        P1_U3129) );
  OAI22_X1 U24096 ( .A1(n22684), .A2(n22528), .B1(n22513), .B2(n22683), .ZN(
        n22491) );
  INV_X1 U24097 ( .A(n22491), .ZN(n22493) );
  AOI22_X1 U24098 ( .A1(n22690), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n22697), .B2(n22525), .ZN(n22492) );
  OAI211_X1 U24099 ( .C1(n22693), .C2(n22519), .A(n22493), .B(n22492), .ZN(
        P1_U3034) );
  OAI22_X1 U24100 ( .A1(n22701), .A2(n22528), .B1(n22513), .B2(n22587), .ZN(
        n22494) );
  INV_X1 U24101 ( .A(n22494), .ZN(n22496) );
  AOI22_X1 U24102 ( .A1(n22704), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n22709), .B2(n22525), .ZN(n22495) );
  OAI211_X1 U24103 ( .C1(n22707), .C2(n22519), .A(n22496), .B(n22495), .ZN(
        P1_U3050) );
  AOI22_X1 U24104 ( .A1(n22709), .A2(n22516), .B1(n22523), .B2(n22708), .ZN(
        n22498) );
  AOI22_X1 U24105 ( .A1(n22710), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n22717), .B2(n22525), .ZN(n22497) );
  OAI211_X1 U24106 ( .C1(n22713), .C2(n22519), .A(n22498), .B(n22497), .ZN(
        P1_U3058) );
  INV_X1 U24107 ( .A(n22499), .ZN(n22722) );
  AOI22_X1 U24108 ( .A1(n22722), .A2(n22524), .B1(n22523), .B2(n22721), .ZN(
        n22501) );
  AOI22_X1 U24109 ( .A1(n22723), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n22730), .B2(n22525), .ZN(n22500) );
  OAI211_X1 U24110 ( .C1(n22528), .C2(n22726), .A(n22501), .B(n22500), .ZN(
        P1_U3074) );
  AOI22_X1 U24111 ( .A1(n22730), .A2(n22516), .B1(n22523), .B2(n22664), .ZN(
        n22503) );
  AOI22_X1 U24112 ( .A1(n22731), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n22738), .B2(n22525), .ZN(n22502) );
  OAI211_X1 U24113 ( .C1(n22734), .C2(n22519), .A(n22503), .B(n22502), .ZN(
        P1_U3082) );
  INV_X1 U24114 ( .A(n22504), .ZN(n22751) );
  AOI22_X1 U24115 ( .A1(n22751), .A2(n22524), .B1(n22523), .B2(n22750), .ZN(
        n22506) );
  AOI22_X1 U24116 ( .A1(n22752), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n22758), .B2(n22525), .ZN(n22505) );
  OAI211_X1 U24117 ( .C1(n22528), .C2(n22755), .A(n22506), .B(n22505), .ZN(
        P1_U3106) );
  OAI22_X1 U24118 ( .A1(n22768), .A2(n22514), .B1(n22756), .B2(n22513), .ZN(
        n22507) );
  INV_X1 U24119 ( .A(n22507), .ZN(n22509) );
  AOI22_X1 U24120 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n22759), .B1(
        n22758), .B2(n22516), .ZN(n22508) );
  OAI211_X1 U24121 ( .C1(n22762), .C2(n22519), .A(n22509), .B(n22508), .ZN(
        P1_U3114) );
  INV_X1 U24122 ( .A(n22510), .ZN(n22764) );
  AOI22_X1 U24123 ( .A1(n22764), .A2(n22524), .B1(n22523), .B2(n22763), .ZN(
        n22512) );
  AOI22_X1 U24124 ( .A1(n22765), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n22772), .B2(n22525), .ZN(n22511) );
  OAI211_X1 U24125 ( .C1(n22528), .C2(n22768), .A(n22512), .B(n22511), .ZN(
        P1_U3122) );
  OAI22_X1 U24126 ( .A1(n22783), .A2(n22514), .B1(n22770), .B2(n22513), .ZN(
        n22515) );
  INV_X1 U24127 ( .A(n22515), .ZN(n22518) );
  AOI22_X1 U24128 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n22773), .B1(
        n22772), .B2(n22516), .ZN(n22517) );
  OAI211_X1 U24129 ( .C1(n22777), .C2(n22519), .A(n22518), .B(n22517), .ZN(
        P1_U3130) );
  INV_X1 U24130 ( .A(n22520), .ZN(n22779) );
  AOI22_X1 U24131 ( .A1(n22779), .A2(n22524), .B1(n22523), .B2(n22778), .ZN(
        n22522) );
  AOI22_X1 U24132 ( .A1(n22780), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n22787), .B2(n22525), .ZN(n22521) );
  OAI211_X1 U24133 ( .C1(n22528), .C2(n22783), .A(n22522), .B(n22521), .ZN(
        P1_U3138) );
  AOI22_X1 U24134 ( .A1(n22795), .A2(n22524), .B1(n22523), .B2(n22793), .ZN(
        n22527) );
  AOI22_X1 U24135 ( .A1(n22798), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n22797), .B2(n22525), .ZN(n22526) );
  OAI211_X1 U24136 ( .C1(n22528), .C2(n22801), .A(n22527), .B(n22526), .ZN(
        P1_U3154) );
  INV_X1 U24137 ( .A(n22549), .ZN(n22560) );
  OAI22_X1 U24138 ( .A1(n22684), .A2(n22560), .B1(n22546), .B2(n22683), .ZN(
        n22529) );
  INV_X1 U24139 ( .A(n22529), .ZN(n22531) );
  INV_X1 U24140 ( .A(n22547), .ZN(n22557) );
  AOI22_X1 U24141 ( .A1(n22690), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n22697), .B2(n22557), .ZN(n22530) );
  OAI211_X1 U24142 ( .C1(n22693), .C2(n22552), .A(n22531), .B(n22530), .ZN(
        P1_U3035) );
  INV_X1 U24143 ( .A(n22587), .ZN(n22702) );
  AOI22_X1 U24144 ( .A1(n22709), .A2(n22557), .B1(n22702), .B2(n22555), .ZN(
        n22533) );
  AOI22_X1 U24145 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n22704), .B1(
        n22703), .B2(n22549), .ZN(n22532) );
  OAI211_X1 U24146 ( .C1(n22707), .C2(n22552), .A(n22533), .B(n22532), .ZN(
        P1_U3051) );
  AOI22_X1 U24147 ( .A1(n22717), .A2(n22557), .B1(n22708), .B2(n22555), .ZN(
        n22535) );
  AOI22_X1 U24148 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n22710), .B1(
        n22709), .B2(n22549), .ZN(n22534) );
  OAI211_X1 U24149 ( .C1(n22713), .C2(n22552), .A(n22535), .B(n22534), .ZN(
        P1_U3059) );
  AOI22_X1 U24150 ( .A1(n22722), .A2(n22556), .B1(n22555), .B2(n22721), .ZN(
        n22537) );
  AOI22_X1 U24151 ( .A1(n22723), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n22730), .B2(n22557), .ZN(n22536) );
  OAI211_X1 U24152 ( .C1(n22560), .C2(n22726), .A(n22537), .B(n22536), .ZN(
        P1_U3075) );
  AOI22_X1 U24153 ( .A1(n22730), .A2(n22549), .B1(n22555), .B2(n22664), .ZN(
        n22539) );
  AOI22_X1 U24154 ( .A1(n22731), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n22738), .B2(n22557), .ZN(n22538) );
  OAI211_X1 U24155 ( .C1(n22734), .C2(n22552), .A(n22539), .B(n22538), .ZN(
        P1_U3083) );
  AOI22_X1 U24156 ( .A1(n22751), .A2(n22556), .B1(n22555), .B2(n22750), .ZN(
        n22541) );
  AOI22_X1 U24157 ( .A1(n22752), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n22758), .B2(n22557), .ZN(n22540) );
  OAI211_X1 U24158 ( .C1(n22560), .C2(n22755), .A(n22541), .B(n22540), .ZN(
        P1_U3107) );
  AOI22_X1 U24159 ( .A1(n22758), .A2(n22549), .B1(n22555), .B2(n22634), .ZN(
        n22543) );
  AOI22_X1 U24160 ( .A1(n22759), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n22635), .B2(n22557), .ZN(n22542) );
  OAI211_X1 U24161 ( .C1(n22762), .C2(n22552), .A(n22543), .B(n22542), .ZN(
        P1_U3115) );
  AOI22_X1 U24162 ( .A1(n22764), .A2(n22556), .B1(n22555), .B2(n22763), .ZN(
        n22545) );
  AOI22_X1 U24163 ( .A1(n22765), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n22772), .B2(n22557), .ZN(n22544) );
  OAI211_X1 U24164 ( .C1(n22560), .C2(n22768), .A(n22545), .B(n22544), .ZN(
        P1_U3123) );
  OAI22_X1 U24165 ( .A1(n22783), .A2(n22547), .B1(n22770), .B2(n22546), .ZN(
        n22548) );
  INV_X1 U24166 ( .A(n22548), .ZN(n22551) );
  AOI22_X1 U24167 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n22773), .B1(
        n22772), .B2(n22549), .ZN(n22550) );
  OAI211_X1 U24168 ( .C1(n22777), .C2(n22552), .A(n22551), .B(n22550), .ZN(
        P1_U3131) );
  AOI22_X1 U24169 ( .A1(n22779), .A2(n22556), .B1(n22555), .B2(n22778), .ZN(
        n22554) );
  AOI22_X1 U24170 ( .A1(n22780), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n22787), .B2(n22557), .ZN(n22553) );
  OAI211_X1 U24171 ( .C1(n22560), .C2(n22783), .A(n22554), .B(n22553), .ZN(
        P1_U3139) );
  AOI22_X1 U24172 ( .A1(n22795), .A2(n22556), .B1(n22555), .B2(n22793), .ZN(
        n22559) );
  AOI22_X1 U24173 ( .A1(n22798), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n22797), .B2(n22557), .ZN(n22558) );
  OAI211_X1 U24174 ( .C1(n22560), .C2(n22801), .A(n22559), .B(n22558), .ZN(
        P1_U3155) );
  OAI22_X1 U24175 ( .A1(n22684), .A2(n22564), .B1(n22683), .B2(n22577), .ZN(
        n22561) );
  INV_X1 U24176 ( .A(n22561), .ZN(n22563) );
  AOI22_X1 U24177 ( .A1(n22690), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n22697), .B2(n22571), .ZN(n22562) );
  OAI211_X1 U24178 ( .C1(n22693), .C2(n22583), .A(n22563), .B(n22562), .ZN(
        P1_U3036) );
  OAI22_X1 U24179 ( .A1(n22701), .A2(n22564), .B1(n22587), .B2(n22577), .ZN(
        n22565) );
  INV_X1 U24180 ( .A(n22565), .ZN(n22567) );
  AOI22_X1 U24181 ( .A1(n22704), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n22709), .B2(n22571), .ZN(n22566) );
  OAI211_X1 U24182 ( .C1(n22707), .C2(n22583), .A(n22567), .B(n22566), .ZN(
        P1_U3052) );
  AOI22_X1 U24183 ( .A1(n22717), .A2(n22571), .B1(n22708), .B2(n22570), .ZN(
        n22569) );
  AOI22_X1 U24184 ( .A1(n22710), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n22709), .B2(n22580), .ZN(n22568) );
  OAI211_X1 U24185 ( .C1(n22713), .C2(n22583), .A(n22569), .B(n22568), .ZN(
        P1_U3060) );
  AOI22_X1 U24186 ( .A1(n22730), .A2(n22580), .B1(n22664), .B2(n22570), .ZN(
        n22573) );
  AOI22_X1 U24187 ( .A1(n22731), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n22738), .B2(n22571), .ZN(n22572) );
  OAI211_X1 U24188 ( .C1(n22734), .C2(n22583), .A(n22573), .B(n22572), .ZN(
        P1_U3084) );
  OAI22_X1 U24189 ( .A1(n22768), .A2(n22578), .B1(n22756), .B2(n22577), .ZN(
        n22574) );
  INV_X1 U24190 ( .A(n22574), .ZN(n22576) );
  AOI22_X1 U24191 ( .A1(n22759), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n22758), .B2(n22580), .ZN(n22575) );
  OAI211_X1 U24192 ( .C1(n22762), .C2(n22583), .A(n22576), .B(n22575), .ZN(
        P1_U3116) );
  OAI22_X1 U24193 ( .A1(n22783), .A2(n22578), .B1(n22770), .B2(n22577), .ZN(
        n22579) );
  INV_X1 U24194 ( .A(n22579), .ZN(n22582) );
  AOI22_X1 U24195 ( .A1(n22773), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n22772), .B2(n22580), .ZN(n22581) );
  OAI211_X1 U24196 ( .C1(n22777), .C2(n22583), .A(n22582), .B(n22581), .ZN(
        P1_U3132) );
  OAI22_X1 U24197 ( .A1(n22684), .A2(n22619), .B1(n22605), .B2(n22683), .ZN(
        n22584) );
  INV_X1 U24198 ( .A(n22584), .ZN(n22586) );
  AOI22_X1 U24199 ( .A1(n22690), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n22697), .B2(n22616), .ZN(n22585) );
  OAI211_X1 U24200 ( .C1(n22693), .C2(n22611), .A(n22586), .B(n22585), .ZN(
        P1_U3037) );
  OAI22_X1 U24201 ( .A1(n22701), .A2(n22619), .B1(n22605), .B2(n22587), .ZN(
        n22588) );
  INV_X1 U24202 ( .A(n22588), .ZN(n22590) );
  AOI22_X1 U24203 ( .A1(n22704), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n22709), .B2(n22616), .ZN(n22589) );
  OAI211_X1 U24204 ( .C1(n22707), .C2(n22611), .A(n22590), .B(n22589), .ZN(
        P1_U3053) );
  AOI22_X1 U24205 ( .A1(n22709), .A2(n22608), .B1(n22614), .B2(n22708), .ZN(
        n22592) );
  AOI22_X1 U24206 ( .A1(n22710), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n22717), .B2(n22616), .ZN(n22591) );
  OAI211_X1 U24207 ( .C1(n22713), .C2(n22611), .A(n22592), .B(n22591), .ZN(
        P1_U3061) );
  AOI22_X1 U24208 ( .A1(n22722), .A2(n22615), .B1(n22614), .B2(n22721), .ZN(
        n22594) );
  AOI22_X1 U24209 ( .A1(n22723), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n22730), .B2(n22616), .ZN(n22593) );
  OAI211_X1 U24210 ( .C1(n22619), .C2(n22726), .A(n22594), .B(n22593), .ZN(
        P1_U3077) );
  OAI22_X1 U24211 ( .A1(n22728), .A2(n22606), .B1(n22727), .B2(n22605), .ZN(
        n22595) );
  INV_X1 U24212 ( .A(n22595), .ZN(n22597) );
  AOI22_X1 U24213 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n22731), .B1(
        n22730), .B2(n22608), .ZN(n22596) );
  OAI211_X1 U24214 ( .C1(n22734), .C2(n22611), .A(n22597), .B(n22596), .ZN(
        P1_U3085) );
  AOI22_X1 U24215 ( .A1(n22751), .A2(n22615), .B1(n22614), .B2(n22750), .ZN(
        n22599) );
  AOI22_X1 U24216 ( .A1(n22752), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n22758), .B2(n22616), .ZN(n22598) );
  OAI211_X1 U24217 ( .C1(n22619), .C2(n22755), .A(n22599), .B(n22598), .ZN(
        P1_U3109) );
  OAI22_X1 U24218 ( .A1(n22768), .A2(n22606), .B1(n22756), .B2(n22605), .ZN(
        n22600) );
  INV_X1 U24219 ( .A(n22600), .ZN(n22602) );
  AOI22_X1 U24220 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n22759), .B1(
        n22758), .B2(n22608), .ZN(n22601) );
  OAI211_X1 U24221 ( .C1(n22762), .C2(n22611), .A(n22602), .B(n22601), .ZN(
        P1_U3117) );
  AOI22_X1 U24222 ( .A1(n22764), .A2(n22615), .B1(n22614), .B2(n22763), .ZN(
        n22604) );
  AOI22_X1 U24223 ( .A1(n22765), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n22772), .B2(n22616), .ZN(n22603) );
  OAI211_X1 U24224 ( .C1(n22619), .C2(n22768), .A(n22604), .B(n22603), .ZN(
        P1_U3125) );
  OAI22_X1 U24225 ( .A1(n22783), .A2(n22606), .B1(n22770), .B2(n22605), .ZN(
        n22607) );
  INV_X1 U24226 ( .A(n22607), .ZN(n22610) );
  AOI22_X1 U24227 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n22773), .B1(
        n22772), .B2(n22608), .ZN(n22609) );
  OAI211_X1 U24228 ( .C1(n22777), .C2(n22611), .A(n22610), .B(n22609), .ZN(
        P1_U3133) );
  AOI22_X1 U24229 ( .A1(n22779), .A2(n22615), .B1(n22614), .B2(n22778), .ZN(
        n22613) );
  AOI22_X1 U24230 ( .A1(n22780), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n22787), .B2(n22616), .ZN(n22612) );
  OAI211_X1 U24231 ( .C1(n22619), .C2(n22783), .A(n22613), .B(n22612), .ZN(
        P1_U3141) );
  AOI22_X1 U24232 ( .A1(n22795), .A2(n22615), .B1(n22614), .B2(n22793), .ZN(
        n22618) );
  AOI22_X1 U24233 ( .A1(n22798), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n22797), .B2(n22616), .ZN(n22617) );
  OAI211_X1 U24234 ( .C1(n22619), .C2(n22801), .A(n22618), .B(n22617), .ZN(
        P1_U3157) );
  INV_X1 U24235 ( .A(n22643), .ZN(n22654) );
  OAI22_X1 U24236 ( .A1(n22684), .A2(n22654), .B1(n22640), .B2(n22683), .ZN(
        n22620) );
  INV_X1 U24237 ( .A(n22620), .ZN(n22622) );
  INV_X1 U24238 ( .A(n22641), .ZN(n22651) );
  AOI22_X1 U24239 ( .A1(n22690), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n22697), .B2(n22651), .ZN(n22621) );
  OAI211_X1 U24240 ( .C1(n22693), .C2(n22646), .A(n22622), .B(n22621), .ZN(
        P1_U3038) );
  AOI22_X1 U24241 ( .A1(n22709), .A2(n22651), .B1(n22702), .B2(n22649), .ZN(
        n22624) );
  AOI22_X1 U24242 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n22704), .B1(
        n22703), .B2(n22643), .ZN(n22623) );
  OAI211_X1 U24243 ( .C1(n22707), .C2(n22646), .A(n22624), .B(n22623), .ZN(
        P1_U3054) );
  AOI22_X1 U24244 ( .A1(n22709), .A2(n22643), .B1(n22649), .B2(n22708), .ZN(
        n22626) );
  AOI22_X1 U24245 ( .A1(n22710), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n22717), .B2(n22651), .ZN(n22625) );
  OAI211_X1 U24246 ( .C1(n22713), .C2(n22646), .A(n22626), .B(n22625), .ZN(
        P1_U3062) );
  AOI22_X1 U24247 ( .A1(n22722), .A2(n22650), .B1(n22649), .B2(n22721), .ZN(
        n22628) );
  AOI22_X1 U24248 ( .A1(n22723), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n22730), .B2(n22651), .ZN(n22627) );
  OAI211_X1 U24249 ( .C1(n22654), .C2(n22726), .A(n22628), .B(n22627), .ZN(
        P1_U3078) );
  OAI22_X1 U24250 ( .A1(n22728), .A2(n22641), .B1(n22727), .B2(n22640), .ZN(
        n22629) );
  INV_X1 U24251 ( .A(n22629), .ZN(n22631) );
  AOI22_X1 U24252 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n22731), .B1(
        n22730), .B2(n22643), .ZN(n22630) );
  OAI211_X1 U24253 ( .C1(n22734), .C2(n22646), .A(n22631), .B(n22630), .ZN(
        P1_U3086) );
  AOI22_X1 U24254 ( .A1(n22751), .A2(n22650), .B1(n22649), .B2(n22750), .ZN(
        n22633) );
  AOI22_X1 U24255 ( .A1(n22752), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n22758), .B2(n22651), .ZN(n22632) );
  OAI211_X1 U24256 ( .C1(n22654), .C2(n22755), .A(n22633), .B(n22632), .ZN(
        P1_U3110) );
  AOI22_X1 U24257 ( .A1(n22758), .A2(n22643), .B1(n22649), .B2(n22634), .ZN(
        n22637) );
  AOI22_X1 U24258 ( .A1(n22759), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n22635), .B2(n22651), .ZN(n22636) );
  OAI211_X1 U24259 ( .C1(n22762), .C2(n22646), .A(n22637), .B(n22636), .ZN(
        P1_U3118) );
  AOI22_X1 U24260 ( .A1(n22764), .A2(n22650), .B1(n22649), .B2(n22763), .ZN(
        n22639) );
  AOI22_X1 U24261 ( .A1(n22765), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n22772), .B2(n22651), .ZN(n22638) );
  OAI211_X1 U24262 ( .C1(n22654), .C2(n22768), .A(n22639), .B(n22638), .ZN(
        P1_U3126) );
  OAI22_X1 U24263 ( .A1(n22783), .A2(n22641), .B1(n22770), .B2(n22640), .ZN(
        n22642) );
  INV_X1 U24264 ( .A(n22642), .ZN(n22645) );
  AOI22_X1 U24265 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n22773), .B1(
        n22772), .B2(n22643), .ZN(n22644) );
  OAI211_X1 U24266 ( .C1(n22777), .C2(n22646), .A(n22645), .B(n22644), .ZN(
        P1_U3134) );
  AOI22_X1 U24267 ( .A1(n22779), .A2(n22650), .B1(n22649), .B2(n22778), .ZN(
        n22648) );
  AOI22_X1 U24268 ( .A1(n22780), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n22787), .B2(n22651), .ZN(n22647) );
  OAI211_X1 U24269 ( .C1(n22654), .C2(n22783), .A(n22648), .B(n22647), .ZN(
        P1_U3142) );
  AOI22_X1 U24270 ( .A1(n22795), .A2(n22650), .B1(n22649), .B2(n22793), .ZN(
        n22653) );
  AOI22_X1 U24271 ( .A1(n22798), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n22797), .B2(n22651), .ZN(n22652) );
  OAI211_X1 U24272 ( .C1(n22654), .C2(n22801), .A(n22653), .B(n22652), .ZN(
        P1_U3158) );
  OAI22_X1 U24273 ( .A1(n22684), .A2(n22655), .B1(n22683), .B2(n22671), .ZN(
        n22656) );
  INV_X1 U24274 ( .A(n22656), .ZN(n22658) );
  AOI22_X1 U24275 ( .A1(n22690), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n22697), .B2(n22665), .ZN(n22657) );
  OAI211_X1 U24276 ( .C1(n22693), .C2(n22677), .A(n22658), .B(n22657), .ZN(
        P1_U3039) );
  AOI22_X1 U24277 ( .A1(n22709), .A2(n22665), .B1(n22702), .B2(n22663), .ZN(
        n22660) );
  AOI22_X1 U24278 ( .A1(n22704), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n22703), .B2(n22674), .ZN(n22659) );
  OAI211_X1 U24279 ( .C1(n22707), .C2(n22677), .A(n22660), .B(n22659), .ZN(
        P1_U3055) );
  AOI22_X1 U24280 ( .A1(n22717), .A2(n22665), .B1(n22708), .B2(n22663), .ZN(
        n22662) );
  AOI22_X1 U24281 ( .A1(n22710), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n22709), .B2(n22674), .ZN(n22661) );
  OAI211_X1 U24282 ( .C1(n22713), .C2(n22677), .A(n22662), .B(n22661), .ZN(
        P1_U3063) );
  AOI22_X1 U24283 ( .A1(n22730), .A2(n22674), .B1(n22664), .B2(n22663), .ZN(
        n22667) );
  AOI22_X1 U24284 ( .A1(n22731), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n22738), .B2(n22665), .ZN(n22666) );
  OAI211_X1 U24285 ( .C1(n22734), .C2(n22677), .A(n22667), .B(n22666), .ZN(
        P1_U3087) );
  OAI22_X1 U24286 ( .A1(n22768), .A2(n22672), .B1(n22756), .B2(n22671), .ZN(
        n22668) );
  INV_X1 U24287 ( .A(n22668), .ZN(n22670) );
  AOI22_X1 U24288 ( .A1(n22759), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n22758), .B2(n22674), .ZN(n22669) );
  OAI211_X1 U24289 ( .C1(n22762), .C2(n22677), .A(n22670), .B(n22669), .ZN(
        P1_U3119) );
  OAI22_X1 U24290 ( .A1(n22783), .A2(n22672), .B1(n22770), .B2(n22671), .ZN(
        n22673) );
  INV_X1 U24291 ( .A(n22673), .ZN(n22676) );
  AOI22_X1 U24292 ( .A1(n22773), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n22772), .B2(n22674), .ZN(n22675) );
  OAI211_X1 U24293 ( .C1(n22777), .C2(n22677), .A(n22676), .B(n22675), .ZN(
        P1_U3135) );
  NOR2_X1 U24294 ( .A1(n22679), .A2(n22678), .ZN(n22794) );
  INV_X1 U24295 ( .A(n22794), .ZN(n22776) );
  INV_X1 U24296 ( .A(DATAI_31_), .ZN(n22681) );
  INV_X1 U24297 ( .A(n22786), .ZN(n22802) );
  NAND2_X1 U24298 ( .A1(n12941), .A2(n22682), .ZN(n22769) );
  OAI22_X1 U24299 ( .A1(n22684), .A2(n22802), .B1(n22769), .B2(n22683), .ZN(
        n22685) );
  INV_X1 U24300 ( .A(n22685), .ZN(n22692) );
  INV_X1 U24301 ( .A(DATAI_23_), .ZN(n22689) );
  OAI22_X1 U24302 ( .A1(n22689), .A2(n22688), .B1(n22687), .B2(n22686), .ZN(
        n22796) );
  AOI22_X1 U24303 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n22690), .B1(
        n22697), .B2(n22796), .ZN(n22691) );
  OAI211_X1 U24304 ( .C1(n22693), .C2(n22776), .A(n22692), .B(n22691), .ZN(
        P1_U3040) );
  INV_X1 U24305 ( .A(n22796), .ZN(n22791) );
  INV_X1 U24306 ( .A(n22694), .ZN(n22696) );
  AOI22_X1 U24307 ( .A1(n22696), .A2(n22794), .B1(n22695), .B2(n22792), .ZN(
        n22700) );
  AOI22_X1 U24308 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n22698), .B1(
        n22697), .B2(n22786), .ZN(n22699) );
  OAI211_X1 U24309 ( .C1(n22791), .C2(n22701), .A(n22700), .B(n22699), .ZN(
        P1_U3048) );
  AOI22_X1 U24310 ( .A1(n22709), .A2(n22796), .B1(n22792), .B2(n22702), .ZN(
        n22706) );
  AOI22_X1 U24311 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n22704), .B1(
        n22703), .B2(n22786), .ZN(n22705) );
  OAI211_X1 U24312 ( .C1(n22707), .C2(n22776), .A(n22706), .B(n22705), .ZN(
        P1_U3056) );
  AOI22_X1 U24313 ( .A1(n22717), .A2(n22796), .B1(n22792), .B2(n22708), .ZN(
        n22712) );
  AOI22_X1 U24314 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n22710), .B1(
        n22709), .B2(n22786), .ZN(n22711) );
  OAI211_X1 U24315 ( .C1(n22713), .C2(n22776), .A(n22712), .B(n22711), .ZN(
        P1_U3064) );
  INV_X1 U24316 ( .A(n22714), .ZN(n22716) );
  AOI22_X1 U24317 ( .A1(n22716), .A2(n22794), .B1(n22715), .B2(n22792), .ZN(
        n22720) );
  AOI22_X1 U24318 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n22718), .B1(
        n22717), .B2(n22786), .ZN(n22719) );
  OAI211_X1 U24319 ( .C1(n22791), .C2(n22726), .A(n22720), .B(n22719), .ZN(
        P1_U3072) );
  AOI22_X1 U24320 ( .A1(n22722), .A2(n22794), .B1(n22721), .B2(n22792), .ZN(
        n22725) );
  AOI22_X1 U24321 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n22723), .B1(
        n22730), .B2(n22796), .ZN(n22724) );
  OAI211_X1 U24322 ( .C1(n22802), .C2(n22726), .A(n22725), .B(n22724), .ZN(
        P1_U3080) );
  OAI22_X1 U24323 ( .A1(n22728), .A2(n22791), .B1(n22769), .B2(n22727), .ZN(
        n22729) );
  INV_X1 U24324 ( .A(n22729), .ZN(n22733) );
  AOI22_X1 U24325 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n22731), .B1(
        n22730), .B2(n22786), .ZN(n22732) );
  OAI211_X1 U24326 ( .C1(n22734), .C2(n22776), .A(n22733), .B(n22732), .ZN(
        P1_U3088) );
  INV_X1 U24327 ( .A(n22735), .ZN(n22736) );
  AOI22_X1 U24328 ( .A1(n22737), .A2(n22794), .B1(n22736), .B2(n22792), .ZN(
        n22741) );
  AOI22_X1 U24329 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n22739), .B1(
        n22738), .B2(n22786), .ZN(n22740) );
  OAI211_X1 U24330 ( .C1(n22791), .C2(n22742), .A(n22741), .B(n22740), .ZN(
        P1_U3096) );
  INV_X1 U24331 ( .A(n22743), .ZN(n22745) );
  AOI22_X1 U24332 ( .A1(n22745), .A2(n22794), .B1(n22744), .B2(n22792), .ZN(
        n22749) );
  AOI22_X1 U24333 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n22747), .B1(
        n22746), .B2(n22786), .ZN(n22748) );
  OAI211_X1 U24334 ( .C1(n22791), .C2(n22755), .A(n22749), .B(n22748), .ZN(
        P1_U3104) );
  AOI22_X1 U24335 ( .A1(n22751), .A2(n22794), .B1(n22750), .B2(n22792), .ZN(
        n22754) );
  AOI22_X1 U24336 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n22752), .B1(
        n22758), .B2(n22796), .ZN(n22753) );
  OAI211_X1 U24337 ( .C1(n22802), .C2(n22755), .A(n22754), .B(n22753), .ZN(
        P1_U3112) );
  OAI22_X1 U24338 ( .A1(n22768), .A2(n22791), .B1(n22769), .B2(n22756), .ZN(
        n22757) );
  INV_X1 U24339 ( .A(n22757), .ZN(n22761) );
  AOI22_X1 U24340 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n22759), .B1(
        n22758), .B2(n22786), .ZN(n22760) );
  OAI211_X1 U24341 ( .C1(n22762), .C2(n22776), .A(n22761), .B(n22760), .ZN(
        P1_U3120) );
  AOI22_X1 U24342 ( .A1(n22764), .A2(n22794), .B1(n22763), .B2(n22792), .ZN(
        n22767) );
  AOI22_X1 U24343 ( .A1(n22765), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n22772), .B2(n22796), .ZN(n22766) );
  OAI211_X1 U24344 ( .C1(n22802), .C2(n22768), .A(n22767), .B(n22766), .ZN(
        P1_U3128) );
  OAI22_X1 U24345 ( .A1(n22783), .A2(n22791), .B1(n22770), .B2(n22769), .ZN(
        n22771) );
  INV_X1 U24346 ( .A(n22771), .ZN(n22775) );
  AOI22_X1 U24347 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n22773), .B1(
        n22772), .B2(n22786), .ZN(n22774) );
  OAI211_X1 U24348 ( .C1(n22777), .C2(n22776), .A(n22775), .B(n22774), .ZN(
        P1_U3136) );
  AOI22_X1 U24349 ( .A1(n22779), .A2(n22794), .B1(n22778), .B2(n22792), .ZN(
        n22782) );
  AOI22_X1 U24350 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n22780), .B1(
        n22787), .B2(n22796), .ZN(n22781) );
  OAI211_X1 U24351 ( .C1(n22802), .C2(n22783), .A(n22782), .B(n22781), .ZN(
        P1_U3144) );
  AOI22_X1 U24352 ( .A1(n22785), .A2(n22794), .B1(n22784), .B2(n22792), .ZN(
        n22790) );
  AOI22_X1 U24353 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n22788), .B1(
        n22787), .B2(n22786), .ZN(n22789) );
  OAI211_X1 U24354 ( .C1(n22791), .C2(n22801), .A(n22790), .B(n22789), .ZN(
        P1_U3152) );
  AOI22_X1 U24355 ( .A1(n22795), .A2(n22794), .B1(n22793), .B2(n22792), .ZN(
        n22800) );
  AOI22_X1 U24356 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n22798), .B1(
        n22797), .B2(n22796), .ZN(n22799) );
  OAI211_X1 U24357 ( .C1(n22802), .C2(n22801), .A(n22800), .B(n22799), .ZN(
        P1_U3160) );
  INV_X1 U24358 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n22806) );
  AOI22_X1 U24359 ( .A1(n22805), .A2(n22806), .B1(n22804), .B2(n22803), .ZN(
        P1_U3486) );
  AOI21_X1 U24360 ( .B1(n22808), .B2(n22807), .A(n22806), .ZN(n22809) );
  OR3_X1 U24361 ( .A1(n22811), .A2(n22810), .A3(n22809), .ZN(P1_U2801) );
  NAND2_X1 U11639 ( .A1(n11162), .A2(n12941), .ZN(n12948) );
  INV_X1 U11522 ( .A(n12933), .ZN(n12957) );
  BUF_X2 U11316 ( .A(n18331), .Z(n11151) );
  NOR2_X2 U11638 ( .A1(n14797), .A2(n12886), .ZN(n12946) );
  AND2_X1 U14556 ( .A1(n12946), .A2(n12945), .ZN(n14421) );
  BUF_X2 U11256 ( .A(n12876), .Z(n11188) );
  CLKBUF_X1 U11257 ( .A(n11666), .Z(n20429) );
  CLKBUF_X2 U11271 ( .A(n13800), .Z(n11156) );
  CLKBUF_X1 U11281 ( .A(n13807), .Z(n18432) );
  INV_X2 U11283 ( .A(n16320), .ZN(n16385) );
  CLKBUF_X1 U11291 ( .A(n16833), .Z(n16834) );
  CLKBUF_X1 U11303 ( .A(n11661), .Z(n16136) );
  AND2_X1 U11317 ( .A1(n11743), .A2(n11742), .ZN(n12286) );
  INV_X1 U11361 ( .A(n16321), .ZN(n16320) );
  CLKBUF_X1 U11363 ( .A(n16744), .Z(n16757) );
  CLKBUF_X1 U11371 ( .A(n17004), .Z(n11165) );
  CLKBUF_X1 U11584 ( .A(n14461), .Z(n11193) );
  CLKBUF_X1 U12103 ( .A(n20860), .Z(n20890) );
  CLKBUF_X1 U12354 ( .A(n19476), .Z(n19811) );
  OR2_X1 U12382 ( .A1(n13725), .A2(n13724), .ZN(n22812) );
  INV_X2 U12807 ( .A(n20831), .ZN(n19015) );
endmodule

