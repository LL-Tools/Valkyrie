

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput63,
         keyinput62, keyinput61, keyinput60, keyinput59, keyinput58,
         keyinput57, keyinput56, keyinput55, keyinput54, keyinput53,
         keyinput52, keyinput51, keyinput50, keyinput49, keyinput48,
         keyinput47, keyinput46, keyinput45, keyinput44, keyinput43,
         keyinput42, keyinput41, keyinput40, keyinput39, keyinput38,
         keyinput37, keyinput36, keyinput35, keyinput34, keyinput33,
         keyinput32, keyinput31, keyinput30, keyinput29, keyinput28,
         keyinput27, keyinput26, keyinput25, keyinput24, keyinput23,
         keyinput22, keyinput21, keyinput20, keyinput19, keyinput18,
         keyinput17, keyinput16, keyinput15, keyinput14, keyinput13,
         keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, keyinput7,
         keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, keyinput1,
         keyinput0;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6431, n6432, n6436, n6437, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7688, n7689, n7690, n7691, n7692, n7693, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15339;

  AND2_X1 U7179 ( .A1(n12710), .A2(n9625), .ZN(n12685) );
  INV_X4 U7180 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NAND2_X2 U7181 ( .A1(n12052), .A2(n12051), .ZN(n13564) );
  NOR2_X1 U7182 ( .A1(n6911), .A2(n6910), .ZN(n13993) );
  INV_X4 U7183 ( .A(n13372), .ZN(n13460) );
  INV_X2 U7184 ( .A(n8800), .ZN(n8806) );
  INV_X1 U7185 ( .A(n12319), .ZN(n12274) );
  AND2_X4 U7186 ( .A1(n10282), .A2(n10281), .ZN(n12319) );
  AND2_X4 U7187 ( .A1(n10282), .A2(n10280), .ZN(n12333) );
  INV_X1 U7188 ( .A(n8076), .ZN(n9921) );
  CLKBUF_X2 U7189 ( .A(n9115), .Z(n9473) );
  CLKBUF_X2 U7190 ( .A(n9339), .Z(n6440) );
  INV_X4 U7192 ( .A(n8088), .ZN(n7750) );
  INV_X1 U7193 ( .A(n8645), .ZN(n8754) );
  INV_X1 U7194 ( .A(n8359), .ZN(n8745) );
  BUF_X1 U7195 ( .A(n9038), .Z(n9231) );
  NAND2_X1 U7197 ( .A1(n7556), .A2(n6820), .ZN(n13142) );
  NAND2_X2 U7198 ( .A1(n7103), .A2(n7728), .ZN(n11869) );
  AND2_X1 U7199 ( .A1(n8909), .A2(n8910), .ZN(n9051) );
  NAND2_X1 U7200 ( .A1(n15085), .A2(n9037), .ZN(n9525) );
  INV_X1 U7201 ( .A(n14963), .ZN(n12641) );
  OR2_X1 U7202 ( .A1(n12772), .A2(n12773), .ZN(n12770) );
  INV_X1 U7203 ( .A(n10398), .ZN(n9633) );
  INV_X1 U7205 ( .A(n9676), .ZN(n12990) );
  INV_X1 U7206 ( .A(n10487), .ZN(n12191) );
  INV_X1 U7209 ( .A(n7951), .ZN(n8076) );
  OAI22_X1 U7210 ( .A1(n12106), .A2(n10196), .B1(n11869), .B2(n11872), .ZN(
        n10650) );
  INV_X2 U7211 ( .A(n8779), .ZN(n8419) );
  NAND2_X1 U7212 ( .A1(n7824), .A2(n7823), .ZN(n11919) );
  XNOR2_X1 U7213 ( .A(n8361), .B(P1_IR_REG_2__SCAN_IN), .ZN(n10343) );
  AND4_X1 U7214 ( .A1(n6988), .A2(n9142), .A3(n9138), .A4(n9091), .ZN(n6431)
         );
  XNOR2_X2 U7215 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n14211) );
  OAI21_X1 U7216 ( .B1(n11172), .B2(n9559), .A(n9561), .ZN(n11227) );
  OAI211_X2 U7217 ( .C1(n12380), .C2(n12360), .A(n6767), .B(n6766), .ZN(n14079) );
  XNOR2_X2 U7218 ( .A(n7584), .B(n9836), .ZN(n7583) );
  AOI21_X1 U7220 ( .B1(n11013), .B2(n11012), .A(n7573), .ZN(n11112) );
  AOI21_X2 U7221 ( .B1(n11457), .B2(n12119), .A(n8238), .ZN(n11601) );
  OAI21_X2 U7222 ( .B1(n11278), .B2(n6476), .A(n7207), .ZN(n11457) );
  XNOR2_X2 U7223 ( .A(n7707), .B(n7706), .ZN(n8222) );
  INV_X1 U7224 ( .A(n6440), .ZN(n6432) );
  NAND2_X1 U7225 ( .A1(n9048), .A2(n9831), .ZN(n9339) );
  AOI21_X2 U7226 ( .B1(n12679), .B2(n12672), .A(n6514), .ZN(n12673) );
  XNOR2_X2 U7227 ( .A(n9033), .B(n9032), .ZN(n10422) );
  AOI21_X2 U7228 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n10295), .A(n10294), .ZN(
        n10298) );
  NOR2_X2 U7229 ( .A1(n14326), .A2(n14325), .ZN(n14324) );
  NOR2_X2 U7230 ( .A1(n13876), .A2(n13875), .ZN(n13878) );
  AND2_X4 U7231 ( .A1(n12950), .A2(n12952), .ZN(n9038) );
  OAI22_X2 U7232 ( .A1(n9158), .A2(n8930), .B1(P2_DATAO_REG_9__SCAN_IN), .B2(
        n15276), .ZN(n9170) );
  NOR2_X2 U7233 ( .A1(n13315), .A2(n13500), .ZN(n13305) );
  OAI21_X2 U7234 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n10055), .A(n10054), .ZN(
        n10181) );
  XNOR2_X2 U7235 ( .A(n9022), .B(P3_IR_REG_2__SCAN_IN), .ZN(n12569) );
  NOR2_X2 U7236 ( .A1(n10834), .A2(n12560), .ZN(n10914) );
  NOR2_X2 U7238 ( .A1(n11703), .A2(n11702), .ZN(n13861) );
  AOI21_X2 U7239 ( .B1(n11700), .B2(P1_REG1_REG_16__SCAN_IN), .A(n11699), .ZN(
        n11703) );
  OR2_X1 U7240 ( .A1(n13283), .A2(n13282), .ZN(n6838) );
  AND2_X1 U7241 ( .A1(n8118), .A2(n8117), .ZN(n13320) );
  NOR2_X1 U7242 ( .A1(n8671), .A2(n8670), .ZN(n8672) );
  NAND2_X1 U7243 ( .A1(n8665), .A2(n8664), .ZN(n14012) );
  NAND2_X1 U7244 ( .A1(n7995), .A2(n7994), .ZN(n11978) );
  NAND2_X1 U7245 ( .A1(n8602), .A2(n8601), .ZN(n14150) );
  NAND2_X1 U7246 ( .A1(n9535), .A2(n9531), .ZN(n7114) );
  NAND2_X1 U7247 ( .A1(n13143), .A2(n11862), .ZN(n10140) );
  INV_X1 U7248 ( .A(n10516), .ZN(n12557) );
  INV_X4 U7249 ( .A(n8349), .ZN(n8800) );
  INV_X2 U7250 ( .A(n10893), .ZN(n12555) );
  INV_X1 U7251 ( .A(n12558), .ZN(n15085) );
  CLKBUF_X2 U7252 ( .A(n7754), .Z(n8150) );
  INV_X1 U7254 ( .A(n10243), .ZN(n8883) );
  NAND2_X2 U7255 ( .A1(n8179), .A2(n13640), .ZN(n7742) );
  NAND2_X2 U7256 ( .A1(n8305), .A2(n14192), .ZN(n8779) );
  OAI21_X1 U7258 ( .B1(n8611), .B2(P1_IR_REG_18__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8318) );
  NAND2_X2 U7259 ( .A1(n8882), .A2(n14197), .ZN(n8343) );
  NAND2_X2 U7260 ( .A1(n12154), .A2(n14192), .ZN(n8788) );
  BUF_X1 U7261 ( .A(n9385), .Z(n6436) );
  AND3_X1 U7262 ( .A1(n8290), .A2(n7320), .A3(n7319), .ZN(n7280) );
  NAND2_X1 U7263 ( .A1(n7743), .A2(n7745), .ZN(n7759) );
  NOR2_X1 U7264 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n8284) );
  NOR2_X1 U7265 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n8285) );
  NOR2_X1 U7266 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n6861) );
  NOR2_X1 U7267 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n8872) );
  OAI21_X1 U7268 ( .B1(n13697), .B2(n6665), .A(n6663), .ZN(n13656) );
  AND2_X1 U7269 ( .A1(n7027), .A2(n6574), .ZN(n8860) );
  INV_X1 U7270 ( .A(n12405), .ZN(n14089) );
  AND2_X1 U7271 ( .A1(n6791), .A2(n6790), .ZN(n13567) );
  AOI21_X1 U7272 ( .B1(n14077), .B2(n14138), .A(n7225), .ZN(n14078) );
  NOR2_X1 U7273 ( .A1(n7371), .A2(n7373), .ZN(n7370) );
  AOI21_X1 U7274 ( .B1(n9395), .B2(n15089), .A(n9394), .ZN(n12431) );
  INV_X1 U7275 ( .A(n7515), .ZN(n7513) );
  NOR2_X2 U7276 ( .A1(n7227), .A2(n13909), .ZN(n13901) );
  NAND2_X1 U7277 ( .A1(n12401), .A2(n12400), .ZN(n12399) );
  NAND2_X1 U7278 ( .A1(n6902), .A2(n13664), .ZN(n13909) );
  NAND2_X1 U7279 ( .A1(n8819), .A2(n8818), .ZN(n8850) );
  AND2_X1 U7280 ( .A1(n7128), .A2(n6481), .ZN(n12676) );
  NAND2_X1 U7281 ( .A1(n6662), .A2(n13759), .ZN(n13665) );
  NAND2_X1 U7282 ( .A1(n8799), .A2(n8798), .ZN(n13900) );
  AOI22_X2 U7283 ( .A1(n13622), .A2(n7750), .B1(n12050), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n12422) );
  NAND2_X1 U7284 ( .A1(n6904), .A2(n6903), .ZN(n13922) );
  XNOR2_X1 U7285 ( .A(n8817), .B(n8816), .ZN(n13622) );
  NOR2_X1 U7286 ( .A1(n12658), .A2(n6992), .ZN(n12660) );
  INV_X1 U7287 ( .A(n13942), .ZN(n6904) );
  XNOR2_X1 U7288 ( .A(n8814), .B(n8796), .ZN(n12152) );
  OAI21_X1 U7289 ( .B1(n8814), .B2(n8813), .A(n8812), .ZN(n8817) );
  NAND2_X1 U7290 ( .A1(n13955), .A2(n12376), .ZN(n13936) );
  NAND2_X1 U7291 ( .A1(n8795), .A2(n8794), .ZN(n8814) );
  OR2_X1 U7292 ( .A1(n13489), .A2(n9793), .ZN(n8170) );
  OR2_X1 U7293 ( .A1(n13965), .A2(n13940), .ZN(n13942) );
  NAND2_X1 U7294 ( .A1(n8760), .A2(n8759), .ZN(n14082) );
  NAND2_X1 U7295 ( .A1(n7219), .A2(n13993), .ZN(n13965) );
  NAND2_X1 U7296 ( .A1(n13988), .A2(n6458), .ZN(n13973) );
  NOR2_X1 U7297 ( .A1(n6784), .A2(n8253), .ZN(n6783) );
  NAND2_X1 U7298 ( .A1(n8159), .A2(n8158), .ZN(n13489) );
  NAND2_X1 U7299 ( .A1(n8747), .A2(n8746), .ZN(n14087) );
  NAND2_X1 U7300 ( .A1(n8718), .A2(n8717), .ZN(n13940) );
  AND2_X1 U7301 ( .A1(n7220), .A2(n14112), .ZN(n7219) );
  AOI21_X1 U7302 ( .B1(n13365), .B2(n8252), .A(n6526), .ZN(n7218) );
  XNOR2_X1 U7303 ( .A(n8157), .B(n8156), .ZN(n14193) );
  NAND2_X1 U7304 ( .A1(n8131), .A2(n8130), .ZN(n13500) );
  NAND2_X1 U7305 ( .A1(n8733), .A2(n8732), .ZN(n13921) );
  AOI21_X1 U7306 ( .B1(n8674), .B2(n8673), .A(n8672), .ZN(n8685) );
  NAND2_X1 U7307 ( .A1(n6753), .A2(n12352), .ZN(n14006) );
  NAND2_X1 U7308 ( .A1(n8698), .A2(n8697), .ZN(n13964) );
  INV_X1 U7309 ( .A(n13348), .ZN(n13587) );
  INV_X1 U7310 ( .A(n8838), .ZN(n14112) );
  NAND2_X1 U7311 ( .A1(n13679), .A2(n12259), .ZN(n13737) );
  AND2_X1 U7312 ( .A1(n8090), .A2(n8089), .ZN(n13348) );
  NAND2_X1 U7313 ( .A1(n8300), .A2(n8299), .ZN(n8838) );
  NAND2_X1 U7314 ( .A1(n13676), .A2(n12254), .ZN(n13679) );
  NAND2_X1 U7315 ( .A1(n8071), .A2(n8070), .ZN(n13591) );
  NAND2_X1 U7316 ( .A1(n14206), .A2(n8343), .ZN(n14119) );
  XNOR2_X1 U7317 ( .A(n8676), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14206) );
  OR2_X1 U7318 ( .A1(n14020), .A2(n12350), .ZN(n14023) );
  OR2_X1 U7319 ( .A1(n8085), .A2(n7662), .ZN(n8087) );
  NAND2_X1 U7320 ( .A1(n13705), .A2(n6459), .ZN(n6658) );
  AND2_X1 U7321 ( .A1(n8057), .A2(n8056), .ZN(n13376) );
  INV_X1 U7322 ( .A(n13387), .ZN(n13603) );
  AND2_X1 U7323 ( .A1(n12230), .A2(n12233), .ZN(n7538) );
  NAND2_X1 U7324 ( .A1(n6933), .A2(n6931), .ZN(n12804) );
  NAND2_X1 U7325 ( .A1(n6786), .A2(n8041), .ZN(n13387) );
  NAND2_X1 U7326 ( .A1(n8658), .A2(n8657), .ZN(n14130) );
  XOR2_X1 U7327 ( .A(n14376), .B(n12648), .Z(n14373) );
  NAND2_X1 U7328 ( .A1(n12647), .A2(n15026), .ZN(n12648) );
  OAI21_X1 U7329 ( .B1(n13749), .B2(n6655), .A(n6653), .ZN(n12227) );
  XNOR2_X1 U7330 ( .A(n8039), .B(n8040), .ZN(n11360) );
  OAI21_X1 U7331 ( .B1(n8039), .B2(n7363), .A(n7656), .ZN(n8051) );
  NAND2_X1 U7332 ( .A1(n8026), .A2(n8025), .ZN(n13537) );
  NAND2_X1 U7333 ( .A1(n11458), .A2(n7922), .ZN(n11461) );
  NAND2_X1 U7334 ( .A1(n6924), .A2(n6506), .ZN(n11753) );
  NAND2_X1 U7335 ( .A1(n14348), .A2(n14347), .ZN(n14346) );
  NAND2_X1 U7336 ( .A1(n8639), .A2(n8638), .ZN(n12381) );
  NAND2_X1 U7337 ( .A1(n15009), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n15008) );
  AND2_X1 U7338 ( .A1(n8008), .A2(n8007), .ZN(n13422) );
  NAND2_X1 U7339 ( .A1(n8614), .A2(n8613), .ZN(n14144) );
  NOR2_X1 U7340 ( .A1(n15006), .A2(n12588), .ZN(n15025) );
  NAND2_X1 U7341 ( .A1(n7087), .A2(n6595), .ZN(n7656) );
  NAND2_X1 U7342 ( .A1(n11286), .A2(n11285), .ZN(n11284) );
  NAND2_X1 U7343 ( .A1(n8593), .A2(n8592), .ZN(n12232) );
  AOI21_X1 U7344 ( .B1(n11227), .B2(n9563), .A(n6921), .ZN(n7546) );
  AOI21_X1 U7345 ( .B1(n7520), .B2(n7519), .A(n7518), .ZN(n7517) );
  NAND2_X1 U7346 ( .A1(n8565), .A2(n8564), .ZN(n12222) );
  NAND2_X1 U7347 ( .A1(n7130), .A2(n9401), .ZN(n11172) );
  NAND2_X1 U7348 ( .A1(n11223), .A2(n11226), .ZN(n11222) );
  NAND2_X1 U7349 ( .A1(n7963), .A2(n7962), .ZN(n13617) );
  NOR2_X1 U7350 ( .A1(n14968), .A2(n12585), .ZN(n14987) );
  AND2_X1 U7351 ( .A1(n7946), .A2(n7945), .ZN(n11968) );
  NAND2_X1 U7352 ( .A1(n8553), .A2(n8552), .ZN(n12214) );
  NOR2_X1 U7353 ( .A1(n14330), .A2(n14292), .ZN(n14333) );
  NAND2_X1 U7354 ( .A1(n7911), .A2(n7910), .ZN(n11961) );
  NAND2_X1 U7355 ( .A1(n10877), .A2(n9128), .ZN(n11044) );
  NAND2_X1 U7356 ( .A1(n6641), .A2(n6639), .ZN(n9276) );
  NAND2_X1 U7357 ( .A1(n7897), .A2(n7896), .ZN(n11953) );
  AOI21_X1 U7358 ( .B1(n7526), .B2(n6448), .A(n7525), .ZN(n7524) );
  OAI21_X1 U7359 ( .B1(n7892), .B2(n6880), .A(n6877), .ZN(n7630) );
  NAND2_X1 U7360 ( .A1(n7864), .A2(n7863), .ZN(n13477) );
  NAND2_X1 U7361 ( .A1(n8495), .A2(n8494), .ZN(n14491) );
  NAND2_X1 U7362 ( .A1(n7616), .A2(n7615), .ZN(n7892) );
  NAND2_X1 U7363 ( .A1(n7843), .A2(n7842), .ZN(n11932) );
  AND2_X1 U7364 ( .A1(n15063), .A2(n9079), .ZN(n10892) );
  NAND2_X1 U7365 ( .A1(n13468), .A2(n8272), .ZN(n13463) );
  OAI21_X1 U7366 ( .B1(n10565), .B2(n10885), .A(n6477), .ZN(n6870) );
  INV_X2 U7367 ( .A(n15096), .ZN(n15075) );
  XNOR2_X1 U7368 ( .A(n10534), .B(n10533), .ZN(n10565) );
  AND2_X1 U7369 ( .A1(n9544), .A2(n9540), .ZN(n10890) );
  AOI21_X1 U7370 ( .B1(n7169), .B2(n7168), .A(n6531), .ZN(n10534) );
  NAND2_X1 U7371 ( .A1(n9527), .A2(n9530), .ZN(n15082) );
  NAND2_X1 U7372 ( .A1(n7771), .A2(n7770), .ZN(n14844) );
  OAI21_X1 U7373 ( .B1(n7599), .B2(n7352), .A(n7351), .ZN(n7798) );
  NAND2_X1 U7374 ( .A1(n7758), .A2(n6447), .ZN(n13141) );
  NAND2_X1 U7375 ( .A1(n7104), .A2(n7751), .ZN(n14837) );
  AND4_X1 U7376 ( .A1(n9070), .A2(n9069), .A3(n9068), .A4(n9067), .ZN(n10893)
         );
  AOI21_X1 U7377 ( .B1(n7063), .B2(n6879), .A(n6878), .ZN(n6877) );
  XNOR2_X2 U7378 ( .A(n10357), .B(n10689), .ZN(n10686) );
  NAND2_X1 U7379 ( .A1(n7766), .A2(n7596), .ZN(n7599) );
  AND2_X1 U7380 ( .A1(n6814), .A2(n6713), .ZN(n11862) );
  OAI22_X1 U7381 ( .A1(n9185), .A2(n8933), .B1(P2_DATAO_REG_11__SCAN_IN), .B2(
        n15289), .ZN(n9195) );
  AND2_X1 U7382 ( .A1(n9063), .A2(n6937), .ZN(n10732) );
  INV_X2 U7383 ( .A(n6827), .ZN(n9917) );
  AOI21_X1 U7384 ( .B1(n7065), .B2(n7068), .A(n7064), .ZN(n7063) );
  INV_X2 U7385 ( .A(n12315), .ZN(n12334) );
  AND2_X2 U7386 ( .A1(n12333), .A2(n14058), .ZN(n10923) );
  INV_X1 U7387 ( .A(n9037), .ZN(n10904) );
  AOI21_X1 U7388 ( .B1(n7069), .B2(n7067), .A(n7066), .ZN(n7065) );
  NAND4_X1 U7389 ( .A1(n9042), .A2(n9041), .A3(n9040), .A4(n9039), .ZN(n12560)
         );
  NAND2_X1 U7390 ( .A1(n8373), .A2(n6473), .ZN(n13811) );
  OAI21_X4 U7391 ( .B1(n10480), .B2(n10479), .A(n10478), .ZN(n10487) );
  AND3_X1 U7392 ( .A1(n9077), .A2(n9076), .A3(n9075), .ZN(n15069) );
  AND2_X1 U7393 ( .A1(n7070), .A2(n7549), .ZN(n7069) );
  AND2_X2 U7394 ( .A1(n10280), .A2(n10245), .ZN(n12315) );
  AND2_X1 U7395 ( .A1(n13629), .A2(n13634), .ZN(n7788) );
  NAND2_X1 U7396 ( .A1(n6761), .A2(n6760), .ZN(n14623) );
  CLKBUF_X3 U7397 ( .A(n7742), .Z(n9892) );
  XNOR2_X1 U7398 ( .A(n9173), .B(n9172), .ZN(n14963) );
  AOI21_X1 U7399 ( .B1(n7367), .B2(n7368), .A(n6534), .ZN(n7364) );
  AND2_X1 U7400 ( .A1(n7715), .A2(n7191), .ZN(n7426) );
  AND2_X1 U7401 ( .A1(n10242), .A2(n11378), .ZN(n10281) );
  XNOR2_X1 U7402 ( .A(n8318), .B(P1_IR_REG_19__SCAN_IN), .ZN(n10243) );
  XNOR2_X1 U7403 ( .A(n7712), .B(n13623), .ZN(n13629) );
  AOI21_X1 U7404 ( .B1(n7836), .B2(n7611), .A(n7855), .ZN(n7367) );
  XNOR2_X1 U7405 ( .A(n7695), .B(P2_IR_REG_22__SCAN_IN), .ZN(n12149) );
  OAI21_X1 U7406 ( .B1(n7708), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7707) );
  XNOR2_X1 U7407 ( .A(n7610), .B(SI_8_), .ZN(n7836) );
  XNOR2_X1 U7408 ( .A(n8876), .B(n8875), .ZN(n10224) );
  NAND2_X1 U7409 ( .A1(n7191), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7712) );
  NAND3_X1 U7410 ( .A1(n14186), .A2(n6815), .A3(n6515), .ZN(n14192) );
  NAND2_X1 U7411 ( .A1(n7102), .A2(n6456), .ZN(n6794) );
  NAND3_X1 U7412 ( .A1(n6793), .A2(n6792), .A3(n6507), .ZN(n13640) );
  OR2_X1 U7413 ( .A1(n15339), .A2(n6797), .ZN(n6793) );
  XNOR2_X1 U7414 ( .A(n7601), .B(n7079), .ZN(n7600) );
  OAI21_X1 U7415 ( .B1(n9058), .B2(n8922), .A(n8923), .ZN(n9072) );
  XNOR2_X1 U7416 ( .A(n7602), .B(SI_6_), .ZN(n7797) );
  XNOR2_X1 U7417 ( .A(n7597), .B(SI_4_), .ZN(n7767) );
  MUX2_X1 U7418 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8295), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n8296) );
  OAI21_X1 U7419 ( .B1(n7279), .B2(n6541), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n8877) );
  INV_X2 U7420 ( .A(n9834), .ZN(n9831) );
  OR2_X1 U7421 ( .A1(n7273), .A2(n7272), .ZN(n6815) );
  OR2_X1 U7422 ( .A1(n8322), .A2(n8589), .ZN(n8320) );
  NAND2_X2 U7423 ( .A1(n9031), .A2(P1_U3086), .ZN(n14204) );
  INV_X2 U7424 ( .A(n7595), .ZN(n9834) );
  OR2_X1 U7425 ( .A1(n7859), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n7991) );
  AND2_X1 U7426 ( .A1(n7318), .A2(n8293), .ZN(n7222) );
  AND2_X1 U7427 ( .A1(n7679), .A2(n6562), .ZN(n6695) );
  AND2_X1 U7428 ( .A1(n6750), .A2(n7679), .ZN(n7857) );
  AND2_X1 U7429 ( .A1(n7541), .A2(n7540), .ZN(n7539) );
  INV_X1 U7430 ( .A(n8287), .ZN(n7318) );
  NOR2_X1 U7431 ( .A1(n7118), .A2(n7116), .ZN(n8899) );
  AND3_X1 U7432 ( .A1(n7682), .A2(n7681), .A3(n7699), .ZN(n7685) );
  AND4_X1 U7433 ( .A1(n8283), .A2(n8412), .A3(n7034), .A4(n7035), .ZN(n7319)
         );
  AND3_X1 U7434 ( .A1(n7698), .A2(n7697), .A3(n7683), .ZN(n7684) );
  AND2_X1 U7435 ( .A1(n8360), .A2(n8282), .ZN(n7320) );
  AND2_X1 U7436 ( .A1(n8917), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9045) );
  NAND4_X1 U7437 ( .A1(n6861), .A2(n7780), .A3(n7818), .A4(n7783), .ZN(n7680)
         );
  AND4_X1 U7438 ( .A1(n8289), .A2(n8288), .A3(n8316), .A4(n8315), .ZN(n8290)
         );
  AND2_X1 U7439 ( .A1(n8894), .A2(n8893), .ZN(n8895) );
  NOR2_X1 U7440 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n7313) );
  CLKBUF_X2 U7441 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n14207) );
  INV_X1 U7442 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n9091) );
  INV_X4 U7443 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X4 U7444 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X2 U7445 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n10417) );
  INV_X1 U7446 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n9142) );
  INV_X1 U7447 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8412) );
  INV_X1 U7448 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n7875) );
  INV_X1 U7449 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7745) );
  NOR2_X1 U7450 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n6988) );
  NOR2_X1 U7451 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n8282) );
  INV_X1 U7452 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7780) );
  NOR2_X1 U7453 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n8894) );
  NOR2_X1 U7454 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8893) );
  INV_X1 U7455 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7783) );
  NOR2_X1 U7456 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n8289) );
  INV_X1 U7457 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7818) );
  INV_X1 U7458 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8898) );
  INV_X1 U7459 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9376) );
  NOR2_X1 U7460 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n7119) );
  NOR2_X1 U7461 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n7120) );
  INV_X1 U7462 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8954) );
  INV_X1 U7463 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8988) );
  OAI21_X2 U7464 ( .B1(n13846), .B2(P1_REG1_REG_14__SCAN_IN), .A(n13847), .ZN(
        n11495) );
  NOR2_X2 U7465 ( .A1(n10406), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n14867) );
  XNOR2_X1 U7467 ( .A(n6991), .B(n8955), .ZN(n9385) );
  AOI21_X2 U7468 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n10188), .A(n10180), .ZN(
        n10157) );
  INV_X4 U7469 ( .A(n9129), .ZN(n9286) );
  INV_X2 U7470 ( .A(n9834), .ZN(n6439) );
  AOI21_X2 U7471 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n13862), .A(n13861), .ZN(
        n13874) );
  OR2_X1 U7472 ( .A1(n8360), .A2(n8589), .ZN(n8361) );
  XNOR2_X2 U7473 ( .A(n8958), .B(n8957), .ZN(n9384) );
  AOI21_X1 U7474 ( .B1(n7565), .B2(n7377), .A(n7376), .ZN(n7375) );
  INV_X1 U7475 ( .A(n7637), .ZN(n7377) );
  INV_X1 U7476 ( .A(n7641), .ZN(n7376) );
  NOR2_X1 U7477 ( .A1(n12679), .A2(n7488), .ZN(n7487) );
  INV_X1 U7478 ( .A(n7490), .ZN(n7488) );
  INV_X1 U7479 ( .A(n13644), .ZN(n8215) );
  INV_X1 U7480 ( .A(n10281), .ZN(n10280) );
  NAND2_X1 U7481 ( .A1(n12804), .A2(n9589), .ZN(n12787) );
  NAND2_X1 U7482 ( .A1(n12809), .A2(n9257), .ZN(n12794) );
  NAND2_X1 U7483 ( .A1(n12944), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8903) );
  NAND2_X1 U7484 ( .A1(n7280), .A2(n7221), .ZN(n8298) );
  AND3_X1 U7485 ( .A1(n7318), .A2(n8293), .A3(n6755), .ZN(n7221) );
  NAND2_X1 U7486 ( .A1(n7039), .A2(n7036), .ZN(n8380) );
  OR2_X1 U7487 ( .A1(n8367), .A2(n8365), .ZN(n7039) );
  INV_X1 U7488 ( .A(n8828), .ZN(n7037) );
  AND2_X1 U7489 ( .A1(n6983), .A2(n10398), .ZN(n6982) );
  NAND2_X1 U7490 ( .A1(n6546), .A2(n9545), .ZN(n6983) );
  INV_X1 U7491 ( .A(n9567), .ZN(n6960) );
  NOR2_X1 U7492 ( .A1(n6471), .A2(n7046), .ZN(n7045) );
  NAND2_X1 U7493 ( .A1(n6537), .A2(n11721), .ZN(n7046) );
  AOI22_X1 U7494 ( .A1(n6972), .A2(n11748), .B1(n6973), .B2(n11748), .ZN(n6969) );
  NAND2_X1 U7495 ( .A1(n12024), .A2(n12025), .ZN(n7415) );
  INV_X1 U7496 ( .A(n6730), .ZN(n6728) );
  NAND2_X1 U7497 ( .A1(n12056), .A2(n12055), .ZN(n12080) );
  AND2_X1 U7498 ( .A1(n8737), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8750) );
  INV_X1 U7499 ( .A(n7628), .ZN(n6878) );
  NAND2_X1 U7500 ( .A1(n7347), .A2(n7346), .ZN(n7584) );
  AND2_X1 U7501 ( .A1(n7143), .A2(n6558), .ZN(n14217) );
  OR2_X1 U7502 ( .A1(n14257), .A2(P1_ADDR_REG_3__SCAN_IN), .ZN(n7143) );
  OAI21_X1 U7503 ( .B1(n9486), .B2(n12539), .A(n9498), .ZN(n9639) );
  AND2_X1 U7504 ( .A1(n12608), .A2(n12643), .ZN(n7017) );
  OR2_X1 U7505 ( .A1(n12423), .A2(n12196), .ZN(n9636) );
  OR2_X1 U7506 ( .A1(n12200), .A2(n12674), .ZN(n9632) );
  NAND2_X1 U7507 ( .A1(n12732), .A2(n7558), .ZN(n12716) );
  OR2_X1 U7508 ( .A1(n12907), .A2(n12747), .ZN(n7558) );
  OR2_X1 U7509 ( .A1(n12925), .A2(n12813), .ZN(n9589) );
  NAND2_X1 U7510 ( .A1(n10891), .A2(n7508), .ZN(n15047) );
  AND2_X1 U7511 ( .A1(n9110), .A2(n9097), .ZN(n7508) );
  INV_X1 U7512 ( .A(n15051), .ZN(n9110) );
  INV_X1 U7513 ( .A(n10714), .ZN(n10724) );
  OAI211_X1 U7514 ( .C1(n9339), .C2(n9836), .A(n9036), .B(n9035), .ZN(n9037)
         );
  NAND2_X1 U7515 ( .A1(n9048), .A2(n6494), .ZN(n9036) );
  INV_X1 U7516 ( .A(n7713), .ZN(n6831) );
  NAND2_X1 U7517 ( .A1(n15339), .A2(n7469), .ZN(n7102) );
  INV_X1 U7518 ( .A(n7973), .ZN(n7186) );
  NOR2_X1 U7519 ( .A1(n12124), .A2(n7188), .ZN(n7187) );
  INV_X1 U7520 ( .A(n7957), .ZN(n7188) );
  INV_X1 U7521 ( .A(n10776), .ZN(n7099) );
  INV_X1 U7522 ( .A(n13119), .ZN(n12042) );
  NAND2_X1 U7523 ( .A1(n7470), .A2(n15339), .ZN(n7713) );
  INV_X1 U7524 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7683) );
  INV_X1 U7525 ( .A(n11412), .ZN(n7522) );
  INV_X1 U7526 ( .A(n14192), .ZN(n8310) );
  INV_X1 U7527 ( .A(n12154), .ZN(n8305) );
  NAND2_X1 U7528 ( .A1(n7335), .A2(n6629), .ZN(n12401) );
  OR2_X1 U7529 ( .A1(n13936), .A2(n7339), .ZN(n6629) );
  AOI21_X1 U7530 ( .B1(n7338), .B2(n7337), .A(n7336), .ZN(n7335) );
  INV_X1 U7531 ( .A(n12379), .ZN(n7336) );
  OR2_X1 U7532 ( .A1(n10244), .A2(n10243), .ZN(n10245) );
  AND4_X1 U7533 ( .A1(n8872), .A2(n8292), .A3(n8291), .A4(n8862), .ZN(n8293)
         );
  AOI21_X1 U7534 ( .B1(n7078), .B2(n7374), .A(n6462), .ZN(n7077) );
  INV_X1 U7535 ( .A(n7644), .ZN(n7647) );
  INV_X1 U7536 ( .A(n7767), .ZN(n7596) );
  XNOR2_X1 U7537 ( .A(n14217), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n14220) );
  OAI22_X1 U7538 ( .A1(n14276), .A2(n14224), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n14274), .ZN(n14225) );
  AND2_X1 U7539 ( .A1(n14274), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n14224) );
  NAND2_X1 U7540 ( .A1(n7283), .A2(n12747), .ZN(n7282) );
  NAND2_X1 U7541 ( .A1(n9038), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n9053) );
  OAI21_X1 U7542 ( .B1(n11066), .B2(n7311), .A(n11065), .ZN(n7310) );
  AND2_X1 U7543 ( .A1(n9486), .A2(n12539), .ZN(n9642) );
  AOI21_X1 U7544 ( .B1(n7025), .B2(n10468), .A(n7024), .ZN(n7023) );
  AND2_X1 U7545 ( .A1(n10470), .A2(n14907), .ZN(n7024) );
  OR2_X1 U7546 ( .A1(n14898), .A2(n6567), .ZN(n6690) );
  NAND2_X1 U7547 ( .A1(n6690), .A2(n14922), .ZN(n6691) );
  OR2_X1 U7548 ( .A1(n14960), .A2(n14959), .ZN(n7174) );
  NAND2_X1 U7549 ( .A1(n6687), .A2(n6686), .ZN(n6871) );
  AOI21_X1 U7550 ( .B1(n12591), .B2(n7170), .A(n6609), .ZN(n6686) );
  NAND2_X1 U7551 ( .A1(n8987), .A2(n7314), .ZN(n9277) );
  AND2_X1 U7552 ( .A1(n7315), .A2(n8988), .ZN(n7314) );
  NAND2_X1 U7553 ( .A1(n7484), .A2(n7483), .ZN(n7482) );
  INV_X1 U7554 ( .A(n7572), .ZN(n7483) );
  NAND2_X1 U7555 ( .A1(n12695), .A2(n7491), .ZN(n7490) );
  INV_X1 U7556 ( .A(n12734), .ZN(n12702) );
  AND2_X1 U7557 ( .A1(n7507), .A2(n12773), .ZN(n7506) );
  NAND2_X1 U7558 ( .A1(n7504), .A2(n6516), .ZN(n7503) );
  NAND2_X1 U7559 ( .A1(n12792), .A2(n7507), .ZN(n12780) );
  AOI21_X1 U7560 ( .B1(n12817), .B2(n7123), .A(n7122), .ZN(n7121) );
  INV_X1 U7561 ( .A(n9586), .ZN(n7123) );
  INV_X1 U7562 ( .A(n9595), .ZN(n7122) );
  NOR2_X1 U7563 ( .A1(n12810), .A2(n6935), .ZN(n6934) );
  NAND2_X1 U7564 ( .A1(n12825), .A2(n9256), .ZN(n12809) );
  OAI21_X1 U7565 ( .B1(n11670), .B2(n6613), .A(n7496), .ZN(n6614) );
  NAND2_X1 U7566 ( .A1(n9238), .A2(n9506), .ZN(n6613) );
  NAND2_X1 U7567 ( .A1(n11671), .A2(n7499), .ZN(n11649) );
  AND2_X1 U7568 ( .A1(n9574), .A2(n9575), .ZN(n11673) );
  OR2_X1 U7569 ( .A1(n12941), .A2(n9809), .ZN(n10396) );
  AND2_X1 U7570 ( .A1(n10585), .A2(n12659), .ZN(n10905) );
  INV_X1 U7571 ( .A(n15136), .ZN(n15078) );
  NAND2_X1 U7572 ( .A1(n9460), .A2(n9496), .ZN(n15089) );
  NAND2_X1 U7573 ( .A1(n9973), .A2(n9438), .ZN(n9440) );
  AOI21_X1 U7574 ( .B1(n7269), .B2(n9354), .A(n6644), .ZN(n9470) );
  AND2_X1 U7575 ( .A1(n14194), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6644) );
  INV_X1 U7576 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7502) );
  OAI21_X1 U7577 ( .B1(n8972), .B2(n8970), .A(n6610), .ZN(n6833) );
  OAI21_X1 U7578 ( .B1(n8986), .B2(n8944), .A(n8945), .ZN(n9259) );
  INV_X1 U7579 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9226) );
  INV_X1 U7580 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U7581 ( .A1(n7435), .A2(n7434), .ZN(n7433) );
  NAND2_X1 U7582 ( .A1(n12986), .A2(n12992), .ZN(n7434) );
  NAND2_X1 U7583 ( .A1(n7437), .A2(n7436), .ZN(n7435) );
  INV_X1 U7584 ( .A(n12992), .ZN(n7436) );
  OR2_X1 U7585 ( .A1(n10141), .A2(n12103), .ZN(n9775) );
  NAND2_X1 U7586 ( .A1(n13088), .A2(n13090), .ZN(n13089) );
  AND2_X1 U7587 ( .A1(n8126), .A2(n8125), .ZN(n13093) );
  AND2_X1 U7588 ( .A1(n8018), .A2(n8017), .ZN(n13028) );
  NAND2_X1 U7589 ( .A1(n7717), .A2(n7426), .ZN(n7754) );
  NAND2_X1 U7590 ( .A1(n13305), .A2(n13286), .ZN(n13285) );
  AOI21_X1 U7591 ( .B1(n7218), .B2(n7216), .A(n6512), .ZN(n7215) );
  INV_X1 U7592 ( .A(n7218), .ZN(n7217) );
  INV_X1 U7593 ( .A(n8252), .ZN(n7216) );
  NAND2_X1 U7594 ( .A1(n6787), .A2(n8065), .ZN(n13364) );
  NAND2_X1 U7595 ( .A1(n8248), .A2(n12129), .ZN(n13384) );
  XNOR2_X1 U7596 ( .A(n13387), .B(n13124), .ZN(n13392) );
  NAND2_X1 U7597 ( .A1(n10848), .A2(n7834), .ZN(n7182) );
  XNOR2_X1 U7598 ( .A(n12089), .B(n12090), .ZN(n8261) );
  OR2_X1 U7599 ( .A1(n11860), .A2(n8178), .ZN(n9796) );
  INV_X1 U7600 ( .A(n13284), .ZN(n6800) );
  INV_X1 U7601 ( .A(n13117), .ZN(n9793) );
  AOI21_X1 U7602 ( .B1(n13265), .B2(n13267), .A(n13266), .ZN(n13269) );
  INV_X1 U7603 ( .A(n7724), .ZN(n12050) );
  AND2_X1 U7604 ( .A1(n8203), .A2(n8215), .ZN(n14827) );
  AND2_X1 U7605 ( .A1(n7550), .A2(n7471), .ZN(n7470) );
  NOR2_X1 U7606 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n7471) );
  INV_X1 U7607 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8191) );
  OR2_X2 U7608 ( .A1(n10221), .A2(n8881), .ZN(n10282) );
  NAND2_X1 U7609 ( .A1(n12278), .A2(n12279), .ZN(n13666) );
  AND2_X1 U7610 ( .A1(n10240), .A2(n10239), .ZN(n10673) );
  NAND2_X1 U7611 ( .A1(n10354), .A2(n10288), .ZN(n10356) );
  NAND2_X1 U7612 ( .A1(n14493), .A2(n14494), .ZN(n14506) );
  XNOR2_X1 U7613 ( .A(n10358), .B(n12334), .ZN(n10360) );
  AOI22_X1 U7614 ( .A1(n12319), .A2(n10357), .B1(n12333), .B2(n10689), .ZN(
        n10358) );
  INV_X1 U7615 ( .A(n10359), .ZN(n10362) );
  XNOR2_X1 U7616 ( .A(n8846), .B(n8883), .ZN(n7074) );
  CLKBUF_X2 U7617 ( .A(n8386), .Z(n8784) );
  AND2_X1 U7618 ( .A1(n12154), .A2(n8310), .ZN(n8386) );
  NOR2_X1 U7619 ( .A1(n13801), .A2(n14087), .ZN(n6832) );
  INV_X1 U7620 ( .A(n13922), .ZN(n6902) );
  NAND2_X1 U7621 ( .A1(n13973), .A2(n6504), .ZN(n13952) );
  NAND2_X1 U7622 ( .A1(n14002), .A2(n14008), .ZN(n7331) );
  NAND2_X1 U7623 ( .A1(n8343), .A2(n9031), .ZN(n8359) );
  NAND2_X1 U7624 ( .A1(n14047), .A2(n12347), .ZN(n12349) );
  NOR2_X1 U7625 ( .A1(n11719), .A2(n7262), .ZN(n7261) );
  NAND2_X1 U7626 ( .A1(n7275), .A2(n7274), .ZN(n10859) );
  AND2_X1 U7627 ( .A1(n10745), .A2(n10863), .ZN(n7274) );
  INV_X1 U7628 ( .A(n14740), .ZN(n14711) );
  OR2_X1 U7629 ( .A1(n14334), .A2(n7160), .ZN(n7158) );
  AOI21_X1 U7630 ( .B1(n14967), .B2(n14233), .A(n14232), .ZN(n14293) );
  NAND2_X1 U7631 ( .A1(n7152), .A2(n7154), .ZN(n7148) );
  NAND2_X1 U7632 ( .A1(n7149), .A2(n7151), .ZN(n7147) );
  AOI21_X1 U7633 ( .B1(n14606), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n14236), .ZN(
        n14249) );
  AND2_X1 U7634 ( .A1(n14251), .A2(n14252), .ZN(n14236) );
  NAND2_X1 U7635 ( .A1(n7564), .A2(n14299), .ZN(n7134) );
  NAND2_X1 U7636 ( .A1(n14421), .A2(n6852), .ZN(n12656) );
  OR2_X1 U7637 ( .A1(n14420), .A2(n12654), .ZN(n6852) );
  NAND2_X1 U7638 ( .A1(n10174), .A2(n10173), .ZN(n10172) );
  AND2_X1 U7639 ( .A1(n9819), .A2(n14197), .ZN(n14591) );
  XNOR2_X1 U7640 ( .A(n14253), .B(n6850), .ZN(n14334) );
  XNOR2_X1 U7641 ( .A(n14967), .B(P1_ADDR_REG_10__SCAN_IN), .ZN(n6850) );
  NAND2_X1 U7642 ( .A1(n14544), .A2(n14792), .ZN(n14543) );
  AND2_X1 U7643 ( .A1(n11871), .A2(n11870), .ZN(n11877) );
  NAND2_X1 U7644 ( .A1(n8399), .A2(n8398), .ZN(n8400) );
  OAI21_X1 U7645 ( .B1(n6747), .B2(n11903), .A(n6746), .ZN(n6745) );
  INV_X1 U7646 ( .A(n7411), .ZN(n6747) );
  NOR2_X1 U7647 ( .A1(n6841), .A2(n11906), .ZN(n6746) );
  INV_X1 U7648 ( .A(n7412), .ZN(n6841) );
  NAND2_X1 U7649 ( .A1(n9541), .A2(n6980), .ZN(n6978) );
  NOR2_X1 U7650 ( .A1(n10398), .A2(n6981), .ZN(n6980) );
  NAND2_X1 U7651 ( .A1(n9545), .A2(n9540), .ZN(n6981) );
  NAND2_X1 U7652 ( .A1(n6982), .A2(n9546), .ZN(n6979) );
  NOR2_X1 U7653 ( .A1(n11055), .A2(n6987), .ZN(n6986) );
  NOR2_X1 U7654 ( .A1(n9549), .A2(n10398), .ZN(n6987) );
  INV_X1 U7655 ( .A(n11956), .ZN(n6727) );
  NAND2_X1 U7656 ( .A1(n7423), .A2(n6511), .ZN(n11957) );
  NOR2_X1 U7657 ( .A1(n6517), .A2(n6724), .ZN(n6723) );
  AND2_X1 U7658 ( .A1(n11956), .A2(n6725), .ZN(n6724) );
  INV_X1 U7659 ( .A(n11958), .ZN(n6725) );
  AOI21_X1 U7660 ( .B1(n6958), .B2(n6960), .A(n9569), .ZN(n6957) );
  INV_X1 U7661 ( .A(n9570), .ZN(n6955) );
  AND2_X1 U7662 ( .A1(n6953), .A2(n6951), .ZN(n9578) );
  AOI21_X1 U7663 ( .B1(n6969), .B2(n6457), .A(n6529), .ZN(n6967) );
  INV_X1 U7664 ( .A(n6969), .ZN(n6968) );
  INV_X1 U7665 ( .A(n9587), .ZN(n6966) );
  INV_X1 U7666 ( .A(n12032), .ZN(n7397) );
  NAND2_X1 U7667 ( .A1(n6739), .A2(n6740), .ZN(n7400) );
  AOI21_X1 U7668 ( .B1(n6548), .B2(n12027), .A(n6463), .ZN(n6740) );
  NAND2_X1 U7669 ( .A1(n12031), .A2(n12032), .ZN(n7399) );
  NAND2_X1 U7670 ( .A1(n12034), .A2(n12033), .ZN(n6733) );
  NAND2_X1 U7671 ( .A1(n8687), .A2(n7062), .ZN(n7061) );
  NOR2_X1 U7672 ( .A1(n6446), .A2(n12035), .ZN(n7401) );
  NOR2_X1 U7673 ( .A1(n6446), .A2(n7403), .ZN(n7402) );
  NAND2_X1 U7674 ( .A1(n6730), .A2(n6729), .ZN(n12038) );
  INV_X1 U7675 ( .A(n12037), .ZN(n7403) );
  AOI22_X1 U7676 ( .A1(n12058), .A2(n11863), .B1(n12085), .B2(n12057), .ZN(
        n12075) );
  INV_X1 U7677 ( .A(n8734), .ZN(n7053) );
  NAND2_X1 U7678 ( .A1(n8719), .A2(n8721), .ZN(n7384) );
  NAND2_X1 U7679 ( .A1(n7051), .A2(n8734), .ZN(n7050) );
  INV_X1 U7680 ( .A(n7663), .ZN(n7083) );
  INV_X1 U7681 ( .A(n9531), .ZN(n7115) );
  INV_X1 U7682 ( .A(n7129), .ZN(n7127) );
  NAND2_X1 U7683 ( .A1(n12377), .A2(n12378), .ZN(n7340) );
  INV_X1 U7684 ( .A(n14037), .ZN(n7223) );
  AND2_X1 U7685 ( .A1(n7652), .A2(n7089), .ZN(n7088) );
  INV_X1 U7686 ( .A(n8022), .ZN(n7089) );
  OAI21_X1 U7687 ( .B1(n7375), .B2(SI_17_), .A(SI_18_), .ZN(n6895) );
  NOR2_X1 U7688 ( .A1(n6889), .A2(n6525), .ZN(n6888) );
  INV_X1 U7689 ( .A(n7632), .ZN(n6889) );
  NOR2_X1 U7690 ( .A1(n7987), .A2(n6898), .ZN(n6893) );
  OR2_X1 U7691 ( .A1(n6441), .A2(n7646), .ZN(n6892) );
  NAND2_X1 U7692 ( .A1(n7638), .A2(n10139), .ZN(n7641) );
  INV_X1 U7693 ( .A(n12459), .ZN(n7297) );
  INV_X1 U7694 ( .A(n9642), .ZN(n9513) );
  OR2_X1 U7695 ( .A1(n6452), .A2(n12627), .ZN(n7001) );
  NOR2_X1 U7696 ( .A1(n14396), .A2(n12627), .ZN(n7000) );
  INV_X1 U7697 ( .A(n9368), .ZN(n11854) );
  AND2_X1 U7698 ( .A1(n12688), .A2(n9625), .ZN(n7129) );
  NAND2_X1 U7699 ( .A1(n7493), .A2(n12703), .ZN(n7492) );
  OR2_X1 U7700 ( .A1(n12774), .A2(n12782), .ZN(n9604) );
  AND2_X1 U7701 ( .A1(n12786), .A2(n9274), .ZN(n7507) );
  NOR2_X1 U7702 ( .A1(n9403), .A2(n6929), .ZN(n6928) );
  INV_X1 U7703 ( .A(n9572), .ZN(n6929) );
  AND2_X1 U7704 ( .A1(n11650), .A2(n9222), .ZN(n7499) );
  AND2_X1 U7705 ( .A1(n9402), .A2(n7476), .ZN(n7475) );
  NAND2_X1 U7706 ( .A1(n9192), .A2(n7477), .ZN(n7476) );
  INV_X1 U7707 ( .A(n9191), .ZN(n7477) );
  INV_X1 U7708 ( .A(n9192), .ZN(n7478) );
  INV_X1 U7709 ( .A(n10962), .ZN(n9457) );
  NOR2_X1 U7710 ( .A1(n7246), .A2(n7243), .ZN(n7242) );
  INV_X1 U7711 ( .A(n8940), .ZN(n7245) );
  INV_X1 U7712 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8939) );
  NAND2_X1 U7713 ( .A1(n6642), .A2(n8934), .ZN(n8936) );
  NAND2_X1 U7714 ( .A1(n9195), .A2(n9193), .ZN(n6642) );
  NAND2_X1 U7715 ( .A1(n13046), .A2(n6705), .ZN(n6703) );
  INV_X1 U7716 ( .A(n12977), .ZN(n6705) );
  AND2_X1 U7717 ( .A1(n9709), .A2(n9703), .ZN(n7467) );
  NOR2_X1 U7718 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n6830) );
  INV_X1 U7719 ( .A(n12067), .ZN(n7394) );
  NAND2_X1 U7720 ( .A1(n7391), .A2(n7388), .ZN(n7392) );
  INV_X1 U7721 ( .A(n13629), .ZN(n7717) );
  AND2_X1 U7722 ( .A1(n8178), .A2(n12149), .ZN(n9890) );
  NOR2_X1 U7723 ( .A1(n6466), .A2(n8101), .ZN(n6784) );
  INV_X1 U7724 ( .A(n9892), .ZN(n6715) );
  OAI21_X1 U7725 ( .B1(n13283), .B2(n7179), .A(n7175), .ZN(n7177) );
  AOI21_X1 U7726 ( .B1(n7178), .B2(n13280), .A(n7176), .ZN(n7175) );
  INV_X1 U7727 ( .A(n8170), .ZN(n7176) );
  NOR2_X1 U7728 ( .A1(n13489), .A2(n13569), .ZN(n7100) );
  NAND2_X1 U7729 ( .A1(n11684), .A2(n11968), .ZN(n11773) );
  NAND2_X1 U7730 ( .A1(n10987), .A2(n7854), .ZN(n11237) );
  NAND2_X1 U7731 ( .A1(n11237), .A2(n11236), .ZN(n11235) );
  NOR2_X1 U7732 ( .A1(n13143), .A2(n11865), .ZN(n10198) );
  INV_X1 U7733 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8188) );
  INV_X1 U7734 ( .A(n11188), .ZN(n7528) );
  AND2_X1 U7735 ( .A1(n12277), .A2(n12276), .ZN(n12279) );
  OR2_X1 U7736 ( .A1(n8779), .A2(n10012), .ZN(n8356) );
  NAND2_X1 U7737 ( .A1(n13974), .A2(n6628), .ZN(n13955) );
  AND2_X1 U7738 ( .A1(n13956), .A2(n12375), .ZN(n6628) );
  NAND2_X1 U7739 ( .A1(n7223), .A2(n6909), .ZN(n6911) );
  NOR2_X1 U7740 ( .A1(n14012), .A2(n14130), .ZN(n6909) );
  XNOR2_X1 U7741 ( .A(n14119), .B(n6899), .ZN(n12372) );
  NAND2_X1 U7742 ( .A1(n7330), .A2(n12362), .ZN(n7329) );
  NOR2_X1 U7743 ( .A1(n14349), .A2(n6464), .ZN(n7324) );
  INV_X1 U7744 ( .A(n11625), .ZN(n6625) );
  INV_X1 U7745 ( .A(n11585), .ZN(n7321) );
  NAND2_X1 U7746 ( .A1(n11584), .A2(n11583), .ZN(n11586) );
  NAND2_X1 U7747 ( .A1(n10973), .A2(n10972), .ZN(n7343) );
  INV_X1 U7748 ( .A(n10755), .ZN(n7326) );
  NAND2_X1 U7749 ( .A1(n8829), .A2(n10749), .ZN(n10738) );
  NAND2_X1 U7750 ( .A1(n13936), .A2(n12378), .ZN(n7334) );
  AOI21_X1 U7751 ( .B1(n6442), .B2(n8102), .A(n6604), .ZN(n7081) );
  INV_X1 U7752 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7543) );
  INV_X1 U7753 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8319) );
  NAND2_X1 U7754 ( .A1(n7634), .A2(n10040), .ZN(n7637) );
  INV_X1 U7755 ( .A(n7624), .ZN(n7066) );
  INV_X1 U7756 ( .A(n7620), .ZN(n7067) );
  INV_X1 U7757 ( .A(n7598), .ZN(n7354) );
  NAND2_X1 U7758 ( .A1(n7594), .A2(n7593), .ZN(n7766) );
  INV_X1 U7759 ( .A(P1_RD_REG_SCAN_IN), .ZN(n6777) );
  INV_X1 U7760 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7576) );
  INV_X1 U7761 ( .A(n7595), .ZN(n9031) );
  AOI21_X1 U7762 ( .B1(n14220), .B2(n14219), .A(n14218), .ZN(n14221) );
  INV_X1 U7763 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14219) );
  XNOR2_X1 U7764 ( .A(n14221), .B(n6849), .ZN(n14256) );
  AOI21_X1 U7765 ( .B1(n14254), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n14226), .ZN(
        n14282) );
  AOI21_X1 U7766 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n14235), .A(n14234), .ZN(
        n14251) );
  NOR2_X1 U7767 ( .A1(n14293), .A2(n14294), .ZN(n14234) );
  OR2_X1 U7768 ( .A1(n14247), .A2(n14246), .ZN(n14238) );
  AND3_X1 U7769 ( .A1(n9127), .A2(n9126), .A3(n9125), .ZN(n11100) );
  NAND2_X1 U7770 ( .A1(n12501), .A2(n6505), .ZN(n7283) );
  INV_X1 U7771 ( .A(n12177), .ZN(n7284) );
  AND2_X1 U7772 ( .A1(n12513), .A2(n6676), .ZN(n6675) );
  NAND2_X1 U7773 ( .A1(n6677), .A2(n12162), .ZN(n6676) );
  INV_X1 U7774 ( .A(n12161), .ZN(n6677) );
  AOI21_X1 U7775 ( .B1(n12434), .B2(n12189), .A(n12193), .ZN(n7291) );
  OAI21_X1 U7776 ( .B1(n11388), .B2(n11343), .A(n7303), .ZN(n7302) );
  NAND2_X1 U7777 ( .A1(n7304), .A2(n14436), .ZN(n7303) );
  NAND2_X1 U7778 ( .A1(n12178), .A2(n12177), .ZN(n12484) );
  NAND2_X1 U7779 ( .A1(n6682), .A2(n6681), .ZN(n7305) );
  INV_X1 U7780 ( .A(n10592), .ZN(n6681) );
  INV_X1 U7781 ( .A(n10593), .ZN(n6682) );
  AND2_X1 U7782 ( .A1(n9130), .A2(n10556), .ZN(n9151) );
  NOR2_X1 U7783 ( .A1(n7310), .A2(n11068), .ZN(n7306) );
  NAND2_X1 U7784 ( .A1(n6444), .A2(n6670), .ZN(n6668) );
  INV_X1 U7785 ( .A(n7545), .ZN(n6670) );
  NAND2_X1 U7786 ( .A1(n7305), .A2(n7308), .ZN(n7307) );
  NOR2_X1 U7787 ( .A1(n11066), .A2(n10806), .ZN(n7308) );
  XNOR2_X1 U7788 ( .A(n11571), .B(n10487), .ZN(n7304) );
  NAND2_X1 U7789 ( .A1(n12469), .A2(n12187), .ZN(n12526) );
  OR2_X1 U7790 ( .A1(n10422), .A2(n14865), .ZN(n7167) );
  NAND2_X1 U7791 ( .A1(n12569), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n6853) );
  OR2_X1 U7792 ( .A1(n14884), .A2(n10468), .ZN(n7026) );
  OR2_X1 U7793 ( .A1(n14916), .A2(n10448), .ZN(n7169) );
  NOR2_X1 U7794 ( .A1(n9106), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n9123) );
  INV_X1 U7795 ( .A(n6847), .ZN(n12582) );
  INV_X1 U7796 ( .A(n14979), .ZN(n7015) );
  NAND2_X1 U7797 ( .A1(n7174), .A2(n7173), .ZN(n7172) );
  NAND2_X1 U7798 ( .A1(n14963), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7173) );
  OR2_X1 U7799 ( .A1(n14987), .A2(n14986), .ZN(n7163) );
  NAND2_X1 U7800 ( .A1(n7015), .A2(n7012), .ZN(n7010) );
  INV_X1 U7801 ( .A(n7017), .ZN(n7012) );
  INV_X1 U7802 ( .A(n12607), .ZN(n7014) );
  INV_X1 U7803 ( .A(n7010), .ZN(n7009) );
  NAND2_X1 U7804 ( .A1(n7163), .A2(n7162), .ZN(n7161) );
  NAND2_X1 U7805 ( .A1(n14323), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7162) );
  NOR2_X1 U7806 ( .A1(n15016), .A2(n15017), .ZN(n15015) );
  AND2_X1 U7807 ( .A1(n12622), .A2(n12621), .ZN(n7005) );
  AOI21_X1 U7808 ( .B1(n7005), .B2(n7004), .A(n6605), .ZN(n7003) );
  NAND2_X1 U7809 ( .A1(n14379), .A2(n7004), .ZN(n7002) );
  INV_X1 U7810 ( .A(n6871), .ZN(n12593) );
  NAND2_X1 U7811 ( .A1(n14422), .A2(n14423), .ZN(n14421) );
  AND2_X1 U7812 ( .A1(n9651), .A2(n9351), .ZN(n12679) );
  NAND2_X1 U7813 ( .A1(n12687), .A2(n7492), .ZN(n7489) );
  NAND2_X1 U7814 ( .A1(n12721), .A2(n7551), .ZN(n12699) );
  AOI21_X1 U7815 ( .B1(n12745), .B2(n9314), .A(n6540), .ZN(n12733) );
  NAND2_X1 U7816 ( .A1(n7109), .A2(n9611), .ZN(n12738) );
  OR2_X1 U7817 ( .A1(n9296), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9298) );
  NAND2_X1 U7818 ( .A1(n12770), .A2(n9604), .ZN(n12761) );
  NAND2_X1 U7819 ( .A1(n12455), .A2(n9290), .ZN(n9291) );
  INV_X1 U7820 ( .A(n12794), .ZN(n9273) );
  NOR2_X1 U7821 ( .A1(n9272), .A2(n6932), .ZN(n6931) );
  INV_X1 U7822 ( .A(n7121), .ZN(n6932) );
  NAND2_X1 U7823 ( .A1(n9255), .A2(n6935), .ZN(n12825) );
  AOI21_X1 U7824 ( .B1(n6928), .B2(n9402), .A(n6926), .ZN(n6925) );
  INV_X1 U7825 ( .A(n9575), .ZN(n6926) );
  INV_X1 U7826 ( .A(n6928), .ZN(n6927) );
  INV_X1 U7827 ( .A(n11670), .ZN(n6612) );
  AND4_X1 U7828 ( .A1(n9207), .A2(n9206), .A3(n9205), .A4(n9204), .ZN(n11675)
         );
  NAND2_X1 U7829 ( .A1(n6615), .A2(n7494), .ZN(n11223) );
  AOI21_X1 U7830 ( .B1(n7495), .B2(n11046), .A(n6484), .ZN(n7494) );
  NAND2_X1 U7831 ( .A1(n11044), .A2(n7495), .ZN(n6615) );
  NAND2_X1 U7832 ( .A1(n11045), .A2(n11046), .ZN(n7130) );
  NAND2_X1 U7833 ( .A1(n15047), .A2(n9112), .ZN(n10878) );
  AND2_X1 U7834 ( .A1(n9549), .A2(n9545), .ZN(n15051) );
  INV_X1 U7835 ( .A(n15089), .ZN(n15049) );
  INV_X1 U7836 ( .A(n10890), .ZN(n9096) );
  AND4_X1 U7837 ( .A1(n9087), .A2(n9086), .A3(n9085), .A4(n9084), .ZN(n15061)
         );
  NAND2_X1 U7838 ( .A1(n10398), .A2(n9386), .ZN(n15084) );
  AND2_X1 U7839 ( .A1(n10398), .A2(n9391), .ZN(n14437) );
  NAND2_X1 U7840 ( .A1(n9367), .A2(n9366), .ZN(n12423) );
  OAI21_X1 U7841 ( .B1(n12949), .B2(n9472), .A(n7267), .ZN(n14452) );
  OR2_X1 U7842 ( .A1(n6440), .A2(n12948), .ZN(n7267) );
  INV_X1 U7843 ( .A(n10732), .ZN(n15108) );
  NOR2_X1 U7844 ( .A1(n10388), .A2(n9633), .ZN(n10376) );
  INV_X1 U7845 ( .A(n14437), .ZN(n15087) );
  AOI21_X1 U7846 ( .B1(n9470), .B2(n9469), .A(n6611), .ZN(n9481) );
  NAND2_X1 U7847 ( .A1(n15193), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7270) );
  AOI21_X1 U7848 ( .B1(n6833), .B2(n8953), .A(n7271), .ZN(n9353) );
  AND2_X1 U7849 ( .A1(n14200), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7271) );
  INV_X1 U7850 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7500) );
  AND2_X1 U7851 ( .A1(n6556), .A2(n6633), .ZN(n8972) );
  NAND2_X1 U7852 ( .A1(n9326), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6633) );
  XNOR2_X1 U7853 ( .A(n8951), .B(n14202), .ZN(n9326) );
  NAND2_X1 U7854 ( .A1(n9303), .A2(n9302), .ZN(n8947) );
  INV_X1 U7855 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9414) );
  OAI21_X1 U7856 ( .B1(n9413), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9415) );
  AND2_X1 U7857 ( .A1(n6636), .A2(n7248), .ZN(n9303) );
  NAND2_X1 U7858 ( .A1(n15178), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7248) );
  NAND2_X1 U7859 ( .A1(n7251), .A2(n6634), .ZN(n6636) );
  NOR2_X1 U7860 ( .A1(n8975), .A2(n6635), .ZN(n6634) );
  NOR2_X1 U7861 ( .A1(n6947), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n6946) );
  NAND2_X1 U7862 ( .A1(n9377), .A2(n9376), .ZN(n9413) );
  INV_X1 U7863 ( .A(n9379), .ZN(n9377) );
  NAND2_X1 U7864 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n7250), .ZN(n7249) );
  NAND2_X1 U7865 ( .A1(n8898), .A2(n7117), .ZN(n6947) );
  NAND2_X1 U7866 ( .A1(n8943), .A2(n8942), .ZN(n8986) );
  OAI21_X1 U7867 ( .B1(n9170), .B2(n8932), .A(n8931), .ZN(n9185) );
  OAI21_X1 U7868 ( .B1(n9186), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9187) );
  AND2_X1 U7869 ( .A1(n15276), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8930) );
  AND2_X1 U7870 ( .A1(n9139), .A2(n9138), .ZN(n9143) );
  INV_X1 U7871 ( .A(n8929), .ZN(n7235) );
  INV_X1 U7872 ( .A(n7234), .ZN(n7233) );
  OAI21_X1 U7873 ( .B1(n7237), .B2(n6443), .A(n7239), .ZN(n7234) );
  NAND2_X1 U7874 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n7240), .ZN(n7239) );
  NOR2_X1 U7875 ( .A1(n9104), .A2(n7238), .ZN(n7237) );
  INV_X1 U7876 ( .A(n8926), .ZN(n7238) );
  NAND2_X1 U7877 ( .A1(n9089), .A2(n9088), .ZN(n8927) );
  XNOR2_X1 U7878 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n9088) );
  NAND2_X1 U7879 ( .A1(n6643), .A2(n8921), .ZN(n9058) );
  NAND2_X1 U7880 ( .A1(n9021), .A2(n8920), .ZN(n6643) );
  INV_X1 U7881 ( .A(n13140), .ZN(n7777) );
  INV_X1 U7882 ( .A(n13121), .ZN(n13040) );
  INV_X1 U7883 ( .A(n6700), .ZN(n6699) );
  OAI21_X1 U7884 ( .B1(n7467), .B2(n6701), .A(n11202), .ZN(n6700) );
  INV_X1 U7885 ( .A(n9710), .ZN(n6701) );
  NAND2_X1 U7886 ( .A1(n7468), .A2(n7467), .ZN(n11127) );
  NAND2_X1 U7887 ( .A1(n8042), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8058) );
  NOR2_X1 U7888 ( .A1(n6510), .A2(n7444), .ZN(n7443) );
  NOR2_X1 U7889 ( .A1(n12976), .A2(n7445), .ZN(n7444) );
  AND2_X1 U7890 ( .A1(n7555), .A2(n7441), .ZN(n7440) );
  NOR2_X1 U7891 ( .A1(n7446), .A2(n13016), .ZN(n7441) );
  NAND2_X1 U7892 ( .A1(n7447), .A2(n13023), .ZN(n7446) );
  NAND2_X1 U7893 ( .A1(n9725), .A2(n9724), .ZN(n11572) );
  INV_X1 U7894 ( .A(n11574), .ZN(n9725) );
  AND4_X1 U7895 ( .A1(n7955), .A2(n7954), .A3(n7953), .A4(n7952), .ZN(n11967)
         );
  BUF_X1 U7896 ( .A(n8079), .Z(n6827) );
  OR2_X1 U7897 ( .A1(n8079), .A2(n7737), .ZN(n7741) );
  INV_X1 U7898 ( .A(n7788), .ZN(n7965) );
  NAND2_X1 U7899 ( .A1(n13634), .A2(n7717), .ZN(n8079) );
  NAND2_X1 U7900 ( .A1(n13283), .A2(n13282), .ZN(n13265) );
  NAND2_X1 U7901 ( .A1(n6782), .A2(n6783), .ZN(n6781) );
  NAND2_X1 U7902 ( .A1(n6788), .A2(n13392), .ZN(n6803) );
  INV_X1 U7903 ( .A(n8038), .ZN(n6788) );
  AOI21_X1 U7904 ( .B1(n13392), .B2(n6805), .A(n6521), .ZN(n6804) );
  INV_X1 U7905 ( .A(n8037), .ZN(n6805) );
  AND2_X1 U7906 ( .A1(n6499), .A2(n8000), .ZN(n7193) );
  NOR2_X1 U7907 ( .A1(n13424), .A2(n7214), .ZN(n7213) );
  INV_X1 U7908 ( .A(n8247), .ZN(n7214) );
  NAND2_X1 U7909 ( .A1(n7742), .A2(n9831), .ZN(n8088) );
  NAND2_X1 U7910 ( .A1(n6807), .A2(n6806), .ZN(n13432) );
  NAND2_X1 U7911 ( .A1(n7185), .A2(n7986), .ZN(n6806) );
  NAND2_X1 U7912 ( .A1(n13432), .A2(n13431), .ZN(n13429) );
  NAND2_X1 U7913 ( .A1(n7958), .A2(n7187), .ZN(n11767) );
  NAND2_X1 U7914 ( .A1(n11284), .A2(n7192), .ZN(n11458) );
  AND2_X1 U7915 ( .A1(n12120), .A2(n7890), .ZN(n7192) );
  NAND2_X1 U7916 ( .A1(n7182), .A2(n7180), .ZN(n10987) );
  NOR2_X1 U7917 ( .A1(n12115), .A2(n7181), .ZN(n7180) );
  INV_X1 U7918 ( .A(n7835), .ZN(n7181) );
  NAND2_X1 U7919 ( .A1(n11029), .A2(n7814), .ZN(n10848) );
  NAND2_X1 U7920 ( .A1(n7098), .A2(n10852), .ZN(n7095) );
  NOR2_X1 U7921 ( .A1(n10776), .A2(n14844), .ZN(n10775) );
  AND2_X1 U7922 ( .A1(n8222), .A2(n8178), .ZN(n12090) );
  XNOR2_X1 U7923 ( .A(n10778), .B(n7777), .ZN(n10769) );
  NAND2_X1 U7924 ( .A1(n10652), .A2(n7752), .ZN(n10347) );
  XNOR2_X1 U7925 ( .A(n13142), .B(n14837), .ZN(n12105) );
  NAND2_X1 U7926 ( .A1(n10653), .A2(n12105), .ZN(n10652) );
  INV_X1 U7927 ( .A(n10140), .ZN(n10196) );
  INV_X1 U7928 ( .A(n7202), .ZN(n7201) );
  NOR2_X1 U7929 ( .A1(n8256), .A2(n7206), .ZN(n7205) );
  INV_X1 U7930 ( .A(n8254), .ZN(n7206) );
  NAND2_X1 U7931 ( .A1(n8251), .A2(n12102), .ZN(n13354) );
  OR2_X1 U7932 ( .A1(n13370), .A2(n8250), .ZN(n8251) );
  OR2_X1 U7933 ( .A1(n13354), .A2(n13365), .ZN(n13355) );
  NAND2_X1 U7934 ( .A1(n13437), .A2(n13436), .ZN(n13435) );
  NOR2_X1 U7935 ( .A1(n7208), .A2(n6500), .ZN(n7207) );
  NOR2_X1 U7936 ( .A1(n6476), .A2(n12117), .ZN(n7208) );
  XNOR2_X1 U7937 ( .A(n8217), .B(n8216), .ZN(n11742) );
  MUX2_X1 U7938 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7714), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n7715) );
  INV_X1 U7939 ( .A(n7691), .ZN(n6751) );
  OR2_X1 U7940 ( .A1(n8196), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n8200) );
  NAND2_X1 U7941 ( .A1(n8189), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8217) );
  INV_X1 U7942 ( .A(n8194), .ZN(n8189) );
  INV_X1 U7943 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8216) );
  INV_X1 U7944 ( .A(n10920), .ZN(n6650) );
  NOR2_X1 U7945 ( .A1(n14567), .A2(n6648), .ZN(n6647) );
  INV_X1 U7946 ( .A(n6816), .ZN(n6648) );
  NOR2_X1 U7947 ( .A1(n11402), .A2(n11401), .ZN(n7525) );
  INV_X1 U7948 ( .A(n11403), .ZN(n7526) );
  AND2_X1 U7949 ( .A1(n8566), .A2(n8307), .ZN(n8582) );
  AND2_X1 U7950 ( .A1(n13694), .A2(n12301), .ZN(n13728) );
  OR2_X1 U7951 ( .A1(n8467), .A2(n8466), .ZN(n8484) );
  AND2_X1 U7952 ( .A1(n10284), .A2(n10283), .ZN(n10288) );
  NAND2_X1 U7953 ( .A1(n10287), .A2(n10286), .ZN(n10354) );
  INV_X1 U7954 ( .A(n11838), .ZN(n7530) );
  AND2_X1 U7955 ( .A1(n11845), .A2(n7534), .ZN(n7533) );
  INV_X1 U7956 ( .A(n7554), .ZN(n7534) );
  OAI21_X1 U7957 ( .B1(n13737), .B2(n7536), .A(n6659), .ZN(n6662) );
  AOI21_X1 U7958 ( .B1(n7535), .B2(n6661), .A(n6660), .ZN(n6659) );
  INV_X1 U7959 ( .A(n13738), .ZN(n6661) );
  AOI21_X1 U7960 ( .B1(n12219), .B2(n6654), .A(n6495), .ZN(n6653) );
  INV_X1 U7961 ( .A(n12219), .ZN(n6655) );
  INV_X2 U7962 ( .A(n10923), .ZN(n12317) );
  AND4_X1 U7963 ( .A1(n8559), .A2(n8558), .A3(n8557), .A4(n8556), .ZN(n13753)
         );
  NAND2_X1 U7964 ( .A1(n6885), .A2(n6882), .ZN(n6621) );
  NAND2_X1 U7965 ( .A1(n14082), .A2(n13660), .ZN(n6881) );
  NAND2_X1 U7966 ( .A1(n6883), .A2(n13800), .ZN(n6882) );
  INV_X1 U7967 ( .A(n7257), .ZN(n7256) );
  NAND2_X1 U7968 ( .A1(n13920), .A2(n12377), .ZN(n7258) );
  OAI21_X1 U7969 ( .B1(n13928), .B2(n7259), .A(n6502), .ZN(n7257) );
  AND2_X1 U7970 ( .A1(n8752), .A2(n8740), .ZN(n13662) );
  NAND2_X1 U7971 ( .A1(n13993), .A2(n14112), .ZN(n13978) );
  NAND2_X1 U7972 ( .A1(n14006), .A2(n12354), .ZN(n13990) );
  INV_X1 U7973 ( .A(n12372), .ZN(n13989) );
  NAND2_X1 U7974 ( .A1(n14023), .A2(n12369), .ZN(n14002) );
  AOI21_X1 U7975 ( .B1(n11723), .B2(n6765), .A(n6522), .ZN(n6763) );
  INV_X1 U7976 ( .A(n6765), .ZN(n6764) );
  NAND2_X1 U7977 ( .A1(n11731), .A2(n11730), .ZN(n11807) );
  AND4_X1 U7978 ( .A1(n8573), .A2(n8572), .A3(n8571), .A4(n8570), .ZN(n12226)
         );
  NAND2_X1 U7979 ( .A1(n8544), .A2(n8543), .ZN(n14343) );
  NAND2_X1 U7980 ( .A1(n11586), .A2(n11585), .ZN(n14350) );
  AND4_X1 U7981 ( .A1(n8510), .A2(n8509), .A3(n8508), .A4(n8507), .ZN(n11833)
         );
  AND4_X1 U7982 ( .A1(n8526), .A2(n8525), .A3(n8524), .A4(n8523), .ZN(n11843)
         );
  AND2_X1 U7983 ( .A1(n11477), .A2(n7254), .ZN(n7253) );
  OR2_X1 U7984 ( .A1(n11153), .A2(n7255), .ZN(n7254) );
  INV_X1 U7985 ( .A(n11329), .ZN(n7255) );
  NAND2_X1 U7986 ( .A1(n11246), .A2(n11146), .ZN(n11147) );
  NAND2_X1 U7987 ( .A1(n11249), .A2(n11152), .ZN(n11154) );
  NAND2_X1 U7988 ( .A1(n11154), .A2(n11153), .ZN(n11330) );
  NAND2_X1 U7989 ( .A1(n11248), .A2(n11247), .ZN(n11246) );
  NAND2_X1 U7990 ( .A1(n11074), .A2(n10978), .ZN(n10980) );
  NAND2_X1 U7991 ( .A1(n10971), .A2(n10970), .ZN(n11080) );
  NAND2_X1 U7992 ( .A1(n10968), .A2(n10967), .ZN(n10971) );
  AND2_X1 U7993 ( .A1(n10870), .A2(n10757), .ZN(n11077) );
  NAND2_X1 U7994 ( .A1(n10823), .A2(n10752), .ZN(n10955) );
  AND4_X1 U7995 ( .A1(n8407), .A2(n8406), .A3(n8405), .A4(n8404), .ZN(n11017)
         );
  INV_X1 U7996 ( .A(n14630), .ZN(n6757) );
  NAND2_X1 U7997 ( .A1(n13813), .A2(n14623), .ZN(n14630) );
  NOR2_X1 U7998 ( .A1(n14058), .A2(n8883), .ZN(n10930) );
  NAND2_X1 U7999 ( .A1(n13910), .A2(n13911), .ZN(n6915) );
  INV_X1 U8000 ( .A(n7230), .ZN(n13910) );
  AOI21_X1 U8001 ( .B1(n14082), .B2(n14740), .A(n14081), .ZN(n6914) );
  INV_X1 U8002 ( .A(n14138), .ZN(n14621) );
  AND2_X1 U8003 ( .A1(n10225), .A2(n10224), .ZN(n10322) );
  INV_X1 U8004 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7345) );
  AND2_X1 U8005 ( .A1(n7319), .A2(n7277), .ZN(n7276) );
  AND2_X1 U8006 ( .A1(n7320), .A2(n8290), .ZN(n7278) );
  NOR2_X1 U8007 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n7277) );
  XNOR2_X1 U8008 ( .A(n8863), .B(n8862), .ZN(n10933) );
  NAND2_X1 U8009 ( .A1(n8325), .A2(n7539), .ZN(n8868) );
  NOR2_X1 U8010 ( .A1(n7279), .A2(n7542), .ZN(n8322) );
  AOI21_X1 U8011 ( .B1(n7959), .B2(n7078), .A(n7076), .ZN(n7075) );
  INV_X1 U8012 ( .A(n7077), .ZN(n7076) );
  INV_X1 U8013 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n14262) );
  NAND2_X1 U8014 ( .A1(n15318), .A2(n14269), .ZN(n14272) );
  AND2_X1 U8015 ( .A1(n7139), .A2(n6490), .ZN(n14286) );
  OAI21_X1 U8016 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n14230), .A(n14229), .ZN(
        n14253) );
  AOI21_X1 U8017 ( .B1(n11640), .B2(n11639), .A(n6671), .ZN(n11713) );
  NOR2_X1 U8018 ( .A1(n11638), .A2(n11637), .ZN(n6671) );
  NAND2_X1 U8019 ( .A1(n10519), .A2(n6683), .ZN(n10589) );
  AND2_X1 U8020 ( .A1(n10520), .A2(n10518), .ZN(n6683) );
  AND3_X1 U8021 ( .A1(n9271), .A2(n9270), .A3(n9269), .ZN(n12813) );
  NAND2_X1 U8022 ( .A1(n12526), .A2(n12527), .ZN(n12525) );
  NAND2_X1 U8023 ( .A1(n9356), .A2(n9355), .ZN(n12200) );
  AND4_X1 U8024 ( .A1(n9119), .A2(n9118), .A3(n9117), .A4(n9116), .ZN(n15046)
         );
  OR2_X1 U8025 ( .A1(n6440), .A2(n10715), .ZN(n8978) );
  AND4_X1 U8026 ( .A1(n9015), .A2(n9014), .A3(n9013), .A4(n9012), .ZN(n12812)
         );
  AND4_X1 U8027 ( .A1(n9056), .A2(n9055), .A3(n9054), .A4(n9053), .ZN(n15086)
         );
  AOI21_X1 U8028 ( .B1(n9052), .B2(P3_REG1_REG_19__SCAN_IN), .A(n6593), .ZN(
        n9288) );
  AND4_X1 U8029 ( .A1(n9237), .A2(n9236), .A3(n9235), .A4(n9234), .ZN(n11751)
         );
  NAND2_X1 U8030 ( .A1(n9245), .A2(n9244), .ZN(n11754) );
  NAND2_X1 U8031 ( .A1(n15081), .A2(n10393), .ZN(n12521) );
  NAND2_X1 U8032 ( .A1(n9644), .A2(n10905), .ZN(n6963) );
  AOI21_X1 U8033 ( .B1(n12666), .B2(n9286), .A(n9362), .ZN(n12674) );
  INV_X1 U8034 ( .A(n12828), .ZN(n12547) );
  NAND2_X1 U8035 ( .A1(n9038), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9221) );
  XNOR2_X1 U8036 ( .A(n9074), .B(P3_IR_REG_4__SCAN_IN), .ZN(n14907) );
  AND2_X1 U8037 ( .A1(n14896), .A2(n14895), .ZN(n14898) );
  XNOR2_X1 U8038 ( .A(n7172), .B(n14975), .ZN(n14969) );
  NOR2_X1 U8039 ( .A1(n14969), .A2(n14970), .ZN(n14968) );
  XNOR2_X1 U8040 ( .A(n7161), .B(n15012), .ZN(n15007) );
  NOR2_X1 U8041 ( .A1(n15007), .A2(n15242), .ZN(n15006) );
  NAND2_X1 U8042 ( .A1(n7166), .A2(n6694), .ZN(n6693) );
  NAND2_X1 U8043 ( .A1(n14430), .A2(n14429), .ZN(n6694) );
  INV_X1 U8044 ( .A(n14912), .ZN(n15035) );
  AND2_X1 U8045 ( .A1(n10415), .A2(n10414), .ZN(n14866) );
  OR2_X1 U8046 ( .A1(n14430), .A2(n14429), .ZN(n7166) );
  NAND2_X1 U8047 ( .A1(n6995), .A2(n6993), .ZN(n6992) );
  AOI21_X1 U8048 ( .B1(n14992), .B2(n12659), .A(n6994), .ZN(n6993) );
  NAND2_X1 U8049 ( .A1(n6996), .A2(n15037), .ZN(n6995) );
  INV_X1 U8050 ( .A(n12633), .ZN(n6994) );
  NAND2_X1 U8051 ( .A1(n9657), .A2(n6591), .ZN(n12665) );
  NAND2_X1 U8052 ( .A1(n8960), .A2(n8959), .ZN(n12695) );
  INV_X1 U8053 ( .A(n9409), .ZN(n12726) );
  NAND2_X1 U8054 ( .A1(n9230), .A2(n9229), .ZN(n14456) );
  INV_X1 U8055 ( .A(n12200), .ZN(n12897) );
  AOI21_X1 U8056 ( .B1(n12669), .B2(n15101), .A(n12665), .ZN(n12895) );
  OR2_X1 U8057 ( .A1(n15142), .A2(n15136), .ZN(n12939) );
  NAND2_X1 U8058 ( .A1(n6936), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8958) );
  NAND2_X1 U8059 ( .A1(n9278), .A2(n8898), .ZN(n9375) );
  INV_X1 U8060 ( .A(n14420), .ZN(n12634) );
  OAI21_X1 U8061 ( .B1(n13286), .B2(n13114), .A(n9803), .ZN(n9804) );
  NOR2_X1 U8062 ( .A1(n6460), .A2(n13070), .ZN(n7430) );
  NAND2_X1 U8063 ( .A1(n7433), .A2(n7438), .ZN(n7432) );
  NAND2_X1 U8064 ( .A1(n7439), .A2(n12992), .ZN(n7438) );
  INV_X1 U8065 ( .A(n9783), .ZN(n7439) );
  NAND2_X1 U8066 ( .A1(n13089), .A2(n9779), .ZN(n9782) );
  INV_X1 U8067 ( .A(n7428), .ZN(n7427) );
  NAND2_X1 U8068 ( .A1(n9674), .A2(n9675), .ZN(n10041) );
  NAND2_X1 U8069 ( .A1(n13505), .A2(n13081), .ZN(n6875) );
  NAND2_X1 U8070 ( .A1(n7459), .A2(n7458), .ZN(n7457) );
  OR2_X1 U8071 ( .A1(n9685), .A2(n9686), .ZN(n9687) );
  INV_X1 U8072 ( .A(n11862), .ZN(n11865) );
  NAND2_X1 U8073 ( .A1(n11360), .A2(n7750), .ZN(n6786) );
  AND2_X1 U8074 ( .A1(n9682), .A2(n9681), .ZN(n10174) );
  INV_X1 U8075 ( .A(n13422), .ZN(n13541) );
  NAND2_X1 U8076 ( .A1(n8139), .A2(n8138), .ZN(n13119) );
  INV_X1 U8077 ( .A(n12023), .ZN(n13124) );
  OR2_X1 U8078 ( .A1(n13273), .A2(n13472), .ZN(n6862) );
  NAND2_X1 U8079 ( .A1(n13279), .A2(n8269), .ZN(n13470) );
  NAND2_X2 U8080 ( .A1(n14835), .A2(n8266), .ZN(n13472) );
  AOI21_X1 U8081 ( .B1(n13283), .B2(n6789), .A(n6543), .ZN(n6790) );
  CLKBUF_X1 U8082 ( .A(n13552), .Z(n14864) );
  INV_X1 U8083 ( .A(n13534), .ZN(n13558) );
  INV_X1 U8084 ( .A(n14864), .ZN(n14862) );
  AND2_X1 U8085 ( .A1(n8278), .A2(n7183), .ZN(n9662) );
  AND2_X1 U8086 ( .A1(n8271), .A2(n7184), .ZN(n7183) );
  NAND2_X1 U8087 ( .A1(n12058), .A2(n14845), .ZN(n7184) );
  NAND2_X1 U8088 ( .A1(n13567), .A2(n14859), .ZN(n6802) );
  NAND2_X1 U8089 ( .A1(n14858), .A2(n13568), .ZN(n6801) );
  NAND2_X1 U8090 ( .A1(n8225), .A2(n8224), .ZN(n14831) );
  NAND2_X1 U8092 ( .A1(n13656), .A2(n13657), .ZN(n13655) );
  AOI21_X1 U8093 ( .B1(n13777), .B2(n6664), .A(n12324), .ZN(n6663) );
  NOR2_X1 U8094 ( .A1(n13664), .A2(n14577), .ZN(n6836) );
  AND4_X1 U8095 ( .A1(n8539), .A2(n8538), .A3(n8537), .A4(n8536), .ZN(n12206)
         );
  AND2_X1 U8096 ( .A1(n8724), .A2(n8710), .ZN(n13945) );
  NAND2_X1 U8097 ( .A1(n6645), .A2(n6472), .ZN(n6651) );
  NAND2_X1 U8098 ( .A1(n14573), .A2(n14574), .ZN(n6645) );
  OR2_X1 U8099 ( .A1(n10279), .A2(n10278), .ZN(n14565) );
  AND2_X1 U8100 ( .A1(n14564), .A2(n14740), .ZN(n13739) );
  INV_X1 U8101 ( .A(n14565), .ZN(n14580) );
  INV_X1 U8102 ( .A(n13792), .ZN(n13803) );
  INV_X1 U8103 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n13893) );
  NAND2_X1 U8104 ( .A1(n12399), .A2(n6884), .ZN(n13917) );
  NOR2_X1 U8105 ( .A1(n12397), .A2(n6813), .ZN(n14090) );
  AND2_X1 U8106 ( .A1(n12398), .A2(n12400), .ZN(n6813) );
  AND2_X1 U8107 ( .A1(n13973), .A2(n12357), .ZN(n13954) );
  NAND2_X1 U8108 ( .A1(n6825), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6824) );
  INV_X1 U8109 ( .A(n14075), .ZN(n7226) );
  INV_X1 U8110 ( .A(n14078), .ZN(n6769) );
  NAND2_X1 U8111 ( .A1(n13906), .A2(n6771), .ZN(n6766) );
  OR2_X1 U8112 ( .A1(n13906), .A2(n12380), .ZN(n6767) );
  NOR2_X1 U8113 ( .A1(n12361), .A2(n6772), .ZN(n6771) );
  AOI21_X1 U8114 ( .B1(n8297), .B2(P1_IR_REG_31__SCAN_IN), .A(n6755), .ZN(
        n6754) );
  NAND2_X1 U8115 ( .A1(n15319), .A2(n15320), .ZN(n15318) );
  NAND2_X1 U8116 ( .A1(n7138), .A2(n7137), .ZN(n6616) );
  NOR2_X1 U8117 ( .A1(n14331), .A2(n14773), .ZN(n14330) );
  NAND2_X1 U8118 ( .A1(n14333), .A2(n7158), .ZN(n7156) );
  OAI21_X1 U8119 ( .B1(n7158), .B2(n7154), .A(n14541), .ZN(n7153) );
  XNOR2_X1 U8120 ( .A(n14296), .B(n6823), .ZN(n14544) );
  INV_X1 U8121 ( .A(n14295), .ZN(n6823) );
  OAI21_X1 U8122 ( .B1(n14546), .B2(n14547), .A(n7131), .ZN(n6618) );
  INV_X1 U8123 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7131) );
  OAI21_X1 U8124 ( .B1(n14560), .B2(n14559), .A(n6822), .ZN(n6617) );
  INV_X1 U8125 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n6822) );
  NAND2_X1 U8126 ( .A1(n11884), .A2(n6496), .ZN(n6749) );
  AND2_X1 U8127 ( .A1(n7411), .A2(n11906), .ZN(n7410) );
  NAND2_X1 U8128 ( .A1(n11901), .A2(n7413), .ZN(n7412) );
  INV_X1 U8129 ( .A(n11902), .ZN(n7413) );
  NAND2_X1 U8130 ( .A1(n8417), .A2(n7056), .ZN(n7055) );
  NAND2_X1 U8131 ( .A1(n8449), .A2(n7033), .ZN(n7032) );
  INV_X1 U8132 ( .A(n7032), .ZN(n7030) );
  NOR2_X1 U8133 ( .A1(n7420), .A2(n7421), .ZN(n7419) );
  NAND2_X1 U8134 ( .A1(n11911), .A2(n6745), .ZN(n11916) );
  INV_X1 U8135 ( .A(n11915), .ZN(n7421) );
  NAND2_X1 U8136 ( .A1(n8482), .A2(n7059), .ZN(n7058) );
  INV_X1 U8137 ( .A(n11963), .ZN(n7408) );
  NOR2_X1 U8138 ( .A1(n6471), .A2(n7043), .ZN(n7042) );
  AND2_X1 U8139 ( .A1(n7047), .A2(n7044), .ZN(n7043) );
  INV_X1 U8140 ( .A(n8610), .ZN(n7044) );
  OR2_X1 U8141 ( .A1(n8581), .A2(n8580), .ZN(n7047) );
  INV_X1 U8142 ( .A(n6957), .ZN(n6956) );
  NOR2_X1 U8143 ( .A1(n6985), .A2(n9147), .ZN(n6984) );
  INV_X1 U8144 ( .A(n9552), .ZN(n6985) );
  AOI21_X1 U8145 ( .B1(n11752), .B2(n6974), .A(n10398), .ZN(n6973) );
  AOI21_X1 U8146 ( .B1(n11752), .B2(n6451), .A(n6549), .ZN(n6972) );
  AOI21_X1 U8147 ( .B1(n6723), .B2(n6726), .A(n6544), .ZN(n6721) );
  NAND2_X1 U8148 ( .A1(n11957), .A2(n6723), .ZN(n6722) );
  AND2_X1 U8149 ( .A1(n11958), .A2(n6727), .ZN(n6726) );
  NOR2_X1 U8150 ( .A1(n6952), .A2(n9573), .ZN(n6951) );
  NOR2_X1 U8151 ( .A1(n6954), .A2(n6475), .ZN(n6952) );
  AOI21_X1 U8152 ( .B1(n6957), .B2(n6959), .A(n6955), .ZN(n6954) );
  INV_X1 U8153 ( .A(n6973), .ZN(n6970) );
  INV_X1 U8154 ( .A(n6972), .ZN(n6971) );
  OR3_X1 U8155 ( .A1(n11999), .A2(n11998), .A3(n11997), .ZN(n12004) );
  OAI22_X1 U8156 ( .A1(n11972), .A2(n11971), .B1(n11989), .B2(n11988), .ZN(
        n11974) );
  AOI21_X1 U8157 ( .B1(n6967), .B2(n6968), .A(n6966), .ZN(n6965) );
  AND2_X1 U8158 ( .A1(n7361), .A2(n7360), .ZN(n8684) );
  OR2_X1 U8159 ( .A1(n6899), .A2(n8806), .ZN(n7360) );
  NAND2_X1 U8160 ( .A1(n14206), .A2(n7362), .ZN(n7361) );
  NOR2_X1 U8161 ( .A1(n8800), .A2(n8637), .ZN(n7362) );
  NAND2_X1 U8162 ( .A1(n7418), .A2(n7417), .ZN(n7416) );
  INV_X1 U8163 ( .A(n7415), .ZN(n6741) );
  OAI21_X1 U8164 ( .B1(n8685), .B2(n8684), .A(n7356), .ZN(n7355) );
  NAND2_X1 U8165 ( .A1(n7358), .A2(n7357), .ZN(n7356) );
  OR2_X1 U8166 ( .A1(n6899), .A2(n8800), .ZN(n7357) );
  NAND2_X1 U8167 ( .A1(n14206), .A2(n7359), .ZN(n7358) );
  NOR2_X1 U8168 ( .A1(n12034), .A2(n12033), .ZN(n6731) );
  NAND2_X1 U8169 ( .A1(n7397), .A2(n12029), .ZN(n7396) );
  NOR2_X1 U8170 ( .A1(n6731), .A2(n12039), .ZN(n6729) );
  NAND2_X1 U8171 ( .A1(n8720), .A2(n7382), .ZN(n7381) );
  INV_X1 U8172 ( .A(n12044), .ZN(n6720) );
  XNOR2_X1 U8173 ( .A(n8883), .B(n8820), .ZN(n8329) );
  INV_X1 U8174 ( .A(n7563), .ZN(n7064) );
  INV_X1 U8175 ( .A(n7065), .ZN(n6879) );
  NAND2_X1 U8176 ( .A1(n6943), .A2(n9630), .ZN(n6942) );
  OAI21_X1 U8177 ( .B1(n9627), .B2(n12708), .A(n6944), .ZN(n6943) );
  AND2_X1 U8178 ( .A1(n12688), .A2(n9626), .ZN(n6944) );
  INV_X1 U8179 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8897) );
  INV_X1 U8180 ( .A(n12078), .ZN(n7389) );
  AOI21_X1 U8181 ( .B1(n6449), .B2(n7052), .A(n6547), .ZN(n7049) );
  AND2_X1 U8182 ( .A1(n8736), .A2(n7053), .ZN(n7052) );
  INV_X1 U8183 ( .A(n12378), .ZN(n7337) );
  NAND2_X1 U8184 ( .A1(n7665), .A2(n7083), .ZN(n7082) );
  OAI21_X1 U8185 ( .B1(n8039), .B2(n6598), .A(n6886), .ZN(n7660) );
  NAND2_X1 U8186 ( .A1(n7092), .A2(n7091), .ZN(n7090) );
  INV_X1 U8187 ( .A(n7653), .ZN(n7092) );
  INV_X1 U8188 ( .A(n7611), .ZN(n7368) );
  OAI21_X1 U8189 ( .B1(n6465), .B2(n7600), .A(n6785), .ZN(n7349) );
  INV_X1 U8190 ( .A(n7797), .ZN(n6785) );
  NOR2_X1 U8191 ( .A1(n7354), .A2(n6465), .ZN(n7353) );
  AND2_X1 U8192 ( .A1(n7146), .A2(n7157), .ZN(n7155) );
  INV_X1 U8193 ( .A(n14541), .ZN(n7146) );
  NAND2_X1 U8194 ( .A1(n6939), .A2(n6938), .ZN(n9638) );
  NAND2_X1 U8195 ( .A1(n6941), .A2(n6940), .ZN(n6939) );
  NAND2_X1 U8196 ( .A1(n12682), .A2(n9631), .ZN(n6940) );
  NAND2_X1 U8197 ( .A1(n6942), .A2(n12679), .ZN(n6941) );
  NAND2_X1 U8198 ( .A1(n10434), .A2(n6855), .ZN(n10436) );
  OR2_X1 U8199 ( .A1(n14907), .A2(n10435), .ZN(n6855) );
  NAND2_X1 U8200 ( .A1(n15038), .A2(n12619), .ZN(n12620) );
  AND2_X1 U8201 ( .A1(n6480), .A2(n7316), .ZN(n7315) );
  INV_X1 U8202 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7316) );
  OR2_X1 U8203 ( .A1(n9357), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9368) );
  NOR2_X1 U8204 ( .A1(n7572), .A2(n7486), .ZN(n7485) );
  INV_X1 U8205 ( .A(n7492), .ZN(n7486) );
  INV_X1 U8206 ( .A(n7487), .ZN(n7484) );
  NAND2_X1 U8207 ( .A1(n12773), .A2(n7505), .ZN(n7504) );
  INV_X1 U8208 ( .A(n9291), .ZN(n7505) );
  AND2_X1 U8209 ( .A1(n9607), .A2(n9608), .ZN(n9606) );
  NOR2_X1 U8210 ( .A1(n9011), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9267) );
  OR2_X1 U8211 ( .A1(n9249), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9011) );
  INV_X1 U8212 ( .A(n7497), .ZN(n7496) );
  OAI21_X1 U8213 ( .B1(n7499), .B2(n7498), .A(n11748), .ZN(n7497) );
  INV_X1 U8214 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n9246) );
  NAND2_X1 U8215 ( .A1(n9247), .A2(n9246), .ZN(n9249) );
  AND2_X1 U8216 ( .A1(n9216), .A2(n9215), .ZN(n9232) );
  NOR2_X1 U8217 ( .A1(n10717), .A2(n7115), .ZN(n7110) );
  NAND2_X1 U8218 ( .A1(n7126), .A2(n7124), .ZN(n9488) );
  INV_X1 U8219 ( .A(n7125), .ZN(n7124) );
  OAI21_X1 U8220 ( .B1(n6481), .B2(n9634), .A(n9632), .ZN(n7125) );
  INV_X1 U8221 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8950) );
  INV_X1 U8222 ( .A(n7249), .ZN(n6635) );
  INV_X1 U8223 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8948) );
  INV_X1 U8224 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n8941) );
  AND2_X1 U8225 ( .A1(n8987), .A2(n7315), .ZN(n8989) );
  NAND2_X1 U8226 ( .A1(n12986), .A2(n9783), .ZN(n7437) );
  NOR2_X1 U8227 ( .A1(n7968), .A2(n13106), .ZN(n7979) );
  NAND2_X1 U8228 ( .A1(n13023), .A2(n13024), .ZN(n7445) );
  INV_X1 U8229 ( .A(n12976), .ZN(n7447) );
  XNOR2_X1 U8230 ( .A(n9676), .B(n11869), .ZN(n9673) );
  NAND2_X1 U8231 ( .A1(n13011), .A2(n9774), .ZN(n7461) );
  INV_X1 U8232 ( .A(n13037), .ZN(n6710) );
  NAND2_X1 U8233 ( .A1(n9774), .A2(n9770), .ZN(n7462) );
  INV_X1 U8234 ( .A(n7462), .ZN(n6712) );
  INV_X1 U8235 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7697) );
  OR2_X1 U8236 ( .A1(n8161), .A2(n8160), .ZN(n8171) );
  NOR2_X1 U8237 ( .A1(n6810), .A2(n6533), .ZN(n6808) );
  INV_X1 U8238 ( .A(n7956), .ZN(n6809) );
  NAND2_X1 U8239 ( .A1(n7880), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7900) );
  INV_X1 U8240 ( .A(n7882), .ZN(n7880) );
  OR2_X1 U8241 ( .A1(n12115), .A2(n7198), .ZN(n7197) );
  NAND2_X1 U8242 ( .A1(n13272), .A2(n13271), .ZN(n6846) );
  NOR2_X1 U8243 ( .A1(n8258), .A2(n7203), .ZN(n7202) );
  INV_X1 U8244 ( .A(n8257), .ZN(n7203) );
  NAND2_X1 U8245 ( .A1(n7202), .A2(n7200), .ZN(n7199) );
  INV_X1 U8246 ( .A(n7205), .ZN(n7200) );
  INV_X1 U8247 ( .A(n8236), .ZN(n7209) );
  AND2_X1 U8248 ( .A1(n8707), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8722) );
  AND2_X1 U8249 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n8691), .ZN(n8707) );
  INV_X1 U8250 ( .A(n13748), .ZN(n6654) );
  NOR2_X1 U8251 ( .A1(n7372), .A2(n8776), .ZN(n7373) );
  INV_X1 U8252 ( .A(n8809), .ZN(n7371) );
  NAND2_X1 U8253 ( .A1(n6538), .A2(n8809), .ZN(n7369) );
  INV_X1 U8254 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8316) );
  INV_X1 U8255 ( .A(n7260), .ZN(n7259) );
  AND2_X1 U8256 ( .A1(n11806), .A2(n6557), .ZN(n6765) );
  NOR2_X1 U8257 ( .A1(n14336), .A2(n6918), .ZN(n6917) );
  NAND2_X1 U8258 ( .A1(n14156), .A2(n6919), .ZN(n6918) );
  INV_X1 U8259 ( .A(n6920), .ZN(n6919) );
  INV_X1 U8260 ( .A(n11626), .ZN(n7262) );
  NAND2_X1 U8261 ( .A1(n11724), .A2(n11723), .ZN(n11812) );
  OR2_X1 U8262 ( .A1(n12222), .A2(n12214), .ZN(n6920) );
  NAND2_X1 U8263 ( .A1(n11486), .A2(n11851), .ZN(n11592) );
  NAND2_X1 U8264 ( .A1(n11153), .A2(n11323), .ZN(n7333) );
  AND2_X1 U8265 ( .A1(n11333), .A2(n14532), .ZN(n11486) );
  NOR2_X1 U8266 ( .A1(n13909), .A2(n14082), .ZN(n7230) );
  NAND2_X1 U8267 ( .A1(n7223), .A2(n12260), .ZN(n14028) );
  NAND2_X1 U8268 ( .A1(n10750), .A2(n10749), .ZN(n10821) );
  AOI21_X1 U8269 ( .B1(n10322), .B2(n10227), .A(n10226), .ZN(n10289) );
  OR2_X1 U8270 ( .A1(n8811), .A2(n12948), .ZN(n8812) );
  INV_X1 U8271 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n7034) );
  INV_X1 U8272 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n7035) );
  INV_X1 U8273 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n7540) );
  NAND2_X1 U8274 ( .A1(n7385), .A2(n7386), .ZN(n7085) );
  INV_X1 U8275 ( .A(n7660), .ZN(n7385) );
  NAND2_X1 U8276 ( .A1(n7660), .A2(SI_22_), .ZN(n7086) );
  XNOR2_X1 U8277 ( .A(n7653), .B(SI_19_), .ZN(n8022) );
  NAND2_X1 U8278 ( .A1(n6890), .A2(n6891), .ZN(n7652) );
  AND2_X1 U8279 ( .A1(n6892), .A2(n6894), .ZN(n6891) );
  INV_X1 U8280 ( .A(n6895), .ZN(n6894) );
  AND2_X1 U8281 ( .A1(n6576), .A2(n7375), .ZN(n7078) );
  INV_X1 U8282 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8315) );
  INV_X1 U8283 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8540) );
  INV_X1 U8284 ( .A(SI_11_), .ZN(n9188) );
  OR2_X1 U8285 ( .A1(n8511), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n8527) );
  INV_X1 U8286 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8283) );
  NOR2_X1 U8287 ( .A1(n14213), .A2(n14212), .ZN(n14215) );
  AND2_X1 U8288 ( .A1(n10333), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n14212) );
  AOI21_X1 U8289 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n14228), .A(n14227), .ZN(
        n14289) );
  AOI21_X1 U8290 ( .B1(n7155), .B2(n7150), .A(P2_ADDR_REG_11__SCAN_IN), .ZN(
        n7149) );
  INV_X1 U8291 ( .A(n7158), .ZN(n7150) );
  INV_X1 U8292 ( .A(n7155), .ZN(n7151) );
  OR2_X1 U8293 ( .A1(n9163), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9178) );
  NOR2_X1 U8294 ( .A1(n9113), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9130) );
  INV_X1 U8295 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10556) );
  NAND2_X1 U8296 ( .A1(n12495), .A2(n12494), .ZN(n7298) );
  NAND2_X1 U8297 ( .A1(n12186), .A2(n12467), .ZN(n12469) );
  AND3_X1 U8298 ( .A1(n9095), .A2(n9094), .A3(n9093), .ZN(n10811) );
  INV_X1 U8299 ( .A(n10808), .ZN(n7311) );
  OR2_X1 U8300 ( .A1(n10807), .A2(n10806), .ZN(n7312) );
  INV_X1 U8301 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9080) );
  OR2_X1 U8302 ( .A1(n9319), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9328) );
  NAND2_X1 U8303 ( .A1(n7307), .A2(n7306), .ZN(n11341) );
  INV_X1 U8304 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n9150) );
  AOI21_X1 U8305 ( .B1(n7295), .B2(n7294), .A(n7293), .ZN(n7292) );
  INV_X1 U8306 ( .A(n12173), .ZN(n7293) );
  INV_X1 U8307 ( .A(n12494), .ZN(n7294) );
  NAND2_X1 U8308 ( .A1(n12175), .A2(n12174), .ZN(n12176) );
  OR2_X1 U8309 ( .A1(n12503), .A2(n12758), .ZN(n12501) );
  NAND2_X1 U8310 ( .A1(n11341), .A2(n7545), .ZN(n11368) );
  XNOR2_X1 U8311 ( .A(n10487), .B(n15077), .ZN(n10517) );
  OR2_X1 U8312 ( .A1(n12476), .A2(n12545), .ZN(n12161) );
  NOR2_X1 U8313 ( .A1(n6638), .A2(n9639), .ZN(n6637) );
  NOR2_X1 U8314 ( .A1(n9515), .A2(n9514), .ZN(n6866) );
  INV_X1 U8315 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10416) );
  INV_X1 U8316 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n14214) );
  NAND2_X1 U8317 ( .A1(n9061), .A2(n9073), .ZN(n9090) );
  INV_X1 U8318 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n9073) );
  XNOR2_X1 U8319 ( .A(n10436), .B(n6854), .ZN(n14927) );
  NAND2_X1 U8320 ( .A1(n7021), .A2(n7022), .ZN(n7018) );
  INV_X1 U8321 ( .A(n10531), .ZN(n7168) );
  NAND2_X1 U8322 ( .A1(n6870), .A2(n6869), .ZN(n12581) );
  INV_X1 U8323 ( .A(n10537), .ZN(n6869) );
  NAND2_X1 U8324 ( .A1(n12581), .A2(n12580), .ZN(n6847) );
  NAND2_X1 U8325 ( .A1(n12606), .A2(n12607), .ZN(n14978) );
  XNOR2_X1 U8326 ( .A(n12645), .B(n12613), .ZN(n15009) );
  INV_X1 U8327 ( .A(n14386), .ZN(n7170) );
  NAND2_X1 U8328 ( .A1(n6689), .A2(n6688), .ZN(n7171) );
  XNOR2_X1 U8329 ( .A(n6998), .B(n6997), .ZN(n6996) );
  INV_X1 U8330 ( .A(n12631), .ZN(n6997) );
  NAND2_X1 U8331 ( .A1(n14424), .A2(n12630), .ZN(n6998) );
  NAND2_X1 U8332 ( .A1(n9038), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n9387) );
  OR2_X1 U8333 ( .A1(n12897), .A2(n12674), .ZN(n7567) );
  AND2_X1 U8334 ( .A1(n9629), .A2(n9628), .ZN(n12688) );
  NAND2_X1 U8335 ( .A1(n12733), .A2(n12737), .ZN(n12732) );
  NAND2_X1 U8336 ( .A1(n12755), .A2(n6817), .ZN(n12745) );
  NAND2_X1 U8337 ( .A1(n6818), .A2(n12769), .ZN(n6817) );
  NAND2_X1 U8338 ( .A1(n9407), .A2(n9607), .ZN(n12749) );
  NAND2_X1 U8339 ( .A1(n12761), .A2(n9608), .ZN(n9407) );
  INV_X1 U8340 ( .A(n9298), .ZN(n8889) );
  INV_X1 U8341 ( .A(n9606), .ZN(n12760) );
  INV_X1 U8342 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n12451) );
  NAND2_X1 U8343 ( .A1(n9284), .A2(n12451), .ZN(n9296) );
  AND2_X1 U8344 ( .A1(n12792), .A2(n9274), .ZN(n12781) );
  AND4_X1 U8345 ( .A1(n9001), .A2(n9000), .A3(n8999), .A4(n8998), .ZN(n12829)
         );
  AOI21_X1 U8346 ( .B1(n7475), .B2(n7478), .A(n6589), .ZN(n7473) );
  INV_X1 U8347 ( .A(n9565), .ZN(n6921) );
  INV_X1 U8348 ( .A(n11044), .ZN(n9148) );
  AND2_X1 U8349 ( .A1(n11042), .A2(n9149), .ZN(n11175) );
  NAND2_X1 U8350 ( .A1(n10717), .A2(n10718), .ZN(n7111) );
  AOI21_X1 U8351 ( .B1(n15083), .B2(n15082), .A(n7548), .ZN(n10726) );
  NAND2_X1 U8352 ( .A1(n10726), .A2(n7114), .ZN(n10725) );
  AND2_X1 U8353 ( .A1(n9412), .A2(n9455), .ZN(n15093) );
  NAND2_X1 U8354 ( .A1(n9341), .A2(n9340), .ZN(n12839) );
  NAND2_X1 U8355 ( .A1(n8974), .A2(n8973), .ZN(n12847) );
  AND2_X1 U8356 ( .A1(n15093), .A2(n15137), .ZN(n14458) );
  INV_X1 U8357 ( .A(n14458), .ZN(n15101) );
  AOI21_X1 U8358 ( .B1(n6680), .B2(n11525), .A(n6679), .ZN(n9973) );
  XNOR2_X1 U8359 ( .A(n11400), .B(P3_B_REG_SCAN_IN), .ZN(n6680) );
  NOR2_X1 U8360 ( .A1(n9225), .A2(n8901), .ZN(n6819) );
  INV_X1 U8361 ( .A(n12944), .ZN(n8905) );
  INV_X1 U8362 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8957) );
  AND3_X1 U8363 ( .A1(n7501), .A2(n8987), .A3(n7500), .ZN(n9416) );
  NAND2_X1 U8364 ( .A1(n7501), .A2(n8987), .ZN(n9418) );
  XNOR2_X1 U8365 ( .A(n6684), .B(P3_IR_REG_24__SCAN_IN), .ZN(n9421) );
  NAND2_X1 U8366 ( .A1(n6685), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6684) );
  NAND2_X1 U8367 ( .A1(n8987), .A2(n8899), .ZN(n6685) );
  NAND2_X1 U8368 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n6640), .ZN(n6639) );
  NAND2_X1 U8369 ( .A1(n9259), .A2(n9258), .ZN(n6641) );
  NAND2_X1 U8370 ( .A1(n8987), .A2(n6480), .ZN(n9005) );
  AOI21_X1 U8371 ( .B1(n7245), .B2(n9239), .A(n6597), .ZN(n7244) );
  XNOR2_X1 U8372 ( .A(n8936), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9208) );
  AND2_X1 U8373 ( .A1(n15289), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8933) );
  OR2_X1 U8374 ( .A1(n9171), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n9186) );
  AOI21_X1 U8375 ( .B1(n7233), .B2(n6454), .A(n6539), .ZN(n7232) );
  AND2_X1 U8376 ( .A1(n9123), .A2(n9122), .ZN(n9139) );
  OR2_X1 U8377 ( .A1(n9090), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n9106) );
  XNOR2_X1 U8378 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n9071) );
  NAND2_X1 U8379 ( .A1(n8919), .A2(n8918), .ZN(n9021) );
  NAND2_X1 U8380 ( .A1(n6851), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9022) );
  XNOR2_X1 U8381 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9030) );
  OAI21_X1 U8382 ( .B1(n11574), .B2(n6532), .A(n7463), .ZN(n11785) );
  NAND2_X1 U8383 ( .A1(n7464), .A2(n9734), .ZN(n7463) );
  INV_X1 U8384 ( .A(n7465), .ZN(n7464) );
  NAND2_X1 U8385 ( .A1(n11785), .A2(n11784), .ZN(n11783) );
  OR2_X1 U8386 ( .A1(n7947), .A2(n11787), .ZN(n7968) );
  NAND2_X1 U8387 ( .A1(n13056), .A2(n9765), .ZN(n9766) );
  NAND2_X1 U8388 ( .A1(n6706), .A2(n6703), .ZN(n6702) );
  INV_X1 U8389 ( .A(n13048), .ZN(n6706) );
  OR2_X1 U8390 ( .A1(n7900), .A2(n7899), .ZN(n7914) );
  NAND2_X1 U8391 ( .A1(n6821), .A2(n9741), .ZN(n7555) );
  INV_X1 U8392 ( .A(n9742), .ZN(n6821) );
  NAND2_X1 U8393 ( .A1(n7979), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7996) );
  INV_X1 U8394 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n13030) );
  XNOR2_X1 U8395 ( .A(n9676), .B(n6828), .ZN(n9684) );
  INV_X1 U8396 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7865) );
  OR2_X1 U8397 ( .A1(n7866), .A2(n7865), .ZN(n7882) );
  NOR2_X1 U8398 ( .A1(n11659), .A2(n7466), .ZN(n7465) );
  INV_X1 U8399 ( .A(n9728), .ZN(n7466) );
  INV_X1 U8400 ( .A(n13122), .ZN(n12030) );
  NAND2_X1 U8401 ( .A1(n7449), .A2(n7448), .ZN(n7442) );
  OR2_X1 U8402 ( .A1(n7996), .A2(n13030), .ZN(n8011) );
  NAND2_X1 U8403 ( .A1(n6711), .A2(n6708), .ZN(n13088) );
  INV_X1 U8404 ( .A(n6709), .ZN(n6708) );
  NAND2_X1 U8405 ( .A1(n13038), .A2(n6712), .ZN(n6711) );
  OAI21_X1 U8406 ( .B1(n7462), .B2(n6710), .A(n7461), .ZN(n6709) );
  INV_X1 U8407 ( .A(n13094), .ZN(n13061) );
  NOR2_X1 U8408 ( .A1(n6831), .A2(n6830), .ZN(n6829) );
  INV_X1 U8409 ( .A(n8222), .ZN(n12103) );
  NAND2_X1 U8410 ( .A1(n6716), .A2(n12088), .ZN(n12098) );
  AND2_X1 U8411 ( .A1(n8064), .A2(n8063), .ZN(n13059) );
  AND2_X1 U8412 ( .A1(n8050), .A2(n8049), .ZN(n12023) );
  OR2_X1 U8413 ( .A1(n14762), .A2(n14761), .ZN(n14764) );
  NAND2_X1 U8414 ( .A1(n6554), .A2(n12060), .ZN(n13255) );
  AND2_X1 U8415 ( .A1(n6783), .A2(n13312), .ZN(n6780) );
  AND2_X1 U8416 ( .A1(n8133), .A2(n8121), .ZN(n13318) );
  NAND2_X1 U8417 ( .A1(n13330), .A2(n13320), .ZN(n13315) );
  NAND2_X1 U8418 ( .A1(n8072), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8093) );
  INV_X1 U8419 ( .A(n8074), .ZN(n8072) );
  NOR2_X1 U8420 ( .A1(n13591), .A2(n13526), .ZN(n7106) );
  NAND2_X1 U8421 ( .A1(n13385), .A2(n13376), .ZN(n13371) );
  OAI21_X1 U8422 ( .B1(n13437), .B2(n7212), .A(n7211), .ZN(n13399) );
  AOI21_X1 U8423 ( .B1(n7213), .B2(n13431), .A(n6524), .ZN(n7211) );
  INV_X1 U8424 ( .A(n7213), .ZN(n7212) );
  NOR2_X1 U8425 ( .A1(n11978), .A2(n13458), .ZN(n13443) );
  NAND2_X1 U8426 ( .A1(n7108), .A2(n7107), .ZN(n13458) );
  NAND2_X1 U8427 ( .A1(n7912), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7929) );
  INV_X1 U8428 ( .A(n7914), .ZN(n7912) );
  OR2_X1 U8429 ( .A1(n7929), .A2(n10315), .ZN(n7947) );
  NAND2_X1 U8430 ( .A1(n11284), .A2(n7890), .ZN(n11445) );
  NAND2_X1 U8431 ( .A1(n11235), .A2(n7872), .ZN(n11286) );
  NAND2_X1 U8432 ( .A1(n10990), .A2(n12115), .ZN(n10989) );
  NAND2_X1 U8433 ( .A1(n10600), .A2(n7796), .ZN(n11030) );
  NAND2_X1 U8434 ( .A1(n11030), .A2(n12111), .ZN(n11029) );
  NAND2_X1 U8435 ( .A1(n10775), .A2(n10707), .ZN(n11036) );
  NOR2_X1 U8436 ( .A1(n11907), .A2(n7097), .ZN(n7096) );
  INV_X1 U8437 ( .A(n7098), .ZN(n7097) );
  NAND2_X1 U8438 ( .A1(n10601), .A2(n12110), .ZN(n10600) );
  INV_X1 U8439 ( .A(n10769), .ZN(n12108) );
  NAND2_X1 U8440 ( .A1(n10345), .A2(n7765), .ZN(n10770) );
  XNOR2_X1 U8441 ( .A(n13141), .B(n6828), .ZN(n10346) );
  NAND2_X1 U8442 ( .A1(n10347), .A2(n10346), .ZN(n10345) );
  NAND2_X1 U8443 ( .A1(n9892), .A2(n13653), .ZN(n6814) );
  NAND2_X1 U8444 ( .A1(n6715), .A2(n6714), .ZN(n6713) );
  INV_X1 U8445 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6714) );
  NAND2_X1 U8446 ( .A1(n12138), .A2(n12089), .ZN(n10141) );
  NOR2_X1 U8447 ( .A1(n13280), .A2(n13454), .ZN(n6789) );
  OAI21_X1 U8448 ( .B1(n11683), .B2(n8242), .A(n8243), .ZN(n11766) );
  NAND2_X1 U8449 ( .A1(n7928), .A2(n7927), .ZN(n11969) );
  INV_X1 U8450 ( .A(n10346), .ZN(n12107) );
  NAND2_X1 U8451 ( .A1(n9668), .A2(n11860), .ZN(n14850) );
  NAND2_X1 U8452 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), 
        .ZN(n6797) );
  OR2_X1 U8453 ( .A1(n7550), .A2(n6797), .ZN(n6796) );
  NAND2_X1 U8454 ( .A1(n7688), .A2(n7711), .ZN(n6795) );
  NAND3_X1 U8455 ( .A1(n7085), .A2(n8066), .A3(n7086), .ZN(n8069) );
  OAI21_X1 U8456 ( .B1(n7991), .B2(n7691), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n7693) );
  NAND2_X1 U8457 ( .A1(n7708), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7709) );
  OR2_X1 U8458 ( .A1(n7942), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n7975) );
  OR2_X1 U8459 ( .A1(n7991), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n7925) );
  NOR2_X1 U8460 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n7425) );
  INV_X1 U8461 ( .A(n7680), .ZN(n7424) );
  INV_X1 U8462 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8917) );
  NAND2_X1 U8463 ( .A1(n7595), .A2(SI_0_), .ZN(n9046) );
  AND2_X1 U8464 ( .A1(n10933), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9806) );
  INV_X1 U8465 ( .A(n12311), .ZN(n6664) );
  INV_X1 U8466 ( .A(n13777), .ZN(n6665) );
  AND2_X1 U8467 ( .A1(n13727), .A2(n12291), .ZN(n13667) );
  INV_X1 U8468 ( .A(n8678), .ZN(n8309) );
  AOI21_X1 U8469 ( .B1(n13657), .B2(n12324), .A(n12332), .ZN(n7515) );
  NAND2_X1 U8470 ( .A1(n11189), .A2(n7527), .ZN(n7523) );
  NAND2_X1 U8471 ( .A1(n13737), .A2(n13738), .ZN(n7537) );
  NAND2_X1 U8472 ( .A1(n14506), .A2(n11838), .ZN(n7532) );
  NAND2_X1 U8473 ( .A1(n13786), .A2(n7538), .ZN(n13705) );
  NAND2_X1 U8474 ( .A1(n12287), .A2(n12288), .ZN(n13727) );
  NOR2_X1 U8475 ( .A1(n15301), .A2(n8309), .ZN(n8691) );
  OAI21_X1 U8476 ( .B1(n6647), .B2(n7562), .A(n6646), .ZN(n11011) );
  OAI21_X1 U8477 ( .B1(n11189), .B2(n7521), .A(n7517), .ZN(n6667) );
  INV_X1 U8478 ( .A(n11552), .ZN(n7518) );
  INV_X1 U8479 ( .A(n7527), .ZN(n7519) );
  AND2_X1 U8480 ( .A1(n8532), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8566) );
  AND2_X1 U8481 ( .A1(n13666), .A2(n12282), .ZN(n13759) );
  INV_X1 U8482 ( .A(n7532), .ZN(n14508) );
  NAND2_X1 U8483 ( .A1(n10356), .A2(n10355), .ZN(n14574) );
  NAND2_X1 U8484 ( .A1(n6658), .A2(n6656), .ZN(n13676) );
  NOR2_X1 U8485 ( .A1(n13768), .A2(n6657), .ZN(n6656) );
  INV_X1 U8486 ( .A(n12242), .ZN(n6657) );
  NAND2_X1 U8487 ( .A1(n12310), .A2(n13695), .ZN(n13697) );
  INV_X1 U8488 ( .A(n10675), .ZN(n7073) );
  OR2_X1 U8489 ( .A1(n8788), .A2(n8354), .ZN(n8355) );
  NAND2_X1 U8490 ( .A1(n6759), .A2(n6758), .ZN(n10357) );
  INV_X1 U8491 ( .A(n6848), .ZN(n6758) );
  NOR2_X2 U8492 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n8360) );
  AOI21_X1 U8493 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n13832), .A(n10009), .ZN(
        n10010) );
  AOI21_X1 U8494 ( .B1(n10159), .B2(P1_REG1_REG_7__SCAN_IN), .A(n10155), .ZN(
        n10060) );
  INV_X1 U8495 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10214) );
  AOI21_X1 U8496 ( .B1(n11269), .B2(P1_REG1_REG_13__SCAN_IN), .A(n11268), .ZN(
        n13848) );
  XNOR2_X1 U8497 ( .A(n11495), .B(n11504), .ZN(n11271) );
  NAND2_X1 U8498 ( .A1(n11271), .A2(n11270), .ZN(n11497) );
  NAND2_X1 U8499 ( .A1(n8317), .A2(n8288), .ZN(n8611) );
  INV_X1 U8500 ( .A(n8599), .ZN(n8317) );
  AND2_X1 U8501 ( .A1(n12385), .A2(n8753), .ZN(n13912) );
  AND2_X1 U8502 ( .A1(n13940), .A2(n13959), .ZN(n7260) );
  NAND2_X1 U8503 ( .A1(n13952), .A2(n12359), .ZN(n13938) );
  NOR2_X1 U8504 ( .A1(n13938), .A2(n13939), .ZN(n13937) );
  AND2_X1 U8505 ( .A1(n13974), .A2(n12375), .ZN(n13957) );
  OR2_X1 U8506 ( .A1(n11747), .A2(n8359), .ZN(n8300) );
  NAND2_X1 U8507 ( .A1(n6619), .A2(n12373), .ZN(n13975) );
  NAND2_X1 U8508 ( .A1(n7331), .A2(n6492), .ZN(n6619) );
  NAND2_X1 U8509 ( .A1(n13975), .A2(n13976), .ZN(n13974) );
  INV_X1 U8510 ( .A(n14119), .ZN(n6910) );
  INV_X1 U8511 ( .A(n14005), .ZN(n6753) );
  NOR2_X1 U8512 ( .A1(n14059), .A2(n14144), .ZN(n14057) );
  NAND2_X1 U8513 ( .A1(n14057), .A2(n14136), .ZN(n14037) );
  NAND2_X1 U8514 ( .A1(n6632), .A2(n6631), .ZN(n7574) );
  NAND2_X1 U8515 ( .A1(n7328), .A2(n12365), .ZN(n6631) );
  OR2_X1 U8516 ( .A1(n8616), .A2(n8308), .ZN(n8641) );
  INV_X1 U8517 ( .A(n12364), .ZN(n14048) );
  NAND2_X1 U8518 ( .A1(n12363), .A2(n12362), .ZN(n14049) );
  NAND2_X1 U8519 ( .A1(n8582), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8616) );
  NAND2_X1 U8520 ( .A1(n11812), .A2(n11811), .ZN(n12363) );
  INV_X1 U8521 ( .A(n6917), .ZN(n11816) );
  NAND2_X1 U8522 ( .A1(n14346), .A2(n7264), .ZN(n7263) );
  NOR2_X1 U8523 ( .A1(n11627), .A2(n7265), .ZN(n7264) );
  INV_X1 U8524 ( .A(n11590), .ZN(n7265) );
  NOR2_X1 U8525 ( .A1(n14336), .A2(n6920), .ZN(n11732) );
  OAI21_X1 U8526 ( .B1(n11586), .B2(n6626), .A(n6624), .ZN(n11720) );
  AOI21_X1 U8527 ( .B1(n7323), .B2(n6503), .A(n6625), .ZN(n6624) );
  NOR2_X1 U8528 ( .A1(n11591), .A2(n7324), .ZN(n7323) );
  OR2_X1 U8529 ( .A1(n11592), .A2(n14343), .ZN(n14336) );
  NAND2_X1 U8530 ( .A1(n6752), .A2(n7252), .ZN(n11476) );
  AOI21_X1 U8531 ( .B1(n7253), .B2(n7255), .A(n6520), .ZN(n7252) );
  NOR2_X1 U8532 ( .A1(n11332), .A2(n14491), .ZN(n11333) );
  NAND2_X1 U8533 ( .A1(n11324), .A2(n11323), .ZN(n11479) );
  OR2_X1 U8534 ( .A1(n11147), .A2(n11153), .ZN(n11324) );
  NAND2_X1 U8535 ( .A1(n6901), .A2(n6900), .ZN(n11332) );
  INV_X1 U8536 ( .A(n11256), .ZN(n6901) );
  NAND2_X1 U8537 ( .A1(n6620), .A2(n7341), .ZN(n11248) );
  NAND2_X1 U8538 ( .A1(n6552), .A2(n6450), .ZN(n7341) );
  NAND2_X1 U8539 ( .A1(n11080), .A2(n6493), .ZN(n6620) );
  AND2_X1 U8540 ( .A1(n11077), .A2(n14712), .ZN(n11155) );
  NAND2_X1 U8541 ( .A1(n10976), .A2(n10975), .ZN(n11075) );
  NAND2_X1 U8542 ( .A1(n7325), .A2(n6627), .ZN(n10968) );
  AOI21_X1 U8543 ( .B1(n7326), .B2(n10862), .A(n6485), .ZN(n7325) );
  NAND2_X1 U8544 ( .A1(n10955), .A2(n6497), .ZN(n6627) );
  NOR2_X1 U8545 ( .A1(n6907), .A2(n10949), .ZN(n10870) );
  NOR2_X1 U8546 ( .A1(n6906), .A2(n11019), .ZN(n6905) );
  NAND2_X1 U8547 ( .A1(n10818), .A2(n10817), .ZN(n10948) );
  OR2_X1 U8548 ( .A1(n10948), .A2(n10949), .ZN(n10946) );
  AND2_X1 U8549 ( .A1(n9812), .A2(n10252), .ZN(n14339) );
  INV_X1 U8550 ( .A(n10738), .ZN(n10737) );
  NAND2_X1 U8551 ( .A1(n10696), .A2(n10737), .ZN(n10750) );
  AOI22_X1 U8552 ( .A1(n6630), .A2(n10695), .B1(n6863), .B2(n14676), .ZN(
        n10696) );
  NAND2_X1 U8553 ( .A1(n14626), .A2(n10689), .ZN(n6630) );
  AND2_X1 U8554 ( .A1(n10282), .A2(n9806), .ZN(n10272) );
  NAND2_X1 U8555 ( .A1(n7229), .A2(n6883), .ZN(n7227) );
  INV_X1 U8556 ( .A(n12360), .ZN(n6772) );
  NAND2_X1 U8557 ( .A1(n7334), .A2(n7338), .ZN(n13926) );
  NAND2_X1 U8558 ( .A1(n8529), .A2(n8528), .ZN(n11616) );
  AND2_X1 U8559 ( .A1(n10276), .A2(n10275), .ZN(n14740) );
  NAND2_X1 U8560 ( .A1(n7327), .A2(n10755), .ZN(n10864) );
  NAND2_X1 U8561 ( .A1(n10955), .A2(n10753), .ZN(n7327) );
  INV_X1 U8562 ( .A(n8301), .ZN(n7273) );
  OAI21_X1 U8563 ( .B1(n8144), .B2(n7672), .A(n7673), .ZN(n8157) );
  XNOR2_X1 U8564 ( .A(n8116), .B(n8115), .ZN(n11858) );
  NAND2_X1 U8565 ( .A1(n8103), .A2(n7665), .ZN(n8114) );
  NAND2_X1 U8566 ( .A1(n8069), .A2(n7086), .ZN(n8085) );
  NAND2_X1 U8567 ( .A1(n8085), .A2(n7662), .ZN(n8086) );
  AND2_X1 U8568 ( .A1(n8324), .A2(n8323), .ZN(n10242) );
  MUX2_X1 U8569 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8321), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n8324) );
  NAND2_X1 U8570 ( .A1(n8325), .A2(n8319), .ZN(n8327) );
  INV_X1 U8571 ( .A(n8002), .ZN(n7650) );
  OR2_X1 U8572 ( .A1(n7959), .A2(n7960), .ZN(n7378) );
  NAND2_X1 U8573 ( .A1(n7366), .A2(n7611), .ZN(n7856) );
  NAND2_X1 U8574 ( .A1(n7837), .A2(n7609), .ZN(n7366) );
  AOI21_X1 U8575 ( .B1(n7600), .B2(n7354), .A(n6465), .ZN(n7351) );
  XNOR2_X1 U8576 ( .A(n7779), .B(n7352), .ZN(n9861) );
  NAND2_X1 U8577 ( .A1(n7599), .A2(n7598), .ZN(n7779) );
  INV_X1 U8578 ( .A(n7747), .ZN(n7749) );
  INV_X1 U8579 ( .A(n7583), .ZN(n7727) );
  INV_X1 U8580 ( .A(n14211), .ZN(n14260) );
  AOI21_X1 U8581 ( .B1(n14211), .B2(n14210), .A(n14209), .ZN(n14259) );
  AND2_X1 U8582 ( .A1(n15191), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n14209) );
  INV_X1 U8583 ( .A(n14261), .ZN(n14210) );
  XNOR2_X1 U8584 ( .A(n14220), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n14267) );
  NAND2_X1 U8585 ( .A1(n15321), .A2(n14273), .ZN(n14278) );
  NOR2_X1 U8586 ( .A1(n14223), .A2(n14222), .ZN(n14276) );
  NOR2_X1 U8587 ( .A1(n14256), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n14222) );
  NAND2_X1 U8588 ( .A1(n14327), .A2(n14287), .ZN(n14290) );
  OAI22_X1 U8589 ( .A1(n14248), .A2(P1_ADDR_REG_13__SCAN_IN), .B1(n14249), 
        .B2(n14237), .ZN(n14246) );
  AND4_X1 U8590 ( .A1(n9103), .A2(n9102), .A3(n9101), .A4(n9100), .ZN(n11102)
         );
  NAND2_X1 U8591 ( .A1(n12525), .A2(n12190), .ZN(n12433) );
  INV_X1 U8592 ( .A(n7282), .ZN(n7281) );
  NAND2_X1 U8593 ( .A1(n12484), .A2(n7283), .ZN(n12441) );
  NAND2_X1 U8594 ( .A1(n9318), .A2(n9317), .ZN(n12446) );
  AOI21_X1 U8595 ( .B1(n6675), .B2(n6678), .A(n6530), .ZN(n6673) );
  INV_X1 U8596 ( .A(n12162), .ZN(n6678) );
  INV_X1 U8597 ( .A(n7291), .ZN(n7287) );
  AND3_X1 U8598 ( .A1(n9301), .A2(n9300), .A3(n9299), .ZN(n12782) );
  NAND2_X1 U8599 ( .A1(n7298), .A2(n12171), .ZN(n12458) );
  NAND2_X1 U8600 ( .A1(n7300), .A2(n7301), .ZN(n11542) );
  INV_X1 U8601 ( .A(n7302), .ZN(n7301) );
  OR2_X1 U8602 ( .A1(n11368), .A2(n11388), .ZN(n7300) );
  OAI21_X1 U8603 ( .B1(n12160), .B2(n12159), .A(n12158), .ZN(n12478) );
  OR2_X1 U8604 ( .A1(n12157), .A2(n12812), .ZN(n12158) );
  AND2_X1 U8605 ( .A1(n8969), .A2(n8968), .ZN(n12719) );
  NAND2_X1 U8606 ( .A1(n9038), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8965) );
  NAND2_X1 U8607 ( .A1(n10589), .A2(n6498), .ZN(n10593) );
  INV_X1 U8608 ( .A(n7305), .ZN(n10807) );
  NAND2_X1 U8609 ( .A1(n7307), .A2(n7309), .ZN(n11067) );
  INV_X1 U8610 ( .A(n7310), .ZN(n7309) );
  NAND2_X1 U8611 ( .A1(n10386), .A2(n10385), .ZN(n12505) );
  NAND2_X1 U8612 ( .A1(n9295), .A2(n9294), .ZN(n12774) );
  AND2_X1 U8613 ( .A1(n6669), .A2(n6575), .ZN(n11640) );
  NAND2_X1 U8614 ( .A1(n9305), .A2(n9304), .ZN(n12510) );
  AND2_X1 U8615 ( .A1(n11368), .A2(n11343), .ZN(n11389) );
  NAND2_X1 U8616 ( .A1(n10501), .A2(n10502), .ZN(n10519) );
  XNOR2_X1 U8617 ( .A(n10517), .B(n12557), .ZN(n10502) );
  NAND2_X1 U8618 ( .A1(n6674), .A2(n12162), .ZN(n12514) );
  NAND2_X1 U8619 ( .A1(n12478), .A2(n12161), .ZN(n6674) );
  INV_X1 U8620 ( .A(n12523), .ZN(n12528) );
  INV_X1 U8621 ( .A(n12516), .ZN(n12535) );
  NAND2_X1 U8622 ( .A1(n10493), .A2(n10492), .ZN(n12508) );
  NAND2_X1 U8623 ( .A1(n10374), .A2(n10373), .ZN(n12523) );
  AND2_X1 U8624 ( .A1(n9478), .A2(n9372), .ZN(n12196) );
  NAND2_X1 U8625 ( .A1(n9335), .A2(n9334), .ZN(n12734) );
  INV_X1 U8626 ( .A(n12782), .ZN(n12757) );
  INV_X1 U8627 ( .A(n12829), .ZN(n12545) );
  NAND2_X1 U8628 ( .A1(n9038), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n9134) );
  INV_X1 U8629 ( .A(n15046), .ZN(n12552) );
  INV_X1 U8630 ( .A(n11102), .ZN(n12553) );
  OR2_X2 U8631 ( .A1(n12941), .A2(n10377), .ZN(n12559) );
  NAND2_X1 U8632 ( .A1(n7167), .A2(n6455), .ZN(n10442) );
  AND2_X1 U8633 ( .A1(n7167), .A2(n10441), .ZN(n10418) );
  OR2_X1 U8634 ( .A1(n9061), .A2(n9225), .ZN(n9062) );
  AND2_X1 U8635 ( .A1(n7026), .A2(n7025), .ZN(n14901) );
  NAND2_X1 U8636 ( .A1(n10447), .A2(n6854), .ZN(n6872) );
  INV_X1 U8637 ( .A(n6690), .ZN(n10447) );
  INV_X1 U8638 ( .A(n7169), .ZN(n10532) );
  INV_X1 U8639 ( .A(n6870), .ZN(n10538) );
  XNOR2_X1 U8640 ( .A(n6847), .B(n14940), .ZN(n14933) );
  INV_X1 U8641 ( .A(n7174), .ZN(n14958) );
  NOR2_X1 U8642 ( .A1(n7016), .A2(n7015), .ZN(n14981) );
  INV_X1 U8643 ( .A(n14978), .ZN(n7016) );
  INV_X1 U8644 ( .A(n7172), .ZN(n12584) );
  INV_X1 U8645 ( .A(n7163), .ZN(n14985) );
  OAI21_X1 U8646 ( .B1(n12606), .B2(n7009), .A(n7007), .ZN(n15000) );
  AOI21_X1 U8647 ( .B1(n7011), .B2(n7010), .A(n7008), .ZN(n7007) );
  INV_X1 U8648 ( .A(n15001), .ZN(n7008) );
  INV_X1 U8649 ( .A(n7006), .ZN(n15002) );
  AOI21_X1 U8650 ( .B1(n12606), .B2(n7013), .A(n7009), .ZN(n7006) );
  INV_X1 U8651 ( .A(n7161), .ZN(n12587) );
  NOR2_X1 U8652 ( .A1(n15015), .A2(n6989), .ZN(n15040) );
  AND2_X1 U8653 ( .A1(n12612), .A2(n12613), .ZN(n6989) );
  NAND2_X1 U8654 ( .A1(n15040), .A2(n15039), .ZN(n15038) );
  INV_X1 U8655 ( .A(n7171), .ZN(n14387) );
  NOR2_X1 U8656 ( .A1(n14379), .A2(n7005), .ZN(n14399) );
  XNOR2_X1 U8657 ( .A(n6871), .B(n14413), .ZN(n14404) );
  AND2_X1 U8658 ( .A1(n6452), .A2(n7002), .ZN(n14409) );
  NAND2_X1 U8659 ( .A1(n7002), .A2(n7003), .ZN(n14410) );
  NAND2_X1 U8660 ( .A1(n12634), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7165) );
  AND2_X1 U8661 ( .A1(n7128), .A2(n9629), .ZN(n12678) );
  NAND2_X1 U8662 ( .A1(n7489), .A2(n7490), .ZN(n12672) );
  NOR2_X1 U8663 ( .A1(n9327), .A2(n9060), .ZN(n12851) );
  NAND2_X1 U8664 ( .A1(n12780), .A2(n9291), .ZN(n12767) );
  NAND2_X1 U8665 ( .A1(n6933), .A2(n7121), .ZN(n12802) );
  NAND2_X1 U8666 ( .A1(n9405), .A2(n9586), .ZN(n12818) );
  NAND2_X1 U8667 ( .A1(n12830), .A2(n12831), .ZN(n9405) );
  AND2_X1 U8668 ( .A1(n12816), .A2(n12815), .ZN(n12882) );
  NAND2_X1 U8669 ( .A1(n11649), .A2(n9238), .ZN(n11749) );
  NAND2_X1 U8670 ( .A1(n6922), .A2(n6925), .ZN(n11648) );
  OR2_X1 U8671 ( .A1(n14442), .A2(n6927), .ZN(n6922) );
  AND2_X1 U8672 ( .A1(n11671), .A2(n9222), .ZN(n11651) );
  NAND2_X1 U8673 ( .A1(n6930), .A2(n9572), .ZN(n11669) );
  NAND2_X1 U8674 ( .A1(n14442), .A2(n14441), .ZN(n6930) );
  NAND2_X1 U8675 ( .A1(n11434), .A2(n9191), .ZN(n7474) );
  NAND2_X1 U8676 ( .A1(n10891), .A2(n9097), .ZN(n15050) );
  OR2_X1 U8677 ( .A1(n10396), .A2(n10390), .ZN(n15081) );
  INV_X1 U8678 ( .A(n12805), .ZN(n14445) );
  INV_X1 U8679 ( .A(n12446), .ZN(n12907) );
  INV_X1 U8680 ( .A(n12510), .ZN(n12911) );
  NAND2_X1 U8681 ( .A1(n9263), .A2(n9262), .ZN(n12925) );
  NAND2_X1 U8682 ( .A1(n8995), .A2(n8994), .ZN(n12929) );
  AOI22_X1 U8683 ( .A1(n6432), .A2(SI_11_), .B1(n9060), .B2(n12643), .ZN(n9189) );
  NAND2_X1 U8684 ( .A1(n10397), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12941) );
  AOI22_X1 U8685 ( .A1(n9481), .A2(n9480), .B1(P1_DATAO_REG_30__SCAN_IN), .B2(
        n12153), .ZN(n9483) );
  XNOR2_X1 U8686 ( .A(n9481), .B(n7268), .ZN(n12949) );
  INV_X1 U8687 ( .A(n9471), .ZN(n7268) );
  NAND2_X1 U8688 ( .A1(n8908), .A2(n8907), .ZN(n12952) );
  NOR2_X1 U8689 ( .A1(n8905), .A2(n8904), .ZN(n8908) );
  NAND2_X1 U8690 ( .A1(n8906), .A2(n6819), .ZN(n8907) );
  NOR2_X1 U8691 ( .A1(P3_IR_REG_29__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8904) );
  INV_X1 U8692 ( .A(n7269), .ZN(n9364) );
  INV_X1 U8693 ( .A(SI_26_), .ZN(n12961) );
  INV_X1 U8694 ( .A(n6833), .ZN(n9337) );
  XNOR2_X1 U8695 ( .A(n9378), .B(P3_IR_REG_22__SCAN_IN), .ZN(n10962) );
  NAND2_X1 U8696 ( .A1(n9413), .A2(n9381), .ZN(n10714) );
  MUX2_X1 U8697 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9380), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n9381) );
  NAND2_X1 U8698 ( .A1(n7251), .A2(n7249), .ZN(n8977) );
  INV_X1 U8699 ( .A(SI_20_), .ZN(n10583) );
  XNOR2_X1 U8700 ( .A(n9383), .B(n9382), .ZN(n10585) );
  NAND2_X1 U8701 ( .A1(n6479), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9383) );
  INV_X1 U8702 ( .A(n6947), .ZN(n6945) );
  INV_X1 U8703 ( .A(SI_16_), .ZN(n10139) );
  INV_X1 U8704 ( .A(n12650), .ZN(n14393) );
  NAND2_X1 U8705 ( .A1(n8987), .A2(n9226), .ZN(n9241) );
  INV_X1 U8706 ( .A(SI_15_), .ZN(n10040) );
  NAND2_X1 U8707 ( .A1(n7247), .A2(n8940), .ZN(n9240) );
  NAND2_X1 U8708 ( .A1(n9224), .A2(n9223), .ZN(n7247) );
  OR2_X1 U8709 ( .A1(n8987), .A2(n9225), .ZN(n9227) );
  INV_X1 U8710 ( .A(n12643), .ZN(n14975) );
  OAI21_X1 U8711 ( .B1(n8927), .B2(n6443), .A(n7233), .ZN(n9137) );
  NAND2_X1 U8712 ( .A1(n7236), .A2(n8929), .ZN(n9121) );
  NAND2_X1 U8713 ( .A1(n8927), .A2(n7237), .ZN(n7236) );
  NAND2_X1 U8714 ( .A1(n8927), .A2(n8926), .ZN(n9105) );
  INV_X1 U8715 ( .A(n10541), .ZN(n10548) );
  NAND2_X1 U8716 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n9032) );
  INV_X1 U8717 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n11787) );
  XNOR2_X1 U8718 ( .A(n9766), .B(n9767), .ZN(n12964) );
  NAND2_X1 U8719 ( .A1(n6698), .A2(n6696), .ZN(n11294) );
  AOI21_X1 U8720 ( .B1(n6699), .B2(n6701), .A(n6697), .ZN(n6696) );
  NAND2_X1 U8721 ( .A1(n7468), .A2(n6699), .ZN(n6698) );
  INV_X1 U8722 ( .A(n9716), .ZN(n6697) );
  NAND2_X1 U8723 ( .A1(n7468), .A2(n9703), .ZN(n11130) );
  OAI21_X1 U8724 ( .B1(n7468), .B2(n6701), .A(n6699), .ZN(n11200) );
  NAND2_X1 U8725 ( .A1(n11127), .A2(n9710), .ZN(n11201) );
  NAND2_X1 U8726 ( .A1(n6707), .A2(n7443), .ZN(n6704) );
  NAND2_X1 U8727 ( .A1(n11572), .A2(n9728), .ZN(n11660) );
  INV_X1 U8728 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n13106) );
  NAND2_X1 U8729 ( .A1(n9795), .A2(n9794), .ZN(n13108) );
  AND2_X1 U8730 ( .A1(n10031), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13110) );
  OR2_X1 U8731 ( .A1(n15339), .A2(n7711), .ZN(n7695) );
  OR2_X1 U8732 ( .A1(n6827), .A2(n10774), .ZN(n7776) );
  OR2_X1 U8733 ( .A1(n7965), .A2(n7738), .ZN(n7556) );
  OR2_X1 U8734 ( .A1(n7754), .A2(n10632), .ZN(n7732) );
  OR2_X1 U8735 ( .A1(n8079), .A2(n7729), .ZN(n7733) );
  INV_X1 U8736 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13254) );
  AND2_X1 U8737 ( .A1(n9902), .A2(n12145), .ZN(n14820) );
  NAND2_X1 U8738 ( .A1(n13265), .A2(n6800), .ZN(n6799) );
  INV_X1 U8739 ( .A(n6838), .ZN(n6798) );
  NAND2_X1 U8740 ( .A1(n6781), .A2(n6811), .ZN(n13311) );
  AOI21_X1 U8741 ( .B1(n13340), .B2(n8101), .A(n6466), .ZN(n13324) );
  NAND2_X1 U8742 ( .A1(n13355), .A2(n8252), .ZN(n13345) );
  NAND2_X1 U8743 ( .A1(n6803), .A2(n6804), .ZN(n13379) );
  NAND2_X1 U8744 ( .A1(n8038), .A2(n8037), .ZN(n13393) );
  NAND2_X1 U8745 ( .A1(n13435), .A2(n8247), .ZN(n13423) );
  NAND2_X1 U8746 ( .A1(n13429), .A2(n8000), .ZN(n13412) );
  NAND2_X1 U8747 ( .A1(n11767), .A2(n7973), .ZN(n13451) );
  NAND2_X1 U8748 ( .A1(n7958), .A2(n7957), .ZN(n11769) );
  NAND2_X1 U8749 ( .A1(n7210), .A2(n8236), .ZN(n11443) );
  NAND2_X1 U8750 ( .A1(n11278), .A2(n12117), .ZN(n7210) );
  NAND2_X1 U8751 ( .A1(n7182), .A2(n7835), .ZN(n10986) );
  INV_X1 U8752 ( .A(n14837), .ZN(n11883) );
  NAND2_X1 U8753 ( .A1(n7879), .A2(n7878), .ZN(n11946) );
  NAND2_X1 U8754 ( .A1(n12152), .A2(n7750), .ZN(n12052) );
  INV_X1 U8755 ( .A(n6868), .ZN(n6867) );
  OAI21_X1 U8756 ( .B1(n13492), .B2(n11860), .A(n13490), .ZN(n6868) );
  NAND2_X1 U8757 ( .A1(n7204), .A2(n8257), .ZN(n13298) );
  NAND2_X1 U8758 ( .A1(n8255), .A2(n7205), .ZN(n7204) );
  NAND2_X1 U8759 ( .A1(n8255), .A2(n8254), .ZN(n13310) );
  INV_X1 U8760 ( .A(n11968), .ZN(n11966) );
  INV_X1 U8761 ( .A(n13602), .ZN(n13616) );
  AND2_X1 U8762 ( .A1(n9807), .A2(n8218), .ZN(n14835) );
  INV_X1 U8763 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13623) );
  AND2_X1 U8764 ( .A1(n7470), .A2(n7190), .ZN(n7189) );
  INV_X1 U8765 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7190) );
  INV_X1 U8766 ( .A(n7426), .ZN(n13634) );
  NAND2_X1 U8767 ( .A1(n8199), .A2(n8202), .ZN(n13644) );
  XNOR2_X1 U8768 ( .A(n8192), .B(n8191), .ZN(n13652) );
  INV_X1 U8769 ( .A(n8221), .ZN(n13249) );
  INV_X1 U8770 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10587) );
  INV_X1 U8771 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10576) );
  INV_X1 U8772 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10424) );
  INV_X1 U8773 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10259) );
  INV_X1 U8774 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9963) );
  INV_X1 U8775 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n15289) );
  INV_X1 U8776 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9925) );
  INV_X1 U8777 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n15276) );
  INV_X1 U8778 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9881) );
  INV_X1 U8779 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9876) );
  INV_X1 U8780 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9868) );
  XNOR2_X1 U8781 ( .A(n7723), .B(n7722), .ZN(n9938) );
  INV_X1 U8782 ( .A(n9806), .ZN(n10323) );
  AOI21_X1 U8783 ( .B1(n11189), .B2(n11188), .A(n6448), .ZN(n11404) );
  NAND2_X1 U8784 ( .A1(n6649), .A2(n6816), .ZN(n14566) );
  NAND2_X1 U8785 ( .A1(n6651), .A2(n6650), .ZN(n6649) );
  INV_X1 U8786 ( .A(n12381), .ZN(n14136) );
  AND4_X1 U8787 ( .A1(n8473), .A2(n8472), .A3(n8471), .A4(n8470), .ZN(n11553)
         );
  NAND2_X1 U8788 ( .A1(n7523), .A2(n7524), .ZN(n11413) );
  AND2_X1 U8789 ( .A1(n10736), .A2(n10673), .ZN(n14584) );
  NAND2_X1 U8790 ( .A1(n7537), .A2(n12266), .ZN(n13687) );
  NOR2_X1 U8791 ( .A1(n14508), .A2(n7554), .ZN(n11846) );
  NAND2_X1 U8792 ( .A1(n7532), .A2(n7533), .ZN(n12205) );
  NAND2_X1 U8793 ( .A1(n12230), .A2(n13786), .ZN(n13707) );
  AND4_X1 U8794 ( .A1(n8716), .A2(n8715), .A3(n8714), .A4(n8713), .ZN(n13779)
         );
  AND4_X1 U8795 ( .A1(n8492), .A2(n8491), .A3(n8490), .A4(n8489), .ZN(n11828)
         );
  NAND2_X1 U8796 ( .A1(n8343), .A2(n14208), .ZN(n6760) );
  OR2_X1 U8797 ( .A1(n8343), .A2(n6762), .ZN(n6761) );
  AOI21_X1 U8798 ( .B1(n7533), .B2(n7530), .A(n6491), .ZN(n7529) );
  INV_X1 U8799 ( .A(n7533), .ZN(n7531) );
  NAND2_X1 U8800 ( .A1(n10937), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14572) );
  NAND2_X1 U8801 ( .A1(n13697), .A2(n12311), .ZN(n13776) );
  NAND2_X1 U8802 ( .A1(n13776), .A2(n13777), .ZN(n13775) );
  AND4_X1 U8803 ( .A1(n8588), .A2(n8587), .A3(n8586), .A4(n8585), .ZN(n13792)
         );
  XNOR2_X1 U8804 ( .A(n12227), .B(n12228), .ZN(n13788) );
  AND2_X1 U8805 ( .A1(n8853), .A2(n8854), .ZN(n7071) );
  NAND2_X1 U8806 ( .A1(n8860), .A2(n8859), .ZN(n8861) );
  NAND2_X1 U8807 ( .A1(n7074), .A2(n7073), .ZN(n7072) );
  INV_X1 U8808 ( .A(n8824), .ZN(n14052) );
  INV_X1 U8809 ( .A(n8827), .ZN(n8828) );
  CLKBUF_X1 U8810 ( .A(n10357), .Z(n6863) );
  CLKBUF_X2 U8811 ( .A(P1_U4016), .Z(n13812) );
  AND2_X1 U8812 ( .A1(n8332), .A2(n8334), .ZN(n6756) );
  INV_X1 U8813 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n15191) );
  NAND2_X1 U8814 ( .A1(n13817), .A2(n6864), .ZN(n13830) );
  OR2_X1 U8815 ( .A1(n13814), .A2(n10008), .ZN(n6864) );
  NAND2_X1 U8816 ( .A1(n13830), .A2(n13831), .ZN(n13829) );
  INV_X1 U8817 ( .A(n8850), .ZN(n14069) );
  INV_X1 U8818 ( .A(n13900), .ZN(n14072) );
  XNOR2_X1 U8819 ( .A(n6623), .B(n12380), .ZN(n14077) );
  OAI21_X1 U8820 ( .B1(n12399), .B2(n6622), .A(n6535), .ZN(n6623) );
  INV_X1 U8821 ( .A(n6882), .ZN(n6622) );
  INV_X1 U8822 ( .A(n6915), .ZN(n14080) );
  OAI21_X1 U8823 ( .B1(n14090), .B2(n14631), .A(n12404), .ZN(n12405) );
  NAND2_X1 U8824 ( .A1(n7331), .A2(n12371), .ZN(n13987) );
  NAND2_X1 U8825 ( .A1(n12349), .A2(n12348), .ZN(n14034) );
  NAND2_X1 U8826 ( .A1(n11807), .A2(n11806), .ZN(n12346) );
  INV_X1 U8827 ( .A(n7322), .ZN(n11624) );
  AOI21_X1 U8828 ( .B1(n14350), .B2(n14349), .A(n6464), .ZN(n7322) );
  NAND2_X1 U8829 ( .A1(n14346), .A2(n11590), .ZN(n11628) );
  CLKBUF_X1 U8830 ( .A(n10243), .Z(n14345) );
  OAI21_X1 U8831 ( .B1(n11154), .B2(n7255), .A(n7253), .ZN(n11475) );
  NAND2_X1 U8832 ( .A1(n11330), .A2(n11329), .ZN(n11331) );
  NAND2_X1 U8833 ( .A1(n7342), .A2(n10973), .ZN(n11145) );
  OR2_X1 U8834 ( .A1(n11080), .A2(n10972), .ZN(n7342) );
  NAND2_X1 U8835 ( .A1(n7275), .A2(n10745), .ZN(n10861) );
  OR2_X1 U8836 ( .A1(n12386), .A2(n14345), .ZN(n14639) );
  INV_X1 U8837 ( .A(n14636), .ZN(n14608) );
  AND2_X1 U8838 ( .A1(n10272), .A2(n10930), .ZN(n14636) );
  AND2_X1 U8839 ( .A1(n14610), .A2(n14138), .ZN(n14045) );
  AND2_X2 U8840 ( .A1(n10736), .A2(n10735), .ZN(n14748) );
  INV_X1 U8841 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6774) );
  OR2_X1 U8842 ( .A1(n14085), .A2(n14153), .ZN(n6916) );
  OR2_X1 U8843 ( .A1(n14109), .A2(n14108), .ZN(n14176) );
  AND2_X2 U8844 ( .A1(n10241), .A2(n10735), .ZN(n15160) );
  INV_X1 U8845 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8302) );
  INV_X1 U8846 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14194) );
  NAND2_X1 U8847 ( .A1(n8298), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8295) );
  INV_X1 U8848 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15193) );
  INV_X1 U8849 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14200) );
  INV_X1 U8850 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11859) );
  INV_X1 U8851 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8870) );
  NAND2_X1 U8852 ( .A1(n8879), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8871) );
  INV_X1 U8853 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n15178) );
  INV_X1 U8854 ( .A(n10242), .ZN(n11492) );
  NAND2_X1 U8855 ( .A1(n8051), .A2(n7658), .ZN(n8054) );
  INV_X1 U8856 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n12155) );
  INV_X1 U8857 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10425) );
  INV_X1 U8858 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9959) );
  INV_X1 U8859 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9926) );
  INV_X1 U8860 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9882) );
  INV_X1 U8861 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9874) );
  INV_X1 U8862 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9862) );
  XNOR2_X1 U8863 ( .A(n14272), .B(n14271), .ZN(n15323) );
  NAND2_X1 U8864 ( .A1(n15323), .A2(n15322), .ZN(n15321) );
  INV_X1 U8865 ( .A(n15327), .ZN(n7135) );
  XNOR2_X1 U8866 ( .A(n14286), .B(n14285), .ZN(n14329) );
  INV_X1 U8867 ( .A(n14284), .ZN(n14285) );
  NAND2_X1 U8868 ( .A1(n14329), .A2(n14328), .ZN(n14327) );
  XNOR2_X1 U8869 ( .A(n14290), .B(n14291), .ZN(n14331) );
  NAND2_X1 U8870 ( .A1(n14543), .A2(n14297), .ZN(n14546) );
  NAND2_X1 U8871 ( .A1(n7134), .A2(n7133), .ZN(n14556) );
  NAND2_X1 U8872 ( .A1(n14556), .A2(n14557), .ZN(n14553) );
  NAND2_X1 U8873 ( .A1(n7132), .A2(n6486), .ZN(n14555) );
  NAND2_X1 U8874 ( .A1(n14553), .A2(n14555), .ZN(n14560) );
  NAND2_X1 U8875 ( .A1(n14309), .A2(n14357), .ZN(n14364) );
  OR2_X1 U8876 ( .A1(n14359), .A2(n14358), .ZN(n14308) );
  NAND2_X1 U8877 ( .A1(n14364), .A2(n14365), .ZN(n14366) );
  OAI21_X1 U8878 ( .B1(n14364), .B2(n14365), .A(n15255), .ZN(n7142) );
  NAND2_X1 U8879 ( .A1(n6693), .A2(n14866), .ZN(n6692) );
  XNOR2_X1 U8880 ( .A(n7164), .B(n12597), .ZN(n12661) );
  NAND2_X1 U8881 ( .A1(n7166), .A2(n7165), .ZN(n7164) );
  OAI211_X1 U8882 ( .C1(n12835), .C2(n9466), .A(n12428), .B(n6478), .ZN(n12429) );
  OAI22_X1 U8883 ( .A1(n12897), .A2(n12894), .B1(n15157), .B2(n15229), .ZN(
        n9658) );
  OAI21_X1 U8884 ( .B1(n12895), .B2(n15142), .A(n7479), .ZN(P3_U3455) );
  INV_X1 U8885 ( .A(n7480), .ZN(n7479) );
  OAI22_X1 U8886 ( .A1(n12897), .A2(n12939), .B1(n15141), .B2(n12896), .ZN(
        n7480) );
  NOR2_X1 U8887 ( .A1(n9782), .A2(n9783), .ZN(n12988) );
  NAND2_X1 U8888 ( .A1(n7432), .A2(n9789), .ZN(n7431) );
  NAND2_X1 U8889 ( .A1(n10030), .A2(n9669), .ZN(n10042) );
  NAND2_X1 U8890 ( .A1(n6875), .A2(n6874), .ZN(n6873) );
  INV_X1 U8891 ( .A(n13013), .ZN(n6874) );
  NAND2_X1 U8892 ( .A1(n7456), .A2(n7457), .ZN(n10510) );
  NAND2_X1 U8893 ( .A1(n8270), .A2(n13470), .ZN(n8281) );
  INV_X1 U8894 ( .A(n8279), .ZN(n8280) );
  INV_X1 U8895 ( .A(n6843), .ZN(n6842) );
  OAI21_X1 U8896 ( .B1(n13492), .B2(n13279), .A(n13278), .ZN(n6843) );
  OAI21_X1 U8897 ( .B1(n9662), .B2(n14862), .A(n8264), .ZN(P2_U3528) );
  INV_X1 U8898 ( .A(n8263), .ZN(n8264) );
  INV_X1 U8899 ( .A(n6858), .ZN(n6857) );
  OAI21_X1 U8900 ( .B1(n13572), .B2(n13561), .A(n13496), .ZN(n6858) );
  OAI21_X1 U8901 ( .B1(n9662), .B2(n14858), .A(n9666), .ZN(P2_U3496) );
  INV_X1 U8902 ( .A(n9665), .ZN(n9666) );
  INV_X1 U8903 ( .A(n6860), .ZN(n6859) );
  NAND2_X1 U8904 ( .A1(n6802), .A2(n6801), .ZN(n13571) );
  OAI21_X1 U8905 ( .B1(n13572), .B2(n13620), .A(n13570), .ZN(n6860) );
  NOR2_X1 U8906 ( .A1(n6836), .A2(n6835), .ZN(n6834) );
  INV_X1 U8907 ( .A(n13663), .ZN(n6835) );
  INV_X1 U8908 ( .A(n6651), .ZN(n10921) );
  MUX2_X1 U8909 ( .A(n13890), .B(n13889), .S(n8883), .Z(n13892) );
  NAND2_X1 U8910 ( .A1(n15160), .A2(n14729), .ZN(n6770) );
  NAND2_X1 U8911 ( .A1(n6769), .A2(n15160), .ZN(n6768) );
  NAND2_X1 U8912 ( .A1(n6913), .A2(n6912), .ZN(P1_U3524) );
  OR2_X1 U8913 ( .A1(n15160), .A2(n15286), .ZN(n6912) );
  NAND2_X1 U8914 ( .A1(n14172), .A2(n15160), .ZN(n6913) );
  NOR2_X1 U8915 ( .A1(n14333), .A2(n14334), .ZN(n14332) );
  OAI21_X1 U8916 ( .B1(n14333), .B2(n7154), .A(n7152), .ZN(n14539) );
  NAND2_X1 U8917 ( .A1(n7156), .A2(n7157), .ZN(n14540) );
  XNOR2_X1 U8918 ( .A(n7141), .B(n7140), .ZN(SUB_1596_U4) );
  XNOR2_X1 U8919 ( .A(n14368), .B(n14367), .ZN(n7140) );
  NAND2_X1 U8920 ( .A1(n7142), .A2(n14366), .ZN(n7141) );
  XNOR2_X1 U8921 ( .A(n7552), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n14367) );
  INV_X1 U8922 ( .A(n14082), .ZN(n6883) );
  AND2_X1 U8923 ( .A1(n7375), .A2(SI_17_), .ZN(n6441) );
  AND2_X1 U8924 ( .A1(n7667), .A2(n7082), .ZN(n6442) );
  INV_X2 U8925 ( .A(n11863), .ZN(n12059) );
  NAND2_X4 U8926 ( .A1(n6744), .A2(n6742), .ZN(n11863) );
  INV_X1 U8927 ( .A(n14922), .ZN(n6854) );
  INV_X1 U8928 ( .A(n7157), .ZN(n7154) );
  NAND2_X1 U8929 ( .A1(n13103), .A2(n6509), .ZN(n7449) );
  OR2_X1 U8930 ( .A1(n9120), .A2(n7235), .ZN(n6443) );
  NOR2_X1 U8931 ( .A1(n7302), .A2(n11541), .ZN(n6444) );
  OR2_X1 U8932 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10407), .ZN(n6445) );
  AND2_X1 U8933 ( .A1(n12041), .A2(n7406), .ZN(n6446) );
  INV_X1 U8934 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7678) );
  AND2_X1 U8935 ( .A1(n7757), .A2(n6508), .ZN(n6447) );
  AND2_X1 U8936 ( .A1(n11187), .A2(n11186), .ZN(n6448) );
  NAND2_X1 U8937 ( .A1(n8343), .A2(n9831), .ZN(n8408) );
  INV_X1 U8938 ( .A(n8408), .ZN(n6825) );
  AND2_X1 U8939 ( .A1(n6545), .A2(n7050), .ZN(n6449) );
  OR2_X1 U8940 ( .A1(n14717), .A2(n11408), .ZN(n6450) );
  OR2_X1 U8941 ( .A1(n6975), .A2(n9633), .ZN(n6451) );
  INV_X1 U8942 ( .A(n13431), .ZN(n13436) );
  AND2_X1 U8943 ( .A1(n7003), .A2(n12626), .ZN(n6452) );
  INV_X1 U8944 ( .A(n6743), .ZN(n11860) );
  AND2_X1 U8945 ( .A1(n7266), .A2(n12348), .ZN(n6453) );
  AND2_X1 U8946 ( .A1(n6443), .A2(n6469), .ZN(n6454) );
  AND2_X1 U8947 ( .A1(n10441), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n6455) );
  INV_X1 U8948 ( .A(n12810), .ZN(n12817) );
  INV_X1 U8949 ( .A(n14087), .ZN(n13664) );
  AND2_X1 U8950 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n6456) );
  INV_X1 U8951 ( .A(n11863), .ZN(n12066) );
  AND2_X1 U8952 ( .A1(n6971), .A2(n6970), .ZN(n6457) );
  AND2_X1 U8953 ( .A1(n12356), .A2(n12355), .ZN(n6458) );
  AND2_X1 U8954 ( .A1(n6594), .A2(n12236), .ZN(n6459) );
  OR2_X1 U8955 ( .A1(n12222), .A2(n12226), .ZN(n11721) );
  AND2_X1 U8956 ( .A1(n7433), .A2(n6482), .ZN(n6460) );
  AND2_X1 U8957 ( .A1(n9594), .A2(n9598), .ZN(n6461) );
  AND2_X1 U8958 ( .A1(n7647), .A2(n6561), .ZN(n6462) );
  AND2_X1 U8959 ( .A1(n6741), .A2(n12026), .ZN(n6463) );
  AND2_X1 U8960 ( .A1(n7690), .A2(n7689), .ZN(n12060) );
  INV_X1 U8961 ( .A(n12060), .ZN(n12058) );
  NAND2_X1 U8962 ( .A1(n7565), .A2(n7379), .ZN(n7374) );
  AOI21_X1 U8963 ( .B1(n6444), .B2(n11388), .A(n6550), .ZN(n7299) );
  NAND2_X1 U8964 ( .A1(n6612), .A2(n9506), .ZN(n11671) );
  INV_X1 U8965 ( .A(n12703), .ZN(n7491) );
  INV_X1 U8966 ( .A(n14004), .ZN(n6899) );
  AND3_X1 U8967 ( .A1(n8983), .A2(n8982), .A3(n8981), .ZN(n12769) );
  INV_X1 U8968 ( .A(SI_17_), .ZN(n6898) );
  INV_X1 U8969 ( .A(n9239), .ZN(n7246) );
  NAND2_X2 U8970 ( .A1(n7978), .A2(n7977), .ZN(n13551) );
  INV_X1 U8971 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9878) );
  NAND2_X1 U8972 ( .A1(n15339), .A2(n7189), .ZN(n7191) );
  NOR2_X1 U8973 ( .A1(n14343), .A2(n12206), .ZN(n6464) );
  AND2_X1 U8974 ( .A1(n7601), .A2(SI_5_), .ZN(n6465) );
  XNOR2_X1 U8975 ( .A(n7709), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8221) );
  AND2_X1 U8976 ( .A1(n13587), .A2(n13040), .ZN(n6466) );
  NAND2_X1 U8977 ( .A1(n7320), .A2(n7319), .ZN(n8456) );
  NAND2_X1 U8978 ( .A1(n7442), .A2(n13023), .ZN(n12972) );
  NAND2_X1 U8979 ( .A1(n7679), .A2(n7678), .ZN(n7768) );
  NAND4_X1 U8980 ( .A1(n9029), .A2(n9028), .A3(n9027), .A4(n9026), .ZN(n12558)
         );
  AND2_X1 U8981 ( .A1(n7281), .A2(n12484), .ZN(n6467) );
  AND2_X1 U8982 ( .A1(n7537), .A2(n7535), .ZN(n6468) );
  INV_X1 U8983 ( .A(n9051), .ZN(n9129) );
  NAND2_X1 U8984 ( .A1(n9882), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n6469) );
  NOR2_X1 U8985 ( .A1(n10263), .A2(n7460), .ZN(n6470) );
  NAND2_X1 U8986 ( .A1(n8609), .A2(n7544), .ZN(n6471) );
  OR2_X1 U8987 ( .A1(n10362), .A2(n10361), .ZN(n6472) );
  AND3_X1 U8988 ( .A1(n8371), .A2(n8370), .A3(n8372), .ZN(n6473) );
  XOR2_X1 U8989 ( .A(n13257), .B(n12422), .Z(n6474) );
  AND2_X1 U8990 ( .A1(n9571), .A2(n10398), .ZN(n6475) );
  OR2_X1 U8991 ( .A1(n8237), .A2(n7209), .ZN(n6476) );
  INV_X1 U8992 ( .A(n12040), .ZN(n7406) );
  INV_X1 U8993 ( .A(n7521), .ZN(n7520) );
  NAND2_X1 U8994 ( .A1(n7524), .A2(n7522), .ZN(n7521) );
  OR2_X1 U8995 ( .A1(n10533), .A2(n10534), .ZN(n6477) );
  OR2_X1 U8996 ( .A1(n12427), .A2(n12805), .ZN(n6478) );
  INV_X1 U8997 ( .A(n7600), .ZN(n7352) );
  NAND2_X1 U8998 ( .A1(n9278), .A2(n6945), .ZN(n6479) );
  NAND2_X1 U8999 ( .A1(n9583), .A2(n9580), .ZN(n11748) );
  OR2_X1 U9000 ( .A1(n12695), .A2(n12703), .ZN(n9629) );
  AND2_X1 U9001 ( .A1(n9226), .A2(n7317), .ZN(n6480) );
  INV_X1 U9002 ( .A(n10951), .ZN(n10949) );
  AND2_X1 U9003 ( .A1(n8393), .A2(n8392), .ZN(n10951) );
  AND2_X1 U9004 ( .A1(n12679), .A2(n9629), .ZN(n6481) );
  NAND2_X1 U9005 ( .A1(n7633), .A2(n7632), .ZN(n7959) );
  NAND2_X1 U9006 ( .A1(n8004), .A2(n7652), .ZN(n8021) );
  OR2_X1 U9007 ( .A1(n12992), .A2(n12987), .ZN(n6482) );
  OR2_X1 U9008 ( .A1(n7033), .A2(n8449), .ZN(n6483) );
  AND2_X1 U9009 ( .A1(n12550), .A2(n11181), .ZN(n6484) );
  AND4_X1 U9010 ( .A1(n9019), .A2(n9018), .A3(n9017), .A4(n9016), .ZN(n10516)
         );
  AND2_X1 U9011 ( .A1(n7763), .A2(n7764), .ZN(n11889) );
  INV_X1 U9012 ( .A(n15077), .ZN(n10504) );
  AND3_X1 U9013 ( .A1(n9025), .A2(n9024), .A3(n9023), .ZN(n15077) );
  INV_X1 U9014 ( .A(n13376), .ZN(n13526) );
  AND2_X1 U9015 ( .A1(n11019), .A2(n11017), .ZN(n6485) );
  XOR2_X1 U9016 ( .A(n14302), .B(n14301), .Z(n6486) );
  INV_X1 U9017 ( .A(n11591), .ZN(n11627) );
  INV_X1 U9018 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7240) );
  NAND2_X1 U9020 ( .A1(n7426), .A2(n13629), .ZN(n7951) );
  XNOR2_X1 U9021 ( .A(n8903), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8909) );
  INV_X1 U9022 ( .A(n13921), .ZN(n6903) );
  OR2_X1 U9023 ( .A1(n7406), .A2(n12041), .ZN(n6487) );
  XNOR2_X1 U9024 ( .A(n9417), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9424) );
  INV_X1 U9025 ( .A(n9424), .ZN(n6679) );
  INV_X1 U9026 ( .A(n12274), .ZN(n12312) );
  AND2_X1 U9027 ( .A1(n8146), .A2(n8145), .ZN(n13286) );
  INV_X1 U9028 ( .A(n13286), .ZN(n13569) );
  OR3_X1 U9029 ( .A1(n11992), .A2(n11991), .A3(n11990), .ZN(n6488) );
  INV_X1 U9030 ( .A(n8749), .ZN(n7380) );
  INV_X1 U9031 ( .A(n8688), .ZN(n7062) );
  INV_X1 U9032 ( .A(n8777), .ZN(n7372) );
  INV_X1 U9033 ( .A(n8418), .ZN(n7056) );
  INV_X1 U9034 ( .A(n8483), .ZN(n7059) );
  NAND2_X1 U9035 ( .A1(n9632), .A2(n9396), .ZN(n12194) );
  INV_X1 U9036 ( .A(n12194), .ZN(n6938) );
  OR2_X1 U9037 ( .A1(n14456), .A2(n11751), .ZN(n9581) );
  INV_X1 U9038 ( .A(n9581), .ZN(n6974) );
  AND2_X1 U9039 ( .A1(n13046), .A2(n7443), .ZN(n6489) );
  INV_X1 U9040 ( .A(n13940), .ZN(n14100) );
  INV_X1 U9041 ( .A(n13657), .ZN(n7516) );
  OR2_X1 U9042 ( .A1(n14281), .A2(n14280), .ZN(n6490) );
  NAND3_X1 U9043 ( .A1(n8362), .A2(n8363), .A3(n6824), .ZN(n10694) );
  INV_X1 U9044 ( .A(n10694), .ZN(n7038) );
  AND2_X1 U9045 ( .A1(n12203), .A2(n12204), .ZN(n6491) );
  INV_X1 U9046 ( .A(n13024), .ZN(n7448) );
  INV_X1 U9047 ( .A(n9402), .ZN(n14441) );
  INV_X1 U9048 ( .A(n11019), .ZN(n6908) );
  AND2_X1 U9049 ( .A1(n12372), .A2(n12371), .ZN(n6492) );
  AND4_X1 U9050 ( .A1(n9183), .A2(n9182), .A3(n9181), .A4(n9180), .ZN(n11394)
         );
  INV_X1 U9051 ( .A(n11394), .ZN(n14436) );
  AND2_X1 U9052 ( .A1(n10973), .A2(n6450), .ZN(n6493) );
  AND2_X1 U9053 ( .A1(n9834), .A2(n9835), .ZN(n6494) );
  AND2_X1 U9054 ( .A1(n12220), .A2(n12221), .ZN(n6495) );
  AND2_X1 U9055 ( .A1(n11881), .A2(n11880), .ZN(n6496) );
  AND2_X1 U9056 ( .A1(n8915), .A2(n8914), .ZN(n12703) );
  AND2_X1 U9057 ( .A1(n10862), .A2(n10753), .ZN(n6497) );
  INV_X1 U9058 ( .A(n6959), .ZN(n6958) );
  OAI21_X1 U9059 ( .B1(n6523), .B2(n6960), .A(n6961), .ZN(n6959) );
  INV_X1 U9060 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7580) );
  OR2_X1 U9061 ( .A1(n10590), .A2(n15086), .ZN(n6498) );
  NAND2_X1 U9062 ( .A1(n13422), .A2(n12981), .ZN(n6499) );
  NOR2_X1 U9063 ( .A1(n11953), .A2(n13133), .ZN(n6500) );
  AND2_X1 U9064 ( .A1(n7387), .A2(n7394), .ZN(n6501) );
  INV_X1 U9065 ( .A(n7339), .ZN(n7338) );
  NAND2_X1 U9066 ( .A1(n13928), .A2(n7340), .ZN(n7339) );
  INV_X1 U9067 ( .A(n11914), .ZN(n7420) );
  AND2_X1 U9068 ( .A1(n9585), .A2(n9586), .ZN(n12831) );
  INV_X1 U9069 ( .A(n12831), .ZN(n6935) );
  OR2_X1 U9070 ( .A1(n6903), .A2(n13701), .ZN(n6502) );
  OR2_X1 U9071 ( .A1(n6464), .A2(n7321), .ZN(n6503) );
  INV_X1 U9072 ( .A(n8736), .ZN(n7051) );
  AND2_X1 U9073 ( .A1(n13953), .A2(n12357), .ZN(n6504) );
  AND2_X1 U9074 ( .A1(n12176), .A2(n7284), .ZN(n6505) );
  AND2_X1 U9075 ( .A1(n6923), .A2(n9579), .ZN(n6506) );
  AND2_X1 U9076 ( .A1(n6796), .A2(n6795), .ZN(n6507) );
  AND2_X1 U9077 ( .A1(n7756), .A2(n7755), .ZN(n6508) );
  AND2_X1 U9078 ( .A1(n7555), .A2(n7450), .ZN(n6509) );
  NAND2_X1 U9079 ( .A1(n12978), .A2(n9753), .ZN(n6510) );
  OR2_X1 U9080 ( .A1(n11947), .A2(n11949), .ZN(n6511) );
  AND2_X1 U9081 ( .A1(n13587), .A2(n13121), .ZN(n6512) );
  OR2_X1 U9082 ( .A1(n8636), .A2(n8635), .ZN(n6513) );
  AND2_X1 U9083 ( .A1(n7489), .A2(n7487), .ZN(n6514) );
  OR2_X1 U9084 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n6515) );
  INV_X1 U9085 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8862) );
  NAND2_X1 U9086 ( .A1(n12774), .A2(n12757), .ZN(n6516) );
  AND2_X1 U9087 ( .A1(n11174), .A2(n9149), .ZN(n7495) );
  INV_X1 U9088 ( .A(n12793), .ZN(n9272) );
  AND2_X1 U9089 ( .A1(n9589), .A2(n9597), .ZN(n12793) );
  NOR2_X1 U9090 ( .A1(n7407), .A2(n7408), .ZN(n6517) );
  OR2_X1 U9091 ( .A1(n6728), .A2(n6731), .ZN(n6518) );
  NOR2_X1 U9092 ( .A1(n12381), .A2(n14051), .ZN(n6519) );
  NOR2_X1 U9093 ( .A1(n11835), .A2(n13804), .ZN(n6520) );
  NOR2_X1 U9094 ( .A1(n13603), .A2(n13124), .ZN(n6521) );
  AND2_X1 U9095 ( .A1(n14150), .A2(n14052), .ZN(n6522) );
  AND2_X1 U9096 ( .A1(n9563), .A2(n9562), .ZN(n6523) );
  AND2_X1 U9097 ( .A1(n13422), .A2(n13028), .ZN(n6524) );
  INV_X1 U9098 ( .A(n7279), .ZN(n8325) );
  NAND2_X1 U9099 ( .A1(n7280), .A2(n7318), .ZN(n7279) );
  INV_X1 U9100 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8955) );
  NAND2_X1 U9101 ( .A1(n7093), .A2(n8775), .ZN(n12382) );
  OR2_X1 U9102 ( .A1(n7374), .A2(n6893), .ZN(n6525) );
  AND2_X1 U9103 ( .A1(n13348), .A2(n13040), .ZN(n6526) );
  OR2_X1 U9104 ( .A1(n8808), .A2(n8807), .ZN(n6527) );
  AND2_X1 U9105 ( .A1(n7028), .A2(n7032), .ZN(n6528) );
  NOR2_X1 U9106 ( .A1(n9584), .A2(n10398), .ZN(n6529) );
  AND2_X1 U9107 ( .A1(n12164), .A2(n12544), .ZN(n6530) );
  AND2_X1 U9108 ( .A1(n10548), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n6531) );
  OR2_X1 U9109 ( .A1(n9735), .A2(n11575), .ZN(n6532) );
  OR2_X1 U9110 ( .A1(n7186), .A2(n6809), .ZN(n6533) );
  AND2_X1 U9111 ( .A1(n7612), .A2(SI_9_), .ZN(n6534) );
  INV_X1 U9112 ( .A(n13920), .ZN(n13928) );
  INV_X1 U9113 ( .A(n7542), .ZN(n7541) );
  NAND2_X1 U9114 ( .A1(n8319), .A2(n7543), .ZN(n7542) );
  INV_X1 U9115 ( .A(n14549), .ZN(n14298) );
  NAND2_X1 U9116 ( .A1(n14550), .A2(n14551), .ZN(n14549) );
  INV_X1 U9117 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7701) );
  AND2_X1 U9118 ( .A1(n6881), .A2(n6621), .ZN(n6535) );
  INV_X1 U9119 ( .A(n7536), .ZN(n7535) );
  NAND2_X1 U9120 ( .A1(n12273), .A2(n12266), .ZN(n7536) );
  AND2_X1 U9121 ( .A1(n6755), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6536) );
  NAND2_X1 U9122 ( .A1(n9283), .A2(n9282), .ZN(n12455) );
  INV_X1 U9123 ( .A(n7084), .ZN(n8675) );
  NAND2_X1 U9124 ( .A1(n7085), .A2(n7086), .ZN(n7084) );
  AND2_X1 U9125 ( .A1(n11627), .A2(n8560), .ZN(n6537) );
  AND2_X1 U9126 ( .A1(n8776), .A2(n7372), .ZN(n6538) );
  AND2_X1 U9127 ( .A1(n9881), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n6539) );
  AND2_X1 U9128 ( .A1(n12911), .A2(n12444), .ZN(n6540) );
  INV_X1 U9129 ( .A(n7562), .ZN(n6652) );
  INV_X1 U9130 ( .A(n9238), .ZN(n7498) );
  NAND2_X1 U9131 ( .A1(n7539), .A2(n8862), .ZN(n6541) );
  OR2_X1 U9132 ( .A1(n13102), .A2(n12042), .ZN(n6542) );
  INV_X1 U9133 ( .A(n6885), .ZN(n6884) );
  NOR2_X1 U9134 ( .A1(n13664), .A2(n13801), .ZN(n6885) );
  NAND2_X1 U9135 ( .A1(n13493), .A2(n6800), .ZN(n6543) );
  NOR2_X1 U9136 ( .A1(n11962), .A2(n11963), .ZN(n6544) );
  OR2_X1 U9137 ( .A1(n7380), .A2(n8748), .ZN(n6545) );
  NAND2_X1 U9138 ( .A1(n9549), .A2(n9544), .ZN(n6546) );
  AND2_X1 U9139 ( .A1(n8748), .A2(n7380), .ZN(n6547) );
  NAND2_X1 U9140 ( .A1(n7415), .A2(n12028), .ZN(n6548) );
  NAND2_X1 U9141 ( .A1(n9586), .A2(n9580), .ZN(n6549) );
  NAND2_X1 U9142 ( .A1(n11902), .A2(n11900), .ZN(n7411) );
  OAI21_X1 U9143 ( .B1(n7187), .B2(n7186), .A(n7985), .ZN(n7185) );
  AND2_X1 U9144 ( .A1(n11544), .A2(n11675), .ZN(n6550) );
  AND3_X1 U9145 ( .A1(n9512), .A2(n12679), .A3(n6938), .ZN(n6551) );
  NAND2_X1 U9146 ( .A1(n7343), .A2(n11144), .ZN(n6552) );
  INV_X1 U9147 ( .A(n13964), .ZN(n7220) );
  OR2_X1 U9148 ( .A1(n12026), .A2(n12027), .ZN(n6553) );
  AND2_X1 U9149 ( .A1(n13305), .A2(n7100), .ZN(n6554) );
  NOR2_X1 U9150 ( .A1(n13937), .A2(n7260), .ZN(n6555) );
  NAND2_X1 U9151 ( .A1(n8105), .A2(n8104), .ZN(n13331) );
  OR2_X1 U9152 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n8951), .ZN(n6556) );
  OR2_X1 U9153 ( .A1(n14150), .A2(n14052), .ZN(n6557) );
  OR2_X1 U9154 ( .A1(n14215), .A2(n14214), .ZN(n6558) );
  AND2_X1 U9155 ( .A1(n6925), .A2(n9581), .ZN(n6559) );
  AND2_X1 U9156 ( .A1(n7550), .A2(n7688), .ZN(n7469) );
  OR2_X1 U9157 ( .A1(n13376), .A2(n13123), .ZN(n6560) );
  OR2_X1 U9158 ( .A1(n7646), .A2(n7645), .ZN(n6561) );
  AND3_X1 U9159 ( .A1(n7875), .A2(n7701), .A3(n7692), .ZN(n6562) );
  NOR2_X1 U9160 ( .A1(n8900), .A2(P3_IR_REG_25__SCAN_IN), .ZN(n6563) );
  NOR2_X1 U9161 ( .A1(n9634), .A2(n7127), .ZN(n6564) );
  INV_X1 U9162 ( .A(n8233), .ZN(n7198) );
  AND2_X1 U9163 ( .A1(n12744), .A2(n9609), .ZN(n6565) );
  AND2_X1 U9164 ( .A1(n11723), .A2(n12362), .ZN(n6566) );
  AND2_X1 U9165 ( .A1(n10446), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6567) );
  AND2_X1 U9166 ( .A1(n13988), .A2(n12355), .ZN(n6568) );
  AND2_X1 U9167 ( .A1(n6483), .A2(n8462), .ZN(n6569) );
  AND2_X1 U9168 ( .A1(n7233), .A2(n6469), .ZN(n6570) );
  AND2_X1 U9169 ( .A1(n6915), .A2(n6914), .ZN(n6571) );
  INV_X1 U9170 ( .A(n6812), .ZN(n6811) );
  NOR2_X1 U9171 ( .A1(n13584), .A2(n13120), .ZN(n6812) );
  OR2_X1 U9172 ( .A1(n7062), .A2(n8687), .ZN(n6572) );
  OR2_X1 U9173 ( .A1(n11933), .A2(n11935), .ZN(n6573) );
  AND2_X1 U9174 ( .A1(n6527), .A2(n7369), .ZN(n6574) );
  AND2_X1 U9175 ( .A1(n7299), .A2(n6668), .ZN(n6575) );
  AND2_X1 U9176 ( .A1(n7575), .A2(SI_18_), .ZN(n6576) );
  OR2_X1 U9177 ( .A1(n8417), .A2(n7056), .ZN(n6577) );
  AND2_X1 U9178 ( .A1(n11478), .A2(n7333), .ZN(n6578) );
  OR2_X1 U9179 ( .A1(n8482), .A2(n7059), .ZN(n6579) );
  AND2_X1 U9180 ( .A1(n7171), .A2(n7170), .ZN(n6580) );
  OR2_X1 U9181 ( .A1(n11934), .A2(n11936), .ZN(n6581) );
  NAND2_X1 U9182 ( .A1(n7685), .A2(n7684), .ZN(n7691) );
  OR2_X1 U9183 ( .A1(n11948), .A2(n11950), .ZN(n6582) );
  AND2_X1 U9184 ( .A1(n6542), .A2(n7199), .ZN(n6583) );
  INV_X1 U9185 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7688) );
  OR2_X1 U9186 ( .A1(n6956), .A2(n6475), .ZN(n6584) );
  AND2_X1 U9187 ( .A1(n6563), .A2(n8902), .ZN(n6585) );
  INV_X1 U9188 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6755) );
  INV_X1 U9189 ( .A(n7296), .ZN(n7295) );
  NAND2_X1 U9190 ( .A1(n7297), .A2(n12171), .ZN(n7296) );
  NAND2_X1 U9191 ( .A1(n13505), .A2(n13093), .ZN(n6586) );
  INV_X1 U9192 ( .A(n7374), .ZN(n6897) );
  INV_X1 U9193 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n9138) );
  OR2_X1 U9194 ( .A1(n7516), .A2(n7514), .ZN(n6587) );
  NAND2_X1 U9195 ( .A1(n11681), .A2(n7956), .ZN(n7958) );
  NAND2_X1 U9196 ( .A1(n13749), .A2(n13748), .ZN(n13747) );
  INV_X1 U9197 ( .A(n8654), .ZN(n8645) );
  AND2_X2 U9198 ( .A1(n10724), .A2(n10962), .ZN(n10398) );
  XNOR2_X1 U9199 ( .A(n8838), .B(n13958), .ZN(n13976) );
  INV_X1 U9200 ( .A(n13976), .ZN(n12356) );
  NAND2_X1 U9201 ( .A1(n11222), .A2(n9177), .ZN(n11434) );
  NAND2_X1 U9202 ( .A1(n7263), .A2(n11626), .ZN(n11726) );
  NAND2_X1 U9203 ( .A1(n6704), .A2(n12977), .ZN(n13045) );
  NAND2_X1 U9204 ( .A1(n13705), .A2(n12236), .ZN(n13715) );
  NAND2_X1 U9205 ( .A1(n7474), .A2(n9192), .ZN(n14434) );
  INV_X1 U9206 ( .A(n14036), .ZN(n7266) );
  INV_X1 U9207 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7117) );
  INV_X1 U9208 ( .A(n7987), .ZN(n7646) );
  NAND2_X1 U9209 ( .A1(n9325), .A2(n9324), .ZN(n12504) );
  NAND2_X1 U9210 ( .A1(n12272), .A2(n12271), .ZN(n13758) );
  INV_X1 U9211 ( .A(n13758), .ZN(n6660) );
  NAND2_X1 U9212 ( .A1(n6658), .A2(n12242), .ZN(n13766) );
  NAND2_X1 U9213 ( .A1(n13747), .A2(n12219), .ZN(n14481) );
  OR2_X1 U9214 ( .A1(n12196), .A2(n15087), .ZN(n6588) );
  AND2_X1 U9215 ( .A1(n14443), .A2(n12548), .ZN(n6589) );
  INV_X1 U9216 ( .A(n7108), .ZN(n13461) );
  NOR2_X1 U9217 ( .A1(n11773), .A2(n13617), .ZN(n7108) );
  AND2_X1 U9218 ( .A1(n13435), .A2(n7213), .ZN(n6590) );
  INV_X1 U9219 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7711) );
  INV_X1 U9220 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n6849) );
  AND2_X1 U9221 ( .A1(n9656), .A2(n6588), .ZN(n6591) );
  NAND2_X1 U9222 ( .A1(n11572), .A2(n7465), .ZN(n6592) );
  AND2_X1 U9223 ( .A1(n9038), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n6593) );
  OR2_X1 U9224 ( .A1(n13717), .A2(n13716), .ZN(n6594) );
  AND2_X1 U9225 ( .A1(n7090), .A2(SI_20_), .ZN(n6595) );
  INV_X1 U9226 ( .A(n7224), .ZN(n14059) );
  AND2_X1 U9227 ( .A1(n6917), .A2(n11819), .ZN(n7224) );
  AND2_X1 U9228 ( .A1(n7298), .A2(n7295), .ZN(n6596) );
  INV_X1 U9229 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9848) );
  INV_X1 U9230 ( .A(n8040), .ZN(n7363) );
  AND2_X1 U9231 ( .A1(n10425), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n6597) );
  OR2_X1 U9232 ( .A1(n8052), .A2(n7363), .ZN(n6598) );
  INV_X1 U9233 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7317) );
  INV_X1 U9234 ( .A(n7960), .ZN(n7379) );
  INV_X1 U9235 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8896) );
  OR2_X1 U9236 ( .A1(n9661), .A2(n9784), .ZN(n14858) );
  AND2_X1 U9237 ( .A1(n8909), .A2(n12952), .ZN(n9115) );
  XNOR2_X1 U9238 ( .A(n8871), .B(n8870), .ZN(n10221) );
  INV_X1 U9239 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6640) );
  INV_X1 U9240 ( .A(n15157), .ZN(n15154) );
  AND2_X1 U9241 ( .A1(n9448), .A2(n9447), .ZN(n15142) );
  INV_X1 U9242 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7250) );
  NAND2_X1 U9243 ( .A1(n8979), .A2(n8978), .ZN(n12762) );
  INV_X1 U9244 ( .A(n12762), .ZN(n6818) );
  INV_X1 U9245 ( .A(n9048), .ZN(n9060) );
  NAND2_X1 U9246 ( .A1(n11117), .A2(n7557), .ZN(n11189) );
  INV_X1 U9247 ( .A(n9223), .ZN(n7243) );
  XNOR2_X1 U9248 ( .A(n8320), .B(P1_IR_REG_22__SCAN_IN), .ZN(n8820) );
  NAND2_X1 U9249 ( .A1(n14334), .A2(n7160), .ZN(n7157) );
  OR2_X1 U9250 ( .A1(n14336), .A2(n12214), .ZN(n6599) );
  NAND2_X1 U9251 ( .A1(n7099), .A2(n7096), .ZN(n6600) );
  AND2_X1 U9252 ( .A1(n8880), .A2(n8879), .ZN(n10222) );
  OAI21_X1 U9253 ( .B1(n13077), .B2(n13076), .A(n9699), .ZN(n10835) );
  XNOR2_X1 U9254 ( .A(n6667), .B(n11822), .ZN(n11824) );
  OAI21_X1 U9255 ( .B1(n11824), .B2(n11823), .A(n6666), .ZN(n14493) );
  NAND2_X1 U9256 ( .A1(n10989), .A2(n8233), .ZN(n11232) );
  AND2_X1 U9257 ( .A1(n7020), .A2(n7023), .ZN(n6601) );
  NAND2_X1 U9258 ( .A1(n11042), .A2(n7495), .ZN(n11173) );
  INV_X1 U9259 ( .A(n13551), .ZN(n7107) );
  AND2_X1 U9260 ( .A1(n7312), .A2(n7311), .ZN(n6602) );
  INV_X1 U9261 ( .A(n14396), .ZN(n7004) );
  NAND2_X1 U9262 ( .A1(n9148), .A2(n9147), .ZN(n11042) );
  AND2_X1 U9263 ( .A1(n7523), .A2(n7520), .ZN(n6603) );
  AND2_X1 U9264 ( .A1(n7669), .A2(n11523), .ZN(n6604) );
  INV_X1 U9265 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11376) );
  NAND2_X1 U9266 ( .A1(n15339), .A2(n7550), .ZN(n8199) );
  INV_X1 U9267 ( .A(n13430), .ZN(n13454) );
  INV_X1 U9268 ( .A(SI_19_), .ZN(n7091) );
  NOR2_X1 U9269 ( .A1(n9661), .A2(n14831), .ZN(n13552) );
  INV_X1 U9270 ( .A(n14739), .ZN(n6900) );
  INV_X1 U9271 ( .A(n7114), .ZN(n10718) );
  INV_X1 U9272 ( .A(n10629), .ZN(n6744) );
  OAI21_X1 U9273 ( .B1(n10686), .B2(n6757), .A(n10685), .ZN(n10739) );
  NAND2_X1 U9274 ( .A1(n10741), .A2(n10740), .ZN(n10816) );
  AND2_X1 U9275 ( .A1(n12624), .A2(n12650), .ZN(n6605) );
  INV_X1 U9276 ( .A(n12651), .ZN(n14413) );
  NAND2_X1 U9277 ( .A1(n8301), .A2(n8296), .ZN(n8882) );
  NOR2_X1 U9278 ( .A1(n7455), .A2(n10509), .ZN(n7454) );
  INV_X1 U9279 ( .A(n7013), .ZN(n7011) );
  NOR2_X1 U9280 ( .A1(n7017), .A2(n7014), .ZN(n7013) );
  AND2_X1 U9281 ( .A1(n6649), .A2(n6647), .ZN(n6606) );
  AND2_X1 U9282 ( .A1(n7456), .A2(n7454), .ZN(n6607) );
  AND2_X1 U9283 ( .A1(n7427), .A2(n9675), .ZN(n6608) );
  AND2_X1 U9284 ( .A1(n14393), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n6609) );
  NAND2_X1 U9285 ( .A1(n11859), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6610) );
  INV_X1 U9286 ( .A(SI_22_), .ZN(n7386) );
  NOR2_X1 U9287 ( .A1(n10629), .A2(n12149), .ZN(n6743) );
  XNOR2_X1 U9288 ( .A(n9279), .B(n7117), .ZN(n12596) );
  AND2_X1 U9289 ( .A1(n13633), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6611) );
  INV_X1 U9290 ( .A(n14207), .ZN(n6762) );
  INV_X1 U9291 ( .A(SI_5_), .ZN(n7079) );
  NOR2_X1 U9292 ( .A1(n8806), .A2(n8637), .ZN(n7359) );
  NAND2_X1 U9293 ( .A1(n6614), .A2(n9254), .ZN(n12824) );
  NAND2_X2 U9294 ( .A1(n10892), .A2(n9096), .ZN(n10891) );
  NAND3_X1 U9295 ( .A1(n7501), .A2(n6585), .A3(n8987), .ZN(n12944) );
  AND4_X4 U9296 ( .A1(n6431), .A2(n9061), .A3(n7313), .A4(n8895), .ZN(n8987)
         );
  AND2_X2 U9297 ( .A1(n10417), .A2(n8892), .ZN(n9061) );
  NAND3_X1 U9298 ( .A1(n7136), .A2(n6616), .A3(n7135), .ZN(n7139) );
  NAND2_X1 U9299 ( .A1(n7136), .A2(n6616), .ZN(n15326) );
  NAND2_X1 U9300 ( .A1(n6617), .A2(n14558), .ZN(n14359) );
  NAND2_X1 U9301 ( .A1(n14560), .A2(n14559), .ZN(n14558) );
  NAND2_X1 U9302 ( .A1(n6618), .A2(n14545), .ZN(n14550) );
  NAND2_X1 U9303 ( .A1(n14546), .A2(n14547), .ZN(n14545) );
  INV_X1 U9304 ( .A(n7323), .ZN(n6626) );
  INV_X1 U9305 ( .A(n8304), .ZN(n14186) );
  NAND3_X1 U9306 ( .A1(n11724), .A2(n12365), .A3(n6566), .ZN(n6632) );
  NAND2_X1 U9307 ( .A1(n7574), .A2(n14036), .ZN(n14035) );
  XNOR2_X1 U9308 ( .A(n6637), .B(n12596), .ZN(n9517) );
  NAND3_X1 U9309 ( .A1(n9513), .A2(n6866), .A3(n6551), .ZN(n6638) );
  NAND3_X1 U9310 ( .A1(n6651), .A2(n6652), .A3(n6650), .ZN(n6646) );
  XNOR2_X1 U9311 ( .A(n10918), .B(n10919), .ZN(n10920) );
  OR2_X1 U9312 ( .A1(n6667), .A2(n11822), .ZN(n6666) );
  NAND3_X1 U9313 ( .A1(n7307), .A2(n6444), .A3(n7306), .ZN(n6669) );
  NAND2_X1 U9314 ( .A1(n12478), .A2(n6675), .ZN(n6672) );
  NAND2_X1 U9315 ( .A1(n6672), .A2(n6673), .ZN(n12450) );
  NAND2_X1 U9316 ( .A1(n12501), .A2(n12176), .ZN(n12178) );
  NAND2_X1 U9317 ( .A1(n14369), .A2(n7170), .ZN(n6687) );
  INV_X1 U9318 ( .A(n12591), .ZN(n6688) );
  INV_X1 U9319 ( .A(n14369), .ZN(n6689) );
  NAND2_X1 U9320 ( .A1(n6872), .A2(n6691), .ZN(n14917) );
  INV_X1 U9321 ( .A(n6691), .ZN(n10448) );
  NAND4_X1 U9322 ( .A1(n6692), .A2(n14432), .A3(n14431), .A4(n14433), .ZN(
        P3_U3200) );
  NAND4_X1 U9323 ( .A1(n9061), .A2(n6431), .A3(n8896), .A4(n8895), .ZN(n9209)
         );
  NAND2_X1 U9324 ( .A1(n7713), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7714) );
  AOI21_X2 U9327 ( .B1(n6707), .B2(n6489), .A(n6702), .ZN(n13000) );
  NAND2_X1 U9328 ( .A1(n7440), .A2(n13103), .ZN(n6707) );
  NOR2_X1 U9329 ( .A1(n13038), .A2(n13037), .ZN(n13036) );
  NAND4_X2 U9330 ( .A1(n7733), .A2(n7732), .A3(n7730), .A4(n7731), .ZN(n13143)
         );
  INV_X1 U9331 ( .A(n12098), .ZN(n12141) );
  OAI21_X1 U9332 ( .B1(n6501), .B2(n6717), .A(n7392), .ZN(n6716) );
  NAND2_X1 U9333 ( .A1(n7395), .A2(n7393), .ZN(n6717) );
  NAND2_X1 U9334 ( .A1(n12069), .A2(n12068), .ZN(n7387) );
  NAND2_X1 U9335 ( .A1(n12046), .A2(n6718), .ZN(n12069) );
  NAND2_X1 U9336 ( .A1(n6719), .A2(n12043), .ZN(n6718) );
  NAND3_X1 U9337 ( .A1(n7405), .A2(n7404), .A3(n6487), .ZN(n12045) );
  NAND4_X1 U9338 ( .A1(n7405), .A2(n7404), .A3(n6487), .A4(n6720), .ZN(n6719)
         );
  NAND2_X1 U9339 ( .A1(n6722), .A2(n6721), .ZN(n11972) );
  NAND2_X1 U9340 ( .A1(n7398), .A2(n6732), .ZN(n6730) );
  AND2_X1 U9341 ( .A1(n6733), .A2(n7396), .ZN(n6732) );
  NAND3_X1 U9342 ( .A1(n6736), .A2(n6582), .A3(n6734), .ZN(n7423) );
  NAND2_X1 U9343 ( .A1(n6735), .A2(n11943), .ZN(n6734) );
  INV_X1 U9344 ( .A(n6738), .ZN(n6735) );
  NAND2_X1 U9345 ( .A1(n6737), .A2(n11941), .ZN(n6736) );
  NAND2_X1 U9346 ( .A1(n6738), .A2(n11942), .ZN(n6737) );
  NAND2_X1 U9347 ( .A1(n7422), .A2(n6573), .ZN(n6738) );
  NAND3_X1 U9348 ( .A1(n7414), .A2(n7416), .A3(n6553), .ZN(n6739) );
  NOR2_X1 U9349 ( .A1(n12149), .A2(n12138), .ZN(n6742) );
  NOR2_X1 U9350 ( .A1(n11884), .A2(n6496), .ZN(n6748) );
  OAI21_X1 U9351 ( .B1(n11885), .B2(n6748), .A(n6749), .ZN(n11892) );
  NAND2_X1 U9352 ( .A1(n11892), .A2(n11893), .ZN(n11891) );
  NOR2_X2 U9353 ( .A1(n7680), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n6750) );
  INV_X2 U9354 ( .A(n7759), .ZN(n7679) );
  NAND2_X1 U9355 ( .A1(n10980), .A2(n10979), .ZN(n11151) );
  NAND2_X1 U9356 ( .A1(n11075), .A2(n11079), .ZN(n11074) );
  NAND2_X1 U9357 ( .A1(n11154), .A2(n7253), .ZN(n6752) );
  NAND2_X1 U9358 ( .A1(n11251), .A2(n11250), .ZN(n11249) );
  NAND2_X2 U9359 ( .A1(n13990), .A2(n13989), .ZN(n13988) );
  OAI21_X2 U9360 ( .B1(n6754), .B2(n6536), .A(n8298), .ZN(n14197) );
  NAND3_X1 U9361 ( .A1(n6756), .A2(n8333), .A3(n8331), .ZN(n13813) );
  AND2_X1 U9362 ( .A1(n8341), .A2(n8340), .ZN(n6759) );
  OAI21_X1 U9363 ( .B1(n13938), .B2(n7258), .A(n7256), .ZN(n12398) );
  OAI21_X2 U9364 ( .B1(n11731), .B2(n6764), .A(n6763), .ZN(n14047) );
  OAI21_X1 U9365 ( .B1(n14079), .B2(n14153), .A(n14078), .ZN(n14171) );
  OAI211_X1 U9366 ( .C1(n6770), .C2(n14079), .A(n6768), .B(n6773), .ZN(
        P1_U3525) );
  OR2_X1 U9367 ( .A1(n15160), .A2(n6774), .ZN(n6773) );
  NAND2_X1 U9368 ( .A1(n6775), .A2(n7591), .ZN(n7594) );
  XNOR2_X1 U9369 ( .A(n6775), .B(n7762), .ZN(n9855) );
  NAND2_X1 U9370 ( .A1(n7590), .A2(n7589), .ZN(n6775) );
  NAND2_X1 U9371 ( .A1(n6776), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n7579) );
  NAND3_X1 U9372 ( .A1(n13254), .A2(n13893), .A3(n6777), .ZN(n6776) );
  NAND2_X1 U9373 ( .A1(n6778), .A2(n6586), .ZN(n6779) );
  NAND2_X1 U9374 ( .A1(n13312), .A2(n6812), .ZN(n6778) );
  AOI21_X1 U9375 ( .B1(n6782), .B2(n6780), .A(n6779), .ZN(n13294) );
  OR2_X1 U9376 ( .A1(n13340), .A2(n6466), .ZN(n6782) );
  MUX2_X1 U9377 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n9834), .Z(n7602) );
  MUX2_X1 U9378 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n9834), .Z(n7601) );
  NAND3_X1 U9379 ( .A1(n6804), .A2(n6803), .A3(n6560), .ZN(n6787) );
  OR2_X1 U9380 ( .A1(n6838), .A2(n13454), .ZN(n6791) );
  NAND2_X1 U9381 ( .A1(n15339), .A2(n7469), .ZN(n6792) );
  NAND2_X2 U9382 ( .A1(n6829), .A2(n6794), .ZN(n8179) );
  OAI22_X1 U9383 ( .A1(n6799), .A2(n6798), .B1(n13430), .B2(n13284), .ZN(
        n13494) );
  NAND2_X1 U9384 ( .A1(n11681), .A2(n6808), .ZN(n6807) );
  INV_X1 U9385 ( .A(n7986), .ZN(n6810) );
  OAI21_X2 U9386 ( .B1(n13294), .B2(n12100), .A(n8140), .ZN(n13283) );
  NAND2_X1 U9387 ( .A1(n10197), .A2(n7736), .ZN(n10653) );
  NAND2_X1 U9388 ( .A1(n10198), .A2(n12106), .ZN(n10197) );
  NAND2_X1 U9389 ( .A1(n11729), .A2(n11728), .ZN(n11731) );
  NAND2_X1 U9390 ( .A1(n11461), .A2(n7923), .ZN(n11607) );
  NAND2_X1 U9391 ( .A1(n11589), .A2(n11588), .ZN(n14348) );
  XNOR2_X2 U9392 ( .A(n13811), .B(n14562), .ZN(n10820) );
  NAND2_X1 U9393 ( .A1(n10859), .A2(n10746), .ZN(n10748) );
  AOI21_X2 U9394 ( .B1(n12349), .B2(n6453), .A(n6519), .ZN(n7570) );
  NOR2_X2 U9395 ( .A1(n12397), .A2(n6832), .ZN(n13908) );
  OR2_X1 U9396 ( .A1(n10918), .A2(n10919), .ZN(n6816) );
  AOI21_X1 U9397 ( .B1(n10816), .B2(n10743), .A(n10742), .ZN(n10945) );
  INV_X1 U9398 ( .A(n6936), .ZN(n8956) );
  NAND2_X1 U9399 ( .A1(n11606), .A2(n7936), .ZN(n11681) );
  NAND2_X1 U9400 ( .A1(n8241), .A2(n8240), .ZN(n11683) );
  OAI21_X1 U9401 ( .B1(n8255), .B2(n7201), .A(n6583), .ZN(n13281) );
  NAND2_X1 U9402 ( .A1(n11766), .A2(n12124), .ZN(n8245) );
  AOI21_X1 U9403 ( .B1(n13364), .B2(n13365), .A(n8083), .ZN(n13340) );
  AND3_X1 U9404 ( .A1(n7739), .A2(n7741), .A3(n7740), .ZN(n6820) );
  NAND2_X1 U9405 ( .A1(n7788), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7720) );
  NAND2_X1 U9406 ( .A1(n10770), .A2(n10769), .ZN(n10768) );
  NAND2_X1 U9407 ( .A1(n7608), .A2(n7607), .ZN(n7837) );
  NAND2_X1 U9408 ( .A1(n6896), .A2(n7375), .ZN(n7989) );
  INV_X1 U9409 ( .A(n11811), .ZN(n7330) );
  NAND2_X1 U9410 ( .A1(n14048), .A2(n7329), .ZN(n7328) );
  OAI22_X2 U9411 ( .A1(n12964), .A2(n12965), .B1(n9767), .B2(n9766), .ZN(
        n13038) );
  NAND2_X1 U9412 ( .A1(n10835), .A2(n10836), .ZN(n7468) );
  NAND2_X1 U9413 ( .A1(n11476), .A2(n11482), .ZN(n11589) );
  INV_X1 U9414 ( .A(n10689), .ZN(n14676) );
  NAND2_X1 U9415 ( .A1(n14308), .A2(n14307), .ZN(n14309) );
  NOR2_X1 U9416 ( .A1(n14298), .A2(n6486), .ZN(n7133) );
  XNOR2_X1 U9417 ( .A(n14278), .B(n14277), .ZN(n14326) );
  OAI21_X1 U9418 ( .B1(n12495), .B2(n7296), .A(n7292), .ZN(n12175) );
  NAND2_X1 U9419 ( .A1(n12433), .A2(n12434), .ZN(n12432) );
  AOI21_X1 U9420 ( .B1(n11800), .B2(n11799), .A(n7559), .ZN(n12160) );
  NAND2_X1 U9421 ( .A1(n13788), .A2(n13787), .ZN(n13786) );
  INV_X4 U9422 ( .A(n8343), .ZN(n8637) );
  NOR2_X2 U9423 ( .A1(n8297), .A2(n7344), .ZN(n8304) );
  NAND2_X1 U9424 ( .A1(n7222), .A2(n7280), .ZN(n8297) );
  XNOR2_X2 U9425 ( .A(n11869), .B(n11872), .ZN(n12106) );
  INV_X1 U9426 ( .A(n11889), .ZN(n6828) );
  OAI211_X1 U9427 ( .C1(n13269), .C2(n13270), .A(n13268), .B(n6846), .ZN(n6845) );
  INV_X1 U9428 ( .A(n6845), .ZN(n13491) );
  NAND2_X1 U9429 ( .A1(n11607), .A2(n12122), .ZN(n11606) );
  NAND2_X1 U9430 ( .A1(n10768), .A2(n7778), .ZN(n10601) );
  INV_X1 U9431 ( .A(n7725), .ZN(n7103) );
  XNOR2_X2 U9432 ( .A(n8303), .B(n8302), .ZN(n12154) );
  NAND2_X1 U9433 ( .A1(n8938), .A2(n8937), .ZN(n9224) );
  OAI21_X2 U9434 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n8950), .A(n8949), .ZN(
        n8951) );
  NAND2_X1 U9435 ( .A1(n9293), .A2(n9292), .ZN(n7251) );
  OAI211_X1 U9436 ( .C1(n9644), .C2(n9459), .A(n9646), .B(n6963), .ZN(n6962)
         );
  NAND2_X1 U9437 ( .A1(n6837), .A2(n6834), .ZN(P1_U3214) );
  NAND2_X1 U9438 ( .A1(n13658), .A2(n14580), .ZN(n6837) );
  AND2_X1 U9439 ( .A1(n11011), .A2(n11010), .ZN(n7573) );
  NAND2_X1 U9440 ( .A1(n6876), .A2(n7577), .ZN(n7578) );
  NAND2_X1 U9441 ( .A1(n7378), .A2(n7637), .ZN(n7974) );
  AOI21_X1 U9442 ( .B1(n12014), .B2(n12013), .A(n12012), .ZN(n12015) );
  OAI21_X1 U9443 ( .B1(n12144), .B2(n12143), .A(n12142), .ZN(n12151) );
  INV_X1 U9444 ( .A(n7457), .ZN(n7455) );
  OAI22_X1 U9445 ( .A1(n11294), .A2(n11293), .B1(n9718), .B2(n9717), .ZN(
        n11424) );
  OAI21_X1 U9446 ( .B1(n6839), .B2(n12988), .A(n9805), .ZN(P2_U3186) );
  NAND2_X1 U9447 ( .A1(n9790), .A2(n9789), .ZN(n6839) );
  NAND2_X1 U9448 ( .A1(n8261), .A2(n13249), .ZN(n9668) );
  OAI211_X1 U9449 ( .C1(n6470), .C2(n7453), .A(n9688), .B(n7451), .ZN(n10621)
         );
  NAND2_X1 U9450 ( .A1(n6518), .A2(n7401), .ZN(n7404) );
  OAI21_X1 U9451 ( .B1(n12022), .B2(n12021), .A(n12020), .ZN(n7414) );
  OR2_X1 U9452 ( .A1(n13012), .A2(n6873), .ZN(P2_U3197) );
  NOR2_X1 U9453 ( .A1(n13009), .A2(n13011), .ZN(n13010) );
  NAND2_X1 U9454 ( .A1(n6844), .A2(n6842), .ZN(P2_U3237) );
  NAND2_X1 U9455 ( .A1(n13274), .A2(n13468), .ZN(n6844) );
  INV_X1 U9456 ( .A(n10417), .ZN(n6851) );
  OAI21_X1 U9457 ( .B1(n8338), .B2(n8779), .A(n8339), .ZN(n6848) );
  INV_X1 U9458 ( .A(n7153), .ZN(n7152) );
  NAND3_X1 U9459 ( .A1(n7147), .A2(n7144), .A3(n7148), .ZN(n14296) );
  NOR2_X1 U9460 ( .A1(n14370), .A2(n14371), .ZN(n14369) );
  NOR2_X1 U9461 ( .A1(n14932), .A2(n12583), .ZN(n14960) );
  NAND2_X1 U9462 ( .A1(n7651), .A2(n7650), .ZN(n8004) );
  NAND2_X1 U9463 ( .A1(n7087), .A2(n7090), .ZN(n7654) );
  AOI21_X1 U9464 ( .B1(n12141), .B2(n6744), .A(n12140), .ZN(n12143) );
  NAND2_X1 U9465 ( .A1(n11151), .A2(n11150), .ZN(n11251) );
  INV_X1 U9466 ( .A(n7069), .ZN(n7068) );
  XNOR2_X1 U9467 ( .A(n7630), .B(SI_14_), .ZN(n7937) );
  NAND2_X1 U9468 ( .A1(n7400), .A2(n7399), .ZN(n7398) );
  NAND2_X1 U9469 ( .A1(n7891), .A2(n7620), .ZN(n7070) );
  NOR2_X1 U9470 ( .A1(n14404), .A2(n14405), .ZN(n14403) );
  NOR2_X1 U9471 ( .A1(n14917), .A2(n14918), .ZN(n14916) );
  INV_X1 U9472 ( .A(n7746), .ZN(n7104) );
  OAI21_X2 U9473 ( .B1(n12650), .B2(n12888), .A(n14388), .ZN(n12652) );
  OAI21_X2 U9474 ( .B1(n12641), .B2(n12640), .A(n14950), .ZN(n12642) );
  NOR2_X2 U9475 ( .A1(n14910), .A2(n14909), .ZN(n14908) );
  OAI21_X1 U9476 ( .B1(n12569), .B2(P3_REG1_REG_2__SCAN_IN), .A(n6853), .ZN(
        n12563) );
  NAND2_X1 U9477 ( .A1(n13497), .A2(n6857), .ZN(P2_U3526) );
  NAND2_X1 U9478 ( .A1(n13571), .A2(n6859), .ZN(P2_U3494) );
  NAND2_X1 U9479 ( .A1(n8020), .A2(n8019), .ZN(n13400) );
  NAND2_X1 U9480 ( .A1(n13491), .A2(n6867), .ZN(n13566) );
  NAND2_X1 U9481 ( .A1(n13491), .A2(n6862), .ZN(n13274) );
  OAI22_X1 U9482 ( .A1(n7724), .A2(n9830), .B1(n7742), .B2(n9938), .ZN(n7725)
         );
  XNOR2_X1 U9483 ( .A(n7177), .B(n12134), .ZN(n8187) );
  XNOR2_X2 U9484 ( .A(n8344), .B(P1_IR_REG_1__SCAN_IN), .ZN(n10013) );
  OAI21_X1 U9485 ( .B1(P1_DATAO_REG_19__SCAN_IN), .B2(n12155), .A(n8946), .ZN(
        n9293) );
  OAI21_X1 U9486 ( .B1(n9353), .B2(n9352), .A(n7270), .ZN(n7269) );
  OAI21_X1 U9487 ( .B1(P1_DATAO_REG_22__SCAN_IN), .B2(n8948), .A(n8947), .ZN(
        n9316) );
  NAND2_X1 U9488 ( .A1(n9072), .A2(n9071), .ZN(n8925) );
  NAND2_X1 U9489 ( .A1(n6865), .A2(n9650), .ZN(P3_U3296) );
  OAI21_X1 U9490 ( .B1(n6962), .B2(n9648), .A(n9647), .ZN(n6865) );
  NAND2_X1 U9491 ( .A1(n12589), .A2(n12618), .ZN(n12590) );
  NOR2_X1 U9492 ( .A1(n14403), .A2(n12594), .ZN(n14430) );
  NAND2_X2 U9493 ( .A1(n7579), .A2(n7578), .ZN(n7595) );
  NAND3_X1 U9494 ( .A1(n7576), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n6876) );
  INV_X1 U9495 ( .A(n7063), .ZN(n6880) );
  INV_X1 U9496 ( .A(n6887), .ZN(n6886) );
  OAI21_X1 U9497 ( .B1(n7656), .B2(n8052), .A(n7659), .ZN(n6887) );
  NAND2_X1 U9498 ( .A1(n7633), .A2(n6888), .ZN(n6890) );
  NAND3_X1 U9499 ( .A1(n7632), .A2(n7633), .A3(n6897), .ZN(n6896) );
  INV_X1 U9500 ( .A(n10817), .ZN(n6906) );
  NAND2_X1 U9501 ( .A1(n10818), .A2(n6905), .ZN(n6907) );
  INV_X1 U9502 ( .A(n6911), .ZN(n14015) );
  NAND3_X1 U9503 ( .A1(n6916), .A2(n14084), .A3(n6571), .ZN(n14172) );
  NAND2_X1 U9504 ( .A1(n14442), .A2(n6559), .ZN(n6924) );
  NAND3_X1 U9505 ( .A1(n6925), .A2(n6927), .A3(n9581), .ZN(n6923) );
  OAI21_X2 U9506 ( .B1(n9409), .B2(n9620), .A(n12700), .ZN(n12710) );
  NOR2_X2 U9507 ( .A1(n12727), .A2(n12728), .ZN(n9409) );
  NAND2_X1 U9508 ( .A1(n12830), .A2(n6934), .ZN(n6933) );
  NAND3_X1 U9509 ( .A1(n7501), .A2(n8987), .A3(n6563), .ZN(n6936) );
  NAND2_X1 U9510 ( .A1(n10732), .A2(n15086), .ZN(n9531) );
  NAND2_X1 U9511 ( .A1(n12556), .A2(n15108), .ZN(n9535) );
  AND2_X1 U9512 ( .A1(n9064), .A2(n9065), .ZN(n6937) );
  NAND2_X1 U9513 ( .A1(n9278), .A2(n6946), .ZN(n9379) );
  NAND2_X1 U9514 ( .A1(n6948), .A2(n6565), .ZN(n9613) );
  NAND3_X1 U9515 ( .A1(n6949), .A2(n9605), .A3(n9606), .ZN(n6948) );
  OAI211_X1 U9516 ( .C1(n9602), .C2(n10398), .A(n9406), .B(n6950), .ZN(n6949)
         );
  NAND2_X1 U9517 ( .A1(n6461), .A2(n10398), .ZN(n6950) );
  OR2_X1 U9518 ( .A1(n9564), .A2(n6584), .ZN(n6953) );
  INV_X1 U9519 ( .A(n11433), .ZN(n6961) );
  NAND2_X1 U9520 ( .A1(n6964), .A2(n6965), .ZN(n9588) );
  NAND2_X1 U9521 ( .A1(n9582), .A2(n6967), .ZN(n6964) );
  INV_X1 U9522 ( .A(n9579), .ZN(n6975) );
  NAND2_X1 U9523 ( .A1(n9547), .A2(n6982), .ZN(n6977) );
  NAND2_X1 U9524 ( .A1(n6976), .A2(n6984), .ZN(n9558) );
  NAND4_X1 U9525 ( .A1(n6978), .A2(n6977), .A3(n6986), .A4(n6979), .ZN(n6976)
         );
  NAND2_X1 U9526 ( .A1(n6990), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6991) );
  NAND4_X1 U9527 ( .A1(n7501), .A2(n8987), .A3(n8954), .A4(n7500), .ZN(n6990)
         );
  NAND2_X1 U9528 ( .A1(n7001), .A2(n6999), .ZN(n12629) );
  NAND2_X1 U9529 ( .A1(n14379), .A2(n7000), .ZN(n6999) );
  NAND2_X1 U9530 ( .A1(n7021), .A2(n14884), .ZN(n7019) );
  NAND3_X1 U9531 ( .A1(n7019), .A2(n7018), .A3(n10472), .ZN(n10543) );
  NAND2_X1 U9532 ( .A1(n14884), .A2(n7025), .ZN(n7020) );
  AOI21_X1 U9533 ( .B1(n7023), .B2(n14902), .A(n14919), .ZN(n7021) );
  INV_X1 U9534 ( .A(n7023), .ZN(n7022) );
  INV_X1 U9535 ( .A(n7026), .ZN(n14903) );
  INV_X1 U9536 ( .A(n14902), .ZN(n7025) );
  NAND3_X1 U9537 ( .A1(n8768), .A2(n8767), .A3(n7370), .ZN(n7027) );
  NAND3_X1 U9538 ( .A1(n8436), .A2(n8435), .A3(n6483), .ZN(n7028) );
  AND2_X1 U9539 ( .A1(n7031), .A2(n7029), .ZN(n8461) );
  NAND2_X1 U9540 ( .A1(n7030), .A2(n8462), .ZN(n7029) );
  NAND3_X1 U9541 ( .A1(n8436), .A2(n8435), .A3(n6569), .ZN(n7031) );
  INV_X1 U9542 ( .A(n8448), .ZN(n7033) );
  MUX2_X1 U9543 ( .A(n7038), .B(n7037), .S(n8800), .Z(n7036) );
  NAND2_X1 U9544 ( .A1(n7040), .A2(n7041), .ZN(n8649) );
  NAND2_X1 U9545 ( .A1(n8561), .A2(n7045), .ZN(n7040) );
  NOR2_X1 U9546 ( .A1(n7042), .A2(n6513), .ZN(n7041) );
  NAND2_X1 U9547 ( .A1(n8735), .A2(n6449), .ZN(n7048) );
  NAND2_X1 U9548 ( .A1(n7048), .A2(n7049), .ZN(n8763) );
  NAND2_X1 U9549 ( .A1(n7054), .A2(n7055), .ZN(n8431) );
  NAND3_X1 U9550 ( .A1(n8401), .A2(n8400), .A3(n6577), .ZN(n7054) );
  NAND2_X1 U9551 ( .A1(n7057), .A2(n7058), .ZN(n8498) );
  NAND3_X1 U9552 ( .A1(n8465), .A2(n6579), .A3(n8464), .ZN(n7057) );
  NAND2_X1 U9553 ( .A1(n7060), .A2(n7061), .ZN(n8701) );
  NAND3_X1 U9554 ( .A1(n7355), .A2(n6572), .A3(n8686), .ZN(n7060) );
  OAI21_X1 U9555 ( .B1(n7892), .B2(n7068), .A(n7065), .ZN(n7924) );
  OAI21_X1 U9556 ( .B1(n7892), .B2(n7891), .A(n7620), .ZN(n7906) );
  NAND3_X1 U9557 ( .A1(n7072), .A2(n8861), .A3(n7071), .ZN(n8866) );
  NAND2_X1 U9558 ( .A1(n7648), .A2(n7075), .ZN(n8001) );
  INV_X1 U9559 ( .A(n8001), .ZN(n7651) );
  NAND2_X1 U9560 ( .A1(n8086), .A2(n6442), .ZN(n7080) );
  NAND2_X1 U9561 ( .A1(n7080), .A2(n7081), .ZN(n8129) );
  NAND2_X1 U9562 ( .A1(n8086), .A2(n7663), .ZN(n8103) );
  NAND2_X1 U9563 ( .A1(n7088), .A2(n8004), .ZN(n7087) );
  MUX2_X1 U9564 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n9834), .Z(n7597) );
  NAND2_X1 U9565 ( .A1(n13632), .A2(n8745), .ZN(n7093) );
  XNOR2_X1 U9566 ( .A(n8792), .B(n8791), .ZN(n13632) );
  NAND2_X1 U9567 ( .A1(n7099), .A2(n7094), .ZN(n10993) );
  NOR2_X1 U9568 ( .A1(n11907), .A2(n7095), .ZN(n7094) );
  NOR2_X1 U9569 ( .A1(n13080), .A2(n14844), .ZN(n7098) );
  INV_X1 U9570 ( .A(n13564), .ZN(n7101) );
  NAND3_X1 U9571 ( .A1(n6554), .A2(n12060), .A3(n7101), .ZN(n13257) );
  AND2_X1 U9572 ( .A1(n11883), .A2(n10656), .ZN(n10657) );
  NOR2_X2 U9573 ( .A1(n11869), .A2(n11862), .ZN(n10656) );
  NAND2_X1 U9574 ( .A1(n13358), .A2(n13348), .ZN(n13347) );
  AND2_X2 U9575 ( .A1(n7106), .A2(n13385), .ZN(n13358) );
  INV_X1 U9576 ( .A(n13347), .ZN(n7105) );
  NAND2_X1 U9577 ( .A1(n7105), .A2(n13584), .ZN(n13317) );
  NOR2_X2 U9578 ( .A1(n11602), .A2(n11969), .ZN(n11684) );
  NAND2_X1 U9579 ( .A1(n12738), .A2(n9615), .ZN(n9408) );
  NAND2_X1 U9580 ( .A1(n12749), .A2(n9610), .ZN(n7109) );
  OAI21_X1 U9581 ( .B1(n7112), .B2(n7110), .A(n9539), .ZN(n10889) );
  NAND2_X1 U9582 ( .A1(n7111), .A2(n9531), .ZN(n15060) );
  NAND2_X1 U9583 ( .A1(n9500), .A2(n7113), .ZN(n7112) );
  NAND2_X1 U9584 ( .A1(n7114), .A2(n9531), .ZN(n7113) );
  NAND4_X1 U9585 ( .A1(n8897), .A2(n8988), .A3(n9382), .A4(n7117), .ZN(n7116)
         );
  NAND4_X1 U9586 ( .A1(n7120), .A2(n7119), .A3(n9376), .A4(n8898), .ZN(n7118)
         );
  NAND2_X1 U9587 ( .A1(n12710), .A2(n6564), .ZN(n7126) );
  NAND2_X1 U9588 ( .A1(n12710), .A2(n7129), .ZN(n7128) );
  INV_X1 U9589 ( .A(n15082), .ZN(n9523) );
  NAND2_X1 U9590 ( .A1(n10504), .A2(n12557), .ZN(n9527) );
  OAI21_X2 U9591 ( .B1(n12787), .B2(n12786), .A(n9598), .ZN(n12772) );
  NAND2_X1 U9592 ( .A1(n14549), .A2(n7134), .ZN(n7132) );
  INV_X1 U9593 ( .A(n14555), .ZN(n14554) );
  NOR2_X1 U9594 ( .A1(n14324), .A2(n14279), .ZN(n14281) );
  OAI21_X1 U9595 ( .B1(n14324), .B2(n14279), .A(P2_ADDR_REG_7__SCAN_IN), .ZN(
        n7136) );
  NOR2_X1 U9596 ( .A1(n14279), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7137) );
  INV_X1 U9597 ( .A(n14324), .ZN(n7138) );
  INV_X1 U9598 ( .A(n7139), .ZN(n15325) );
  NAND2_X1 U9599 ( .A1(n7145), .A2(n14333), .ZN(n7144) );
  OR2_X1 U9600 ( .A1(n7149), .A2(n7152), .ZN(n7145) );
  INV_X1 U9601 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7159) );
  INV_X1 U9602 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7160) );
  MUX2_X1 U9603 ( .A(n12963), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  MUX2_X1 U9604 ( .A(P3_IR_REG_0__SCAN_IN), .B(n12963), .S(n9048), .Z(n10802)
         );
  MUX2_X1 U9605 ( .A(n15033), .B(n14869), .S(n10416), .Z(n14872) );
  NAND2_X1 U9606 ( .A1(n13265), .A2(n7178), .ZN(n13264) );
  INV_X1 U9607 ( .A(n7179), .ZN(n7178) );
  NAND2_X1 U9608 ( .A1(n13266), .A2(n13267), .ZN(n7179) );
  NAND2_X1 U9609 ( .A1(n13429), .A2(n7193), .ZN(n8020) );
  NAND2_X1 U9610 ( .A1(n7194), .A2(n8226), .ZN(n10351) );
  NAND2_X1 U9611 ( .A1(n10649), .A2(n10650), .ZN(n7194) );
  OAI21_X1 U9612 ( .B1(n10650), .B2(n10649), .A(n7194), .ZN(n10651) );
  INV_X1 U9613 ( .A(n8232), .ZN(n10990) );
  NAND2_X1 U9614 ( .A1(n7195), .A2(n7196), .ZN(n8235) );
  NAND2_X1 U9615 ( .A1(n8232), .A2(n8233), .ZN(n7195) );
  AND2_X1 U9616 ( .A1(n7197), .A2(n12116), .ZN(n7196) );
  OAI21_X2 U9617 ( .B1(n13384), .B2(n13392), .A(n8249), .ZN(n13370) );
  OAI21_X1 U9618 ( .B1(n13354), .B2(n7217), .A(n7215), .ZN(n13328) );
  NAND2_X1 U9619 ( .A1(n7656), .A2(n7655), .ZN(n8039) );
  NAND2_X1 U9620 ( .A1(n7365), .A2(n7364), .ZN(n7874) );
  NAND2_X1 U9621 ( .A1(n13450), .A2(n8246), .ZN(n13437) );
  NAND2_X1 U9622 ( .A1(n10766), .A2(n12108), .ZN(n10765) );
  NAND2_X1 U9623 ( .A1(n11028), .A2(n11027), .ZN(n11026) );
  NOR2_X1 U9624 ( .A1(n7228), .A2(n13901), .ZN(n14076) );
  OAI21_X1 U9625 ( .B1(n7228), .B2(n13901), .A(n7226), .ZN(n7225) );
  OAI21_X1 U9626 ( .B1(n7230), .B2(n7229), .A(n14637), .ZN(n7228) );
  INV_X1 U9627 ( .A(n12382), .ZN(n7229) );
  NAND2_X1 U9628 ( .A1(n8927), .A2(n6570), .ZN(n7231) );
  NAND2_X1 U9629 ( .A1(n7231), .A2(n7232), .ZN(n9158) );
  NAND2_X1 U9630 ( .A1(n9224), .A2(n7242), .ZN(n7241) );
  NAND2_X1 U9631 ( .A1(n7241), .A2(n7244), .ZN(n9004) );
  NOR2_X1 U9632 ( .A1(n12398), .A2(n12400), .ZN(n12397) );
  NAND2_X1 U9633 ( .A1(n7263), .A2(n7261), .ZN(n11729) );
  NAND2_X1 U9634 ( .A1(n7570), .A2(n12350), .ZN(n14024) );
  INV_X1 U9635 ( .A(n14452), .ZN(n12664) );
  NAND2_X1 U9636 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), 
        .ZN(n7272) );
  NAND2_X1 U9637 ( .A1(n10945), .A2(n10744), .ZN(n7275) );
  NAND4_X1 U9638 ( .A1(n7318), .A2(n7278), .A3(n8293), .A4(n7276), .ZN(n8301)
         );
  NAND2_X1 U9639 ( .A1(n7282), .A2(n12484), .ZN(n12182) );
  OAI211_X1 U9640 ( .C1(n12525), .C2(n7290), .A(n7288), .B(n7285), .ZN(n12202)
         );
  NAND2_X1 U9641 ( .A1(n12525), .A2(n7286), .ZN(n7285) );
  NOR2_X1 U9642 ( .A1(n7287), .A2(n12195), .ZN(n7286) );
  OAI21_X1 U9643 ( .B1(n12195), .B2(n7291), .A(n7289), .ZN(n7288) );
  OAI21_X1 U9644 ( .B1(n12195), .B2(n12434), .A(n7291), .ZN(n7289) );
  NAND2_X1 U9645 ( .A1(n12195), .A2(n12434), .ZN(n7290) );
  INV_X1 U9646 ( .A(n7312), .ZN(n10809) );
  NAND3_X1 U9647 ( .A1(n6431), .A2(n9061), .A3(n8895), .ZN(n9196) );
  NAND4_X1 U9648 ( .A1(n8286), .A2(n8284), .A3(n8285), .A4(n8540), .ZN(n8287)
         );
  NAND2_X1 U9649 ( .A1(n8360), .A2(n8283), .ZN(n8374) );
  NAND2_X1 U9650 ( .A1(n7332), .A2(n6578), .ZN(n11481) );
  NAND2_X1 U9651 ( .A1(n11147), .A2(n11323), .ZN(n7332) );
  OAI21_X1 U9652 ( .B1(n13936), .B2(n12377), .A(n12378), .ZN(n13927) );
  NAND3_X1 U9653 ( .A1(n8294), .A2(n6755), .A3(n7345), .ZN(n7344) );
  OR2_X2 U9654 ( .A1(n8304), .A2(n8589), .ZN(n8303) );
  NAND3_X1 U9655 ( .A1(n7579), .A2(n7578), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n7346) );
  NAND2_X1 U9656 ( .A1(n7595), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7347) );
  NAND2_X1 U9657 ( .A1(n7350), .A2(n7348), .ZN(n7604) );
  INV_X1 U9658 ( .A(n7349), .ZN(n7348) );
  NAND2_X1 U9659 ( .A1(n7599), .A2(n7353), .ZN(n7350) );
  NAND2_X1 U9660 ( .A1(n7837), .A2(n7367), .ZN(n7365) );
  NAND3_X1 U9661 ( .A1(n8706), .A2(n8705), .A3(n7381), .ZN(n7383) );
  INV_X1 U9662 ( .A(n8719), .ZN(n7382) );
  NAND2_X1 U9663 ( .A1(n7383), .A2(n7384), .ZN(n8735) );
  NAND2_X1 U9664 ( .A1(n8675), .A2(n9834), .ZN(n8676) );
  NAND3_X1 U9665 ( .A1(n7390), .A2(n12083), .A3(n7389), .ZN(n7388) );
  INV_X1 U9666 ( .A(n12070), .ZN(n7390) );
  NAND2_X1 U9667 ( .A1(n12077), .A2(n12083), .ZN(n7391) );
  NOR2_X1 U9668 ( .A1(n12077), .A2(n12065), .ZN(n7393) );
  NAND2_X1 U9669 ( .A1(n12048), .A2(n12047), .ZN(n7395) );
  NAND2_X1 U9670 ( .A1(n12038), .A2(n7402), .ZN(n7405) );
  INV_X1 U9671 ( .A(n11962), .ZN(n7407) );
  NAND2_X1 U9672 ( .A1(n7410), .A2(n7409), .ZN(n11910) );
  NAND2_X1 U9673 ( .A1(n11903), .A2(n7412), .ZN(n7409) );
  INV_X1 U9674 ( .A(n12025), .ZN(n7417) );
  INV_X1 U9675 ( .A(n12024), .ZN(n7418) );
  OAI22_X1 U9676 ( .A1(n11916), .A2(n7419), .B1(n11915), .B2(n11914), .ZN(
        n11924) );
  NAND2_X1 U9677 ( .A1(n11924), .A2(n11925), .ZN(n11923) );
  NAND3_X1 U9678 ( .A1(n11929), .A2(n11928), .A3(n6581), .ZN(n7422) );
  NAND3_X1 U9679 ( .A1(n7679), .A2(n7425), .A3(n7424), .ZN(n7859) );
  NAND2_X1 U9680 ( .A1(n7428), .A2(n9675), .ZN(n10173) );
  NAND3_X1 U9681 ( .A1(n10030), .A2(n9674), .A3(n9669), .ZN(n7428) );
  NAND2_X1 U9682 ( .A1(n9782), .A2(n7430), .ZN(n7429) );
  OAI211_X1 U9683 ( .C1(n9782), .C2(n7431), .A(n12998), .B(n7429), .ZN(
        P2_U3192) );
  NAND2_X1 U9684 ( .A1(n13103), .A2(n7555), .ZN(n13015) );
  INV_X1 U9685 ( .A(n7449), .ZN(n13014) );
  INV_X1 U9686 ( .A(n13016), .ZN(n7450) );
  NAND2_X1 U9687 ( .A1(n7452), .A2(n7454), .ZN(n7451) );
  INV_X1 U9688 ( .A(n10172), .ZN(n7452) );
  INV_X1 U9689 ( .A(n7454), .ZN(n7453) );
  NAND2_X1 U9690 ( .A1(n6470), .A2(n10172), .ZN(n7456) );
  NAND2_X1 U9691 ( .A1(n10172), .A2(n9682), .ZN(n10262) );
  INV_X1 U9692 ( .A(n9683), .ZN(n7458) );
  INV_X1 U9693 ( .A(n9684), .ZN(n7459) );
  INV_X1 U9694 ( .A(n9682), .ZN(n7460) );
  NOR2_X1 U9695 ( .A1(n13036), .A2(n9771), .ZN(n13009) );
  NAND2_X2 U9696 ( .A1(n9385), .A2(n9384), .ZN(n9048) );
  NAND2_X1 U9697 ( .A1(n11434), .A2(n7475), .ZN(n7472) );
  NAND2_X1 U9698 ( .A1(n7472), .A2(n7473), .ZN(n11670) );
  NAND2_X1 U9699 ( .A1(n12687), .A2(n7485), .ZN(n7481) );
  NAND2_X1 U9700 ( .A1(n7481), .A2(n7482), .ZN(n9655) );
  INV_X1 U9701 ( .A(n12695), .ZN(n7493) );
  AND2_X2 U9702 ( .A1(n8899), .A2(n7502), .ZN(n7501) );
  AOI21_X1 U9703 ( .B1(n12792), .B2(n7506), .A(n7503), .ZN(n12756) );
  OAI211_X1 U9704 ( .C1(n13775), .C2(n6587), .A(n7511), .B(n7509), .ZN(n12345)
         );
  NAND2_X1 U9705 ( .A1(n13775), .A2(n7510), .ZN(n7509) );
  NOR2_X1 U9706 ( .A1(n7513), .A2(n12338), .ZN(n7510) );
  OAI22_X1 U9707 ( .A1(n7513), .A2(n7512), .B1(n12338), .B2(n7515), .ZN(n7511)
         );
  NOR2_X1 U9708 ( .A1(n12338), .A2(n13657), .ZN(n7512) );
  INV_X1 U9709 ( .A(n12338), .ZN(n7514) );
  NOR2_X1 U9710 ( .A1(n11403), .A2(n7528), .ZN(n7527) );
  OAI21_X2 U9711 ( .B1(n14506), .B2(n7531), .A(n7529), .ZN(n13749) );
  NOR2_X1 U9712 ( .A1(n8456), .A2(n8287), .ZN(n8562) );
  AOI21_X1 U9713 ( .B1(n12943), .B2(n6437), .A(n9484), .ZN(n9486) );
  NAND2_X1 U9714 ( .A1(n9004), .A2(n9002), .ZN(n8943) );
  AOI21_X1 U9715 ( .B1(n8187), .B2(n13430), .A(n8186), .ZN(n8278) );
  OAI21_X1 U9716 ( .B1(n8278), .B2(n13428), .A(n8277), .ZN(n8279) );
  INV_X1 U9717 ( .A(n8051), .ZN(n8053) );
  INV_X1 U9718 ( .A(n12080), .ZN(n12081) );
  OAI22_X1 U9719 ( .A1(n9664), .A2(n13620), .B1(n14859), .B2(n9663), .ZN(n9665) );
  OAI22_X1 U9720 ( .A1(n9664), .A2(n13561), .B1(n13552), .B2(n8262), .ZN(n8263) );
  NAND2_X1 U9721 ( .A1(n8766), .A2(n8765), .ZN(n8767) );
  NOR2_X1 U9722 ( .A1(n11974), .A2(n11973), .ZN(n12011) );
  NOR2_X1 U9723 ( .A1(n12019), .A2(n12018), .ZN(n12022) );
  AOI21_X1 U9724 ( .B1(n12017), .B2(n12016), .A(n12015), .ZN(n12019) );
  INV_X1 U9725 ( .A(n8178), .ZN(n12138) );
  OR2_X1 U9726 ( .A1(n8779), .A2(n10681), .ZN(n8331) );
  NAND2_X1 U9727 ( .A1(n13564), .A2(n12085), .ZN(n12056) );
  OAI211_X2 U9728 ( .C1(n8359), .C2(n9832), .A(n8346), .B(n8345), .ZN(n10689)
         );
  NAND2_X1 U9729 ( .A1(n13813), .A2(n12319), .ZN(n10287) );
  NAND2_X1 U9730 ( .A1(n10923), .A2(n13813), .ZN(n10284) );
  AND4_X2 U9731 ( .A1(n8358), .A2(n8357), .A3(n8356), .A4(n8355), .ZN(n8827)
         );
  NAND2_X1 U9732 ( .A1(n8877), .A2(n8869), .ZN(n8879) );
  NAND2_X1 U9733 ( .A1(n9782), .A2(n9783), .ZN(n9790) );
  INV_X2 U9734 ( .A(n8788), .ZN(n8369) );
  INV_X1 U9735 ( .A(n8909), .ZN(n12950) );
  INV_X1 U9736 ( .A(n9060), .ZN(n9280) );
  NAND2_X1 U9737 ( .A1(n9060), .A2(n9034), .ZN(n9035) );
  OR2_X1 U9738 ( .A1(n9416), .A2(n9225), .ZN(n9417) );
  NOR2_X1 U9739 ( .A1(n12070), .A2(n12061), .ZN(n12077) );
  XNOR2_X1 U9740 ( .A(n10360), .B(n10362), .ZN(n14573) );
  AOI22_X1 U9741 ( .A1(n12333), .A2(n14623), .B1(n10285), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n10286) );
  AOI22_X1 U9742 ( .A1(n12319), .A2(n14623), .B1(n14207), .B2(n10285), .ZN(
        n10283) );
  OR2_X1 U9743 ( .A1(n8826), .A2(n8800), .ZN(n7544) );
  NOR2_X1 U9744 ( .A1(n11371), .A2(n11366), .ZN(n7545) );
  NOR2_X1 U9745 ( .A1(n10882), .A2(n15136), .ZN(n12801) );
  NAND2_X1 U9746 ( .A1(n10729), .A2(n15081), .ZN(n15096) );
  OR2_X1 U9747 ( .A1(n9466), .A2(n12894), .ZN(n7547) );
  AND2_X1 U9748 ( .A1(n10516), .A2(n10504), .ZN(n7548) );
  AND2_X1 U9749 ( .A1(n7624), .A2(n7623), .ZN(n7549) );
  INV_X1 U9750 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7692) );
  AND4_X1 U9751 ( .A1(n7686), .A2(n8188), .A3(n8191), .A4(n8216), .ZN(n7550)
         );
  OR2_X1 U9752 ( .A1(n12493), .A2(n12702), .ZN(n7551) );
  XOR2_X1 U9753 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n7552) );
  AND2_X1 U9754 ( .A1(n9761), .A2(n9760), .ZN(n7553) );
  AND2_X1 U9755 ( .A1(n11841), .A2(n11840), .ZN(n7554) );
  OR2_X1 U9756 ( .A1(n11116), .A2(n11115), .ZN(n7557) );
  AND2_X1 U9757 ( .A1(n11798), .A2(n12547), .ZN(n7559) );
  NOR2_X1 U9758 ( .A1(n15141), .A2(n9450), .ZN(n7560) );
  OR2_X1 U9759 ( .A1(n7585), .A2(n9836), .ZN(n7561) );
  AND2_X1 U9760 ( .A1(n10927), .A2(n10926), .ZN(n7562) );
  INV_X1 U9761 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8589) );
  NAND2_X1 U9762 ( .A1(n9795), .A2(n9788), .ZN(n13070) );
  INV_X1 U9763 ( .A(n13070), .ZN(n9789) );
  AND2_X1 U9764 ( .A1(n7628), .A2(n7627), .ZN(n7563) );
  OR2_X1 U9765 ( .A1(n14551), .A2(n14550), .ZN(n7564) );
  INV_X1 U9766 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8288) );
  INV_X1 U9767 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8466) );
  AND2_X1 U9768 ( .A1(n7641), .A2(n7640), .ZN(n7565) );
  INV_X1 U9769 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14280) );
  INV_X1 U9770 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14255) );
  INV_X1 U9771 ( .A(n9052), .ZN(n8964) );
  INV_X1 U9772 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7642) );
  INV_X1 U9773 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8437) );
  INV_X1 U9774 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7577) );
  INV_X1 U9775 ( .A(n12367), .ZN(n12350) );
  NOR2_X1 U9776 ( .A1(n8520), .A2(n8532), .ZN(n7566) );
  AND2_X1 U9777 ( .A1(n11865), .A2(n11864), .ZN(n7568) );
  AND2_X1 U9778 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7569) );
  OR2_X1 U9779 ( .A1(n12427), .A2(n14458), .ZN(n7571) );
  AND2_X1 U9780 ( .A1(n12682), .A2(n12690), .ZN(n7572) );
  INV_X1 U9781 ( .A(n13468), .ZN(n13428) );
  INV_X1 U9782 ( .A(n11046), .ZN(n9147) );
  AND3_X1 U9783 ( .A1(n9289), .A2(n9288), .A3(n9287), .ZN(n12796) );
  INV_X1 U9784 ( .A(n12796), .ZN(n9290) );
  INV_X1 U9785 ( .A(n12773), .ZN(n9406) );
  OR2_X1 U9786 ( .A1(n7646), .A2(SI_17_), .ZN(n7575) );
  AND2_X1 U9787 ( .A1(n8365), .A2(n10694), .ZN(n8366) );
  NAND2_X1 U9788 ( .A1(n11897), .A2(n11896), .ZN(n11903) );
  INV_X1 U9789 ( .A(n11908), .ZN(n11909) );
  NAND2_X1 U9790 ( .A1(n11938), .A2(n11937), .ZN(n11942) );
  INV_X1 U9791 ( .A(n11942), .ZN(n11943) );
  INV_X1 U9792 ( .A(n11949), .ZN(n11950) );
  NAND2_X1 U9793 ( .A1(n11952), .A2(n11951), .ZN(n11958) );
  OAI21_X1 U9794 ( .B1(n12059), .B2(n11955), .A(n11954), .ZN(n11956) );
  NAND2_X1 U9795 ( .A1(n11983), .A2(n11982), .ZN(n11999) );
  AOI21_X1 U9796 ( .B1(n12011), .B2(n12010), .A(n12009), .ZN(n12014) );
  NAND2_X1 U9797 ( .A1(n12019), .A2(n12018), .ZN(n12020) );
  AOI22_X1 U9798 ( .A1(n13587), .A2(n11863), .B1(n12085), .B2(n13121), .ZN(
        n12034) );
  XNOR2_X1 U9799 ( .A(n12422), .B(n12412), .ZN(n12070) );
  OR4_X1 U9800 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_22__SCAN_IN), .ZN(n9432) );
  INV_X1 U9801 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8901) );
  INV_X1 U9802 ( .A(SI_12_), .ZN(n9198) );
  INV_X1 U9803 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9215) );
  INV_X1 U9804 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n11642) );
  NAND2_X1 U9805 ( .A1(n8889), .A2(n8888), .ZN(n9306) );
  AND2_X1 U9806 ( .A1(n9267), .A2(n9266), .ZN(n9284) );
  AND2_X1 U9807 ( .A1(n9232), .A2(n11642), .ZN(n9247) );
  AND2_X1 U9808 ( .A1(n8901), .A2(n8957), .ZN(n8902) );
  INV_X1 U9809 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n8935) );
  INV_X1 U9810 ( .A(n8011), .ZN(n8009) );
  INV_X1 U9811 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7899) );
  AOI22_X1 U9812 ( .A1(n13117), .A2(n13050), .B1(n12411), .B2(n13116), .ZN(
        n8185) );
  OR2_X1 U9813 ( .A1(n8120), .A2(n8119), .ZN(n8133) );
  INV_X1 U9814 ( .A(n8044), .ZN(n8042) );
  AND2_X1 U9815 ( .A1(n8722), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8737) );
  INV_X1 U9816 ( .A(n13943), .ZN(n12358) );
  INV_X1 U9817 ( .A(n14008), .ZN(n12352) );
  INV_X1 U9818 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8294) );
  INV_X1 U9819 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8869) );
  OR2_X1 U9820 ( .A1(n8963), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9343) );
  INV_X1 U9821 ( .A(n10485), .ZN(n10486) );
  NOR2_X1 U9822 ( .A1(n9328), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8961) );
  AND2_X1 U9823 ( .A1(n11543), .A2(n12548), .ZN(n11541) );
  AND2_X1 U9824 ( .A1(n9453), .A2(n9444), .ZN(n10492) );
  OR2_X1 U9825 ( .A1(n9306), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9319) );
  INV_X1 U9826 ( .A(n12952), .ZN(n8910) );
  OR2_X1 U9827 ( .A1(n9178), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9202) );
  INV_X1 U9828 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9450) );
  AND2_X1 U9829 ( .A1(n9926), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8932) );
  OR2_X1 U9830 ( .A1(n9778), .A2(n9777), .ZN(n9779) );
  INV_X1 U9831 ( .A(n11129), .ZN(n9709) );
  NAND2_X1 U9832 ( .A1(n8009), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8028) );
  OR2_X1 U9833 ( .A1(n8106), .A2(n13041), .ZN(n8120) );
  OR2_X1 U9834 ( .A1(n8028), .A2(n8027), .ZN(n8044) );
  OR2_X1 U9835 ( .A1(n10079), .A2(n10078), .ZN(n10129) );
  NAND2_X1 U9836 ( .A1(n8091), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8106) );
  AND2_X1 U9837 ( .A1(n15339), .A2(n8188), .ZN(n8194) );
  AND3_X1 U9838 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n8420) );
  NOR2_X1 U9839 ( .A1(n8641), .A2(n8640), .ZN(n8652) );
  AND2_X1 U9840 ( .A1(n8739), .A2(n8725), .ZN(n13924) );
  NAND2_X1 U9841 ( .A1(n7220), .A2(n12358), .ZN(n12359) );
  AND2_X1 U9842 ( .A1(n8652), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8666) );
  INV_X1 U9843 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8875) );
  NOR2_X1 U9844 ( .A1(n14282), .A2(n14283), .ZN(n14227) );
  INV_X1 U9845 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14307) );
  NAND2_X1 U9846 ( .A1(n12560), .A2(n10802), .ZN(n10906) );
  NAND2_X1 U9847 ( .A1(n9151), .A2(n9150), .ZN(n9163) );
  NAND2_X1 U9848 ( .A1(n11342), .A2(n12549), .ZN(n11343) );
  OR2_X1 U9849 ( .A1(n10389), .A2(n10388), .ZN(n12516) );
  AND2_X1 U9850 ( .A1(n9424), .A2(n9420), .ZN(n9809) );
  AND2_X1 U9851 ( .A1(n10400), .A2(n10399), .ZN(n10415) );
  INV_X1 U9852 ( .A(n9514), .ZN(n9373) );
  NOR2_X1 U9853 ( .A1(n9202), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9216) );
  OR2_X1 U9854 ( .A1(n9098), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9113) );
  AND2_X1 U9855 ( .A1(n9887), .A2(n10479), .ZN(n9453) );
  NOR2_X1 U9856 ( .A1(n9437), .A2(n9436), .ZN(n9454) );
  OR2_X1 U9857 ( .A1(n6440), .A2(n11110), .ZN(n9317) );
  NOR2_X1 U9858 ( .A1(n9441), .A2(n10479), .ZN(n10391) );
  INV_X1 U9859 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9225) );
  OR2_X1 U9860 ( .A1(n8058), .A2(n13003), .ZN(n8074) );
  INV_X1 U9861 ( .A(n13110), .ZN(n13097) );
  AND2_X1 U9862 ( .A1(n8171), .A2(n8162), .ZN(n13263) );
  INV_X1 U9863 ( .A(n8150), .ZN(n8175) );
  INV_X1 U9864 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10315) );
  OR2_X1 U9865 ( .A1(n9901), .A2(n12145), .ZN(n14750) );
  INV_X1 U9866 ( .A(n13050), .ZN(n13092) );
  NAND2_X1 U9867 ( .A1(n7750), .A2(n8342), .ZN(n7728) );
  INV_X1 U9868 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7706) );
  NOR2_X1 U9869 ( .A1(n8518), .A2(n8306), .ZN(n8532) );
  AND2_X1 U9870 ( .A1(n12311), .A2(n12309), .ZN(n13695) );
  NOR2_X1 U9871 ( .A1(n15165), .A2(n8679), .ZN(n8678) );
  AND2_X1 U9872 ( .A1(n8750), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8770) );
  AND4_X1 U9873 ( .A1(n8622), .A2(n8621), .A3(n8620), .A4(n8619), .ZN(n13681)
         );
  AOI21_X1 U9874 ( .B1(n12403), .B2(n14138), .A(n12402), .ZN(n12404) );
  AND2_X1 U9875 ( .A1(n8823), .A2(n12366), .ZN(n14036) );
  INV_X1 U9876 ( .A(n13813), .ZN(n14627) );
  XNOR2_X1 U9877 ( .A(n14087), .B(n13801), .ZN(n12400) );
  INV_X1 U9878 ( .A(n14339), .ZN(n14622) );
  INV_X1 U9879 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14274) );
  OAI21_X1 U9880 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n14239), .A(n14238), .ZN(
        n14302) );
  INV_X1 U9881 ( .A(n11571), .ZN(n11348) );
  INV_X1 U9882 ( .A(n12508), .ZN(n12530) );
  OAI22_X1 U9883 ( .A1(n11713), .A2(n11712), .B1(n11751), .B2(n11711), .ZN(
        n11800) );
  AND2_X1 U9884 ( .A1(n9350), .A2(n9349), .ZN(n12690) );
  AND4_X1 U9885 ( .A1(n9253), .A2(n9252), .A3(n9251), .A4(n9250), .ZN(n12828)
         );
  INV_X1 U9886 ( .A(n15018), .ZN(n15037) );
  INV_X1 U9887 ( .A(n12596), .ZN(n12659) );
  INV_X1 U9888 ( .A(n15084), .ZN(n14435) );
  INV_X1 U9889 ( .A(n15081), .ZN(n15071) );
  INV_X1 U9890 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9465) );
  NOR3_X1 U9891 ( .A1(n10396), .A2(n9454), .A3(n9453), .ZN(n10722) );
  INV_X1 U9892 ( .A(n15137), .ZN(n15133) );
  NAND2_X1 U9893 ( .A1(n9457), .A2(n10714), .ZN(n15136) );
  NAND2_X1 U9894 ( .A1(n9440), .A2(n9439), .ZN(n10479) );
  XNOR2_X1 U9895 ( .A(n9415), .B(n9414), .ZN(n10397) );
  INV_X1 U9896 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9382) );
  AND2_X1 U9897 ( .A1(n9831), .A2(P3_U3151), .ZN(n14319) );
  INV_X1 U9898 ( .A(n13320), .ZN(n13505) );
  AND2_X1 U9899 ( .A1(n8155), .A2(n8154), .ZN(n13095) );
  AND2_X1 U9900 ( .A1(n9908), .A2(n9900), .ZN(n14818) );
  NAND2_X1 U9901 ( .A1(n8177), .A2(n8176), .ZN(n13430) );
  INV_X1 U9902 ( .A(n13463), .ZN(n13476) );
  INV_X1 U9903 ( .A(n14853), .ZN(n14845) );
  INV_X1 U9904 ( .A(n14831), .ZN(n9784) );
  AND2_X1 U9905 ( .A1(n11742), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8218) );
  NAND2_X1 U9906 ( .A1(n10279), .A2(n14608), .ZN(n14564) );
  AND2_X1 U9907 ( .A1(n8692), .A2(n8709), .ZN(n13967) );
  OR2_X1 U9908 ( .A1(n8484), .A2(n10214), .ZN(n8518) );
  AND4_X1 U9909 ( .A1(n8731), .A2(n8730), .A3(n8729), .A4(n8728), .ZN(n13701)
         );
  INV_X1 U9910 ( .A(n13681), .ZN(n14038) );
  AND4_X1 U9911 ( .A1(n8598), .A2(n8597), .A3(n8596), .A4(n8595), .ZN(n8824)
         );
  INV_X1 U9912 ( .A(n14591), .ZN(n11701) );
  INV_X1 U9913 ( .A(n14596), .ZN(n13887) );
  INV_X1 U9914 ( .A(n14058), .ZN(n14637) );
  INV_X1 U9915 ( .A(n12380), .ZN(n12361) );
  INV_X1 U9916 ( .A(n12377), .ZN(n13939) );
  INV_X1 U9917 ( .A(n11727), .ZN(n11719) );
  NAND2_X1 U9918 ( .A1(n10250), .A2(n10249), .ZN(n14138) );
  INV_X1 U9919 ( .A(n14639), .ZN(n14060) );
  NAND2_X1 U9920 ( .A1(n12386), .A2(n14608), .ZN(n14610) );
  AND2_X1 U9921 ( .A1(n10672), .A2(n10289), .ZN(n10736) );
  AND2_X1 U9922 ( .A1(n14631), .A2(n14743), .ZN(n14153) );
  INV_X1 U9923 ( .A(n14153), .ZN(n14729) );
  NOR2_X1 U9924 ( .A1(n10673), .A2(n10930), .ZN(n10735) );
  INV_X1 U9925 ( .A(n10272), .ZN(n10321) );
  INV_X1 U9926 ( .A(n8322), .ZN(n8323) );
  AND2_X1 U9927 ( .A1(n8414), .A2(n8444), .ZN(n10055) );
  AND2_X1 U9928 ( .A1(n10401), .A2(n10400), .ZN(n15030) );
  INV_X1 U9929 ( .A(n12839), .ZN(n12682) );
  INV_X1 U9930 ( .A(n12505), .ZN(n12532) );
  INV_X1 U9931 ( .A(n12521), .ZN(n12538) );
  INV_X1 U9932 ( .A(n12690), .ZN(n12541) );
  INV_X1 U9933 ( .A(n12813), .ZN(n12544) );
  INV_X1 U9934 ( .A(n14992), .ZN(n15033) );
  OR2_X1 U9935 ( .A1(n12559), .A2(n10402), .ZN(n15018) );
  INV_X1 U9936 ( .A(n15030), .ZN(n14996) );
  INV_X1 U9937 ( .A(n14866), .ZN(n15043) );
  AND2_X1 U9938 ( .A1(n12785), .A2(n12784), .ZN(n12872) );
  NAND2_X1 U9939 ( .A1(n10913), .A2(n15096), .ZN(n12805) );
  INV_X1 U9940 ( .A(n12801), .ZN(n12835) );
  NAND2_X1 U9941 ( .A1(n15157), .A2(n15078), .ZN(n12894) );
  AND2_X2 U9942 ( .A1(n10722), .A2(n9463), .ZN(n15157) );
  NAND2_X1 U9943 ( .A1(n9464), .A2(n15141), .ZN(n9452) );
  INV_X1 U9944 ( .A(n12455), .ZN(n12922) );
  AND2_X1 U9945 ( .A1(n9190), .A2(n9189), .ZN(n11571) );
  INV_X2 U9946 ( .A(n15142), .ZN(n15141) );
  CLKBUF_X1 U9947 ( .A(n9975), .Z(n10001) );
  INV_X1 U9948 ( .A(n12960), .ZN(n14320) );
  INV_X1 U9949 ( .A(SI_18_), .ZN(n10370) );
  INV_X1 U9950 ( .A(SI_13_), .ZN(n9957) );
  INV_X1 U9951 ( .A(n14791), .ZN(n14812) );
  INV_X1 U9952 ( .A(n11907), .ZN(n10707) );
  INV_X1 U9953 ( .A(n13477), .ZN(n11242) );
  NAND2_X1 U9954 ( .A1(n8168), .A2(n8167), .ZN(n13117) );
  INV_X1 U9955 ( .A(n13059), .ZN(n13123) );
  INV_X1 U9956 ( .A(n11967), .ZN(n13129) );
  INV_X1 U9957 ( .A(n14818), .ZN(n14769) );
  OR2_X1 U9958 ( .A1(n9908), .A2(P2_U3088), .ZN(n14791) );
  INV_X1 U9959 ( .A(n13470), .ZN(n13467) );
  INV_X1 U9960 ( .A(n13331), .ZN(n13584) );
  NAND2_X1 U9961 ( .A1(n14859), .A2(n14845), .ZN(n13602) );
  NAND2_X1 U9962 ( .A1(n14859), .A2(n14850), .ZN(n13620) );
  NOR2_X1 U9963 ( .A1(n14832), .A2(n14827), .ZN(n14828) );
  INV_X1 U9964 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13633) );
  INV_X1 U9965 ( .A(n12149), .ZN(n12089) );
  INV_X1 U9966 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10036) );
  INV_X1 U9967 ( .A(n11616), .ZN(n11851) );
  INV_X1 U9968 ( .A(n14343), .ZN(n14526) );
  INV_X1 U9969 ( .A(n13739), .ZN(n14577) );
  INV_X1 U9970 ( .A(n13779), .ZN(n13959) );
  INV_X1 U9971 ( .A(n11833), .ZN(n13804) );
  OR2_X1 U9972 ( .A1(n10150), .A2(n10252), .ZN(n14601) );
  INV_X1 U9973 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14606) );
  INV_X1 U9974 ( .A(n14045), .ZN(n14351) );
  NAND2_X1 U9975 ( .A1(n14610), .A2(n10676), .ZN(n14352) );
  INV_X2 U9976 ( .A(n14610), .ZN(n14646) );
  INV_X1 U9977 ( .A(n14748), .ZN(n14746) );
  INV_X1 U9978 ( .A(n15160), .ZN(n15158) );
  NOR2_X2 U9979 ( .A1(n10322), .A2(n10321), .ZN(n14660) );
  CLKBUF_X1 U9980 ( .A(n14660), .Z(n14673) );
  INV_X1 U9981 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9967) );
  INV_X1 U9982 ( .A(n12559), .ZN(P3_U3897) );
  NAND2_X1 U9983 ( .A1(n9452), .A2(n9451), .ZN(P3_U3456) );
  INV_X1 U9984 ( .A(n13132), .ZN(P2_U3947) );
  NAND2_X1 U9985 ( .A1(n8281), .A2(n8280), .ZN(P2_U3236) );
  NOR2_X1 U9986 ( .A1(n10282), .A2(n10323), .ZN(P1_U4016) );
  INV_X1 U9987 ( .A(n9046), .ZN(n7581) );
  NAND2_X1 U9988 ( .A1(n7581), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7735) );
  AND2_X1 U9989 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n7582) );
  NAND2_X1 U9990 ( .A1(n9031), .A2(n7582), .ZN(n8337) );
  NAND2_X1 U9991 ( .A1(n7735), .A2(n8337), .ZN(n7726) );
  NAND2_X1 U9992 ( .A1(n7583), .A2(n7726), .ZN(n7586) );
  INV_X1 U9993 ( .A(n7584), .ZN(n7585) );
  INV_X1 U9994 ( .A(SI_1_), .ZN(n9836) );
  NAND2_X1 U9995 ( .A1(n7586), .A2(n7561), .ZN(n7747) );
  INV_X1 U9996 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9866) );
  MUX2_X1 U9997 ( .A(n9848), .B(n9866), .S(n7595), .Z(n7587) );
  XNOR2_X1 U9998 ( .A(n7587), .B(SI_2_), .ZN(n7748) );
  NAND2_X1 U9999 ( .A1(n7747), .A2(n7748), .ZN(n7590) );
  INV_X1 U10000 ( .A(n7587), .ZN(n7588) );
  NAND2_X1 U10001 ( .A1(n7588), .A2(SI_2_), .ZN(n7589) );
  MUX2_X1 U10002 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n7595), .Z(n7592) );
  XNOR2_X1 U10003 ( .A(n7592), .B(SI_3_), .ZN(n7762) );
  INV_X1 U10004 ( .A(n7762), .ZN(n7591) );
  NAND2_X1 U10005 ( .A1(n7592), .A2(SI_3_), .ZN(n7593) );
  NAND2_X1 U10006 ( .A1(n7597), .A2(SI_4_), .ZN(n7598) );
  NAND2_X1 U10007 ( .A1(n7602), .A2(SI_6_), .ZN(n7603) );
  NAND2_X1 U10008 ( .A1(n7604), .A2(n7603), .ZN(n7816) );
  MUX2_X1 U10009 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9831), .Z(n7606) );
  XNOR2_X1 U10010 ( .A(n7606), .B(SI_7_), .ZN(n7815) );
  INV_X1 U10011 ( .A(n7815), .ZN(n7605) );
  NAND2_X1 U10012 ( .A1(n7816), .A2(n7605), .ZN(n7608) );
  NAND2_X1 U10013 ( .A1(n7606), .A2(SI_7_), .ZN(n7607) );
  MUX2_X1 U10014 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9831), .Z(n7610) );
  INV_X1 U10015 ( .A(n7836), .ZN(n7609) );
  NAND2_X1 U10016 ( .A1(n7610), .A2(SI_8_), .ZN(n7611) );
  MUX2_X1 U10017 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9831), .Z(n7612) );
  XNOR2_X1 U10018 ( .A(n7612), .B(SI_9_), .ZN(n7855) );
  MUX2_X1 U10019 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9831), .Z(n7614) );
  XNOR2_X1 U10020 ( .A(n7614), .B(SI_10_), .ZN(n7873) );
  INV_X1 U10021 ( .A(n7873), .ZN(n7613) );
  NAND2_X1 U10022 ( .A1(n7874), .A2(n7613), .ZN(n7616) );
  NAND2_X1 U10023 ( .A1(n7614), .A2(SI_10_), .ZN(n7615) );
  MUX2_X1 U10024 ( .A(n9959), .B(n15289), .S(n6439), .Z(n7617) );
  NAND2_X1 U10025 ( .A1(n7617), .A2(n9188), .ZN(n7620) );
  INV_X1 U10026 ( .A(n7617), .ZN(n7618) );
  NAND2_X1 U10027 ( .A1(n7618), .A2(SI_11_), .ZN(n7619) );
  NAND2_X1 U10028 ( .A1(n7620), .A2(n7619), .ZN(n7891) );
  MUX2_X1 U10029 ( .A(n9967), .B(n9963), .S(n9831), .Z(n7621) );
  NAND2_X1 U10030 ( .A1(n7621), .A2(n9198), .ZN(n7624) );
  INV_X1 U10031 ( .A(n7621), .ZN(n7622) );
  NAND2_X1 U10032 ( .A1(n7622), .A2(SI_12_), .ZN(n7623) );
  MUX2_X1 U10033 ( .A(n8935), .B(n10036), .S(n6439), .Z(n7625) );
  NAND2_X1 U10034 ( .A1(n7625), .A2(n9957), .ZN(n7628) );
  INV_X1 U10035 ( .A(n7625), .ZN(n7626) );
  NAND2_X1 U10036 ( .A1(n7626), .A2(SI_13_), .ZN(n7627) );
  MUX2_X1 U10037 ( .A(n8939), .B(n10259), .S(n6439), .Z(n7938) );
  INV_X1 U10038 ( .A(n7938), .ZN(n7629) );
  NAND2_X1 U10039 ( .A1(n7937), .A2(n7629), .ZN(n7633) );
  INV_X1 U10040 ( .A(n7630), .ZN(n7631) );
  NAND2_X1 U10041 ( .A1(n7631), .A2(SI_14_), .ZN(n7632) );
  MUX2_X1 U10042 ( .A(n10425), .B(n10424), .S(n9831), .Z(n7634) );
  INV_X1 U10043 ( .A(n7634), .ZN(n7635) );
  NAND2_X1 U10044 ( .A1(n7635), .A2(SI_15_), .ZN(n7636) );
  NAND2_X1 U10045 ( .A1(n7637), .A2(n7636), .ZN(n7960) );
  MUX2_X1 U10046 ( .A(n8941), .B(n10576), .S(n9831), .Z(n7638) );
  INV_X1 U10047 ( .A(n7638), .ZN(n7639) );
  NAND2_X1 U10048 ( .A1(n7639), .A2(SI_16_), .ZN(n7640) );
  MUX2_X1 U10049 ( .A(n7642), .B(n10587), .S(n6439), .Z(n7987) );
  AOI21_X1 U10050 ( .B1(n7646), .B2(SI_17_), .A(SI_18_), .ZN(n7643) );
  NAND2_X1 U10051 ( .A1(n7989), .A2(n7643), .ZN(n7648) );
  AOI21_X1 U10052 ( .B1(SI_17_), .B2(SI_18_), .A(n7987), .ZN(n7644) );
  NOR2_X1 U10053 ( .A1(SI_18_), .A2(SI_17_), .ZN(n7645) );
  INV_X1 U10054 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7649) );
  MUX2_X1 U10055 ( .A(n7649), .B(n6640), .S(n6439), .Z(n8002) );
  MUX2_X1 U10056 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9831), .Z(n7653) );
  NAND2_X1 U10057 ( .A1(n7654), .A2(n10583), .ZN(n7655) );
  MUX2_X1 U10058 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n9831), .Z(n8040) );
  MUX2_X1 U10059 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n6439), .Z(n7657) );
  NAND2_X1 U10060 ( .A1(n7657), .A2(SI_21_), .ZN(n7659) );
  OAI21_X1 U10061 ( .B1(SI_21_), .B2(n7657), .A(n7659), .ZN(n8052) );
  INV_X1 U10062 ( .A(n8052), .ZN(n7658) );
  MUX2_X1 U10063 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n6439), .Z(n8066) );
  MUX2_X1 U10064 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9831), .Z(n7661) );
  NAND2_X1 U10065 ( .A1(n7661), .A2(SI_23_), .ZN(n7663) );
  OAI21_X1 U10066 ( .B1(SI_23_), .B2(n7661), .A(n7663), .ZN(n8084) );
  INV_X1 U10067 ( .A(n8084), .ZN(n7662) );
  MUX2_X1 U10068 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n6439), .Z(n7664) );
  NAND2_X1 U10069 ( .A1(n7664), .A2(SI_24_), .ZN(n8113) );
  OAI21_X1 U10070 ( .B1(SI_24_), .B2(n7664), .A(n8113), .ZN(n8102) );
  INV_X1 U10071 ( .A(n8102), .ZN(n7665) );
  MUX2_X1 U10072 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n6439), .Z(n7668) );
  XNOR2_X1 U10073 ( .A(n7668), .B(SI_25_), .ZN(n8115) );
  INV_X1 U10074 ( .A(n8115), .ZN(n7666) );
  AND2_X1 U10075 ( .A1(n7666), .A2(n8113), .ZN(n7667) );
  INV_X1 U10076 ( .A(n7668), .ZN(n7669) );
  INV_X1 U10077 ( .A(SI_25_), .ZN(n11523) );
  INV_X1 U10078 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13643) );
  MUX2_X1 U10079 ( .A(n14200), .B(n13643), .S(n6439), .Z(n8127) );
  INV_X1 U10080 ( .A(n8127), .ZN(n7670) );
  NOR2_X1 U10081 ( .A1(n7670), .A2(SI_26_), .ZN(n7671) );
  OAI22_X1 U10082 ( .A1(n8129), .A2(n7671), .B1(n8127), .B2(n12961), .ZN(n8144) );
  INV_X1 U10083 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13641) );
  MUX2_X1 U10084 ( .A(n15193), .B(n13641), .S(n6439), .Z(n8141) );
  INV_X1 U10085 ( .A(SI_27_), .ZN(n12394) );
  NOR2_X1 U10086 ( .A1(n8141), .A2(n12394), .ZN(n7672) );
  NAND2_X1 U10087 ( .A1(n8141), .A2(n12394), .ZN(n7673) );
  INV_X1 U10088 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13638) );
  MUX2_X1 U10089 ( .A(n14194), .B(n13638), .S(n6439), .Z(n7674) );
  XNOR2_X1 U10090 ( .A(n7674), .B(SI_28_), .ZN(n8156) );
  NAND2_X1 U10091 ( .A1(n8157), .A2(n8156), .ZN(n7676) );
  INV_X1 U10092 ( .A(SI_28_), .ZN(n12957) );
  NAND2_X1 U10093 ( .A1(n7674), .A2(n12957), .ZN(n7675) );
  NAND2_X1 U10094 ( .A1(n7676), .A2(n7675), .ZN(n8792) );
  INV_X1 U10095 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7677) );
  MUX2_X1 U10096 ( .A(n7677), .B(n13633), .S(n9831), .Z(n8793) );
  XNOR2_X1 U10097 ( .A(n8793), .B(SI_29_), .ZN(n8791) );
  NOR2_X2 U10098 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7743) );
  NOR2_X1 U10099 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), 
        .ZN(n7682) );
  NOR2_X1 U10100 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n7681) );
  NOR2_X2 U10101 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), 
        .ZN(n7699) );
  NOR2_X2 U10102 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), 
        .ZN(n7698) );
  NOR2_X1 U10103 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n7686) );
  NAND2_X1 U10104 ( .A1(n13632), .A2(n7750), .ZN(n7690) );
  NAND2_X1 U10105 ( .A1(n12050), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7689) );
  XNOR2_X1 U10106 ( .A(n7693), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8178) );
  INV_X1 U10107 ( .A(n10141), .ZN(n7710) );
  INV_X1 U10108 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7696) );
  NAND4_X1 U10109 ( .A1(n7699), .A2(n7698), .A3(n7697), .A4(n7696), .ZN(n7990)
         );
  INV_X1 U10110 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7700) );
  NAND3_X1 U10111 ( .A1(n7875), .A2(n7701), .A3(n7700), .ZN(n7702) );
  NOR2_X1 U10112 ( .A1(n7990), .A2(n7702), .ZN(n7703) );
  NAND2_X1 U10113 ( .A1(n7857), .A2(n7703), .ZN(n8005) );
  INV_X1 U10114 ( .A(n8005), .ZN(n7705) );
  INV_X1 U10115 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7704) );
  NAND2_X1 U10116 ( .A1(n7705), .A2(n7704), .ZN(n7708) );
  NAND2_X1 U10117 ( .A1(n8222), .A2(n13249), .ZN(n12053) );
  NAND2_X1 U10118 ( .A1(n7710), .A2(n12053), .ZN(n14853) );
  INV_X1 U10119 ( .A(n8079), .ZN(n7716) );
  NAND2_X1 U10120 ( .A1(n7716), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7721) );
  INV_X1 U10121 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10666) );
  OR2_X1 U10122 ( .A1(n7754), .A2(n10666), .ZN(n7719) );
  NAND2_X1 U10123 ( .A1(n8076), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7718) );
  INV_X1 U10124 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9830) );
  INV_X1 U10125 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7723) );
  NAND2_X1 U10126 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n7722) );
  XNOR2_X1 U10127 ( .A(n7726), .B(n7727), .ZN(n8342) );
  INV_X1 U10128 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7729) );
  INV_X1 U10129 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10632) );
  NAND2_X1 U10130 ( .A1(n7788), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7731) );
  NAND2_X1 U10131 ( .A1(n8076), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7730) );
  NAND2_X1 U10132 ( .A1(n9046), .A2(n8917), .ZN(n7734) );
  NAND2_X1 U10133 ( .A1(n7735), .A2(n7734), .ZN(n13653) );
  INV_X1 U10134 ( .A(n11872), .ZN(n10176) );
  NAND2_X1 U10135 ( .A1(n10176), .A2(n11869), .ZN(n7736) );
  INV_X1 U10136 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7737) );
  INV_X1 U10137 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n7738) );
  INV_X1 U10138 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n13144) );
  OR2_X1 U10139 ( .A1(n7754), .A2(n13144), .ZN(n7740) );
  INV_X1 U10140 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9939) );
  OR2_X1 U10141 ( .A1(n7951), .A2(n9939), .ZN(n7739) );
  OR2_X1 U10142 ( .A1(n7743), .A2(n7711), .ZN(n7744) );
  XNOR2_X1 U10143 ( .A(n7745), .B(n7744), .ZN(n13152) );
  OAI22_X1 U10144 ( .A1(n7724), .A2(n9866), .B1(n9892), .B2(n13152), .ZN(n7746) );
  XNOR2_X1 U10145 ( .A(n7749), .B(n7748), .ZN(n9847) );
  NAND2_X1 U10146 ( .A1(n7750), .A2(n9847), .ZN(n7751) );
  INV_X1 U10147 ( .A(n13142), .ZN(n10264) );
  NAND2_X1 U10148 ( .A1(n10264), .A2(n14837), .ZN(n7752) );
  NAND2_X1 U10149 ( .A1(n9917), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7758) );
  INV_X1 U10150 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7753) );
  OR2_X1 U10151 ( .A1(n7965), .A2(n7753), .ZN(n7757) );
  OR2_X1 U10152 ( .A1(n7754), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7756) );
  INV_X1 U10153 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9942) );
  OR2_X1 U10154 ( .A1(n7951), .A2(n9942), .ZN(n7755) );
  NAND2_X1 U10155 ( .A1(n7759), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7760) );
  XNOR2_X1 U10156 ( .A(n7760), .B(n7678), .ZN(n13166) );
  OAI22_X1 U10157 ( .A1(n7724), .A2(n9868), .B1(n9892), .B2(n13166), .ZN(n7761) );
  INV_X1 U10158 ( .A(n7761), .ZN(n7764) );
  NAND2_X1 U10159 ( .A1(n7750), .A2(n9855), .ZN(n7763) );
  INV_X1 U10160 ( .A(n13141), .ZN(n10512) );
  NAND2_X1 U10161 ( .A1(n10512), .A2(n6828), .ZN(n7765) );
  XNOR2_X1 U10162 ( .A(n7767), .B(n7766), .ZN(n9857) );
  NAND2_X1 U10163 ( .A1(n9857), .A2(n7750), .ZN(n7771) );
  INV_X1 U10164 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9870) );
  NAND2_X1 U10165 ( .A1(n7768), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7781) );
  XNOR2_X1 U10166 ( .A(n7780), .B(n7781), .ZN(n13181) );
  OAI22_X1 U10167 ( .A1(n7724), .A2(n9870), .B1(n9892), .B2(n13181), .ZN(n7769) );
  INV_X1 U10168 ( .A(n7769), .ZN(n7770) );
  INV_X1 U10169 ( .A(n14844), .ZN(n10778) );
  INV_X1 U10170 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n7772) );
  OR2_X1 U10171 ( .A1(n7965), .A2(n7772), .ZN(n7775) );
  NAND2_X1 U10172 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n7790) );
  OAI21_X1 U10173 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n7790), .ZN(n10777) );
  OR2_X1 U10174 ( .A1(n8150), .A2(n10777), .ZN(n7774) );
  INV_X1 U10175 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9945) );
  OR2_X1 U10176 ( .A1(n7951), .A2(n9945), .ZN(n7773) );
  NAND4_X1 U10177 ( .A1(n7776), .A2(n7775), .A3(n7774), .A4(n7773), .ZN(n13140) );
  NAND2_X1 U10178 ( .A1(n7777), .A2(n14844), .ZN(n7778) );
  NAND2_X1 U10179 ( .A1(n9861), .A2(n7750), .ZN(n7787) );
  INV_X1 U10180 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9872) );
  NAND2_X1 U10181 ( .A1(n7781), .A2(n7780), .ZN(n7782) );
  NAND2_X1 U10182 ( .A1(n7782), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7784) );
  XNOR2_X1 U10183 ( .A(n7784), .B(n7783), .ZN(n10081) );
  OAI22_X1 U10184 ( .A1(n7724), .A2(n9872), .B1(n9892), .B2(n10081), .ZN(n7785) );
  INV_X1 U10185 ( .A(n7785), .ZN(n7786) );
  NAND2_X1 U10186 ( .A1(n7787), .A2(n7786), .ZN(n11907) );
  NAND2_X1 U10187 ( .A1(n9918), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7795) );
  INV_X1 U10188 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10704) );
  OR2_X1 U10189 ( .A1(n6827), .A2(n10704), .ZN(n7794) );
  INV_X1 U10190 ( .A(n7790), .ZN(n7789) );
  NAND2_X1 U10191 ( .A1(n7789), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7808) );
  INV_X1 U10192 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n15290) );
  NAND2_X1 U10193 ( .A1(n7790), .A2(n15290), .ZN(n7791) );
  NAND2_X1 U10194 ( .A1(n7808), .A2(n7791), .ZN(n10706) );
  OR2_X1 U10195 ( .A1(n8150), .A2(n10706), .ZN(n7793) );
  INV_X1 U10196 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9949) );
  OR2_X1 U10197 ( .A1(n7951), .A2(n9949), .ZN(n7792) );
  NAND4_X1 U10198 ( .A1(n7795), .A2(n7794), .A3(n7793), .A4(n7792), .ZN(n13139) );
  XNOR2_X1 U10199 ( .A(n11907), .B(n13139), .ZN(n12110) );
  INV_X1 U10200 ( .A(n13139), .ZN(n10511) );
  NAND2_X1 U10201 ( .A1(n11907), .A2(n10511), .ZN(n7796) );
  XNOR2_X1 U10202 ( .A(n7798), .B(n7797), .ZN(n9873) );
  NAND2_X1 U10203 ( .A1(n9873), .A2(n7750), .ZN(n7804) );
  INV_X1 U10204 ( .A(n7768), .ZN(n7800) );
  NOR2_X1 U10205 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n7799) );
  NAND2_X1 U10206 ( .A1(n7800), .A2(n7799), .ZN(n7817) );
  NAND2_X1 U10207 ( .A1(n7817), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7801) );
  XNOR2_X1 U10208 ( .A(n7801), .B(n7818), .ZN(n13196) );
  OAI22_X1 U10209 ( .A1(n7724), .A2(n9876), .B1(n9892), .B2(n13196), .ZN(n7802) );
  INV_X1 U10210 ( .A(n7802), .ZN(n7803) );
  NAND2_X1 U10212 ( .A1(n9917), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7813) );
  INV_X1 U10213 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7805) );
  OR2_X1 U10214 ( .A1(n7965), .A2(n7805), .ZN(n7812) );
  INV_X1 U10215 ( .A(n7808), .ZN(n7806) );
  NAND2_X1 U10216 ( .A1(n7806), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7828) );
  INV_X1 U10217 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7807) );
  NAND2_X1 U10218 ( .A1(n7808), .A2(n7807), .ZN(n7809) );
  NAND2_X1 U10219 ( .A1(n7828), .A2(n7809), .ZN(n13082) );
  OR2_X1 U10220 ( .A1(n8150), .A2(n13082), .ZN(n7811) );
  INV_X1 U10221 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10067) );
  OR2_X1 U10222 ( .A1(n9921), .A2(n10067), .ZN(n7810) );
  NAND4_X1 U10223 ( .A1(n7813), .A2(n7812), .A3(n7811), .A4(n7810), .ZN(n13138) );
  XNOR2_X1 U10224 ( .A(n13080), .B(n13138), .ZN(n12111) );
  INV_X1 U10225 ( .A(n13138), .ZN(n10602) );
  NAND2_X1 U10226 ( .A1(n13080), .A2(n10602), .ZN(n7814) );
  XNOR2_X1 U10227 ( .A(n7816), .B(n7815), .ZN(n9877) );
  NAND2_X1 U10228 ( .A1(n9877), .A2(n7750), .ZN(n7824) );
  INV_X1 U10229 ( .A(n7817), .ZN(n7819) );
  NAND2_X1 U10230 ( .A1(n7819), .A2(n7818), .ZN(n7838) );
  NAND2_X1 U10231 ( .A1(n7838), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7821) );
  INV_X1 U10232 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n7820) );
  XNOR2_X1 U10233 ( .A(n7821), .B(n7820), .ZN(n13210) );
  OAI22_X1 U10234 ( .A1(n7724), .A2(n9878), .B1(n9892), .B2(n13210), .ZN(n7822) );
  INV_X1 U10235 ( .A(n7822), .ZN(n7823) );
  NAND2_X1 U10236 ( .A1(n9917), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7833) );
  INV_X1 U10237 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7825) );
  OR2_X1 U10238 ( .A1(n7965), .A2(n7825), .ZN(n7832) );
  INV_X1 U10239 ( .A(n7828), .ZN(n7826) );
  NAND2_X1 U10240 ( .A1(n7826), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7847) );
  INV_X1 U10241 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7827) );
  NAND2_X1 U10242 ( .A1(n7828), .A2(n7827), .ZN(n7829) );
  NAND2_X1 U10243 ( .A1(n7847), .A2(n7829), .ZN(n10853) );
  OR2_X1 U10244 ( .A1(n8150), .A2(n10853), .ZN(n7831) );
  INV_X1 U10245 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10070) );
  OR2_X1 U10246 ( .A1(n9921), .A2(n10070), .ZN(n7830) );
  NAND4_X1 U10247 ( .A1(n7833), .A2(n7832), .A3(n7831), .A4(n7830), .ZN(n13137) );
  INV_X1 U10248 ( .A(n13137), .ZN(n11921) );
  OR2_X1 U10249 ( .A1(n11919), .A2(n11921), .ZN(n7834) );
  NAND2_X1 U10250 ( .A1(n11919), .A2(n11921), .ZN(n7835) );
  XNOR2_X1 U10251 ( .A(n7837), .B(n7836), .ZN(n9880) );
  NAND2_X1 U10252 ( .A1(n9880), .A2(n7750), .ZN(n7843) );
  OAI21_X1 U10253 ( .B1(n7838), .B2(P2_IR_REG_7__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7840) );
  INV_X1 U10254 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7839) );
  XNOR2_X1 U10255 ( .A(n7840), .B(n7839), .ZN(n13227) );
  OAI22_X1 U10256 ( .A1(n7724), .A2(n9881), .B1(n9892), .B2(n13227), .ZN(n7841) );
  INV_X1 U10257 ( .A(n7841), .ZN(n7842) );
  NAND2_X1 U10258 ( .A1(n9917), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7852) );
  INV_X1 U10259 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7844) );
  OR2_X1 U10260 ( .A1(n7965), .A2(n7844), .ZN(n7851) );
  INV_X1 U10261 ( .A(n7847), .ZN(n7845) );
  NAND2_X1 U10262 ( .A1(n7845), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7866) );
  INV_X1 U10263 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7846) );
  NAND2_X1 U10264 ( .A1(n7847), .A2(n7846), .ZN(n7848) );
  NAND2_X1 U10265 ( .A1(n7866), .A2(n7848), .ZN(n11133) );
  OR2_X1 U10266 ( .A1(n8150), .A2(n11133), .ZN(n7850) );
  OR2_X1 U10267 ( .A1(n9921), .A2(n13221), .ZN(n7849) );
  NAND4_X1 U10268 ( .A1(n7852), .A2(n7851), .A3(n7850), .A4(n7849), .ZN(n13136) );
  INV_X1 U10269 ( .A(n13136), .ZN(n7853) );
  XNOR2_X1 U10270 ( .A(n11932), .B(n7853), .ZN(n12115) );
  OR2_X1 U10271 ( .A1(n11932), .A2(n7853), .ZN(n7854) );
  XNOR2_X1 U10272 ( .A(n7856), .B(n7855), .ZN(n9884) );
  NAND2_X1 U10273 ( .A1(n9884), .A2(n7750), .ZN(n7864) );
  NOR2_X1 U10274 ( .A1(n7857), .A2(n7711), .ZN(n7858) );
  MUX2_X1 U10275 ( .A(n7711), .B(n7858), .S(P2_IR_REG_9__SCAN_IN), .Z(n7861)
         );
  INV_X1 U10276 ( .A(n7859), .ZN(n7860) );
  OR2_X1 U10277 ( .A1(n7861), .A2(n7860), .ZN(n14768) );
  OAI22_X1 U10278 ( .A1(n7724), .A2(n15276), .B1(n9892), .B2(n14768), .ZN(
        n7862) );
  INV_X1 U10279 ( .A(n7862), .ZN(n7863) );
  NAND2_X1 U10280 ( .A1(n9918), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7871) );
  INV_X1 U10281 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n13474) );
  OR2_X1 U10282 ( .A1(n6827), .A2(n13474), .ZN(n7870) );
  NAND2_X1 U10283 ( .A1(n7866), .A2(n7865), .ZN(n7867) );
  NAND2_X1 U10284 ( .A1(n7882), .A2(n7867), .ZN(n13473) );
  OR2_X1 U10285 ( .A1(n8150), .A2(n13473), .ZN(n7869) );
  INV_X1 U10286 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10076) );
  OR2_X1 U10287 ( .A1(n9921), .A2(n10076), .ZN(n7868) );
  NAND4_X1 U10288 ( .A1(n7871), .A2(n7870), .A3(n7869), .A4(n7868), .ZN(n13135) );
  INV_X1 U10289 ( .A(n13135), .ZN(n11940) );
  XNOR2_X1 U10290 ( .A(n13477), .B(n11940), .ZN(n12116) );
  INV_X1 U10291 ( .A(n12116), .ZN(n11236) );
  OR2_X1 U10292 ( .A1(n13477), .A2(n11940), .ZN(n7872) );
  XNOR2_X1 U10293 ( .A(n7874), .B(n7873), .ZN(n9924) );
  NAND2_X1 U10294 ( .A1(n9924), .A2(n7750), .ZN(n7879) );
  NAND2_X1 U10295 ( .A1(n7859), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7876) );
  XNOR2_X1 U10296 ( .A(n7876), .B(n7875), .ZN(n10123) );
  OAI22_X1 U10297 ( .A1(n7724), .A2(n9925), .B1(n9892), .B2(n10123), .ZN(n7877) );
  INV_X1 U10298 ( .A(n7877), .ZN(n7878) );
  NAND2_X1 U10299 ( .A1(n9918), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7888) );
  INV_X1 U10300 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11281) );
  OR2_X1 U10301 ( .A1(n6827), .A2(n11281), .ZN(n7887) );
  INV_X1 U10302 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7881) );
  NAND2_X1 U10303 ( .A1(n7882), .A2(n7881), .ZN(n7883) );
  NAND2_X1 U10304 ( .A1(n7900), .A2(n7883), .ZN(n11297) );
  OR2_X1 U10305 ( .A1(n8150), .A2(n11297), .ZN(n7886) );
  INV_X1 U10306 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7884) );
  OR2_X1 U10307 ( .A1(n9921), .A2(n7884), .ZN(n7885) );
  NAND4_X1 U10308 ( .A1(n7888), .A2(n7887), .A3(n7886), .A4(n7885), .ZN(n13134) );
  INV_X1 U10309 ( .A(n13134), .ZN(n7889) );
  XNOR2_X1 U10310 ( .A(n11946), .B(n7889), .ZN(n12117) );
  INV_X1 U10311 ( .A(n12117), .ZN(n11285) );
  OR2_X1 U10312 ( .A1(n11946), .A2(n7889), .ZN(n7890) );
  XNOR2_X1 U10313 ( .A(n7892), .B(n7891), .ZN(n9958) );
  NAND2_X1 U10314 ( .A1(n9958), .A2(n7750), .ZN(n7897) );
  NAND2_X1 U10315 ( .A1(n7991), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7894) );
  INV_X1 U10316 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n7893) );
  XNOR2_X1 U10317 ( .A(n7894), .B(n7893), .ZN(n10311) );
  OAI22_X1 U10318 ( .A1(n7724), .A2(n15289), .B1(n9892), .B2(n10311), .ZN(
        n7895) );
  INV_X1 U10319 ( .A(n7895), .ZN(n7896) );
  NAND2_X1 U10320 ( .A1(n9917), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7905) );
  INV_X1 U10321 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7898) );
  OR2_X1 U10322 ( .A1(n7965), .A2(n7898), .ZN(n7904) );
  NAND2_X1 U10323 ( .A1(n7900), .A2(n7899), .ZN(n7901) );
  NAND2_X1 U10324 ( .A1(n7914), .A2(n7901), .ZN(n11451) );
  OR2_X1 U10325 ( .A1(n8150), .A2(n11451), .ZN(n7903) );
  INV_X1 U10326 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10124) );
  OR2_X1 U10327 ( .A1(n7951), .A2(n10124), .ZN(n7902) );
  NAND4_X1 U10328 ( .A1(n7905), .A2(n7904), .A3(n7903), .A4(n7902), .ZN(n13133) );
  XNOR2_X1 U10329 ( .A(n11953), .B(n13133), .ZN(n12120) );
  INV_X1 U10330 ( .A(n12120), .ZN(n11444) );
  XNOR2_X1 U10331 ( .A(n7906), .B(n7549), .ZN(n9962) );
  NAND2_X1 U10332 ( .A1(n9962), .A2(n7750), .ZN(n7911) );
  NAND2_X1 U10333 ( .A1(n7925), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7908) );
  INV_X1 U10334 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7907) );
  XNOR2_X1 U10335 ( .A(n7908), .B(n7907), .ZN(n14779) );
  OAI22_X1 U10336 ( .A1(n7724), .A2(n9963), .B1(n9892), .B2(n14779), .ZN(n7909) );
  INV_X1 U10337 ( .A(n7909), .ZN(n7910) );
  NAND2_X1 U10338 ( .A1(n9918), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7919) );
  INV_X1 U10339 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11469) );
  OR2_X1 U10340 ( .A1(n6827), .A2(n11469), .ZN(n7918) );
  INV_X1 U10341 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7913) );
  NAND2_X1 U10342 ( .A1(n7914), .A2(n7913), .ZN(n7915) );
  NAND2_X1 U10343 ( .A1(n7929), .A2(n7915), .ZN(n11579) );
  OR2_X1 U10344 ( .A1(n8150), .A2(n11579), .ZN(n7917) );
  INV_X1 U10345 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10307) );
  OR2_X1 U10346 ( .A1(n7951), .A2(n10307), .ZN(n7916) );
  NAND4_X1 U10347 ( .A1(n7919), .A2(n7918), .A3(n7917), .A4(n7916), .ZN(n13131) );
  INV_X1 U10348 ( .A(n13131), .ZN(n7920) );
  OR2_X1 U10349 ( .A1(n11961), .A2(n7920), .ZN(n7923) );
  NAND2_X1 U10350 ( .A1(n11961), .A2(n7920), .ZN(n7921) );
  NAND2_X1 U10351 ( .A1(n7923), .A2(n7921), .ZN(n12119) );
  INV_X1 U10352 ( .A(n13133), .ZN(n11955) );
  AND2_X1 U10353 ( .A1(n11953), .A2(n11955), .ZN(n11459) );
  NOR2_X1 U10354 ( .A1(n12119), .A2(n11459), .ZN(n7922) );
  XNOR2_X1 U10355 ( .A(n7924), .B(n7563), .ZN(n9969) );
  NAND2_X1 U10356 ( .A1(n9969), .A2(n7750), .ZN(n7928) );
  NOR2_X1 U10357 ( .A1(n7925), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n7940) );
  OR2_X1 U10358 ( .A1(n7940), .A2(n7711), .ZN(n7926) );
  XNOR2_X1 U10359 ( .A(n7926), .B(P2_IR_REG_13__SCAN_IN), .ZN(n10312) );
  AOI22_X1 U10360 ( .A1(n12050), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6715), 
        .B2(n10312), .ZN(n7927) );
  NAND2_X1 U10361 ( .A1(n9917), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7934) );
  INV_X1 U10362 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n15190) );
  OR2_X1 U10363 ( .A1(n7965), .A2(n15190), .ZN(n7933) );
  NAND2_X1 U10364 ( .A1(n7929), .A2(n10315), .ZN(n7930) );
  NAND2_X1 U10365 ( .A1(n7947), .A2(n7930), .ZN(n11662) );
  OR2_X1 U10366 ( .A1(n8150), .A2(n11662), .ZN(n7932) );
  INV_X1 U10367 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n15221) );
  OR2_X1 U10368 ( .A1(n7951), .A2(n15221), .ZN(n7931) );
  NAND4_X1 U10369 ( .A1(n7934), .A2(n7933), .A3(n7932), .A4(n7931), .ZN(n13130) );
  XNOR2_X1 U10370 ( .A(n11969), .B(n13130), .ZN(n12122) );
  INV_X1 U10371 ( .A(n13130), .ZN(n7935) );
  OR2_X1 U10372 ( .A1(n11969), .A2(n7935), .ZN(n7936) );
  XNOR2_X1 U10373 ( .A(n7937), .B(n7938), .ZN(n10257) );
  NAND2_X1 U10374 ( .A1(n10257), .A2(n7750), .ZN(n7946) );
  INV_X1 U10375 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7939) );
  NAND2_X1 U10376 ( .A1(n7940), .A2(n7939), .ZN(n7942) );
  NAND2_X1 U10377 ( .A1(n7942), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7941) );
  MUX2_X1 U10378 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7941), .S(
        P2_IR_REG_14__SCAN_IN), .Z(n7943) );
  NAND2_X1 U10379 ( .A1(n7943), .A2(n7975), .ZN(n11310) );
  OAI22_X1 U10380 ( .A1(n11310), .A2(n9892), .B1(n7724), .B2(n10259), .ZN(
        n7944) );
  INV_X1 U10381 ( .A(n7944), .ZN(n7945) );
  NAND2_X1 U10382 ( .A1(n7947), .A2(n11787), .ZN(n7948) );
  AND2_X1 U10383 ( .A1(n7968), .A2(n7948), .ZN(n11790) );
  NAND2_X1 U10384 ( .A1(n8175), .A2(n11790), .ZN(n7955) );
  INV_X1 U10385 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7949) );
  OR2_X1 U10386 ( .A1(n7965), .A2(n7949), .ZN(n7954) );
  INV_X1 U10387 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7950) );
  OR2_X1 U10388 ( .A1(n6827), .A2(n7950), .ZN(n7953) );
  INV_X1 U10389 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11303) );
  OR2_X1 U10390 ( .A1(n7951), .A2(n11303), .ZN(n7952) );
  OR2_X1 U10391 ( .A1(n11968), .A2(n13129), .ZN(n7956) );
  NAND2_X1 U10392 ( .A1(n11968), .A2(n13129), .ZN(n7957) );
  XNOR2_X1 U10393 ( .A(n7959), .B(n7960), .ZN(n10423) );
  NAND2_X1 U10394 ( .A1(n10423), .A2(n7750), .ZN(n7963) );
  NAND2_X1 U10395 ( .A1(n7975), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7961) );
  XNOR2_X1 U10396 ( .A(n7961), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14805) );
  AOI22_X1 U10397 ( .A1(n14805), .A2(n6715), .B1(n12050), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n7962) );
  INV_X1 U10398 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n13557) );
  INV_X1 U10399 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7964) );
  OR2_X1 U10400 ( .A1(n6827), .A2(n7964), .ZN(n7967) );
  INV_X1 U10401 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n13615) );
  OR2_X1 U10402 ( .A1(n7965), .A2(n13615), .ZN(n7966) );
  AND2_X1 U10403 ( .A1(n7967), .A2(n7966), .ZN(n7971) );
  INV_X1 U10404 ( .A(n7979), .ZN(n7981) );
  NAND2_X1 U10405 ( .A1(n7968), .A2(n13106), .ZN(n7969) );
  NAND2_X1 U10406 ( .A1(n7981), .A2(n7969), .ZN(n11774) );
  OR2_X1 U10407 ( .A1(n11774), .A2(n8150), .ZN(n7970) );
  OAI211_X1 U10408 ( .C1(n9921), .C2(n13557), .A(n7971), .B(n7970), .ZN(n13128) );
  INV_X1 U10409 ( .A(n13128), .ZN(n9740) );
  NAND2_X1 U10410 ( .A1(n13617), .A2(n9740), .ZN(n7973) );
  OR2_X1 U10411 ( .A1(n13617), .A2(n9740), .ZN(n7972) );
  NAND2_X1 U10412 ( .A1(n7973), .A2(n7972), .ZN(n12124) );
  XNOR2_X1 U10413 ( .A(n7974), .B(n7565), .ZN(n10527) );
  NAND2_X1 U10414 ( .A1(n10527), .A2(n7750), .ZN(n7978) );
  OAI21_X1 U10415 ( .B1(n7975), .B2(P2_IR_REG_15__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7976) );
  XNOR2_X1 U10416 ( .A(n7976), .B(P2_IR_REG_16__SCAN_IN), .ZN(n11316) );
  AOI22_X1 U10417 ( .A1(n11316), .A2(n6715), .B1(n12050), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n7977) );
  INV_X1 U10418 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n13553) );
  INV_X1 U10419 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7980) );
  NAND2_X1 U10420 ( .A1(n7981), .A2(n7980), .ZN(n7982) );
  NAND2_X1 U10421 ( .A1(n7996), .A2(n7982), .ZN(n13456) );
  OR2_X1 U10422 ( .A1(n13456), .A2(n8150), .ZN(n7984) );
  AOI22_X1 U10423 ( .A1(n9917), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n9918), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n7983) );
  OAI211_X1 U10424 ( .C1(n9921), .C2(n13553), .A(n7984), .B(n7983), .ZN(n13127) );
  INV_X1 U10425 ( .A(n13127), .ZN(n13027) );
  OR2_X1 U10426 ( .A1(n13551), .A2(n13027), .ZN(n7985) );
  NAND2_X1 U10427 ( .A1(n13551), .A2(n13027), .ZN(n7986) );
  XNOR2_X1 U10428 ( .A(n7987), .B(SI_17_), .ZN(n7988) );
  XNOR2_X1 U10429 ( .A(n7989), .B(n7988), .ZN(n10586) );
  NAND2_X1 U10430 ( .A1(n10586), .A2(n7750), .ZN(n7995) );
  OAI21_X1 U10431 ( .B1(n7991), .B2(n7990), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n7992) );
  XNOR2_X1 U10432 ( .A(n7992), .B(P2_IR_REG_17__SCAN_IN), .ZN(n14817) );
  INV_X1 U10433 ( .A(n14817), .ZN(n11534) );
  OAI22_X1 U10434 ( .A1(n7724), .A2(n10587), .B1(n9892), .B2(n11534), .ZN(
        n7993) );
  INV_X1 U10435 ( .A(n7993), .ZN(n7994) );
  NAND2_X1 U10436 ( .A1(n7996), .A2(n13030), .ZN(n7997) );
  NAND2_X1 U10437 ( .A1(n8011), .A2(n7997), .ZN(n13438) );
  AOI22_X1 U10438 ( .A1(n8076), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n9918), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n7999) );
  INV_X1 U10439 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13439) );
  OR2_X1 U10440 ( .A1(n6827), .A2(n13439), .ZN(n7998) );
  OAI211_X1 U10441 ( .C1(n13438), .C2(n8150), .A(n7999), .B(n7998), .ZN(n13126) );
  XNOR2_X1 U10442 ( .A(n11978), .B(n13126), .ZN(n13431) );
  INV_X1 U10443 ( .A(n13126), .ZN(n13066) );
  OR2_X1 U10444 ( .A1(n11978), .A2(n13066), .ZN(n8000) );
  NAND2_X1 U10445 ( .A1(n8001), .A2(n8002), .ZN(n8003) );
  NAND2_X1 U10446 ( .A1(n8004), .A2(n8003), .ZN(n10966) );
  OR2_X1 U10447 ( .A1(n10966), .A2(n8088), .ZN(n8008) );
  NAND2_X1 U10448 ( .A1(n8005), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8006) );
  XNOR2_X1 U10449 ( .A(n8006), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13241) );
  AOI22_X1 U10450 ( .A1(n12050), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6715), 
        .B2(n13241), .ZN(n8007) );
  INV_X1 U10451 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8010) );
  NAND2_X1 U10452 ( .A1(n8011), .A2(n8010), .ZN(n8012) );
  NAND2_X1 U10453 ( .A1(n8028), .A2(n8012), .ZN(n13418) );
  OR2_X1 U10454 ( .A1(n13418), .A2(n8150), .ZN(n8018) );
  INV_X1 U10455 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8015) );
  NAND2_X1 U10456 ( .A1(n9918), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8014) );
  NAND2_X1 U10457 ( .A1(n9917), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8013) );
  OAI211_X1 U10458 ( .C1(n9921), .C2(n8015), .A(n8014), .B(n8013), .ZN(n8016)
         );
  INV_X1 U10459 ( .A(n8016), .ZN(n8017) );
  INV_X1 U10460 ( .A(n13028), .ZN(n12981) );
  NAND2_X1 U10461 ( .A1(n13541), .A2(n13028), .ZN(n8019) );
  XNOR2_X1 U10462 ( .A(n8021), .B(n8022), .ZN(n11162) );
  NAND2_X1 U10463 ( .A1(n11162), .A2(n7750), .ZN(n8026) );
  INV_X1 U10464 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8023) );
  OAI22_X1 U10465 ( .A1(n7724), .A2(n8023), .B1(n13249), .B2(n9892), .ZN(n8024) );
  INV_X1 U10466 ( .A(n8024), .ZN(n8025) );
  INV_X1 U10467 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8027) );
  NAND2_X1 U10468 ( .A1(n8028), .A2(n8027), .ZN(n8029) );
  AND2_X1 U10469 ( .A1(n8044), .A2(n8029), .ZN(n13405) );
  NAND2_X1 U10470 ( .A1(n13405), .A2(n8175), .ZN(n8035) );
  INV_X1 U10471 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U10472 ( .A1(n9917), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8031) );
  NAND2_X1 U10473 ( .A1(n9918), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8030) );
  OAI211_X1 U10474 ( .C1(n8032), .C2(n9921), .A(n8031), .B(n8030), .ZN(n8033)
         );
  INV_X1 U10475 ( .A(n8033), .ZN(n8034) );
  NAND2_X1 U10476 ( .A1(n8035), .A2(n8034), .ZN(n13125) );
  INV_X1 U10477 ( .A(n13125), .ZN(n13067) );
  OR2_X1 U10478 ( .A1(n13537), .A2(n13067), .ZN(n8036) );
  NAND2_X1 U10479 ( .A1(n13400), .A2(n8036), .ZN(n8038) );
  NAND2_X1 U10480 ( .A1(n13537), .A2(n13067), .ZN(n8037) );
  NAND2_X1 U10481 ( .A1(n12050), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8041) );
  INV_X1 U10482 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8043) );
  NAND2_X1 U10483 ( .A1(n8044), .A2(n8043), .ZN(n8045) );
  NAND2_X1 U10484 ( .A1(n8058), .A2(n8045), .ZN(n13389) );
  OR2_X1 U10485 ( .A1(n13389), .A2(n8150), .ZN(n8050) );
  INV_X1 U10486 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n13388) );
  NAND2_X1 U10487 ( .A1(n8076), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8047) );
  NAND2_X1 U10488 ( .A1(n9918), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8046) );
  OAI211_X1 U10489 ( .C1(n6827), .C2(n13388), .A(n8047), .B(n8046), .ZN(n8048)
         );
  INV_X1 U10490 ( .A(n8048), .ZN(n8049) );
  NAND2_X1 U10491 ( .A1(n8053), .A2(n8052), .ZN(n8055) );
  NAND2_X1 U10492 ( .A1(n8055), .A2(n8054), .ZN(n11857) );
  OR2_X1 U10493 ( .A1(n11857), .A2(n8088), .ZN(n8057) );
  NAND2_X1 U10494 ( .A1(n12050), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8056) );
  INV_X1 U10495 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13003) );
  NAND2_X1 U10496 ( .A1(n8058), .A2(n13003), .ZN(n8059) );
  AND2_X1 U10497 ( .A1(n8074), .A2(n8059), .ZN(n13374) );
  NAND2_X1 U10498 ( .A1(n13374), .A2(n8175), .ZN(n8064) );
  INV_X1 U10499 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13527) );
  NAND2_X1 U10500 ( .A1(n9917), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8061) );
  NAND2_X1 U10501 ( .A1(n9918), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8060) );
  OAI211_X1 U10502 ( .C1(n13527), .C2(n9921), .A(n8061), .B(n8060), .ZN(n8062)
         );
  INV_X1 U10503 ( .A(n8062), .ZN(n8063) );
  NAND2_X1 U10504 ( .A1(n13376), .A2(n13123), .ZN(n8065) );
  INV_X1 U10505 ( .A(n8066), .ZN(n8067) );
  NAND2_X1 U10506 ( .A1(n7084), .A2(n8067), .ZN(n8068) );
  AND2_X1 U10507 ( .A1(n8069), .A2(n8068), .ZN(n11708) );
  NAND2_X1 U10508 ( .A1(n11708), .A2(n7750), .ZN(n8071) );
  NAND2_X1 U10509 ( .A1(n12050), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8070) );
  INV_X1 U10510 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8073) );
  NAND2_X1 U10511 ( .A1(n8074), .A2(n8073), .ZN(n8075) );
  NAND2_X1 U10512 ( .A1(n8093), .A2(n8075), .ZN(n13361) );
  OR2_X1 U10513 ( .A1(n13361), .A2(n8150), .ZN(n8082) );
  INV_X1 U10514 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13360) );
  NAND2_X1 U10515 ( .A1(n8076), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8078) );
  NAND2_X1 U10516 ( .A1(n9918), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8077) );
  OAI211_X1 U10517 ( .C1(n6827), .C2(n13360), .A(n8078), .B(n8077), .ZN(n8080)
         );
  INV_X1 U10518 ( .A(n8080), .ZN(n8081) );
  NAND2_X1 U10519 ( .A1(n8082), .A2(n8081), .ZN(n13122) );
  XNOR2_X1 U10520 ( .A(n13591), .B(n12030), .ZN(n13356) );
  INV_X1 U10521 ( .A(n13356), .ZN(n13365) );
  NOR2_X1 U10522 ( .A1(n13591), .A2(n12030), .ZN(n8083) );
  NAND2_X1 U10523 ( .A1(n8087), .A2(n8086), .ZN(n11747) );
  OR2_X1 U10524 ( .A1(n11747), .A2(n8088), .ZN(n8090) );
  NAND2_X1 U10525 ( .A1(n12050), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8089) );
  INV_X1 U10526 ( .A(n8093), .ZN(n8091) );
  INV_X1 U10527 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8092) );
  NAND2_X1 U10528 ( .A1(n8093), .A2(n8092), .ZN(n8094) );
  NAND2_X1 U10529 ( .A1(n8106), .A2(n8094), .ZN(n12967) );
  OR2_X1 U10530 ( .A1(n12967), .A2(n8150), .ZN(n8100) );
  INV_X1 U10531 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8097) );
  NAND2_X1 U10532 ( .A1(n9917), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8096) );
  NAND2_X1 U10533 ( .A1(n9918), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8095) );
  OAI211_X1 U10534 ( .C1(n8097), .C2(n9921), .A(n8096), .B(n8095), .ZN(n8098)
         );
  INV_X1 U10535 ( .A(n8098), .ZN(n8099) );
  NAND2_X1 U10536 ( .A1(n8100), .A2(n8099), .ZN(n13121) );
  NAND2_X1 U10537 ( .A1(n13348), .A2(n13121), .ZN(n8101) );
  XNOR2_X1 U10538 ( .A(n8103), .B(n8102), .ZN(n13649) );
  NAND2_X1 U10539 ( .A1(n13649), .A2(n7750), .ZN(n8105) );
  NAND2_X1 U10540 ( .A1(n12050), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8104) );
  INV_X1 U10541 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13041) );
  NAND2_X1 U10542 ( .A1(n8106), .A2(n13041), .ZN(n8107) );
  NAND2_X1 U10543 ( .A1(n8120), .A2(n8107), .ZN(n13332) );
  OR2_X1 U10544 ( .A1(n13332), .A2(n8150), .ZN(n8112) );
  INV_X1 U10545 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n13510) );
  NAND2_X1 U10546 ( .A1(n9917), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8109) );
  NAND2_X1 U10547 ( .A1(n9918), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8108) );
  OAI211_X1 U10548 ( .C1(n13510), .C2(n9921), .A(n8109), .B(n8108), .ZN(n8110)
         );
  INV_X1 U10549 ( .A(n8110), .ZN(n8111) );
  NAND2_X1 U10550 ( .A1(n8112), .A2(n8111), .ZN(n13120) );
  XNOR2_X1 U10551 ( .A(n13331), .B(n13120), .ZN(n13329) );
  INV_X1 U10552 ( .A(n13329), .ZN(n8253) );
  NAND2_X1 U10553 ( .A1(n8114), .A2(n8113), .ZN(n8116) );
  NAND2_X1 U10554 ( .A1(n11858), .A2(n7750), .ZN(n8118) );
  NAND2_X1 U10555 ( .A1(n12050), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8117) );
  INV_X1 U10556 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8119) );
  NAND2_X1 U10557 ( .A1(n8120), .A2(n8119), .ZN(n8121) );
  NAND2_X1 U10558 ( .A1(n13318), .A2(n8175), .ZN(n8126) );
  INV_X1 U10559 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n15194) );
  NAND2_X1 U10560 ( .A1(n9917), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8123) );
  NAND2_X1 U10561 ( .A1(n9918), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8122) );
  OAI211_X1 U10562 ( .C1(n15194), .C2(n9921), .A(n8123), .B(n8122), .ZN(n8124)
         );
  INV_X1 U10563 ( .A(n8124), .ZN(n8125) );
  INV_X1 U10564 ( .A(n13093), .ZN(n10638) );
  XNOR2_X1 U10565 ( .A(n13505), .B(n10638), .ZN(n13312) );
  XNOR2_X1 U10566 ( .A(n8127), .B(SI_26_), .ZN(n8128) );
  XNOR2_X1 U10567 ( .A(n8129), .B(n8128), .ZN(n13642) );
  NAND2_X1 U10568 ( .A1(n13642), .A2(n7750), .ZN(n8131) );
  NAND2_X1 U10569 ( .A1(n12050), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8130) );
  INV_X1 U10570 ( .A(n8133), .ZN(n8132) );
  NAND2_X1 U10571 ( .A1(n8132), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8148) );
  INV_X1 U10572 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13096) );
  NAND2_X1 U10573 ( .A1(n8133), .A2(n13096), .ZN(n8134) );
  NAND2_X1 U10574 ( .A1(n8148), .A2(n8134), .ZN(n13301) );
  OR2_X1 U10575 ( .A1(n13301), .A2(n8150), .ZN(n8139) );
  INV_X1 U10576 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n13501) );
  NAND2_X1 U10577 ( .A1(n9918), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8136) );
  NAND2_X1 U10578 ( .A1(n9917), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8135) );
  OAI211_X1 U10579 ( .C1(n9921), .C2(n13501), .A(n8136), .B(n8135), .ZN(n8137)
         );
  INV_X1 U10580 ( .A(n8137), .ZN(n8138) );
  NOR2_X1 U10581 ( .A1(n13500), .A2(n12042), .ZN(n12100) );
  AND2_X1 U10582 ( .A1(n13500), .A2(n12042), .ZN(n12099) );
  INV_X1 U10583 ( .A(n12099), .ZN(n8140) );
  INV_X1 U10584 ( .A(n8141), .ZN(n8142) );
  XNOR2_X1 U10585 ( .A(n8142), .B(SI_27_), .ZN(n8143) );
  XNOR2_X1 U10586 ( .A(n8144), .B(n8143), .ZN(n13639) );
  NAND2_X1 U10587 ( .A1(n13639), .A2(n7750), .ZN(n8146) );
  NAND2_X1 U10588 ( .A1(n12050), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8145) );
  INV_X1 U10589 ( .A(n8148), .ZN(n8147) );
  NAND2_X1 U10590 ( .A1(n8147), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8161) );
  INV_X1 U10591 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9801) );
  NAND2_X1 U10592 ( .A1(n8148), .A2(n9801), .ZN(n8149) );
  NAND2_X1 U10593 ( .A1(n8161), .A2(n8149), .ZN(n13288) );
  OR2_X1 U10594 ( .A1(n13288), .A2(n8150), .ZN(n8155) );
  INV_X1 U10595 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n13495) );
  NAND2_X1 U10596 ( .A1(n9918), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8152) );
  NAND2_X1 U10597 ( .A1(n9917), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8151) );
  OAI211_X1 U10598 ( .C1(n13495), .C2(n9921), .A(n8152), .B(n8151), .ZN(n8153)
         );
  INV_X1 U10599 ( .A(n8153), .ZN(n8154) );
  XNOR2_X1 U10600 ( .A(n13569), .B(n13095), .ZN(n13280) );
  INV_X1 U10601 ( .A(n13280), .ZN(n13282) );
  NAND2_X1 U10602 ( .A1(n14193), .A2(n7750), .ZN(n8159) );
  NAND2_X1 U10603 ( .A1(n12050), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8158) );
  INV_X1 U10604 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8160) );
  NAND2_X1 U10605 ( .A1(n8161), .A2(n8160), .ZN(n8162) );
  NAND2_X1 U10606 ( .A1(n13263), .A2(n8175), .ZN(n8168) );
  INV_X1 U10607 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8165) );
  NAND2_X1 U10608 ( .A1(n9917), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8164) );
  NAND2_X1 U10609 ( .A1(n9918), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8163) );
  OAI211_X1 U10610 ( .C1(n8165), .C2(n9921), .A(n8164), .B(n8163), .ZN(n8166)
         );
  INV_X1 U10611 ( .A(n8166), .ZN(n8167) );
  NAND2_X1 U10612 ( .A1(n13489), .A2(n9793), .ZN(n8169) );
  NAND2_X1 U10613 ( .A1(n8170), .A2(n8169), .ZN(n13261) );
  INV_X1 U10614 ( .A(n13261), .ZN(n13266) );
  NAND2_X1 U10615 ( .A1(n13569), .A2(n13095), .ZN(n13267) );
  INV_X1 U10616 ( .A(n8171), .ZN(n8273) );
  INV_X1 U10617 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8262) );
  NAND2_X1 U10618 ( .A1(n9918), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8173) );
  NAND2_X1 U10619 ( .A1(n9917), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8172) );
  OAI211_X1 U10620 ( .C1(n8262), .C2(n9921), .A(n8173), .B(n8172), .ZN(n8174)
         );
  AOI21_X1 U10621 ( .B1(n8273), .B2(n8175), .A(n8174), .ZN(n12993) );
  XNOR2_X1 U10622 ( .A(n12058), .B(n12993), .ZN(n12134) );
  OR2_X1 U10623 ( .A1(n12138), .A2(n8222), .ZN(n8177) );
  NAND2_X1 U10624 ( .A1(n8221), .A2(n12149), .ZN(n8176) );
  INV_X1 U10625 ( .A(n9890), .ZN(n9787) );
  NOR2_X2 U10626 ( .A1(n9787), .A2(n8179), .ZN(n13050) );
  NAND2_X1 U10627 ( .A1(n8179), .A2(n9890), .ZN(n13094) );
  INV_X1 U10628 ( .A(P2_B_REG_SCAN_IN), .ZN(n8180) );
  NOR2_X1 U10629 ( .A1(n13640), .A2(n8180), .ZN(n8181) );
  NOR2_X1 U10630 ( .A1(n13094), .A2(n8181), .ZN(n12411) );
  INV_X1 U10631 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8184) );
  NAND2_X1 U10632 ( .A1(n9917), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8183) );
  NAND2_X1 U10633 ( .A1(n9918), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8182) );
  OAI211_X1 U10634 ( .C1(n9921), .C2(n8184), .A(n8183), .B(n8182), .ZN(n13116)
         );
  INV_X1 U10635 ( .A(n8185), .ZN(n8186) );
  NAND2_X1 U10636 ( .A1(n10657), .A2(n11889), .ZN(n10776) );
  NOR2_X1 U10637 ( .A1(n10993), .A2(n11932), .ZN(n11233) );
  AND2_X2 U10638 ( .A1(n11233), .A2(n11242), .ZN(n11279) );
  INV_X1 U10639 ( .A(n11946), .ZN(n11383) );
  AND2_X2 U10640 ( .A1(n11279), .A2(n11383), .ZN(n11450) );
  INV_X1 U10641 ( .A(n11953), .ZN(n14854) );
  NAND2_X1 U10642 ( .A1(n11450), .A2(n14854), .ZN(n11467) );
  OR2_X2 U10643 ( .A1(n11467), .A2(n11961), .ZN(n11602) );
  NAND2_X1 U10644 ( .A1(n13422), .A2(n13443), .ZN(n13415) );
  NOR2_X2 U10645 ( .A1(n13537), .A2(n13415), .ZN(n13404) );
  AND2_X1 U10646 ( .A1(n13603), .A2(n13404), .ZN(n13385) );
  INV_X1 U10647 ( .A(n13317), .ZN(n13330) );
  INV_X2 U10648 ( .A(n9775), .ZN(n13372) );
  OAI211_X1 U10649 ( .C1(n12060), .C2(n6554), .A(n13372), .B(n13255), .ZN(
        n8271) );
  NAND2_X1 U10650 ( .A1(n8217), .A2(n8216), .ZN(n8190) );
  NAND2_X1 U10651 ( .A1(n8190), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8192) );
  XNOR2_X1 U10652 ( .A(n13652), .B(P2_B_REG_SCAN_IN), .ZN(n8198) );
  NOR2_X1 U10653 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .ZN(n8193) );
  NAND2_X1 U10654 ( .A1(n8194), .A2(n8193), .ZN(n8196) );
  NAND2_X1 U10655 ( .A1(n8196), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8195) );
  MUX2_X1 U10656 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8195), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8197) );
  NAND2_X1 U10657 ( .A1(n8197), .A2(n8200), .ZN(n13646) );
  NAND2_X1 U10658 ( .A1(n8198), .A2(n13646), .ZN(n8203) );
  NAND2_X1 U10659 ( .A1(n8200), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8201) );
  MUX2_X1 U10660 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8201), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8202) );
  NOR4_X1 U10661 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n8212) );
  OR4_X1 U10662 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n8209) );
  NOR4_X1 U10663 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8207) );
  NOR4_X1 U10664 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n8206) );
  NOR4_X1 U10665 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8205) );
  NOR4_X1 U10666 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8204) );
  NAND4_X1 U10667 ( .A1(n8207), .A2(n8206), .A3(n8205), .A4(n8204), .ZN(n8208)
         );
  NOR4_X1 U10668 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n8209), .A4(n8208), .ZN(n8211) );
  NOR4_X1 U10669 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n8210) );
  NAND3_X1 U10670 ( .A1(n8212), .A2(n8211), .A3(n8210), .ZN(n8213) );
  AND2_X1 U10671 ( .A1(n14827), .A2(n8213), .ZN(n8265) );
  INV_X1 U10672 ( .A(n8265), .ZN(n8223) );
  NOR2_X1 U10673 ( .A1(n13646), .A2(n13652), .ZN(n8214) );
  NAND2_X1 U10674 ( .A1(n8215), .A2(n8214), .ZN(n9807) );
  NAND2_X1 U10675 ( .A1(n9890), .A2(n12053), .ZN(n9798) );
  AND2_X1 U10676 ( .A1(n14835), .A2(n9798), .ZN(n12146) );
  INV_X1 U10677 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14833) );
  NAND2_X1 U10678 ( .A1(n14827), .A2(n14833), .ZN(n8220) );
  NAND2_X1 U10679 ( .A1(n13644), .A2(n13646), .ZN(n8219) );
  NAND2_X1 U10680 ( .A1(n8220), .A2(n8219), .ZN(n14834) );
  NAND2_X1 U10681 ( .A1(n8222), .A2(n8221), .ZN(n10629) );
  NAND4_X1 U10682 ( .A1(n8223), .A2(n12146), .A3(n14834), .A4(n9796), .ZN(
        n9661) );
  INV_X1 U10683 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14830) );
  NAND2_X1 U10684 ( .A1(n14827), .A2(n14830), .ZN(n8225) );
  NAND2_X1 U10685 ( .A1(n13644), .A2(n13652), .ZN(n8224) );
  INV_X1 U10686 ( .A(n12105), .ZN(n10649) );
  NAND2_X1 U10687 ( .A1(n10264), .A2(n11883), .ZN(n8226) );
  NAND2_X1 U10688 ( .A1(n10351), .A2(n12107), .ZN(n10350) );
  NAND2_X1 U10689 ( .A1(n10512), .A2(n11889), .ZN(n8227) );
  NAND2_X1 U10690 ( .A1(n10350), .A2(n8227), .ZN(n10766) );
  NAND2_X1 U10691 ( .A1(n7777), .A2(n10778), .ZN(n8228) );
  NAND2_X1 U10692 ( .A1(n10765), .A2(n8228), .ZN(n10605) );
  INV_X1 U10693 ( .A(n12110), .ZN(n10604) );
  NAND2_X1 U10694 ( .A1(n10605), .A2(n10604), .ZN(n10607) );
  OR2_X1 U10695 ( .A1(n13139), .A2(n11907), .ZN(n8229) );
  NAND2_X1 U10696 ( .A1(n10607), .A2(n8229), .ZN(n11028) );
  INV_X1 U10697 ( .A(n12111), .ZN(n11027) );
  OR2_X1 U10698 ( .A1(n13080), .A2(n13138), .ZN(n8230) );
  NAND2_X1 U10699 ( .A1(n11026), .A2(n8230), .ZN(n10846) );
  XNOR2_X1 U10700 ( .A(n11919), .B(n13137), .ZN(n12113) );
  INV_X1 U10701 ( .A(n12113), .ZN(n10847) );
  NAND2_X1 U10702 ( .A1(n10846), .A2(n10847), .ZN(n10845) );
  OR2_X1 U10703 ( .A1(n11919), .A2(n13137), .ZN(n8231) );
  NAND2_X1 U10704 ( .A1(n10845), .A2(n8231), .ZN(n8232) );
  NAND2_X1 U10705 ( .A1(n11932), .A2(n13136), .ZN(n8233) );
  NAND2_X1 U10706 ( .A1(n13477), .A2(n13135), .ZN(n8234) );
  NAND2_X1 U10707 ( .A1(n8235), .A2(n8234), .ZN(n11278) );
  NAND2_X1 U10708 ( .A1(n11946), .A2(n13134), .ZN(n8236) );
  AND2_X1 U10709 ( .A1(n11953), .A2(n13133), .ZN(n8237) );
  NOR2_X1 U10710 ( .A1(n11961), .A2(n13131), .ZN(n8238) );
  OR2_X1 U10711 ( .A1(n11969), .A2(n13130), .ZN(n8239) );
  NAND2_X1 U10712 ( .A1(n11601), .A2(n8239), .ZN(n8241) );
  NAND2_X1 U10713 ( .A1(n11969), .A2(n13130), .ZN(n8240) );
  NOR2_X1 U10714 ( .A1(n11968), .A2(n11967), .ZN(n8242) );
  NAND2_X1 U10715 ( .A1(n11968), .A2(n11967), .ZN(n8243) );
  OR2_X1 U10716 ( .A1(n13617), .A2(n13128), .ZN(n8244) );
  NAND2_X1 U10717 ( .A1(n8245), .A2(n8244), .ZN(n13448) );
  XNOR2_X1 U10718 ( .A(n13551), .B(n13127), .ZN(n13452) );
  NAND2_X1 U10720 ( .A1(n13551), .A2(n13127), .ZN(n8246) );
  NAND2_X1 U10721 ( .A1(n11978), .A2(n13126), .ZN(n8247) );
  XNOR2_X1 U10722 ( .A(n13541), .B(n13028), .ZN(n13411) );
  INV_X1 U10723 ( .A(n13411), .ZN(n13424) );
  NAND2_X1 U10724 ( .A1(n13537), .A2(n13125), .ZN(n12128) );
  NAND2_X1 U10725 ( .A1(n13399), .A2(n12128), .ZN(n8248) );
  OR2_X1 U10726 ( .A1(n13537), .A2(n13125), .ZN(n12129) );
  OR2_X1 U10727 ( .A1(n13603), .A2(n12023), .ZN(n8249) );
  NAND2_X1 U10728 ( .A1(n13526), .A2(n13123), .ZN(n12101) );
  INV_X1 U10729 ( .A(n12101), .ZN(n8250) );
  NAND2_X1 U10730 ( .A1(n13376), .A2(n13059), .ZN(n12102) );
  NAND2_X1 U10731 ( .A1(n13591), .A2(n13122), .ZN(n8252) );
  NAND2_X1 U10732 ( .A1(n13328), .A2(n8253), .ZN(n8255) );
  NAND2_X1 U10733 ( .A1(n13331), .A2(n13120), .ZN(n8254) );
  NOR2_X1 U10734 ( .A1(n13320), .A2(n13093), .ZN(n8256) );
  NAND2_X1 U10735 ( .A1(n13320), .A2(n13093), .ZN(n8257) );
  NOR2_X1 U10736 ( .A1(n13500), .A2(n13119), .ZN(n8258) );
  INV_X1 U10737 ( .A(n13500), .ZN(n13102) );
  NOR2_X1 U10738 ( .A1(n13286), .A2(n13095), .ZN(n8259) );
  AOI21_X1 U10739 ( .B1(n13281), .B2(n13280), .A(n8259), .ZN(n13262) );
  INV_X1 U10740 ( .A(n13489), .ZN(n13276) );
  OAI22_X1 U10741 ( .A1(n13262), .A2(n13266), .B1(n9793), .B2(n13276), .ZN(
        n8260) );
  XNOR2_X1 U10742 ( .A(n8260), .B(n12134), .ZN(n9664) );
  NAND2_X1 U10743 ( .A1(n14864), .A2(n14850), .ZN(n13561) );
  INV_X1 U10744 ( .A(n9664), .ZN(n8270) );
  NOR2_X1 U10745 ( .A1(n14834), .A2(n8265), .ZN(n9785) );
  NAND3_X1 U10746 ( .A1(n9785), .A2(n12146), .A3(n14831), .ZN(n8267) );
  INV_X1 U10747 ( .A(n9796), .ZN(n8266) );
  NAND2_X2 U10748 ( .A1(n8267), .A2(n13472), .ZN(n13468) );
  AND2_X1 U10749 ( .A1(n12090), .A2(n8221), .ZN(n8268) );
  NAND2_X1 U10750 ( .A1(n13468), .A2(n8268), .ZN(n13279) );
  INV_X1 U10751 ( .A(n9668), .ZN(n13271) );
  NAND2_X1 U10752 ( .A1(n13468), .A2(n13271), .ZN(n8269) );
  NAND2_X1 U10753 ( .A1(n13468), .A2(n13249), .ZN(n13350) );
  NOR2_X1 U10754 ( .A1(n8271), .A2(n13350), .ZN(n8276) );
  OR2_X1 U10755 ( .A1(n10141), .A2(n8222), .ZN(n9791) );
  INV_X1 U10756 ( .A(n9791), .ZN(n8272) );
  INV_X1 U10757 ( .A(n13472), .ZN(n13419) );
  AOI22_X1 U10758 ( .A1(n8273), .A2(n13419), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n13428), .ZN(n8274) );
  OAI21_X1 U10759 ( .B1(n12060), .B2(n13463), .A(n8274), .ZN(n8275) );
  NOR2_X1 U10760 ( .A1(n8276), .A2(n8275), .ZN(n8277) );
  NOR2_X1 U10761 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8286) );
  NOR2_X1 U10762 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), 
        .ZN(n8292) );
  NOR2_X1 U10763 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .ZN(n8291) );
  INV_X2 U10764 ( .A(n8408), .ZN(n8797) );
  NAND2_X1 U10765 ( .A1(n8797), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8299) );
  NAND2_X1 U10766 ( .A1(n8769), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8314) );
  NAND2_X1 U10767 ( .A1(n8419), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8313) );
  AND2_X2 U10768 ( .A1(n8305), .A2(n8310), .ZN(n8654) );
  INV_X1 U10769 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n15301) );
  INV_X1 U10770 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n15165) );
  NAND2_X1 U10771 ( .A1(n8420), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8438) );
  NOR2_X1 U10772 ( .A1(n8438), .A2(n8437), .ZN(n8450) );
  NAND2_X1 U10773 ( .A1(n8450), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U10774 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n8306) );
  AND2_X1 U10775 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_REG3_REG_14__SCAN_IN), 
        .ZN(n8307) );
  NAND2_X1 U10776 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n8308) );
  INV_X1 U10777 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8640) );
  NAND2_X1 U10778 ( .A1(n8666), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8679) );
  AOI21_X1 U10779 ( .B1(n15301), .B2(n8309), .A(n8691), .ZN(n13980) );
  NAND2_X1 U10780 ( .A1(n8754), .A2(n13980), .ZN(n8312) );
  NAND2_X1 U10781 ( .A1(n8784), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8311) );
  NAND4_X1 U10782 ( .A1(n8314), .A2(n8313), .A3(n8312), .A4(n8311), .ZN(n13958) );
  AND2_X1 U10783 ( .A1(n8562), .A2(n8315), .ZN(n8590) );
  NAND2_X1 U10784 ( .A1(n8590), .A2(n8316), .ZN(n8599) );
  NAND2_X1 U10785 ( .A1(n8327), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U10786 ( .A1(n8329), .A2(n11492), .ZN(n8803) );
  NAND2_X1 U10787 ( .A1(n7279), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8326) );
  MUX2_X1 U10788 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8326), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n8328) );
  NAND2_X1 U10789 ( .A1(n8328), .A2(n8327), .ZN(n11378) );
  INV_X1 U10790 ( .A(n11378), .ZN(n8847) );
  NAND2_X1 U10791 ( .A1(n10242), .A2(n8847), .ZN(n10249) );
  NAND2_X1 U10792 ( .A1(n8803), .A2(n10249), .ZN(n8783) );
  NAND2_X1 U10793 ( .A1(n8329), .A2(n8847), .ZN(n8330) );
  NAND2_X2 U10794 ( .A1(n8783), .A2(n8330), .ZN(n8349) );
  MUX2_X1 U10795 ( .A(n8838), .B(n13958), .S(n8806), .Z(n8688) );
  NAND2_X1 U10796 ( .A1(n8369), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n8333) );
  NAND2_X1 U10797 ( .A1(n8654), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n8332) );
  NAND2_X1 U10798 ( .A1(n8386), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n8334) );
  INV_X1 U10799 ( .A(SI_0_), .ZN(n8335) );
  INV_X1 U10800 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9043) );
  OAI21_X1 U10801 ( .B1(n9831), .B2(n8335), .A(n9043), .ZN(n8336) );
  AND2_X1 U10802 ( .A1(n8337), .A2(n8336), .ZN(n14208) );
  NAND2_X1 U10803 ( .A1(n14627), .A2(n14623), .ZN(n10695) );
  XNOR2_X1 U10804 ( .A(n10695), .B(n8349), .ZN(n8348) );
  NAND2_X1 U10805 ( .A1(n8386), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8339) );
  INV_X1 U10806 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n8338) );
  NAND2_X1 U10807 ( .A1(n8369), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8341) );
  NAND2_X1 U10808 ( .A1(n8654), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n8340) );
  INV_X1 U10809 ( .A(n8342), .ZN(n9832) );
  NAND2_X1 U10810 ( .A1(n6825), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8346) );
  NAND2_X1 U10811 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n14207), .ZN(n8344) );
  NAND2_X1 U10812 ( .A1(n8637), .A2(n10013), .ZN(n8345) );
  OAI21_X1 U10813 ( .B1(n13813), .B2(n14623), .A(n14630), .ZN(n10251) );
  NAND2_X1 U10814 ( .A1(n10251), .A2(n10281), .ZN(n8347) );
  NAND3_X1 U10815 ( .A1(n8348), .A2(n10686), .A3(n8347), .ZN(n8353) );
  NAND2_X1 U10816 ( .A1(n6863), .A2(n8349), .ZN(n8351) );
  INV_X1 U10817 ( .A(n10357), .ZN(n14626) );
  NAND2_X1 U10818 ( .A1(n14626), .A2(n8800), .ZN(n8350) );
  MUX2_X1 U10819 ( .A(n8351), .B(n8350), .S(n10689), .Z(n8352) );
  NAND2_X1 U10820 ( .A1(n8353), .A2(n8352), .ZN(n8367) );
  NAND2_X1 U10821 ( .A1(n8654), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n8358) );
  NAND2_X1 U10822 ( .A1(n8386), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8357) );
  INV_X1 U10823 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10012) );
  INV_X1 U10824 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n8354) );
  INV_X2 U10825 ( .A(n8359), .ZN(n8474) );
  NAND2_X1 U10826 ( .A1(n8474), .A2(n9847), .ZN(n8363) );
  NAND2_X1 U10827 ( .A1(n8637), .A2(n10343), .ZN(n8362) );
  NAND2_X1 U10828 ( .A1(n8800), .A2(n10694), .ZN(n8364) );
  NAND2_X1 U10829 ( .A1(n8827), .A2(n8364), .ZN(n8365) );
  NAND2_X1 U10830 ( .A1(n8367), .A2(n8366), .ZN(n8379) );
  NAND2_X1 U10831 ( .A1(n8419), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8373) );
  INV_X1 U10832 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8368) );
  NAND2_X1 U10833 ( .A1(n8654), .A2(n8368), .ZN(n8372) );
  NAND2_X1 U10834 ( .A1(n8386), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8371) );
  NAND2_X1 U10835 ( .A1(n8369), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8370) );
  NAND2_X1 U10836 ( .A1(n8374), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8376) );
  INV_X1 U10837 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8375) );
  XNOR2_X1 U10838 ( .A(n8376), .B(n8375), .ZN(n13814) );
  NAND2_X1 U10839 ( .A1(n9855), .A2(n8474), .ZN(n8378) );
  NAND2_X1 U10840 ( .A1(n6825), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8377) );
  OAI211_X1 U10841 ( .C1(n8343), .C2(n13814), .A(n8378), .B(n8377), .ZN(n14562) );
  NAND3_X1 U10842 ( .A1(n8380), .A2(n8379), .A3(n10820), .ZN(n8384) );
  NAND2_X1 U10843 ( .A1(n8349), .A2(n14562), .ZN(n8382) );
  INV_X1 U10844 ( .A(n14562), .ZN(n10817) );
  NAND2_X1 U10845 ( .A1(n8800), .A2(n10817), .ZN(n8381) );
  MUX2_X1 U10846 ( .A(n8382), .B(n8381), .S(n13811), .Z(n8383) );
  NAND2_X1 U10847 ( .A1(n8384), .A2(n8383), .ZN(n8396) );
  NAND2_X1 U10848 ( .A1(n8769), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8390) );
  NAND2_X1 U10849 ( .A1(n8419), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n8389) );
  INV_X1 U10850 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n8385) );
  XNOR2_X1 U10851 ( .A(n8385), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n10938) );
  NAND2_X1 U10852 ( .A1(n8754), .A2(n10938), .ZN(n8388) );
  NAND2_X1 U10853 ( .A1(n8784), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8387) );
  NAND4_X1 U10854 ( .A1(n8390), .A2(n8389), .A3(n8388), .A4(n8387), .ZN(n13810) );
  NAND2_X1 U10855 ( .A1(n9857), .A2(n8745), .ZN(n8393) );
  OR2_X1 U10856 ( .A1(n8374), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n8409) );
  NAND2_X1 U10857 ( .A1(n8409), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8391) );
  XNOR2_X1 U10858 ( .A(n8391), .B(P1_IR_REG_4__SCAN_IN), .ZN(n13832) );
  AOI22_X1 U10859 ( .A1(n8797), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n8637), .B2(
        n13832), .ZN(n8392) );
  MUX2_X1 U10860 ( .A(n13810), .B(n10949), .S(n8349), .Z(n8397) );
  NAND2_X1 U10861 ( .A1(n8396), .A2(n8397), .ZN(n8395) );
  MUX2_X1 U10862 ( .A(n13810), .B(n10949), .S(n8800), .Z(n8394) );
  NAND2_X1 U10863 ( .A1(n8395), .A2(n8394), .ZN(n8401) );
  INV_X1 U10864 ( .A(n8396), .ZN(n8399) );
  INV_X1 U10865 ( .A(n8397), .ZN(n8398) );
  AOI21_X1 U10866 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8402) );
  NOR2_X1 U10867 ( .A1(n8402), .A2(n8420), .ZN(n10871) );
  NAND2_X1 U10868 ( .A1(n8754), .A2(n10871), .ZN(n8407) );
  NAND2_X1 U10869 ( .A1(n8784), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n8406) );
  INV_X1 U10870 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n8403) );
  OR2_X1 U10871 ( .A1(n8788), .A2(n8403), .ZN(n8405) );
  INV_X1 U10872 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10869) );
  OR2_X1 U10873 ( .A1(n8779), .A2(n10869), .ZN(n8404) );
  INV_X1 U10874 ( .A(n11017), .ZN(n13809) );
  NAND2_X1 U10875 ( .A1(n9861), .A2(n8474), .ZN(n8416) );
  NOR2_X1 U10876 ( .A1(n8409), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n8413) );
  INV_X1 U10877 ( .A(n8413), .ZN(n8410) );
  NAND2_X1 U10878 ( .A1(n8410), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8411) );
  MUX2_X1 U10879 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8411), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n8414) );
  NAND2_X1 U10880 ( .A1(n8413), .A2(n8412), .ZN(n8444) );
  AOI22_X1 U10881 ( .A1(n8797), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8637), .B2(
        n10055), .ZN(n8415) );
  NAND2_X1 U10882 ( .A1(n8416), .A2(n8415), .ZN(n11019) );
  MUX2_X1 U10883 ( .A(n13809), .B(n11019), .S(n8800), .Z(n8418) );
  MUX2_X1 U10884 ( .A(n13809), .B(n11019), .S(n8349), .Z(n8417) );
  NAND2_X1 U10885 ( .A1(n8769), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8425) );
  NAND2_X1 U10886 ( .A1(n8419), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n8424) );
  OAI21_X1 U10887 ( .B1(n8420), .B2(P1_REG3_REG_6__SCAN_IN), .A(n8438), .ZN(
        n14609) );
  INV_X1 U10888 ( .A(n14609), .ZN(n8421) );
  NAND2_X1 U10889 ( .A1(n8654), .A2(n8421), .ZN(n8423) );
  NAND2_X1 U10890 ( .A1(n8784), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8422) );
  NAND4_X1 U10891 ( .A1(n8425), .A2(n8424), .A3(n8423), .A4(n8422), .ZN(n13808) );
  NAND2_X1 U10892 ( .A1(n9873), .A2(n8474), .ZN(n8428) );
  NAND2_X1 U10893 ( .A1(n8444), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8426) );
  XNOR2_X1 U10894 ( .A(n8426), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10188) );
  AOI22_X1 U10895 ( .A1(n8797), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8637), .B2(
        n10188), .ZN(n8427) );
  NAND2_X1 U10896 ( .A1(n8428), .A2(n8427), .ZN(n14612) );
  MUX2_X1 U10897 ( .A(n13808), .B(n14612), .S(n8349), .Z(n8432) );
  NAND2_X1 U10898 ( .A1(n8431), .A2(n8432), .ZN(n8430) );
  MUX2_X1 U10899 ( .A(n13808), .B(n14612), .S(n8800), .Z(n8429) );
  NAND2_X1 U10900 ( .A1(n8430), .A2(n8429), .ZN(n8436) );
  INV_X1 U10901 ( .A(n8431), .ZN(n8434) );
  INV_X1 U10902 ( .A(n8432), .ZN(n8433) );
  NAND2_X1 U10903 ( .A1(n8434), .A2(n8433), .ZN(n8435) );
  NAND2_X1 U10904 ( .A1(n8769), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8443) );
  NAND2_X1 U10905 ( .A1(n8419), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8442) );
  AND2_X1 U10906 ( .A1(n8438), .A2(n8437), .ZN(n8439) );
  NOR2_X1 U10907 ( .A1(n8450), .A2(n8439), .ZN(n11197) );
  NAND2_X1 U10908 ( .A1(n8754), .A2(n11197), .ZN(n8441) );
  NAND2_X1 U10909 ( .A1(n8784), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8440) );
  NAND4_X1 U10910 ( .A1(n8443), .A2(n8442), .A3(n8441), .A4(n8440), .ZN(n13807) );
  NAND2_X1 U10911 ( .A1(n9877), .A2(n8474), .ZN(n8447) );
  OAI21_X1 U10912 ( .B1(n8444), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8445) );
  XNOR2_X1 U10913 ( .A(n8445), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10159) );
  AOI22_X1 U10914 ( .A1(n8797), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8637), .B2(
        n10159), .ZN(n8446) );
  NAND2_X1 U10915 ( .A1(n8447), .A2(n8446), .ZN(n11193) );
  MUX2_X1 U10916 ( .A(n13807), .B(n11193), .S(n8800), .Z(n8448) );
  MUX2_X1 U10917 ( .A(n13807), .B(n11193), .S(n8349), .Z(n8449) );
  NAND2_X1 U10918 ( .A1(n8769), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8455) );
  NAND2_X1 U10919 ( .A1(n8419), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8454) );
  OR2_X1 U10920 ( .A1(n8450), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8451) );
  AND2_X1 U10921 ( .A1(n8467), .A2(n8451), .ZN(n11419) );
  NAND2_X1 U10922 ( .A1(n8754), .A2(n11419), .ZN(n8453) );
  NAND2_X1 U10923 ( .A1(n8784), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8452) );
  NAND4_X1 U10924 ( .A1(n8455), .A2(n8454), .A3(n8453), .A4(n8452), .ZN(n13806) );
  NAND2_X1 U10925 ( .A1(n9880), .A2(n8474), .ZN(n8459) );
  NAND2_X1 U10926 ( .A1(n8456), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8457) );
  XNOR2_X1 U10927 ( .A(n8457), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10102) );
  AOI22_X1 U10928 ( .A1(n8797), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8637), .B2(
        n10102), .ZN(n8458) );
  NAND2_X1 U10929 ( .A1(n8459), .A2(n8458), .ZN(n14717) );
  MUX2_X1 U10930 ( .A(n13806), .B(n14717), .S(n8349), .Z(n8462) );
  MUX2_X1 U10931 ( .A(n13806), .B(n14717), .S(n8800), .Z(n8460) );
  NAND2_X1 U10932 ( .A1(n8461), .A2(n8460), .ZN(n8465) );
  INV_X1 U10933 ( .A(n8462), .ZN(n8463) );
  NAND2_X1 U10934 ( .A1(n6528), .A2(n8463), .ZN(n8464) );
  NAND2_X1 U10935 ( .A1(n8784), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8473) );
  NAND2_X1 U10936 ( .A1(n8467), .A2(n8466), .ZN(n8468) );
  AND2_X1 U10937 ( .A1(n8484), .A2(n8468), .ZN(n11561) );
  NAND2_X1 U10938 ( .A1(n8654), .A2(n11561), .ZN(n8472) );
  INV_X1 U10939 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10107) );
  OR2_X1 U10940 ( .A1(n8779), .A2(n10107), .ZN(n8471) );
  INV_X1 U10941 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n8469) );
  OR2_X1 U10942 ( .A1(n8788), .A2(n8469), .ZN(n8470) );
  INV_X1 U10943 ( .A(n11553), .ZN(n13805) );
  NAND2_X1 U10944 ( .A1(n9884), .A2(n8474), .ZN(n8481) );
  NOR2_X1 U10945 ( .A1(n8456), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n8477) );
  NOR2_X1 U10946 ( .A1(n8477), .A2(n8589), .ZN(n8475) );
  MUX2_X1 U10947 ( .A(n8589), .B(n8475), .S(P1_IR_REG_9__SCAN_IN), .Z(n8479)
         );
  INV_X1 U10948 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8476) );
  NAND2_X1 U10949 ( .A1(n8477), .A2(n8476), .ZN(n8511) );
  INV_X1 U10950 ( .A(n8511), .ZN(n8478) );
  NOR2_X1 U10951 ( .A1(n8479), .A2(n8478), .ZN(n10209) );
  AOI22_X1 U10952 ( .A1(n8797), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8637), .B2(
        n10209), .ZN(n8480) );
  NAND2_X1 U10953 ( .A1(n8481), .A2(n8480), .ZN(n14739) );
  MUX2_X1 U10954 ( .A(n13805), .B(n14739), .S(n8800), .Z(n8483) );
  MUX2_X1 U10955 ( .A(n13805), .B(n14739), .S(n8806), .Z(n8482) );
  NAND2_X1 U10956 ( .A1(n8484), .A2(n10214), .ZN(n8485) );
  NAND2_X1 U10957 ( .A1(n8518), .A2(n8485), .ZN(n14503) );
  INV_X1 U10958 ( .A(n14503), .ZN(n8486) );
  NAND2_X1 U10959 ( .A1(n8754), .A2(n8486), .ZN(n8492) );
  NAND2_X1 U10960 ( .A1(n8784), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8491) );
  INV_X1 U10961 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n8487) );
  OR2_X1 U10962 ( .A1(n8788), .A2(n8487), .ZN(n8490) );
  INV_X1 U10963 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n8488) );
  OR2_X1 U10964 ( .A1(n8779), .A2(n8488), .ZN(n8489) );
  INV_X1 U10965 ( .A(n11828), .ZN(n14509) );
  NAND2_X1 U10966 ( .A1(n9924), .A2(n8745), .ZN(n8495) );
  NAND2_X1 U10967 ( .A1(n8511), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8493) );
  XNOR2_X1 U10968 ( .A(n8493), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10295) );
  AOI22_X1 U10969 ( .A1(n8797), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8637), 
        .B2(n10295), .ZN(n8494) );
  MUX2_X1 U10970 ( .A(n14509), .B(n14491), .S(n8349), .Z(n8499) );
  NAND2_X1 U10971 ( .A1(n8498), .A2(n8499), .ZN(n8497) );
  MUX2_X1 U10972 ( .A(n14509), .B(n14491), .S(n8800), .Z(n8496) );
  NAND2_X1 U10973 ( .A1(n8497), .A2(n8496), .ZN(n8503) );
  INV_X1 U10974 ( .A(n8498), .ZN(n8501) );
  INV_X1 U10975 ( .A(n8499), .ZN(n8500) );
  NAND2_X1 U10976 ( .A1(n8501), .A2(n8500), .ZN(n8502) );
  NAND2_X1 U10977 ( .A1(n8503), .A2(n8502), .ZN(n8517) );
  INV_X1 U10978 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8504) );
  XNOR2_X1 U10979 ( .A(n8518), .B(n8504), .ZN(n14518) );
  INV_X1 U10980 ( .A(n14518), .ZN(n8505) );
  NAND2_X1 U10981 ( .A1(n8754), .A2(n8505), .ZN(n8510) );
  NAND2_X1 U10982 ( .A1(n8784), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8509) );
  INV_X1 U10983 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n8506) );
  OR2_X1 U10984 ( .A1(n8788), .A2(n8506), .ZN(n8508) );
  INV_X1 U10985 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11334) );
  OR2_X1 U10986 ( .A1(n8779), .A2(n11334), .ZN(n8507) );
  NAND2_X1 U10987 ( .A1(n9958), .A2(n8745), .ZN(n8514) );
  NAND2_X1 U10988 ( .A1(n8527), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8512) );
  XNOR2_X1 U10989 ( .A(n8512), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10790) );
  AOI22_X1 U10990 ( .A1(n8797), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8637), 
        .B2(n10790), .ZN(n8513) );
  NAND2_X1 U10991 ( .A1(n8514), .A2(n8513), .ZN(n11835) );
  MUX2_X1 U10992 ( .A(n13804), .B(n11835), .S(n8800), .Z(n8516) );
  INV_X1 U10993 ( .A(n11835), .ZN(n14532) );
  MUX2_X1 U10994 ( .A(n11833), .B(n14532), .S(n8806), .Z(n8515) );
  AOI21_X1 U10995 ( .B1(n8517), .B2(n8516), .A(n8515), .ZN(n8531) );
  NOR2_X1 U10996 ( .A1(n8517), .A2(n8516), .ZN(n8530) );
  INV_X1 U10997 ( .A(n8518), .ZN(n8519) );
  AOI21_X1 U10998 ( .B1(n8519), .B2(P1_REG3_REG_11__SCAN_IN), .A(
        P1_REG3_REG_12__SCAN_IN), .ZN(n8520) );
  NAND2_X1 U10999 ( .A1(n8654), .A2(n7566), .ZN(n8526) );
  NAND2_X1 U11000 ( .A1(n8784), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8525) );
  INV_X1 U11001 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n8521) );
  OR2_X1 U11002 ( .A1(n8779), .A2(n8521), .ZN(n8524) );
  INV_X1 U11003 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n8522) );
  OR2_X1 U11004 ( .A1(n8788), .A2(n8522), .ZN(n8523) );
  NAND2_X1 U11005 ( .A1(n9962), .A2(n8745), .ZN(n8529) );
  OAI21_X1 U11006 ( .B1(n8527), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8541) );
  XNOR2_X1 U11007 ( .A(n8541), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10795) );
  AOI22_X1 U11008 ( .A1(n8797), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n8637), 
        .B2(n10795), .ZN(n8528) );
  MUX2_X1 U11009 ( .A(n11843), .B(n11851), .S(n8800), .Z(n8546) );
  INV_X1 U11010 ( .A(n11843), .ZN(n14511) );
  MUX2_X1 U11011 ( .A(n14511), .B(n11616), .S(n8806), .Z(n8545) );
  OAI22_X1 U11012 ( .A1(n8531), .A2(n8530), .B1(n8546), .B2(n8545), .ZN(n8561)
         );
  NOR2_X1 U11013 ( .A1(n8532), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8533) );
  OR2_X1 U11014 ( .A1(n8566), .A2(n8533), .ZN(n14340) );
  INV_X1 U11015 ( .A(n14340), .ZN(n8534) );
  NAND2_X1 U11016 ( .A1(n8654), .A2(n8534), .ZN(n8539) );
  NAND2_X1 U11017 ( .A1(n8784), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8538) );
  INV_X1 U11018 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10797) );
  OR2_X1 U11019 ( .A1(n8779), .A2(n10797), .ZN(n8537) );
  INV_X1 U11020 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n8535) );
  OR2_X1 U11021 ( .A1(n8788), .A2(n8535), .ZN(n8536) );
  NAND2_X1 U11022 ( .A1(n9969), .A2(n8745), .ZN(n8544) );
  NAND2_X1 U11023 ( .A1(n8541), .A2(n8540), .ZN(n8542) );
  NAND2_X1 U11024 ( .A1(n8542), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8549) );
  XNOR2_X1 U11025 ( .A(n8549), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11269) );
  AOI22_X1 U11026 ( .A1(n8797), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n8637), 
        .B2(n11269), .ZN(n8543) );
  MUX2_X1 U11027 ( .A(n12206), .B(n14526), .S(n8800), .Z(n8574) );
  INV_X1 U11028 ( .A(n12206), .ZN(n14483) );
  MUX2_X1 U11029 ( .A(n14483), .B(n14343), .S(n8806), .Z(n8547) );
  AOI22_X1 U11030 ( .A1(n8574), .A2(n8547), .B1(n8546), .B2(n8545), .ZN(n8560)
         );
  NAND2_X1 U11031 ( .A1(n10257), .A2(n8745), .ZN(n8553) );
  INV_X1 U11032 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U11033 ( .A1(n8549), .A2(n8548), .ZN(n8550) );
  NAND2_X1 U11034 ( .A1(n8550), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8551) );
  XNOR2_X1 U11035 ( .A(n8551), .B(P1_IR_REG_14__SCAN_IN), .ZN(n13846) );
  AOI22_X1 U11036 ( .A1(n13846), .A2(n8637), .B1(n8797), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8552) );
  XNOR2_X1 U11037 ( .A(n8566), .B(P1_REG3_REG_14__SCAN_IN), .ZN(n14490) );
  INV_X1 U11038 ( .A(n14490), .ZN(n8554) );
  NAND2_X1 U11039 ( .A1(n8754), .A2(n8554), .ZN(n8559) );
  NAND2_X1 U11040 ( .A1(n8784), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8558) );
  INV_X1 U11041 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11594) );
  OR2_X1 U11042 ( .A1(n8779), .A2(n11594), .ZN(n8557) );
  INV_X1 U11043 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n8555) );
  OR2_X1 U11044 ( .A1(n8788), .A2(n8555), .ZN(n8556) );
  XNOR2_X1 U11045 ( .A(n12214), .B(n13753), .ZN(n11591) );
  INV_X1 U11046 ( .A(n12214), .ZN(n14520) );
  INV_X1 U11047 ( .A(n13753), .ZN(n14338) );
  NAND2_X1 U11048 ( .A1(n10423), .A2(n8745), .ZN(n8565) );
  OR2_X1 U11049 ( .A1(n8562), .A2(n8589), .ZN(n8563) );
  XNOR2_X1 U11050 ( .A(n8563), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U11051 ( .A1(n8797), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8637), 
        .B2(n11504), .ZN(n8564) );
  AOI21_X1 U11052 ( .B1(n8566), .B2(P1_REG3_REG_14__SCAN_IN), .A(
        P1_REG3_REG_15__SCAN_IN), .ZN(n8567) );
  OR2_X1 U11053 ( .A1(n8582), .A2(n8567), .ZN(n11631) );
  INV_X1 U11054 ( .A(n11631), .ZN(n13795) );
  NAND2_X1 U11055 ( .A1(n8754), .A2(n13795), .ZN(n8573) );
  NAND2_X1 U11056 ( .A1(n8784), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n8572) );
  INV_X1 U11057 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n8568) );
  OR2_X1 U11058 ( .A1(n8788), .A2(n8568), .ZN(n8571) );
  INV_X1 U11059 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8569) );
  OR2_X1 U11060 ( .A1(n8779), .A2(n8569), .ZN(n8570) );
  NAND2_X1 U11061 ( .A1(n12222), .A2(n12226), .ZN(n8826) );
  OAI21_X1 U11062 ( .B1(n14520), .B2(n14338), .A(n8826), .ZN(n8579) );
  INV_X1 U11063 ( .A(n8574), .ZN(n8577) );
  AND2_X1 U11064 ( .A1(n8800), .A2(n14483), .ZN(n8575) );
  AOI21_X1 U11065 ( .B1(n14343), .B2(n8806), .A(n8575), .ZN(n8576) );
  AND2_X1 U11066 ( .A1(n8577), .A2(n8576), .ZN(n8578) );
  AOI22_X1 U11067 ( .A1(n8579), .A2(n8800), .B1(n8578), .B2(n11627), .ZN(n8581) );
  INV_X1 U11068 ( .A(n11721), .ZN(n8580) );
  OR2_X1 U11069 ( .A1(n12214), .A2(n13753), .ZN(n11625) );
  AOI21_X1 U11070 ( .B1(n11721), .B2(n11625), .A(n8800), .ZN(n8610) );
  OR2_X1 U11071 ( .A1(n8582), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8583) );
  AND2_X1 U11072 ( .A1(n8583), .A2(n8616), .ZN(n13712) );
  NAND2_X1 U11073 ( .A1(n8654), .A2(n13712), .ZN(n8588) );
  NAND2_X1 U11074 ( .A1(n8784), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8587) );
  INV_X1 U11075 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11737) );
  OR2_X1 U11076 ( .A1(n8779), .A2(n11737), .ZN(n8586) );
  INV_X1 U11077 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n8584) );
  OR2_X1 U11078 ( .A1(n8788), .A2(n8584), .ZN(n8585) );
  NAND2_X1 U11079 ( .A1(n10527), .A2(n8745), .ZN(n8593) );
  OR2_X1 U11080 ( .A1(n8590), .A2(n8589), .ZN(n8591) );
  XNOR2_X1 U11081 ( .A(n8591), .B(P1_IR_REG_16__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U11082 ( .A1(n8797), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8637), 
        .B2(n11700), .ZN(n8592) );
  MUX2_X1 U11083 ( .A(n13803), .B(n12232), .S(n8800), .Z(n8632) );
  XNOR2_X1 U11084 ( .A(n8616), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n13720) );
  NAND2_X1 U11085 ( .A1(n8754), .A2(n13720), .ZN(n8598) );
  NAND2_X1 U11086 ( .A1(n8784), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8597) );
  INV_X1 U11087 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n8594) );
  OR2_X1 U11088 ( .A1(n8788), .A2(n8594), .ZN(n8596) );
  INV_X1 U11089 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n13868) );
  OR2_X1 U11090 ( .A1(n8779), .A2(n13868), .ZN(n8595) );
  NAND2_X1 U11091 ( .A1(n8632), .A2(n14052), .ZN(n8603) );
  NAND2_X1 U11092 ( .A1(n13792), .A2(n8800), .ZN(n8623) );
  NAND2_X1 U11093 ( .A1(n10586), .A2(n8745), .ZN(n8602) );
  NAND2_X1 U11094 ( .A1(n8599), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8600) );
  XNOR2_X1 U11095 ( .A(n8600), .B(P1_IR_REG_17__SCAN_IN), .ZN(n13862) );
  AOI22_X1 U11096 ( .A1(n8797), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8637), 
        .B2(n13862), .ZN(n8601) );
  INV_X1 U11097 ( .A(n14150), .ZN(n11819) );
  AOI21_X1 U11098 ( .B1(n8603), .B2(n8623), .A(n11819), .ZN(n8608) );
  NAND2_X1 U11099 ( .A1(n8632), .A2(n8824), .ZN(n8604) );
  OR2_X1 U11100 ( .A1(n12232), .A2(n8800), .ZN(n8630) );
  AOI21_X1 U11101 ( .B1(n8604), .B2(n8630), .A(n14150), .ZN(n8607) );
  NAND2_X1 U11102 ( .A1(n14052), .A2(n8806), .ZN(n8633) );
  OR2_X1 U11103 ( .A1(n12232), .A2(n8633), .ZN(n8606) );
  NAND3_X1 U11104 ( .A1(n13792), .A2(n8824), .A3(n8800), .ZN(n8605) );
  NAND2_X1 U11105 ( .A1(n8606), .A2(n8605), .ZN(n8627) );
  OR3_X1 U11106 ( .A1(n8608), .A2(n8607), .A3(n8627), .ZN(n8609) );
  OR2_X1 U11107 ( .A1(n10966), .A2(n8359), .ZN(n8614) );
  NAND2_X1 U11108 ( .A1(n8611), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8612) );
  XNOR2_X1 U11109 ( .A(n8612), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13880) );
  AOI22_X1 U11110 ( .A1(n8797), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8637), 
        .B2(n13880), .ZN(n8613) );
  INV_X1 U11111 ( .A(n14144), .ZN(n14064) );
  INV_X1 U11112 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11696) );
  INV_X1 U11113 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8615) );
  OAI21_X1 U11114 ( .B1(n8616), .B2(n11696), .A(n8615), .ZN(n8617) );
  AND2_X1 U11115 ( .A1(n8617), .A2(n8641), .ZN(n14061) );
  NAND2_X1 U11116 ( .A1(n14061), .A2(n8654), .ZN(n8622) );
  NAND2_X1 U11117 ( .A1(n8769), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8621) );
  NAND2_X1 U11118 ( .A1(n8784), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8620) );
  INV_X1 U11119 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8618) );
  OR2_X1 U11120 ( .A1(n8779), .A2(n8618), .ZN(n8619) );
  NAND2_X1 U11121 ( .A1(n14064), .A2(n14038), .ZN(n12365) );
  NAND2_X1 U11122 ( .A1(n14144), .A2(n13681), .ZN(n8646) );
  INV_X1 U11123 ( .A(n8623), .ZN(n8624) );
  NAND2_X1 U11124 ( .A1(n8632), .A2(n8624), .ZN(n8625) );
  OAI21_X1 U11125 ( .B1(n14052), .B2(n8806), .A(n8625), .ZN(n8626) );
  NAND2_X1 U11126 ( .A1(n8626), .A2(n14150), .ZN(n8629) );
  NAND2_X1 U11127 ( .A1(n8632), .A2(n8627), .ZN(n8628) );
  NAND4_X1 U11128 ( .A1(n12365), .A2(n8646), .A3(n8629), .A4(n8628), .ZN(n8636) );
  INV_X1 U11129 ( .A(n8630), .ZN(n8631) );
  NAND2_X1 U11130 ( .A1(n8632), .A2(n8631), .ZN(n8634) );
  AOI21_X1 U11131 ( .B1(n8634), .B2(n8633), .A(n14150), .ZN(n8635) );
  NAND2_X1 U11132 ( .A1(n11162), .A2(n8745), .ZN(n8639) );
  AOI22_X1 U11133 ( .A1(n8797), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8637), 
        .B2(n14345), .ZN(n8638) );
  AND2_X1 U11134 ( .A1(n8641), .A2(n8640), .ZN(n8642) );
  OR2_X1 U11135 ( .A1(n8642), .A2(n8652), .ZN(n14040) );
  AOI22_X1 U11136 ( .A1(n8419), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n8784), .B2(
        P1_REG1_REG_19__SCAN_IN), .ZN(n8644) );
  NAND2_X1 U11137 ( .A1(n8769), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8643) );
  OAI211_X1 U11138 ( .C1(n14040), .C2(n8645), .A(n8644), .B(n8643), .ZN(n14051) );
  INV_X1 U11139 ( .A(n14051), .ZN(n13770) );
  NAND2_X1 U11140 ( .A1(n12381), .A2(n13770), .ZN(n12366) );
  AND2_X1 U11141 ( .A1(n12366), .A2(n8646), .ZN(n8647) );
  MUX2_X1 U11142 ( .A(n12365), .B(n8647), .S(n8806), .Z(n8648) );
  OR2_X1 U11143 ( .A1(n12381), .A2(n13770), .ZN(n8823) );
  NAND3_X1 U11144 ( .A1(n8649), .A2(n8648), .A3(n8823), .ZN(n8651) );
  MUX2_X1 U11145 ( .A(n12366), .B(n8823), .S(n8806), .Z(n8650) );
  NAND2_X1 U11146 ( .A1(n8651), .A2(n8650), .ZN(n8661) );
  NOR2_X1 U11147 ( .A1(n8652), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8653) );
  OR2_X1 U11148 ( .A1(n8666), .A2(n8653), .ZN(n14025) );
  AOI22_X1 U11149 ( .A1(n8769), .A2(P1_REG0_REG_20__SCAN_IN), .B1(n8419), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n8656) );
  NAND2_X1 U11150 ( .A1(n8784), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8655) );
  OAI211_X1 U11151 ( .C1(n14025), .C2(n8645), .A(n8656), .B(n8655), .ZN(n14039) );
  INV_X1 U11152 ( .A(n14039), .ZN(n12368) );
  NAND2_X1 U11153 ( .A1(n11360), .A2(n8745), .ZN(n8658) );
  NAND2_X1 U11154 ( .A1(n8797), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8657) );
  INV_X1 U11155 ( .A(n14130), .ZN(n12260) );
  MUX2_X1 U11156 ( .A(n12368), .B(n12260), .S(n8806), .Z(n8660) );
  MUX2_X1 U11157 ( .A(n14039), .B(n14130), .S(n8800), .Z(n8659) );
  OAI21_X1 U11158 ( .B1(n8661), .B2(n8660), .A(n8659), .ZN(n8663) );
  NAND2_X1 U11159 ( .A1(n8661), .A2(n8660), .ZN(n8662) );
  NAND2_X1 U11160 ( .A1(n8663), .A2(n8662), .ZN(n8671) );
  OR2_X1 U11161 ( .A1(n11857), .A2(n8359), .ZN(n8665) );
  NAND2_X1 U11162 ( .A1(n8797), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8664) );
  OR2_X1 U11163 ( .A1(n8666), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U11164 ( .A1(n8667), .A2(n8679), .ZN(n14009) );
  AOI22_X1 U11165 ( .A1(n8769), .A2(P1_REG0_REG_21__SCAN_IN), .B1(n8419), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n8669) );
  NAND2_X1 U11166 ( .A1(n8784), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8668) );
  OAI211_X1 U11167 ( .C1(n14009), .C2(n8645), .A(n8669), .B(n8668), .ZN(n13802) );
  MUX2_X1 U11168 ( .A(n14012), .B(n13802), .S(n8806), .Z(n8670) );
  NAND2_X1 U11169 ( .A1(n8671), .A2(n8670), .ZN(n8674) );
  MUX2_X1 U11170 ( .A(n14012), .B(n13802), .S(n8800), .Z(n8673) );
  NAND2_X1 U11171 ( .A1(n8769), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8683) );
  INV_X1 U11172 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n8677) );
  OR2_X1 U11173 ( .A1(n8779), .A2(n8677), .ZN(n8682) );
  AOI21_X1 U11174 ( .B1(n15165), .B2(n8679), .A(n8678), .ZN(n13994) );
  NAND2_X1 U11175 ( .A1(n8754), .A2(n13994), .ZN(n8681) );
  NAND2_X1 U11176 ( .A1(n8784), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8680) );
  NAND4_X1 U11177 ( .A1(n8683), .A2(n8682), .A3(n8681), .A4(n8680), .ZN(n14004) );
  NAND2_X1 U11178 ( .A1(n8685), .A2(n8684), .ZN(n8686) );
  MUX2_X1 U11179 ( .A(n13958), .B(n8838), .S(n8806), .Z(n8687) );
  NAND2_X1 U11180 ( .A1(n8419), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8696) );
  NAND2_X1 U11181 ( .A1(n8769), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8695) );
  INV_X1 U11182 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8690) );
  INV_X1 U11183 ( .A(n8691), .ZN(n8689) );
  NAND2_X1 U11184 ( .A1(n8690), .A2(n8689), .ZN(n8692) );
  INV_X1 U11185 ( .A(n8707), .ZN(n8709) );
  NAND2_X1 U11186 ( .A1(n8754), .A2(n13967), .ZN(n8694) );
  NAND2_X1 U11187 ( .A1(n8784), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8693) );
  NAND4_X1 U11188 ( .A1(n8696), .A2(n8695), .A3(n8694), .A4(n8693), .ZN(n13943) );
  NAND2_X1 U11189 ( .A1(n13649), .A2(n8745), .ZN(n8698) );
  NAND2_X1 U11190 ( .A1(n8797), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8697) );
  MUX2_X1 U11191 ( .A(n13943), .B(n13964), .S(n8806), .Z(n8702) );
  NAND2_X1 U11192 ( .A1(n8701), .A2(n8702), .ZN(n8700) );
  MUX2_X1 U11193 ( .A(n13943), .B(n13964), .S(n8800), .Z(n8699) );
  NAND2_X1 U11194 ( .A1(n8700), .A2(n8699), .ZN(n8706) );
  INV_X1 U11195 ( .A(n8701), .ZN(n8704) );
  INV_X1 U11196 ( .A(n8702), .ZN(n8703) );
  NAND2_X1 U11197 ( .A1(n8704), .A2(n8703), .ZN(n8705) );
  INV_X1 U11198 ( .A(n8722), .ZN(n8724) );
  INV_X1 U11199 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8708) );
  NAND2_X1 U11200 ( .A1(n8709), .A2(n8708), .ZN(n8710) );
  NAND2_X1 U11201 ( .A1(n8754), .A2(n13945), .ZN(n8716) );
  NAND2_X1 U11202 ( .A1(n8784), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8715) );
  INV_X1 U11203 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n8711) );
  OR2_X1 U11204 ( .A1(n8788), .A2(n8711), .ZN(n8714) );
  INV_X1 U11205 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n8712) );
  OR2_X1 U11206 ( .A1(n8779), .A2(n8712), .ZN(n8713) );
  NAND2_X1 U11207 ( .A1(n11858), .A2(n8745), .ZN(n8718) );
  NAND2_X1 U11208 ( .A1(n8797), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8717) );
  MUX2_X1 U11209 ( .A(n13959), .B(n13940), .S(n8800), .Z(n8720) );
  MUX2_X1 U11210 ( .A(n13959), .B(n13940), .S(n8806), .Z(n8719) );
  INV_X1 U11211 ( .A(n8720), .ZN(n8721) );
  INV_X1 U11212 ( .A(n8737), .ZN(n8739) );
  INV_X1 U11213 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U11214 ( .A1(n8724), .A2(n8723), .ZN(n8725) );
  NAND2_X1 U11215 ( .A1(n8754), .A2(n13924), .ZN(n8731) );
  NAND2_X1 U11216 ( .A1(n8784), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8730) );
  INV_X1 U11217 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n8726) );
  OR2_X1 U11218 ( .A1(n8788), .A2(n8726), .ZN(n8729) );
  INV_X1 U11219 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n8727) );
  OR2_X1 U11220 ( .A1(n8779), .A2(n8727), .ZN(n8728) );
  INV_X1 U11221 ( .A(n13701), .ZN(n13944) );
  NAND2_X1 U11222 ( .A1(n13642), .A2(n8745), .ZN(n8733) );
  NAND2_X1 U11223 ( .A1(n8797), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8732) );
  MUX2_X1 U11224 ( .A(n13944), .B(n13921), .S(n8806), .Z(n8736) );
  MUX2_X1 U11225 ( .A(n13944), .B(n13921), .S(n8800), .Z(n8734) );
  NAND2_X1 U11226 ( .A1(n8769), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8744) );
  NAND2_X1 U11227 ( .A1(n8419), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8743) );
  INV_X1 U11228 ( .A(n8750), .ZN(n8752) );
  INV_X1 U11229 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8738) );
  NAND2_X1 U11230 ( .A1(n8739), .A2(n8738), .ZN(n8740) );
  NAND2_X1 U11231 ( .A1(n8754), .A2(n13662), .ZN(n8742) );
  NAND2_X1 U11232 ( .A1(n8784), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8741) );
  NAND4_X1 U11233 ( .A1(n8744), .A2(n8743), .A3(n8742), .A4(n8741), .ZN(n13801) );
  NAND2_X1 U11234 ( .A1(n13639), .A2(n8745), .ZN(n8747) );
  NAND2_X1 U11235 ( .A1(n8797), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8746) );
  MUX2_X1 U11236 ( .A(n13801), .B(n14087), .S(n8800), .Z(n8749) );
  MUX2_X1 U11237 ( .A(n13801), .B(n14087), .S(n8806), .Z(n8748) );
  INV_X1 U11238 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n15286) );
  OR2_X1 U11239 ( .A1(n8788), .A2(n15286), .ZN(n8758) );
  NAND2_X1 U11240 ( .A1(n8419), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8757) );
  INV_X1 U11241 ( .A(n8770), .ZN(n12385) );
  INV_X1 U11242 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8751) );
  NAND2_X1 U11243 ( .A1(n8752), .A2(n8751), .ZN(n8753) );
  NAND2_X1 U11244 ( .A1(n8754), .A2(n13912), .ZN(n8756) );
  NAND2_X1 U11245 ( .A1(n8784), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8755) );
  NAND4_X1 U11246 ( .A1(n8758), .A2(n8757), .A3(n8756), .A4(n8755), .ZN(n13800) );
  NAND2_X1 U11247 ( .A1(n14193), .A2(n8745), .ZN(n8760) );
  NAND2_X1 U11248 ( .A1(n8797), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8759) );
  MUX2_X1 U11249 ( .A(n13800), .B(n14082), .S(n8806), .Z(n8764) );
  NAND2_X1 U11250 ( .A1(n8763), .A2(n8764), .ZN(n8762) );
  MUX2_X1 U11251 ( .A(n13800), .B(n14082), .S(n8800), .Z(n8761) );
  NAND2_X1 U11252 ( .A1(n8762), .A2(n8761), .ZN(n8768) );
  INV_X1 U11253 ( .A(n8763), .ZN(n8766) );
  INV_X1 U11254 ( .A(n8764), .ZN(n8765) );
  NAND2_X1 U11255 ( .A1(n8769), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8774) );
  NAND2_X1 U11256 ( .A1(n8419), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8773) );
  NAND2_X1 U11257 ( .A1(n8754), .A2(n8770), .ZN(n8772) );
  NAND2_X1 U11258 ( .A1(n8784), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8771) );
  NAND4_X1 U11259 ( .A1(n8774), .A2(n8773), .A3(n8772), .A4(n8771), .ZN(n13799) );
  NAND2_X1 U11260 ( .A1(n8797), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8775) );
  MUX2_X1 U11261 ( .A(n13799), .B(n12382), .S(n8800), .Z(n8777) );
  MUX2_X1 U11262 ( .A(n13799), .B(n12382), .S(n8806), .Z(n8776) );
  INV_X1 U11263 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8782) );
  NAND2_X1 U11264 ( .A1(n8784), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8781) );
  INV_X1 U11265 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8778) );
  OR2_X1 U11266 ( .A1(n8779), .A2(n8778), .ZN(n8780) );
  OAI211_X1 U11267 ( .C1(n8788), .C2(n8782), .A(n8781), .B(n8780), .ZN(n13897)
         );
  INV_X1 U11268 ( .A(n8783), .ZN(n8789) );
  INV_X1 U11269 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n8787) );
  NAND2_X1 U11270 ( .A1(n8419), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8786) );
  NAND2_X1 U11271 ( .A1(n8784), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8785) );
  OAI211_X1 U11272 ( .C1(n8788), .C2(n8787), .A(n8786), .B(n8785), .ZN(n13798)
         );
  OAI21_X1 U11273 ( .B1(n13897), .B2(n8789), .A(n13798), .ZN(n8790) );
  INV_X1 U11274 ( .A(n8790), .ZN(n8801) );
  NAND2_X1 U11275 ( .A1(n8792), .A2(n8791), .ZN(n8795) );
  INV_X1 U11276 ( .A(SI_29_), .ZN(n12954) );
  NAND2_X1 U11277 ( .A1(n8793), .A2(n12954), .ZN(n8794) );
  MUX2_X1 U11278 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6439), .Z(n8810) );
  XNOR2_X1 U11279 ( .A(n8810), .B(SI_30_), .ZN(n8813) );
  INV_X1 U11280 ( .A(n8813), .ZN(n8796) );
  NAND2_X1 U11281 ( .A1(n12152), .A2(n8745), .ZN(n8799) );
  NAND2_X1 U11282 ( .A1(n8797), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8798) );
  MUX2_X1 U11283 ( .A(n8801), .B(n13900), .S(n8800), .Z(n8808) );
  NAND2_X1 U11284 ( .A1(n8800), .A2(n13897), .ZN(n8804) );
  INV_X1 U11285 ( .A(n13798), .ZN(n8802) );
  AOI21_X1 U11286 ( .B1(n8804), .B2(n8803), .A(n8802), .ZN(n8805) );
  AOI21_X1 U11287 ( .B1(n13900), .B2(n8806), .A(n8805), .ZN(n8807) );
  NAND2_X1 U11288 ( .A1(n8808), .A2(n8807), .ZN(n8809) );
  INV_X1 U11289 ( .A(n8810), .ZN(n8811) );
  INV_X1 U11290 ( .A(SI_30_), .ZN(n12948) );
  MUX2_X1 U11291 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9831), .Z(n8815) );
  XNOR2_X1 U11292 ( .A(n8815), .B(SI_31_), .ZN(n8816) );
  NAND2_X1 U11293 ( .A1(n13622), .A2(n8745), .ZN(n8819) );
  NAND2_X1 U11294 ( .A1(n8797), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8818) );
  XOR2_X1 U11295 ( .A(n13897), .B(n8850), .Z(n8845) );
  NAND2_X1 U11296 ( .A1(n10281), .A2(n14345), .ZN(n10687) );
  NAND2_X1 U11297 ( .A1(n8820), .A2(n10242), .ZN(n10277) );
  INV_X1 U11298 ( .A(n8820), .ZN(n10244) );
  NAND2_X1 U11299 ( .A1(n10244), .A2(n11378), .ZN(n10247) );
  NAND2_X1 U11300 ( .A1(n10277), .A2(n10247), .ZN(n8821) );
  NAND2_X1 U11301 ( .A1(n10687), .A2(n8821), .ZN(n8851) );
  NOR3_X1 U11302 ( .A1(n8860), .A2(n8845), .A3(n8851), .ZN(n8867) );
  XOR2_X1 U11303 ( .A(n13798), .B(n13900), .Z(n8844) );
  XNOR2_X1 U11304 ( .A(n12382), .B(n13799), .ZN(n12380) );
  NAND2_X1 U11305 ( .A1(n13921), .A2(n13701), .ZN(n12379) );
  OR2_X1 U11306 ( .A1(n13921), .A2(n13701), .ZN(n8822) );
  NAND2_X1 U11307 ( .A1(n12379), .A2(n8822), .ZN(n13920) );
  XNOR2_X1 U11308 ( .A(n13940), .B(n13779), .ZN(n12377) );
  XNOR2_X1 U11309 ( .A(n13964), .B(n13943), .ZN(n13956) );
  XNOR2_X1 U11310 ( .A(n14012), .B(n13802), .ZN(n14008) );
  XNOR2_X1 U11311 ( .A(n14144), .B(n13681), .ZN(n12364) );
  OR2_X1 U11312 ( .A1(n14150), .A2(n8824), .ZN(n12362) );
  NAND2_X1 U11313 ( .A1(n14150), .A2(n8824), .ZN(n8825) );
  NAND2_X1 U11314 ( .A1(n12362), .A2(n8825), .ZN(n11810) );
  NAND2_X1 U11315 ( .A1(n11721), .A2(n8826), .ZN(n11727) );
  XNOR2_X1 U11316 ( .A(n11616), .B(n11843), .ZN(n11482) );
  XNOR2_X1 U11317 ( .A(n14343), .B(n12206), .ZN(n14347) );
  XNOR2_X1 U11318 ( .A(n11835), .B(n11833), .ZN(n11477) );
  XNOR2_X1 U11319 ( .A(n14491), .B(n11828), .ZN(n11153) );
  XNOR2_X1 U11320 ( .A(n14739), .B(n11553), .ZN(n11250) );
  XNOR2_X1 U11321 ( .A(n14717), .B(n13806), .ZN(n11144) );
  NAND2_X1 U11322 ( .A1(n8827), .A2(n10694), .ZN(n10749) );
  NAND2_X1 U11323 ( .A1(n8828), .A2(n7038), .ZN(n8829) );
  NAND4_X1 U11324 ( .A1(n10737), .A2(n10686), .A3(n10251), .A4(n10820), .ZN(
        n8830) );
  XNOR2_X1 U11325 ( .A(n11019), .B(n11017), .ZN(n10863) );
  XNOR2_X1 U11326 ( .A(n13810), .B(n10951), .ZN(n10954) );
  NOR3_X1 U11327 ( .A1(n8830), .A2(n10863), .A3(n10954), .ZN(n8831) );
  XNOR2_X1 U11328 ( .A(n11193), .B(n13807), .ZN(n10977) );
  XNOR2_X1 U11329 ( .A(n14612), .B(n13808), .ZN(n10967) );
  NAND4_X1 U11330 ( .A1(n11144), .A2(n8831), .A3(n10977), .A4(n10967), .ZN(
        n8832) );
  OR4_X1 U11331 ( .A1(n11477), .A2(n11153), .A3(n11250), .A4(n8832), .ZN(n8833) );
  OR4_X1 U11332 ( .A1(n11727), .A2(n11482), .A3(n14347), .A4(n8833), .ZN(n8834) );
  XNOR2_X1 U11333 ( .A(n12232), .B(n13792), .ZN(n11730) );
  OR4_X1 U11334 ( .A1(n11810), .A2(n8834), .A3(n11591), .A4(n11730), .ZN(n8835) );
  NOR2_X1 U11335 ( .A1(n12364), .A2(n8835), .ZN(n8836) );
  XNOR2_X1 U11336 ( .A(n14130), .B(n14039), .ZN(n12367) );
  NAND4_X1 U11337 ( .A1(n14008), .A2(n14036), .A3(n8836), .A4(n12367), .ZN(
        n8837) );
  NOR2_X1 U11338 ( .A1(n13989), .A2(n8837), .ZN(n8839) );
  NAND3_X1 U11339 ( .A1(n13956), .A2(n8839), .A3(n13976), .ZN(n8840) );
  NOR3_X1 U11340 ( .A1(n13920), .A2(n12377), .A3(n8840), .ZN(n8842) );
  NAND2_X1 U11341 ( .A1(n14082), .A2(n13800), .ZN(n12360) );
  OR2_X1 U11342 ( .A1(n14082), .A2(n13800), .ZN(n8841) );
  NAND2_X1 U11343 ( .A1(n12360), .A2(n8841), .ZN(n13916) );
  NAND4_X1 U11344 ( .A1(n12380), .A2(n8842), .A3(n12400), .A4(n13916), .ZN(
        n8843) );
  NOR3_X1 U11345 ( .A1(n8845), .A2(n8844), .A3(n8843), .ZN(n8846) );
  NAND2_X1 U11346 ( .A1(n11492), .A2(n8847), .ZN(n10675) );
  NAND2_X1 U11347 ( .A1(n8851), .A2(n10675), .ZN(n8857) );
  NOR3_X1 U11348 ( .A1(n14069), .A2(n13897), .A3(n8857), .ZN(n8849) );
  NAND2_X1 U11349 ( .A1(n8850), .A2(n8800), .ZN(n8855) );
  NOR3_X1 U11350 ( .A1(n8855), .A2(n13897), .A3(n8851), .ZN(n8848) );
  AOI21_X1 U11351 ( .B1(n8849), .B2(n8855), .A(n8848), .ZN(n8854) );
  NOR2_X1 U11352 ( .A1(n8850), .A2(n8800), .ZN(n8858) );
  XOR2_X1 U11353 ( .A(n8851), .B(n8858), .Z(n8852) );
  NAND3_X1 U11354 ( .A1(n8852), .A2(n14069), .A3(n13897), .ZN(n8853) );
  NOR2_X1 U11355 ( .A1(n8855), .A2(n13897), .ZN(n8856) );
  AOI211_X1 U11356 ( .C1(n8858), .C2(n13897), .A(n8857), .B(n8856), .ZN(n8859)
         );
  NAND2_X1 U11357 ( .A1(n8868), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8863) );
  INV_X1 U11358 ( .A(n10933), .ZN(n8864) );
  NAND2_X1 U11359 ( .A1(n8864), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11746) );
  INV_X1 U11360 ( .A(n11746), .ZN(n8865) );
  OAI21_X1 U11361 ( .B1(n8867), .B2(n8866), .A(n8865), .ZN(n8887) );
  INV_X1 U11362 ( .A(n8872), .ZN(n8873) );
  NAND2_X1 U11363 ( .A1(n8873), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8874) );
  NAND2_X1 U11364 ( .A1(n8877), .A2(n8874), .ZN(n8876) );
  INV_X1 U11365 ( .A(n8877), .ZN(n8878) );
  NAND2_X1 U11366 ( .A1(n8878), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n8880) );
  NAND2_X1 U11367 ( .A1(n10224), .A2(n10222), .ZN(n8881) );
  INV_X1 U11368 ( .A(n10277), .ZN(n9812) );
  INV_X1 U11369 ( .A(n8882), .ZN(n10252) );
  NAND2_X1 U11370 ( .A1(n8883), .A2(n11378), .ZN(n10275) );
  NAND2_X1 U11371 ( .A1(n10275), .A2(n9812), .ZN(n10932) );
  NAND3_X1 U11372 ( .A1(n10272), .A2(n14339), .A3(n10932), .ZN(n14575) );
  NOR2_X1 U11373 ( .A1(n14575), .A2(n14197), .ZN(n8885) );
  OAI21_X1 U11374 ( .B1(n11746), .B2(n8820), .A(P1_B_REG_SCAN_IN), .ZN(n8884)
         );
  OR2_X1 U11375 ( .A1(n8885), .A2(n8884), .ZN(n8886) );
  NAND2_X1 U11376 ( .A1(n8887), .A2(n8886), .ZN(P1_U3242) );
  NOR2_X1 U11377 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n9081) );
  NAND2_X1 U11378 ( .A1(n9081), .A2(n9080), .ZN(n9098) );
  INV_X1 U11379 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n9266) );
  INV_X1 U11380 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8888) );
  INV_X1 U11381 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8890) );
  NAND2_X1 U11382 ( .A1(n8961), .A2(n8890), .ZN(n8963) );
  NAND2_X1 U11383 ( .A1(n8963), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8891) );
  NAND2_X1 U11384 ( .A1(n9343), .A2(n8891), .ZN(n12691) );
  NAND2_X1 U11385 ( .A1(n8955), .A2(n8954), .ZN(n8900) );
  NAND2_X1 U11386 ( .A1(n8956), .A2(n8957), .ZN(n8906) );
  NAND2_X1 U11387 ( .A1(n12691), .A2(n9286), .ZN(n8915) );
  INV_X1 U11388 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12693) );
  INV_X1 U11389 ( .A(n9115), .ZN(n9361) );
  AND2_X2 U11390 ( .A1(n12950), .A2(n8910), .ZN(n9052) );
  NAND2_X1 U11391 ( .A1(n9083), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8912) );
  NAND2_X1 U11392 ( .A1(n9231), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8911) );
  OAI211_X1 U11393 ( .C1(n12693), .C2(n9361), .A(n8912), .B(n8911), .ZN(n8913)
         );
  INV_X1 U11394 ( .A(n8913), .ZN(n8914) );
  INV_X1 U11395 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8916) );
  AOI22_X1 U11396 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n8916), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n8950), .ZN(n9315) );
  INV_X1 U11397 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U11398 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n11709), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n8948), .ZN(n9302) );
  AOI22_X1 U11399 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n7250), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n11376), .ZN(n9292) );
  AOI22_X1 U11400 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n8023), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n12155), .ZN(n9275) );
  AOI22_X1 U11401 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n6640), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n7649), .ZN(n9258) );
  NAND2_X1 U11402 ( .A1(n9030), .A2(n9045), .ZN(n8919) );
  NAND2_X1 U11403 ( .A1(n9830), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8918) );
  NAND2_X1 U11404 ( .A1(n9848), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8920) );
  NAND2_X1 U11405 ( .A1(n9866), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8921) );
  AND2_X1 U11406 ( .A1(n9868), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8922) );
  INV_X1 U11407 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9856) );
  NAND2_X1 U11408 ( .A1(n9856), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8923) );
  INV_X1 U11409 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9858) );
  NAND2_X1 U11410 ( .A1(n9858), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8924) );
  NAND2_X1 U11411 ( .A1(n8925), .A2(n8924), .ZN(n9089) );
  NAND2_X1 U11412 ( .A1(n9862), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8926) );
  NAND2_X1 U11413 ( .A1(n9876), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8929) );
  NAND2_X1 U11414 ( .A1(n9874), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8928) );
  NAND2_X1 U11415 ( .A1(n8929), .A2(n8928), .ZN(n9104) );
  XNOR2_X1 U11416 ( .A(n7240), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n9120) );
  NAND2_X1 U11417 ( .A1(n9925), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8931) );
  XNOR2_X1 U11418 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n9193) );
  NAND2_X1 U11419 ( .A1(n9967), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8934) );
  NAND2_X1 U11420 ( .A1(n9208), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n8938) );
  NAND2_X1 U11421 ( .A1(n8936), .A2(n8935), .ZN(n8937) );
  XNOR2_X1 U11422 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n9223) );
  NAND2_X1 U11423 ( .A1(n8939), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8940) );
  XNOR2_X1 U11424 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n9239) );
  XNOR2_X1 U11425 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n9002) );
  NAND2_X1 U11426 ( .A1(n8941), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8942) );
  NOR2_X1 U11427 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n10587), .ZN(n8944) );
  NAND2_X1 U11428 ( .A1(n10587), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8945) );
  NAND2_X1 U11429 ( .A1(n9275), .A2(n9276), .ZN(n8946) );
  INV_X1 U11430 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11856) );
  AOI22_X1 U11431 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(
        P1_DATAO_REG_21__SCAN_IN), .B1(n11856), .B2(n15178), .ZN(n8975) );
  NAND2_X1 U11432 ( .A1(n9315), .A2(n9316), .ZN(n8949) );
  INV_X1 U11433 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8952) );
  INV_X1 U11434 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n14202) );
  INV_X1 U11435 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13648) );
  AOI22_X1 U11436 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n13648), .B2(n11859), .ZN(n8970) );
  AOI22_X1 U11437 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(
        P1_DATAO_REG_26__SCAN_IN), .B1(n13643), .B2(n14200), .ZN(n9336) );
  INV_X1 U11438 ( .A(n9336), .ZN(n8953) );
  XNOR2_X1 U11439 ( .A(n9337), .B(n8953), .ZN(n12958) );
  NAND2_X1 U11440 ( .A1(n12958), .A2(n6437), .ZN(n8960) );
  OR2_X1 U11441 ( .A1(n6440), .A2(n12961), .ZN(n8959) );
  INV_X1 U11442 ( .A(n8961), .ZN(n9330) );
  NAND2_X1 U11443 ( .A1(n9330), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8962) );
  NAND2_X1 U11444 ( .A1(n8963), .A2(n8962), .ZN(n12711) );
  NAND2_X1 U11445 ( .A1(n12711), .A2(n9286), .ZN(n8969) );
  NAND2_X1 U11446 ( .A1(n9473), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8967) );
  NAND2_X1 U11447 ( .A1(n9083), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8966) );
  AND3_X1 U11448 ( .A1(n8967), .A2(n8966), .A3(n8965), .ZN(n8968) );
  INV_X1 U11449 ( .A(n8970), .ZN(n8971) );
  XNOR2_X1 U11450 ( .A(n8972), .B(n8971), .ZN(n11522) );
  NAND2_X1 U11451 ( .A1(n11522), .A2(n9059), .ZN(n8974) );
  OR2_X1 U11452 ( .A1(n6440), .A2(n11523), .ZN(n8973) );
  INV_X1 U11453 ( .A(n12847), .ZN(n12713) );
  INV_X1 U11454 ( .A(n8975), .ZN(n8976) );
  XNOR2_X1 U11455 ( .A(n8977), .B(n8976), .ZN(n10713) );
  NAND2_X1 U11456 ( .A1(n10713), .A2(n9059), .ZN(n8979) );
  INV_X1 U11457 ( .A(SI_21_), .ZN(n10715) );
  NAND2_X1 U11458 ( .A1(n9298), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8980) );
  NAND2_X1 U11459 ( .A1(n9306), .A2(n8980), .ZN(n12763) );
  NAND2_X1 U11460 ( .A1(n12763), .A2(n9286), .ZN(n8983) );
  AOI22_X1 U11461 ( .A1(n9473), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n9231), .B2(
        P3_REG0_REG_21__SCAN_IN), .ZN(n8982) );
  INV_X2 U11462 ( .A(n8964), .ZN(n9083) );
  NAND2_X1 U11463 ( .A1(n9083), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8981) );
  INV_X1 U11464 ( .A(n12769), .ZN(n12543) );
  AOI22_X1 U11465 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n10587), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n7642), .ZN(n8984) );
  INV_X1 U11466 ( .A(n8984), .ZN(n8985) );
  XNOR2_X1 U11467 ( .A(n8986), .B(n8985), .ZN(n10194) );
  NAND2_X1 U11468 ( .A1(n10194), .A2(n6437), .ZN(n8995) );
  NOR2_X1 U11469 ( .A1(n8989), .A2(n9225), .ZN(n8990) );
  MUX2_X1 U11470 ( .A(n9225), .B(n8990), .S(P3_IR_REG_17__SCAN_IN), .Z(n8991)
         );
  INV_X1 U11471 ( .A(n8991), .ZN(n8992) );
  AND2_X1 U11472 ( .A1(n9277), .A2(n8992), .ZN(n12651) );
  OAI22_X1 U11473 ( .A1(n6440), .A2(n6898), .B1(n9280), .B2(n14413), .ZN(n8993) );
  INV_X1 U11474 ( .A(n8993), .ZN(n8994) );
  INV_X1 U11475 ( .A(n9267), .ZN(n8997) );
  NAND2_X1 U11476 ( .A1(n9011), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8996) );
  NAND2_X1 U11477 ( .A1(n8997), .A2(n8996), .ZN(n12819) );
  NAND2_X1 U11478 ( .A1(n12819), .A2(n9286), .ZN(n9001) );
  NAND2_X1 U11479 ( .A1(n9083), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9000) );
  NAND2_X1 U11480 ( .A1(n9231), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8999) );
  NAND2_X1 U11481 ( .A1(n9473), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8998) );
  OR2_X1 U11482 ( .A1(n12929), .A2(n12829), .ZN(n9590) );
  NAND2_X1 U11483 ( .A1(n12929), .A2(n12829), .ZN(n9595) );
  NAND2_X1 U11484 ( .A1(n9590), .A2(n9595), .ZN(n12810) );
  INV_X1 U11485 ( .A(n9002), .ZN(n9003) );
  XNOR2_X1 U11486 ( .A(n9004), .B(n9003), .ZN(n10137) );
  NAND2_X1 U11487 ( .A1(n10137), .A2(n9059), .ZN(n9009) );
  NAND2_X1 U11488 ( .A1(n9005), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9006) );
  XNOR2_X1 U11489 ( .A(n9006), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12650) );
  OAI22_X1 U11490 ( .A1(n6440), .A2(n10139), .B1(n9280), .B2(n14393), .ZN(
        n9007) );
  INV_X1 U11491 ( .A(n9007), .ZN(n9008) );
  NAND2_X1 U11492 ( .A1(n9009), .A2(n9008), .ZN(n12832) );
  NAND2_X1 U11493 ( .A1(n9083), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n9015) );
  NAND2_X1 U11494 ( .A1(n9231), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n9014) );
  NAND2_X1 U11495 ( .A1(n9249), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9010) );
  NAND2_X1 U11496 ( .A1(n9011), .A2(n9010), .ZN(n12833) );
  NAND2_X1 U11497 ( .A1(n9286), .A2(n12833), .ZN(n9013) );
  NAND2_X1 U11498 ( .A1(n9473), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n9012) );
  INV_X1 U11499 ( .A(n12812), .ZN(n12546) );
  OR2_X1 U11500 ( .A1(n12832), .A2(n12546), .ZN(n12808) );
  AND2_X1 U11501 ( .A1(n12810), .A2(n12808), .ZN(n9256) );
  NAND2_X1 U11502 ( .A1(n9051), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n9019) );
  NAND2_X1 U11503 ( .A1(n9052), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n9018) );
  NAND2_X1 U11504 ( .A1(n9115), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n9017) );
  NAND2_X1 U11505 ( .A1(n9038), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n9016) );
  XNOR2_X1 U11506 ( .A(n9866), .B(P2_DATAO_REG_2__SCAN_IN), .ZN(n9020) );
  XNOR2_X1 U11507 ( .A(n9021), .B(n9020), .ZN(n9844) );
  NAND2_X1 U11508 ( .A1(n9059), .A2(n9844), .ZN(n9025) );
  OR2_X1 U11509 ( .A1(n9339), .A2(SI_2_), .ZN(n9024) );
  OR2_X1 U11510 ( .A1(n9048), .A2(n12569), .ZN(n9023) );
  NAND2_X1 U11511 ( .A1(n10516), .A2(n15077), .ZN(n9530) );
  NAND2_X1 U11512 ( .A1(n9115), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n9029) );
  NAND2_X1 U11513 ( .A1(n9052), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U11514 ( .A1(n9051), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n9027) );
  NAND2_X1 U11515 ( .A1(n9038), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n9026) );
  XNOR2_X1 U11516 ( .A(n9030), .B(n9045), .ZN(n9835) );
  INV_X1 U11517 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n9033) );
  INV_X1 U11518 ( .A(n10422), .ZN(n9034) );
  NAND2_X1 U11519 ( .A1(n10904), .A2(n12558), .ZN(n9521) );
  NAND2_X1 U11520 ( .A1(n9525), .A2(n9521), .ZN(n9502) );
  NAND2_X1 U11521 ( .A1(n9038), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9042) );
  NAND2_X1 U11522 ( .A1(n9051), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9041) );
  NAND2_X1 U11523 ( .A1(n9115), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9040) );
  NAND2_X1 U11524 ( .A1(n9052), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n9039) );
  AND2_X1 U11525 ( .A1(n9043), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9044) );
  NOR2_X1 U11526 ( .A1(n9045), .A2(n9044), .ZN(n9047) );
  OAI21_X1 U11527 ( .B1(n9831), .B2(n9047), .A(n9046), .ZN(n12963) );
  NAND2_X1 U11528 ( .A1(n9502), .A2(n10906), .ZN(n9050) );
  NAND2_X1 U11529 ( .A1(n15085), .A2(n10904), .ZN(n9049) );
  NAND2_X1 U11530 ( .A1(n9050), .A2(n9049), .ZN(n15083) );
  INV_X1 U11531 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10522) );
  NAND2_X1 U11532 ( .A1(n9286), .A2(n10522), .ZN(n9056) );
  NAND2_X1 U11533 ( .A1(n9115), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9055) );
  NAND2_X1 U11534 ( .A1(n9052), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n9054) );
  XNOR2_X1 U11535 ( .A(n9868), .B(P2_DATAO_REG_3__SCAN_IN), .ZN(n9057) );
  XNOR2_X1 U11536 ( .A(n9058), .B(n9057), .ZN(n9842) );
  NAND2_X1 U11537 ( .A1(n9059), .A2(n9842), .ZN(n9065) );
  OR2_X1 U11538 ( .A1(n9339), .A2(SI_3_), .ZN(n9064) );
  XNOR2_X1 U11539 ( .A(n9062), .B(P3_IR_REG_3__SCAN_IN), .ZN(n14889) );
  OR2_X1 U11540 ( .A1(n9280), .A2(n14889), .ZN(n9063) );
  INV_X1 U11541 ( .A(n15086), .ZN(n12556) );
  NAND2_X1 U11542 ( .A1(n12556), .A2(n10732), .ZN(n9066) );
  NAND2_X1 U11543 ( .A1(n10725), .A2(n9066), .ZN(n15065) );
  NAND2_X1 U11544 ( .A1(n9231), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n9070) );
  NAND2_X1 U11545 ( .A1(n9083), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n9069) );
  OR2_X1 U11546 ( .A1(n7569), .A2(n9081), .ZN(n15070) );
  NAND2_X1 U11547 ( .A1(n9286), .A2(n15070), .ZN(n9068) );
  NAND2_X1 U11548 ( .A1(n9115), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9067) );
  XNOR2_X1 U11549 ( .A(n9072), .B(n9071), .ZN(n9849) );
  NAND2_X1 U11550 ( .A1(n9059), .A2(n9849), .ZN(n9077) );
  OR2_X1 U11551 ( .A1(n9339), .A2(SI_4_), .ZN(n9076) );
  NAND2_X1 U11552 ( .A1(n9090), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9074) );
  OR2_X1 U11553 ( .A1(n9280), .A2(n14907), .ZN(n9075) );
  NAND2_X1 U11554 ( .A1(n10893), .A2(n15069), .ZN(n9539) );
  INV_X1 U11555 ( .A(n15069), .ZN(n9078) );
  NAND2_X1 U11556 ( .A1(n12555), .A2(n9078), .ZN(n9542) );
  NAND2_X1 U11557 ( .A1(n9539), .A2(n9542), .ZN(n15064) );
  NAND2_X1 U11558 ( .A1(n15065), .A2(n15064), .ZN(n15063) );
  NAND2_X1 U11559 ( .A1(n12555), .A2(n15069), .ZN(n9079) );
  NAND2_X1 U11560 ( .A1(n9231), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n9087) );
  NAND2_X1 U11561 ( .A1(n9473), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n9086) );
  OR2_X1 U11562 ( .A1(n9081), .A2(n9080), .ZN(n9082) );
  NAND2_X1 U11563 ( .A1(n9098), .A2(n9082), .ZN(n10899) );
  NAND2_X1 U11564 ( .A1(n9286), .A2(n10899), .ZN(n9085) );
  NAND2_X1 U11565 ( .A1(n9083), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n9084) );
  XNOR2_X1 U11566 ( .A(n9089), .B(n9088), .ZN(n9851) );
  NAND2_X1 U11567 ( .A1(n6437), .A2(n9851), .ZN(n9095) );
  OR2_X1 U11568 ( .A1(n6440), .A2(SI_5_), .ZN(n9094) );
  NAND2_X1 U11569 ( .A1(n9106), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9092) );
  XNOR2_X1 U11570 ( .A(n9092), .B(n9091), .ZN(n14922) );
  OR2_X1 U11571 ( .A1(n9280), .A2(n6854), .ZN(n9093) );
  NAND2_X1 U11572 ( .A1(n15061), .A2(n10811), .ZN(n9544) );
  INV_X1 U11573 ( .A(n15061), .ZN(n12554) );
  INV_X1 U11574 ( .A(n10811), .ZN(n10898) );
  NAND2_X1 U11575 ( .A1(n12554), .A2(n10898), .ZN(n9540) );
  NAND2_X1 U11576 ( .A1(n15061), .A2(n10898), .ZN(n9097) );
  NAND2_X1 U11577 ( .A1(n9098), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9099) );
  NAND2_X1 U11578 ( .A1(n9113), .A2(n9099), .ZN(n15055) );
  NAND2_X1 U11579 ( .A1(n9286), .A2(n15055), .ZN(n9103) );
  NAND2_X1 U11580 ( .A1(n9083), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n9102) );
  NAND2_X1 U11581 ( .A1(n9473), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9101) );
  NAND2_X1 U11582 ( .A1(n9231), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n9100) );
  INV_X1 U11583 ( .A(SI_6_), .ZN(n9839) );
  XNOR2_X1 U11584 ( .A(n9105), .B(n9104), .ZN(n9838) );
  NAND2_X1 U11585 ( .A1(n9059), .A2(n9838), .ZN(n9109) );
  OR2_X1 U11586 ( .A1(n9123), .A2(n9225), .ZN(n9107) );
  XNOR2_X1 U11587 ( .A(n9107), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10541) );
  OR2_X1 U11588 ( .A1(n9280), .A2(n10548), .ZN(n9108) );
  OAI211_X1 U11589 ( .C1(n6440), .C2(n9839), .A(n9109), .B(n9108), .ZN(n9111)
         );
  NAND2_X1 U11590 ( .A1(n11102), .A2(n9111), .ZN(n9549) );
  INV_X1 U11591 ( .A(n9111), .ZN(n15056) );
  NAND2_X1 U11592 ( .A1(n12553), .A2(n15056), .ZN(n9545) );
  NAND2_X1 U11593 ( .A1(n12553), .A2(n9111), .ZN(n9112) );
  NAND2_X1 U11594 ( .A1(n9231), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n9119) );
  NAND2_X1 U11595 ( .A1(n9052), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n9118) );
  AND2_X1 U11596 ( .A1(n9113), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9114) );
  OR2_X1 U11597 ( .A1(n9114), .A2(n9130), .ZN(n11104) );
  NAND2_X1 U11598 ( .A1(n9286), .A2(n11104), .ZN(n9117) );
  NAND2_X1 U11599 ( .A1(n9473), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n9116) );
  XNOR2_X1 U11600 ( .A(n9121), .B(n9120), .ZN(n9846) );
  NAND2_X1 U11601 ( .A1(n6437), .A2(n9846), .ZN(n9127) );
  OR2_X1 U11602 ( .A1(n6440), .A2(SI_7_), .ZN(n9126) );
  INV_X1 U11603 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9122) );
  OR2_X1 U11604 ( .A1(n9139), .A2(n9225), .ZN(n9124) );
  XNOR2_X1 U11605 ( .A(n9124), .B(n9138), .ZN(n10571) );
  INV_X1 U11606 ( .A(n10571), .ZN(n10533) );
  OR2_X1 U11607 ( .A1(n9280), .A2(n10533), .ZN(n9125) );
  NAND2_X1 U11608 ( .A1(n15046), .A2(n11100), .ZN(n9550) );
  INV_X1 U11609 ( .A(n11100), .ZN(n10883) );
  NAND2_X1 U11610 ( .A1(n12552), .A2(n10883), .ZN(n9551) );
  NAND2_X1 U11611 ( .A1(n9550), .A2(n9551), .ZN(n11055) );
  NAND2_X1 U11612 ( .A1(n10878), .A2(n11055), .ZN(n10877) );
  NAND2_X1 U11613 ( .A1(n12552), .A2(n11100), .ZN(n9128) );
  NAND2_X1 U11614 ( .A1(n9083), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n9135) );
  NOR2_X1 U11615 ( .A1(n9130), .A2(n10556), .ZN(n9131) );
  OR2_X1 U11616 ( .A1(n9151), .A2(n9131), .ZN(n11219) );
  NAND2_X1 U11617 ( .A1(n9286), .A2(n11219), .ZN(n9133) );
  NAND2_X1 U11618 ( .A1(n9115), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9132) );
  NAND4_X1 U11619 ( .A1(n9135), .A2(n9134), .A3(n9133), .A4(n9132), .ZN(n12551) );
  INV_X1 U11620 ( .A(SI_8_), .ZN(n9854) );
  XNOR2_X1 U11621 ( .A(n9881), .B(P2_DATAO_REG_8__SCAN_IN), .ZN(n9136) );
  XNOR2_X1 U11622 ( .A(n9137), .B(n9136), .ZN(n9852) );
  NAND2_X1 U11623 ( .A1(n9059), .A2(n9852), .ZN(n9146) );
  NOR2_X1 U11624 ( .A1(n9143), .A2(n9225), .ZN(n9140) );
  MUX2_X1 U11625 ( .A(n9225), .B(n9140), .S(P3_IR_REG_8__SCAN_IN), .Z(n9141)
         );
  INV_X1 U11626 ( .A(n9141), .ZN(n9144) );
  NAND2_X1 U11627 ( .A1(n9143), .A2(n9142), .ZN(n9171) );
  NAND2_X1 U11628 ( .A1(n9144), .A2(n9171), .ZN(n12635) );
  OR2_X1 U11629 ( .A1(n9280), .A2(n12635), .ZN(n9145) );
  OAI211_X1 U11630 ( .C1(n6440), .C2(n9854), .A(n9146), .B(n9145), .ZN(n9553)
         );
  XNOR2_X1 U11631 ( .A(n12551), .B(n9553), .ZN(n11046) );
  INV_X1 U11632 ( .A(n12551), .ZN(n11097) );
  INV_X1 U11633 ( .A(n9553), .ZN(n11214) );
  NAND2_X1 U11634 ( .A1(n11097), .A2(n11214), .ZN(n9149) );
  NAND2_X1 U11635 ( .A1(n9231), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n9156) );
  NAND2_X1 U11636 ( .A1(n9083), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n9155) );
  OR2_X1 U11637 ( .A1(n9151), .A2(n9150), .ZN(n9152) );
  NAND2_X1 U11638 ( .A1(n9163), .A2(n9152), .ZN(n11178) );
  NAND2_X1 U11639 ( .A1(n9286), .A2(n11178), .ZN(n9154) );
  NAND2_X1 U11640 ( .A1(n9473), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n9153) );
  NAND4_X1 U11641 ( .A1(n9156), .A2(n9155), .A3(n9154), .A4(n9153), .ZN(n12550) );
  XNOR2_X1 U11642 ( .A(n15276), .B(P2_DATAO_REG_9__SCAN_IN), .ZN(n9157) );
  XNOR2_X1 U11643 ( .A(n9158), .B(n9157), .ZN(n9860) );
  NAND2_X1 U11644 ( .A1(n6437), .A2(n9860), .ZN(n9162) );
  NAND2_X1 U11645 ( .A1(n9171), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9160) );
  INV_X1 U11646 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9159) );
  XNOR2_X1 U11647 ( .A(n9160), .B(n9159), .ZN(n14940) );
  INV_X1 U11648 ( .A(n14940), .ZN(n12603) );
  OR2_X1 U11649 ( .A1(n9280), .A2(n12603), .ZN(n9161) );
  OAI211_X1 U11650 ( .C1(n6440), .C2(SI_9_), .A(n9162), .B(n9161), .ZN(n15135)
         );
  XNOR2_X1 U11651 ( .A(n12550), .B(n15135), .ZN(n11174) );
  INV_X1 U11652 ( .A(n15135), .ZN(n11181) );
  NAND2_X1 U11653 ( .A1(n9083), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9168) );
  NAND2_X1 U11654 ( .A1(n9231), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n9167) );
  NAND2_X1 U11655 ( .A1(n9163), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9164) );
  NAND2_X1 U11656 ( .A1(n9178), .A2(n9164), .ZN(n11374) );
  NAND2_X1 U11657 ( .A1(n9286), .A2(n11374), .ZN(n9166) );
  NAND2_X1 U11658 ( .A1(n9473), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n9165) );
  NAND4_X1 U11659 ( .A1(n9168), .A2(n9167), .A3(n9166), .A4(n9165), .ZN(n12549) );
  XNOR2_X1 U11660 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n9169) );
  XNOR2_X1 U11661 ( .A(n9170), .B(n9169), .ZN(n9863) );
  NAND2_X1 U11662 ( .A1(n9863), .A2(n9059), .ZN(n9176) );
  NAND2_X1 U11663 ( .A1(n9186), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9173) );
  INV_X1 U11664 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9172) );
  OAI22_X1 U11665 ( .A1(n6440), .A2(SI_10_), .B1(n12641), .B2(n9280), .ZN(
        n9174) );
  INV_X1 U11666 ( .A(n9174), .ZN(n9175) );
  NAND2_X1 U11667 ( .A1(n9176), .A2(n9175), .ZN(n11356) );
  XNOR2_X1 U11668 ( .A(n12549), .B(n11356), .ZN(n11226) );
  INV_X1 U11669 ( .A(n11356), .ZN(n11362) );
  NAND2_X1 U11670 ( .A1(n12549), .A2(n11362), .ZN(n9177) );
  NAND2_X1 U11671 ( .A1(n9083), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n9183) );
  NAND2_X1 U11672 ( .A1(n9038), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n9182) );
  NAND2_X1 U11673 ( .A1(n9178), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9179) );
  NAND2_X1 U11674 ( .A1(n9202), .A2(n9179), .ZN(n11438) );
  NAND2_X1 U11675 ( .A1(n9286), .A2(n11438), .ZN(n9181) );
  NAND2_X1 U11676 ( .A1(n9473), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n9180) );
  XNOR2_X1 U11677 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9184) );
  XNOR2_X1 U11678 ( .A(n9185), .B(n9184), .ZN(n14317) );
  NAND2_X1 U11679 ( .A1(n14317), .A2(n9059), .ZN(n9190) );
  XNOR2_X1 U11680 ( .A(n9187), .B(P3_IR_REG_11__SCAN_IN), .ZN(n12643) );
  NAND2_X1 U11681 ( .A1(n11394), .A2(n11571), .ZN(n9191) );
  NAND2_X1 U11682 ( .A1(n11348), .A2(n14436), .ZN(n9192) );
  INV_X1 U11683 ( .A(n9193), .ZN(n9194) );
  XNOR2_X1 U11684 ( .A(n9195), .B(n9194), .ZN(n14321) );
  NAND2_X1 U11685 ( .A1(n14321), .A2(n6437), .ZN(n9201) );
  NAND2_X1 U11686 ( .A1(n9196), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9197) );
  XNOR2_X1 U11687 ( .A(n9197), .B(P3_IR_REG_12__SCAN_IN), .ZN(n14991) );
  INV_X1 U11688 ( .A(n14991), .ZN(n14323) );
  OAI22_X1 U11689 ( .A1(n6440), .A2(n9198), .B1(n9280), .B2(n14323), .ZN(n9199) );
  INV_X1 U11690 ( .A(n9199), .ZN(n9200) );
  NAND2_X1 U11691 ( .A1(n9201), .A2(n9200), .ZN(n14443) );
  NAND2_X1 U11692 ( .A1(n9231), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n9207) );
  AND2_X1 U11693 ( .A1(n9202), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9203) );
  OR2_X1 U11694 ( .A1(n9203), .A2(n9216), .ZN(n14440) );
  NAND2_X1 U11695 ( .A1(n9286), .A2(n14440), .ZN(n9206) );
  NAND2_X1 U11696 ( .A1(n9473), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U11697 ( .A1(n9083), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n9204) );
  OR2_X1 U11698 ( .A1(n14443), .A2(n11675), .ZN(n9570) );
  NAND2_X1 U11699 ( .A1(n14443), .A2(n11675), .ZN(n9572) );
  NAND2_X1 U11700 ( .A1(n9570), .A2(n9572), .ZN(n9402) );
  INV_X1 U11701 ( .A(n11675), .ZN(n12548) );
  XNOR2_X1 U11702 ( .A(n9208), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n9956) );
  NAND2_X1 U11703 ( .A1(n9956), .A2(n6437), .ZN(n9214) );
  NAND2_X1 U11704 ( .A1(n9209), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9211) );
  INV_X1 U11705 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n9210) );
  XNOR2_X1 U11706 ( .A(n9211), .B(n9210), .ZN(n15012) );
  INV_X1 U11707 ( .A(n15012), .ZN(n12613) );
  OAI22_X1 U11708 ( .A1(n6440), .A2(SI_13_), .B1(n12613), .B2(n9280), .ZN(
        n9212) );
  INV_X1 U11709 ( .A(n9212), .ZN(n9213) );
  NAND2_X1 U11710 ( .A1(n9214), .A2(n9213), .ZN(n14457) );
  NAND2_X1 U11711 ( .A1(n9473), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n9220) );
  NOR2_X1 U11712 ( .A1(n9216), .A2(n9215), .ZN(n9217) );
  OR2_X1 U11713 ( .A1(n9232), .A2(n9217), .ZN(n11546) );
  NAND2_X1 U11714 ( .A1(n9286), .A2(n11546), .ZN(n9219) );
  NAND2_X1 U11715 ( .A1(n9083), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n9218) );
  NAND4_X1 U11716 ( .A1(n9221), .A2(n9220), .A3(n9219), .A4(n9218), .ZN(n14438) );
  OR2_X1 U11717 ( .A1(n14457), .A2(n14438), .ZN(n9574) );
  NAND2_X1 U11718 ( .A1(n14457), .A2(n14438), .ZN(n9575) );
  INV_X1 U11719 ( .A(n14438), .ZN(n11637) );
  NAND2_X1 U11720 ( .A1(n14457), .A2(n11637), .ZN(n9222) );
  XNOR2_X1 U11721 ( .A(n9224), .B(n7243), .ZN(n9964) );
  NAND2_X1 U11722 ( .A1(n9964), .A2(n6437), .ZN(n9230) );
  INV_X1 U11723 ( .A(SI_14_), .ZN(n9966) );
  XNOR2_X1 U11724 ( .A(n9227), .B(n9226), .ZN(n15032) );
  OAI22_X1 U11725 ( .A1(n6440), .A2(n9966), .B1(n9280), .B2(n15032), .ZN(n9228) );
  INV_X1 U11726 ( .A(n9228), .ZN(n9229) );
  NAND2_X1 U11727 ( .A1(n9083), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9237) );
  NAND2_X1 U11728 ( .A1(n9231), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n9236) );
  NOR2_X1 U11729 ( .A1(n9232), .A2(n11642), .ZN(n9233) );
  OR2_X1 U11730 ( .A1(n9247), .A2(n9233), .ZN(n11641) );
  NAND2_X1 U11731 ( .A1(n9286), .A2(n11641), .ZN(n9235) );
  NAND2_X1 U11732 ( .A1(n9473), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9234) );
  NAND2_X1 U11733 ( .A1(n14456), .A2(n11751), .ZN(n9579) );
  NAND2_X1 U11734 ( .A1(n9581), .A2(n9579), .ZN(n11650) );
  INV_X1 U11735 ( .A(n11751), .ZN(n9971) );
  NAND2_X1 U11736 ( .A1(n14456), .A2(n9971), .ZN(n9238) );
  XNOR2_X1 U11737 ( .A(n9240), .B(n7246), .ZN(n10038) );
  NAND2_X1 U11738 ( .A1(n10038), .A2(n9059), .ZN(n9245) );
  NAND2_X1 U11739 ( .A1(n9241), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9242) );
  XNOR2_X1 U11740 ( .A(n9242), .B(n7317), .ZN(n14376) );
  OAI22_X1 U11741 ( .A1(n6440), .A2(n10040), .B1(n9280), .B2(n14376), .ZN(
        n9243) );
  INV_X1 U11742 ( .A(n9243), .ZN(n9244) );
  NAND2_X1 U11743 ( .A1(n9083), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n9253) );
  NAND2_X1 U11744 ( .A1(n9231), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9252) );
  OR2_X1 U11745 ( .A1(n9247), .A2(n9246), .ZN(n9248) );
  NAND2_X1 U11746 ( .A1(n9249), .A2(n9248), .ZN(n11755) );
  NAND2_X1 U11747 ( .A1(n9286), .A2(n11755), .ZN(n9251) );
  NAND2_X1 U11748 ( .A1(n9473), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n9250) );
  OR2_X1 U11749 ( .A1(n11754), .A2(n12828), .ZN(n9583) );
  NAND2_X1 U11750 ( .A1(n11754), .A2(n12828), .ZN(n9580) );
  NAND2_X1 U11751 ( .A1(n11754), .A2(n12547), .ZN(n9254) );
  INV_X1 U11752 ( .A(n12824), .ZN(n9255) );
  OR2_X1 U11753 ( .A1(n12832), .A2(n12812), .ZN(n9585) );
  NAND2_X1 U11754 ( .A1(n12832), .A2(n12812), .ZN(n9586) );
  NAND2_X1 U11755 ( .A1(n12929), .A2(n12545), .ZN(n9257) );
  XNOR2_X1 U11756 ( .A(n9259), .B(n9258), .ZN(n10368) );
  NAND2_X1 U11757 ( .A1(n10368), .A2(n6437), .ZN(n9263) );
  NAND2_X1 U11758 ( .A1(n9277), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9260) );
  XNOR2_X1 U11759 ( .A(n9260), .B(P3_IR_REG_18__SCAN_IN), .ZN(n14420) );
  OAI22_X1 U11760 ( .A1(n6440), .A2(n10370), .B1(n9280), .B2(n12634), .ZN(
        n9261) );
  INV_X1 U11761 ( .A(n9261), .ZN(n9262) );
  NAND2_X1 U11762 ( .A1(n9083), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9265) );
  NAND2_X1 U11763 ( .A1(n9038), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n9264) );
  AND2_X1 U11764 ( .A1(n9265), .A2(n9264), .ZN(n9271) );
  NOR2_X1 U11765 ( .A1(n9267), .A2(n9266), .ZN(n9268) );
  OR2_X1 U11766 ( .A1(n9284), .A2(n9268), .ZN(n12515) );
  NAND2_X1 U11767 ( .A1(n12515), .A2(n9286), .ZN(n9270) );
  NAND2_X1 U11768 ( .A1(n9473), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9269) );
  NAND2_X1 U11769 ( .A1(n12925), .A2(n12813), .ZN(n9597) );
  NAND2_X1 U11770 ( .A1(n9273), .A2(n9272), .ZN(n12792) );
  OR2_X1 U11771 ( .A1(n12925), .A2(n12544), .ZN(n9274) );
  XNOR2_X1 U11772 ( .A(n9276), .B(n9275), .ZN(n10428) );
  NAND2_X1 U11773 ( .A1(n10428), .A2(n9059), .ZN(n9283) );
  INV_X1 U11774 ( .A(n9277), .ZN(n9278) );
  NAND2_X1 U11775 ( .A1(n9375), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9279) );
  OAI22_X1 U11776 ( .A1(n6440), .A2(n7091), .B1(n12596), .B2(n9280), .ZN(n9281) );
  INV_X1 U11777 ( .A(n9281), .ZN(n9282) );
  OR2_X1 U11778 ( .A1(n9284), .A2(n12451), .ZN(n9285) );
  NAND2_X1 U11779 ( .A1(n9296), .A2(n9285), .ZN(n12788) );
  NAND2_X1 U11780 ( .A1(n12788), .A2(n9286), .ZN(n9289) );
  NAND2_X1 U11781 ( .A1(n9473), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n9287) );
  OR2_X1 U11782 ( .A1(n12455), .A2(n12796), .ZN(n9599) );
  NAND2_X1 U11783 ( .A1(n12455), .A2(n12796), .ZN(n9598) );
  NAND2_X1 U11784 ( .A1(n9599), .A2(n9598), .ZN(n12786) );
  XNOR2_X1 U11785 ( .A(n9293), .B(n9292), .ZN(n10582) );
  NAND2_X1 U11786 ( .A1(n10582), .A2(n6437), .ZN(n9295) );
  OR2_X1 U11787 ( .A1(n6440), .A2(n10583), .ZN(n9294) );
  NAND2_X1 U11788 ( .A1(n9296), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9297) );
  NAND2_X1 U11789 ( .A1(n9298), .A2(n9297), .ZN(n12775) );
  NAND2_X1 U11790 ( .A1(n12775), .A2(n9286), .ZN(n9301) );
  AOI22_X1 U11791 ( .A1(n9473), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n9083), .B2(
        P3_REG1_REG_20__SCAN_IN), .ZN(n9300) );
  NAND2_X1 U11792 ( .A1(n9038), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n9299) );
  NAND2_X1 U11793 ( .A1(n12774), .A2(n12782), .ZN(n9603) );
  NAND2_X1 U11794 ( .A1(n9604), .A2(n9603), .ZN(n12773) );
  OR2_X1 U11795 ( .A1(n12762), .A2(n12769), .ZN(n9607) );
  NAND2_X1 U11796 ( .A1(n12762), .A2(n12769), .ZN(n9608) );
  NAND2_X1 U11797 ( .A1(n12756), .A2(n12760), .ZN(n12755) );
  XNOR2_X1 U11798 ( .A(n9303), .B(n9302), .ZN(n10961) );
  NAND2_X1 U11799 ( .A1(n10961), .A2(n6437), .ZN(n9305) );
  OR2_X1 U11800 ( .A1(n6440), .A2(n7386), .ZN(n9304) );
  NAND2_X1 U11801 ( .A1(n9306), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9307) );
  NAND2_X1 U11802 ( .A1(n9319), .A2(n9307), .ZN(n12750) );
  NAND2_X1 U11803 ( .A1(n12750), .A2(n9286), .ZN(n9313) );
  INV_X1 U11804 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n9310) );
  NAND2_X1 U11805 ( .A1(n9083), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9309) );
  NAND2_X1 U11806 ( .A1(n9231), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n9308) );
  OAI211_X1 U11807 ( .C1(n9310), .C2(n9361), .A(n9309), .B(n9308), .ZN(n9311)
         );
  INV_X1 U11808 ( .A(n9311), .ZN(n9312) );
  NAND2_X1 U11809 ( .A1(n9313), .A2(n9312), .ZN(n12758) );
  NAND2_X1 U11810 ( .A1(n12510), .A2(n12758), .ZN(n9314) );
  INV_X1 U11811 ( .A(n12758), .ZN(n12444) );
  XNOR2_X1 U11812 ( .A(n9316), .B(n9315), .ZN(n11107) );
  NAND2_X1 U11813 ( .A1(n11107), .A2(n9059), .ZN(n9318) );
  INV_X1 U11814 ( .A(SI_23_), .ZN(n11110) );
  NAND2_X1 U11815 ( .A1(n9319), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9320) );
  NAND2_X1 U11816 ( .A1(n9328), .A2(n9320), .ZN(n12739) );
  NAND2_X1 U11817 ( .A1(n12739), .A2(n9286), .ZN(n9325) );
  NAND2_X1 U11818 ( .A1(n9473), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9323) );
  NAND2_X1 U11819 ( .A1(n9083), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9322) );
  NAND2_X1 U11820 ( .A1(n9038), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n9321) );
  AND3_X1 U11821 ( .A1(n9323), .A2(n9322), .A3(n9321), .ZN(n9324) );
  XNOR2_X1 U11822 ( .A(n12446), .B(n12504), .ZN(n9615) );
  INV_X1 U11823 ( .A(n9615), .ZN(n12737) );
  INV_X1 U11824 ( .A(n12504), .ZN(n12747) );
  XOR2_X1 U11825 ( .A(n8952), .B(n9326), .Z(n11399) );
  INV_X1 U11826 ( .A(SI_24_), .ZN(n11398) );
  MUX2_X1 U11827 ( .A(n11399), .B(n11398), .S(n9831), .Z(n9327) );
  INV_X1 U11828 ( .A(n12851), .ZN(n12493) );
  NAND2_X1 U11829 ( .A1(n9328), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9329) );
  NAND2_X1 U11830 ( .A1(n9330), .A2(n9329), .ZN(n12723) );
  NAND2_X1 U11831 ( .A1(n12723), .A2(n9286), .ZN(n9335) );
  INV_X1 U11832 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12724) );
  NAND2_X1 U11833 ( .A1(n9083), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9332) );
  NAND2_X1 U11834 ( .A1(n9038), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n9331) );
  OAI211_X1 U11835 ( .C1(n12724), .C2(n9361), .A(n9332), .B(n9331), .ZN(n9333)
         );
  INV_X1 U11836 ( .A(n9333), .ZN(n9334) );
  NAND2_X1 U11837 ( .A1(n12493), .A2(n12734), .ZN(n9618) );
  NAND2_X1 U11838 ( .A1(n12851), .A2(n12702), .ZN(n12707) );
  NAND2_X1 U11839 ( .A1(n9618), .A2(n12707), .ZN(n12728) );
  NAND2_X1 U11840 ( .A1(n12716), .A2(n12728), .ZN(n12721) );
  XNOR2_X1 U11841 ( .A(n12847), .B(n12719), .ZN(n12708) );
  NAND2_X1 U11842 ( .A1(n12699), .A2(n12708), .ZN(n12705) );
  OAI21_X2 U11843 ( .B1(n12719), .B2(n12713), .A(n12705), .ZN(n12687) );
  AOI22_X1 U11844 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n13641), .B2(n15193), .ZN(n9352) );
  INV_X1 U11845 ( .A(n9352), .ZN(n9338) );
  XNOR2_X1 U11846 ( .A(n9353), .B(n9338), .ZN(n12393) );
  NAND2_X1 U11847 ( .A1(n12393), .A2(n6437), .ZN(n9341) );
  OR2_X1 U11848 ( .A1(n6440), .A2(n12394), .ZN(n9340) );
  INV_X1 U11849 ( .A(n9343), .ZN(n9342) );
  INV_X1 U11850 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n12436) );
  NAND2_X1 U11851 ( .A1(n9342), .A2(n12436), .ZN(n9357) );
  NAND2_X1 U11852 ( .A1(n9343), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9344) );
  NAND2_X1 U11853 ( .A1(n9357), .A2(n9344), .ZN(n12680) );
  NAND2_X1 U11854 ( .A1(n12680), .A2(n9286), .ZN(n9350) );
  INV_X1 U11855 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n9347) );
  NAND2_X1 U11856 ( .A1(n9231), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n9346) );
  NAND2_X1 U11857 ( .A1(n9083), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9345) );
  OAI211_X1 U11858 ( .C1(n9361), .C2(n9347), .A(n9346), .B(n9345), .ZN(n9348)
         );
  INV_X1 U11859 ( .A(n9348), .ZN(n9349) );
  NAND2_X1 U11860 ( .A1(n12839), .A2(n12690), .ZN(n9651) );
  OR2_X1 U11861 ( .A1(n12839), .A2(n12690), .ZN(n9351) );
  AOI22_X1 U11862 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(
        P1_DATAO_REG_28__SCAN_IN), .B1(n13638), .B2(n14194), .ZN(n9363) );
  INV_X1 U11863 ( .A(n9363), .ZN(n9354) );
  XNOR2_X1 U11864 ( .A(n9364), .B(n9354), .ZN(n12955) );
  NAND2_X1 U11865 ( .A1(n12955), .A2(n9059), .ZN(n9356) );
  OR2_X1 U11866 ( .A1(n6440), .A2(n12957), .ZN(n9355) );
  NAND2_X1 U11867 ( .A1(n9357), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9358) );
  NAND2_X1 U11868 ( .A1(n9368), .A2(n9358), .ZN(n12666) );
  INV_X1 U11869 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n15295) );
  NAND2_X1 U11870 ( .A1(n9083), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9360) );
  NAND2_X1 U11871 ( .A1(n9038), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n9359) );
  OAI211_X1 U11872 ( .C1(n15295), .C2(n9361), .A(n9360), .B(n9359), .ZN(n9362)
         );
  NAND2_X1 U11873 ( .A1(n12200), .A2(n12674), .ZN(n9396) );
  NAND2_X1 U11874 ( .A1(n9655), .A2(n12194), .ZN(n9654) );
  NAND2_X1 U11875 ( .A1(n9654), .A2(n7567), .ZN(n9374) );
  AOI22_X1 U11876 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n13633), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n7677), .ZN(n9365) );
  XNOR2_X1 U11877 ( .A(n9470), .B(n9365), .ZN(n12951) );
  NAND2_X1 U11878 ( .A1(n12951), .A2(n9059), .ZN(n9367) );
  OR2_X1 U11879 ( .A1(n6440), .A2(n12954), .ZN(n9366) );
  NAND2_X1 U11880 ( .A1(n11854), .A2(n9286), .ZN(n9478) );
  NAND2_X1 U11881 ( .A1(n9473), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9370) );
  NAND2_X1 U11882 ( .A1(n9038), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9369) );
  OAI211_X1 U11883 ( .C1(n9465), .C2(n8964), .A(n9370), .B(n9369), .ZN(n9371)
         );
  INV_X1 U11884 ( .A(n9371), .ZN(n9372) );
  NAND2_X1 U11885 ( .A1(n12423), .A2(n12196), .ZN(n9491) );
  NAND2_X1 U11886 ( .A1(n9636), .A2(n9491), .ZN(n9514) );
  XNOR2_X1 U11887 ( .A(n9374), .B(n9373), .ZN(n9395) );
  NAND2_X1 U11888 ( .A1(n9413), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9378) );
  NAND2_X1 U11889 ( .A1(n10962), .A2(n12659), .ZN(n9460) );
  NAND2_X1 U11890 ( .A1(n9379), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9380) );
  INV_X1 U11891 ( .A(n10585), .ZN(n9442) );
  NAND2_X1 U11892 ( .A1(n10724), .A2(n9442), .ZN(n9496) );
  OR2_X1 U11893 ( .A1(n9384), .A2(n12628), .ZN(n10413) );
  NAND2_X1 U11894 ( .A1(n10413), .A2(n9280), .ZN(n9391) );
  INV_X1 U11895 ( .A(n9391), .ZN(n9386) );
  NAND2_X1 U11896 ( .A1(n9473), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9389) );
  NAND2_X1 U11897 ( .A1(n9083), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9388) );
  AND3_X1 U11898 ( .A1(n9389), .A2(n9388), .A3(n9387), .ZN(n9390) );
  AND2_X1 U11899 ( .A1(n9478), .A2(n9390), .ZN(n9490) );
  INV_X1 U11900 ( .A(P3_B_REG_SCAN_IN), .ZN(n9392) );
  OR2_X1 U11901 ( .A1(n9384), .A2(n9392), .ZN(n9393) );
  NAND2_X1 U11902 ( .A1(n14437), .A2(n9393), .ZN(n11852) );
  OAI22_X1 U11903 ( .A1(n12674), .A2(n15084), .B1(n9490), .B2(n11852), .ZN(
        n9394) );
  NAND2_X1 U11904 ( .A1(n9396), .A2(n9651), .ZN(n9634) );
  INV_X1 U11905 ( .A(n10802), .ZN(n10834) );
  NAND2_X1 U11906 ( .A1(n10914), .A2(n9521), .ZN(n10483) );
  NAND2_X1 U11907 ( .A1(n10483), .A2(n9525), .ZN(n15076) );
  NAND2_X1 U11908 ( .A1(n15076), .A2(n9523), .ZN(n9397) );
  NAND2_X1 U11909 ( .A1(n9397), .A2(n9530), .ZN(n10717) );
  INV_X1 U11910 ( .A(n15064), .ZN(n9500) );
  NAND2_X1 U11911 ( .A1(n10889), .A2(n10890), .ZN(n9398) );
  NAND2_X1 U11912 ( .A1(n9398), .A2(n9544), .ZN(n15045) );
  NAND2_X1 U11913 ( .A1(n15045), .A2(n15051), .ZN(n9399) );
  NAND2_X1 U11914 ( .A1(n9399), .A2(n9549), .ZN(n10876) );
  INV_X1 U11915 ( .A(n11055), .ZN(n9548) );
  NAND2_X1 U11916 ( .A1(n10876), .A2(n9548), .ZN(n9400) );
  NAND2_X1 U11917 ( .A1(n9400), .A2(n9550), .ZN(n11045) );
  NAND2_X1 U11918 ( .A1(n11097), .A2(n9553), .ZN(n9401) );
  NOR2_X1 U11919 ( .A1(n12550), .A2(n15135), .ZN(n9559) );
  NAND2_X1 U11920 ( .A1(n12550), .A2(n15135), .ZN(n9561) );
  INV_X1 U11921 ( .A(n11226), .ZN(n9563) );
  NAND2_X1 U11922 ( .A1(n12549), .A2(n11356), .ZN(n9565) );
  XNOR2_X1 U11923 ( .A(n11571), .B(n14436), .ZN(n11433) );
  NAND2_X1 U11924 ( .A1(n7546), .A2(n6961), .ZN(n11437) );
  NAND2_X1 U11925 ( .A1(n11394), .A2(n11348), .ZN(n9568) );
  NAND2_X2 U11926 ( .A1(n11437), .A2(n9568), .ZN(n14442) );
  INV_X1 U11927 ( .A(n9574), .ZN(n9403) );
  INV_X1 U11928 ( .A(n11748), .ZN(n11752) );
  NAND2_X1 U11929 ( .A1(n11753), .A2(n11752), .ZN(n9404) );
  NAND2_X1 U11930 ( .A1(n9404), .A2(n9580), .ZN(n12830) );
  NAND2_X1 U11931 ( .A1(n12510), .A2(n12444), .ZN(n9610) );
  OR2_X1 U11932 ( .A1(n12510), .A2(n12444), .ZN(n9611) );
  NAND2_X1 U11933 ( .A1(n12907), .A2(n12504), .ZN(n9617) );
  NAND2_X1 U11934 ( .A1(n9408), .A2(n9617), .ZN(n12727) );
  INV_X1 U11935 ( .A(n12708), .ZN(n12700) );
  NAND2_X1 U11936 ( .A1(n12847), .A2(n12719), .ZN(n9625) );
  NAND2_X1 U11937 ( .A1(n12695), .A2(n12703), .ZN(n9628) );
  XOR2_X1 U11938 ( .A(n9488), .B(n9514), .Z(n12427) );
  NAND2_X1 U11939 ( .A1(n10714), .A2(n10585), .ZN(n9456) );
  XNOR2_X1 U11940 ( .A(n9456), .B(n10962), .ZN(n9411) );
  NAND2_X1 U11941 ( .A1(n10714), .A2(n12596), .ZN(n9410) );
  NAND2_X1 U11942 ( .A1(n9411), .A2(n9410), .ZN(n10380) );
  AND2_X1 U11943 ( .A1(n10380), .A2(n15136), .ZN(n10614) );
  NAND2_X1 U11944 ( .A1(n10585), .A2(n12596), .ZN(n9459) );
  INV_X1 U11945 ( .A(n9459), .ZN(n9645) );
  NAND2_X1 U11946 ( .A1(n10614), .A2(n9645), .ZN(n9412) );
  OR3_X1 U11947 ( .A1(n9457), .A2(n12659), .A3(n10585), .ZN(n9455) );
  NAND2_X1 U11948 ( .A1(n9457), .A2(n10905), .ZN(n15137) );
  NAND2_X1 U11949 ( .A1(n12431), .A2(n7571), .ZN(n9464) );
  NAND2_X1 U11950 ( .A1(n9418), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9419) );
  XNOR2_X1 U11951 ( .A(n9419), .B(P3_IR_REG_25__SCAN_IN), .ZN(n9422) );
  AND2_X1 U11952 ( .A1(n9422), .A2(n9421), .ZN(n9420) );
  OR2_X1 U11953 ( .A1(n10396), .A2(n9459), .ZN(n10388) );
  INV_X1 U11954 ( .A(n9421), .ZN(n11400) );
  INV_X1 U11955 ( .A(n9422), .ZN(n11525) );
  INV_X1 U11956 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9423) );
  NAND2_X1 U11957 ( .A1(n9973), .A2(n9423), .ZN(n9426) );
  NAND2_X1 U11958 ( .A1(n6679), .A2(n11525), .ZN(n9425) );
  NAND2_X1 U11959 ( .A1(n9426), .A2(n9425), .ZN(n9887) );
  INV_X1 U11960 ( .A(n9973), .ZN(n9437) );
  NOR4_X1 U11961 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n9435) );
  NOR4_X1 U11962 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n9430) );
  NOR4_X1 U11963 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n9429) );
  NOR4_X1 U11964 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9428) );
  NOR4_X1 U11965 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n9427) );
  NAND4_X1 U11966 ( .A1(n9430), .A2(n9429), .A3(n9428), .A4(n9427), .ZN(n9431)
         );
  NOR4_X1 U11967 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        n9432), .A4(n9431), .ZN(n9434) );
  NOR4_X1 U11968 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n9433) );
  AND3_X1 U11969 ( .A1(n9435), .A2(n9434), .A3(n9433), .ZN(n9436) );
  OR2_X1 U11970 ( .A1(n9887), .A2(n9454), .ZN(n9441) );
  INV_X1 U11971 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9438) );
  NAND2_X1 U11972 ( .A1(n6679), .A2(n11400), .ZN(n9439) );
  NAND2_X1 U11973 ( .A1(n10376), .A2(n10391), .ZN(n9448) );
  INV_X1 U11974 ( .A(n9460), .ZN(n9443) );
  NAND2_X1 U11975 ( .A1(n10714), .A2(n9442), .ZN(n10480) );
  INV_X1 U11976 ( .A(n10480), .ZN(n9516) );
  NAND2_X1 U11977 ( .A1(n9443), .A2(n9516), .ZN(n10383) );
  INV_X1 U11978 ( .A(n10391), .ZN(n10379) );
  INV_X1 U11979 ( .A(n9454), .ZN(n9444) );
  NAND2_X1 U11980 ( .A1(n10380), .A2(n10492), .ZN(n9445) );
  OAI21_X1 U11981 ( .B1(n10383), .B2(n10379), .A(n9445), .ZN(n9446) );
  INV_X1 U11982 ( .A(n10396), .ZN(n10373) );
  NAND2_X1 U11983 ( .A1(n9446), .A2(n10373), .ZN(n9447) );
  INV_X1 U11984 ( .A(n12423), .ZN(n9466) );
  NOR2_X1 U11985 ( .A1(n9466), .A2(n12939), .ZN(n9449) );
  NOR2_X1 U11986 ( .A1(n9449), .A2(n7560), .ZN(n9451) );
  NAND2_X1 U11987 ( .A1(n10398), .A2(n9459), .ZN(n10378) );
  NAND2_X1 U11988 ( .A1(n9633), .A2(n9455), .ZN(n10719) );
  NAND2_X1 U11989 ( .A1(n10378), .A2(n10719), .ZN(n10721) );
  INV_X1 U11990 ( .A(n10479), .ZN(n12942) );
  NAND2_X1 U11991 ( .A1(n9457), .A2(n9456), .ZN(n9458) );
  NAND3_X1 U11992 ( .A1(n9460), .A2(n9459), .A3(n9458), .ZN(n9461) );
  NAND3_X1 U11993 ( .A1(n9461), .A2(n9633), .A3(n9887), .ZN(n9462) );
  OAI21_X1 U11994 ( .B1(n10721), .B2(n12942), .A(n9462), .ZN(n9463) );
  NAND2_X1 U11995 ( .A1(n9464), .A2(n15157), .ZN(n9468) );
  OR2_X1 U11996 ( .A1(n15157), .A2(n9465), .ZN(n9467) );
  NAND3_X1 U11997 ( .A1(n9468), .A2(n9467), .A3(n7547), .ZN(P3_U3488) );
  INV_X1 U11998 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13630) );
  INV_X1 U11999 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12153) );
  AOI22_X1 U12000 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(
        P1_DATAO_REG_30__SCAN_IN), .B1(n13630), .B2(n12153), .ZN(n9471) );
  NAND2_X1 U12001 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n7677), .ZN(n9469) );
  INV_X1 U12002 ( .A(n6437), .ZN(n9472) );
  INV_X1 U12003 ( .A(n9490), .ZN(n12540) );
  NAND2_X1 U12004 ( .A1(n12664), .A2(n12540), .ZN(n9498) );
  INV_X1 U12005 ( .A(n9498), .ZN(n9479) );
  NAND2_X1 U12006 ( .A1(n9473), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n9476) );
  NAND2_X1 U12007 ( .A1(n9083), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n9475) );
  NAND2_X1 U12008 ( .A1(n9038), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n9474) );
  AND3_X1 U12009 ( .A1(n9476), .A2(n9475), .A3(n9474), .ZN(n9477) );
  NAND2_X1 U12010 ( .A1(n9478), .A2(n9477), .ZN(n12539) );
  INV_X1 U12011 ( .A(n12539), .ZN(n9485) );
  NOR2_X1 U12012 ( .A1(n9479), .A2(n9485), .ZN(n9494) );
  NAND2_X1 U12013 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n13630), .ZN(n9480) );
  INV_X1 U12014 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13625) );
  INV_X1 U12015 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9923) );
  AOI22_X1 U12016 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(n13625), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(n9923), .ZN(n9482) );
  XNOR2_X1 U12017 ( .A(n9483), .B(n9482), .ZN(n12943) );
  INV_X1 U12018 ( .A(SI_31_), .ZN(n12947) );
  NOR2_X1 U12019 ( .A1(n6440), .A2(n12947), .ZN(n9484) );
  INV_X1 U12020 ( .A(n9636), .ZN(n9489) );
  NAND2_X1 U12021 ( .A1(n14452), .A2(n9485), .ZN(n9487) );
  OAI211_X1 U12022 ( .C1(n9489), .C2(n9488), .A(n9487), .B(n9513), .ZN(n9493)
         );
  NAND2_X1 U12023 ( .A1(n14452), .A2(n9490), .ZN(n9499) );
  AND2_X1 U12024 ( .A1(n9499), .A2(n9491), .ZN(n9641) );
  INV_X1 U12025 ( .A(n9641), .ZN(n9492) );
  OAI22_X1 U12026 ( .A1(n9494), .A2(n9486), .B1(n9493), .B2(n9492), .ZN(n9495)
         );
  XNOR2_X1 U12027 ( .A(n9495), .B(n12596), .ZN(n9497) );
  NOR2_X1 U12028 ( .A1(n9497), .A2(n9496), .ZN(n9648) );
  INV_X1 U12029 ( .A(n9499), .ZN(n9515) );
  NAND2_X1 U12030 ( .A1(n9611), .A2(n9610), .ZN(n12748) );
  NAND4_X1 U12031 ( .A1(n9523), .A2(n9500), .A3(n9548), .A4(n10890), .ZN(n9504) );
  NAND2_X1 U12032 ( .A1(n12560), .A2(n10834), .ZN(n9518) );
  INV_X1 U12033 ( .A(n9518), .ZN(n9501) );
  NOR2_X1 U12034 ( .A1(n10914), .A2(n9501), .ZN(n10616) );
  INV_X1 U12035 ( .A(n9502), .ZN(n10915) );
  NAND4_X1 U12036 ( .A1(n10616), .A2(n10915), .A3(n10718), .A4(n15051), .ZN(
        n9503) );
  NOR4_X1 U12037 ( .A1(n9504), .A2(n9503), .A3(n9147), .A4(n11174), .ZN(n9505)
         );
  NAND4_X1 U12038 ( .A1(n9505), .A2(n9563), .A3(n14441), .A4(n6961), .ZN(n9507) );
  INV_X1 U12039 ( .A(n11673), .ZN(n9506) );
  NOR4_X1 U12040 ( .A1(n11748), .A2(n11650), .A3(n9507), .A4(n9506), .ZN(n9508) );
  NAND4_X1 U12041 ( .A1(n12793), .A2(n12831), .A3(n12817), .A4(n9508), .ZN(
        n9509) );
  NOR4_X1 U12042 ( .A1(n12773), .A2(n12786), .A3(n12748), .A4(n9509), .ZN(
        n9510) );
  NAND4_X1 U12043 ( .A1(n9615), .A2(n9606), .A3(n12688), .A4(n9510), .ZN(n9511) );
  NOR3_X1 U12044 ( .A1(n9511), .A2(n12708), .A3(n12728), .ZN(n9512) );
  NAND2_X1 U12045 ( .A1(n9517), .A2(n9516), .ZN(n9646) );
  AND2_X1 U12046 ( .A1(n9521), .A2(n9518), .ZN(n9520) );
  OAI21_X1 U12047 ( .B1(n10914), .B2(n10724), .A(n9518), .ZN(n9519) );
  MUX2_X1 U12048 ( .A(n9520), .B(n9519), .S(n9633), .Z(n9526) );
  MUX2_X1 U12049 ( .A(n9521), .B(n9525), .S(n10398), .Z(n9522) );
  NAND2_X1 U12050 ( .A1(n9523), .A2(n9522), .ZN(n9524) );
  AOI21_X1 U12051 ( .B1(n9526), .B2(n9525), .A(n9524), .ZN(n9529) );
  AOI21_X1 U12052 ( .B1(n9535), .B2(n9527), .A(n9633), .ZN(n9528) );
  OAI21_X1 U12053 ( .B1(n9529), .B2(n9528), .A(n9531), .ZN(n9534) );
  NAND2_X1 U12054 ( .A1(n9531), .A2(n9530), .ZN(n9532) );
  NAND2_X1 U12055 ( .A1(n9532), .A2(n9633), .ZN(n9533) );
  NAND2_X1 U12056 ( .A1(n9534), .A2(n9533), .ZN(n9538) );
  NOR2_X1 U12057 ( .A1(n9535), .A2(n10398), .ZN(n9536) );
  NOR2_X1 U12058 ( .A1(n15064), .A2(n9536), .ZN(n9537) );
  NAND2_X1 U12059 ( .A1(n9538), .A2(n9537), .ZN(n9543) );
  NAND3_X1 U12060 ( .A1(n9543), .A2(n10890), .A3(n9539), .ZN(n9541) );
  NAND3_X1 U12061 ( .A1(n9543), .A2(n10890), .A3(n9542), .ZN(n9547) );
  INV_X1 U12062 ( .A(n9545), .ZN(n9546) );
  MUX2_X1 U12063 ( .A(n9551), .B(n9550), .S(n10398), .Z(n9552) );
  INV_X1 U12064 ( .A(n11174), .ZN(n9557) );
  NAND2_X1 U12065 ( .A1(n9633), .A2(n9553), .ZN(n9555) );
  NAND2_X1 U12066 ( .A1(n10398), .A2(n11214), .ZN(n9554) );
  MUX2_X1 U12067 ( .A(n9555), .B(n9554), .S(n12551), .Z(n9556) );
  NAND3_X1 U12068 ( .A1(n9558), .A2(n9557), .A3(n9556), .ZN(n9564) );
  INV_X1 U12069 ( .A(n9559), .ZN(n9560) );
  MUX2_X1 U12070 ( .A(n9561), .B(n9560), .S(n10398), .Z(n9562) );
  INV_X1 U12071 ( .A(n12549), .ZN(n11436) );
  NAND2_X1 U12072 ( .A1(n11436), .A2(n11362), .ZN(n9566) );
  MUX2_X1 U12073 ( .A(n9566), .B(n9565), .S(n10398), .Z(n9567) );
  AOI21_X1 U12074 ( .B1(n9572), .B2(n9568), .A(n10398), .ZN(n9569) );
  OAI21_X1 U12075 ( .B1(n11394), .B2(n11348), .A(n9570), .ZN(n9571) );
  OAI21_X1 U12076 ( .B1(n9572), .B2(n9633), .A(n11673), .ZN(n9573) );
  MUX2_X1 U12077 ( .A(n9575), .B(n9574), .S(n9633), .Z(n9576) );
  INV_X1 U12078 ( .A(n9576), .ZN(n9577) );
  OR3_X1 U12079 ( .A1(n9578), .A2(n9577), .A3(n11650), .ZN(n9582) );
  AND2_X1 U12080 ( .A1(n9585), .A2(n9583), .ZN(n9584) );
  MUX2_X1 U12081 ( .A(n9586), .B(n9585), .S(n10398), .Z(n9587) );
  NAND2_X1 U12082 ( .A1(n9588), .A2(n12817), .ZN(n9596) );
  INV_X1 U12083 ( .A(n9597), .ZN(n9591) );
  OAI211_X1 U12084 ( .C1(n9591), .C2(n9590), .A(n9599), .B(n9589), .ZN(n9592)
         );
  INV_X1 U12085 ( .A(n9592), .ZN(n9593) );
  OAI21_X1 U12086 ( .B1(n9596), .B2(n9272), .A(n9593), .ZN(n9594) );
  AOI21_X1 U12087 ( .B1(n9596), .B2(n9595), .A(n9272), .ZN(n9601) );
  NAND2_X1 U12088 ( .A1(n9598), .A2(n9597), .ZN(n9600) );
  OAI21_X1 U12089 ( .B1(n9601), .B2(n9600), .A(n9599), .ZN(n9602) );
  MUX2_X1 U12090 ( .A(n9604), .B(n9603), .S(n10398), .Z(n9605) );
  INV_X1 U12091 ( .A(n12748), .ZN(n12744) );
  MUX2_X1 U12092 ( .A(n9608), .B(n9607), .S(n10398), .Z(n9609) );
  MUX2_X1 U12093 ( .A(n9611), .B(n9610), .S(n10398), .Z(n9612) );
  NAND2_X1 U12094 ( .A1(n9613), .A2(n9612), .ZN(n9616) );
  NOR2_X1 U12095 ( .A1(n12504), .A2(n9633), .ZN(n9614) );
  AOI22_X1 U12096 ( .A1(n9616), .A2(n9615), .B1(n9614), .B2(n12446), .ZN(n9623) );
  NAND2_X1 U12097 ( .A1(n9618), .A2(n9617), .ZN(n9619) );
  NAND3_X1 U12098 ( .A1(n9619), .A2(n12707), .A3(n9633), .ZN(n9622) );
  INV_X1 U12099 ( .A(n12707), .ZN(n9620) );
  NAND2_X1 U12100 ( .A1(n9620), .A2(n10398), .ZN(n9621) );
  OAI211_X1 U12101 ( .C1(n12728), .C2(n9623), .A(n9622), .B(n9621), .ZN(n9627)
         );
  OR2_X1 U12102 ( .A1(n12847), .A2(n12719), .ZN(n9624) );
  MUX2_X1 U12103 ( .A(n9625), .B(n9624), .S(n10398), .Z(n9626) );
  MUX2_X1 U12104 ( .A(n9629), .B(n9628), .S(n10398), .Z(n9630) );
  NOR2_X1 U12105 ( .A1(n12690), .A2(n10398), .ZN(n9631) );
  OAI21_X1 U12106 ( .B1(n9634), .B2(n9633), .A(n9632), .ZN(n9635) );
  NAND2_X1 U12107 ( .A1(n9635), .A2(n9638), .ZN(n9637) );
  OAI211_X1 U12108 ( .C1(n10398), .C2(n9638), .A(n9637), .B(n9636), .ZN(n9640)
         );
  AOI21_X1 U12109 ( .B1(n9641), .B2(n9640), .A(n9639), .ZN(n9643) );
  NOR2_X1 U12110 ( .A1(n9643), .A2(n9642), .ZN(n9644) );
  OR2_X1 U12111 ( .A1(n10397), .A2(P3_U3151), .ZN(n11108) );
  INV_X1 U12112 ( .A(n11108), .ZN(n9647) );
  NOR2_X1 U12113 ( .A1(n10388), .A2(n15084), .ZN(n10493) );
  INV_X1 U12114 ( .A(n9384), .ZN(n10402) );
  NAND2_X1 U12115 ( .A1(n10493), .A2(n10402), .ZN(n9649) );
  OAI211_X1 U12116 ( .C1(n10962), .C2(n11108), .A(n9649), .B(P3_B_REG_SCAN_IN), 
        .ZN(n9650) );
  INV_X1 U12117 ( .A(n9651), .ZN(n9652) );
  NOR2_X1 U12118 ( .A1(n12676), .A2(n9652), .ZN(n9653) );
  XNOR2_X1 U12119 ( .A(n9653), .B(n12194), .ZN(n12669) );
  OAI211_X1 U12120 ( .C1(n9655), .C2(n12194), .A(n9654), .B(n15089), .ZN(n9657) );
  NAND2_X1 U12121 ( .A1(n12541), .A2(n14435), .ZN(n9656) );
  OR2_X1 U12122 ( .A1(n12895), .A2(n15154), .ZN(n9660) );
  INV_X1 U12123 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n15229) );
  INV_X1 U12124 ( .A(n9658), .ZN(n9659) );
  NAND2_X1 U12125 ( .A1(n9660), .A2(n9659), .ZN(P3_U3487) );
  INV_X2 U12126 ( .A(n14858), .ZN(n14859) );
  INV_X1 U12127 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n9663) );
  NAND2_X1 U12128 ( .A1(n10196), .A2(n9775), .ZN(n10030) );
  INV_X1 U12129 ( .A(n12090), .ZN(n9667) );
  AND2_X2 U12130 ( .A1(n9668), .A2(n9667), .ZN(n9676) );
  NAND2_X1 U12131 ( .A1(n11865), .A2(n9676), .ZN(n9669) );
  INV_X1 U12132 ( .A(n9673), .ZN(n9671) );
  NAND2_X1 U12133 ( .A1(n11872), .A2(n9775), .ZN(n9672) );
  INV_X1 U12134 ( .A(n9672), .ZN(n9670) );
  NAND2_X1 U12135 ( .A1(n9671), .A2(n9670), .ZN(n9674) );
  NAND2_X1 U12136 ( .A1(n9673), .A2(n9672), .ZN(n9675) );
  XNOR2_X1 U12137 ( .A(n9676), .B(n14837), .ZN(n9678) );
  NAND2_X1 U12138 ( .A1(n13142), .A2(n9775), .ZN(n9677) );
  NAND2_X1 U12139 ( .A1(n9678), .A2(n9677), .ZN(n9682) );
  INV_X1 U12140 ( .A(n9677), .ZN(n9680) );
  INV_X1 U12141 ( .A(n9678), .ZN(n9679) );
  NAND2_X1 U12142 ( .A1(n9680), .A2(n9679), .ZN(n9681) );
  NAND2_X1 U12143 ( .A1(n13141), .A2(n9775), .ZN(n9683) );
  XNOR2_X1 U12144 ( .A(n9684), .B(n9683), .ZN(n10263) );
  XNOR2_X1 U12145 ( .A(n14844), .B(n9676), .ZN(n9685) );
  NAND2_X1 U12146 ( .A1(n13140), .A2(n9775), .ZN(n9686) );
  NAND2_X1 U12147 ( .A1(n9685), .A2(n9686), .ZN(n9688) );
  NAND2_X1 U12148 ( .A1(n9688), .A2(n9687), .ZN(n10509) );
  XNOR2_X1 U12149 ( .A(n11907), .B(n9676), .ZN(n9689) );
  NAND2_X1 U12150 ( .A1(n13139), .A2(n9775), .ZN(n9690) );
  NAND2_X1 U12151 ( .A1(n9689), .A2(n9690), .ZN(n9694) );
  INV_X1 U12152 ( .A(n9689), .ZN(n9692) );
  INV_X1 U12153 ( .A(n9690), .ZN(n9691) );
  NAND2_X1 U12154 ( .A1(n9692), .A2(n9691), .ZN(n9693) );
  AND2_X1 U12155 ( .A1(n9694), .A2(n9693), .ZN(n10622) );
  NAND2_X1 U12156 ( .A1(n10621), .A2(n10622), .ZN(n10620) );
  NAND2_X1 U12157 ( .A1(n10620), .A2(n9694), .ZN(n13077) );
  XNOR2_X1 U12158 ( .A(n13080), .B(n6840), .ZN(n9695) );
  NAND2_X1 U12159 ( .A1(n13138), .A2(n9775), .ZN(n9696) );
  XNOR2_X1 U12160 ( .A(n9695), .B(n9696), .ZN(n13076) );
  INV_X1 U12161 ( .A(n9695), .ZN(n9698) );
  INV_X1 U12162 ( .A(n9696), .ZN(n9697) );
  NAND2_X1 U12163 ( .A1(n9698), .A2(n9697), .ZN(n9699) );
  XNOR2_X1 U12164 ( .A(n11919), .B(n12990), .ZN(n9702) );
  NAND2_X1 U12165 ( .A1(n13137), .A2(n9775), .ZN(n9700) );
  XNOR2_X1 U12166 ( .A(n9702), .B(n9700), .ZN(n10836) );
  INV_X1 U12167 ( .A(n9700), .ZN(n9701) );
  NAND2_X1 U12168 ( .A1(n9702), .A2(n9701), .ZN(n9703) );
  XNOR2_X1 U12169 ( .A(n11932), .B(n6840), .ZN(n9704) );
  NAND2_X1 U12170 ( .A1(n13136), .A2(n9775), .ZN(n9705) );
  NAND2_X1 U12171 ( .A1(n9704), .A2(n9705), .ZN(n9710) );
  INV_X1 U12172 ( .A(n9704), .ZN(n9707) );
  INV_X1 U12173 ( .A(n9705), .ZN(n9706) );
  NAND2_X1 U12174 ( .A1(n9707), .A2(n9706), .ZN(n9708) );
  NAND2_X1 U12175 ( .A1(n9710), .A2(n9708), .ZN(n11129) );
  XNOR2_X1 U12176 ( .A(n13477), .B(n6840), .ZN(n9711) );
  NAND2_X1 U12177 ( .A1(n13135), .A2(n13460), .ZN(n9712) );
  NAND2_X1 U12178 ( .A1(n9711), .A2(n9712), .ZN(n9716) );
  INV_X1 U12179 ( .A(n9711), .ZN(n9714) );
  INV_X1 U12180 ( .A(n9712), .ZN(n9713) );
  NAND2_X1 U12181 ( .A1(n9714), .A2(n9713), .ZN(n9715) );
  AND2_X1 U12182 ( .A1(n9716), .A2(n9715), .ZN(n11202) );
  XNOR2_X1 U12183 ( .A(n11946), .B(n6840), .ZN(n9718) );
  NAND2_X1 U12184 ( .A1(n13134), .A2(n13460), .ZN(n9717) );
  XNOR2_X1 U12185 ( .A(n9718), .B(n9717), .ZN(n11293) );
  XNOR2_X1 U12186 ( .A(n11953), .B(n6840), .ZN(n9719) );
  NAND2_X1 U12187 ( .A1(n13133), .A2(n13460), .ZN(n9720) );
  NAND2_X1 U12188 ( .A1(n9719), .A2(n9720), .ZN(n11423) );
  NAND2_X1 U12189 ( .A1(n11424), .A2(n11423), .ZN(n9723) );
  INV_X1 U12190 ( .A(n9719), .ZN(n9722) );
  INV_X1 U12191 ( .A(n9720), .ZN(n9721) );
  NAND2_X1 U12192 ( .A1(n9722), .A2(n9721), .ZN(n11422) );
  NAND2_X1 U12193 ( .A1(n9723), .A2(n11422), .ZN(n11574) );
  XNOR2_X1 U12194 ( .A(n11961), .B(n6840), .ZN(n9727) );
  NAND2_X1 U12195 ( .A1(n13131), .A2(n13460), .ZN(n9726) );
  XNOR2_X1 U12196 ( .A(n9727), .B(n9726), .ZN(n11575) );
  INV_X1 U12197 ( .A(n11575), .ZN(n9724) );
  NAND2_X1 U12198 ( .A1(n9727), .A2(n9726), .ZN(n9728) );
  XNOR2_X1 U12199 ( .A(n11969), .B(n12990), .ZN(n9729) );
  AND2_X1 U12200 ( .A1(n13130), .A2(n13460), .ZN(n9730) );
  NAND2_X1 U12201 ( .A1(n9729), .A2(n9730), .ZN(n9734) );
  INV_X1 U12202 ( .A(n9729), .ZN(n9732) );
  INV_X1 U12203 ( .A(n9730), .ZN(n9731) );
  NAND2_X1 U12204 ( .A1(n9732), .A2(n9731), .ZN(n9733) );
  NAND2_X1 U12205 ( .A1(n9734), .A2(n9733), .ZN(n11659) );
  INV_X1 U12206 ( .A(n9734), .ZN(n9735) );
  XNOR2_X1 U12207 ( .A(n11968), .B(n12990), .ZN(n9738) );
  NOR2_X1 U12208 ( .A1(n11967), .A2(n13372), .ZN(n9736) );
  XNOR2_X1 U12209 ( .A(n9738), .B(n9736), .ZN(n11784) );
  INV_X1 U12210 ( .A(n9736), .ZN(n9737) );
  NAND2_X1 U12211 ( .A1(n9738), .A2(n9737), .ZN(n9739) );
  NAND2_X1 U12212 ( .A1(n11783), .A2(n9739), .ZN(n9742) );
  XNOR2_X1 U12213 ( .A(n13617), .B(n12990), .ZN(n9741) );
  XNOR2_X1 U12214 ( .A(n9742), .B(n9741), .ZN(n13105) );
  NOR2_X1 U12215 ( .A1(n9740), .A2(n13372), .ZN(n13104) );
  NAND2_X1 U12216 ( .A1(n13105), .A2(n13104), .ZN(n13103) );
  NAND2_X1 U12217 ( .A1(n13127), .A2(n13460), .ZN(n9743) );
  XNOR2_X1 U12218 ( .A(n13551), .B(n12990), .ZN(n9745) );
  XOR2_X1 U12219 ( .A(n9743), .B(n9745), .Z(n13016) );
  INV_X1 U12220 ( .A(n9743), .ZN(n9744) );
  NOR2_X1 U12221 ( .A1(n9745), .A2(n9744), .ZN(n13024) );
  XNOR2_X1 U12222 ( .A(n11978), .B(n12990), .ZN(n9747) );
  NAND2_X1 U12223 ( .A1(n13126), .A2(n13460), .ZN(n9748) );
  XNOR2_X1 U12224 ( .A(n9747), .B(n9748), .ZN(n13023) );
  XNOR2_X1 U12225 ( .A(n13422), .B(n12990), .ZN(n12975) );
  INV_X1 U12226 ( .A(n12975), .ZN(n9746) );
  NOR2_X1 U12227 ( .A1(n13028), .A2(n13372), .ZN(n9750) );
  AND2_X1 U12228 ( .A1(n9746), .A2(n9750), .ZN(n12976) );
  XNOR2_X1 U12229 ( .A(n13537), .B(n6840), .ZN(n9754) );
  NAND2_X1 U12230 ( .A1(n13125), .A2(n13460), .ZN(n9755) );
  NAND2_X1 U12231 ( .A1(n9754), .A2(n9755), .ZN(n12978) );
  INV_X1 U12232 ( .A(n9747), .ZN(n9749) );
  NAND2_X1 U12233 ( .A1(n9749), .A2(n9748), .ZN(n12973) );
  NAND2_X1 U12234 ( .A1(n12973), .A2(n9750), .ZN(n9752) );
  INV_X1 U12235 ( .A(n12973), .ZN(n9751) );
  INV_X1 U12236 ( .A(n9750), .ZN(n12974) );
  AOI22_X1 U12237 ( .A1(n12975), .A2(n9752), .B1(n9751), .B2(n12974), .ZN(
        n9753) );
  INV_X1 U12238 ( .A(n9754), .ZN(n9757) );
  INV_X1 U12239 ( .A(n9755), .ZN(n9756) );
  NAND2_X1 U12240 ( .A1(n9757), .A2(n9756), .ZN(n12977) );
  XNOR2_X1 U12241 ( .A(n13603), .B(n12990), .ZN(n9759) );
  NAND2_X1 U12242 ( .A1(n13124), .A2(n13460), .ZN(n9758) );
  NAND2_X1 U12243 ( .A1(n9759), .A2(n9758), .ZN(n13046) );
  NOR2_X1 U12244 ( .A1(n9759), .A2(n9758), .ZN(n13048) );
  XNOR2_X1 U12245 ( .A(n13526), .B(n12990), .ZN(n9761) );
  NOR2_X1 U12246 ( .A1(n13059), .A2(n13372), .ZN(n9760) );
  XNOR2_X1 U12247 ( .A(n9761), .B(n9760), .ZN(n13001) );
  NOR2_X1 U12248 ( .A1(n13000), .A2(n13001), .ZN(n12999) );
  NOR2_X1 U12249 ( .A1(n12999), .A2(n7553), .ZN(n9764) );
  XNOR2_X1 U12250 ( .A(n13591), .B(n12990), .ZN(n9762) );
  XNOR2_X1 U12251 ( .A(n9764), .B(n9762), .ZN(n13058) );
  NOR2_X1 U12252 ( .A1(n12030), .A2(n13372), .ZN(n13057) );
  NAND2_X1 U12253 ( .A1(n13058), .A2(n13057), .ZN(n13056) );
  INV_X1 U12254 ( .A(n9762), .ZN(n9763) );
  OR2_X1 U12255 ( .A1(n9764), .A2(n9763), .ZN(n9765) );
  XNOR2_X1 U12256 ( .A(n13587), .B(n12990), .ZN(n9767) );
  NOR2_X1 U12257 ( .A1(n13040), .A2(n13372), .ZN(n12965) );
  XNOR2_X1 U12258 ( .A(n13331), .B(n12990), .ZN(n9769) );
  AND2_X1 U12259 ( .A1(n13120), .A2(n13460), .ZN(n9768) );
  NAND2_X1 U12260 ( .A1(n9769), .A2(n9768), .ZN(n9770) );
  OAI21_X1 U12261 ( .B1(n9769), .B2(n9768), .A(n9770), .ZN(n13037) );
  INV_X1 U12262 ( .A(n9770), .ZN(n9771) );
  XNOR2_X1 U12263 ( .A(n13320), .B(n6840), .ZN(n9773) );
  NOR2_X1 U12264 ( .A1(n13093), .A2(n13372), .ZN(n9772) );
  NAND2_X1 U12265 ( .A1(n9773), .A2(n9772), .ZN(n9774) );
  OAI21_X1 U12266 ( .B1(n9773), .B2(n9772), .A(n9774), .ZN(n13011) );
  XNOR2_X1 U12267 ( .A(n13500), .B(n12990), .ZN(n9778) );
  NAND2_X1 U12268 ( .A1(n13119), .A2(n13460), .ZN(n9776) );
  XNOR2_X1 U12269 ( .A(n9778), .B(n9776), .ZN(n13090) );
  INV_X1 U12270 ( .A(n9776), .ZN(n9777) );
  XNOR2_X1 U12271 ( .A(n13286), .B(n6840), .ZN(n9781) );
  NOR2_X1 U12272 ( .A1(n13095), .A2(n13372), .ZN(n9780) );
  NAND2_X1 U12273 ( .A1(n9781), .A2(n9780), .ZN(n12986) );
  OAI21_X1 U12274 ( .B1(n9781), .B2(n9780), .A(n12986), .ZN(n9783) );
  NAND2_X1 U12275 ( .A1(n9785), .A2(n9784), .ZN(n9797) );
  INV_X1 U12276 ( .A(n9797), .ZN(n9786) );
  AND2_X1 U12277 ( .A1(n9786), .A2(n14835), .ZN(n9795) );
  AND2_X1 U12278 ( .A1(n14853), .A2(n9787), .ZN(n9788) );
  INV_X1 U12279 ( .A(n9795), .ZN(n9792) );
  OAI21_X2 U12280 ( .B1(n9792), .B2(n9791), .A(n13472), .ZN(n13081) );
  INV_X1 U12281 ( .A(n13081), .ZN(n13114) );
  OAI22_X1 U12282 ( .A1(n9793), .A2(n13094), .B1(n12042), .B2(n13092), .ZN(
        n13284) );
  INV_X1 U12283 ( .A(n12053), .ZN(n9794) );
  INV_X1 U12284 ( .A(n13108), .ZN(n13099) );
  NAND2_X1 U12285 ( .A1(n9797), .A2(n9796), .ZN(n9800) );
  AND3_X1 U12286 ( .A1(n9807), .A2(n11742), .A3(n9798), .ZN(n9799) );
  NAND2_X1 U12287 ( .A1(n9800), .A2(n9799), .ZN(n10031) );
  OAI22_X1 U12288 ( .A1(n13288), .A2(n13097), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9801), .ZN(n9802) );
  AOI21_X1 U12289 ( .B1(n13284), .B2(n13099), .A(n9802), .ZN(n9803) );
  INV_X1 U12290 ( .A(n9804), .ZN(n9805) );
  INV_X1 U12291 ( .A(n9807), .ZN(n9808) );
  NAND2_X1 U12292 ( .A1(n9808), .A2(n11742), .ZN(n9894) );
  OR2_X2 U12293 ( .A1(n9894), .A2(P2_U3088), .ZN(n13132) );
  INV_X1 U12294 ( .A(n9809), .ZN(n10377) );
  AND2_X1 U12295 ( .A1(n14207), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9810) );
  INV_X1 U12296 ( .A(n9810), .ZN(n10329) );
  MUX2_X1 U12297 ( .A(n8338), .B(P1_REG2_REG_1__SCAN_IN), .S(n10013), .Z(n9817) );
  MUX2_X1 U12298 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n8338), .S(n10013), .Z(n9811) );
  NAND2_X1 U12299 ( .A1(n9811), .A2(n9810), .ZN(n10015) );
  INV_X1 U12300 ( .A(n10015), .ZN(n9816) );
  NAND2_X1 U12301 ( .A1(n10321), .A2(n11746), .ZN(n9824) );
  NAND2_X1 U12302 ( .A1(n9812), .A2(n10933), .ZN(n9813) );
  NAND2_X1 U12303 ( .A1(n9813), .A2(n8343), .ZN(n9823) );
  INV_X1 U12304 ( .A(n9823), .ZN(n9814) );
  NAND2_X1 U12305 ( .A1(n9824), .A2(n9814), .ZN(n10150) );
  INV_X1 U12306 ( .A(n14197), .ZN(n12383) );
  NAND2_X1 U12307 ( .A1(n10252), .A2(n12383), .ZN(n9815) );
  OR2_X1 U12308 ( .A1(n10150), .A2(n9815), .ZN(n14596) );
  AOI211_X1 U12309 ( .C1(n10329), .C2(n9817), .A(n9816), .B(n14596), .ZN(n9829) );
  NAND2_X1 U12310 ( .A1(n14207), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9822) );
  INV_X1 U12311 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n15162) );
  MUX2_X1 U12312 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n15162), .S(n10013), .Z(
        n9818) );
  INV_X1 U12313 ( .A(n9818), .ZN(n9821) );
  NAND3_X1 U12314 ( .A1(n9818), .A2(n14207), .A3(P1_REG1_REG_0__SCAN_IN), .ZN(
        n10004) );
  INV_X1 U12315 ( .A(n10004), .ZN(n9820) );
  INV_X1 U12316 ( .A(n10150), .ZN(n9819) );
  AOI211_X1 U12317 ( .C1(n9822), .C2(n9821), .A(n9820), .B(n11701), .ZN(n9828)
         );
  INV_X1 U12318 ( .A(n10013), .ZN(n10005) );
  NOR2_X1 U12319 ( .A1(n14601), .A2(n10005), .ZN(n9827) );
  NAND2_X1 U12320 ( .A1(n9824), .A2(n9823), .ZN(n14605) );
  INV_X1 U12321 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9825) );
  OAI22_X1 U12322 ( .A1(n14605), .A2(n15191), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9825), .ZN(n9826) );
  OR4_X1 U12323 ( .A1(n9829), .A2(n9828), .A3(n9827), .A4(n9826), .ZN(P1_U3244) );
  NAND2_X1 U12324 ( .A1(n9834), .A2(P2_U3088), .ZN(n13650) );
  NAND2_X1 U12325 ( .A1(n6439), .A2(P2_U3088), .ZN(n13651) );
  OAI222_X1 U12326 ( .A1(n13650), .A2(n9830), .B1(n13651), .B2(n9832), .C1(
        P2_U3088), .C2(n9938), .ZN(P2_U3326) );
  NAND2_X2 U12327 ( .A1(n6439), .A2(P1_U3086), .ZN(n14201) );
  OAI222_X1 U12328 ( .A1(n10005), .A2(P1_U3086), .B1(n14204), .B2(n9832), .C1(
        n7580), .C2(n14201), .ZN(P1_U3354) );
  NAND2_X1 U12329 ( .A1(n9834), .A2(P3_U3151), .ZN(n12960) );
  INV_X1 U12330 ( .A(n14320), .ZN(n12396) );
  INV_X1 U12331 ( .A(n9835), .ZN(n9837) );
  INV_X2 U12332 ( .A(n14319), .ZN(n12962) );
  OAI222_X1 U12333 ( .A1(n12396), .A2(n9837), .B1(n12962), .B2(n9836), .C1(
        P3_U3151), .C2(n10422), .ZN(P3_U3294) );
  INV_X1 U12334 ( .A(n9838), .ZN(n9840) );
  OAI222_X1 U12335 ( .A1(P3_U3151), .A2(n10548), .B1(n12960), .B2(n9840), .C1(
        n9839), .C2(n12962), .ZN(P3_U3289) );
  INV_X1 U12336 ( .A(n14889), .ZN(n10464) );
  INV_X1 U12337 ( .A(SI_3_), .ZN(n9841) );
  OAI222_X1 U12338 ( .A1(n10464), .A2(P3_U3151), .B1(n12960), .B2(n9842), .C1(
        n9841), .C2(n12962), .ZN(P3_U3292) );
  INV_X1 U12339 ( .A(n12569), .ZN(n10459) );
  INV_X1 U12340 ( .A(SI_2_), .ZN(n9843) );
  OAI222_X1 U12341 ( .A1(n10459), .A2(P3_U3151), .B1(n12960), .B2(n9844), .C1(
        n9843), .C2(n12962), .ZN(P3_U3293) );
  INV_X1 U12342 ( .A(SI_7_), .ZN(n9845) );
  OAI222_X1 U12343 ( .A1(n10571), .A2(P3_U3151), .B1(n12396), .B2(n9846), .C1(
        n9845), .C2(n12962), .ZN(P3_U3288) );
  INV_X1 U12344 ( .A(n10343), .ZN(n10006) );
  INV_X1 U12345 ( .A(n9847), .ZN(n9865) );
  OAI222_X1 U12346 ( .A1(n10006), .A2(P1_U3086), .B1(n14204), .B2(n9865), .C1(
        n9848), .C2(n14201), .ZN(P1_U3353) );
  INV_X1 U12347 ( .A(n14907), .ZN(n10446) );
  INV_X1 U12348 ( .A(SI_4_), .ZN(n9850) );
  OAI222_X1 U12349 ( .A1(P3_U3151), .A2(n10446), .B1(n12962), .B2(n9850), .C1(
        n12396), .C2(n9849), .ZN(P3_U3291) );
  OAI222_X1 U12350 ( .A1(P3_U3151), .A2(n14922), .B1(n12962), .B2(n7079), .C1(
        n12396), .C2(n9851), .ZN(P3_U3290) );
  INV_X1 U12351 ( .A(n9852), .ZN(n9853) );
  OAI222_X1 U12352 ( .A1(P3_U3151), .A2(n12635), .B1(n12962), .B2(n9854), .C1(
        n12396), .C2(n9853), .ZN(P3_U3287) );
  INV_X1 U12353 ( .A(n9855), .ZN(n9867) );
  OAI222_X1 U12354 ( .A1(n13814), .A2(P1_U3086), .B1(n14204), .B2(n9867), .C1(
        n9856), .C2(n14201), .ZN(P1_U3352) );
  INV_X1 U12355 ( .A(n13832), .ZN(n13826) );
  INV_X1 U12356 ( .A(n9857), .ZN(n9869) );
  OAI222_X1 U12357 ( .A1(n13826), .A2(P1_U3086), .B1(n14204), .B2(n9869), .C1(
        n9858), .C2(n14201), .ZN(P1_U3351) );
  INV_X1 U12358 ( .A(SI_9_), .ZN(n9859) );
  OAI222_X1 U12359 ( .A1(n14940), .A2(P3_U3151), .B1(n12396), .B2(n9860), .C1(
        n9859), .C2(n12962), .ZN(P3_U3286) );
  INV_X1 U12360 ( .A(n10055), .ZN(n10029) );
  INV_X1 U12361 ( .A(n9861), .ZN(n9871) );
  OAI222_X1 U12362 ( .A1(n10029), .A2(P1_U3086), .B1(n14204), .B2(n9871), .C1(
        n9862), .C2(n14201), .ZN(P1_U3350) );
  INV_X1 U12363 ( .A(SI_10_), .ZN(n9864) );
  OAI222_X1 U12364 ( .A1(P3_U3151), .A2(n14963), .B1(n12962), .B2(n9864), .C1(
        n12396), .C2(n9863), .ZN(P3_U3285) );
  INV_X1 U12365 ( .A(n13650), .ZN(n11743) );
  INV_X1 U12366 ( .A(n11743), .ZN(n13624) );
  INV_X1 U12367 ( .A(n13651), .ZN(n13635) );
  INV_X1 U12368 ( .A(n13635), .ZN(n13645) );
  OAI222_X1 U12369 ( .A1(n13624), .A2(n9866), .B1(n13645), .B2(n9865), .C1(
        P2_U3088), .C2(n13152), .ZN(P2_U3325) );
  OAI222_X1 U12370 ( .A1(n13624), .A2(n9868), .B1(n13645), .B2(n9867), .C1(
        P2_U3088), .C2(n13166), .ZN(P2_U3324) );
  OAI222_X1 U12371 ( .A1(n13624), .A2(n9870), .B1(n13645), .B2(n9869), .C1(
        P2_U3088), .C2(n13181), .ZN(P2_U3323) );
  OAI222_X1 U12372 ( .A1(n13624), .A2(n9872), .B1(n13645), .B2(n9871), .C1(
        P2_U3088), .C2(n10081), .ZN(P2_U3322) );
  INV_X1 U12373 ( .A(n10188), .ZN(n10048) );
  INV_X1 U12374 ( .A(n9873), .ZN(n9875) );
  OAI222_X1 U12375 ( .A1(n10048), .A2(P1_U3086), .B1(n14204), .B2(n9875), .C1(
        n9874), .C2(n14201), .ZN(P1_U3349) );
  OAI222_X1 U12376 ( .A1(n13624), .A2(n9876), .B1(n13645), .B2(n9875), .C1(
        P2_U3088), .C2(n13196), .ZN(P2_U3321) );
  INV_X1 U12377 ( .A(n9877), .ZN(n9879) );
  OAI222_X1 U12378 ( .A1(n13624), .A2(n9878), .B1(n13645), .B2(n9879), .C1(
        P2_U3088), .C2(n13210), .ZN(P2_U3320) );
  INV_X1 U12379 ( .A(n10159), .ZN(n10167) );
  OAI222_X1 U12380 ( .A1(n10167), .A2(P1_U3086), .B1(n14204), .B2(n9879), .C1(
        n7240), .C2(n14201), .ZN(P1_U3348) );
  INV_X1 U12381 ( .A(n9880), .ZN(n9883) );
  OAI222_X1 U12382 ( .A1(n13624), .A2(n9881), .B1(n13645), .B2(n9883), .C1(
        P2_U3088), .C2(n13227), .ZN(P2_U3319) );
  INV_X1 U12383 ( .A(n10102), .ZN(n10106) );
  OAI222_X1 U12384 ( .A1(n10106), .A2(P1_U3086), .B1(n14204), .B2(n9883), .C1(
        n9882), .C2(n14201), .ZN(P1_U3347) );
  INV_X1 U12385 ( .A(n9884), .ZN(n9886) );
  OAI222_X1 U12386 ( .A1(n13624), .A2(n15276), .B1(n13645), .B2(n9886), .C1(
        P2_U3088), .C2(n14768), .ZN(P2_U3318) );
  INV_X1 U12387 ( .A(n10209), .ZN(n10114) );
  INV_X1 U12388 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9885) );
  OAI222_X1 U12389 ( .A1(n10114), .A2(P1_U3086), .B1(n14204), .B2(n9886), .C1(
        n9885), .C2(n14201), .ZN(P1_U3346) );
  INV_X1 U12390 ( .A(n12941), .ZN(n9889) );
  INV_X1 U12391 ( .A(n9887), .ZN(n10720) );
  NAND2_X1 U12392 ( .A1(n9889), .A2(n10720), .ZN(n9888) );
  OAI21_X1 U12393 ( .B1(n9889), .B2(n9423), .A(n9888), .ZN(P3_U3377) );
  NAND2_X1 U12394 ( .A1(n9890), .A2(n11742), .ZN(n9891) );
  NAND2_X1 U12395 ( .A1(n9892), .A2(n9891), .ZN(n9893) );
  NAND2_X1 U12396 ( .A1(n9894), .A2(n9893), .ZN(n9908) );
  INV_X1 U12397 ( .A(n8179), .ZN(n9899) );
  NAND2_X1 U12398 ( .A1(n9899), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13636) );
  INV_X1 U12399 ( .A(n13636), .ZN(n9895) );
  NAND2_X1 U12400 ( .A1(n9908), .A2(n9895), .ZN(n9901) );
  INV_X1 U12401 ( .A(n13640), .ZN(n12145) );
  INV_X1 U12402 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9896) );
  NOR2_X1 U12403 ( .A1(n14750), .A2(n9896), .ZN(n14749) );
  INV_X1 U12404 ( .A(n14750), .ZN(n14814) );
  MUX2_X1 U12405 ( .A(n9937), .B(P2_REG1_REG_1__SCAN_IN), .S(n9938), .Z(n9898)
         );
  AOI22_X1 U12406 ( .A1(n14749), .A2(P2_IR_REG_0__SCAN_IN), .B1(n14814), .B2(
        n9898), .ZN(n9916) );
  AND2_X1 U12407 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9897) );
  NAND2_X1 U12408 ( .A1(n9898), .A2(n9897), .ZN(n13149) );
  INV_X1 U12409 ( .A(n13149), .ZN(n9915) );
  NOR2_X1 U12410 ( .A1(n9899), .A2(P2_U3088), .ZN(n9900) );
  INV_X1 U12411 ( .A(n9901), .ZN(n9902) );
  INV_X1 U12412 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10664) );
  MUX2_X1 U12413 ( .A(n10664), .B(P2_REG2_REG_1__SCAN_IN), .S(n9938), .Z(n9903) );
  AND2_X1 U12414 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9904) );
  NAND2_X1 U12415 ( .A1(n9903), .A2(n9904), .ZN(n13154) );
  MUX2_X1 U12416 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10664), .S(n9938), .Z(n9906) );
  INV_X1 U12417 ( .A(n9904), .ZN(n9905) );
  NAND2_X1 U12418 ( .A1(n9906), .A2(n9905), .ZN(n9907) );
  NAND3_X1 U12419 ( .A1(n14820), .A2(n13154), .A3(n9907), .ZN(n9912) );
  INV_X1 U12420 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9909) );
  OAI22_X1 U12421 ( .A1(n14791), .A2(n9909), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10666), .ZN(n9910) );
  INV_X1 U12422 ( .A(n9910), .ZN(n9911) );
  OAI211_X1 U12423 ( .C1(n14769), .C2(n9938), .A(n9912), .B(n9911), .ZN(n9913)
         );
  INV_X1 U12424 ( .A(n9913), .ZN(n9914) );
  OAI21_X1 U12425 ( .B1(n9916), .B2(n9915), .A(n9914), .ZN(P2_U3215) );
  INV_X1 U12426 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n12416) );
  NAND2_X1 U12427 ( .A1(n9917), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9920) );
  NAND2_X1 U12428 ( .A1(n9918), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9919) );
  OAI211_X1 U12429 ( .C1(n9921), .C2(n12416), .A(n9920), .B(n9919), .ZN(n12412) );
  NAND2_X1 U12430 ( .A1(P2_U3947), .A2(n12412), .ZN(n9922) );
  OAI21_X1 U12431 ( .B1(P2_U3947), .B2(n9923), .A(n9922), .ZN(P2_U3562) );
  INV_X1 U12432 ( .A(n9924), .ZN(n9927) );
  OAI222_X1 U12433 ( .A1(n13624), .A2(n9925), .B1(n13645), .B2(n9927), .C1(
        P2_U3088), .C2(n10123), .ZN(P2_U3317) );
  INV_X1 U12434 ( .A(n10295), .ZN(n10217) );
  OAI222_X1 U12435 ( .A1(n10217), .A2(P1_U3086), .B1(n14204), .B2(n9927), .C1(
        n9926), .C2(n14201), .ZN(P1_U3345) );
  MUX2_X1 U12436 ( .A(n7737), .B(P2_REG2_REG_2__SCAN_IN), .S(n13152), .Z(n9929) );
  OR2_X1 U12437 ( .A1(n9938), .A2(n10664), .ZN(n13153) );
  NAND2_X1 U12438 ( .A1(n13154), .A2(n13153), .ZN(n9928) );
  NAND2_X1 U12439 ( .A1(n9929), .A2(n9928), .ZN(n13169) );
  INV_X1 U12440 ( .A(n13152), .ZN(n13147) );
  NAND2_X1 U12441 ( .A1(n13147), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n13167) );
  NAND2_X1 U12442 ( .A1(n13169), .A2(n13167), .ZN(n9931) );
  INV_X1 U12443 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10642) );
  MUX2_X1 U12444 ( .A(n10642), .B(P2_REG2_REG_3__SCAN_IN), .S(n13166), .Z(
        n9930) );
  NAND2_X1 U12445 ( .A1(n9931), .A2(n9930), .ZN(n13184) );
  OR2_X1 U12446 ( .A1(n13166), .A2(n10642), .ZN(n13183) );
  NAND2_X1 U12447 ( .A1(n13184), .A2(n13183), .ZN(n9933) );
  INV_X1 U12448 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10774) );
  MUX2_X1 U12449 ( .A(n10774), .B(P2_REG2_REG_4__SCAN_IN), .S(n13181), .Z(
        n9932) );
  NAND2_X1 U12450 ( .A1(n9933), .A2(n9932), .ZN(n13186) );
  OR2_X1 U12451 ( .A1(n13181), .A2(n10774), .ZN(n9934) );
  NAND2_X1 U12452 ( .A1(n13186), .A2(n9934), .ZN(n9936) );
  MUX2_X1 U12453 ( .A(n10704), .B(P2_REG2_REG_5__SCAN_IN), .S(n10081), .Z(
        n9935) );
  NAND2_X1 U12454 ( .A1(n9936), .A2(n9935), .ZN(n13199) );
  OAI211_X1 U12455 ( .C1(n9936), .C2(n9935), .A(n14820), .B(n13199), .ZN(n9953) );
  INV_X1 U12456 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9937) );
  OR2_X1 U12457 ( .A1(n9938), .A2(n9937), .ZN(n13148) );
  NAND2_X1 U12458 ( .A1(n13149), .A2(n13148), .ZN(n9941) );
  MUX2_X1 U12459 ( .A(n9939), .B(P2_REG1_REG_2__SCAN_IN), .S(n13152), .Z(n9940) );
  NAND2_X1 U12460 ( .A1(n9941), .A2(n9940), .ZN(n13164) );
  NAND2_X1 U12461 ( .A1(n13147), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n13163) );
  NAND2_X1 U12462 ( .A1(n13164), .A2(n13163), .ZN(n9944) );
  MUX2_X1 U12463 ( .A(n9942), .B(P2_REG1_REG_3__SCAN_IN), .S(n13166), .Z(n9943) );
  NAND2_X1 U12464 ( .A1(n9944), .A2(n9943), .ZN(n13178) );
  OR2_X1 U12465 ( .A1(n13166), .A2(n9942), .ZN(n13177) );
  NAND2_X1 U12466 ( .A1(n13178), .A2(n13177), .ZN(n9947) );
  MUX2_X1 U12467 ( .A(n9945), .B(P2_REG1_REG_4__SCAN_IN), .S(n13181), .Z(n9946) );
  NAND2_X1 U12468 ( .A1(n9947), .A2(n9946), .ZN(n13180) );
  OR2_X1 U12469 ( .A1(n13181), .A2(n9945), .ZN(n9948) );
  NAND2_X1 U12470 ( .A1(n13180), .A2(n9948), .ZN(n9951) );
  MUX2_X1 U12471 ( .A(n9949), .B(P2_REG1_REG_5__SCAN_IN), .S(n10081), .Z(n9950) );
  NAND2_X1 U12472 ( .A1(n9951), .A2(n9950), .ZN(n13194) );
  OAI211_X1 U12473 ( .C1(n9951), .C2(n9950), .A(n14814), .B(n13194), .ZN(n9952) );
  NAND2_X1 U12474 ( .A1(n9953), .A2(n9952), .ZN(n9954) );
  AND2_X1 U12475 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10625) );
  AOI211_X1 U12476 ( .C1(n14812), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n9954), .B(
        n10625), .ZN(n9955) );
  OAI21_X1 U12477 ( .B1(n10081), .B2(n14769), .A(n9955), .ZN(P2_U3219) );
  OAI222_X1 U12478 ( .A1(P3_U3151), .A2(n15012), .B1(n12962), .B2(n9957), .C1(
        n12396), .C2(n9956), .ZN(P3_U3282) );
  INV_X1 U12479 ( .A(n9958), .ZN(n9960) );
  OAI222_X1 U12480 ( .A1(n13624), .A2(n15289), .B1(n13645), .B2(n9960), .C1(
        P2_U3088), .C2(n10311), .ZN(P2_U3316) );
  INV_X1 U12481 ( .A(n10790), .ZN(n10300) );
  OAI222_X1 U12482 ( .A1(n10300), .A2(P1_U3086), .B1(n14204), .B2(n9960), .C1(
        n9959), .C2(n14201), .ZN(P1_U3344) );
  NAND2_X1 U12483 ( .A1(n12981), .A2(P2_U3947), .ZN(n9961) );
  OAI21_X1 U12484 ( .B1(n7649), .B2(P2_U3947), .A(n9961), .ZN(P2_U3549) );
  INV_X1 U12485 ( .A(n9962), .ZN(n9968) );
  OAI222_X1 U12486 ( .A1(n13651), .A2(n9968), .B1(n14779), .B2(P2_U3088), .C1(
        n9963), .C2(n13624), .ZN(P2_U3315) );
  INV_X1 U12487 ( .A(n9964), .ZN(n9965) );
  OAI222_X1 U12488 ( .A1(P3_U3151), .A2(n15032), .B1(n12962), .B2(n9966), .C1(
        n12396), .C2(n9965), .ZN(P3_U3281) );
  INV_X1 U12489 ( .A(n10795), .ZN(n14600) );
  OAI222_X1 U12490 ( .A1(P1_U3086), .A2(n14600), .B1(n14204), .B2(n9968), .C1(
        n9967), .C2(n14201), .ZN(P1_U3343) );
  INV_X1 U12491 ( .A(n9969), .ZN(n10037) );
  INV_X1 U12492 ( .A(n14201), .ZN(n14188) );
  AOI22_X1 U12493 ( .A1(n11269), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n14188), .ZN(n9970) );
  OAI21_X1 U12494 ( .B1(n10037), .B2(n14204), .A(n9970), .ZN(P1_U3342) );
  INV_X1 U12495 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n15216) );
  NAND2_X1 U12496 ( .A1(n9971), .A2(P3_U3897), .ZN(n9972) );
  OAI21_X1 U12497 ( .B1(P3_U3897), .B2(n15216), .A(n9972), .ZN(P3_U3505) );
  NOR2_X1 U12498 ( .A1(n12941), .A2(n9973), .ZN(n9975) );
  INV_X1 U12499 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9974) );
  NOR2_X1 U12500 ( .A1(n10001), .A2(n9974), .ZN(P3_U3262) );
  INV_X1 U12501 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9976) );
  NOR2_X1 U12502 ( .A1(n10001), .A2(n9976), .ZN(P3_U3263) );
  INV_X1 U12503 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9977) );
  NOR2_X1 U12504 ( .A1(n10001), .A2(n9977), .ZN(P3_U3257) );
  INV_X1 U12505 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n15219) );
  NOR2_X1 U12506 ( .A1(n10001), .A2(n15219), .ZN(P3_U3256) );
  INV_X1 U12507 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9978) );
  NOR2_X1 U12508 ( .A1(n10001), .A2(n9978), .ZN(P3_U3255) );
  INV_X1 U12509 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9979) );
  NOR2_X1 U12510 ( .A1(n10001), .A2(n9979), .ZN(P3_U3254) );
  INV_X1 U12511 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9980) );
  NOR2_X1 U12512 ( .A1(n10001), .A2(n9980), .ZN(P3_U3261) );
  INV_X1 U12513 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n9981) );
  NOR2_X1 U12514 ( .A1(n9975), .A2(n9981), .ZN(P3_U3260) );
  INV_X1 U12515 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9982) );
  NOR2_X1 U12516 ( .A1(n10001), .A2(n9982), .ZN(P3_U3259) );
  INV_X1 U12517 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9983) );
  NOR2_X1 U12518 ( .A1(n9975), .A2(n9983), .ZN(P3_U3258) );
  INV_X1 U12519 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9984) );
  NOR2_X1 U12520 ( .A1(n10001), .A2(n9984), .ZN(P3_U3251) );
  INV_X1 U12521 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9985) );
  NOR2_X1 U12522 ( .A1(n10001), .A2(n9985), .ZN(P3_U3249) );
  INV_X1 U12523 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9986) );
  NOR2_X1 U12524 ( .A1(n10001), .A2(n9986), .ZN(P3_U3248) );
  INV_X1 U12525 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9987) );
  NOR2_X1 U12526 ( .A1(n10001), .A2(n9987), .ZN(P3_U3247) );
  INV_X1 U12527 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9988) );
  NOR2_X1 U12528 ( .A1(n10001), .A2(n9988), .ZN(P3_U3253) );
  INV_X1 U12529 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9989) );
  NOR2_X1 U12530 ( .A1(n10001), .A2(n9989), .ZN(P3_U3252) );
  INV_X1 U12531 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9990) );
  NOR2_X1 U12532 ( .A1(n10001), .A2(n9990), .ZN(P3_U3246) );
  INV_X1 U12533 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9991) );
  NOR2_X1 U12534 ( .A1(n9975), .A2(n9991), .ZN(P3_U3245) );
  INV_X1 U12535 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9992) );
  NOR2_X1 U12536 ( .A1(n9975), .A2(n9992), .ZN(P3_U3244) );
  INV_X1 U12537 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9993) );
  NOR2_X1 U12538 ( .A1(n9975), .A2(n9993), .ZN(P3_U3243) );
  INV_X1 U12539 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9994) );
  NOR2_X1 U12540 ( .A1(n9975), .A2(n9994), .ZN(P3_U3242) );
  INV_X1 U12541 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n9995) );
  NOR2_X1 U12542 ( .A1(n9975), .A2(n9995), .ZN(P3_U3241) );
  INV_X1 U12543 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9996) );
  NOR2_X1 U12544 ( .A1(n9975), .A2(n9996), .ZN(P3_U3240) );
  INV_X1 U12545 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9997) );
  NOR2_X1 U12546 ( .A1(n9975), .A2(n9997), .ZN(P3_U3239) );
  INV_X1 U12547 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9998) );
  NOR2_X1 U12548 ( .A1(n9975), .A2(n9998), .ZN(P3_U3238) );
  INV_X1 U12549 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9999) );
  NOR2_X1 U12550 ( .A1(n9975), .A2(n9999), .ZN(P3_U3237) );
  INV_X1 U12551 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10000) );
  NOR2_X1 U12552 ( .A1(n10001), .A2(n10000), .ZN(P3_U3250) );
  INV_X1 U12553 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10002) );
  NOR2_X1 U12554 ( .A1(n10001), .A2(n10002), .ZN(P3_U3236) );
  INV_X1 U12555 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10003) );
  NOR2_X1 U12556 ( .A1(n10001), .A2(n10003), .ZN(P3_U3235) );
  INV_X1 U12557 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n15181) );
  NOR2_X1 U12558 ( .A1(n10001), .A2(n15181), .ZN(P3_U3234) );
  XOR2_X1 U12559 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10055), .Z(n10011) );
  INV_X1 U12560 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10008) );
  INV_X1 U12561 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10007) );
  OAI21_X1 U12562 ( .B1(n10005), .B2(n15162), .A(n10004), .ZN(n10337) );
  MUX2_X1 U12563 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10007), .S(n10343), .Z(
        n10338) );
  NAND2_X1 U12564 ( .A1(n10337), .A2(n10338), .ZN(n10336) );
  OAI21_X1 U12565 ( .B1(n10007), .B2(n10006), .A(n10336), .ZN(n13818) );
  MUX2_X1 U12566 ( .A(n10008), .B(P1_REG1_REG_3__SCAN_IN), .S(n13814), .Z(
        n13819) );
  NAND2_X1 U12567 ( .A1(n13818), .A2(n13819), .ZN(n13817) );
  INV_X1 U12568 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n15244) );
  MUX2_X1 U12569 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n15244), .S(n13832), .Z(
        n13831) );
  INV_X1 U12570 ( .A(n13829), .ZN(n10009) );
  NAND2_X1 U12571 ( .A1(n10010), .A2(n10011), .ZN(n10054) );
  OAI21_X1 U12572 ( .B1(n10011), .B2(n10010), .A(n10054), .ZN(n10025) );
  MUX2_X1 U12573 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10012), .S(n10343), .Z(
        n10335) );
  NAND2_X1 U12574 ( .A1(n10013), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10014) );
  NAND2_X1 U12575 ( .A1(n10015), .A2(n10014), .ZN(n10334) );
  AOI22_X1 U12576 ( .A1(n10335), .A2(n10334), .B1(n10343), .B2(
        P1_REG2_REG_2__SCAN_IN), .ZN(n13821) );
  INV_X1 U12577 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10016) );
  MUX2_X1 U12578 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10016), .S(n13814), .Z(
        n13820) );
  NOR2_X1 U12579 ( .A1(n13821), .A2(n13820), .ZN(n13838) );
  NOR2_X1 U12580 ( .A1(n13814), .A2(n10016), .ZN(n13833) );
  INV_X1 U12581 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10017) );
  MUX2_X1 U12582 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10017), .S(n13832), .Z(
        n10018) );
  OAI21_X1 U12583 ( .B1(n13838), .B2(n13833), .A(n10018), .ZN(n13836) );
  INV_X1 U12584 ( .A(n13836), .ZN(n10021) );
  NOR2_X1 U12585 ( .A1(n13826), .A2(n10017), .ZN(n10020) );
  MUX2_X1 U12586 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10869), .S(n10055), .Z(
        n10019) );
  OAI21_X1 U12587 ( .B1(n10021), .B2(n10020), .A(n10019), .ZN(n10185) );
  INV_X1 U12588 ( .A(n10185), .ZN(n10023) );
  NOR3_X1 U12589 ( .A1(n10021), .A2(n10020), .A3(n10019), .ZN(n10022) );
  NOR3_X1 U12590 ( .A1(n14596), .A2(n10023), .A3(n10022), .ZN(n10024) );
  AOI21_X1 U12591 ( .B1(n14591), .B2(n10025), .A(n10024), .ZN(n10028) );
  INV_X1 U12592 ( .A(n14605), .ZN(n13852) );
  AND2_X1 U12593 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10026) );
  AOI21_X1 U12594 ( .B1(n13852), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10026), .ZN(
        n10027) );
  OAI211_X1 U12595 ( .C1(n10029), .C2(n14601), .A(n10028), .B(n10027), .ZN(
        P1_U3248) );
  AOI21_X1 U12596 ( .B1(n9789), .B2(n10030), .A(n13081), .ZN(n10035) );
  OR2_X1 U12597 ( .A1(n10031), .A2(P2_U3088), .ZN(n10177) );
  NAND2_X1 U12598 ( .A1(n11872), .A2(n13061), .ZN(n10142) );
  NAND4_X1 U12599 ( .A1(n10140), .A2(n13143), .A3(n9789), .A4(n13460), .ZN(
        n10032) );
  OAI21_X1 U12600 ( .B1(n13108), .B2(n10142), .A(n10032), .ZN(n10033) );
  AOI21_X1 U12601 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n10177), .A(n10033), .ZN(
        n10034) );
  OAI21_X1 U12602 ( .B1(n10035), .B2(n11865), .A(n10034), .ZN(P2_U3204) );
  INV_X1 U12603 ( .A(n10312), .ZN(n11309) );
  OAI222_X1 U12604 ( .A1(n13651), .A2(n10037), .B1(n11309), .B2(P2_U3088), 
        .C1(n10036), .C2(n13650), .ZN(P2_U3314) );
  INV_X1 U12605 ( .A(n10038), .ZN(n10039) );
  OAI222_X1 U12606 ( .A1(P3_U3151), .A2(n14376), .B1(n12962), .B2(n10040), 
        .C1(n12396), .C2(n10039), .ZN(P3_U3280) );
  AOI21_X1 U12607 ( .B1(n10042), .B2(n10041), .A(n6608), .ZN(n10046) );
  INV_X1 U12608 ( .A(n10177), .ZN(n10043) );
  AOI22_X1 U12609 ( .A1(n13050), .A2(n13143), .B1(n13142), .B2(n13061), .ZN(
        n10200) );
  OAI22_X1 U12610 ( .A1(n10043), .A2(n10666), .B1(n13108), .B2(n10200), .ZN(
        n10044) );
  AOI21_X1 U12611 ( .B1(n11869), .B2(n13081), .A(n10044), .ZN(n10045) );
  OAI21_X1 U12612 ( .B1(n10046), .B2(n13070), .A(n10045), .ZN(P2_U3194) );
  NAND2_X1 U12613 ( .A1(n10055), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10184) );
  INV_X1 U12614 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10047) );
  MUX2_X1 U12615 ( .A(n10047), .B(P1_REG2_REG_6__SCAN_IN), .S(n10188), .Z(
        n10183) );
  AOI21_X1 U12616 ( .B1(n10185), .B2(n10184), .A(n10183), .ZN(n10187) );
  NOR2_X1 U12617 ( .A1(n10048), .A2(n10047), .ZN(n10158) );
  INV_X1 U12618 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10049) );
  MUX2_X1 U12619 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10049), .S(n10159), .Z(
        n10050) );
  OAI21_X1 U12620 ( .B1(n10187), .B2(n10158), .A(n10050), .ZN(n10162) );
  NAND2_X1 U12621 ( .A1(n10159), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10052) );
  INV_X1 U12622 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10105) );
  MUX2_X1 U12623 ( .A(n10105), .B(P1_REG2_REG_8__SCAN_IN), .S(n10102), .Z(
        n10051) );
  AOI21_X1 U12624 ( .B1(n10162), .B2(n10052), .A(n10051), .ZN(n10110) );
  NAND3_X1 U12625 ( .A1(n10162), .A2(n10052), .A3(n10051), .ZN(n10053) );
  NAND2_X1 U12626 ( .A1(n13887), .A2(n10053), .ZN(n10066) );
  INV_X1 U12627 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10056) );
  MUX2_X1 U12628 ( .A(n10056), .B(P1_REG1_REG_6__SCAN_IN), .S(n10188), .Z(
        n10182) );
  NOR2_X1 U12629 ( .A1(n10181), .A2(n10182), .ZN(n10180) );
  INV_X1 U12630 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10057) );
  MUX2_X1 U12631 ( .A(n10057), .B(P1_REG1_REG_7__SCAN_IN), .S(n10159), .Z(
        n10156) );
  NOR2_X1 U12632 ( .A1(n10157), .A2(n10156), .ZN(n10155) );
  INV_X1 U12633 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10058) );
  MUX2_X1 U12634 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10058), .S(n10102), .Z(
        n10059) );
  NAND2_X1 U12635 ( .A1(n10060), .A2(n10059), .ZN(n10101) );
  OAI21_X1 U12636 ( .B1(n10060), .B2(n10059), .A(n10101), .ZN(n10061) );
  NAND2_X1 U12637 ( .A1(n10061), .A2(n14591), .ZN(n10065) );
  NAND2_X1 U12638 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11414) );
  INV_X1 U12639 ( .A(n11414), .ZN(n10063) );
  NOR2_X1 U12640 ( .A1(n14601), .A2(n10106), .ZN(n10062) );
  AOI211_X1 U12641 ( .C1(n13852), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10063), .B(
        n10062), .ZN(n10064) );
  OAI211_X1 U12642 ( .C1(n10110), .C2(n10066), .A(n10065), .B(n10064), .ZN(
        P1_U3251) );
  MUX2_X1 U12643 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7884), .S(n10123), .Z(
        n10078) );
  OR2_X1 U12644 ( .A1(n10081), .A2(n9949), .ZN(n13193) );
  NAND2_X1 U12645 ( .A1(n13194), .A2(n13193), .ZN(n10069) );
  MUX2_X1 U12646 ( .A(n10067), .B(P2_REG1_REG_6__SCAN_IN), .S(n13196), .Z(
        n10068) );
  NAND2_X1 U12647 ( .A1(n10069), .A2(n10068), .ZN(n13208) );
  OR2_X1 U12648 ( .A1(n13196), .A2(n10067), .ZN(n13207) );
  NAND2_X1 U12649 ( .A1(n13208), .A2(n13207), .ZN(n10072) );
  MUX2_X1 U12650 ( .A(n10070), .B(P2_REG1_REG_7__SCAN_IN), .S(n13210), .Z(
        n10071) );
  NAND2_X1 U12651 ( .A1(n10072), .A2(n10071), .ZN(n13224) );
  OR2_X1 U12652 ( .A1(n13210), .A2(n10070), .ZN(n13223) );
  NAND2_X1 U12653 ( .A1(n13224), .A2(n13223), .ZN(n10074) );
  MUX2_X1 U12654 ( .A(n13221), .B(P2_REG1_REG_8__SCAN_IN), .S(n13227), .Z(
        n10073) );
  NAND2_X1 U12655 ( .A1(n10074), .A2(n10073), .ZN(n13226) );
  INV_X1 U12656 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n13221) );
  OR2_X1 U12657 ( .A1(n13227), .A2(n13221), .ZN(n10075) );
  NAND2_X1 U12658 ( .A1(n13226), .A2(n10075), .ZN(n14757) );
  MUX2_X1 U12659 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10076), .S(n14768), .Z(
        n14756) );
  OR2_X1 U12660 ( .A1(n14757), .A2(n14756), .ZN(n14759) );
  NAND2_X1 U12661 ( .A1(n14768), .A2(n10076), .ZN(n10077) );
  NAND2_X1 U12662 ( .A1(n14759), .A2(n10077), .ZN(n10079) );
  AOI21_X1 U12663 ( .B1(n10078), .B2(n10079), .A(n14750), .ZN(n10080) );
  NAND2_X1 U12664 ( .A1(n10080), .A2(n10129), .ZN(n10095) );
  MUX2_X1 U12665 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n11281), .S(n10123), .Z(
        n10092) );
  INV_X1 U12666 ( .A(n14768), .ZN(n10090) );
  OR2_X1 U12667 ( .A1(n10081), .A2(n10704), .ZN(n13198) );
  NAND2_X1 U12668 ( .A1(n13199), .A2(n13198), .ZN(n10083) );
  INV_X1 U12669 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11035) );
  MUX2_X1 U12670 ( .A(n11035), .B(P2_REG2_REG_6__SCAN_IN), .S(n13196), .Z(
        n10082) );
  NAND2_X1 U12671 ( .A1(n10083), .A2(n10082), .ZN(n13213) );
  OR2_X1 U12672 ( .A1(n13196), .A2(n11035), .ZN(n13212) );
  NAND2_X1 U12673 ( .A1(n13213), .A2(n13212), .ZN(n10086) );
  INV_X1 U12674 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10084) );
  MUX2_X1 U12675 ( .A(n10084), .B(P2_REG2_REG_7__SCAN_IN), .S(n13210), .Z(
        n10085) );
  NAND2_X1 U12676 ( .A1(n10086), .A2(n10085), .ZN(n13230) );
  OR2_X1 U12677 ( .A1(n13210), .A2(n10084), .ZN(n13229) );
  NAND2_X1 U12678 ( .A1(n13230), .A2(n13229), .ZN(n10088) );
  INV_X1 U12679 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10991) );
  MUX2_X1 U12680 ( .A(n10991), .B(P2_REG2_REG_8__SCAN_IN), .S(n13227), .Z(
        n10087) );
  NAND2_X1 U12681 ( .A1(n10088), .A2(n10087), .ZN(n13232) );
  OR2_X1 U12682 ( .A1(n13227), .A2(n10991), .ZN(n10089) );
  NAND2_X1 U12683 ( .A1(n13232), .A2(n10089), .ZN(n14762) );
  MUX2_X1 U12684 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n13474), .S(n14768), .Z(
        n14761) );
  OAI21_X1 U12685 ( .B1(n10090), .B2(P2_REG2_REG_9__SCAN_IN), .A(n14764), .ZN(
        n10091) );
  NOR2_X1 U12686 ( .A1(n10091), .A2(n10092), .ZN(n10119) );
  INV_X1 U12687 ( .A(n14820), .ZN(n14751) );
  AOI211_X1 U12688 ( .C1(n10092), .C2(n10091), .A(n10119), .B(n14751), .ZN(
        n10093) );
  INV_X1 U12689 ( .A(n10093), .ZN(n10094) );
  NAND2_X1 U12690 ( .A1(n10095), .A2(n10094), .ZN(n10097) );
  NAND2_X1 U12691 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11295)
         );
  INV_X1 U12692 ( .A(n11295), .ZN(n10096) );
  AOI211_X1 U12693 ( .C1(n14812), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n10097), 
        .B(n10096), .ZN(n10098) );
  OAI21_X1 U12694 ( .B1(n10123), .B2(n14769), .A(n10098), .ZN(P2_U3224) );
  INV_X1 U12695 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10099) );
  MUX2_X1 U12696 ( .A(n10099), .B(P1_REG1_REG_9__SCAN_IN), .S(n10209), .Z(
        n10100) );
  INV_X1 U12697 ( .A(n10100), .ZN(n10104) );
  OAI21_X1 U12698 ( .B1(n10102), .B2(P1_REG1_REG_8__SCAN_IN), .A(n10101), .ZN(
        n10103) );
  NAND2_X1 U12699 ( .A1(n10103), .A2(n10104), .ZN(n10206) );
  OAI21_X1 U12700 ( .B1(n10104), .B2(n10103), .A(n10206), .ZN(n10117) );
  NOR2_X1 U12701 ( .A1(n10106), .A2(n10105), .ZN(n10109) );
  MUX2_X1 U12702 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10107), .S(n10209), .Z(
        n10108) );
  OAI21_X1 U12703 ( .B1(n10110), .B2(n10109), .A(n10108), .ZN(n10212) );
  INV_X1 U12704 ( .A(n10212), .ZN(n10112) );
  NOR3_X1 U12705 ( .A1(n10110), .A2(n10109), .A3(n10108), .ZN(n10111) );
  NOR3_X1 U12706 ( .A1(n10112), .A2(n10111), .A3(n14596), .ZN(n10116) );
  NOR2_X1 U12707 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8466), .ZN(n11556) );
  AOI21_X1 U12708 ( .B1(n13852), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n11556), .ZN(
        n10113) );
  OAI21_X1 U12709 ( .B1(n10114), .B2(n14601), .A(n10113), .ZN(n10115) );
  AOI211_X1 U12710 ( .C1(n10117), .C2(n14591), .A(n10116), .B(n10115), .ZN(
        n10118) );
  INV_X1 U12711 ( .A(n10118), .ZN(P1_U3252) );
  INV_X1 U12712 ( .A(n10123), .ZN(n10120) );
  AOI21_X1 U12713 ( .B1(n10120), .B2(P2_REG2_REG_10__SCAN_IN), .A(n10119), 
        .ZN(n10122) );
  INV_X1 U12714 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10310) );
  MUX2_X1 U12715 ( .A(n10310), .B(P2_REG2_REG_11__SCAN_IN), .S(n10311), .Z(
        n10121) );
  NAND2_X1 U12716 ( .A1(n10122), .A2(n10121), .ZN(n14783) );
  OAI21_X1 U12717 ( .B1(n10122), .B2(n10121), .A(n14783), .ZN(n10135) );
  OR2_X1 U12718 ( .A1(n10123), .A2(n7884), .ZN(n10128) );
  NAND2_X1 U12719 ( .A1(n10129), .A2(n10128), .ZN(n10126) );
  MUX2_X1 U12720 ( .A(n10124), .B(P2_REG1_REG_11__SCAN_IN), .S(n10311), .Z(
        n10125) );
  NAND2_X1 U12721 ( .A1(n10126), .A2(n10125), .ZN(n14775) );
  MUX2_X1 U12722 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n10124), .S(n10311), .Z(
        n10127) );
  NAND3_X1 U12723 ( .A1(n10129), .A2(n10128), .A3(n10127), .ZN(n10130) );
  AND3_X1 U12724 ( .A1(n14775), .A2(n14814), .A3(n10130), .ZN(n10134) );
  INV_X1 U12725 ( .A(n10311), .ZN(n10131) );
  NAND2_X1 U12726 ( .A1(n14818), .A2(n10131), .ZN(n10132) );
  NAND2_X1 U12727 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11428)
         );
  OAI211_X1 U12728 ( .C1(n14791), .C2(n7159), .A(n10132), .B(n11428), .ZN(
        n10133) );
  AOI211_X1 U12729 ( .C1(n10135), .C2(n14820), .A(n10134), .B(n10133), .ZN(
        n10136) );
  INV_X1 U12730 ( .A(n10136), .ZN(P2_U3225) );
  INV_X1 U12731 ( .A(n10137), .ZN(n10138) );
  OAI222_X1 U12732 ( .A1(P3_U3151), .A2(n14393), .B1(n12962), .B2(n10139), 
        .C1(n12396), .C2(n10138), .ZN(P3_U3279) );
  INV_X1 U12733 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10145) );
  OAI21_X1 U12734 ( .B1(n13143), .B2(n11862), .A(n10140), .ZN(n12104) );
  INV_X1 U12735 ( .A(n12104), .ZN(n10143) );
  NOR2_X1 U12736 ( .A1(n11865), .A2(n10141), .ZN(n10631) );
  OAI21_X1 U12737 ( .B1(n12104), .B2(n13454), .A(n10142), .ZN(n10630) );
  AOI211_X1 U12738 ( .C1(n10143), .C2(n14850), .A(n10631), .B(n10630), .ZN(
        n10530) );
  OR2_X1 U12739 ( .A1(n10530), .A2(n14858), .ZN(n10144) );
  OAI21_X1 U12740 ( .B1(n14859), .B2(n10145), .A(n10144), .ZN(P2_U3430) );
  NOR2_X1 U12741 ( .A1(n13852), .A2(n13812), .ZN(P1_U3085) );
  NAND2_X1 U12742 ( .A1(n12383), .A2(n10681), .ZN(n10146) );
  NAND2_X1 U12743 ( .A1(n10252), .A2(n10146), .ZN(n10330) );
  INV_X1 U12744 ( .A(n10330), .ZN(n10147) );
  OAI21_X1 U12745 ( .B1(n12383), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10147), .ZN(
        n10148) );
  MUX2_X1 U12746 ( .A(n10148), .B(n10147), .S(n14207), .Z(n10149) );
  INV_X1 U12747 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10292) );
  OAI22_X1 U12748 ( .A1(n10150), .A2(n10149), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10292), .ZN(n10152) );
  NOR3_X1 U12749 ( .A1(n11701), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n6762), .ZN(
        n10151) );
  AOI211_X1 U12750 ( .C1(n13852), .C2(P1_ADDR_REG_0__SCAN_IN), .A(n10152), .B(
        n10151), .ZN(n10153) );
  INV_X1 U12751 ( .A(n10153), .ZN(P1_U3243) );
  NAND2_X1 U12752 ( .A1(P1_U4016), .A2(n13897), .ZN(n10154) );
  OAI21_X1 U12753 ( .B1(n13812), .B2(n13625), .A(n10154), .ZN(P1_U3591) );
  AOI211_X1 U12754 ( .C1(n10157), .C2(n10156), .A(n11701), .B(n10155), .ZN(
        n10169) );
  INV_X1 U12755 ( .A(n10158), .ZN(n10161) );
  MUX2_X1 U12756 ( .A(n10049), .B(P1_REG2_REG_7__SCAN_IN), .S(n10159), .Z(
        n10160) );
  NAND2_X1 U12757 ( .A1(n10161), .A2(n10160), .ZN(n10163) );
  OAI211_X1 U12758 ( .C1(n10187), .C2(n10163), .A(n13887), .B(n10162), .ZN(
        n10166) );
  NOR2_X1 U12759 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8437), .ZN(n10164) );
  AOI21_X1 U12760 ( .B1(n13852), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n10164), .ZN(
        n10165) );
  OAI211_X1 U12761 ( .C1(n14601), .C2(n10167), .A(n10166), .B(n10165), .ZN(
        n10168) );
  OR2_X1 U12762 ( .A1(n10169), .A2(n10168), .ZN(P1_U3250) );
  NAND2_X1 U12763 ( .A1(n14051), .A2(P1_U4016), .ZN(n10170) );
  OAI21_X1 U12764 ( .B1(n8023), .B2(n13812), .A(n10170), .ZN(P1_U3579) );
  NAND2_X1 U12765 ( .A1(n14039), .A2(P1_U4016), .ZN(n10171) );
  OAI21_X1 U12766 ( .B1(n7250), .B2(n13812), .A(n10171), .ZN(P1_U3580) );
  OAI21_X1 U12767 ( .B1(n10174), .B2(n10173), .A(n10172), .ZN(n10175) );
  NAND2_X1 U12768 ( .A1(n10175), .A2(n9789), .ZN(n10179) );
  OAI22_X1 U12769 ( .A1(n10176), .A2(n13092), .B1(n10512), .B2(n13094), .ZN(
        n10654) );
  AOI22_X1 U12770 ( .A1(n13099), .A2(n10654), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n10177), .ZN(n10178) );
  OAI211_X1 U12771 ( .C1(n11883), .C2(n13114), .A(n10179), .B(n10178), .ZN(
        P2_U3209) );
  AOI211_X1 U12772 ( .C1(n10182), .C2(n10181), .A(n10180), .B(n11701), .ZN(
        n10193) );
  AND3_X1 U12773 ( .A1(n10185), .A2(n10184), .A3(n10183), .ZN(n10186) );
  NOR3_X1 U12774 ( .A1(n14596), .A2(n10187), .A3(n10186), .ZN(n10192) );
  INV_X1 U12775 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10190) );
  INV_X1 U12776 ( .A(n14601), .ZN(n13860) );
  NAND2_X1 U12777 ( .A1(n13860), .A2(n10188), .ZN(n10189) );
  NAND2_X1 U12778 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n11123) );
  OAI211_X1 U12779 ( .C1(n14605), .C2(n10190), .A(n10189), .B(n11123), .ZN(
        n10191) );
  OR3_X1 U12780 ( .A1(n10193), .A2(n10192), .A3(n10191), .ZN(P1_U3249) );
  INV_X1 U12781 ( .A(n10194), .ZN(n10195) );
  OAI222_X1 U12782 ( .A1(n14413), .A2(P3_U3151), .B1(n12396), .B2(n10195), 
        .C1(n6898), .C2(n12962), .ZN(P3_U3278) );
  XNOR2_X1 U12783 ( .A(n12106), .B(n10196), .ZN(n10662) );
  OAI21_X1 U12784 ( .B1(n10198), .B2(n12106), .A(n10197), .ZN(n10199) );
  NAND2_X1 U12785 ( .A1(n10199), .A2(n13430), .ZN(n10201) );
  NAND2_X1 U12786 ( .A1(n10201), .A2(n10200), .ZN(n10663) );
  AOI211_X1 U12787 ( .C1(n11862), .C2(n11869), .A(n13460), .B(n10656), .ZN(
        n10668) );
  AOI211_X1 U12788 ( .C1(n10662), .C2(n14850), .A(n10663), .B(n10668), .ZN(
        n10637) );
  INV_X1 U12789 ( .A(n11869), .ZN(n11874) );
  INV_X1 U12790 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10202) );
  OAI22_X1 U12791 ( .A1(n13602), .A2(n11874), .B1(n14859), .B2(n10202), .ZN(
        n10203) );
  INV_X1 U12792 ( .A(n10203), .ZN(n10204) );
  OAI21_X1 U12793 ( .B1(n10637), .B2(n14858), .A(n10204), .ZN(P2_U3433) );
  INV_X1 U12794 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10205) );
  MUX2_X1 U12795 ( .A(n10205), .B(P1_REG1_REG_10__SCAN_IN), .S(n10295), .Z(
        n10208) );
  OAI21_X1 U12796 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n10209), .A(n10206), .ZN(
        n10207) );
  NOR2_X1 U12797 ( .A1(n10207), .A2(n10208), .ZN(n10294) );
  AOI211_X1 U12798 ( .C1(n10208), .C2(n10207), .A(n11701), .B(n10294), .ZN(
        n10220) );
  NAND2_X1 U12799 ( .A1(n10209), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10211) );
  MUX2_X1 U12800 ( .A(n8488), .B(P1_REG2_REG_10__SCAN_IN), .S(n10295), .Z(
        n10210) );
  AOI21_X1 U12801 ( .B1(n10212), .B2(n10211), .A(n10210), .ZN(n10293) );
  AND3_X1 U12802 ( .A1(n10212), .A2(n10211), .A3(n10210), .ZN(n10213) );
  NOR3_X1 U12803 ( .A1(n10293), .A2(n10213), .A3(n14596), .ZN(n10219) );
  NOR2_X1 U12804 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10214), .ZN(n10215) );
  AOI21_X1 U12805 ( .B1(n13852), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n10215), 
        .ZN(n10216) );
  OAI21_X1 U12806 ( .B1(n10217), .B2(n14601), .A(n10216), .ZN(n10218) );
  OR3_X1 U12807 ( .A1(n10220), .A2(n10219), .A3(n10218), .ZN(P1_U3253) );
  NAND2_X1 U12808 ( .A1(n10221), .A2(P1_B_REG_SCAN_IN), .ZN(n10223) );
  MUX2_X1 U12809 ( .A(n10223), .B(P1_B_REG_SCAN_IN), .S(n10222), .Z(n10225) );
  INV_X1 U12810 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10227) );
  NOR2_X1 U12811 ( .A1(n10224), .A2(n10222), .ZN(n10226) );
  INV_X1 U12812 ( .A(n10289), .ZN(n10674) );
  NOR4_X1 U12813 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n10231) );
  NOR4_X1 U12814 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n10230) );
  NOR4_X1 U12815 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n10229) );
  NOR4_X1 U12816 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n10228) );
  NAND4_X1 U12817 ( .A1(n10231), .A2(n10230), .A3(n10229), .A4(n10228), .ZN(
        n10236) );
  NOR2_X1 U12818 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n15275) );
  NOR4_X1 U12819 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n10234) );
  NOR4_X1 U12820 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n10233) );
  NOR4_X1 U12821 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n10232) );
  NAND4_X1 U12822 ( .A1(n15275), .A2(n10234), .A3(n10233), .A4(n10232), .ZN(
        n10235) );
  OAI21_X1 U12823 ( .B1(n10236), .B2(n10235), .A(n10322), .ZN(n10270) );
  AND2_X1 U12824 ( .A1(n10272), .A2(n10932), .ZN(n10237) );
  AND2_X1 U12825 ( .A1(n10270), .A2(n10237), .ZN(n10672) );
  AND2_X1 U12826 ( .A1(n10674), .A2(n10672), .ZN(n10241) );
  INV_X1 U12827 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10238) );
  NAND2_X1 U12828 ( .A1(n10322), .A2(n10238), .ZN(n10240) );
  INV_X1 U12829 ( .A(n10224), .ZN(n14199) );
  NAND2_X1 U12830 ( .A1(n10221), .A2(n14199), .ZN(n10239) );
  OR2_X2 U12831 ( .A1(n10247), .A2(n10242), .ZN(n14058) );
  INV_X1 U12832 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10256) );
  OR2_X1 U12833 ( .A1(n8820), .A2(n10242), .ZN(n10274) );
  INV_X1 U12834 ( .A(n14623), .ZN(n10684) );
  AND2_X1 U12835 ( .A1(n10281), .A2(n8820), .ZN(n10246) );
  NOR2_X1 U12836 ( .A1(n12315), .A2(n10246), .ZN(n10676) );
  NAND2_X1 U12837 ( .A1(n10676), .A2(n8883), .ZN(n14631) );
  INV_X1 U12838 ( .A(n10247), .ZN(n10248) );
  NAND2_X1 U12839 ( .A1(n10248), .A2(n14345), .ZN(n14743) );
  NAND2_X1 U12840 ( .A1(n14345), .A2(n8820), .ZN(n10250) );
  INV_X1 U12841 ( .A(n10251), .ZN(n10677) );
  OAI21_X1 U12842 ( .B1(n14729), .B2(n14138), .A(n10677), .ZN(n10254) );
  NOR2_X2 U12843 ( .A1(n10252), .A2(n10277), .ZN(n14050) );
  INV_X1 U12844 ( .A(n14050), .ZN(n14583) );
  NOR2_X1 U12845 ( .A1(n14626), .A2(n14583), .ZN(n10678) );
  INV_X1 U12846 ( .A(n10678), .ZN(n10253) );
  OAI211_X1 U12847 ( .C1(n10274), .C2(n10684), .A(n10254), .B(n10253), .ZN(
        n14168) );
  NAND2_X1 U12848 ( .A1(n15160), .A2(n14168), .ZN(n10255) );
  OAI21_X1 U12849 ( .B1(n15160), .B2(n10256), .A(n10255), .ZN(P1_U3459) );
  INV_X1 U12850 ( .A(n10257), .ZN(n10260) );
  AOI22_X1 U12851 ( .A1(n13846), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n14188), .ZN(n10258) );
  OAI21_X1 U12852 ( .B1(n10260), .B2(n14204), .A(n10258), .ZN(P1_U3341) );
  OAI222_X1 U12853 ( .A1(n13651), .A2(n10260), .B1(n11310), .B2(P2_U3088), 
        .C1(n10259), .C2(n13624), .ZN(P2_U3313) );
  NAND2_X1 U12854 ( .A1(n13812), .A2(n13943), .ZN(n10261) );
  OAI21_X1 U12855 ( .B1(n13812), .B2(n8952), .A(n10261), .ZN(P1_U3584) );
  XNOR2_X1 U12856 ( .A(n10262), .B(n10263), .ZN(n10268) );
  OAI22_X1 U12857 ( .A1(n10264), .A2(n13092), .B1(n7777), .B2(n13094), .ZN(
        n10348) );
  AND2_X1 U12858 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n13161) );
  AOI21_X1 U12859 ( .B1(n13099), .B2(n10348), .A(n13161), .ZN(n10267) );
  INV_X1 U12860 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10265) );
  AOI22_X1 U12861 ( .A1(n13081), .A2(n6828), .B1(n13110), .B2(n10265), .ZN(
        n10266) );
  OAI211_X1 U12862 ( .C1(n10268), .C2(n13070), .A(n10267), .B(n10266), .ZN(
        P2_U3190) );
  NAND2_X1 U12863 ( .A1(n14038), .A2(n13812), .ZN(n10269) );
  OAI21_X1 U12864 ( .B1(n13812), .B2(n6640), .A(n10269), .ZN(P1_U3578) );
  NAND3_X1 U12865 ( .A1(n10673), .A2(n10289), .A3(n10270), .ZN(n14576) );
  INV_X1 U12866 ( .A(n14576), .ZN(n10271) );
  NAND2_X1 U12867 ( .A1(n10271), .A2(n10272), .ZN(n10279) );
  INV_X1 U12868 ( .A(n14564), .ZN(n13782) );
  INV_X1 U12869 ( .A(n10932), .ZN(n10273) );
  NOR2_X1 U12870 ( .A1(n13782), .A2(n10273), .ZN(n14582) );
  INV_X1 U12871 ( .A(n10274), .ZN(n10276) );
  NAND2_X1 U12872 ( .A1(n14711), .A2(n10277), .ZN(n10278) );
  INV_X1 U12873 ( .A(n10282), .ZN(n10285) );
  OAI21_X1 U12874 ( .B1(n10288), .B2(n10354), .A(n10356), .ZN(n10328) );
  NAND2_X1 U12875 ( .A1(n14584), .A2(n14050), .ZN(n13791) );
  INV_X1 U12876 ( .A(n13791), .ZN(n14512) );
  AOI22_X1 U12877 ( .A1(n14580), .A2(n10328), .B1(n14512), .B2(n6863), .ZN(
        n10291) );
  NAND2_X1 U12878 ( .A1(n13739), .A2(n14623), .ZN(n10290) );
  OAI211_X1 U12879 ( .C1(n14582), .C2(n10292), .A(n10291), .B(n10290), .ZN(
        P1_U3232) );
  AOI21_X1 U12880 ( .B1(n10295), .B2(P1_REG2_REG_10__SCAN_IN), .A(n10293), 
        .ZN(n10792) );
  MUX2_X1 U12881 ( .A(n11334), .B(P1_REG2_REG_11__SCAN_IN), .S(n10790), .Z(
        n10791) );
  XNOR2_X1 U12882 ( .A(n10792), .B(n10791), .ZN(n10305) );
  INV_X1 U12883 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10296) );
  MUX2_X1 U12884 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10296), .S(n10790), .Z(
        n10297) );
  NAND2_X1 U12885 ( .A1(n10298), .A2(n10297), .ZN(n10784) );
  OAI21_X1 U12886 ( .B1(n10298), .B2(n10297), .A(n10784), .ZN(n10299) );
  NAND2_X1 U12887 ( .A1(n10299), .A2(n14591), .ZN(n10304) );
  NAND2_X1 U12888 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14516)
         );
  INV_X1 U12889 ( .A(n14516), .ZN(n10302) );
  NOR2_X1 U12890 ( .A1(n14601), .A2(n10300), .ZN(n10301) );
  AOI211_X1 U12891 ( .C1(n13852), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10302), 
        .B(n10301), .ZN(n10303) );
  OAI211_X1 U12892 ( .C1(n14596), .C2(n10305), .A(n10304), .B(n10303), .ZN(
        P1_U3254) );
  XNOR2_X1 U12893 ( .A(n14779), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n14777) );
  OR2_X1 U12894 ( .A1(n10311), .A2(n10124), .ZN(n14774) );
  AND2_X1 U12895 ( .A1(n14777), .A2(n14774), .ZN(n10306) );
  NAND2_X1 U12896 ( .A1(n14775), .A2(n10306), .ZN(n14776) );
  NAND2_X1 U12897 ( .A1(n14779), .A2(n10307), .ZN(n10308) );
  XNOR2_X1 U12898 ( .A(n10312), .B(n15221), .ZN(n10309) );
  AOI21_X1 U12899 ( .B1(n14776), .B2(n10308), .A(n10309), .ZN(n10320) );
  NAND3_X1 U12900 ( .A1(n14776), .A2(n10309), .A3(n10308), .ZN(n11302) );
  NAND2_X1 U12901 ( .A1(n11302), .A2(n14814), .ZN(n10319) );
  NAND2_X1 U12902 ( .A1(n10311), .A2(n10310), .ZN(n14781) );
  MUX2_X1 U12903 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11469), .S(n14779), .Z(
        n14782) );
  AOI21_X1 U12904 ( .B1(n14783), .B2(n14781), .A(n14782), .ZN(n14780) );
  AOI21_X1 U12905 ( .B1(n11469), .B2(n14779), .A(n14780), .ZN(n10314) );
  INV_X1 U12906 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11603) );
  MUX2_X1 U12907 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n11603), .S(n10312), .Z(
        n10313) );
  NAND2_X1 U12908 ( .A1(n10314), .A2(n10313), .ZN(n11308) );
  OAI211_X1 U12909 ( .C1(n10314), .C2(n10313), .A(n11308), .B(n14820), .ZN(
        n10318) );
  NOR2_X1 U12910 ( .A1(n10315), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11664) );
  NOR2_X1 U12911 ( .A1(n14769), .A2(n11309), .ZN(n10316) );
  AOI211_X1 U12912 ( .C1(n14812), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n11664), 
        .B(n10316), .ZN(n10317) );
  OAI211_X1 U12913 ( .C1(n10320), .C2(n10319), .A(n10318), .B(n10317), .ZN(
        P2_U3227) );
  INV_X1 U12914 ( .A(n10221), .ZN(n10324) );
  OR2_X1 U12915 ( .A1(n10323), .A2(n10224), .ZN(n10326) );
  OAI22_X1 U12916 ( .A1(n14673), .A2(P1_D_REG_1__SCAN_IN), .B1(n10324), .B2(
        n10326), .ZN(n10325) );
  INV_X1 U12917 ( .A(n10325), .ZN(P1_U3446) );
  OAI22_X1 U12918 ( .A1(n14673), .A2(P1_D_REG_0__SCAN_IN), .B1(n10222), .B2(
        n10326), .ZN(n10327) );
  INV_X1 U12919 ( .A(n10327), .ZN(P1_U3445) );
  MUX2_X1 U12920 ( .A(n10329), .B(n10328), .S(n14197), .Z(n10332) );
  NAND2_X1 U12921 ( .A1(n10330), .A2(n6762), .ZN(n10331) );
  OAI211_X1 U12922 ( .C1(n10332), .C2(n8882), .A(n13812), .B(n10331), .ZN(
        n13842) );
  INV_X1 U12923 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n10333) );
  INV_X1 U12924 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10691) );
  OAI22_X1 U12925 ( .A1(n14605), .A2(n10333), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10691), .ZN(n10342) );
  XNOR2_X1 U12926 ( .A(n10335), .B(n10334), .ZN(n10340) );
  OAI211_X1 U12927 ( .C1(n10338), .C2(n10337), .A(n14591), .B(n10336), .ZN(
        n10339) );
  OAI21_X1 U12928 ( .B1(n10340), .B2(n14596), .A(n10339), .ZN(n10341) );
  AOI211_X1 U12929 ( .C1(n10343), .C2(n13860), .A(n10342), .B(n10341), .ZN(
        n10344) );
  NAND2_X1 U12930 ( .A1(n13842), .A2(n10344), .ZN(P1_U3245) );
  OAI21_X1 U12931 ( .B1(n10347), .B2(n10346), .A(n10345), .ZN(n10349) );
  AOI21_X1 U12932 ( .B1(n10349), .B2(n13430), .A(n10348), .ZN(n10641) );
  OAI211_X1 U12933 ( .C1(n10657), .C2(n11889), .A(n13372), .B(n10776), .ZN(
        n10643) );
  AND2_X1 U12934 ( .A1(n10641), .A2(n10643), .ZN(n10581) );
  OAI21_X1 U12935 ( .B1(n10351), .B2(n12107), .A(n10350), .ZN(n10640) );
  INV_X1 U12936 ( .A(n13620), .ZN(n11514) );
  OAI22_X1 U12937 ( .A1(n13602), .A2(n11889), .B1(n14859), .B2(n7753), .ZN(
        n10352) );
  AOI21_X1 U12938 ( .B1(n10640), .B2(n11514), .A(n10352), .ZN(n10353) );
  OAI21_X1 U12939 ( .B1(n10581), .B2(n14858), .A(n10353), .ZN(P2_U3439) );
  OR2_X1 U12940 ( .A1(n10354), .A2(n12315), .ZN(n10355) );
  AOI22_X1 U12941 ( .A1(n10923), .A2(n10357), .B1(n10689), .B2(n12319), .ZN(
        n10359) );
  INV_X1 U12942 ( .A(n10360), .ZN(n10361) );
  OAI22_X1 U12943 ( .A1(n12317), .A2(n8827), .B1(n7038), .B2(n12274), .ZN(
        n10918) );
  INV_X1 U12944 ( .A(n12333), .ZN(n11842) );
  OAI22_X1 U12945 ( .A1(n8827), .A2(n12274), .B1(n7038), .B2(n11842), .ZN(
        n10363) );
  XNOR2_X1 U12946 ( .A(n10363), .B(n12334), .ZN(n10919) );
  XOR2_X1 U12947 ( .A(n10920), .B(n10921), .Z(n10367) );
  AND2_X1 U12948 ( .A1(n14584), .A2(n14339), .ZN(n14510) );
  AOI22_X1 U12949 ( .A1(n14512), .A2(n13811), .B1(n14510), .B2(n6863), .ZN(
        n10364) );
  OAI21_X1 U12950 ( .B1(n14582), .B2(n10691), .A(n10364), .ZN(n10365) );
  AOI21_X1 U12951 ( .B1(n13739), .B2(n10694), .A(n10365), .ZN(n10366) );
  OAI21_X1 U12952 ( .B1(n10367), .B2(n14565), .A(n10366), .ZN(P1_U3237) );
  INV_X1 U12953 ( .A(n10368), .ZN(n10369) );
  OAI222_X1 U12954 ( .A1(P3_U3151), .A2(n12634), .B1(n12962), .B2(n10370), 
        .C1(n12396), .C2(n10369), .ZN(P3_U3277) );
  NAND2_X1 U12955 ( .A1(n10614), .A2(n10391), .ZN(n10372) );
  INV_X1 U12956 ( .A(n10492), .ZN(n10375) );
  OR2_X1 U12957 ( .A1(n10383), .A2(n10375), .ZN(n10371) );
  NAND2_X1 U12958 ( .A1(n10372), .A2(n10371), .ZN(n10374) );
  NAND2_X1 U12959 ( .A1(n10376), .A2(n10375), .ZN(n10386) );
  AND3_X1 U12960 ( .A1(n10378), .A2(n10377), .A3(n10397), .ZN(n10382) );
  NAND2_X1 U12961 ( .A1(n10380), .A2(n10379), .ZN(n10381) );
  OAI211_X1 U12962 ( .C1(n10492), .C2(n10383), .A(n10382), .B(n10381), .ZN(
        n10384) );
  NAND2_X1 U12963 ( .A1(n10384), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10385) );
  NOR2_X1 U12964 ( .A1(n12505), .A2(P3_U3151), .ZN(n10508) );
  INV_X1 U12965 ( .A(n10508), .ZN(n10387) );
  NAND2_X1 U12966 ( .A1(n10387), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10395) );
  NAND2_X1 U12967 ( .A1(n14437), .A2(n10492), .ZN(n10389) );
  NAND2_X1 U12968 ( .A1(n15078), .A2(n10905), .ZN(n10390) );
  NAND2_X1 U12969 ( .A1(n15078), .A2(n10391), .ZN(n10392) );
  OR2_X1 U12970 ( .A1(n10396), .A2(n10392), .ZN(n10393) );
  AOI22_X1 U12971 ( .A1(n12535), .A2(n12558), .B1(n10802), .B2(n12521), .ZN(
        n10394) );
  OAI211_X1 U12972 ( .C1(n10616), .C2(n12523), .A(n10395), .B(n10394), .ZN(
        P3_U3172) );
  NAND2_X1 U12973 ( .A1(n10396), .A2(n11108), .ZN(n10400) );
  AOI21_X1 U12974 ( .B1(n10398), .B2(n10397), .A(n9060), .ZN(n10399) );
  MUX2_X1 U12975 ( .A(P3_U3897), .B(n10415), .S(n9384), .Z(n14992) );
  INV_X1 U12976 ( .A(n10399), .ZN(n10401) );
  MUX2_X1 U12977 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n12628), .Z(n14868) );
  OR2_X1 U12978 ( .A1(n14868), .A2(n10416), .ZN(n14875) );
  INV_X1 U12979 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10911) );
  INV_X1 U12980 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10408) );
  MUX2_X1 U12981 ( .A(n10911), .B(n10408), .S(n12628), .Z(n10403) );
  NAND2_X1 U12982 ( .A1(n10403), .A2(n9034), .ZN(n10455) );
  OAI21_X1 U12983 ( .B1(n10403), .B2(n9034), .A(n10455), .ZN(n10404) );
  NOR2_X1 U12984 ( .A1(n10404), .A2(n14875), .ZN(n12572) );
  AOI21_X1 U12985 ( .B1(n14875), .B2(n10404), .A(n12572), .ZN(n10405) );
  INV_X1 U12986 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10497) );
  OAI22_X1 U12987 ( .A1(n15018), .A2(n10405), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10497), .ZN(n10412) );
  INV_X1 U12988 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10406) );
  INV_X1 U12989 ( .A(n14867), .ZN(n10407) );
  OAI21_X1 U12990 ( .B1(n10422), .B2(n14867), .A(n6445), .ZN(n10409) );
  OR2_X1 U12991 ( .A1(n10409), .A2(n10408), .ZN(n10430) );
  NAND2_X1 U12992 ( .A1(n10409), .A2(n10408), .ZN(n10410) );
  NAND2_X1 U12993 ( .A1(n10415), .A2(n6436), .ZN(n14912) );
  AOI21_X1 U12994 ( .B1(n10430), .B2(n10410), .A(n14912), .ZN(n10411) );
  AOI211_X1 U12995 ( .C1(n15030), .C2(P3_ADDR_REG_1__SCAN_IN), .A(n10412), .B(
        n10411), .ZN(n10421) );
  INV_X1 U12996 ( .A(n10413), .ZN(n10414) );
  AND2_X1 U12997 ( .A1(n10416), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n14865) );
  NAND2_X1 U12998 ( .A1(n10417), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10441) );
  OAI21_X1 U12999 ( .B1(n10418), .B2(P3_REG2_REG_1__SCAN_IN), .A(n10442), .ZN(
        n10419) );
  NAND2_X1 U13000 ( .A1(n14866), .A2(n10419), .ZN(n10420) );
  OAI211_X1 U13001 ( .C1(n15033), .C2(n10422), .A(n10421), .B(n10420), .ZN(
        P3_U3183) );
  INV_X1 U13002 ( .A(n10423), .ZN(n10426) );
  INV_X1 U13003 ( .A(n14805), .ZN(n11314) );
  OAI222_X1 U13004 ( .A1(n13624), .A2(n10424), .B1(n13645), .B2(n10426), .C1(
        P2_U3088), .C2(n11314), .ZN(P2_U3312) );
  INV_X1 U13005 ( .A(n11504), .ZN(n11496) );
  OAI222_X1 U13006 ( .A1(n11496), .A2(P1_U3086), .B1(n14204), .B2(n10426), 
        .C1(n10425), .C2(n14201), .ZN(P1_U3340) );
  INV_X1 U13007 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n15177) );
  NAND2_X1 U13008 ( .A1(n12504), .A2(P3_U3897), .ZN(n10427) );
  OAI21_X1 U13009 ( .B1(P3_U3897), .B2(n15177), .A(n10427), .ZN(P3_U3514) );
  INV_X1 U13010 ( .A(n10428), .ZN(n10429) );
  OAI222_X1 U13011 ( .A1(n12962), .A2(n7091), .B1(n12396), .B2(n10429), .C1(
        n12596), .C2(P3_U3151), .ZN(P3_U3276) );
  INV_X1 U13012 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15149) );
  AOI22_X1 U13013 ( .A1(n10541), .A2(n15149), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n10548), .ZN(n10439) );
  INV_X1 U13014 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10435) );
  INV_X1 U13015 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10456) );
  NAND2_X1 U13016 ( .A1(n10430), .A2(n6445), .ZN(n12562) );
  NAND2_X1 U13017 ( .A1(n12563), .A2(n12562), .ZN(n12561) );
  NAND2_X1 U13018 ( .A1(n10459), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10431) );
  NAND2_X1 U13019 ( .A1(n12561), .A2(n10431), .ZN(n10432) );
  XNOR2_X1 U13020 ( .A(n10432), .B(n14889), .ZN(n14890) );
  AND2_X1 U13021 ( .A1(n10432), .A2(n10464), .ZN(n10433) );
  AOI21_X1 U13022 ( .B1(n14890), .B2(P3_REG1_REG_3__SCAN_IN), .A(n10433), .ZN(
        n14910) );
  MUX2_X1 U13023 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n10435), .S(n14907), .Z(
        n14909) );
  INV_X1 U13024 ( .A(n14908), .ZN(n10434) );
  NAND2_X1 U13025 ( .A1(n14922), .A2(n10436), .ZN(n10437) );
  NAND2_X1 U13026 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n14927), .ZN(n14926) );
  NAND2_X1 U13027 ( .A1(n10437), .A2(n14926), .ZN(n10438) );
  NAND2_X1 U13028 ( .A1(n10439), .A2(n10438), .ZN(n10549) );
  OAI21_X1 U13029 ( .B1(n10439), .B2(n10438), .A(n10549), .ZN(n10440) );
  INV_X1 U13030 ( .A(n10440), .ZN(n10454) );
  XNOR2_X1 U13031 ( .A(n12569), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n12566) );
  NAND2_X1 U13032 ( .A1(n10442), .A2(n10441), .ZN(n12565) );
  NAND2_X1 U13033 ( .A1(n12566), .A2(n12565), .ZN(n12564) );
  NAND2_X1 U13034 ( .A1(n10459), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10443) );
  NAND2_X1 U13035 ( .A1(n12564), .A2(n10443), .ZN(n10444) );
  XNOR2_X1 U13036 ( .A(n10444), .B(n14889), .ZN(n14877) );
  INV_X1 U13037 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10730) );
  NAND2_X1 U13038 ( .A1(n14877), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n14879) );
  NAND2_X1 U13039 ( .A1(n10444), .A2(n10464), .ZN(n10445) );
  NAND2_X1 U13040 ( .A1(n14879), .A2(n10445), .ZN(n14896) );
  XNOR2_X1 U13041 ( .A(n14907), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n14895) );
  INV_X1 U13042 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n14918) );
  NAND2_X1 U13043 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n10548), .ZN(n10449) );
  OAI21_X1 U13044 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n10548), .A(n10449), .ZN(
        n10531) );
  XNOR2_X1 U13045 ( .A(n10532), .B(n10531), .ZN(n10450) );
  NAND2_X1 U13046 ( .A1(n14866), .A2(n10450), .ZN(n10453) );
  INV_X1 U13047 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10451) );
  NOR2_X1 U13048 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10451), .ZN(n11004) );
  AOI21_X1 U13049 ( .B1(n15030), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11004), .ZN(
        n10452) );
  OAI211_X1 U13050 ( .C1(n14912), .C2(n10454), .A(n10453), .B(n10452), .ZN(
        n10475) );
  MUX2_X1 U13051 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12628), .Z(n10539) );
  XNOR2_X1 U13052 ( .A(n10539), .B(n10541), .ZN(n10542) );
  MUX2_X1 U13053 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12628), .Z(n10469) );
  INV_X1 U13054 ( .A(n10469), .ZN(n10470) );
  INV_X1 U13055 ( .A(n10455), .ZN(n12571) );
  INV_X1 U13056 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10457) );
  MUX2_X1 U13057 ( .A(n10457), .B(n10456), .S(n12628), .Z(n10458) );
  NAND2_X1 U13058 ( .A1(n10458), .A2(n12569), .ZN(n14881) );
  INV_X1 U13059 ( .A(n10458), .ZN(n10460) );
  NAND2_X1 U13060 ( .A1(n10460), .A2(n10459), .ZN(n10461) );
  AND2_X1 U13061 ( .A1(n14881), .A2(n10461), .ZN(n12570) );
  OAI21_X1 U13062 ( .B1(n12572), .B2(n12571), .A(n12570), .ZN(n14882) );
  INV_X1 U13063 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10462) );
  MUX2_X1 U13064 ( .A(n10730), .B(n10462), .S(n12628), .Z(n10463) );
  NAND2_X1 U13065 ( .A1(n10463), .A2(n14889), .ZN(n10467) );
  INV_X1 U13066 ( .A(n10463), .ZN(n10465) );
  NAND2_X1 U13067 ( .A1(n10465), .A2(n10464), .ZN(n10466) );
  NAND2_X1 U13068 ( .A1(n10467), .A2(n10466), .ZN(n14880) );
  AOI21_X1 U13069 ( .B1(n14882), .B2(n14881), .A(n14880), .ZN(n14884) );
  INV_X1 U13070 ( .A(n10467), .ZN(n10468) );
  XOR2_X1 U13071 ( .A(n14907), .B(n10469), .Z(n14902) );
  MUX2_X1 U13072 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12628), .Z(n10471) );
  AND2_X1 U13073 ( .A1(n10471), .A2(n14922), .ZN(n14919) );
  NOR2_X1 U13074 ( .A1(n10471), .A2(n14922), .ZN(n14920) );
  INV_X1 U13075 ( .A(n14920), .ZN(n10472) );
  XOR2_X1 U13076 ( .A(n10542), .B(n10543), .Z(n10473) );
  NOR2_X1 U13077 ( .A1(n10473), .A2(n15018), .ZN(n10474) );
  AOI211_X1 U13078 ( .C1(n14992), .C2(n10541), .A(n10475), .B(n10474), .ZN(
        n10476) );
  INV_X1 U13079 ( .A(n10476), .ZN(P3_U3188) );
  NAND2_X1 U13080 ( .A1(n10714), .A2(n12659), .ZN(n10477) );
  NAND2_X1 U13081 ( .A1(n10477), .A2(n10585), .ZN(n10478) );
  XNOR2_X1 U13082 ( .A(n10487), .B(n10904), .ZN(n10481) );
  NOR2_X1 U13083 ( .A1(n12558), .A2(n10481), .ZN(n10498) );
  NOR3_X1 U13084 ( .A1(n15085), .A2(n10904), .A3(n10487), .ZN(n10482) );
  NOR2_X1 U13085 ( .A1(n10498), .A2(n10482), .ZN(n10490) );
  INV_X1 U13086 ( .A(n10483), .ZN(n10484) );
  OAI21_X1 U13087 ( .B1(n10484), .B2(n12191), .A(n10906), .ZN(n10485) );
  NAND2_X1 U13088 ( .A1(n10490), .A2(n10486), .ZN(n10500) );
  INV_X1 U13089 ( .A(n10914), .ZN(n10488) );
  NAND3_X1 U13090 ( .A1(n10488), .A2(n9502), .A3(n10487), .ZN(n10489) );
  OAI211_X1 U13091 ( .C1(n10490), .C2(n10906), .A(n10500), .B(n10489), .ZN(
        n10491) );
  NAND2_X1 U13092 ( .A1(n10491), .A2(n12528), .ZN(n10496) );
  OAI22_X1 U13093 ( .A1(n12538), .A2(n10904), .B1(n12516), .B2(n10516), .ZN(
        n10494) );
  AOI21_X1 U13094 ( .B1(n12530), .B2(n12560), .A(n10494), .ZN(n10495) );
  OAI211_X1 U13095 ( .C1(n10508), .C2(n10497), .A(n10496), .B(n10495), .ZN(
        P3_U3162) );
  INV_X1 U13096 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15258) );
  INV_X1 U13097 ( .A(n10498), .ZN(n10499) );
  NAND2_X1 U13098 ( .A1(n10500), .A2(n10499), .ZN(n10501) );
  OAI21_X1 U13099 ( .B1(n10502), .B2(n10501), .A(n10519), .ZN(n10503) );
  NAND2_X1 U13100 ( .A1(n10503), .A2(n12528), .ZN(n10507) );
  OAI22_X1 U13101 ( .A1(n12538), .A2(n10504), .B1(n12516), .B2(n15086), .ZN(
        n10505) );
  AOI21_X1 U13102 ( .B1(n12530), .B2(n12558), .A(n10505), .ZN(n10506) );
  OAI211_X1 U13103 ( .C1(n10508), .C2(n15258), .A(n10507), .B(n10506), .ZN(
        P3_U3177) );
  AOI21_X1 U13104 ( .B1(n10510), .B2(n10509), .A(n6607), .ZN(n10515) );
  OAI22_X1 U13105 ( .A1(n10512), .A2(n13092), .B1(n10511), .B2(n13094), .ZN(
        n10772) );
  AND2_X1 U13106 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n13175) );
  OAI22_X1 U13107 ( .A1(n13114), .A2(n10778), .B1(n13097), .B2(n10777), .ZN(
        n10513) );
  AOI211_X1 U13108 ( .C1(n13099), .C2(n10772), .A(n13175), .B(n10513), .ZN(
        n10514) );
  OAI21_X1 U13109 ( .B1(n10515), .B2(n13070), .A(n10514), .ZN(P2_U3202) );
  NAND2_X1 U13110 ( .A1(n10517), .A2(n10516), .ZN(n10518) );
  AND2_X1 U13111 ( .A1(n10519), .A2(n10518), .ZN(n10521) );
  XNOR2_X1 U13112 ( .A(n10487), .B(n15108), .ZN(n10588) );
  XNOR2_X1 U13113 ( .A(n10588), .B(n15086), .ZN(n10520) );
  OAI211_X1 U13114 ( .C1(n10521), .C2(n10520), .A(n12528), .B(n10589), .ZN(
        n10526) );
  NOR2_X1 U13115 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10522), .ZN(n14885) );
  AOI21_X1 U13116 ( .B1(n12535), .B2(n12555), .A(n14885), .ZN(n10523) );
  OAI21_X1 U13117 ( .B1(n12538), .B2(n15108), .A(n10523), .ZN(n10524) );
  AOI21_X1 U13118 ( .B1(n12530), .B2(n12557), .A(n10524), .ZN(n10525) );
  OAI211_X1 U13119 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12532), .A(n10526), .B(
        n10525), .ZN(P3_U3158) );
  INV_X1 U13120 ( .A(n10527), .ZN(n10577) );
  AOI22_X1 U13121 ( .A1(n11700), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n14188), .ZN(n10528) );
  OAI21_X1 U13122 ( .B1(n10577), .B2(n14204), .A(n10528), .ZN(P1_U3339) );
  NAND2_X1 U13123 ( .A1(n14862), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10529) );
  OAI21_X1 U13124 ( .B1(n10530), .B2(n14862), .A(n10529), .ZN(P2_U3499) );
  INV_X1 U13125 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10885) );
  NAND2_X1 U13126 ( .A1(n12635), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n12580) );
  OR2_X1 U13127 ( .A1(n12635), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n10535) );
  NAND2_X1 U13128 ( .A1(n12580), .A2(n10535), .ZN(n10537) );
  INV_X1 U13129 ( .A(n12581), .ZN(n10536) );
  AOI21_X1 U13130 ( .B1(n10538), .B2(n10537), .A(n10536), .ZN(n10562) );
  INV_X1 U13131 ( .A(n10539), .ZN(n10540) );
  AOI22_X1 U13132 ( .A1(n10543), .A2(n10542), .B1(n10541), .B2(n10540), .ZN(
        n10563) );
  MUX2_X1 U13133 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12628), .Z(n10544) );
  XNOR2_X1 U13134 ( .A(n10544), .B(n10571), .ZN(n10564) );
  OAI22_X1 U13135 ( .A1(n10563), .A2(n10564), .B1(n10544), .B2(n10571), .ZN(
        n10546) );
  MUX2_X1 U13136 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12628), .Z(n12600) );
  XOR2_X1 U13137 ( .A(n12635), .B(n12600), .Z(n10545) );
  NAND2_X1 U13138 ( .A1(n10546), .A2(n10545), .ZN(n12601) );
  OAI21_X1 U13139 ( .B1(n10546), .B2(n10545), .A(n12601), .ZN(n10547) );
  NAND2_X1 U13140 ( .A1(n10547), .A2(n15037), .ZN(n10561) );
  NAND2_X1 U13141 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n10548), .ZN(n10550) );
  NAND2_X1 U13142 ( .A1(n10550), .A2(n10549), .ZN(n10551) );
  NAND2_X1 U13143 ( .A1(n10571), .A2(n10551), .ZN(n10552) );
  XOR2_X1 U13144 ( .A(n10551), .B(n10571), .Z(n10567) );
  NAND2_X1 U13145 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n10567), .ZN(n10566) );
  NAND2_X1 U13146 ( .A1(n10552), .A2(n10566), .ZN(n10555) );
  INV_X1 U13147 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n10553) );
  MUX2_X1 U13148 ( .A(P3_REG1_REG_8__SCAN_IN), .B(n10553), .S(n12635), .Z(
        n10554) );
  NAND2_X1 U13149 ( .A1(n10554), .A2(n10555), .ZN(n12636) );
  OAI21_X1 U13150 ( .B1(n10555), .B2(n10554), .A(n12636), .ZN(n10559) );
  NOR2_X1 U13151 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10556), .ZN(n11216) );
  AOI21_X1 U13152 ( .B1(n15030), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11216), .ZN(
        n10557) );
  OAI21_X1 U13153 ( .B1(n15033), .B2(n12635), .A(n10557), .ZN(n10558) );
  AOI21_X1 U13154 ( .B1(n15035), .B2(n10559), .A(n10558), .ZN(n10560) );
  OAI211_X1 U13155 ( .C1(n10562), .C2(n15043), .A(n10561), .B(n10560), .ZN(
        P3_U3190) );
  XOR2_X1 U13156 ( .A(n10564), .B(n10563), .Z(n10575) );
  XOR2_X1 U13157 ( .A(P3_REG2_REG_7__SCAN_IN), .B(n10565), .Z(n10573) );
  AND2_X1 U13158 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11099) );
  AOI21_X1 U13159 ( .B1(n15030), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11099), .ZN(
        n10570) );
  OAI21_X1 U13160 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n10567), .A(n10566), .ZN(
        n10568) );
  NAND2_X1 U13161 ( .A1(n10568), .A2(n15035), .ZN(n10569) );
  OAI211_X1 U13162 ( .C1(n15033), .C2(n10571), .A(n10570), .B(n10569), .ZN(
        n10572) );
  AOI21_X1 U13163 ( .B1(n14866), .B2(n10573), .A(n10572), .ZN(n10574) );
  OAI21_X1 U13164 ( .B1(n10575), .B2(n15018), .A(n10574), .ZN(P3_U3189) );
  INV_X1 U13165 ( .A(n11316), .ZN(n11533) );
  OAI222_X1 U13166 ( .A1(n13651), .A2(n10577), .B1(n11533), .B2(P2_U3088), 
        .C1(n10576), .C2(n13624), .ZN(P2_U3311) );
  INV_X1 U13167 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n15231) );
  NAND2_X1 U13168 ( .A1(n12734), .A2(P3_U3897), .ZN(n10578) );
  OAI21_X1 U13169 ( .B1(P3_U3897), .B2(n15231), .A(n10578), .ZN(P3_U3515) );
  INV_X1 U13170 ( .A(n13561), .ZN(n11517) );
  NAND2_X1 U13171 ( .A1(n14864), .A2(n14845), .ZN(n13534) );
  OAI22_X1 U13172 ( .A1(n13534), .A2(n11889), .B1(n13552), .B2(n9942), .ZN(
        n10579) );
  AOI21_X1 U13173 ( .B1(n10640), .B2(n11517), .A(n10579), .ZN(n10580) );
  OAI21_X1 U13174 ( .B1(n10581), .B2(n14862), .A(n10580), .ZN(P2_U3502) );
  INV_X1 U13175 ( .A(n10582), .ZN(n10584) );
  OAI222_X1 U13176 ( .A1(P3_U3151), .A2(n10585), .B1(n12396), .B2(n10584), 
        .C1(n10583), .C2(n12962), .ZN(P3_U3275) );
  INV_X1 U13177 ( .A(n10586), .ZN(n10613) );
  OAI222_X1 U13178 ( .A1(n13651), .A2(n10613), .B1(n11534), .B2(P2_U3088), 
        .C1(n10587), .C2(n13650), .ZN(P2_U3310) );
  INV_X1 U13179 ( .A(n10588), .ZN(n10590) );
  XNOR2_X1 U13180 ( .A(n10487), .B(n15069), .ZN(n10591) );
  NAND2_X1 U13181 ( .A1(n10591), .A2(n10893), .ZN(n10805) );
  OAI21_X1 U13182 ( .B1(n10591), .B2(n10893), .A(n10805), .ZN(n10592) );
  AOI21_X1 U13183 ( .B1(n10593), .B2(n10592), .A(n10807), .ZN(n10599) );
  INV_X1 U13184 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10594) );
  NOR2_X1 U13185 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10594), .ZN(n14899) );
  NOR2_X1 U13186 ( .A1(n12516), .A2(n15061), .ZN(n10595) );
  AOI211_X1 U13187 ( .C1(n15069), .C2(n12521), .A(n14899), .B(n10595), .ZN(
        n10596) );
  OAI21_X1 U13188 ( .B1(n15086), .B2(n12508), .A(n10596), .ZN(n10597) );
  AOI21_X1 U13189 ( .B1(n15070), .B2(n12505), .A(n10597), .ZN(n10598) );
  OAI21_X1 U13190 ( .B1(n10599), .B2(n12523), .A(n10598), .ZN(P3_U3170) );
  OAI21_X1 U13191 ( .B1(n10601), .B2(n12110), .A(n10600), .ZN(n10603) );
  OAI22_X1 U13192 ( .A1(n7777), .A2(n13092), .B1(n10602), .B2(n13094), .ZN(
        n10626) );
  AOI21_X1 U13193 ( .B1(n10603), .B2(n13430), .A(n10626), .ZN(n10703) );
  OAI211_X1 U13194 ( .C1(n10775), .C2(n10707), .A(n11036), .B(n13372), .ZN(
        n10705) );
  AND2_X1 U13195 ( .A1(n10703), .A2(n10705), .ZN(n10612) );
  OR2_X1 U13196 ( .A1(n10605), .A2(n10604), .ZN(n10606) );
  NAND2_X1 U13197 ( .A1(n10607), .A2(n10606), .ZN(n10702) );
  INV_X1 U13198 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15167) );
  OAI22_X1 U13199 ( .A1(n13602), .A2(n10707), .B1(n14859), .B2(n15167), .ZN(
        n10608) );
  AOI21_X1 U13200 ( .B1(n10702), .B2(n11514), .A(n10608), .ZN(n10609) );
  OAI21_X1 U13201 ( .B1(n10612), .B2(n14858), .A(n10609), .ZN(P2_U3445) );
  OAI22_X1 U13202 ( .A1(n13534), .A2(n10707), .B1(n14864), .B2(n9949), .ZN(
        n10610) );
  AOI21_X1 U13203 ( .B1(n10702), .B2(n11517), .A(n10610), .ZN(n10611) );
  OAI21_X1 U13204 ( .B1(n10612), .B2(n14862), .A(n10611), .ZN(P2_U3504) );
  INV_X1 U13205 ( .A(n13862), .ZN(n13867) );
  OAI222_X1 U13206 ( .A1(n13867), .A2(P1_U3086), .B1(n14201), .B2(n7642), .C1(
        n10613), .C2(n14204), .ZN(P1_U3338) );
  NOR2_X1 U13207 ( .A1(n10614), .A2(n15089), .ZN(n10615) );
  OAI22_X1 U13208 ( .A1(n10616), .A2(n10615), .B1(n15085), .B2(n15087), .ZN(
        n10830) );
  INV_X1 U13209 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10617) );
  NOR2_X1 U13210 ( .A1(n15141), .A2(n10617), .ZN(n10618) );
  AOI21_X1 U13211 ( .B1(n15141), .B2(n10830), .A(n10618), .ZN(n10619) );
  OAI21_X1 U13212 ( .B1(n10834), .B2(n12939), .A(n10619), .ZN(P3_U3390) );
  OAI21_X1 U13213 ( .B1(n10622), .B2(n10621), .A(n10620), .ZN(n10623) );
  NAND2_X1 U13214 ( .A1(n10623), .A2(n9789), .ZN(n10628) );
  NOR2_X1 U13215 ( .A1(n13097), .A2(n10706), .ZN(n10624) );
  AOI211_X1 U13216 ( .C1(n13099), .C2(n10626), .A(n10625), .B(n10624), .ZN(
        n10627) );
  OAI211_X1 U13217 ( .C1(n10707), .C2(n13114), .A(n10628), .B(n10627), .ZN(
        P2_U3199) );
  AOI21_X1 U13218 ( .B1(n10631), .B2(n10629), .A(n10630), .ZN(n10633) );
  OAI22_X1 U13219 ( .A1(n10633), .A2(n13428), .B1(n10632), .B2(n13472), .ZN(
        n10634) );
  AOI21_X1 U13220 ( .B1(n13428), .B2(P2_REG2_REG_0__SCAN_IN), .A(n10634), .ZN(
        n10635) );
  OAI21_X1 U13221 ( .B1(n13467), .B2(n12104), .A(n10635), .ZN(P2_U3265) );
  AOI22_X1 U13222 ( .A1(n13558), .A2(n11869), .B1(n14862), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n10636) );
  OAI21_X1 U13223 ( .B1(n10637), .B2(n14862), .A(n10636), .ZN(P2_U3500) );
  NAND2_X1 U13224 ( .A1(n10638), .A2(P2_U3947), .ZN(n10639) );
  OAI21_X1 U13225 ( .B1(n11859), .B2(P2_U3947), .A(n10639), .ZN(P2_U3556) );
  INV_X1 U13226 ( .A(n10640), .ZN(n10648) );
  MUX2_X1 U13227 ( .A(n10642), .B(n10641), .S(n13468), .Z(n10647) );
  INV_X2 U13228 ( .A(n13350), .ZN(n13478) );
  INV_X1 U13229 ( .A(n10643), .ZN(n10645) );
  OAI22_X1 U13230 ( .A1(n13463), .A2(n11889), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13472), .ZN(n10644) );
  AOI21_X1 U13231 ( .B1(n13478), .B2(n10645), .A(n10644), .ZN(n10646) );
  OAI211_X1 U13232 ( .C1(n13467), .C2(n10648), .A(n10647), .B(n10646), .ZN(
        P2_U3262) );
  INV_X1 U13233 ( .A(n10651), .ZN(n14840) );
  OAI21_X1 U13234 ( .B1(n10653), .B2(n12105), .A(n10652), .ZN(n10655) );
  AOI21_X1 U13235 ( .B1(n10655), .B2(n13430), .A(n10654), .ZN(n14838) );
  MUX2_X1 U13236 ( .A(n7737), .B(n14838), .S(n13468), .Z(n10661) );
  INV_X1 U13237 ( .A(n10656), .ZN(n10658) );
  AOI211_X1 U13238 ( .C1(n14837), .C2(n10658), .A(n13460), .B(n10657), .ZN(
        n14836) );
  OAI22_X1 U13239 ( .A1(n13463), .A2(n11883), .B1(n13144), .B2(n13472), .ZN(
        n10659) );
  AOI21_X1 U13240 ( .B1(n14836), .B2(n13478), .A(n10659), .ZN(n10660) );
  OAI211_X1 U13241 ( .C1(n13467), .C2(n14840), .A(n10661), .B(n10660), .ZN(
        P2_U3263) );
  INV_X1 U13242 ( .A(n10662), .ZN(n10671) );
  INV_X1 U13243 ( .A(n10663), .ZN(n10665) );
  MUX2_X1 U13244 ( .A(n10665), .B(n10664), .S(n13428), .Z(n10670) );
  OAI22_X1 U13245 ( .A1(n13463), .A2(n11874), .B1(n13472), .B2(n10666), .ZN(
        n10667) );
  AOI21_X1 U13246 ( .B1(n13478), .B2(n10668), .A(n10667), .ZN(n10669) );
  OAI211_X1 U13247 ( .C1(n13467), .C2(n10671), .A(n10670), .B(n10669), .ZN(
        P2_U3264) );
  NAND3_X1 U13248 ( .A1(n10674), .A2(n10673), .A3(n10672), .ZN(n12386) );
  NOR2_X1 U13249 ( .A1(n10675), .A2(n8820), .ZN(n14342) );
  NAND2_X1 U13250 ( .A1(n14610), .A2(n14342), .ZN(n14640) );
  INV_X1 U13251 ( .A(n14352), .ZN(n14618) );
  OAI21_X1 U13252 ( .B1(n14618), .B2(n14045), .A(n10677), .ZN(n10683) );
  INV_X1 U13253 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10681) );
  NOR3_X1 U13254 ( .A1(n10684), .A2(n14345), .A3(n14058), .ZN(n10679) );
  AOI211_X1 U13255 ( .C1(n14636), .C2(P1_REG3_REG_0__SCAN_IN), .A(n10679), .B(
        n10678), .ZN(n10680) );
  MUX2_X1 U13256 ( .A(n10681), .B(n10680), .S(n14610), .Z(n10682) );
  OAI211_X1 U13257 ( .C1(n14640), .C2(n10684), .A(n10683), .B(n10682), .ZN(
        P1_U3293) );
  NAND2_X1 U13258 ( .A1(n14626), .A2(n14676), .ZN(n10685) );
  XNOR2_X1 U13259 ( .A(n10737), .B(n10739), .ZN(n14682) );
  INV_X1 U13260 ( .A(n10687), .ZN(n10688) );
  NAND2_X1 U13261 ( .A1(n14610), .A2(n10688), .ZN(n14641) );
  INV_X1 U13262 ( .A(n14640), .ZN(n14613) );
  NOR2_X1 U13263 ( .A1(n14610), .A2(n10012), .ZN(n10693) );
  NOR2_X1 U13264 ( .A1(n10689), .A2(n14623), .ZN(n14625) );
  AND2_X1 U13265 ( .A1(n14625), .A2(n7038), .ZN(n10818) );
  OAI21_X1 U13266 ( .B1(n14625), .B2(n7038), .A(n14637), .ZN(n10690) );
  OR2_X1 U13267 ( .A1(n10818), .A2(n10690), .ZN(n14683) );
  OAI22_X1 U13268 ( .A1(n14639), .A2(n14683), .B1(n10691), .B2(n14608), .ZN(
        n10692) );
  AOI211_X1 U13269 ( .C1(n14613), .C2(n10694), .A(n10693), .B(n10692), .ZN(
        n10701) );
  OAI21_X1 U13270 ( .B1(n10737), .B2(n10696), .A(n10750), .ZN(n10698) );
  INV_X1 U13271 ( .A(n13811), .ZN(n10751) );
  OAI22_X1 U13272 ( .A1(n14626), .A2(n14622), .B1(n10751), .B2(n14583), .ZN(
        n10697) );
  AOI21_X1 U13273 ( .B1(n10698), .B2(n14138), .A(n10697), .ZN(n10699) );
  OAI21_X1 U13274 ( .B1(n14682), .B2(n14631), .A(n10699), .ZN(n14684) );
  NAND2_X1 U13275 ( .A1(n14684), .A2(n14610), .ZN(n10700) );
  OAI211_X1 U13276 ( .C1(n14682), .C2(n14641), .A(n10701), .B(n10700), .ZN(
        P1_U3291) );
  INV_X1 U13277 ( .A(n10702), .ZN(n10712) );
  MUX2_X1 U13278 ( .A(n10704), .B(n10703), .S(n13468), .Z(n10711) );
  INV_X1 U13279 ( .A(n10705), .ZN(n10709) );
  OAI22_X1 U13280 ( .A1(n13463), .A2(n10707), .B1(n13472), .B2(n10706), .ZN(
        n10708) );
  AOI21_X1 U13281 ( .B1(n10709), .B2(n13478), .A(n10708), .ZN(n10710) );
  OAI211_X1 U13282 ( .C1(n13467), .C2(n10712), .A(n10711), .B(n10710), .ZN(
        P2_U3260) );
  INV_X1 U13283 ( .A(n10713), .ZN(n10716) );
  OAI222_X1 U13284 ( .A1(n12396), .A2(n10716), .B1(n12962), .B2(n10715), .C1(
        P3_U3151), .C2(n10714), .ZN(P3_U3274) );
  XNOR2_X1 U13285 ( .A(n10717), .B(n7114), .ZN(n15107) );
  AOI22_X1 U13286 ( .A1(n10721), .A2(n12942), .B1(n10720), .B2(n10719), .ZN(
        n10723) );
  NAND2_X1 U13287 ( .A1(n10723), .A2(n10722), .ZN(n10729) );
  NAND2_X1 U13288 ( .A1(n10724), .A2(n10905), .ZN(n10912) );
  INV_X1 U13289 ( .A(n10912), .ZN(n15095) );
  NAND2_X1 U13290 ( .A1(n15096), .A2(n15095), .ZN(n11184) );
  AOI22_X1 U13291 ( .A1(n14435), .A2(n12557), .B1(n12555), .B2(n14437), .ZN(
        n10728) );
  OAI211_X1 U13292 ( .C1(n10726), .C2(n7114), .A(n15089), .B(n10725), .ZN(
        n10727) );
  OAI211_X1 U13293 ( .C1(n15107), .C2(n15093), .A(n10728), .B(n10727), .ZN(
        n15109) );
  NAND2_X1 U13294 ( .A1(n15109), .A2(n15096), .ZN(n10734) );
  OR2_X1 U13295 ( .A1(n10729), .A2(n10905), .ZN(n10882) );
  OAI22_X1 U13296 ( .A1(n15096), .A2(n10730), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n15081), .ZN(n10731) );
  AOI21_X1 U13297 ( .B1(n12801), .B2(n10732), .A(n10731), .ZN(n10733) );
  OAI211_X1 U13298 ( .C1(n15107), .C2(n11184), .A(n10734), .B(n10733), .ZN(
        P3_U3230) );
  NAND2_X1 U13299 ( .A1(n10739), .A2(n10738), .ZN(n10741) );
  NAND2_X1 U13300 ( .A1(n8827), .A2(n7038), .ZN(n10740) );
  INV_X1 U13301 ( .A(n10820), .ZN(n10743) );
  NOR2_X1 U13302 ( .A1(n13811), .A2(n14562), .ZN(n10742) );
  INV_X1 U13303 ( .A(n13810), .ZN(n10754) );
  NAND2_X1 U13304 ( .A1(n10754), .A2(n10951), .ZN(n10744) );
  NAND2_X1 U13305 ( .A1(n10949), .A2(n13810), .ZN(n10745) );
  INV_X1 U13306 ( .A(n10863), .ZN(n10862) );
  NAND2_X1 U13307 ( .A1(n6908), .A2(n11017), .ZN(n10746) );
  INV_X1 U13308 ( .A(n10967), .ZN(n10747) );
  NAND2_X1 U13309 ( .A1(n10748), .A2(n10747), .ZN(n10976) );
  OAI21_X1 U13310 ( .B1(n10748), .B2(n10747), .A(n10976), .ZN(n14617) );
  INV_X1 U13311 ( .A(n14617), .ZN(n10760) );
  NAND2_X1 U13312 ( .A1(n10821), .A2(n10820), .ZN(n10823) );
  NAND2_X1 U13313 ( .A1(n10751), .A2(n6906), .ZN(n10752) );
  NAND2_X1 U13314 ( .A1(n10951), .A2(n13810), .ZN(n10753) );
  NAND2_X1 U13315 ( .A1(n10949), .A2(n10754), .ZN(n10755) );
  XNOR2_X1 U13316 ( .A(n10968), .B(n10967), .ZN(n10756) );
  INV_X1 U13317 ( .A(n13807), .ZN(n11191) );
  OAI22_X1 U13318 ( .A1(n11191), .A2(n14583), .B1(n11017), .B2(n14622), .ZN(
        n11121) );
  AOI21_X1 U13319 ( .B1(n10756), .B2(n14138), .A(n11121), .ZN(n14620) );
  INV_X1 U13320 ( .A(n10870), .ZN(n10758) );
  INV_X1 U13321 ( .A(n14612), .ZN(n10757) );
  AOI211_X1 U13322 ( .C1(n14612), .C2(n10758), .A(n14058), .B(n11077), .ZN(
        n14607) );
  AOI21_X1 U13323 ( .B1(n14740), .B2(n14612), .A(n14607), .ZN(n10759) );
  OAI211_X1 U13324 ( .C1(n10760), .C2(n14153), .A(n14620), .B(n10759), .ZN(
        n10762) );
  NAND2_X1 U13325 ( .A1(n10762), .A2(n14748), .ZN(n10761) );
  OAI21_X1 U13326 ( .B1(n14748), .B2(n10056), .A(n10761), .ZN(P1_U3534) );
  INV_X1 U13327 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10764) );
  NAND2_X1 U13328 ( .A1(n10762), .A2(n15160), .ZN(n10763) );
  OAI21_X1 U13329 ( .B1(n15160), .B2(n10764), .A(n10763), .ZN(P1_U3477) );
  OAI21_X1 U13330 ( .B1(n10766), .B2(n12108), .A(n10765), .ZN(n10767) );
  INV_X1 U13331 ( .A(n10767), .ZN(n14848) );
  OAI21_X1 U13332 ( .B1(n10770), .B2(n10769), .A(n10768), .ZN(n10773) );
  NOR2_X1 U13333 ( .A1(n14848), .A2(n9668), .ZN(n10771) );
  AOI211_X1 U13334 ( .C1(n13430), .C2(n10773), .A(n10772), .B(n10771), .ZN(
        n14847) );
  MUX2_X1 U13335 ( .A(n10774), .B(n14847), .S(n13468), .Z(n10781) );
  AOI211_X1 U13336 ( .C1(n14844), .C2(n10776), .A(n13460), .B(n10775), .ZN(
        n14843) );
  OAI22_X1 U13337 ( .A1(n13463), .A2(n10778), .B1(n10777), .B2(n13472), .ZN(
        n10779) );
  AOI21_X1 U13338 ( .B1(n14843), .B2(n13478), .A(n10779), .ZN(n10780) );
  OAI211_X1 U13339 ( .C1(n14848), .C2(n13279), .A(n10781), .B(n10780), .ZN(
        P2_U3261) );
  INV_X1 U13340 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10782) );
  NOR2_X1 U13341 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10782), .ZN(n13750) );
  AOI21_X1 U13342 ( .B1(n13852), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n13750), 
        .ZN(n10783) );
  INV_X1 U13343 ( .A(n10783), .ZN(n10789) );
  INV_X1 U13344 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11621) );
  AOI22_X1 U13345 ( .A1(n10795), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n11621), 
        .B2(n14600), .ZN(n14590) );
  OAI21_X1 U13346 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n10790), .A(n10784), 
        .ZN(n14589) );
  NAND2_X1 U13347 ( .A1(n14590), .A2(n14589), .ZN(n14588) );
  OAI21_X1 U13348 ( .B1(n10795), .B2(P1_REG1_REG_12__SCAN_IN), .A(n14588), 
        .ZN(n10787) );
  INV_X1 U13349 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10785) );
  MUX2_X1 U13350 ( .A(n10785), .B(P1_REG1_REG_13__SCAN_IN), .S(n11269), .Z(
        n10786) );
  NOR2_X1 U13351 ( .A1(n10787), .A2(n10786), .ZN(n11268) );
  AOI211_X1 U13352 ( .C1(n10787), .C2(n10786), .A(n11268), .B(n11701), .ZN(
        n10788) );
  AOI211_X1 U13353 ( .C1(n13860), .C2(n11269), .A(n10789), .B(n10788), .ZN(
        n10801) );
  AOI22_X1 U13354 ( .A1(n10795), .A2(n8521), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n14600), .ZN(n14595) );
  NAND2_X1 U13355 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n10790), .ZN(n10794) );
  OR2_X1 U13356 ( .A1(n10792), .A2(n10791), .ZN(n10793) );
  NAND2_X1 U13357 ( .A1(n10794), .A2(n10793), .ZN(n14594) );
  NOR2_X1 U13358 ( .A1(n14595), .A2(n14594), .ZN(n14593) );
  NOR2_X1 U13359 ( .A1(n10795), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10796) );
  NOR2_X1 U13360 ( .A1(n14593), .A2(n10796), .ZN(n10799) );
  MUX2_X1 U13361 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n10797), .S(n11269), .Z(
        n10798) );
  NAND2_X1 U13362 ( .A1(n10798), .A2(n10799), .ZN(n11263) );
  OAI211_X1 U13363 ( .C1(n10799), .C2(n10798), .A(n13887), .B(n11263), .ZN(
        n10800) );
  NAND2_X1 U13364 ( .A1(n10801), .A2(n10800), .ZN(P1_U3256) );
  INV_X1 U13365 ( .A(n10830), .ZN(n10804) );
  INV_X1 U13366 ( .A(n12894), .ZN(n12884) );
  AOI22_X1 U13367 ( .A1(n12884), .A2(n10802), .B1(n15154), .B2(
        P3_REG1_REG_0__SCAN_IN), .ZN(n10803) );
  OAI21_X1 U13368 ( .B1(n10804), .B2(n15154), .A(n10803), .ZN(P3_U3459) );
  INV_X1 U13369 ( .A(n10805), .ZN(n10806) );
  XNOR2_X1 U13370 ( .A(n10487), .B(n10811), .ZN(n11000) );
  XNOR2_X1 U13371 ( .A(n11000), .B(n15061), .ZN(n10808) );
  AOI21_X1 U13372 ( .B1(n10809), .B2(n10808), .A(n6602), .ZN(n10815) );
  AND2_X1 U13373 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n14925) );
  NOR2_X1 U13374 ( .A1(n12516), .A2(n11102), .ZN(n10810) );
  AOI211_X1 U13375 ( .C1(n10811), .C2(n12521), .A(n14925), .B(n10810), .ZN(
        n10812) );
  OAI21_X1 U13376 ( .B1(n10893), .B2(n12508), .A(n10812), .ZN(n10813) );
  AOI21_X1 U13377 ( .B1(n10899), .B2(n12505), .A(n10813), .ZN(n10814) );
  OAI21_X1 U13378 ( .B1(n10815), .B2(n12523), .A(n10814), .ZN(P3_U3167) );
  OAI21_X1 U13379 ( .B1(n14646), .B2(n14631), .A(n14641), .ZN(n11086) );
  INV_X1 U13380 ( .A(n11086), .ZN(n10875) );
  XNOR2_X1 U13381 ( .A(n10816), .B(n10820), .ZN(n14688) );
  OAI211_X1 U13382 ( .C1(n10818), .C2(n10817), .A(n14637), .B(n10948), .ZN(
        n14690) );
  OAI22_X1 U13383 ( .A1(n14639), .A2(n14690), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14608), .ZN(n10819) );
  AOI21_X1 U13384 ( .B1(n14613), .B2(n6906), .A(n10819), .ZN(n10829) );
  OR2_X1 U13385 ( .A1(n10821), .A2(n10820), .ZN(n10822) );
  NAND2_X1 U13386 ( .A1(n10823), .A2(n10822), .ZN(n10824) );
  NAND2_X1 U13387 ( .A1(n10824), .A2(n14138), .ZN(n14692) );
  NAND2_X1 U13388 ( .A1(n13810), .A2(n14050), .ZN(n10825) );
  OAI21_X1 U13389 ( .B1(n8827), .B2(n14622), .A(n10825), .ZN(n14569) );
  INV_X1 U13390 ( .A(n14569), .ZN(n14691) );
  NAND2_X1 U13391 ( .A1(n14692), .A2(n14691), .ZN(n10826) );
  MUX2_X1 U13392 ( .A(n10826), .B(P1_REG2_REG_3__SCAN_IN), .S(n14646), .Z(
        n10827) );
  INV_X1 U13393 ( .A(n10827), .ZN(n10828) );
  OAI211_X1 U13394 ( .C1(n10875), .C2(n14688), .A(n10829), .B(n10828), .ZN(
        P1_U3290) );
  INV_X1 U13395 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10832) );
  AOI21_X1 U13396 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n15071), .A(n10830), .ZN(
        n10831) );
  MUX2_X1 U13397 ( .A(n10832), .B(n10831), .S(n15096), .Z(n10833) );
  OAI21_X1 U13398 ( .B1(n10834), .B2(n12835), .A(n10833), .ZN(P3_U3233) );
  XNOR2_X1 U13399 ( .A(n10835), .B(n10836), .ZN(n10843) );
  INV_X1 U13400 ( .A(n10853), .ZN(n10840) );
  AND2_X1 U13401 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n13205) );
  NAND2_X1 U13402 ( .A1(n13138), .A2(n13050), .ZN(n10838) );
  NAND2_X1 U13403 ( .A1(n13136), .A2(n13061), .ZN(n10837) );
  AND2_X1 U13404 ( .A1(n10838), .A2(n10837), .ZN(n10849) );
  NOR2_X1 U13405 ( .A1(n13108), .A2(n10849), .ZN(n10839) );
  AOI211_X1 U13406 ( .C1(n13110), .C2(n10840), .A(n13205), .B(n10839), .ZN(
        n10842) );
  NAND2_X1 U13407 ( .A1(n13081), .A2(n11919), .ZN(n10841) );
  OAI211_X1 U13408 ( .C1(n10843), .C2(n13070), .A(n10842), .B(n10841), .ZN(
        P2_U3185) );
  NAND2_X1 U13409 ( .A1(n12559), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n10844) );
  OAI21_X1 U13410 ( .B1(n12674), .B2(n12559), .A(n10844), .ZN(P3_U3519) );
  OAI21_X1 U13411 ( .B1(n10846), .B2(n10847), .A(n10845), .ZN(n11090) );
  INV_X1 U13412 ( .A(n11090), .ZN(n10858) );
  XNOR2_X1 U13413 ( .A(n10848), .B(n10847), .ZN(n10850) );
  OAI21_X1 U13414 ( .B1(n10850), .B2(n13454), .A(n10849), .ZN(n11088) );
  NAND2_X1 U13415 ( .A1(n11088), .A2(n13468), .ZN(n10857) );
  INV_X1 U13416 ( .A(n10993), .ZN(n10851) );
  AOI211_X1 U13417 ( .C1(n11919), .C2(n6600), .A(n13460), .B(n10851), .ZN(
        n11089) );
  INV_X1 U13418 ( .A(n11919), .ZN(n10852) );
  NOR2_X1 U13419 ( .A1(n10852), .A2(n13463), .ZN(n10855) );
  OAI22_X1 U13420 ( .A1(n13468), .A2(n10084), .B1(n10853), .B2(n13472), .ZN(
        n10854) );
  AOI211_X1 U13421 ( .C1(n11089), .C2(n13478), .A(n10855), .B(n10854), .ZN(
        n10856) );
  OAI211_X1 U13422 ( .C1(n13467), .C2(n10858), .A(n10857), .B(n10856), .ZN(
        P2_U3258) );
  INV_X1 U13423 ( .A(n10859), .ZN(n10860) );
  AOI21_X1 U13424 ( .B1(n10862), .B2(n10861), .A(n10860), .ZN(n14703) );
  XNOR2_X1 U13425 ( .A(n10864), .B(n10863), .ZN(n10865) );
  NOR2_X1 U13426 ( .A1(n10865), .A2(n14621), .ZN(n14708) );
  NAND2_X1 U13427 ( .A1(n13810), .A2(n14339), .ZN(n10867) );
  NAND2_X1 U13428 ( .A1(n13808), .A2(n14050), .ZN(n10866) );
  NAND2_X1 U13429 ( .A1(n10867), .A2(n10866), .ZN(n14704) );
  NOR2_X1 U13430 ( .A1(n14708), .A2(n14704), .ZN(n10868) );
  INV_X1 U13431 ( .A(n14646), .ZN(n11595) );
  MUX2_X1 U13432 ( .A(n10869), .B(n10868), .S(n11595), .Z(n10874) );
  AOI211_X1 U13433 ( .C1(n11019), .C2(n10946), .A(n14058), .B(n10870), .ZN(
        n14706) );
  INV_X1 U13434 ( .A(n10871), .ZN(n11022) );
  OAI22_X1 U13435 ( .A1(n14640), .A2(n6908), .B1(n11022), .B2(n14608), .ZN(
        n10872) );
  AOI21_X1 U13436 ( .B1(n14706), .B2(n14060), .A(n10872), .ZN(n10873) );
  OAI211_X1 U13437 ( .C1(n10875), .C2(n14703), .A(n10874), .B(n10873), .ZN(
        P1_U3288) );
  XNOR2_X1 U13438 ( .A(n10876), .B(n11055), .ZN(n10881) );
  OAI211_X1 U13439 ( .C1(n10878), .C2(n11055), .A(n10877), .B(n15089), .ZN(
        n10880) );
  AOI22_X1 U13440 ( .A1(n12553), .A2(n14435), .B1(n14437), .B2(n12551), .ZN(
        n10879) );
  OAI211_X1 U13441 ( .C1(n15093), .C2(n10881), .A(n10880), .B(n10879), .ZN(
        n15126) );
  INV_X1 U13442 ( .A(n15126), .ZN(n10888) );
  INV_X1 U13443 ( .A(n10881), .ZN(n15128) );
  INV_X1 U13444 ( .A(n11184), .ZN(n15057) );
  INV_X1 U13445 ( .A(n10882), .ZN(n15072) );
  NOR2_X1 U13446 ( .A1(n10883), .A2(n15136), .ZN(n15127) );
  AOI22_X1 U13447 ( .A1(n15072), .A2(n15127), .B1(n15071), .B2(n11104), .ZN(
        n10884) );
  OAI21_X1 U13448 ( .B1(n10885), .B2(n15096), .A(n10884), .ZN(n10886) );
  AOI21_X1 U13449 ( .B1(n15128), .B2(n15057), .A(n10886), .ZN(n10887) );
  OAI21_X1 U13450 ( .B1(n10888), .B2(n15075), .A(n10887), .ZN(P3_U3226) );
  XNOR2_X1 U13451 ( .A(n10889), .B(n9096), .ZN(n10897) );
  OAI21_X1 U13452 ( .B1(n10892), .B2(n9096), .A(n10891), .ZN(n10895) );
  OAI22_X1 U13453 ( .A1(n15087), .A2(n11102), .B1(n10893), .B2(n15084), .ZN(
        n10894) );
  AOI21_X1 U13454 ( .B1(n10895), .B2(n15089), .A(n10894), .ZN(n10896) );
  OAI21_X1 U13455 ( .B1(n15093), .B2(n10897), .A(n10896), .ZN(n15117) );
  INV_X1 U13456 ( .A(n15117), .ZN(n10903) );
  INV_X1 U13457 ( .A(n10897), .ZN(n15119) );
  NOR2_X1 U13458 ( .A1(n10898), .A2(n15136), .ZN(n15118) );
  AOI22_X1 U13459 ( .A1(n15072), .A2(n15118), .B1(n15071), .B2(n10899), .ZN(
        n10900) );
  OAI21_X1 U13460 ( .B1(n14918), .B2(n15096), .A(n10900), .ZN(n10901) );
  AOI21_X1 U13461 ( .B1(n15119), .B2(n15057), .A(n10901), .ZN(n10902) );
  OAI21_X1 U13462 ( .B1(n10903), .B2(n15075), .A(n10902), .ZN(P3_U3228) );
  NOR2_X1 U13463 ( .A1(n10904), .A2(n15136), .ZN(n15099) );
  INV_X1 U13464 ( .A(n10905), .ZN(n15079) );
  XNOR2_X1 U13465 ( .A(n9502), .B(n10906), .ZN(n10907) );
  NAND2_X1 U13466 ( .A1(n10907), .A2(n15089), .ZN(n10909) );
  AOI22_X1 U13467 ( .A1(n12557), .A2(n14437), .B1(n14435), .B2(n12560), .ZN(
        n10908) );
  NAND2_X1 U13468 ( .A1(n10909), .A2(n10908), .ZN(n15098) );
  AOI21_X1 U13469 ( .B1(n15099), .B2(n15079), .A(n15098), .ZN(n10910) );
  MUX2_X1 U13470 ( .A(n10911), .B(n10910), .S(n15096), .Z(n10917) );
  NAND2_X1 U13471 ( .A1(n15093), .A2(n10912), .ZN(n10913) );
  XNOR2_X1 U13472 ( .A(n10915), .B(n10914), .ZN(n15100) );
  AOI22_X1 U13473 ( .A1(n14445), .A2(n15100), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15071), .ZN(n10916) );
  NAND2_X1 U13474 ( .A1(n10917), .A2(n10916), .ZN(P3_U3232) );
  AOI22_X1 U13475 ( .A1(n12319), .A2(n13811), .B1(n12333), .B2(n14562), .ZN(
        n10922) );
  XNOR2_X1 U13476 ( .A(n10922), .B(n12334), .ZN(n10924) );
  AOI22_X1 U13477 ( .A1(n10923), .A2(n13811), .B1(n12319), .B2(n14562), .ZN(
        n10925) );
  XNOR2_X1 U13478 ( .A(n10924), .B(n10925), .ZN(n14567) );
  INV_X1 U13479 ( .A(n10924), .ZN(n10927) );
  INV_X1 U13480 ( .A(n10925), .ZN(n10926) );
  AOI22_X1 U13481 ( .A1(n10923), .A2(n13810), .B1(n10949), .B2(n12312), .ZN(
        n11010) );
  INV_X1 U13482 ( .A(n11010), .ZN(n10928) );
  XNOR2_X1 U13483 ( .A(n11011), .B(n10928), .ZN(n11013) );
  AOI22_X1 U13484 ( .A1(n10949), .A2(n12333), .B1(n12319), .B2(n13810), .ZN(
        n10929) );
  XNOR2_X1 U13485 ( .A(n10929), .B(n12334), .ZN(n11012) );
  XNOR2_X1 U13486 ( .A(n11013), .B(n11012), .ZN(n10943) );
  INV_X1 U13487 ( .A(n10930), .ZN(n10931) );
  NAND2_X1 U13488 ( .A1(n14576), .A2(n10931), .ZN(n10936) );
  AND3_X1 U13489 ( .A1(n10282), .A2(n10933), .A3(n10932), .ZN(n10935) );
  NAND2_X1 U13490 ( .A1(n10936), .A2(n10935), .ZN(n10937) );
  INV_X1 U13491 ( .A(n10938), .ZN(n10950) );
  NAND2_X1 U13492 ( .A1(n13811), .A2(n14339), .ZN(n10939) );
  OAI21_X1 U13493 ( .B1(n11017), .B2(n14583), .A(n10939), .ZN(n14696) );
  AND2_X1 U13494 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n13828) );
  AOI21_X1 U13495 ( .B1(n14584), .B2(n14696), .A(n13828), .ZN(n10941) );
  NOR2_X1 U13496 ( .A1(n10951), .A2(n14711), .ZN(n14698) );
  NAND2_X1 U13497 ( .A1(n14564), .A2(n14698), .ZN(n10940) );
  OAI211_X1 U13498 ( .C1(n14572), .C2(n10950), .A(n10941), .B(n10940), .ZN(
        n10942) );
  AOI21_X1 U13499 ( .B1(n10943), .B2(n14580), .A(n10942), .ZN(n10944) );
  INV_X1 U13500 ( .A(n10944), .ZN(P1_U3230) );
  XOR2_X1 U13501 ( .A(n10945), .B(n10954), .Z(n14701) );
  INV_X1 U13502 ( .A(n14701), .ZN(n10959) );
  INV_X1 U13503 ( .A(n10946), .ZN(n10947) );
  AOI211_X1 U13504 ( .C1(n10949), .C2(n10948), .A(n14058), .B(n10947), .ZN(
        n14697) );
  OAI22_X1 U13505 ( .A1(n14610), .A2(n10017), .B1(n10950), .B2(n14608), .ZN(
        n10953) );
  NOR2_X1 U13506 ( .A1(n14640), .A2(n10951), .ZN(n10952) );
  AOI211_X1 U13507 ( .C1(n14060), .C2(n14697), .A(n10953), .B(n10952), .ZN(
        n10958) );
  XNOR2_X1 U13508 ( .A(n10955), .B(n10954), .ZN(n10956) );
  NOR2_X1 U13509 ( .A1(n10956), .A2(n14621), .ZN(n14699) );
  OAI21_X1 U13510 ( .B1(n14699), .B2(n14696), .A(n11595), .ZN(n10957) );
  OAI211_X1 U13511 ( .C1(n10959), .C2(n14352), .A(n10958), .B(n10957), .ZN(
        P1_U3289) );
  INV_X1 U13512 ( .A(n12993), .ZN(n12057) );
  NAND2_X1 U13513 ( .A1(n12057), .A2(P2_U3947), .ZN(n10960) );
  OAI21_X1 U13514 ( .B1(n7677), .B2(P2_U3947), .A(n10960), .ZN(P2_U3560) );
  INV_X1 U13515 ( .A(n10961), .ZN(n10964) );
  OAI22_X1 U13516 ( .A1(n10962), .A2(P3_U3151), .B1(SI_22_), .B2(n12962), .ZN(
        n10963) );
  AOI21_X1 U13517 ( .B1(n10964), .B2(n14320), .A(n10963), .ZN(P3_U3273) );
  INV_X1 U13518 ( .A(n13880), .ZN(n13873) );
  OAI222_X1 U13519 ( .A1(n13873), .A2(P1_U3086), .B1(n14201), .B2(n7649), .C1(
        n10966), .C2(n14204), .ZN(P1_U3337) );
  NAND2_X1 U13520 ( .A1(n12559), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n10965) );
  OAI21_X1 U13521 ( .B1(n12196), .B2(n12559), .A(n10965), .ZN(P3_U3520) );
  INV_X1 U13522 ( .A(n13241), .ZN(n11531) );
  OAI222_X1 U13523 ( .A1(n13650), .A2(n6640), .B1(n11531), .B2(P2_U3088), .C1(
        n13651), .C2(n10966), .ZN(P2_U3309) );
  INV_X1 U13524 ( .A(n13808), .ZN(n10969) );
  NAND2_X1 U13525 ( .A1(n14612), .A2(n10969), .ZN(n10970) );
  AND2_X1 U13526 ( .A1(n11193), .A2(n11191), .ZN(n10972) );
  OR2_X1 U13527 ( .A1(n11193), .A2(n11191), .ZN(n10973) );
  INV_X1 U13528 ( .A(n11144), .ZN(n10979) );
  XNOR2_X1 U13529 ( .A(n11145), .B(n10979), .ZN(n10974) );
  NAND2_X1 U13530 ( .A1(n10974), .A2(n14138), .ZN(n14719) );
  OR2_X1 U13531 ( .A1(n14612), .A2(n13808), .ZN(n10975) );
  INV_X1 U13532 ( .A(n10977), .ZN(n11079) );
  OR2_X1 U13533 ( .A1(n11193), .A2(n13807), .ZN(n10978) );
  OAI21_X1 U13534 ( .B1(n10980), .B2(n10979), .A(n11151), .ZN(n14718) );
  INV_X1 U13535 ( .A(n14717), .ZN(n11416) );
  INV_X1 U13536 ( .A(n11193), .ZN(n14712) );
  XNOR2_X1 U13537 ( .A(n11155), .B(n11416), .ZN(n10981) );
  OAI222_X1 U13538 ( .A1(n10981), .A2(n14058), .B1(n14583), .B2(n11553), .C1(
        n14622), .C2(n11191), .ZN(n14722) );
  AND2_X1 U13539 ( .A1(n14610), .A2(n8883), .ZN(n13991) );
  NAND2_X1 U13540 ( .A1(n14722), .A2(n13991), .ZN(n10983) );
  AOI22_X1 U13541 ( .A1(n14646), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n11419), 
        .B2(n14636), .ZN(n10982) );
  OAI211_X1 U13542 ( .C1(n11416), .C2(n14640), .A(n10983), .B(n10982), .ZN(
        n10984) );
  AOI21_X1 U13543 ( .B1(n14718), .B2(n14618), .A(n10984), .ZN(n10985) );
  OAI21_X1 U13544 ( .B1(n14646), .B2(n14719), .A(n10985), .ZN(P1_U3285) );
  AOI21_X1 U13545 ( .B1(n10986), .B2(n12115), .A(n13454), .ZN(n10988) );
  OAI22_X1 U13546 ( .A1(n11921), .A2(n13092), .B1(n11940), .B2(n13094), .ZN(
        n11131) );
  AOI21_X1 U13547 ( .B1(n10988), .B2(n10987), .A(n11131), .ZN(n11139) );
  OAI21_X1 U13548 ( .B1(n10990), .B2(n12115), .A(n10989), .ZN(n11140) );
  OAI22_X1 U13549 ( .A1(n13468), .A2(n10991), .B1(n11133), .B2(n13472), .ZN(
        n10992) );
  AOI21_X1 U13550 ( .B1(n11932), .B2(n13476), .A(n10992), .ZN(n10997) );
  NAND2_X1 U13551 ( .A1(n10993), .A2(n11932), .ZN(n10994) );
  NAND2_X1 U13552 ( .A1(n10994), .A2(n13372), .ZN(n10995) );
  NOR2_X1 U13553 ( .A1(n11233), .A2(n10995), .ZN(n11137) );
  NAND2_X1 U13554 ( .A1(n11137), .A2(n13478), .ZN(n10996) );
  OAI211_X1 U13555 ( .C1(n11140), .C2(n13467), .A(n10997), .B(n10996), .ZN(
        n10998) );
  INV_X1 U13556 ( .A(n10998), .ZN(n10999) );
  OAI21_X1 U13557 ( .B1(n13428), .B2(n11139), .A(n10999), .ZN(P2_U3257) );
  INV_X1 U13558 ( .A(n15055), .ZN(n11009) );
  NAND2_X1 U13559 ( .A1(n11000), .A2(n15061), .ZN(n11058) );
  INV_X1 U13560 ( .A(n11058), .ZN(n11001) );
  NOR2_X1 U13561 ( .A1(n6602), .A2(n11001), .ZN(n11003) );
  XNOR2_X1 U13562 ( .A(n10487), .B(n15056), .ZN(n11059) );
  XNOR2_X1 U13563 ( .A(n11059), .B(n11102), .ZN(n11002) );
  NAND2_X1 U13564 ( .A1(n11003), .A2(n11002), .ZN(n11096) );
  OAI211_X1 U13565 ( .C1(n11003), .C2(n11002), .A(n11096), .B(n12528), .ZN(
        n11008) );
  AOI21_X1 U13566 ( .B1(n12535), .B2(n12552), .A(n11004), .ZN(n11005) );
  OAI21_X1 U13567 ( .B1(n15056), .B2(n12538), .A(n11005), .ZN(n11006) );
  AOI21_X1 U13568 ( .B1(n12530), .B2(n12554), .A(n11006), .ZN(n11007) );
  OAI211_X1 U13569 ( .C1(n11009), .C2(n12532), .A(n11008), .B(n11007), .ZN(
        P3_U3179) );
  NAND2_X1 U13570 ( .A1(n11019), .A2(n12333), .ZN(n11014) );
  OAI21_X1 U13571 ( .B1(n11017), .B2(n12274), .A(n11014), .ZN(n11015) );
  XNOR2_X1 U13572 ( .A(n11015), .B(n12334), .ZN(n11114) );
  NAND2_X1 U13573 ( .A1(n11019), .A2(n12312), .ZN(n11016) );
  OAI21_X1 U13574 ( .B1(n12317), .B2(n11017), .A(n11016), .ZN(n11113) );
  XNOR2_X1 U13575 ( .A(n11114), .B(n11113), .ZN(n11018) );
  XNOR2_X1 U13576 ( .A(n11112), .B(n11018), .ZN(n11024) );
  AOI22_X1 U13577 ( .A1(n14584), .A2(n14704), .B1(P1_REG3_REG_5__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11021) );
  AND2_X1 U13578 ( .A1(n11019), .A2(n14740), .ZN(n14705) );
  NAND2_X1 U13579 ( .A1(n14564), .A2(n14705), .ZN(n11020) );
  OAI211_X1 U13580 ( .C1(n14572), .C2(n11022), .A(n11021), .B(n11020), .ZN(
        n11023) );
  AOI21_X1 U13581 ( .B1(n11024), .B2(n14580), .A(n11023), .ZN(n11025) );
  INV_X1 U13582 ( .A(n11025), .ZN(P1_U3227) );
  OAI21_X1 U13583 ( .B1(n11028), .B2(n11027), .A(n11026), .ZN(n11166) );
  INV_X1 U13584 ( .A(n11166), .ZN(n11041) );
  OAI21_X1 U13585 ( .B1(n11030), .B2(n12111), .A(n11029), .ZN(n11034) );
  NAND2_X1 U13586 ( .A1(n13137), .A2(n13061), .ZN(n11032) );
  NAND2_X1 U13587 ( .A1(n13139), .A2(n13050), .ZN(n11031) );
  NAND2_X1 U13588 ( .A1(n11032), .A2(n11031), .ZN(n13079) );
  NOR2_X1 U13589 ( .A1(n11041), .A2(n9668), .ZN(n11033) );
  AOI211_X1 U13590 ( .C1(n13430), .C2(n11034), .A(n13079), .B(n11033), .ZN(
        n11163) );
  MUX2_X1 U13591 ( .A(n11035), .B(n11163), .S(n13468), .Z(n11040) );
  AOI21_X1 U13592 ( .B1(n11036), .B2(n13080), .A(n13460), .ZN(n11037) );
  AND2_X1 U13593 ( .A1(n11037), .A2(n6600), .ZN(n11165) );
  INV_X1 U13594 ( .A(n13080), .ZN(n11167) );
  OAI22_X1 U13595 ( .A1(n13463), .A2(n11167), .B1(n13082), .B2(n13472), .ZN(
        n11038) );
  AOI21_X1 U13596 ( .B1(n11165), .B2(n13478), .A(n11038), .ZN(n11039) );
  OAI211_X1 U13597 ( .C1(n11041), .C2(n13279), .A(n11040), .B(n11039), .ZN(
        P2_U3259) );
  INV_X1 U13598 ( .A(n11042), .ZN(n11043) );
  AOI21_X1 U13599 ( .B1(n11046), .B2(n11044), .A(n11043), .ZN(n11049) );
  AOI22_X1 U13600 ( .A1(n12552), .A2(n14435), .B1(n14437), .B2(n12550), .ZN(
        n11048) );
  XNOR2_X1 U13601 ( .A(n11045), .B(n11046), .ZN(n15132) );
  INV_X1 U13602 ( .A(n15093), .ZN(n15054) );
  NAND2_X1 U13603 ( .A1(n15132), .A2(n15054), .ZN(n11047) );
  OAI211_X1 U13604 ( .C1(n11049), .C2(n15049), .A(n11048), .B(n11047), .ZN(
        n15130) );
  INV_X1 U13605 ( .A(n15130), .ZN(n11054) );
  INV_X1 U13606 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11051) );
  NOR2_X1 U13607 ( .A1(n11214), .A2(n15136), .ZN(n15131) );
  AOI22_X1 U13608 ( .A1(n15072), .A2(n15131), .B1(n15071), .B2(n11219), .ZN(
        n11050) );
  OAI21_X1 U13609 ( .B1(n11051), .B2(n15096), .A(n11050), .ZN(n11052) );
  AOI21_X1 U13610 ( .B1(n15132), .B2(n15057), .A(n11052), .ZN(n11053) );
  OAI21_X1 U13611 ( .B1(n11054), .B2(n15075), .A(n11053), .ZN(P3_U3225) );
  XNOR2_X1 U13612 ( .A(n10487), .B(n15135), .ZN(n11340) );
  XNOR2_X1 U13613 ( .A(n11340), .B(n12550), .ZN(n11068) );
  XNOR2_X1 U13614 ( .A(n11055), .B(n12191), .ZN(n11210) );
  XNOR2_X1 U13615 ( .A(n10487), .B(n11214), .ZN(n11062) );
  XNOR2_X1 U13616 ( .A(n11062), .B(n12551), .ZN(n11061) );
  INV_X1 U13617 ( .A(n11061), .ZN(n11212) );
  INV_X1 U13618 ( .A(n11059), .ZN(n11056) );
  NAND2_X1 U13619 ( .A1(n11056), .A2(n11102), .ZN(n11057) );
  NAND4_X1 U13620 ( .A1(n11210), .A2(n11212), .A3(n11058), .A4(n11057), .ZN(
        n11066) );
  NAND2_X1 U13621 ( .A1(n11059), .A2(n12553), .ZN(n11095) );
  OAI21_X1 U13622 ( .B1(n11061), .B2(n11095), .A(n11210), .ZN(n11064) );
  INV_X1 U13623 ( .A(n11210), .ZN(n11060) );
  OAI21_X1 U13624 ( .B1(n11061), .B2(n15046), .A(n11060), .ZN(n11063) );
  AOI22_X1 U13625 ( .A1(n11064), .A2(n11063), .B1(n11062), .B2(n12551), .ZN(
        n11065) );
  INV_X1 U13626 ( .A(n11341), .ZN(n11367) );
  AOI21_X1 U13627 ( .B1(n11068), .B2(n11067), .A(n11367), .ZN(n11073) );
  AND2_X1 U13628 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n14943) );
  NOR2_X1 U13629 ( .A1(n12516), .A2(n11436), .ZN(n11069) );
  AOI211_X1 U13630 ( .C1(n11181), .C2(n12521), .A(n14943), .B(n11069), .ZN(
        n11070) );
  OAI21_X1 U13631 ( .B1(n11097), .B2(n12508), .A(n11070), .ZN(n11071) );
  AOI21_X1 U13632 ( .B1(n11178), .B2(n12505), .A(n11071), .ZN(n11072) );
  OAI21_X1 U13633 ( .B1(n11073), .B2(n12523), .A(n11072), .ZN(P3_U3171) );
  OAI21_X1 U13634 ( .B1(n11075), .B2(n11079), .A(n11074), .ZN(n14715) );
  INV_X1 U13635 ( .A(n11155), .ZN(n11076) );
  OAI211_X1 U13636 ( .C1(n14712), .C2(n11077), .A(n11076), .B(n14637), .ZN(
        n14710) );
  AOI22_X1 U13637 ( .A1(n14613), .A2(n11193), .B1(n11197), .B2(n14636), .ZN(
        n11078) );
  OAI21_X1 U13638 ( .B1(n14710), .B2(n14639), .A(n11078), .ZN(n11085) );
  XNOR2_X1 U13639 ( .A(n11080), .B(n11079), .ZN(n11083) );
  NAND2_X1 U13640 ( .A1(n13808), .A2(n14339), .ZN(n11082) );
  NAND2_X1 U13641 ( .A1(n13806), .A2(n14050), .ZN(n11081) );
  AND2_X1 U13642 ( .A1(n11082), .A2(n11081), .ZN(n11194) );
  OAI21_X1 U13643 ( .B1(n11083), .B2(n14621), .A(n11194), .ZN(n14713) );
  MUX2_X1 U13644 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n14713), .S(n14610), .Z(
        n11084) );
  AOI211_X1 U13645 ( .C1(n11086), .C2(n14715), .A(n11085), .B(n11084), .ZN(
        n11087) );
  INV_X1 U13646 ( .A(n11087), .ZN(P1_U3286) );
  AOI211_X1 U13647 ( .C1(n14850), .C2(n11090), .A(n11089), .B(n11088), .ZN(
        n11094) );
  NOR2_X1 U13648 ( .A1(n14859), .A2(n7825), .ZN(n11091) );
  AOI21_X1 U13649 ( .B1(n13616), .B2(n11919), .A(n11091), .ZN(n11092) );
  OAI21_X1 U13650 ( .B1(n11094), .B2(n14858), .A(n11092), .ZN(P2_U3451) );
  AOI22_X1 U13651 ( .A1(n13558), .A2(n11919), .B1(n14862), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n11093) );
  OAI21_X1 U13652 ( .B1(n11094), .B2(n14862), .A(n11093), .ZN(P2_U3506) );
  NAND2_X1 U13653 ( .A1(n11096), .A2(n11095), .ZN(n11211) );
  XNOR2_X1 U13654 ( .A(n11211), .B(n11210), .ZN(n11106) );
  NOR2_X1 U13655 ( .A1(n12516), .A2(n11097), .ZN(n11098) );
  AOI211_X1 U13656 ( .C1(n11100), .C2(n12521), .A(n11099), .B(n11098), .ZN(
        n11101) );
  OAI21_X1 U13657 ( .B1(n11102), .B2(n12508), .A(n11101), .ZN(n11103) );
  AOI21_X1 U13658 ( .B1(n11104), .B2(n12505), .A(n11103), .ZN(n11105) );
  OAI21_X1 U13659 ( .B1(n11106), .B2(n12523), .A(n11105), .ZN(P3_U3153) );
  NAND2_X1 U13660 ( .A1(n11107), .A2(n14320), .ZN(n11109) );
  OAI211_X1 U13661 ( .C1(n11110), .C2(n12962), .A(n11109), .B(n11108), .ZN(
        P3_U3272) );
  OR2_X1 U13662 ( .A1(n11113), .A2(n11114), .ZN(n11111) );
  NAND2_X1 U13663 ( .A1(n11112), .A2(n11111), .ZN(n11117) );
  INV_X1 U13664 ( .A(n11113), .ZN(n11116) );
  INV_X1 U13665 ( .A(n11114), .ZN(n11115) );
  NAND2_X1 U13666 ( .A1(n14612), .A2(n12333), .ZN(n11119) );
  NAND2_X1 U13667 ( .A1(n12319), .A2(n13808), .ZN(n11118) );
  NAND2_X1 U13668 ( .A1(n11119), .A2(n11118), .ZN(n11120) );
  XNOR2_X1 U13669 ( .A(n11120), .B(n12334), .ZN(n11186) );
  AOI22_X1 U13670 ( .A1(n14612), .A2(n12312), .B1(n10923), .B2(n13808), .ZN(
        n11185) );
  XNOR2_X1 U13671 ( .A(n11186), .B(n11185), .ZN(n11188) );
  XNOR2_X1 U13672 ( .A(n11189), .B(n11188), .ZN(n11126) );
  NAND2_X1 U13673 ( .A1(n14584), .A2(n11121), .ZN(n11122) );
  OAI211_X1 U13674 ( .C1(n14572), .C2(n14609), .A(n11123), .B(n11122), .ZN(
        n11124) );
  AOI21_X1 U13675 ( .B1(n13739), .B2(n14612), .A(n11124), .ZN(n11125) );
  OAI21_X1 U13676 ( .B1(n11126), .B2(n14565), .A(n11125), .ZN(P1_U3239) );
  INV_X1 U13677 ( .A(n11127), .ZN(n11128) );
  AOI21_X1 U13678 ( .B1(n11130), .B2(n11129), .A(n11128), .ZN(n11136) );
  NAND2_X1 U13679 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n13218) );
  NAND2_X1 U13680 ( .A1(n13099), .A2(n11131), .ZN(n11132) );
  OAI211_X1 U13681 ( .C1(n13097), .C2(n11133), .A(n13218), .B(n11132), .ZN(
        n11134) );
  AOI21_X1 U13682 ( .B1(n11932), .B2(n13081), .A(n11134), .ZN(n11135) );
  OAI21_X1 U13683 ( .B1(n11136), .B2(n13070), .A(n11135), .ZN(P2_U3193) );
  INV_X1 U13684 ( .A(n14850), .ZN(n14841) );
  AOI21_X1 U13685 ( .B1(n14845), .B2(n11932), .A(n11137), .ZN(n11138) );
  OAI211_X1 U13686 ( .C1(n11140), .C2(n14841), .A(n11139), .B(n11138), .ZN(
        n11142) );
  NAND2_X1 U13687 ( .A1(n11142), .A2(n14859), .ZN(n11141) );
  OAI21_X1 U13688 ( .B1(n14859), .B2(n7844), .A(n11141), .ZN(P2_U3454) );
  NAND2_X1 U13689 ( .A1(n11142), .A2(n14864), .ZN(n11143) );
  OAI21_X1 U13690 ( .B1(n14864), .B2(n13221), .A(n11143), .ZN(P2_U3507) );
  INV_X1 U13691 ( .A(n13806), .ZN(n11408) );
  INV_X1 U13692 ( .A(n11250), .ZN(n11247) );
  NAND2_X1 U13693 ( .A1(n14739), .A2(n11553), .ZN(n11146) );
  AOI21_X1 U13694 ( .B1(n11147), .B2(n11153), .A(n14621), .ZN(n11149) );
  NAND2_X1 U13695 ( .A1(n13805), .A2(n14339), .ZN(n14498) );
  INV_X1 U13696 ( .A(n14498), .ZN(n11148) );
  AOI21_X1 U13697 ( .B1(n11149), .B2(n11324), .A(n11148), .ZN(n14726) );
  OR2_X1 U13698 ( .A1(n14717), .A2(n13806), .ZN(n11150) );
  OR2_X1 U13699 ( .A1(n14739), .A2(n13805), .ZN(n11152) );
  OAI21_X1 U13700 ( .B1(n11154), .B2(n11153), .A(n11330), .ZN(n14728) );
  NAND2_X1 U13701 ( .A1(n11155), .A2(n11416), .ZN(n11256) );
  XOR2_X1 U13702 ( .A(n14491), .B(n11332), .Z(n11157) );
  NAND2_X1 U13703 ( .A1(n13804), .A2(n14050), .ZN(n14497) );
  INV_X1 U13704 ( .A(n14497), .ZN(n11156) );
  AOI21_X1 U13705 ( .B1(n11157), .B2(n14637), .A(n11156), .ZN(n14725) );
  OAI22_X1 U13706 ( .A1(n14610), .A2(n8488), .B1(n14503), .B2(n14608), .ZN(
        n11158) );
  AOI21_X1 U13707 ( .B1(n14613), .B2(n14491), .A(n11158), .ZN(n11159) );
  OAI21_X1 U13708 ( .B1(n14725), .B2(n14639), .A(n11159), .ZN(n11160) );
  AOI21_X1 U13709 ( .B1(n14728), .B2(n14618), .A(n11160), .ZN(n11161) );
  OAI21_X1 U13710 ( .B1(n14646), .B2(n14726), .A(n11161), .ZN(P1_U3283) );
  INV_X1 U13711 ( .A(n11162), .ZN(n12156) );
  OAI222_X1 U13712 ( .A1(n13249), .A2(P2_U3088), .B1(n13651), .B2(n12156), 
        .C1(n13650), .C2(n8023), .ZN(P2_U3308) );
  INV_X1 U13713 ( .A(n11163), .ZN(n11164) );
  AOI211_X1 U13714 ( .C1(n6743), .C2(n11166), .A(n11165), .B(n11164), .ZN(
        n11171) );
  OAI22_X1 U13715 ( .A1(n13602), .A2(n11167), .B1(n14859), .B2(n7805), .ZN(
        n11168) );
  INV_X1 U13716 ( .A(n11168), .ZN(n11169) );
  OAI21_X1 U13717 ( .B1(n11171), .B2(n14858), .A(n11169), .ZN(P2_U3448) );
  AOI22_X1 U13718 ( .A1(n13558), .A2(n13080), .B1(n14862), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n11170) );
  OAI21_X1 U13719 ( .B1(n11171), .B2(n14862), .A(n11170), .ZN(P2_U3505) );
  XNOR2_X1 U13720 ( .A(n11172), .B(n11174), .ZN(n15138) );
  OAI211_X1 U13721 ( .C1(n11175), .C2(n11174), .A(n11173), .B(n15089), .ZN(
        n11177) );
  AOI22_X1 U13722 ( .A1(n14435), .A2(n12551), .B1(n14437), .B2(n12549), .ZN(
        n11176) );
  OAI211_X1 U13723 ( .C1(n15093), .C2(n15138), .A(n11177), .B(n11176), .ZN(
        n15140) );
  NAND2_X1 U13724 ( .A1(n15140), .A2(n15096), .ZN(n11183) );
  INV_X1 U13725 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n14934) );
  INV_X1 U13726 ( .A(n11178), .ZN(n11179) );
  OAI22_X1 U13727 ( .A1(n15096), .A2(n14934), .B1(n11179), .B2(n15081), .ZN(
        n11180) );
  AOI21_X1 U13728 ( .B1(n12801), .B2(n11181), .A(n11180), .ZN(n11182) );
  OAI211_X1 U13729 ( .C1(n15138), .C2(n11184), .A(n11183), .B(n11182), .ZN(
        P3_U3224) );
  INV_X1 U13730 ( .A(n11185), .ZN(n11187) );
  AOI22_X1 U13731 ( .A1(n11193), .A2(n12333), .B1(n12319), .B2(n13807), .ZN(
        n11190) );
  XNOR2_X1 U13732 ( .A(n11190), .B(n12334), .ZN(n11401) );
  NOR2_X1 U13733 ( .A1(n12317), .A2(n11191), .ZN(n11192) );
  AOI21_X1 U13734 ( .B1(n11193), .B2(n12312), .A(n11192), .ZN(n11402) );
  XNOR2_X1 U13735 ( .A(n11401), .B(n11402), .ZN(n11403) );
  XNOR2_X1 U13736 ( .A(n11404), .B(n11403), .ZN(n11199) );
  INV_X1 U13737 ( .A(n14572), .ZN(n13794) );
  INV_X1 U13738 ( .A(n14584), .ZN(n14496) );
  OAI22_X1 U13739 ( .A1(n14496), .A2(n11194), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8437), .ZN(n11196) );
  NOR2_X1 U13740 ( .A1(n14577), .A2(n14712), .ZN(n11195) );
  AOI211_X1 U13741 ( .C1(n13794), .C2(n11197), .A(n11196), .B(n11195), .ZN(
        n11198) );
  OAI21_X1 U13742 ( .B1(n11199), .B2(n14565), .A(n11198), .ZN(P1_U3213) );
  OAI21_X1 U13743 ( .B1(n11202), .B2(n11201), .A(n11200), .ZN(n11203) );
  NAND2_X1 U13744 ( .A1(n11203), .A2(n9789), .ZN(n11209) );
  INV_X1 U13745 ( .A(n13473), .ZN(n11207) );
  NAND2_X1 U13746 ( .A1(n13136), .A2(n13050), .ZN(n11205) );
  NAND2_X1 U13747 ( .A1(n13134), .A2(n13061), .ZN(n11204) );
  AND2_X1 U13748 ( .A1(n11205), .A2(n11204), .ZN(n11238) );
  NAND2_X1 U13749 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n14771) );
  OAI21_X1 U13750 ( .B1(n13108), .B2(n11238), .A(n14771), .ZN(n11206) );
  AOI21_X1 U13751 ( .B1(n11207), .B2(n13110), .A(n11206), .ZN(n11208) );
  OAI211_X1 U13752 ( .C1(n11242), .C2(n13114), .A(n11209), .B(n11208), .ZN(
        P2_U3203) );
  MUX2_X1 U13753 ( .A(n12552), .B(n11211), .S(n11210), .Z(n11213) );
  XNOR2_X1 U13754 ( .A(n11213), .B(n11212), .ZN(n11221) );
  NOR2_X1 U13755 ( .A1(n12538), .A2(n11214), .ZN(n11215) );
  AOI211_X1 U13756 ( .C1(n12535), .C2(n12550), .A(n11216), .B(n11215), .ZN(
        n11217) );
  OAI21_X1 U13757 ( .B1(n15046), .B2(n12508), .A(n11217), .ZN(n11218) );
  AOI21_X1 U13758 ( .B1(n11219), .B2(n12505), .A(n11218), .ZN(n11220) );
  OAI21_X1 U13759 ( .B1(n11221), .B2(n12523), .A(n11220), .ZN(P3_U3161) );
  OAI211_X1 U13760 ( .C1(n11223), .C2(n11226), .A(n11222), .B(n15089), .ZN(
        n11225) );
  AOI22_X1 U13761 ( .A1(n14436), .A2(n14437), .B1(n14435), .B2(n12550), .ZN(
        n11224) );
  NAND2_X1 U13762 ( .A1(n11225), .A2(n11224), .ZN(n11351) );
  INV_X1 U13763 ( .A(n11351), .ZN(n11231) );
  XNOR2_X1 U13764 ( .A(n11227), .B(n11226), .ZN(n11352) );
  AOI22_X1 U13765 ( .A1(n15075), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n15071), 
        .B2(n11374), .ZN(n11228) );
  OAI21_X1 U13766 ( .B1(n12835), .B2(n11356), .A(n11228), .ZN(n11229) );
  AOI21_X1 U13767 ( .B1(n11352), .B2(n14445), .A(n11229), .ZN(n11230) );
  OAI21_X1 U13768 ( .B1(n11231), .B2(n15075), .A(n11230), .ZN(P3_U3223) );
  XNOR2_X1 U13769 ( .A(n11232), .B(n11236), .ZN(n13471) );
  OAI21_X1 U13770 ( .B1(n11233), .B2(n11242), .A(n13372), .ZN(n11234) );
  NOR2_X1 U13771 ( .A1(n11234), .A2(n11279), .ZN(n13479) );
  OAI211_X1 U13772 ( .C1(n11237), .C2(n11236), .A(n11235), .B(n13430), .ZN(
        n11239) );
  NAND2_X1 U13773 ( .A1(n11239), .A2(n11238), .ZN(n13469) );
  AOI211_X1 U13774 ( .C1(n14850), .C2(n13471), .A(n13479), .B(n13469), .ZN(
        n11245) );
  AOI22_X1 U13775 ( .A1(n13477), .A2(n13558), .B1(n14862), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11240) );
  OAI21_X1 U13776 ( .B1(n11245), .B2(n14862), .A(n11240), .ZN(P2_U3508) );
  INV_X1 U13777 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11241) );
  OAI22_X1 U13778 ( .A1(n11242), .A2(n13602), .B1(n14859), .B2(n11241), .ZN(
        n11243) );
  INV_X1 U13779 ( .A(n11243), .ZN(n11244) );
  OAI21_X1 U13780 ( .B1(n11245), .B2(n14858), .A(n11244), .ZN(P2_U3457) );
  OAI21_X1 U13781 ( .B1(n11248), .B2(n11247), .A(n11246), .ZN(n11254) );
  OAI22_X1 U13782 ( .A1(n11408), .A2(n14622), .B1(n11828), .B2(n14583), .ZN(
        n11253) );
  OAI21_X1 U13783 ( .B1(n11251), .B2(n11250), .A(n11249), .ZN(n11260) );
  INV_X1 U13784 ( .A(n11260), .ZN(n14744) );
  NOR2_X1 U13785 ( .A1(n14744), .A2(n14631), .ZN(n11252) );
  AOI211_X1 U13786 ( .C1(n14138), .C2(n11254), .A(n11253), .B(n11252), .ZN(
        n14742) );
  INV_X1 U13787 ( .A(n14641), .ZN(n14066) );
  INV_X1 U13788 ( .A(n11332), .ZN(n11255) );
  AOI211_X1 U13789 ( .C1(n14739), .C2(n11256), .A(n14058), .B(n11255), .ZN(
        n14738) );
  NAND2_X1 U13790 ( .A1(n14738), .A2(n14060), .ZN(n11258) );
  AOI22_X1 U13791 ( .A1(n14646), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n11561), 
        .B2(n14636), .ZN(n11257) );
  OAI211_X1 U13792 ( .C1(n6900), .C2(n14640), .A(n11258), .B(n11257), .ZN(
        n11259) );
  AOI21_X1 U13793 ( .B1(n11260), .B2(n14066), .A(n11259), .ZN(n11261) );
  OAI21_X1 U13794 ( .B1(n14742), .B2(n14646), .A(n11261), .ZN(P1_U3284) );
  NAND2_X1 U13795 ( .A1(n13846), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11265) );
  MUX2_X1 U13796 ( .A(n11594), .B(P1_REG2_REG_14__SCAN_IN), .S(n13846), .Z(
        n11262) );
  INV_X1 U13797 ( .A(n11262), .ZN(n13844) );
  INV_X1 U13798 ( .A(n11269), .ZN(n11264) );
  OAI21_X1 U13799 ( .B1(n11264), .B2(n10797), .A(n11263), .ZN(n13845) );
  NAND2_X1 U13800 ( .A1(n13844), .A2(n13845), .ZN(n13843) );
  NAND2_X1 U13801 ( .A1(n11265), .A2(n13843), .ZN(n11503) );
  XNOR2_X1 U13802 ( .A(n11504), .B(n11503), .ZN(n11266) );
  NOR2_X1 U13803 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n11266), .ZN(n11505) );
  AOI21_X1 U13804 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n11266), .A(n11505), 
        .ZN(n11277) );
  INV_X1 U13805 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11267) );
  MUX2_X1 U13806 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n11267), .S(n13846), .Z(
        n13849) );
  NAND2_X1 U13807 ( .A1(n13849), .A2(n13848), .ZN(n13847) );
  INV_X1 U13808 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11270) );
  OAI21_X1 U13809 ( .B1(n11271), .B2(n11270), .A(n11497), .ZN(n11272) );
  NAND2_X1 U13810 ( .A1(n11272), .A2(n14591), .ZN(n11276) );
  INV_X1 U13811 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n11273) );
  NAND2_X1 U13812 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n13789)
         );
  OAI21_X1 U13813 ( .B1(n14605), .B2(n11273), .A(n13789), .ZN(n11274) );
  AOI21_X1 U13814 ( .B1(n11504), .B2(n13860), .A(n11274), .ZN(n11275) );
  OAI211_X1 U13815 ( .C1(n11277), .C2(n14596), .A(n11276), .B(n11275), .ZN(
        P1_U3258) );
  XNOR2_X1 U13816 ( .A(n11278), .B(n11285), .ZN(n11381) );
  INV_X1 U13817 ( .A(n11381), .ZN(n11292) );
  INV_X1 U13818 ( .A(n11279), .ZN(n11280) );
  AOI211_X1 U13819 ( .C1(n11946), .C2(n11280), .A(n13460), .B(n11450), .ZN(
        n11380) );
  NOR2_X1 U13820 ( .A1(n11383), .A2(n13463), .ZN(n11283) );
  OAI22_X1 U13821 ( .A1(n13468), .A2(n11281), .B1(n11297), .B2(n13472), .ZN(
        n11282) );
  AOI211_X1 U13822 ( .C1(n11380), .C2(n13478), .A(n11283), .B(n11282), .ZN(
        n11291) );
  OAI211_X1 U13823 ( .C1(n11286), .C2(n11285), .A(n11284), .B(n13430), .ZN(
        n11289) );
  NAND2_X1 U13824 ( .A1(n13135), .A2(n13050), .ZN(n11288) );
  NAND2_X1 U13825 ( .A1(n13133), .A2(n13061), .ZN(n11287) );
  AND2_X1 U13826 ( .A1(n11288), .A2(n11287), .ZN(n11296) );
  NAND2_X1 U13827 ( .A1(n11289), .A2(n11296), .ZN(n11379) );
  NAND2_X1 U13828 ( .A1(n11379), .A2(n13468), .ZN(n11290) );
  OAI211_X1 U13829 ( .C1(n11292), .C2(n13467), .A(n11291), .B(n11290), .ZN(
        P2_U3255) );
  XNOR2_X1 U13830 ( .A(n11294), .B(n11293), .ZN(n11301) );
  OAI21_X1 U13831 ( .B1(n13108), .B2(n11296), .A(n11295), .ZN(n11299) );
  NOR2_X1 U13832 ( .A1(n13097), .A2(n11297), .ZN(n11298) );
  AOI211_X1 U13833 ( .C1(n11946), .C2(n13081), .A(n11299), .B(n11298), .ZN(
        n11300) );
  OAI21_X1 U13834 ( .B1(n11301), .B2(n13070), .A(n11300), .ZN(P2_U3189) );
  OAI21_X1 U13835 ( .B1(n15221), .B2(n11309), .A(n11302), .ZN(n14798) );
  XNOR2_X1 U13836 ( .A(n11310), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n14797) );
  NAND2_X1 U13837 ( .A1(n14798), .A2(n14797), .ZN(n14796) );
  OAI21_X1 U13838 ( .B1(n11310), .B2(n11303), .A(n14796), .ZN(n11304) );
  NAND2_X1 U13839 ( .A1(n14805), .A2(n11304), .ZN(n11305) );
  XNOR2_X1 U13840 ( .A(n11314), .B(n11304), .ZN(n14807) );
  NAND2_X1 U13841 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n14807), .ZN(n14806) );
  NAND2_X1 U13842 ( .A1(n11305), .A2(n14806), .ZN(n11307) );
  XNOR2_X1 U13843 ( .A(n11316), .B(n13553), .ZN(n11306) );
  NAND2_X1 U13844 ( .A1(n11306), .A2(n11307), .ZN(n11532) );
  OAI211_X1 U13845 ( .C1(n11307), .C2(n11306), .A(n14814), .B(n11532), .ZN(
        n11322) );
  NAND2_X1 U13846 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n13018)
         );
  INV_X1 U13847 ( .A(n11310), .ZN(n14793) );
  OAI21_X1 U13848 ( .B1(n11603), .B2(n11309), .A(n11308), .ZN(n11311) );
  NAND2_X1 U13849 ( .A1(n14793), .A2(n11311), .ZN(n11312) );
  XNOR2_X1 U13850 ( .A(n11311), .B(n11310), .ZN(n14795) );
  NAND2_X1 U13851 ( .A1(n14795), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n14794) );
  NAND2_X1 U13852 ( .A1(n11312), .A2(n14794), .ZN(n11313) );
  NAND2_X1 U13853 ( .A1(n14805), .A2(n11313), .ZN(n11315) );
  XNOR2_X1 U13854 ( .A(n11314), .B(n11313), .ZN(n14804) );
  NAND2_X1 U13855 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14804), .ZN(n14803) );
  NAND2_X1 U13856 ( .A1(n11315), .A2(n14803), .ZN(n11318) );
  INV_X1 U13857 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13462) );
  MUX2_X1 U13858 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n13462), .S(n11316), .Z(
        n11317) );
  NAND2_X1 U13859 ( .A1(n11317), .A2(n11318), .ZN(n11527) );
  OAI211_X1 U13860 ( .C1(n11318), .C2(n11317), .A(n14820), .B(n11527), .ZN(
        n11319) );
  NAND2_X1 U13861 ( .A1(n13018), .A2(n11319), .ZN(n11320) );
  AOI21_X1 U13862 ( .B1(n14812), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n11320), 
        .ZN(n11321) );
  OAI211_X1 U13863 ( .C1(n14769), .C2(n11533), .A(n11322), .B(n11321), .ZN(
        P2_U3230) );
  OR2_X1 U13864 ( .A1(n14491), .A2(n11828), .ZN(n11323) );
  XNOR2_X1 U13865 ( .A(n11479), .B(n11477), .ZN(n11325) );
  NAND2_X1 U13866 ( .A1(n11325), .A2(n14138), .ZN(n11328) );
  OAI22_X1 U13867 ( .A1(n11828), .A2(n14622), .B1(n11843), .B2(n14583), .ZN(
        n11326) );
  INV_X1 U13868 ( .A(n11326), .ZN(n11327) );
  NAND2_X1 U13869 ( .A1(n11328), .A2(n11327), .ZN(n14533) );
  INV_X1 U13870 ( .A(n14533), .ZN(n11339) );
  OR2_X1 U13871 ( .A1(n14491), .A2(n14509), .ZN(n11329) );
  OAI21_X1 U13872 ( .B1(n11331), .B2(n11477), .A(n11475), .ZN(n14535) );
  INV_X1 U13873 ( .A(n11486), .ZN(n11487) );
  OAI211_X1 U13874 ( .C1(n14532), .C2(n11333), .A(n11487), .B(n14637), .ZN(
        n14531) );
  OAI22_X1 U13875 ( .A1(n11595), .A2(n11334), .B1(n14518), .B2(n14608), .ZN(
        n11335) );
  AOI21_X1 U13876 ( .B1(n11835), .B2(n14613), .A(n11335), .ZN(n11336) );
  OAI21_X1 U13877 ( .B1(n14531), .B2(n14639), .A(n11336), .ZN(n11337) );
  AOI21_X1 U13878 ( .B1(n14535), .B2(n14618), .A(n11337), .ZN(n11338) );
  OAI21_X1 U13879 ( .B1(n11339), .B2(n14646), .A(n11338), .ZN(P1_U3282) );
  XNOR2_X1 U13880 ( .A(n10487), .B(n11356), .ZN(n11342) );
  XNOR2_X1 U13881 ( .A(n11342), .B(n12549), .ZN(n11371) );
  NOR2_X1 U13882 ( .A1(n11340), .A2(n12550), .ZN(n11366) );
  XNOR2_X1 U13883 ( .A(n7304), .B(n14436), .ZN(n11344) );
  XNOR2_X1 U13884 ( .A(n11389), .B(n11344), .ZN(n11350) );
  NAND2_X1 U13885 ( .A1(n12505), .A2(n11438), .ZN(n11346) );
  AND2_X1 U13886 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n14973) );
  AOI21_X1 U13887 ( .B1(n12535), .B2(n12548), .A(n14973), .ZN(n11345) );
  OAI211_X1 U13888 ( .C1(n11436), .C2(n12508), .A(n11346), .B(n11345), .ZN(
        n11347) );
  AOI21_X1 U13889 ( .B1(n11348), .B2(n12521), .A(n11347), .ZN(n11349) );
  OAI21_X1 U13890 ( .B1(n11350), .B2(n12523), .A(n11349), .ZN(P3_U3176) );
  AOI21_X1 U13891 ( .B1(n15101), .B2(n11352), .A(n11351), .ZN(n11359) );
  INV_X1 U13892 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n12640) );
  OAI22_X1 U13893 ( .A1(n12894), .A2(n11356), .B1(n15157), .B2(n12640), .ZN(
        n11353) );
  INV_X1 U13894 ( .A(n11353), .ZN(n11354) );
  OAI21_X1 U13895 ( .B1(n11359), .B2(n15154), .A(n11354), .ZN(P3_U3469) );
  INV_X1 U13896 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n11355) );
  OAI22_X1 U13897 ( .A1(n11356), .A2(n12939), .B1(n15141), .B2(n11355), .ZN(
        n11357) );
  INV_X1 U13898 ( .A(n11357), .ZN(n11358) );
  OAI21_X1 U13899 ( .B1(n11359), .B2(n15142), .A(n11358), .ZN(P3_U3420) );
  INV_X1 U13900 ( .A(n11360), .ZN(n11377) );
  OAI222_X1 U13901 ( .A1(n13651), .A2(n11377), .B1(n13624), .B2(n7250), .C1(
        P2_U3088), .C2(n8222), .ZN(P2_U3307) );
  INV_X1 U13902 ( .A(n12550), .ZN(n11365) );
  INV_X1 U13903 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11361) );
  NOR2_X1 U13904 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11361), .ZN(n14953) );
  AOI21_X1 U13905 ( .B1(n12535), .B2(n14436), .A(n14953), .ZN(n11364) );
  NAND2_X1 U13906 ( .A1(n12521), .A2(n11362), .ZN(n11363) );
  OAI211_X1 U13907 ( .C1(n12508), .C2(n11365), .A(n11364), .B(n11363), .ZN(
        n11373) );
  OR2_X1 U13908 ( .A1(n11367), .A2(n11366), .ZN(n11370) );
  INV_X1 U13909 ( .A(n11368), .ZN(n11369) );
  AOI211_X1 U13910 ( .C1(n11371), .C2(n11370), .A(n12523), .B(n11369), .ZN(
        n11372) );
  AOI211_X1 U13911 ( .C1(n11374), .C2(n12505), .A(n11373), .B(n11372), .ZN(
        n11375) );
  INV_X1 U13912 ( .A(n11375), .ZN(P3_U3157) );
  OAI222_X1 U13913 ( .A1(P1_U3086), .A2(n11378), .B1(n14204), .B2(n11377), 
        .C1(n11376), .C2(n14201), .ZN(P1_U3335) );
  AOI211_X1 U13914 ( .C1(n14850), .C2(n11381), .A(n11380), .B(n11379), .ZN(
        n11387) );
  INV_X1 U13915 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11382) );
  OAI22_X1 U13916 ( .A1(n11383), .A2(n13602), .B1(n14859), .B2(n11382), .ZN(
        n11384) );
  INV_X1 U13917 ( .A(n11384), .ZN(n11385) );
  OAI21_X1 U13918 ( .B1(n11387), .B2(n14858), .A(n11385), .ZN(P2_U3460) );
  AOI22_X1 U13919 ( .A1(n11946), .A2(n13558), .B1(n14862), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n11386) );
  OAI21_X1 U13920 ( .B1(n11387), .B2(n14862), .A(n11386), .ZN(P2_U3509) );
  NOR2_X1 U13921 ( .A1(n7304), .A2(n14436), .ZN(n11388) );
  XNOR2_X1 U13922 ( .A(n14443), .B(n12191), .ZN(n11543) );
  XNOR2_X1 U13923 ( .A(n11543), .B(n11675), .ZN(n11390) );
  XNOR2_X1 U13924 ( .A(n11542), .B(n11390), .ZN(n11397) );
  NAND2_X1 U13925 ( .A1(n12505), .A2(n14440), .ZN(n11393) );
  INV_X1 U13926 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11391) );
  NOR2_X1 U13927 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11391), .ZN(n14993) );
  AOI21_X1 U13928 ( .B1(n12535), .B2(n14438), .A(n14993), .ZN(n11392) );
  OAI211_X1 U13929 ( .C1(n11394), .C2(n12508), .A(n11393), .B(n11392), .ZN(
        n11395) );
  AOI21_X1 U13930 ( .B1(n14443), .B2(n12521), .A(n11395), .ZN(n11396) );
  OAI21_X1 U13931 ( .B1(n11397), .B2(n12523), .A(n11396), .ZN(P3_U3164) );
  OAI222_X1 U13932 ( .A1(n11400), .A2(P3_U3151), .B1(n12396), .B2(n11399), 
        .C1(n11398), .C2(n12962), .ZN(P3_U3271) );
  NAND2_X1 U13933 ( .A1(n14717), .A2(n12333), .ZN(n11406) );
  NAND2_X1 U13934 ( .A1(n12319), .A2(n13806), .ZN(n11405) );
  NAND2_X1 U13935 ( .A1(n11406), .A2(n11405), .ZN(n11407) );
  XNOR2_X1 U13936 ( .A(n11407), .B(n12315), .ZN(n11411) );
  NOR2_X1 U13937 ( .A1(n12317), .A2(n11408), .ZN(n11409) );
  AOI21_X1 U13938 ( .B1(n14717), .B2(n12312), .A(n11409), .ZN(n11410) );
  NAND2_X1 U13939 ( .A1(n11411), .A2(n11410), .ZN(n11552) );
  OAI21_X1 U13940 ( .B1(n11411), .B2(n11410), .A(n11552), .ZN(n11412) );
  AOI21_X1 U13941 ( .B1(n11413), .B2(n11412), .A(n6603), .ZN(n11421) );
  NAND2_X1 U13942 ( .A1(n14510), .A2(n13807), .ZN(n11415) );
  OAI211_X1 U13943 ( .C1(n11553), .C2(n13791), .A(n11415), .B(n11414), .ZN(
        n11418) );
  NOR2_X1 U13944 ( .A1(n14577), .A2(n11416), .ZN(n11417) );
  AOI211_X1 U13945 ( .C1(n13794), .C2(n11419), .A(n11418), .B(n11417), .ZN(
        n11420) );
  OAI21_X1 U13946 ( .B1(n11421), .B2(n14565), .A(n11420), .ZN(P1_U3221) );
  NAND2_X1 U13947 ( .A1(n11423), .A2(n11422), .ZN(n11425) );
  XOR2_X1 U13948 ( .A(n11425), .B(n11424), .Z(n11432) );
  NOR2_X1 U13949 ( .A1(n13097), .A2(n11451), .ZN(n11430) );
  NAND2_X1 U13950 ( .A1(n13131), .A2(n13061), .ZN(n11427) );
  NAND2_X1 U13951 ( .A1(n13134), .A2(n13050), .ZN(n11426) );
  AND2_X1 U13952 ( .A1(n11427), .A2(n11426), .ZN(n11448) );
  OAI21_X1 U13953 ( .B1(n13108), .B2(n11448), .A(n11428), .ZN(n11429) );
  AOI211_X1 U13954 ( .C1(n11953), .C2(n13081), .A(n11430), .B(n11429), .ZN(
        n11431) );
  OAI21_X1 U13955 ( .B1(n11432), .B2(n13070), .A(n11431), .ZN(P2_U3208) );
  XNOR2_X1 U13956 ( .A(n11434), .B(n11433), .ZN(n11435) );
  OAI222_X1 U13957 ( .A1(n15087), .A2(n11675), .B1(n15084), .B2(n11436), .C1(
        n15049), .C2(n11435), .ZN(n11564) );
  INV_X1 U13958 ( .A(n11564), .ZN(n11442) );
  OAI21_X1 U13959 ( .B1(n7546), .B2(n6961), .A(n11437), .ZN(n11565) );
  AOI22_X1 U13960 ( .A1(n15075), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n15071), 
        .B2(n11438), .ZN(n11439) );
  OAI21_X1 U13961 ( .B1(n12835), .B2(n11571), .A(n11439), .ZN(n11440) );
  AOI21_X1 U13962 ( .B1(n11565), .B2(n14445), .A(n11440), .ZN(n11441) );
  OAI21_X1 U13963 ( .B1(n11442), .B2(n15075), .A(n11441), .ZN(P3_U3222) );
  XNOR2_X1 U13964 ( .A(n11443), .B(n12120), .ZN(n14851) );
  INV_X1 U13965 ( .A(n14851), .ZN(n11456) );
  NAND2_X1 U13966 ( .A1(n11445), .A2(n11444), .ZN(n11446) );
  NAND2_X1 U13967 ( .A1(n11458), .A2(n11446), .ZN(n11447) );
  NAND2_X1 U13968 ( .A1(n11447), .A2(n13430), .ZN(n11449) );
  NAND2_X1 U13969 ( .A1(n11449), .A2(n11448), .ZN(n14856) );
  OAI211_X1 U13970 ( .C1(n11450), .C2(n14854), .A(n13372), .B(n11467), .ZN(
        n14852) );
  OAI22_X1 U13971 ( .A1(n13468), .A2(n10310), .B1(n11451), .B2(n13472), .ZN(
        n11452) );
  AOI21_X1 U13972 ( .B1(n11953), .B2(n13476), .A(n11452), .ZN(n11453) );
  OAI21_X1 U13973 ( .B1(n14852), .B2(n13350), .A(n11453), .ZN(n11454) );
  AOI21_X1 U13974 ( .B1(n14856), .B2(n13468), .A(n11454), .ZN(n11455) );
  OAI21_X1 U13975 ( .B1(n13467), .B2(n11456), .A(n11455), .ZN(P2_U3254) );
  XNOR2_X1 U13976 ( .A(n11457), .B(n12119), .ZN(n11518) );
  INV_X1 U13977 ( .A(n11518), .ZN(n11474) );
  INV_X1 U13978 ( .A(n11458), .ZN(n11460) );
  OAI21_X1 U13979 ( .B1(n11460), .B2(n11459), .A(n12119), .ZN(n11462) );
  NAND3_X1 U13980 ( .A1(n11462), .A2(n13430), .A3(n11461), .ZN(n11465) );
  NAND2_X1 U13981 ( .A1(n13130), .A2(n13061), .ZN(n11464) );
  NAND2_X1 U13982 ( .A1(n13133), .A2(n13050), .ZN(n11463) );
  AND2_X1 U13983 ( .A1(n11464), .A2(n11463), .ZN(n11576) );
  NAND2_X1 U13984 ( .A1(n11465), .A2(n11576), .ZN(n11513) );
  NAND2_X1 U13985 ( .A1(n11513), .A2(n13468), .ZN(n11473) );
  INV_X1 U13986 ( .A(n11602), .ZN(n11466) );
  AOI211_X1 U13987 ( .C1(n11961), .C2(n11467), .A(n13460), .B(n11466), .ZN(
        n11512) );
  INV_X1 U13988 ( .A(n11961), .ZN(n11468) );
  NOR2_X1 U13989 ( .A1(n11468), .A2(n13463), .ZN(n11471) );
  OAI22_X1 U13990 ( .A1(n13468), .A2(n11469), .B1(n11579), .B2(n13472), .ZN(
        n11470) );
  AOI211_X1 U13991 ( .C1(n11512), .C2(n13478), .A(n11471), .B(n11470), .ZN(
        n11472) );
  OAI211_X1 U13992 ( .C1(n11474), .C2(n13467), .A(n11473), .B(n11472), .ZN(
        P2_U3253) );
  INV_X1 U13993 ( .A(n14631), .ZN(n14056) );
  OAI21_X1 U13994 ( .B1(n11476), .B2(n11482), .A(n11589), .ZN(n11614) );
  OAI22_X1 U13995 ( .A1(n11833), .A2(n14622), .B1(n12206), .B2(n14583), .ZN(
        n11485) );
  INV_X1 U13996 ( .A(n11477), .ZN(n11478) );
  OR2_X1 U13997 ( .A1(n11835), .A2(n11833), .ZN(n11480) );
  NAND2_X1 U13998 ( .A1(n11481), .A2(n11480), .ZN(n11584) );
  INV_X1 U13999 ( .A(n11482), .ZN(n11583) );
  XNOR2_X1 U14000 ( .A(n11584), .B(n11583), .ZN(n11483) );
  NOR2_X1 U14001 ( .A1(n11483), .A2(n14621), .ZN(n11484) );
  AOI211_X1 U14002 ( .C1(n14056), .C2(n11614), .A(n11485), .B(n11484), .ZN(
        n11618) );
  INV_X1 U14003 ( .A(n11592), .ZN(n14337) );
  AOI211_X1 U14004 ( .C1(n11616), .C2(n11487), .A(n14058), .B(n14337), .ZN(
        n11615) );
  NAND2_X1 U14005 ( .A1(n11615), .A2(n14060), .ZN(n11489) );
  AOI22_X1 U14006 ( .A1(n14646), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7566), 
        .B2(n14636), .ZN(n11488) );
  OAI211_X1 U14007 ( .C1(n11851), .C2(n14640), .A(n11489), .B(n11488), .ZN(
        n11490) );
  AOI21_X1 U14008 ( .B1(n11614), .B2(n14066), .A(n11490), .ZN(n11491) );
  OAI21_X1 U14009 ( .B1(n11618), .B2(n14646), .A(n11491), .ZN(P1_U3281) );
  OAI222_X1 U14010 ( .A1(P1_U3086), .A2(n11492), .B1(n14204), .B2(n11857), 
        .C1(n15178), .C2(n14201), .ZN(P1_U3334) );
  INV_X1 U14011 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n13709) );
  NOR2_X1 U14012 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13709), .ZN(n11493) );
  AOI21_X1 U14013 ( .B1(n13852), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11493), 
        .ZN(n11494) );
  INV_X1 U14014 ( .A(n11494), .ZN(n11502) );
  NAND2_X1 U14015 ( .A1(n11496), .A2(n11495), .ZN(n11498) );
  NAND2_X1 U14016 ( .A1(n11498), .A2(n11497), .ZN(n11500) );
  XNOR2_X1 U14017 ( .A(n11700), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11499) );
  NOR2_X1 U14018 ( .A1(n11499), .A2(n11500), .ZN(n11699) );
  AOI211_X1 U14019 ( .C1(n11500), .C2(n11499), .A(n11699), .B(n11701), .ZN(
        n11501) );
  AOI211_X1 U14020 ( .C1(n13860), .C2(n11700), .A(n11502), .B(n11501), .ZN(
        n11511) );
  NOR2_X1 U14021 ( .A1(n11504), .A2(n11503), .ZN(n11506) );
  NOR2_X1 U14022 ( .A1(n11506), .A2(n11505), .ZN(n11509) );
  MUX2_X1 U14023 ( .A(n11737), .B(P1_REG2_REG_16__SCAN_IN), .S(n11700), .Z(
        n11507) );
  INV_X1 U14024 ( .A(n11507), .ZN(n11508) );
  NAND2_X1 U14025 ( .A1(n11508), .A2(n11509), .ZN(n11692) );
  OAI211_X1 U14026 ( .C1(n11509), .C2(n11508), .A(n13887), .B(n11692), .ZN(
        n11510) );
  NAND2_X1 U14027 ( .A1(n11511), .A2(n11510), .ZN(P1_U3259) );
  NOR2_X1 U14028 ( .A1(n11513), .A2(n11512), .ZN(n11521) );
  AOI22_X1 U14029 ( .A1(n11961), .A2(n13616), .B1(P2_REG0_REG_12__SCAN_IN), 
        .B2(n14858), .ZN(n11516) );
  NAND2_X1 U14030 ( .A1(n11518), .A2(n11514), .ZN(n11515) );
  OAI211_X1 U14031 ( .C1(n11521), .C2(n14858), .A(n11516), .B(n11515), .ZN(
        P2_U3466) );
  AOI22_X1 U14032 ( .A1(n11961), .A2(n13558), .B1(P2_REG1_REG_12__SCAN_IN), 
        .B2(n14862), .ZN(n11520) );
  NAND2_X1 U14033 ( .A1(n11518), .A2(n11517), .ZN(n11519) );
  OAI211_X1 U14034 ( .C1(n11521), .C2(n14862), .A(n11520), .B(n11519), .ZN(
        P2_U3511) );
  INV_X1 U14035 ( .A(n11522), .ZN(n11524) );
  OAI222_X1 U14036 ( .A1(P3_U3151), .A2(n11525), .B1(n12396), .B2(n11524), 
        .C1(n11523), .C2(n12962), .ZN(P3_U3270) );
  NAND2_X1 U14037 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n14817), .ZN(n11528) );
  INV_X1 U14038 ( .A(n11528), .ZN(n11526) );
  AOI21_X1 U14039 ( .B1(n13439), .B2(n11534), .A(n11526), .ZN(n14821) );
  OAI21_X1 U14040 ( .B1(n11533), .B2(n13462), .A(n11527), .ZN(n14822) );
  NAND2_X1 U14041 ( .A1(n14821), .A2(n14822), .ZN(n14819) );
  NAND2_X1 U14042 ( .A1(n11528), .A2(n14819), .ZN(n13236) );
  XNOR2_X1 U14043 ( .A(n13241), .B(n13236), .ZN(n11529) );
  NOR2_X1 U14044 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n11529), .ZN(n13238) );
  AOI21_X1 U14045 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n11529), .A(n13238), 
        .ZN(n11540) );
  NAND2_X1 U14046 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3088), .ZN(n11530)
         );
  OAI21_X1 U14047 ( .B1(n14769), .B2(n11531), .A(n11530), .ZN(n11538) );
  INV_X1 U14048 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13547) );
  XNOR2_X1 U14049 ( .A(n14817), .B(n13547), .ZN(n14815) );
  OAI21_X1 U14050 ( .B1(n11533), .B2(n13553), .A(n11532), .ZN(n14816) );
  NAND2_X1 U14051 ( .A1(n14815), .A2(n14816), .ZN(n14813) );
  OAI21_X1 U14052 ( .B1(n11534), .B2(n13547), .A(n14813), .ZN(n13240) );
  XOR2_X1 U14053 ( .A(n13241), .B(n13240), .Z(n11535) );
  NAND2_X1 U14054 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n11535), .ZN(n13243) );
  OAI21_X1 U14055 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n11535), .A(n13243), 
        .ZN(n11536) );
  NOR2_X1 U14056 ( .A1(n11536), .A2(n14750), .ZN(n11537) );
  AOI211_X1 U14057 ( .C1(n14812), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n11538), 
        .B(n11537), .ZN(n11539) );
  OAI21_X1 U14058 ( .B1(n11540), .B2(n14751), .A(n11539), .ZN(P2_U3232) );
  INV_X1 U14059 ( .A(n11543), .ZN(n11544) );
  XOR2_X1 U14060 ( .A(n10487), .B(n14457), .Z(n11638) );
  XNOR2_X1 U14061 ( .A(n11638), .B(n14438), .ZN(n11545) );
  XNOR2_X1 U14062 ( .A(n11640), .B(n11545), .ZN(n11551) );
  INV_X1 U14063 ( .A(n14457), .ZN(n11678) );
  INV_X1 U14064 ( .A(n11546), .ZN(n11676) );
  AND2_X1 U14065 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n15010) );
  NOR2_X1 U14066 ( .A1(n12516), .A2(n11751), .ZN(n11547) );
  AOI211_X1 U14067 ( .C1(n12530), .C2(n12548), .A(n15010), .B(n11547), .ZN(
        n11548) );
  OAI21_X1 U14068 ( .B1(n11676), .B2(n12532), .A(n11548), .ZN(n11549) );
  AOI21_X1 U14069 ( .B1(n11678), .B2(n12521), .A(n11549), .ZN(n11550) );
  OAI21_X1 U14070 ( .B1(n11551), .B2(n12523), .A(n11550), .ZN(P3_U3174) );
  NOR2_X1 U14071 ( .A1(n12317), .A2(n11553), .ZN(n11554) );
  AOI21_X1 U14072 ( .B1(n14739), .B2(n12319), .A(n11554), .ZN(n11822) );
  AOI22_X1 U14073 ( .A1(n14739), .A2(n12333), .B1(n12319), .B2(n13805), .ZN(
        n11555) );
  XNOR2_X1 U14074 ( .A(n11555), .B(n12334), .ZN(n11823) );
  XNOR2_X1 U14075 ( .A(n11824), .B(n11823), .ZN(n11563) );
  NAND2_X1 U14076 ( .A1(n14510), .A2(n13806), .ZN(n11558) );
  INV_X1 U14077 ( .A(n11556), .ZN(n11557) );
  OAI211_X1 U14078 ( .C1(n11828), .C2(n13791), .A(n11558), .B(n11557), .ZN(
        n11560) );
  NOR2_X1 U14079 ( .A1(n14577), .A2(n6900), .ZN(n11559) );
  AOI211_X1 U14080 ( .C1(n13794), .C2(n11561), .A(n11560), .B(n11559), .ZN(
        n11562) );
  OAI21_X1 U14081 ( .B1(n11563), .B2(n14565), .A(n11562), .ZN(P1_U3231) );
  INV_X1 U14082 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n11566) );
  AOI21_X1 U14083 ( .B1(n15101), .B2(n11565), .A(n11564), .ZN(n11568) );
  MUX2_X1 U14084 ( .A(n11566), .B(n11568), .S(n15157), .Z(n11567) );
  OAI21_X1 U14085 ( .B1(n11571), .B2(n12894), .A(n11567), .ZN(P3_U3470) );
  INV_X1 U14086 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n11569) );
  MUX2_X1 U14087 ( .A(n11569), .B(n11568), .S(n15141), .Z(n11570) );
  OAI21_X1 U14088 ( .B1(n11571), .B2(n12939), .A(n11570), .ZN(P3_U3423) );
  INV_X1 U14089 ( .A(n11572), .ZN(n11573) );
  AOI21_X1 U14090 ( .B1(n11575), .B2(n11574), .A(n11573), .ZN(n11582) );
  INV_X1 U14091 ( .A(n11576), .ZN(n11577) );
  AOI22_X1 U14092 ( .A1(n13099), .A2(n11577), .B1(P2_REG3_REG_12__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11578) );
  OAI21_X1 U14093 ( .B1(n11579), .B2(n13097), .A(n11578), .ZN(n11580) );
  AOI21_X1 U14094 ( .B1(n11961), .B2(n13081), .A(n11580), .ZN(n11581) );
  OAI21_X1 U14095 ( .B1(n11582), .B2(n13070), .A(n11581), .ZN(P2_U3196) );
  OR2_X1 U14096 ( .A1(n11616), .A2(n11843), .ZN(n11585) );
  INV_X1 U14097 ( .A(n14347), .ZN(n14349) );
  XNOR2_X1 U14098 ( .A(n11624), .B(n11627), .ZN(n11587) );
  OAI222_X1 U14099 ( .A1(n14583), .A2(n12226), .B1(n11587), .B2(n14621), .C1(
        n14622), .C2(n12206), .ZN(n14521) );
  INV_X1 U14100 ( .A(n14521), .ZN(n11600) );
  OR2_X1 U14101 ( .A1(n11616), .A2(n14511), .ZN(n11588) );
  OR2_X1 U14102 ( .A1(n14343), .A2(n14483), .ZN(n11590) );
  XNOR2_X1 U14103 ( .A(n11628), .B(n11591), .ZN(n14523) );
  AOI21_X1 U14104 ( .B1(n12214), .B2(n14336), .A(n14058), .ZN(n11593) );
  NAND2_X1 U14105 ( .A1(n11593), .A2(n6599), .ZN(n14519) );
  OAI22_X1 U14106 ( .A1(n11595), .A2(n11594), .B1(n14490), .B2(n14608), .ZN(
        n11596) );
  AOI21_X1 U14107 ( .B1(n12214), .B2(n14613), .A(n11596), .ZN(n11597) );
  OAI21_X1 U14108 ( .B1(n14519), .B2(n14639), .A(n11597), .ZN(n11598) );
  AOI21_X1 U14109 ( .B1(n14523), .B2(n14618), .A(n11598), .ZN(n11599) );
  OAI21_X1 U14110 ( .B1(n11600), .B2(n14646), .A(n11599), .ZN(P1_U3279) );
  XOR2_X1 U14111 ( .A(n12122), .B(n11601), .Z(n11796) );
  AOI211_X1 U14112 ( .C1(n11969), .C2(n11602), .A(n13460), .B(n11684), .ZN(
        n11780) );
  INV_X1 U14113 ( .A(n11969), .ZN(n11668) );
  NOR2_X1 U14114 ( .A1(n11668), .A2(n13463), .ZN(n11605) );
  OAI22_X1 U14115 ( .A1(n13468), .A2(n11603), .B1(n11662), .B2(n13472), .ZN(
        n11604) );
  AOI211_X1 U14116 ( .C1(n11780), .C2(n13478), .A(n11605), .B(n11604), .ZN(
        n11613) );
  OAI211_X1 U14117 ( .C1(n11607), .C2(n12122), .A(n11606), .B(n13430), .ZN(
        n11611) );
  OR2_X1 U14118 ( .A1(n11967), .A2(n13094), .ZN(n11609) );
  NAND2_X1 U14119 ( .A1(n13131), .A2(n13050), .ZN(n11608) );
  NAND2_X1 U14120 ( .A1(n11609), .A2(n11608), .ZN(n11665) );
  INV_X1 U14121 ( .A(n11665), .ZN(n11610) );
  NAND2_X1 U14122 ( .A1(n11611), .A2(n11610), .ZN(n11779) );
  NAND2_X1 U14123 ( .A1(n11779), .A2(n13468), .ZN(n11612) );
  OAI211_X1 U14124 ( .C1(n11796), .C2(n13467), .A(n11613), .B(n11612), .ZN(
        P2_U3252) );
  INV_X1 U14125 ( .A(n11614), .ZN(n11619) );
  AOI21_X1 U14126 ( .B1(n14740), .B2(n11616), .A(n11615), .ZN(n11617) );
  OAI211_X1 U14127 ( .C1(n11619), .C2(n14743), .A(n11618), .B(n11617), .ZN(
        n11622) );
  NAND2_X1 U14128 ( .A1(n11622), .A2(n14748), .ZN(n11620) );
  OAI21_X1 U14129 ( .B1(n14748), .B2(n11621), .A(n11620), .ZN(P1_U3540) );
  NAND2_X1 U14130 ( .A1(n11622), .A2(n15160), .ZN(n11623) );
  OAI21_X1 U14131 ( .B1(n15160), .B2(n8522), .A(n11623), .ZN(P1_U3495) );
  XNOR2_X1 U14132 ( .A(n11720), .B(n11719), .ZN(n14167) );
  NAND2_X1 U14133 ( .A1(n12214), .A2(n14338), .ZN(n11626) );
  XNOR2_X1 U14134 ( .A(n11726), .B(n11719), .ZN(n14165) );
  NAND2_X1 U14135 ( .A1(n14165), .A2(n14618), .ZN(n11636) );
  NAND2_X1 U14136 ( .A1(n12222), .A2(n6599), .ZN(n11629) );
  NAND2_X1 U14137 ( .A1(n11629), .A2(n14637), .ZN(n11630) );
  NOR2_X1 U14138 ( .A1(n11732), .A2(n11630), .ZN(n14164) );
  INV_X1 U14139 ( .A(n12222), .ZN(n14162) );
  AOI22_X1 U14140 ( .A1(n14339), .A2(n14338), .B1(n13803), .B2(n14050), .ZN(
        n14161) );
  OAI22_X1 U14141 ( .A1(n14646), .A2(n14161), .B1(n11631), .B2(n14608), .ZN(
        n11632) );
  AOI21_X1 U14142 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14646), .A(n11632), 
        .ZN(n11633) );
  OAI21_X1 U14143 ( .B1(n14162), .B2(n14640), .A(n11633), .ZN(n11634) );
  AOI21_X1 U14144 ( .B1(n14164), .B2(n14060), .A(n11634), .ZN(n11635) );
  OAI211_X1 U14145 ( .C1(n14167), .C2(n14351), .A(n11636), .B(n11635), .ZN(
        P1_U3278) );
  NAND2_X1 U14146 ( .A1(n11638), .A2(n11637), .ZN(n11639) );
  XNOR2_X1 U14147 ( .A(n14456), .B(n10487), .ZN(n11711) );
  XNOR2_X1 U14148 ( .A(n11711), .B(n11751), .ZN(n11712) );
  XNOR2_X1 U14149 ( .A(n11713), .B(n11712), .ZN(n11647) );
  INV_X1 U14150 ( .A(n11641), .ZN(n11654) );
  NOR2_X1 U14151 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11642), .ZN(n15029) );
  NOR2_X1 U14152 ( .A1(n12516), .A2(n12828), .ZN(n11643) );
  AOI211_X1 U14153 ( .C1(n12530), .C2(n14438), .A(n15029), .B(n11643), .ZN(
        n11644) );
  OAI21_X1 U14154 ( .B1(n11654), .B2(n12532), .A(n11644), .ZN(n11645) );
  AOI21_X1 U14155 ( .B1(n14456), .B2(n12521), .A(n11645), .ZN(n11646) );
  OAI21_X1 U14156 ( .B1(n11647), .B2(n12523), .A(n11646), .ZN(P3_U3155) );
  XOR2_X1 U14157 ( .A(n11650), .B(n11648), .Z(n14453) );
  OAI211_X1 U14158 ( .C1(n11651), .C2(n11650), .A(n11649), .B(n15089), .ZN(
        n11653) );
  AOI22_X1 U14159 ( .A1(n12547), .A2(n14437), .B1(n14435), .B2(n14438), .ZN(
        n11652) );
  NAND2_X1 U14160 ( .A1(n11653), .A2(n11652), .ZN(n14454) );
  NAND2_X1 U14161 ( .A1(n14454), .A2(n15096), .ZN(n11658) );
  INV_X1 U14162 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n11655) );
  OAI22_X1 U14163 ( .A1(n15096), .A2(n11655), .B1(n11654), .B2(n15081), .ZN(
        n11656) );
  AOI21_X1 U14164 ( .B1(n14456), .B2(n12801), .A(n11656), .ZN(n11657) );
  OAI211_X1 U14165 ( .C1(n14453), .C2(n12805), .A(n11658), .B(n11657), .ZN(
        P3_U3219) );
  AOI21_X1 U14166 ( .B1(n11660), .B2(n11659), .A(n13070), .ZN(n11661) );
  NAND2_X1 U14167 ( .A1(n11661), .A2(n6592), .ZN(n11667) );
  NOR2_X1 U14168 ( .A1(n13097), .A2(n11662), .ZN(n11663) );
  AOI211_X1 U14169 ( .C1(n13099), .C2(n11665), .A(n11664), .B(n11663), .ZN(
        n11666) );
  OAI211_X1 U14170 ( .C1(n11668), .C2(n13114), .A(n11667), .B(n11666), .ZN(
        P2_U3206) );
  XOR2_X1 U14171 ( .A(n11669), .B(n11673), .Z(n14459) );
  INV_X1 U14172 ( .A(n11671), .ZN(n11672) );
  AOI21_X1 U14173 ( .B1(n11673), .B2(n11670), .A(n11672), .ZN(n11674) );
  OAI222_X1 U14174 ( .A1(n15087), .A2(n11751), .B1(n15084), .B2(n11675), .C1(
        n15049), .C2(n11674), .ZN(n14461) );
  NAND2_X1 U14175 ( .A1(n14461), .A2(n15096), .ZN(n11680) );
  INV_X1 U14176 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n15242) );
  OAI22_X1 U14177 ( .A1(n15096), .A2(n15242), .B1(n11676), .B2(n15081), .ZN(
        n11677) );
  AOI21_X1 U14178 ( .B1(n11678), .B2(n12801), .A(n11677), .ZN(n11679) );
  OAI211_X1 U14179 ( .C1(n12805), .C2(n14459), .A(n11680), .B(n11679), .ZN(
        P3_U3220) );
  XNOR2_X1 U14180 ( .A(n11966), .B(n13129), .ZN(n12125) );
  XNOR2_X1 U14181 ( .A(n11681), .B(n12125), .ZN(n11682) );
  AOI22_X1 U14182 ( .A1(n13128), .A2(n13061), .B1(n13130), .B2(n13050), .ZN(
        n11788) );
  OAI21_X1 U14183 ( .B1(n11682), .B2(n13454), .A(n11788), .ZN(n11760) );
  INV_X1 U14184 ( .A(n11760), .ZN(n11691) );
  XNOR2_X1 U14185 ( .A(n11683), .B(n12125), .ZN(n11762) );
  INV_X1 U14186 ( .A(n11684), .ZN(n11686) );
  INV_X1 U14187 ( .A(n11773), .ZN(n11685) );
  AOI211_X1 U14188 ( .C1(n11966), .C2(n11686), .A(n13460), .B(n11685), .ZN(
        n11761) );
  NAND2_X1 U14189 ( .A1(n11761), .A2(n13478), .ZN(n11688) );
  AOI22_X1 U14190 ( .A1(n13428), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11790), 
        .B2(n13419), .ZN(n11687) );
  OAI211_X1 U14191 ( .C1(n11968), .C2(n13463), .A(n11688), .B(n11687), .ZN(
        n11689) );
  AOI21_X1 U14192 ( .B1(n11762), .B2(n13470), .A(n11689), .ZN(n11690) );
  OAI21_X1 U14193 ( .B1(n11691), .B2(n13428), .A(n11690), .ZN(P2_U3251) );
  NAND2_X1 U14194 ( .A1(n11700), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11693) );
  NAND2_X1 U14195 ( .A1(n11693), .A2(n11692), .ZN(n11695) );
  XNOR2_X1 U14196 ( .A(n13867), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n11694) );
  NAND2_X1 U14197 ( .A1(n11694), .A2(n11695), .ZN(n13866) );
  OAI211_X1 U14198 ( .C1(n11695), .C2(n11694), .A(n13887), .B(n13866), .ZN(
        n11707) );
  INV_X1 U14199 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n11698) );
  NOR2_X1 U14200 ( .A1(n11696), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13719) );
  INV_X1 U14201 ( .A(n13719), .ZN(n11697) );
  OAI21_X1 U14202 ( .B1(n14605), .B2(n11698), .A(n11697), .ZN(n11705) );
  XNOR2_X1 U14203 ( .A(n13862), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n11702) );
  AOI211_X1 U14204 ( .C1(n11703), .C2(n11702), .A(n13861), .B(n11701), .ZN(
        n11704) );
  AOI211_X1 U14205 ( .C1(n13860), .C2(n13862), .A(n11705), .B(n11704), .ZN(
        n11706) );
  NAND2_X1 U14206 ( .A1(n11707), .A2(n11706), .ZN(P1_U3260) );
  INV_X1 U14207 ( .A(n11708), .ZN(n11710) );
  OAI222_X1 U14208 ( .A1(n13651), .A2(n11710), .B1(n12089), .B2(P2_U3088), 
        .C1(n11709), .C2(n13624), .ZN(P2_U3305) );
  XNOR2_X1 U14209 ( .A(n11754), .B(n10487), .ZN(n11797) );
  XNOR2_X1 U14210 ( .A(n11797), .B(n12547), .ZN(n11799) );
  XNOR2_X1 U14211 ( .A(n11800), .B(n11799), .ZN(n11718) );
  NAND2_X1 U14212 ( .A1(n12505), .A2(n11755), .ZN(n11715) );
  AND2_X1 U14213 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n14374) );
  AOI21_X1 U14214 ( .B1(n12535), .B2(n12546), .A(n14374), .ZN(n11714) );
  OAI211_X1 U14215 ( .C1(n11751), .C2(n12508), .A(n11715), .B(n11714), .ZN(
        n11716) );
  AOI21_X1 U14216 ( .B1(n11754), .B2(n12521), .A(n11716), .ZN(n11717) );
  OAI21_X1 U14217 ( .B1(n11718), .B2(n12523), .A(n11717), .ZN(P3_U3181) );
  NAND2_X1 U14218 ( .A1(n11720), .A2(n11719), .ZN(n11722) );
  NAND2_X1 U14219 ( .A1(n11722), .A2(n11721), .ZN(n11725) );
  INV_X1 U14220 ( .A(n11725), .ZN(n11724) );
  INV_X1 U14221 ( .A(n11730), .ZN(n11723) );
  INV_X1 U14222 ( .A(n11812), .ZN(n11808) );
  AOI21_X1 U14223 ( .B1(n11730), .B2(n11725), .A(n11808), .ZN(n14160) );
  INV_X1 U14224 ( .A(n12226), .ZN(n14484) );
  OR2_X1 U14225 ( .A1(n12222), .A2(n14484), .ZN(n11728) );
  OAI21_X1 U14226 ( .B1(n11731), .B2(n11730), .A(n11807), .ZN(n14158) );
  INV_X1 U14227 ( .A(n12232), .ZN(n14156) );
  OAI211_X1 U14228 ( .C1(n14156), .C2(n11732), .A(n14637), .B(n11816), .ZN(
        n14155) );
  NAND2_X1 U14229 ( .A1(n14052), .A2(n14050), .ZN(n11734) );
  NAND2_X1 U14230 ( .A1(n14484), .A2(n14339), .ZN(n11733) );
  AND2_X1 U14231 ( .A1(n11734), .A2(n11733), .ZN(n14154) );
  INV_X1 U14232 ( .A(n14154), .ZN(n11735) );
  AOI22_X1 U14233 ( .A1(n14610), .A2(n11735), .B1(n13712), .B2(n14636), .ZN(
        n11736) );
  OAI21_X1 U14234 ( .B1(n11737), .B2(n14610), .A(n11736), .ZN(n11738) );
  AOI21_X1 U14235 ( .B1(n12232), .B2(n14613), .A(n11738), .ZN(n11739) );
  OAI21_X1 U14236 ( .B1(n14155), .B2(n14639), .A(n11739), .ZN(n11740) );
  AOI21_X1 U14237 ( .B1(n14158), .B2(n14618), .A(n11740), .ZN(n11741) );
  OAI21_X1 U14238 ( .B1(n14160), .B2(n14351), .A(n11741), .ZN(P1_U3277) );
  OR2_X1 U14239 ( .A1(n11742), .A2(P2_U3088), .ZN(n12148) );
  INV_X1 U14240 ( .A(n12148), .ZN(n12142) );
  AOI21_X1 U14241 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n11743), .A(n12142), 
        .ZN(n11744) );
  OAI21_X1 U14242 ( .B1(n11747), .B2(n13645), .A(n11744), .ZN(P2_U3304) );
  NAND2_X1 U14243 ( .A1(n14188), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11745) );
  OAI211_X1 U14244 ( .C1(n11747), .C2(n14204), .A(n11746), .B(n11745), .ZN(
        P1_U3332) );
  XNOR2_X1 U14245 ( .A(n11749), .B(n11748), .ZN(n11750) );
  OAI222_X1 U14246 ( .A1(n15087), .A2(n12812), .B1(n15084), .B2(n11751), .C1(
        n11750), .C2(n15049), .ZN(n12890) );
  INV_X1 U14247 ( .A(n12890), .ZN(n11759) );
  XNOR2_X1 U14248 ( .A(n11753), .B(n11752), .ZN(n12891) );
  INV_X1 U14249 ( .A(n11754), .ZN(n12940) );
  AOI22_X1 U14250 ( .A1(n15075), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15071), 
        .B2(n11755), .ZN(n11756) );
  OAI21_X1 U14251 ( .B1(n12940), .B2(n12835), .A(n11756), .ZN(n11757) );
  AOI21_X1 U14252 ( .B1(n12891), .B2(n14445), .A(n11757), .ZN(n11758) );
  OAI21_X1 U14253 ( .B1(n11759), .B2(n15075), .A(n11758), .ZN(P3_U3218) );
  AOI211_X1 U14254 ( .C1(n14850), .C2(n11762), .A(n11761), .B(n11760), .ZN(
        n11765) );
  AOI22_X1 U14255 ( .A1(n11966), .A2(n13558), .B1(P2_REG1_REG_14__SCAN_IN), 
        .B2(n14862), .ZN(n11763) );
  OAI21_X1 U14256 ( .B1(n11765), .B2(n14862), .A(n11763), .ZN(P2_U3513) );
  AOI22_X1 U14257 ( .A1(n11966), .A2(n13616), .B1(P2_REG0_REG_14__SCAN_IN), 
        .B2(n14858), .ZN(n11764) );
  OAI21_X1 U14258 ( .B1(n11765), .B2(n14858), .A(n11764), .ZN(P2_U3472) );
  XOR2_X1 U14259 ( .A(n11766), .B(n12124), .Z(n13621) );
  INV_X1 U14260 ( .A(n11767), .ZN(n11768) );
  AOI21_X1 U14261 ( .B1(n12124), .B2(n11769), .A(n11768), .ZN(n11772) );
  OR2_X1 U14262 ( .A1(n11967), .A2(n13092), .ZN(n11771) );
  NAND2_X1 U14263 ( .A1(n13127), .A2(n13061), .ZN(n11770) );
  AND2_X1 U14264 ( .A1(n11771), .A2(n11770), .ZN(n13107) );
  OAI21_X1 U14265 ( .B1(n11772), .B2(n13454), .A(n13107), .ZN(n13556) );
  INV_X1 U14266 ( .A(n13617), .ZN(n13115) );
  AOI211_X1 U14267 ( .C1(n13617), .C2(n11773), .A(n13460), .B(n7108), .ZN(
        n13555) );
  NAND2_X1 U14268 ( .A1(n13555), .A2(n13478), .ZN(n11776) );
  INV_X1 U14269 ( .A(n11774), .ZN(n13111) );
  AOI22_X1 U14270 ( .A1(n13428), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n13111), 
        .B2(n13419), .ZN(n11775) );
  OAI211_X1 U14271 ( .C1(n13115), .C2(n13463), .A(n11776), .B(n11775), .ZN(
        n11777) );
  AOI21_X1 U14272 ( .B1(n13556), .B2(n13468), .A(n11777), .ZN(n11778) );
  OAI21_X1 U14273 ( .B1(n13467), .B2(n13621), .A(n11778), .ZN(P2_U3250) );
  AOI211_X1 U14274 ( .C1(n14845), .C2(n11969), .A(n11780), .B(n11779), .ZN(
        n11793) );
  NOR2_X1 U14275 ( .A1(n11793), .A2(n14862), .ZN(n11781) );
  AOI21_X1 U14276 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n14862), .A(n11781), 
        .ZN(n11782) );
  OAI21_X1 U14277 ( .B1(n13561), .B2(n11796), .A(n11782), .ZN(P2_U3512) );
  OAI21_X1 U14278 ( .B1(n11785), .B2(n11784), .A(n11783), .ZN(n11786) );
  NAND2_X1 U14279 ( .A1(n11786), .A2(n9789), .ZN(n11792) );
  OAI22_X1 U14280 ( .A1(n13108), .A2(n11788), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11787), .ZN(n11789) );
  AOI21_X1 U14281 ( .B1(n11790), .B2(n13110), .A(n11789), .ZN(n11791) );
  OAI211_X1 U14282 ( .C1(n11968), .C2(n13114), .A(n11792), .B(n11791), .ZN(
        P2_U3187) );
  NOR2_X1 U14283 ( .A1(n11793), .A2(n14858), .ZN(n11794) );
  AOI21_X1 U14284 ( .B1(P2_REG0_REG_13__SCAN_IN), .B2(n14858), .A(n11794), 
        .ZN(n11795) );
  OAI21_X1 U14285 ( .B1(n13620), .B2(n11796), .A(n11795), .ZN(P2_U3469) );
  INV_X1 U14286 ( .A(n11797), .ZN(n11798) );
  XNOR2_X1 U14287 ( .A(n12832), .B(n10487), .ZN(n12157) );
  XNOR2_X1 U14288 ( .A(n12157), .B(n12812), .ZN(n12159) );
  XNOR2_X1 U14289 ( .A(n12160), .B(n12159), .ZN(n11805) );
  NAND2_X1 U14290 ( .A1(n12505), .A2(n12833), .ZN(n11802) );
  INV_X1 U14291 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n15303) );
  NOR2_X1 U14292 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15303), .ZN(n14391) );
  AOI21_X1 U14293 ( .B1(n12535), .B2(n12545), .A(n14391), .ZN(n11801) );
  OAI211_X1 U14294 ( .C1(n12828), .C2(n12508), .A(n11802), .B(n11801), .ZN(
        n11803) );
  AOI21_X1 U14295 ( .B1(n12832), .B2(n12521), .A(n11803), .ZN(n11804) );
  OAI21_X1 U14296 ( .B1(n11805), .B2(n12523), .A(n11804), .ZN(P3_U3166) );
  OR2_X1 U14297 ( .A1(n12232), .A2(n13803), .ZN(n11806) );
  XOR2_X1 U14298 ( .A(n12346), .B(n11810), .Z(n14152) );
  AND2_X1 U14299 ( .A1(n12232), .A2(n13792), .ZN(n11809) );
  OAI21_X1 U14300 ( .B1(n11808), .B2(n11809), .A(n11810), .ZN(n11813) );
  NOR2_X1 U14301 ( .A1(n11810), .A2(n11809), .ZN(n11811) );
  NAND3_X1 U14302 ( .A1(n11813), .A2(n12363), .A3(n14138), .ZN(n11815) );
  AOI22_X1 U14303 ( .A1(n14050), .A2(n14038), .B1(n13803), .B2(n14339), .ZN(
        n11814) );
  NAND2_X1 U14304 ( .A1(n11815), .A2(n11814), .ZN(n14148) );
  AOI211_X1 U14305 ( .C1(n14150), .C2(n11816), .A(n14058), .B(n7224), .ZN(
        n14149) );
  NAND2_X1 U14306 ( .A1(n14149), .A2(n13991), .ZN(n11818) );
  AOI22_X1 U14307 ( .A1(n14646), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n13720), 
        .B2(n14636), .ZN(n11817) );
  OAI211_X1 U14308 ( .C1(n11819), .C2(n14640), .A(n11818), .B(n11817), .ZN(
        n11820) );
  AOI21_X1 U14309 ( .B1(n14148), .B2(n14610), .A(n11820), .ZN(n11821) );
  OAI21_X1 U14310 ( .B1(n14152), .B2(n14352), .A(n11821), .ZN(P1_U3276) );
  NAND2_X1 U14311 ( .A1(n14491), .A2(n12333), .ZN(n11826) );
  NAND2_X1 U14312 ( .A1(n14509), .A2(n12312), .ZN(n11825) );
  NAND2_X1 U14313 ( .A1(n11826), .A2(n11825), .ZN(n11827) );
  XNOR2_X1 U14314 ( .A(n11827), .B(n12315), .ZN(n11837) );
  NOR2_X1 U14315 ( .A1(n12317), .A2(n11828), .ZN(n11829) );
  AOI21_X1 U14316 ( .B1(n14491), .B2(n12312), .A(n11829), .ZN(n11836) );
  NAND2_X1 U14317 ( .A1(n11837), .A2(n11836), .ZN(n14494) );
  NAND2_X1 U14318 ( .A1(n11835), .A2(n12333), .ZN(n11831) );
  NAND2_X1 U14319 ( .A1(n13804), .A2(n12312), .ZN(n11830) );
  NAND2_X1 U14320 ( .A1(n11831), .A2(n11830), .ZN(n11832) );
  XNOR2_X1 U14321 ( .A(n11832), .B(n12334), .ZN(n11839) );
  NOR2_X1 U14322 ( .A1(n12317), .A2(n11833), .ZN(n11834) );
  AOI21_X1 U14323 ( .B1(n11835), .B2(n12319), .A(n11834), .ZN(n11840) );
  XNOR2_X1 U14324 ( .A(n11839), .B(n11840), .ZN(n14504) );
  OR2_X1 U14325 ( .A1(n11837), .A2(n11836), .ZN(n14505) );
  AND2_X1 U14326 ( .A1(n14504), .A2(n14505), .ZN(n11838) );
  INV_X1 U14327 ( .A(n11839), .ZN(n11841) );
  OAI22_X1 U14328 ( .A1(n11851), .A2(n12274), .B1(n11843), .B2(n12317), .ZN(
        n12204) );
  OAI22_X1 U14329 ( .A1(n11851), .A2(n11842), .B1(n11843), .B2(n12274), .ZN(
        n11844) );
  XNOR2_X1 U14330 ( .A(n11844), .B(n12334), .ZN(n12203) );
  XOR2_X1 U14331 ( .A(n12204), .B(n12203), .Z(n11845) );
  OAI211_X1 U14332 ( .C1(n11846), .C2(n11845), .A(n12205), .B(n14580), .ZN(
        n11850) );
  NAND2_X1 U14333 ( .A1(n14510), .A2(n13804), .ZN(n11847) );
  NAND2_X1 U14334 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n14603)
         );
  OAI211_X1 U14335 ( .C1(n12206), .C2(n13791), .A(n11847), .B(n14603), .ZN(
        n11848) );
  AOI21_X1 U14336 ( .B1(n7566), .B2(n13794), .A(n11848), .ZN(n11849) );
  OAI211_X1 U14337 ( .C1(n11851), .C2(n14577), .A(n11850), .B(n11849), .ZN(
        P1_U3224) );
  INV_X1 U14338 ( .A(n11852), .ZN(n11853) );
  NAND2_X1 U14339 ( .A1(n12539), .A2(n11853), .ZN(n14448) );
  NAND2_X1 U14340 ( .A1(n11854), .A2(n15071), .ZN(n12424) );
  OAI21_X1 U14341 ( .B1(n15075), .B2(n14448), .A(n12424), .ZN(n12662) );
  AOI21_X1 U14342 ( .B1(n15075), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12662), 
        .ZN(n11855) );
  OAI21_X1 U14343 ( .B1(n9486), .B2(n12835), .A(n11855), .ZN(P3_U3202) );
  OAI222_X1 U14344 ( .A1(n13651), .A2(n11857), .B1(n12138), .B2(P2_U3088), 
        .C1(n11856), .C2(n13650), .ZN(P2_U3306) );
  INV_X1 U14345 ( .A(n11858), .ZN(n13647) );
  OAI222_X1 U14346 ( .A1(P1_U3086), .A2(n10221), .B1(n14204), .B2(n13647), 
        .C1(n14201), .C2(n11859), .ZN(P1_U3330) );
  INV_X2 U14347 ( .A(n11863), .ZN(n12085) );
  OAI22_X1 U14348 ( .A1(n13320), .A2(n11863), .B1(n12085), .B2(n13093), .ZN(
        n12041) );
  OAI22_X1 U14349 ( .A1(n13422), .A2(n11863), .B1(n12085), .B2(n13028), .ZN(
        n12013) );
  INV_X1 U14350 ( .A(n12013), .ZN(n12017) );
  INV_X1 U14351 ( .A(n13143), .ZN(n11861) );
  NAND2_X1 U14352 ( .A1(n11860), .A2(n12090), .ZN(n11864) );
  NAND2_X1 U14353 ( .A1(n11861), .A2(n7568), .ZN(n11868) );
  NAND2_X1 U14354 ( .A1(n11862), .A2(n12059), .ZN(n11867) );
  OAI211_X1 U14355 ( .C1(n11865), .C2(n11864), .A(n13143), .B(n11863), .ZN(
        n11866) );
  NAND3_X1 U14356 ( .A1(n11868), .A2(n11867), .A3(n11866), .ZN(n11876) );
  NAND2_X1 U14357 ( .A1(n11872), .A2(n12059), .ZN(n11871) );
  NAND2_X1 U14358 ( .A1(n11869), .A2(n11863), .ZN(n11870) );
  NAND2_X1 U14359 ( .A1(n11872), .A2(n11863), .ZN(n11873) );
  OAI21_X1 U14360 ( .B1(n11874), .B2(n11863), .A(n11873), .ZN(n11875) );
  OAI21_X1 U14361 ( .B1(n11876), .B2(n11877), .A(n11875), .ZN(n11879) );
  NAND2_X1 U14362 ( .A1(n11877), .A2(n11876), .ZN(n11878) );
  NAND2_X1 U14363 ( .A1(n11879), .A2(n11878), .ZN(n11885) );
  NAND2_X1 U14364 ( .A1(n13142), .A2(n11863), .ZN(n11881) );
  NAND2_X1 U14365 ( .A1(n14837), .A2(n12066), .ZN(n11880) );
  NAND2_X1 U14366 ( .A1(n13142), .A2(n12066), .ZN(n11882) );
  OAI21_X1 U14367 ( .B1(n12059), .B2(n11883), .A(n11882), .ZN(n11884) );
  NAND2_X1 U14368 ( .A1(n13141), .A2(n12059), .ZN(n11887) );
  NAND2_X1 U14369 ( .A1(n6828), .A2(n11863), .ZN(n11886) );
  NAND2_X1 U14370 ( .A1(n11887), .A2(n11886), .ZN(n11893) );
  NAND2_X1 U14371 ( .A1(n13141), .A2(n11863), .ZN(n11888) );
  OAI21_X1 U14372 ( .B1(n11889), .B2(n11863), .A(n11888), .ZN(n11890) );
  NAND2_X1 U14373 ( .A1(n11891), .A2(n11890), .ZN(n11897) );
  INV_X1 U14374 ( .A(n11892), .ZN(n11895) );
  INV_X1 U14375 ( .A(n11893), .ZN(n11894) );
  NAND2_X1 U14376 ( .A1(n11895), .A2(n11894), .ZN(n11896) );
  NAND2_X1 U14377 ( .A1(n13140), .A2(n11863), .ZN(n11899) );
  NAND2_X1 U14378 ( .A1(n14844), .A2(n12066), .ZN(n11898) );
  NAND2_X1 U14379 ( .A1(n11899), .A2(n11898), .ZN(n11902) );
  AOI22_X1 U14380 ( .A1(n12085), .A2(n13140), .B1(n14844), .B2(n11863), .ZN(
        n11900) );
  INV_X1 U14381 ( .A(n11900), .ZN(n11901) );
  NAND2_X1 U14382 ( .A1(n11907), .A2(n11863), .ZN(n11905) );
  NAND2_X1 U14383 ( .A1(n13139), .A2(n12066), .ZN(n11904) );
  NAND2_X1 U14384 ( .A1(n11905), .A2(n11904), .ZN(n11906) );
  AOI22_X1 U14385 ( .A1(n11907), .A2(n12059), .B1(n11863), .B2(n13139), .ZN(
        n11908) );
  NAND2_X1 U14386 ( .A1(n11910), .A2(n11909), .ZN(n11911) );
  NAND2_X1 U14387 ( .A1(n13080), .A2(n12066), .ZN(n11913) );
  NAND2_X1 U14388 ( .A1(n13138), .A2(n11863), .ZN(n11912) );
  NAND2_X1 U14389 ( .A1(n11913), .A2(n11912), .ZN(n11915) );
  AOI22_X1 U14390 ( .A1(n13080), .A2(n11863), .B1(n12085), .B2(n13138), .ZN(
        n11914) );
  NAND2_X1 U14391 ( .A1(n11919), .A2(n11863), .ZN(n11918) );
  NAND2_X1 U14392 ( .A1(n13137), .A2(n12059), .ZN(n11917) );
  NAND2_X1 U14393 ( .A1(n11918), .A2(n11917), .ZN(n11925) );
  NAND2_X1 U14394 ( .A1(n11919), .A2(n12066), .ZN(n11920) );
  OAI21_X1 U14395 ( .B1(n12059), .B2(n11921), .A(n11920), .ZN(n11922) );
  NAND2_X1 U14396 ( .A1(n11923), .A2(n11922), .ZN(n11929) );
  INV_X1 U14397 ( .A(n11924), .ZN(n11927) );
  INV_X1 U14398 ( .A(n11925), .ZN(n11926) );
  NAND2_X1 U14399 ( .A1(n11927), .A2(n11926), .ZN(n11928) );
  NAND2_X1 U14400 ( .A1(n11932), .A2(n12066), .ZN(n11931) );
  NAND2_X1 U14401 ( .A1(n13136), .A2(n11863), .ZN(n11930) );
  NAND2_X1 U14402 ( .A1(n11931), .A2(n11930), .ZN(n11935) );
  AOI22_X1 U14403 ( .A1(n11932), .A2(n11863), .B1(n12085), .B2(n13136), .ZN(
        n11933) );
  INV_X1 U14404 ( .A(n11933), .ZN(n11934) );
  INV_X1 U14405 ( .A(n11935), .ZN(n11936) );
  NAND2_X1 U14406 ( .A1(n13477), .A2(n11863), .ZN(n11938) );
  NAND2_X1 U14407 ( .A1(n13135), .A2(n12059), .ZN(n11937) );
  NAND2_X1 U14408 ( .A1(n13477), .A2(n12085), .ZN(n11939) );
  OAI21_X1 U14409 ( .B1(n12085), .B2(n11940), .A(n11939), .ZN(n11941) );
  NAND2_X1 U14410 ( .A1(n11946), .A2(n12085), .ZN(n11945) );
  NAND2_X1 U14411 ( .A1(n13134), .A2(n11863), .ZN(n11944) );
  NAND2_X1 U14412 ( .A1(n11945), .A2(n11944), .ZN(n11949) );
  AOI22_X1 U14413 ( .A1(n11946), .A2(n11863), .B1(n12085), .B2(n13134), .ZN(
        n11947) );
  INV_X1 U14414 ( .A(n11947), .ZN(n11948) );
  NAND2_X1 U14415 ( .A1(n11953), .A2(n11863), .ZN(n11952) );
  NAND2_X1 U14416 ( .A1(n13133), .A2(n12066), .ZN(n11951) );
  NAND2_X1 U14417 ( .A1(n11953), .A2(n12085), .ZN(n11954) );
  NAND2_X1 U14418 ( .A1(n11961), .A2(n12085), .ZN(n11960) );
  NAND2_X1 U14419 ( .A1(n13131), .A2(n11863), .ZN(n11959) );
  NAND2_X1 U14420 ( .A1(n11960), .A2(n11959), .ZN(n11963) );
  AOI22_X1 U14421 ( .A1(n11961), .A2(n11863), .B1(n12085), .B2(n13131), .ZN(
        n11962) );
  NAND2_X1 U14422 ( .A1(n11969), .A2(n11863), .ZN(n11965) );
  NAND2_X1 U14423 ( .A1(n13130), .A2(n12085), .ZN(n11964) );
  NAND2_X1 U14424 ( .A1(n11965), .A2(n11964), .ZN(n11971) );
  AOI22_X1 U14425 ( .A1(n11966), .A2(n12085), .B1(n11863), .B2(n13129), .ZN(
        n11989) );
  OAI22_X1 U14426 ( .A1(n11968), .A2(n12085), .B1(n11967), .B2(n11863), .ZN(
        n11988) );
  AOI22_X1 U14427 ( .A1(n11969), .A2(n12059), .B1(n11863), .B2(n13130), .ZN(
        n11970) );
  AOI21_X1 U14428 ( .B1(n11972), .B2(n11971), .A(n11970), .ZN(n11973) );
  NAND2_X1 U14429 ( .A1(n11978), .A2(n12085), .ZN(n11976) );
  NAND2_X1 U14430 ( .A1(n13126), .A2(n11863), .ZN(n11975) );
  NAND2_X1 U14431 ( .A1(n11976), .A2(n11975), .ZN(n12000) );
  AND2_X1 U14432 ( .A1(n13126), .A2(n12085), .ZN(n11977) );
  AOI21_X1 U14433 ( .B1(n11978), .B2(n11863), .A(n11977), .ZN(n12006) );
  NAND2_X1 U14434 ( .A1(n12000), .A2(n12006), .ZN(n11983) );
  AND2_X1 U14435 ( .A1(n13127), .A2(n12085), .ZN(n11979) );
  AOI21_X1 U14436 ( .B1(n13551), .B2(n11863), .A(n11979), .ZN(n11994) );
  NAND2_X1 U14437 ( .A1(n13551), .A2(n12085), .ZN(n11981) );
  NAND2_X1 U14438 ( .A1(n13127), .A2(n11863), .ZN(n11980) );
  NAND2_X1 U14439 ( .A1(n11981), .A2(n11980), .ZN(n11993) );
  NAND2_X1 U14440 ( .A1(n11994), .A2(n11993), .ZN(n11982) );
  AND2_X1 U14441 ( .A1(n13128), .A2(n12085), .ZN(n11984) );
  AOI21_X1 U14442 ( .B1(n13617), .B2(n11863), .A(n11984), .ZN(n11997) );
  NAND2_X1 U14443 ( .A1(n13617), .A2(n12085), .ZN(n11986) );
  NAND2_X1 U14444 ( .A1(n13128), .A2(n11863), .ZN(n11985) );
  NAND2_X1 U14445 ( .A1(n11986), .A2(n11985), .ZN(n11998) );
  AND2_X1 U14446 ( .A1(n11997), .A2(n11998), .ZN(n11987) );
  OR2_X1 U14447 ( .A1(n11999), .A2(n11987), .ZN(n11992) );
  INV_X1 U14448 ( .A(n11992), .ZN(n12010) );
  INV_X1 U14449 ( .A(n11988), .ZN(n11991) );
  INV_X1 U14450 ( .A(n11989), .ZN(n11990) );
  INV_X1 U14451 ( .A(n11993), .ZN(n11996) );
  INV_X1 U14452 ( .A(n11994), .ZN(n11995) );
  NAND2_X1 U14453 ( .A1(n11996), .A2(n11995), .ZN(n12005) );
  INV_X1 U14454 ( .A(n11978), .ZN(n13035) );
  NAND3_X1 U14455 ( .A1(n12005), .A2(n13035), .A3(n13066), .ZN(n12002) );
  INV_X1 U14456 ( .A(n12000), .ZN(n12001) );
  NAND2_X1 U14457 ( .A1(n12002), .A2(n12001), .ZN(n12003) );
  OAI211_X1 U14458 ( .C1(n12006), .C2(n12005), .A(n12004), .B(n12003), .ZN(
        n12007) );
  INV_X1 U14459 ( .A(n12007), .ZN(n12008) );
  NAND2_X1 U14460 ( .A1(n6488), .A2(n12008), .ZN(n12009) );
  INV_X1 U14461 ( .A(n12014), .ZN(n12016) );
  AOI22_X1 U14462 ( .A1(n13541), .A2(n11863), .B1(n12085), .B2(n12981), .ZN(
        n12012) );
  AOI22_X1 U14463 ( .A1(n13537), .A2(n11863), .B1(n12085), .B2(n13125), .ZN(
        n12018) );
  AOI22_X1 U14464 ( .A1(n13537), .A2(n12085), .B1(n11863), .B2(n13125), .ZN(
        n12021) );
  OAI22_X1 U14465 ( .A1(n13603), .A2(n11863), .B1(n12085), .B2(n12023), .ZN(
        n12025) );
  AOI22_X1 U14466 ( .A1(n13387), .A2(n11863), .B1(n12085), .B2(n13124), .ZN(
        n12024) );
  OAI22_X1 U14467 ( .A1(n13376), .A2(n12085), .B1(n13059), .B2(n11863), .ZN(
        n12028) );
  INV_X1 U14468 ( .A(n12028), .ZN(n12026) );
  OAI22_X1 U14469 ( .A1(n13376), .A2(n11863), .B1(n12085), .B2(n13059), .ZN(
        n12027) );
  AOI22_X1 U14470 ( .A1(n13591), .A2(n12085), .B1(n11863), .B2(n13122), .ZN(
        n12031) );
  INV_X1 U14471 ( .A(n12031), .ZN(n12029) );
  INV_X1 U14472 ( .A(n13591), .ZN(n13359) );
  OAI22_X1 U14473 ( .A1(n13359), .A2(n12085), .B1(n12030), .B2(n11863), .ZN(
        n12032) );
  OAI22_X1 U14474 ( .A1(n13348), .A2(n11863), .B1(n12085), .B2(n13040), .ZN(
        n12033) );
  AOI22_X1 U14475 ( .A1(n13331), .A2(n12085), .B1(n11863), .B2(n13120), .ZN(
        n12039) );
  INV_X1 U14476 ( .A(n12039), .ZN(n12035) );
  INV_X1 U14477 ( .A(n13120), .ZN(n12036) );
  OAI22_X1 U14478 ( .A1(n13584), .A2(n12085), .B1(n12036), .B2(n11863), .ZN(
        n12037) );
  OAI22_X1 U14479 ( .A1(n13320), .A2(n12085), .B1(n13093), .B2(n11863), .ZN(
        n12040) );
  AOI22_X1 U14480 ( .A1(n13500), .A2(n12059), .B1(n11863), .B2(n13119), .ZN(
        n12044) );
  OAI22_X1 U14481 ( .A1(n13102), .A2(n12085), .B1(n12042), .B2(n11863), .ZN(
        n12043) );
  NAND2_X1 U14482 ( .A1(n12045), .A2(n12044), .ZN(n12046) );
  INV_X1 U14483 ( .A(n12069), .ZN(n12048) );
  OAI22_X1 U14484 ( .A1(n13286), .A2(n12059), .B1(n13095), .B2(n11863), .ZN(
        n12068) );
  INV_X1 U14485 ( .A(n12068), .ZN(n12047) );
  NAND2_X1 U14486 ( .A1(n12050), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12051) );
  NAND2_X1 U14487 ( .A1(n12412), .A2(n11863), .ZN(n12084) );
  NAND2_X1 U14488 ( .A1(n6744), .A2(n12149), .ZN(n12094) );
  NAND4_X1 U14489 ( .A1(n12084), .A2(n8178), .A3(n12053), .A4(n12094), .ZN(
        n12054) );
  NAND2_X1 U14490 ( .A1(n12054), .A2(n13116), .ZN(n12055) );
  AOI22_X1 U14491 ( .A1(n13564), .A2(n11863), .B1(n12085), .B2(n13116), .ZN(
        n12079) );
  OAI22_X1 U14492 ( .A1(n12060), .A2(n11863), .B1(n12059), .B2(n12993), .ZN(
        n12076) );
  AOI22_X1 U14493 ( .A1(n12080), .A2(n12079), .B1(n12075), .B2(n12076), .ZN(
        n12061) );
  NAND2_X1 U14494 ( .A1(n13489), .A2(n11863), .ZN(n12063) );
  NAND2_X1 U14495 ( .A1(n13117), .A2(n12085), .ZN(n12062) );
  NAND2_X1 U14496 ( .A1(n12063), .A2(n12062), .ZN(n12071) );
  AND2_X1 U14497 ( .A1(n13117), .A2(n11863), .ZN(n12064) );
  AOI21_X1 U14498 ( .B1(n13489), .B2(n12085), .A(n12064), .ZN(n12072) );
  NOR2_X1 U14499 ( .A1(n12071), .A2(n12072), .ZN(n12065) );
  INV_X1 U14500 ( .A(n13095), .ZN(n13118) );
  AOI22_X1 U14501 ( .A1(n13569), .A2(n12066), .B1(n11863), .B2(n13118), .ZN(
        n12067) );
  INV_X1 U14502 ( .A(n12071), .ZN(n12074) );
  INV_X1 U14503 ( .A(n12072), .ZN(n12073) );
  OAI22_X1 U14504 ( .A1(n12076), .A2(n12075), .B1(n12074), .B2(n12073), .ZN(
        n12078) );
  INV_X1 U14505 ( .A(n12079), .ZN(n12082) );
  NAND2_X1 U14506 ( .A1(n12082), .A2(n12081), .ZN(n12083) );
  NAND2_X1 U14507 ( .A1(n12084), .A2(n11863), .ZN(n12087) );
  NAND2_X1 U14508 ( .A1(n12412), .A2(n12085), .ZN(n12086) );
  MUX2_X1 U14509 ( .A(n12087), .B(n12086), .S(n12422), .Z(n12088) );
  AOI21_X1 U14510 ( .B1(n12090), .B2(n12089), .A(n13249), .ZN(n12091) );
  AOI21_X1 U14511 ( .B1(n12103), .B2(n12138), .A(n12091), .ZN(n12092) );
  INV_X1 U14512 ( .A(n12092), .ZN(n12097) );
  NAND3_X1 U14513 ( .A1(n8178), .A2(n12103), .A3(n8221), .ZN(n12093) );
  NAND2_X1 U14514 ( .A1(n12094), .A2(n12093), .ZN(n12095) );
  NAND2_X1 U14515 ( .A1(n12098), .A2(n12095), .ZN(n12096) );
  OAI21_X1 U14516 ( .B1(n12098), .B2(n12097), .A(n12096), .ZN(n12144) );
  NOR2_X1 U14517 ( .A1(n12100), .A2(n12099), .ZN(n13299) );
  XNOR2_X1 U14518 ( .A(n13587), .B(n13040), .ZN(n13339) );
  NAND2_X1 U14519 ( .A1(n12102), .A2(n12101), .ZN(n13378) );
  NAND4_X1 U14520 ( .A1(n12105), .A2(n12106), .A3(n12104), .A4(n12103), .ZN(
        n12109) );
  NOR3_X1 U14521 ( .A1(n12109), .A2(n12108), .A3(n12107), .ZN(n12112) );
  NAND4_X1 U14522 ( .A1(n12113), .A2(n12112), .A3(n12111), .A4(n12110), .ZN(
        n12114) );
  OR4_X1 U14523 ( .A1(n12117), .A2(n12116), .A3(n12115), .A4(n12114), .ZN(
        n12118) );
  NOR2_X1 U14524 ( .A1(n12119), .A2(n12118), .ZN(n12121) );
  NAND3_X1 U14525 ( .A1(n12122), .A2(n12121), .A3(n12120), .ZN(n12123) );
  NOR2_X1 U14526 ( .A1(n12124), .A2(n12123), .ZN(n12126) );
  NAND4_X1 U14527 ( .A1(n13431), .A2(n12126), .A3(n13452), .A4(n12125), .ZN(
        n12127) );
  NOR2_X1 U14528 ( .A1(n13411), .A2(n12127), .ZN(n12130) );
  NAND2_X1 U14529 ( .A1(n12129), .A2(n12128), .ZN(n13401) );
  NAND4_X1 U14530 ( .A1(n13378), .A2(n12130), .A3(n13392), .A4(n13401), .ZN(
        n12131) );
  NOR3_X1 U14531 ( .A1(n13339), .A2(n13356), .A3(n12131), .ZN(n12132) );
  NAND4_X1 U14532 ( .A1(n13299), .A2(n12132), .A3(n13312), .A4(n13329), .ZN(
        n12133) );
  NOR4_X1 U14533 ( .A1(n12134), .A2(n13280), .A3(n13261), .A4(n12133), .ZN(
        n12136) );
  XNOR2_X1 U14534 ( .A(n13564), .B(n13116), .ZN(n12135) );
  NAND3_X1 U14535 ( .A1(n7390), .A2(n12136), .A3(n12135), .ZN(n12137) );
  XNOR2_X1 U14536 ( .A(n12137), .B(n8221), .ZN(n12139) );
  NAND2_X1 U14537 ( .A1(n12139), .A2(n12138), .ZN(n12140) );
  NAND3_X1 U14538 ( .A1(n12146), .A2(n12145), .A3(n13050), .ZN(n12147) );
  OAI211_X1 U14539 ( .C1(n12149), .C2(n12148), .A(n12147), .B(P2_B_REG_SCAN_IN), .ZN(n12150) );
  NAND2_X1 U14540 ( .A1(n12151), .A2(n12150), .ZN(P2_U3328) );
  INV_X1 U14541 ( .A(n12152), .ZN(n13631) );
  OAI222_X1 U14542 ( .A1(P1_U3086), .A2(n12154), .B1(n14204), .B2(n13631), 
        .C1(n12153), .C2(n14201), .ZN(P1_U3325) );
  OAI222_X1 U14543 ( .A1(n8883), .A2(P1_U3086), .B1(n14204), .B2(n12156), .C1(
        n12155), .C2(n14201), .ZN(P1_U3336) );
  XNOR2_X1 U14544 ( .A(n12929), .B(n12191), .ZN(n12476) );
  NAND2_X1 U14545 ( .A1(n12476), .A2(n12545), .ZN(n12162) );
  XNOR2_X1 U14546 ( .A(n12925), .B(n10487), .ZN(n12163) );
  XNOR2_X1 U14547 ( .A(n12163), .B(n12544), .ZN(n12513) );
  INV_X1 U14548 ( .A(n12163), .ZN(n12164) );
  XNOR2_X1 U14549 ( .A(n12455), .B(n10487), .ZN(n12165) );
  XOR2_X1 U14550 ( .A(n12796), .B(n12165), .Z(n12449) );
  NAND2_X1 U14551 ( .A1(n12450), .A2(n12449), .ZN(n12168) );
  INV_X1 U14552 ( .A(n12165), .ZN(n12166) );
  NAND2_X1 U14553 ( .A1(n12166), .A2(n9290), .ZN(n12167) );
  NAND2_X1 U14554 ( .A1(n12168), .A2(n12167), .ZN(n12495) );
  XNOR2_X1 U14555 ( .A(n12774), .B(n10487), .ZN(n12169) );
  XNOR2_X1 U14556 ( .A(n12169), .B(n12757), .ZN(n12494) );
  INV_X1 U14557 ( .A(n12169), .ZN(n12170) );
  NAND2_X1 U14558 ( .A1(n12170), .A2(n12757), .ZN(n12171) );
  XNOR2_X1 U14559 ( .A(n12762), .B(n10487), .ZN(n12172) );
  NAND2_X1 U14560 ( .A1(n12172), .A2(n12769), .ZN(n12173) );
  OAI21_X1 U14561 ( .B1(n12172), .B2(n12769), .A(n12173), .ZN(n12459) );
  XNOR2_X1 U14562 ( .A(n12510), .B(n10487), .ZN(n12174) );
  OAI21_X1 U14563 ( .B1(n12175), .B2(n12174), .A(n12176), .ZN(n12503) );
  XNOR2_X1 U14564 ( .A(n12446), .B(n10487), .ZN(n12177) );
  XNOR2_X1 U14565 ( .A(n12851), .B(n10487), .ZN(n12179) );
  NAND2_X1 U14566 ( .A1(n12179), .A2(n12702), .ZN(n12466) );
  INV_X1 U14567 ( .A(n12179), .ZN(n12180) );
  NAND2_X1 U14568 ( .A1(n12180), .A2(n12734), .ZN(n12181) );
  AND2_X1 U14569 ( .A1(n12466), .A2(n12181), .ZN(n12485) );
  NAND2_X1 U14570 ( .A1(n12182), .A2(n12485), .ZN(n12465) );
  NAND2_X1 U14571 ( .A1(n12465), .A2(n12466), .ZN(n12186) );
  XNOR2_X1 U14572 ( .A(n12847), .B(n10487), .ZN(n12183) );
  NAND2_X1 U14573 ( .A1(n12183), .A2(n12719), .ZN(n12187) );
  INV_X1 U14574 ( .A(n12183), .ZN(n12184) );
  INV_X1 U14575 ( .A(n12719), .ZN(n12542) );
  NAND2_X1 U14576 ( .A1(n12184), .A2(n12542), .ZN(n12185) );
  AND2_X1 U14577 ( .A1(n12187), .A2(n12185), .ZN(n12467) );
  XNOR2_X1 U14578 ( .A(n12695), .B(n12191), .ZN(n12188) );
  NOR2_X1 U14579 ( .A1(n12188), .A2(n7491), .ZN(n12189) );
  AOI21_X1 U14580 ( .B1(n12188), .B2(n7491), .A(n12189), .ZN(n12527) );
  INV_X1 U14581 ( .A(n12189), .ZN(n12190) );
  XNOR2_X1 U14582 ( .A(n12839), .B(n12191), .ZN(n12192) );
  NOR2_X1 U14583 ( .A1(n12192), .A2(n12541), .ZN(n12193) );
  AOI21_X1 U14584 ( .B1(n12192), .B2(n12541), .A(n12193), .ZN(n12434) );
  XNOR2_X1 U14585 ( .A(n12194), .B(n10487), .ZN(n12195) );
  NOR2_X1 U14586 ( .A1(n12196), .A2(n12516), .ZN(n12199) );
  AOI22_X1 U14587 ( .A1(n12666), .A2(n12505), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12197) );
  OAI21_X1 U14588 ( .B1(n12690), .B2(n12508), .A(n12197), .ZN(n12198) );
  AOI211_X1 U14589 ( .C1(n12200), .C2(n12521), .A(n12199), .B(n12198), .ZN(
        n12201) );
  OAI21_X1 U14590 ( .B1(n12202), .B2(n12523), .A(n12201), .ZN(P3_U3160) );
  OAI22_X1 U14591 ( .A1(n14526), .A2(n12274), .B1(n12206), .B2(n12317), .ZN(
        n12216) );
  NAND2_X1 U14592 ( .A1(n14343), .A2(n12333), .ZN(n12208) );
  NAND2_X1 U14593 ( .A1(n14483), .A2(n12312), .ZN(n12207) );
  NAND2_X1 U14594 ( .A1(n12208), .A2(n12207), .ZN(n12209) );
  XNOR2_X1 U14595 ( .A(n12209), .B(n12334), .ZN(n12215) );
  XOR2_X1 U14596 ( .A(n12216), .B(n12215), .Z(n13748) );
  NAND2_X1 U14597 ( .A1(n12214), .A2(n12333), .ZN(n12211) );
  NAND2_X1 U14598 ( .A1(n14338), .A2(n12319), .ZN(n12210) );
  NAND2_X1 U14599 ( .A1(n12211), .A2(n12210), .ZN(n12212) );
  XNOR2_X1 U14600 ( .A(n12212), .B(n12315), .ZN(n12220) );
  NOR2_X1 U14601 ( .A1(n12317), .A2(n13753), .ZN(n12213) );
  AOI21_X1 U14602 ( .B1(n12214), .B2(n12312), .A(n12213), .ZN(n12221) );
  XNOR2_X1 U14603 ( .A(n12220), .B(n12221), .ZN(n14478) );
  INV_X1 U14604 ( .A(n12215), .ZN(n12218) );
  INV_X1 U14605 ( .A(n12216), .ZN(n12217) );
  NOR2_X1 U14606 ( .A1(n12218), .A2(n12217), .ZN(n14479) );
  NOR2_X1 U14607 ( .A1(n14478), .A2(n14479), .ZN(n12219) );
  NAND2_X1 U14608 ( .A1(n12222), .A2(n12333), .ZN(n12224) );
  NAND2_X1 U14609 ( .A1(n14484), .A2(n12319), .ZN(n12223) );
  NAND2_X1 U14610 ( .A1(n12224), .A2(n12223), .ZN(n12225) );
  XNOR2_X1 U14611 ( .A(n12225), .B(n12334), .ZN(n12228) );
  OAI22_X1 U14612 ( .A1(n14162), .A2(n12274), .B1(n12226), .B2(n12317), .ZN(
        n13787) );
  INV_X1 U14613 ( .A(n12227), .ZN(n12229) );
  NAND2_X1 U14614 ( .A1(n12229), .A2(n12228), .ZN(n12230) );
  AOI22_X1 U14615 ( .A1(n12232), .A2(n12333), .B1(n12319), .B2(n13803), .ZN(
        n12231) );
  XNOR2_X1 U14616 ( .A(n12231), .B(n12334), .ZN(n12235) );
  AOI22_X1 U14617 ( .A1(n12232), .A2(n12319), .B1(n10923), .B2(n13803), .ZN(
        n12234) );
  XNOR2_X1 U14618 ( .A(n12235), .B(n12234), .ZN(n13708) );
  INV_X1 U14619 ( .A(n13708), .ZN(n12233) );
  NAND2_X1 U14620 ( .A1(n12235), .A2(n12234), .ZN(n12236) );
  NAND2_X1 U14621 ( .A1(n14150), .A2(n12333), .ZN(n12238) );
  NAND2_X1 U14622 ( .A1(n14052), .A2(n12319), .ZN(n12237) );
  NAND2_X1 U14623 ( .A1(n12238), .A2(n12237), .ZN(n12239) );
  XNOR2_X1 U14624 ( .A(n12239), .B(n12334), .ZN(n13717) );
  NAND2_X1 U14625 ( .A1(n14150), .A2(n12312), .ZN(n12241) );
  NAND2_X1 U14626 ( .A1(n10923), .A2(n14052), .ZN(n12240) );
  NAND2_X1 U14627 ( .A1(n12241), .A2(n12240), .ZN(n13716) );
  NAND2_X1 U14628 ( .A1(n13717), .A2(n13716), .ZN(n12242) );
  NOR2_X1 U14629 ( .A1(n12317), .A2(n13681), .ZN(n12243) );
  AOI21_X1 U14630 ( .B1(n14144), .B2(n12319), .A(n12243), .ZN(n12252) );
  NAND2_X1 U14631 ( .A1(n14144), .A2(n12333), .ZN(n12245) );
  NAND2_X1 U14632 ( .A1(n14038), .A2(n12312), .ZN(n12244) );
  NAND2_X1 U14633 ( .A1(n12245), .A2(n12244), .ZN(n12246) );
  XNOR2_X1 U14634 ( .A(n12246), .B(n12334), .ZN(n12251) );
  XOR2_X1 U14635 ( .A(n12252), .B(n12251), .Z(n13768) );
  NAND2_X1 U14636 ( .A1(n12381), .A2(n12333), .ZN(n12248) );
  NAND2_X1 U14637 ( .A1(n14051), .A2(n12312), .ZN(n12247) );
  NAND2_X1 U14638 ( .A1(n12248), .A2(n12247), .ZN(n12249) );
  XNOR2_X1 U14639 ( .A(n12249), .B(n12315), .ZN(n12255) );
  AND2_X1 U14640 ( .A1(n10923), .A2(n14051), .ZN(n12250) );
  AOI21_X1 U14641 ( .B1(n12381), .B2(n12319), .A(n12250), .ZN(n12256) );
  XNOR2_X1 U14642 ( .A(n12255), .B(n12256), .ZN(n13677) );
  INV_X1 U14643 ( .A(n12251), .ZN(n12253) );
  AND2_X1 U14644 ( .A1(n12253), .A2(n12252), .ZN(n13678) );
  NOR2_X1 U14645 ( .A1(n13677), .A2(n13678), .ZN(n12254) );
  INV_X1 U14646 ( .A(n12255), .ZN(n12258) );
  INV_X1 U14647 ( .A(n12256), .ZN(n12257) );
  NAND2_X1 U14648 ( .A1(n12258), .A2(n12257), .ZN(n12259) );
  OAI22_X1 U14649 ( .A1(n12260), .A2(n12274), .B1(n12368), .B2(n12317), .ZN(
        n12264) );
  NAND2_X1 U14650 ( .A1(n14130), .A2(n12333), .ZN(n12262) );
  NAND2_X1 U14651 ( .A1(n14039), .A2(n12312), .ZN(n12261) );
  NAND2_X1 U14652 ( .A1(n12262), .A2(n12261), .ZN(n12263) );
  XNOR2_X1 U14653 ( .A(n12263), .B(n12334), .ZN(n12265) );
  XOR2_X1 U14654 ( .A(n12264), .B(n12265), .Z(n13738) );
  NAND2_X1 U14655 ( .A1(n12265), .A2(n12264), .ZN(n12266) );
  NAND2_X1 U14656 ( .A1(n14012), .A2(n12333), .ZN(n12268) );
  NAND2_X1 U14657 ( .A1(n13802), .A2(n12312), .ZN(n12267) );
  NAND2_X1 U14658 ( .A1(n12268), .A2(n12267), .ZN(n12269) );
  XNOR2_X1 U14659 ( .A(n12269), .B(n12315), .ZN(n12272) );
  AND2_X1 U14660 ( .A1(n13802), .A2(n10923), .ZN(n12270) );
  AOI21_X1 U14661 ( .B1(n14012), .B2(n12319), .A(n12270), .ZN(n12271) );
  OAI21_X1 U14662 ( .B1(n12272), .B2(n12271), .A(n13758), .ZN(n13686) );
  INV_X1 U14663 ( .A(n13686), .ZN(n12273) );
  OAI22_X1 U14664 ( .A1(n14119), .A2(n11842), .B1(n6899), .B2(n12274), .ZN(
        n12275) );
  XNOR2_X1 U14665 ( .A(n12275), .B(n12315), .ZN(n12278) );
  OR2_X1 U14666 ( .A1(n14119), .A2(n12274), .ZN(n12277) );
  NAND2_X1 U14667 ( .A1(n10923), .A2(n14004), .ZN(n12276) );
  INV_X1 U14668 ( .A(n12278), .ZN(n12281) );
  INV_X1 U14669 ( .A(n12279), .ZN(n12280) );
  NAND2_X1 U14670 ( .A1(n12281), .A2(n12280), .ZN(n12282) );
  NAND2_X1 U14671 ( .A1(n13665), .A2(n13666), .ZN(n12292) );
  NAND2_X1 U14672 ( .A1(n8838), .A2(n12333), .ZN(n12284) );
  NAND2_X1 U14673 ( .A1(n12319), .A2(n13958), .ZN(n12283) );
  NAND2_X1 U14674 ( .A1(n12284), .A2(n12283), .ZN(n12285) );
  XNOR2_X1 U14675 ( .A(n12285), .B(n12315), .ZN(n12287) );
  INV_X1 U14676 ( .A(n13958), .ZN(n12374) );
  NOR2_X1 U14677 ( .A1(n12317), .A2(n12374), .ZN(n12286) );
  AOI21_X1 U14678 ( .B1(n8838), .B2(n12319), .A(n12286), .ZN(n12288) );
  INV_X1 U14679 ( .A(n12287), .ZN(n12290) );
  INV_X1 U14680 ( .A(n12288), .ZN(n12289) );
  NAND2_X1 U14681 ( .A1(n12290), .A2(n12289), .ZN(n12291) );
  NAND2_X1 U14682 ( .A1(n12292), .A2(n13667), .ZN(n13669) );
  NAND2_X1 U14683 ( .A1(n13669), .A2(n13727), .ZN(n12302) );
  NAND2_X1 U14684 ( .A1(n13964), .A2(n12333), .ZN(n12294) );
  NAND2_X1 U14685 ( .A1(n12319), .A2(n13943), .ZN(n12293) );
  NAND2_X1 U14686 ( .A1(n12294), .A2(n12293), .ZN(n12295) );
  XNOR2_X1 U14687 ( .A(n12295), .B(n12315), .ZN(n12297) );
  NOR2_X1 U14688 ( .A1(n12317), .A2(n12358), .ZN(n12296) );
  AOI21_X1 U14689 ( .B1(n13964), .B2(n12319), .A(n12296), .ZN(n12298) );
  NAND2_X1 U14690 ( .A1(n12297), .A2(n12298), .ZN(n13694) );
  INV_X1 U14691 ( .A(n12297), .ZN(n12300) );
  INV_X1 U14692 ( .A(n12298), .ZN(n12299) );
  NAND2_X1 U14693 ( .A1(n12300), .A2(n12299), .ZN(n12301) );
  NAND2_X1 U14694 ( .A1(n12302), .A2(n13728), .ZN(n13693) );
  NAND2_X1 U14695 ( .A1(n13693), .A2(n13694), .ZN(n12310) );
  NAND2_X1 U14696 ( .A1(n13940), .A2(n12333), .ZN(n12304) );
  NAND2_X1 U14697 ( .A1(n13959), .A2(n12312), .ZN(n12303) );
  NAND2_X1 U14698 ( .A1(n12304), .A2(n12303), .ZN(n12305) );
  XNOR2_X1 U14699 ( .A(n12305), .B(n12315), .ZN(n12308) );
  NOR2_X1 U14700 ( .A1(n12317), .A2(n13779), .ZN(n12306) );
  AOI21_X1 U14701 ( .B1(n13940), .B2(n12319), .A(n12306), .ZN(n12307) );
  NAND2_X1 U14702 ( .A1(n12308), .A2(n12307), .ZN(n12311) );
  OR2_X1 U14703 ( .A1(n12308), .A2(n12307), .ZN(n12309) );
  NAND2_X1 U14704 ( .A1(n13921), .A2(n12333), .ZN(n12314) );
  NAND2_X1 U14705 ( .A1(n13944), .A2(n12312), .ZN(n12313) );
  NAND2_X1 U14706 ( .A1(n12314), .A2(n12313), .ZN(n12316) );
  XNOR2_X1 U14707 ( .A(n12316), .B(n12315), .ZN(n12321) );
  INV_X1 U14708 ( .A(n12321), .ZN(n12323) );
  NOR2_X1 U14709 ( .A1(n12317), .A2(n13701), .ZN(n12318) );
  AOI21_X1 U14710 ( .B1(n13921), .B2(n12319), .A(n12318), .ZN(n12320) );
  INV_X1 U14711 ( .A(n12320), .ZN(n12322) );
  AND2_X1 U14712 ( .A1(n12321), .A2(n12320), .ZN(n12324) );
  AOI21_X1 U14713 ( .B1(n12323), .B2(n12322), .A(n12324), .ZN(n13777) );
  NAND2_X1 U14714 ( .A1(n14087), .A2(n12333), .ZN(n12326) );
  NAND2_X1 U14715 ( .A1(n12312), .A2(n13801), .ZN(n12325) );
  NAND2_X1 U14716 ( .A1(n12326), .A2(n12325), .ZN(n12327) );
  XNOR2_X1 U14717 ( .A(n12327), .B(n12334), .ZN(n12331) );
  NAND2_X1 U14718 ( .A1(n14087), .A2(n12319), .ZN(n12329) );
  NAND2_X1 U14719 ( .A1(n10923), .A2(n13801), .ZN(n12328) );
  NAND2_X1 U14720 ( .A1(n12329), .A2(n12328), .ZN(n12330) );
  NOR2_X1 U14721 ( .A1(n12331), .A2(n12330), .ZN(n12332) );
  AOI21_X1 U14722 ( .B1(n12331), .B2(n12330), .A(n12332), .ZN(n13657) );
  AOI22_X1 U14723 ( .A1(n14082), .A2(n12333), .B1(n12319), .B2(n13800), .ZN(
        n12335) );
  XNOR2_X1 U14724 ( .A(n12335), .B(n12334), .ZN(n12337) );
  AOI22_X1 U14725 ( .A1(n14082), .A2(n12319), .B1(n10923), .B2(n13800), .ZN(
        n12336) );
  XNOR2_X1 U14726 ( .A(n12337), .B(n12336), .ZN(n12338) );
  INV_X1 U14727 ( .A(n13912), .ZN(n12342) );
  NAND2_X1 U14728 ( .A1(n13799), .A2(n14050), .ZN(n12340) );
  NAND2_X1 U14729 ( .A1(n13801), .A2(n14339), .ZN(n12339) );
  NAND2_X1 U14730 ( .A1(n12340), .A2(n12339), .ZN(n14081) );
  AOI22_X1 U14731 ( .A1(n14584), .A2(n14081), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12341) );
  OAI21_X1 U14732 ( .B1(n12342), .B2(n14572), .A(n12341), .ZN(n12343) );
  AOI21_X1 U14733 ( .B1(n14082), .B2(n13739), .A(n12343), .ZN(n12344) );
  OAI21_X1 U14734 ( .B1(n12345), .B2(n14565), .A(n12344), .ZN(P1_U3220) );
  OR2_X1 U14735 ( .A1(n14144), .A2(n14038), .ZN(n12347) );
  NAND2_X1 U14736 ( .A1(n14144), .A2(n14038), .ZN(n12348) );
  NAND2_X1 U14737 ( .A1(n14130), .A2(n14039), .ZN(n12351) );
  NAND2_X1 U14738 ( .A1(n14024), .A2(n12351), .ZN(n14005) );
  INV_X1 U14739 ( .A(n14012), .ZN(n12370) );
  INV_X1 U14740 ( .A(n13802), .ZN(n12353) );
  NAND2_X1 U14741 ( .A1(n12370), .A2(n12353), .ZN(n12354) );
  NAND2_X1 U14742 ( .A1(n14119), .A2(n6899), .ZN(n12355) );
  NAND2_X1 U14743 ( .A1(n8838), .A2(n13958), .ZN(n12357) );
  INV_X1 U14744 ( .A(n13956), .ZN(n13953) );
  INV_X1 U14745 ( .A(n13916), .ZN(n13907) );
  NAND2_X1 U14746 ( .A1(n13908), .A2(n13907), .ZN(n13906) );
  INV_X1 U14747 ( .A(n13800), .ZN(n13660) );
  NAND2_X1 U14748 ( .A1(n14035), .A2(n12366), .ZN(n14020) );
  OR2_X1 U14749 ( .A1(n14130), .A2(n12368), .ZN(n12369) );
  NAND2_X1 U14750 ( .A1(n12370), .A2(n13802), .ZN(n12371) );
  OR2_X1 U14751 ( .A1(n14119), .A2(n14004), .ZN(n12373) );
  NAND2_X1 U14752 ( .A1(n8838), .A2(n12374), .ZN(n12375) );
  OR2_X1 U14753 ( .A1(n13964), .A2(n12358), .ZN(n12376) );
  NAND2_X1 U14754 ( .A1(n13940), .A2(n13779), .ZN(n12378) );
  NAND2_X1 U14755 ( .A1(n14076), .A2(n14060), .ZN(n12390) );
  NAND2_X1 U14756 ( .A1(n12383), .A2(P1_B_REG_SCAN_IN), .ZN(n12384) );
  AND2_X1 U14757 ( .A1(n14050), .A2(n12384), .ZN(n13896) );
  NAND2_X1 U14758 ( .A1(n13798), .A2(n13896), .ZN(n14074) );
  OAI22_X1 U14759 ( .A1(n12386), .A2(n14074), .B1(n12385), .B2(n14608), .ZN(
        n12388) );
  NAND2_X1 U14760 ( .A1(n13800), .A2(n14339), .ZN(n14073) );
  NOR2_X1 U14761 ( .A1(n14646), .A2(n14073), .ZN(n12387) );
  AOI211_X1 U14762 ( .C1(n14646), .C2(P1_REG2_REG_29__SCAN_IN), .A(n12388), 
        .B(n12387), .ZN(n12389) );
  OAI211_X1 U14763 ( .C1(n7229), .C2(n14640), .A(n12390), .B(n12389), .ZN(
        n12391) );
  AOI21_X1 U14764 ( .B1(n14045), .B2(n14077), .A(n12391), .ZN(n12392) );
  OAI21_X1 U14765 ( .B1(n14079), .B2(n14352), .A(n12392), .ZN(P1_U3356) );
  INV_X1 U14766 ( .A(n12393), .ZN(n12395) );
  OAI222_X1 U14767 ( .A1(n12396), .A2(n12395), .B1(n12962), .B2(n12394), .C1(
        P3_U3151), .C2(n6436), .ZN(P3_U3268) );
  OAI21_X1 U14768 ( .B1(n12401), .B2(n12400), .A(n12399), .ZN(n12403) );
  OAI22_X1 U14769 ( .A1(n13660), .A2(n14583), .B1(n13701), .B2(n14622), .ZN(
        n12402) );
  INV_X1 U14770 ( .A(n13909), .ZN(n12406) );
  AOI211_X1 U14771 ( .C1(n14087), .C2(n13922), .A(n14058), .B(n12406), .ZN(
        n14086) );
  AOI22_X1 U14772 ( .A1(n14646), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13662), 
        .B2(n14636), .ZN(n12407) );
  OAI21_X1 U14773 ( .B1(n13664), .B2(n14640), .A(n12407), .ZN(n12409) );
  NOR2_X1 U14774 ( .A1(n14090), .A2(n14641), .ZN(n12408) );
  AOI211_X1 U14775 ( .C1(n14086), .C2(n14060), .A(n12409), .B(n12408), .ZN(
        n12410) );
  OAI21_X1 U14776 ( .B1(n14089), .B2(n14646), .A(n12410), .ZN(P1_U3266) );
  INV_X1 U14777 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n12413) );
  NOR2_X2 U14778 ( .A1(n6474), .A2(n13460), .ZN(n12418) );
  AND2_X1 U14779 ( .A1(n12412), .A2(n12411), .ZN(n12419) );
  NOR2_X1 U14780 ( .A1(n12418), .A2(n12419), .ZN(n12415) );
  MUX2_X1 U14781 ( .A(n12413), .B(n12415), .S(n14859), .Z(n12414) );
  OAI21_X1 U14782 ( .B1(n12422), .B2(n13602), .A(n12414), .ZN(P2_U3498) );
  MUX2_X1 U14783 ( .A(n12416), .B(n12415), .S(n14864), .Z(n12417) );
  OAI21_X1 U14784 ( .B1(n12422), .B2(n13534), .A(n12417), .ZN(P2_U3530) );
  NAND2_X1 U14785 ( .A1(n12418), .A2(n13478), .ZN(n12421) );
  INV_X1 U14786 ( .A(n12419), .ZN(n13484) );
  NOR2_X1 U14787 ( .A1(n13428), .A2(n13484), .ZN(n13258) );
  AOI21_X1 U14788 ( .B1(n13428), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13258), 
        .ZN(n12420) );
  OAI211_X1 U14789 ( .C1(n12422), .C2(n13463), .A(n12421), .B(n12420), .ZN(
        P2_U3234) );
  INV_X1 U14790 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n12425) );
  OAI21_X1 U14791 ( .B1(n15096), .B2(n12425), .A(n12424), .ZN(n12426) );
  INV_X1 U14792 ( .A(n12426), .ZN(n12428) );
  INV_X1 U14793 ( .A(n12429), .ZN(n12430) );
  OAI21_X1 U14794 ( .B1(n12431), .B2(n15075), .A(n12430), .ZN(P3_U3204) );
  OAI21_X1 U14795 ( .B1(n12434), .B2(n12433), .A(n12432), .ZN(n12435) );
  NAND2_X1 U14796 ( .A1(n12435), .A2(n12528), .ZN(n12440) );
  OAI22_X1 U14797 ( .A1(n12703), .A2(n12508), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12436), .ZN(n12438) );
  NOR2_X1 U14798 ( .A1(n12674), .A2(n12516), .ZN(n12437) );
  AOI211_X1 U14799 ( .C1(n12680), .C2(n12505), .A(n12438), .B(n12437), .ZN(
        n12439) );
  OAI211_X1 U14800 ( .C1(n12682), .C2(n12538), .A(n12440), .B(n12439), .ZN(
        P3_U3154) );
  AOI21_X1 U14801 ( .B1(n12504), .B2(n12441), .A(n6467), .ZN(n12448) );
  AOI22_X1 U14802 ( .A1(n12734), .A2(n12535), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12443) );
  NAND2_X1 U14803 ( .A1(n12505), .A2(n12739), .ZN(n12442) );
  OAI211_X1 U14804 ( .C1(n12444), .C2(n12508), .A(n12443), .B(n12442), .ZN(
        n12445) );
  AOI21_X1 U14805 ( .B1(n12446), .B2(n12521), .A(n12445), .ZN(n12447) );
  OAI21_X1 U14806 ( .B1(n12448), .B2(n12523), .A(n12447), .ZN(P3_U3156) );
  XNOR2_X1 U14807 ( .A(n12450), .B(n12449), .ZN(n12457) );
  NAND2_X1 U14808 ( .A1(n12505), .A2(n12788), .ZN(n12453) );
  NOR2_X1 U14809 ( .A1(n12451), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12632) );
  AOI21_X1 U14810 ( .B1(n12757), .B2(n12535), .A(n12632), .ZN(n12452) );
  OAI211_X1 U14811 ( .C1(n12813), .C2(n12508), .A(n12453), .B(n12452), .ZN(
        n12454) );
  AOI21_X1 U14812 ( .B1(n12455), .B2(n12521), .A(n12454), .ZN(n12456) );
  OAI21_X1 U14813 ( .B1(n12457), .B2(n12523), .A(n12456), .ZN(P3_U3159) );
  AOI21_X1 U14814 ( .B1(n12459), .B2(n12458), .A(n6596), .ZN(n12464) );
  AOI22_X1 U14815 ( .A1(n12758), .A2(n12535), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12461) );
  NAND2_X1 U14816 ( .A1(n12505), .A2(n12763), .ZN(n12460) );
  OAI211_X1 U14817 ( .C1(n12782), .C2(n12508), .A(n12461), .B(n12460), .ZN(
        n12462) );
  AOI21_X1 U14818 ( .B1(n12762), .B2(n12521), .A(n12462), .ZN(n12463) );
  OAI21_X1 U14819 ( .B1(n12464), .B2(n12523), .A(n12463), .ZN(P3_U3163) );
  INV_X1 U14820 ( .A(n12465), .ZN(n12487) );
  INV_X1 U14821 ( .A(n12466), .ZN(n12468) );
  NOR3_X1 U14822 ( .A1(n12487), .A2(n12468), .A3(n12467), .ZN(n12471) );
  INV_X1 U14823 ( .A(n12469), .ZN(n12470) );
  OAI21_X1 U14824 ( .B1(n12471), .B2(n12470), .A(n12528), .ZN(n12475) );
  AOI22_X1 U14825 ( .A1(n12734), .A2(n12530), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12472) );
  OAI21_X1 U14826 ( .B1(n12703), .B2(n12516), .A(n12472), .ZN(n12473) );
  AOI21_X1 U14827 ( .B1(n12711), .B2(n12505), .A(n12473), .ZN(n12474) );
  OAI211_X1 U14828 ( .C1(n12713), .C2(n12538), .A(n12475), .B(n12474), .ZN(
        P3_U3165) );
  XNOR2_X1 U14829 ( .A(n12476), .B(n12829), .ZN(n12477) );
  XNOR2_X1 U14830 ( .A(n12478), .B(n12477), .ZN(n12483) );
  NAND2_X1 U14831 ( .A1(n12505), .A2(n12819), .ZN(n12480) );
  AND2_X1 U14832 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n14417) );
  AOI21_X1 U14833 ( .B1(n12535), .B2(n12544), .A(n14417), .ZN(n12479) );
  OAI211_X1 U14834 ( .C1(n12812), .C2(n12508), .A(n12480), .B(n12479), .ZN(
        n12481) );
  AOI21_X1 U14835 ( .B1(n12929), .B2(n12521), .A(n12481), .ZN(n12482) );
  OAI21_X1 U14836 ( .B1(n12483), .B2(n12523), .A(n12482), .ZN(P3_U3168) );
  INV_X1 U14837 ( .A(n12484), .ZN(n12486) );
  NOR3_X1 U14838 ( .A1(n6467), .A2(n12486), .A3(n12485), .ZN(n12488) );
  OAI21_X1 U14839 ( .B1(n12488), .B2(n12487), .A(n12528), .ZN(n12492) );
  AOI22_X1 U14840 ( .A1(n12504), .A2(n12530), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12489) );
  OAI21_X1 U14841 ( .B1(n12719), .B2(n12516), .A(n12489), .ZN(n12490) );
  AOI21_X1 U14842 ( .B1(n12723), .B2(n12505), .A(n12490), .ZN(n12491) );
  OAI211_X1 U14843 ( .C1(n12538), .C2(n12493), .A(n12492), .B(n12491), .ZN(
        P3_U3169) );
  XNOR2_X1 U14844 ( .A(n12495), .B(n12494), .ZN(n12500) );
  AOI22_X1 U14845 ( .A1(n12543), .A2(n12535), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12497) );
  NAND2_X1 U14846 ( .A1(n12505), .A2(n12775), .ZN(n12496) );
  OAI211_X1 U14847 ( .C1(n12796), .C2(n12508), .A(n12497), .B(n12496), .ZN(
        n12498) );
  AOI21_X1 U14848 ( .B1(n12774), .B2(n12521), .A(n12498), .ZN(n12499) );
  OAI21_X1 U14849 ( .B1(n12500), .B2(n12523), .A(n12499), .ZN(P3_U3173) );
  INV_X1 U14850 ( .A(n12501), .ZN(n12502) );
  AOI21_X1 U14851 ( .B1(n12758), .B2(n12503), .A(n12502), .ZN(n12512) );
  AOI22_X1 U14852 ( .A1(n12504), .A2(n12535), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12507) );
  NAND2_X1 U14853 ( .A1(n12505), .A2(n12750), .ZN(n12506) );
  OAI211_X1 U14854 ( .C1(n12769), .C2(n12508), .A(n12507), .B(n12506), .ZN(
        n12509) );
  AOI21_X1 U14855 ( .B1(n12510), .B2(n12521), .A(n12509), .ZN(n12511) );
  OAI21_X1 U14856 ( .B1(n12512), .B2(n12523), .A(n12511), .ZN(P3_U3175) );
  XNOR2_X1 U14857 ( .A(n12514), .B(n12513), .ZN(n12524) );
  INV_X1 U14858 ( .A(n12515), .ZN(n12799) );
  NAND2_X1 U14859 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n14431)
         );
  INV_X1 U14860 ( .A(n14431), .ZN(n12518) );
  NOR2_X1 U14861 ( .A1(n12516), .A2(n12796), .ZN(n12517) );
  AOI211_X1 U14862 ( .C1(n12530), .C2(n12545), .A(n12518), .B(n12517), .ZN(
        n12519) );
  OAI21_X1 U14863 ( .B1(n12799), .B2(n12532), .A(n12519), .ZN(n12520) );
  AOI21_X1 U14864 ( .B1(n12925), .B2(n12521), .A(n12520), .ZN(n12522) );
  OAI21_X1 U14865 ( .B1(n12524), .B2(n12523), .A(n12522), .ZN(P3_U3178) );
  OAI21_X1 U14866 ( .B1(n12527), .B2(n12526), .A(n12525), .ZN(n12529) );
  NAND2_X1 U14867 ( .A1(n12529), .A2(n12528), .ZN(n12537) );
  INV_X1 U14868 ( .A(n12691), .ZN(n12533) );
  AOI22_X1 U14869 ( .A1(n12542), .A2(n12530), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12531) );
  OAI21_X1 U14870 ( .B1(n12533), .B2(n12532), .A(n12531), .ZN(n12534) );
  AOI21_X1 U14871 ( .B1(n12535), .B2(n12541), .A(n12534), .ZN(n12536) );
  OAI211_X1 U14872 ( .C1(n7493), .C2(n12538), .A(n12537), .B(n12536), .ZN(
        P3_U3180) );
  MUX2_X1 U14873 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12539), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14874 ( .A(n12540), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12559), .Z(
        P3_U3521) );
  MUX2_X1 U14875 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12541), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14876 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n7491), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14877 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12542), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14878 ( .A(n12758), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12559), .Z(
        P3_U3513) );
  MUX2_X1 U14879 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12543), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14880 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12757), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14881 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n9290), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14882 ( .A(n12544), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12559), .Z(
        P3_U3509) );
  MUX2_X1 U14883 ( .A(n12545), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12559), .Z(
        P3_U3508) );
  MUX2_X1 U14884 ( .A(n12546), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12559), .Z(
        P3_U3507) );
  MUX2_X1 U14885 ( .A(n12547), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12559), .Z(
        P3_U3506) );
  MUX2_X1 U14886 ( .A(n14438), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12559), .Z(
        P3_U3504) );
  MUX2_X1 U14887 ( .A(n12548), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12559), .Z(
        P3_U3503) );
  MUX2_X1 U14888 ( .A(n14436), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12559), .Z(
        P3_U3502) );
  MUX2_X1 U14889 ( .A(n12549), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12559), .Z(
        P3_U3501) );
  MUX2_X1 U14890 ( .A(n12550), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12559), .Z(
        P3_U3500) );
  MUX2_X1 U14891 ( .A(n12551), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12559), .Z(
        P3_U3499) );
  MUX2_X1 U14892 ( .A(n12552), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12559), .Z(
        P3_U3498) );
  MUX2_X1 U14893 ( .A(n12553), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12559), .Z(
        P3_U3497) );
  MUX2_X1 U14894 ( .A(n12554), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12559), .Z(
        P3_U3496) );
  MUX2_X1 U14895 ( .A(n12555), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12559), .Z(
        P3_U3495) );
  MUX2_X1 U14896 ( .A(n12556), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12559), .Z(
        P3_U3494) );
  MUX2_X1 U14897 ( .A(n12557), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12559), .Z(
        P3_U3493) );
  MUX2_X1 U14898 ( .A(n12558), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12559), .Z(
        P3_U3492) );
  MUX2_X1 U14899 ( .A(n12560), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12559), .Z(
        P3_U3491) );
  OAI21_X1 U14900 ( .B1(n12563), .B2(n12562), .A(n12561), .ZN(n12568) );
  OAI21_X1 U14901 ( .B1(n12566), .B2(n12565), .A(n12564), .ZN(n12567) );
  AOI22_X1 U14902 ( .A1(n15035), .A2(n12568), .B1(n14866), .B2(n12567), .ZN(
        n12578) );
  AOI22_X1 U14903 ( .A1(n15030), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n12577) );
  NAND2_X1 U14904 ( .A1(n14992), .A2(n12569), .ZN(n12576) );
  INV_X1 U14905 ( .A(n14882), .ZN(n12574) );
  NOR3_X1 U14906 ( .A1(n12572), .A2(n12571), .A3(n12570), .ZN(n12573) );
  OAI21_X1 U14907 ( .B1(n12574), .B2(n12573), .A(n15037), .ZN(n12575) );
  NAND4_X1 U14908 ( .A1(n12578), .A2(n12577), .A3(n12576), .A4(n12575), .ZN(
        P3_U3184) );
  INV_X1 U14909 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12579) );
  MUX2_X1 U14910 ( .A(n12579), .B(P3_REG2_REG_19__SCAN_IN), .S(n12596), .Z(
        n12597) );
  NAND2_X1 U14911 ( .A1(n15032), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12618) );
  NOR2_X1 U14912 ( .A1(n12603), .A2(n12582), .ZN(n12583) );
  NOR2_X1 U14913 ( .A1(n14934), .A2(n14933), .ZN(n14932) );
  INV_X1 U14914 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n15299) );
  AOI22_X1 U14915 ( .A1(n12641), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n15299), 
        .B2(n14963), .ZN(n14959) );
  NOR2_X1 U14916 ( .A1(n12643), .A2(n12584), .ZN(n12585) );
  INV_X1 U14917 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n14970) );
  INV_X1 U14918 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12586) );
  AOI22_X1 U14919 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n14991), .B1(n14323), 
        .B2(n12586), .ZN(n14986) );
  NOR2_X1 U14920 ( .A1(n12613), .A2(n12587), .ZN(n12588) );
  OAI21_X1 U14921 ( .B1(n15032), .B2(P3_REG2_REG_14__SCAN_IN), .A(n12618), 
        .ZN(n15024) );
  NOR2_X1 U14922 ( .A1(n15025), .A2(n15024), .ZN(n15023) );
  INV_X1 U14923 ( .A(n15023), .ZN(n12589) );
  AND2_X1 U14924 ( .A1(n14376), .A2(n12590), .ZN(n12591) );
  INV_X1 U14925 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14371) );
  XNOR2_X1 U14926 ( .A(n14376), .B(n12590), .ZN(n14370) );
  INV_X1 U14927 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12592) );
  AOI22_X1 U14928 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12650), .B1(n14393), 
        .B2(n12592), .ZN(n14386) );
  NOR2_X1 U14929 ( .A1(n12651), .A2(n12593), .ZN(n12594) );
  INV_X1 U14930 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14405) );
  INV_X1 U14931 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12595) );
  AOI22_X1 U14932 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n14420), .B1(n12634), 
        .B2(n12595), .ZN(n14429) );
  XNOR2_X1 U14933 ( .A(n12596), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12655) );
  MUX2_X1 U14934 ( .A(n12597), .B(n12655), .S(n6436), .Z(n12631) );
  INV_X1 U14935 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12598) );
  MUX2_X1 U14936 ( .A(n14405), .B(n12598), .S(n12628), .Z(n12625) );
  NOR2_X1 U14937 ( .A1(n12625), .A2(n12651), .ZN(n12627) );
  MUX2_X1 U14938 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12628), .Z(n12611) );
  INV_X1 U14939 ( .A(n12611), .ZN(n12612) );
  MUX2_X1 U14940 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12628), .Z(n12609) );
  INV_X1 U14941 ( .A(n12609), .ZN(n12610) );
  MUX2_X1 U14942 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12628), .Z(n12599) );
  INV_X1 U14943 ( .A(n12599), .ZN(n12608) );
  XNOR2_X1 U14944 ( .A(n12599), .B(n12643), .ZN(n14979) );
  MUX2_X1 U14945 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12628), .Z(n12605) );
  OR2_X1 U14946 ( .A1(n12605), .A2(n14963), .ZN(n12607) );
  INV_X1 U14947 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15155) );
  MUX2_X1 U14948 ( .A(n14934), .B(n15155), .S(n12628), .Z(n12604) );
  OR2_X1 U14949 ( .A1(n12604), .A2(n12603), .ZN(n14936) );
  OR2_X1 U14950 ( .A1(n12600), .A2(n12635), .ZN(n12602) );
  NAND2_X1 U14951 ( .A1(n12602), .A2(n12601), .ZN(n14939) );
  AND2_X1 U14952 ( .A1(n12604), .A2(n12603), .ZN(n14935) );
  AOI21_X1 U14953 ( .B1(n14936), .B2(n14939), .A(n14935), .ZN(n14957) );
  XNOR2_X1 U14954 ( .A(n12605), .B(n14963), .ZN(n14956) );
  NOR2_X1 U14955 ( .A1(n14957), .A2(n14956), .ZN(n14955) );
  INV_X1 U14956 ( .A(n14955), .ZN(n12606) );
  XNOR2_X1 U14957 ( .A(n12609), .B(n14991), .ZN(n15001) );
  OAI21_X1 U14958 ( .B1(n14991), .B2(n12610), .A(n15000), .ZN(n15016) );
  XNOR2_X1 U14959 ( .A(n12611), .B(n15012), .ZN(n15017) );
  INV_X1 U14960 ( .A(n15024), .ZN(n12617) );
  INV_X1 U14961 ( .A(n15032), .ZN(n12616) );
  INV_X1 U14962 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12615) );
  NAND2_X1 U14963 ( .A1(n15032), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12647) );
  INV_X1 U14964 ( .A(n12647), .ZN(n12614) );
  AOI21_X1 U14965 ( .B1(n12616), .B2(n12615), .A(n12614), .ZN(n15028) );
  MUX2_X1 U14966 ( .A(n12617), .B(n15028), .S(n12628), .Z(n15039) );
  MUX2_X1 U14967 ( .A(n12618), .B(n12647), .S(n6436), .Z(n12619) );
  INV_X1 U14968 ( .A(n12620), .ZN(n12622) );
  INV_X1 U14969 ( .A(n14376), .ZN(n12621) );
  XNOR2_X1 U14970 ( .A(n12620), .B(n14376), .ZN(n14380) );
  MUX2_X1 U14971 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n6436), .Z(n14381) );
  NOR2_X1 U14972 ( .A1(n14380), .A2(n14381), .ZN(n14379) );
  MUX2_X1 U14973 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n6436), .Z(n12623) );
  AND2_X1 U14974 ( .A1(n12623), .A2(n14393), .ZN(n14396) );
  INV_X1 U14975 ( .A(n12623), .ZN(n12624) );
  AOI21_X1 U14976 ( .B1(n12651), .B2(n12625), .A(n12627), .ZN(n12626) );
  INV_X1 U14977 ( .A(n12626), .ZN(n14411) );
  XNOR2_X1 U14978 ( .A(n12634), .B(n12629), .ZN(n14426) );
  INV_X1 U14979 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12654) );
  MUX2_X1 U14980 ( .A(n12595), .B(n12654), .S(n12628), .Z(n14425) );
  NAND2_X1 U14981 ( .A1(n14426), .A2(n14425), .ZN(n14424) );
  NAND2_X1 U14982 ( .A1(n14420), .A2(n12629), .ZN(n12630) );
  AOI21_X1 U14983 ( .B1(n15030), .B2(P3_ADDR_REG_19__SCAN_IN), .A(n12632), 
        .ZN(n12633) );
  AOI22_X1 U14984 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n12634), .B1(n14420), 
        .B2(n12654), .ZN(n14423) );
  INV_X1 U14985 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12888) );
  AOI22_X1 U14986 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n14393), .B1(n12650), 
        .B2(n12888), .ZN(n14390) );
  INV_X1 U14987 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14467) );
  AOI22_X1 U14988 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n14323), .B1(n14991), 
        .B2(n14467), .ZN(n14990) );
  AOI22_X1 U14989 ( .A1(n12641), .A2(n12640), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n14963), .ZN(n14952) );
  NAND2_X1 U14990 ( .A1(n12635), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n12637) );
  NAND2_X1 U14991 ( .A1(n12637), .A2(n12636), .ZN(n12638) );
  NAND2_X1 U14992 ( .A1(n14940), .A2(n12638), .ZN(n12639) );
  XOR2_X1 U14993 ( .A(n12638), .B(n14940), .Z(n14945) );
  NAND2_X1 U14994 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n14945), .ZN(n14944) );
  NAND2_X1 U14995 ( .A1(n12639), .A2(n14944), .ZN(n14951) );
  NAND2_X1 U14996 ( .A1(n14952), .A2(n14951), .ZN(n14950) );
  NAND2_X1 U14997 ( .A1(n14975), .A2(n12642), .ZN(n12644) );
  XNOR2_X1 U14998 ( .A(n12643), .B(n12642), .ZN(n14972) );
  NAND2_X1 U14999 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n14972), .ZN(n14971) );
  NAND2_X1 U15000 ( .A1(n12644), .A2(n14971), .ZN(n14989) );
  NAND2_X1 U15001 ( .A1(n14990), .A2(n14989), .ZN(n14988) );
  OAI21_X1 U15002 ( .B1(n14991), .B2(n14467), .A(n14988), .ZN(n12645) );
  NAND2_X1 U15003 ( .A1(n15012), .A2(n12645), .ZN(n12646) );
  NAND2_X1 U15004 ( .A1(n12646), .A2(n15008), .ZN(n15027) );
  NAND2_X1 U15005 ( .A1(n15028), .A2(n15027), .ZN(n15026) );
  NAND2_X1 U15006 ( .A1(n14376), .A2(n12648), .ZN(n12649) );
  NAND2_X1 U15007 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n14373), .ZN(n14372) );
  NAND2_X1 U15008 ( .A1(n12649), .A2(n14372), .ZN(n14389) );
  NAND2_X1 U15009 ( .A1(n14390), .A2(n14389), .ZN(n14388) );
  NAND2_X1 U15010 ( .A1(n14413), .A2(n12652), .ZN(n12653) );
  XNOR2_X1 U15011 ( .A(n12652), .B(n12651), .ZN(n14407) );
  NAND2_X1 U15012 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n14407), .ZN(n14406) );
  NAND2_X1 U15013 ( .A1(n12653), .A2(n14406), .ZN(n14422) );
  XNOR2_X1 U15014 ( .A(n12656), .B(n12655), .ZN(n12657) );
  NOR2_X1 U15015 ( .A1(n12657), .A2(n14912), .ZN(n12658) );
  OAI21_X1 U15016 ( .B1(n12661), .B2(n15043), .A(n12660), .ZN(P3_U3201) );
  AOI21_X1 U15017 ( .B1(n15075), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12662), 
        .ZN(n12663) );
  OAI21_X1 U15018 ( .B1(n12664), .B2(n12835), .A(n12663), .ZN(P3_U3203) );
  INV_X1 U15019 ( .A(n12665), .ZN(n12671) );
  AOI22_X1 U15020 ( .A1(n12666), .A2(n15071), .B1(n15075), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12667) );
  OAI21_X1 U15021 ( .B1(n12897), .B2(n12835), .A(n12667), .ZN(n12668) );
  AOI21_X1 U15022 ( .B1(n12669), .B2(n14445), .A(n12668), .ZN(n12670) );
  OAI21_X1 U15023 ( .B1(n12671), .B2(n15075), .A(n12670), .ZN(P3_U3205) );
  OAI222_X1 U15024 ( .A1(n15087), .A2(n12674), .B1(n15084), .B2(n12703), .C1(
        n15049), .C2(n12673), .ZN(n12675) );
  INV_X1 U15025 ( .A(n12675), .ZN(n12842) );
  INV_X1 U15026 ( .A(n12676), .ZN(n12677) );
  OAI21_X1 U15027 ( .B1(n12679), .B2(n12678), .A(n12677), .ZN(n12840) );
  AOI22_X1 U15028 ( .A1(n12680), .A2(n15071), .B1(n15075), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12681) );
  OAI21_X1 U15029 ( .B1(n12682), .B2(n12835), .A(n12681), .ZN(n12683) );
  AOI21_X1 U15030 ( .B1(n12840), .B2(n14445), .A(n12683), .ZN(n12684) );
  OAI21_X1 U15031 ( .B1(n12842), .B2(n15075), .A(n12684), .ZN(P3_U3206) );
  INV_X1 U15032 ( .A(n12688), .ZN(n12686) );
  XNOR2_X1 U15033 ( .A(n12686), .B(n12685), .ZN(n12844) );
  INV_X1 U15034 ( .A(n12844), .ZN(n12698) );
  XOR2_X1 U15035 ( .A(n12688), .B(n12687), .Z(n12689) );
  OAI222_X1 U15036 ( .A1(n15087), .A2(n12690), .B1(n15084), .B2(n12719), .C1(
        n12689), .C2(n15049), .ZN(n12843) );
  NAND2_X1 U15037 ( .A1(n12843), .A2(n15096), .ZN(n12697) );
  NAND2_X1 U15038 ( .A1(n12691), .A2(n15071), .ZN(n12692) );
  OAI21_X1 U15039 ( .B1(n15096), .B2(n12693), .A(n12692), .ZN(n12694) );
  AOI21_X1 U15040 ( .B1(n12695), .B2(n12801), .A(n12694), .ZN(n12696) );
  OAI211_X1 U15041 ( .C1(n12698), .C2(n12805), .A(n12697), .B(n12696), .ZN(
        P3_U3207) );
  INV_X1 U15042 ( .A(n12699), .ZN(n12701) );
  AOI21_X1 U15043 ( .B1(n12701), .B2(n12700), .A(n15049), .ZN(n12706) );
  OAI22_X1 U15044 ( .A1(n12703), .A2(n15087), .B1(n12702), .B2(n15084), .ZN(
        n12704) );
  AOI21_X1 U15045 ( .B1(n12706), .B2(n12705), .A(n12704), .ZN(n12850) );
  NAND3_X1 U15046 ( .A1(n12726), .A2(n12708), .A3(n12707), .ZN(n12709) );
  NAND2_X1 U15047 ( .A1(n12710), .A2(n12709), .ZN(n12848) );
  AOI22_X1 U15048 ( .A1(n12711), .A2(n15071), .B1(n15075), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12712) );
  OAI21_X1 U15049 ( .B1(n12713), .B2(n12835), .A(n12712), .ZN(n12714) );
  AOI21_X1 U15050 ( .B1(n12848), .B2(n14445), .A(n12714), .ZN(n12715) );
  OAI21_X1 U15051 ( .B1(n12850), .B2(n15075), .A(n12715), .ZN(P3_U3208) );
  INV_X1 U15052 ( .A(n12716), .ZN(n12718) );
  INV_X1 U15053 ( .A(n12728), .ZN(n12717) );
  AOI21_X1 U15054 ( .B1(n12718), .B2(n12717), .A(n15049), .ZN(n12722) );
  OAI22_X1 U15055 ( .A1(n12719), .A2(n15087), .B1(n12747), .B2(n15084), .ZN(
        n12720) );
  AOI21_X1 U15056 ( .B1(n12722), .B2(n12721), .A(n12720), .ZN(n12853) );
  INV_X1 U15057 ( .A(n12723), .ZN(n12725) );
  OAI22_X1 U15058 ( .A1(n12725), .A2(n15081), .B1(n15096), .B2(n12724), .ZN(
        n12730) );
  AOI21_X1 U15059 ( .B1(n12728), .B2(n12727), .A(n9409), .ZN(n12854) );
  NOR2_X1 U15060 ( .A1(n12854), .A2(n12805), .ZN(n12729) );
  AOI211_X1 U15061 ( .C1(n12801), .C2(n12851), .A(n12730), .B(n12729), .ZN(
        n12731) );
  OAI21_X1 U15062 ( .B1(n12853), .B2(n15075), .A(n12731), .ZN(P3_U3209) );
  OAI211_X1 U15063 ( .C1(n12733), .C2(n12737), .A(n12732), .B(n15089), .ZN(
        n12736) );
  AOI22_X1 U15064 ( .A1(n12734), .A2(n14437), .B1(n14435), .B2(n12758), .ZN(
        n12735) );
  NAND2_X1 U15065 ( .A1(n12736), .A2(n12735), .ZN(n12855) );
  INV_X1 U15066 ( .A(n12855), .ZN(n12743) );
  XNOR2_X1 U15067 ( .A(n12738), .B(n12737), .ZN(n12856) );
  AOI22_X1 U15068 ( .A1(n15075), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15071), 
        .B2(n12739), .ZN(n12740) );
  OAI21_X1 U15069 ( .B1(n12907), .B2(n12835), .A(n12740), .ZN(n12741) );
  AOI21_X1 U15070 ( .B1(n12856), .B2(n14445), .A(n12741), .ZN(n12742) );
  OAI21_X1 U15071 ( .B1(n12743), .B2(n15075), .A(n12742), .ZN(P3_U3210) );
  XNOR2_X1 U15072 ( .A(n12745), .B(n12744), .ZN(n12746) );
  OAI222_X1 U15073 ( .A1(n15084), .A2(n12769), .B1(n15087), .B2(n12747), .C1(
        n15049), .C2(n12746), .ZN(n12858) );
  INV_X1 U15074 ( .A(n12858), .ZN(n12754) );
  XNOR2_X1 U15075 ( .A(n12749), .B(n12748), .ZN(n12859) );
  AOI22_X1 U15076 ( .A1(n15075), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15071), 
        .B2(n12750), .ZN(n12751) );
  OAI21_X1 U15077 ( .B1(n12911), .B2(n12835), .A(n12751), .ZN(n12752) );
  AOI21_X1 U15078 ( .B1(n12859), .B2(n14445), .A(n12752), .ZN(n12753) );
  OAI21_X1 U15079 ( .B1(n12754), .B2(n15075), .A(n12753), .ZN(P3_U3211) );
  OAI21_X1 U15080 ( .B1(n12756), .B2(n12760), .A(n12755), .ZN(n12759) );
  AOI222_X1 U15081 ( .A1(n15089), .A2(n12759), .B1(n12758), .B2(n14437), .C1(
        n12757), .C2(n14435), .ZN(n12862) );
  XNOR2_X1 U15082 ( .A(n12761), .B(n12760), .ZN(n12864) );
  AOI22_X1 U15083 ( .A1(n15075), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15071), 
        .B2(n12763), .ZN(n12764) );
  OAI21_X1 U15084 ( .B1(n6818), .B2(n12835), .A(n12764), .ZN(n12765) );
  AOI21_X1 U15085 ( .B1(n12864), .B2(n14445), .A(n12765), .ZN(n12766) );
  OAI21_X1 U15086 ( .B1(n12862), .B2(n15075), .A(n12766), .ZN(P3_U3212) );
  XNOR2_X1 U15087 ( .A(n12767), .B(n12773), .ZN(n12768) );
  OAI222_X1 U15088 ( .A1(n15087), .A2(n12769), .B1(n15084), .B2(n12796), .C1(
        n12768), .C2(n15049), .ZN(n12867) );
  INV_X1 U15089 ( .A(n12867), .ZN(n12779) );
  INV_X1 U15090 ( .A(n12770), .ZN(n12771) );
  AOI21_X1 U15091 ( .B1(n12773), .B2(n12772), .A(n12771), .ZN(n12868) );
  INV_X1 U15092 ( .A(n12774), .ZN(n12918) );
  AOI22_X1 U15093 ( .A1(n15075), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15071), 
        .B2(n12775), .ZN(n12776) );
  OAI21_X1 U15094 ( .B1(n12918), .B2(n12835), .A(n12776), .ZN(n12777) );
  AOI21_X1 U15095 ( .B1(n12868), .B2(n14445), .A(n12777), .ZN(n12778) );
  OAI21_X1 U15096 ( .B1(n12779), .B2(n15075), .A(n12778), .ZN(P3_U3213) );
  OAI211_X1 U15097 ( .C1(n12781), .C2(n12786), .A(n12780), .B(n15089), .ZN(
        n12785) );
  OAI22_X1 U15098 ( .A1(n12782), .A2(n15087), .B1(n12813), .B2(n15084), .ZN(
        n12783) );
  INV_X1 U15099 ( .A(n12783), .ZN(n12784) );
  XNOR2_X1 U15100 ( .A(n12787), .B(n12786), .ZN(n12870) );
  AOI22_X1 U15101 ( .A1(n15075), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15071), 
        .B2(n12788), .ZN(n12789) );
  OAI21_X1 U15102 ( .B1(n12922), .B2(n12835), .A(n12789), .ZN(n12790) );
  AOI21_X1 U15103 ( .B1(n12870), .B2(n14445), .A(n12790), .ZN(n12791) );
  OAI21_X1 U15104 ( .B1(n12872), .B2(n15075), .A(n12791), .ZN(P3_U3214) );
  NAND2_X1 U15105 ( .A1(n12794), .A2(n12793), .ZN(n12795) );
  NAND2_X1 U15106 ( .A1(n12792), .A2(n12795), .ZN(n12798) );
  OAI22_X1 U15107 ( .A1(n12796), .A2(n15087), .B1(n12829), .B2(n15084), .ZN(
        n12797) );
  AOI21_X1 U15108 ( .B1(n12798), .B2(n15089), .A(n12797), .ZN(n12877) );
  OAI22_X1 U15109 ( .A1(n15096), .A2(n12595), .B1(n12799), .B2(n15081), .ZN(
        n12800) );
  AOI21_X1 U15110 ( .B1(n12925), .B2(n12801), .A(n12800), .ZN(n12807) );
  NAND2_X1 U15111 ( .A1(n12802), .A2(n9272), .ZN(n12803) );
  NAND2_X1 U15112 ( .A1(n12804), .A2(n12803), .ZN(n12875) );
  OR2_X1 U15113 ( .A1(n12875), .A2(n12805), .ZN(n12806) );
  OAI211_X1 U15114 ( .C1(n12877), .C2(n15075), .A(n12807), .B(n12806), .ZN(
        P3_U3215) );
  AND2_X1 U15115 ( .A1(n12825), .A2(n12808), .ZN(n12811) );
  OAI211_X1 U15116 ( .C1(n12811), .C2(n12810), .A(n12809), .B(n15089), .ZN(
        n12816) );
  OAI22_X1 U15117 ( .A1(n15087), .A2(n12813), .B1(n12812), .B2(n15084), .ZN(
        n12814) );
  INV_X1 U15118 ( .A(n12814), .ZN(n12815) );
  XNOR2_X1 U15119 ( .A(n12818), .B(n12817), .ZN(n12880) );
  INV_X1 U15120 ( .A(n12929), .ZN(n12821) );
  AOI22_X1 U15121 ( .A1(n15075), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15071), 
        .B2(n12819), .ZN(n12820) );
  OAI21_X1 U15122 ( .B1(n12821), .B2(n12835), .A(n12820), .ZN(n12822) );
  AOI21_X1 U15123 ( .B1(n12880), .B2(n14445), .A(n12822), .ZN(n12823) );
  OAI21_X1 U15124 ( .B1(n12882), .B2(n15075), .A(n12823), .ZN(P3_U3216) );
  INV_X1 U15125 ( .A(n12825), .ZN(n12826) );
  AOI21_X1 U15126 ( .B1(n12831), .B2(n12824), .A(n12826), .ZN(n12827) );
  OAI222_X1 U15127 ( .A1(n15087), .A2(n12829), .B1(n15084), .B2(n12828), .C1(
        n15049), .C2(n12827), .ZN(n12886) );
  INV_X1 U15128 ( .A(n12886), .ZN(n12838) );
  XNOR2_X1 U15129 ( .A(n12830), .B(n12831), .ZN(n12887) );
  INV_X1 U15130 ( .A(n12832), .ZN(n12935) );
  AOI22_X1 U15131 ( .A1(n15075), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15071), 
        .B2(n12833), .ZN(n12834) );
  OAI21_X1 U15132 ( .B1(n12935), .B2(n12835), .A(n12834), .ZN(n12836) );
  AOI21_X1 U15133 ( .B1(n12887), .B2(n14445), .A(n12836), .ZN(n12837) );
  OAI21_X1 U15134 ( .B1(n12838), .B2(n15075), .A(n12837), .ZN(P3_U3217) );
  AOI22_X1 U15135 ( .A1(n12840), .A2(n15101), .B1(n15078), .B2(n12839), .ZN(
        n12841) );
  NAND2_X1 U15136 ( .A1(n12842), .A2(n12841), .ZN(n12898) );
  MUX2_X1 U15137 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n12898), .S(n15157), .Z(
        P3_U3486) );
  INV_X1 U15138 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12845) );
  AOI21_X1 U15139 ( .B1(n12844), .B2(n15101), .A(n12843), .ZN(n12899) );
  MUX2_X1 U15140 ( .A(n12845), .B(n12899), .S(n15157), .Z(n12846) );
  OAI21_X1 U15141 ( .B1(n7493), .B2(n12894), .A(n12846), .ZN(P3_U3485) );
  AOI22_X1 U15142 ( .A1(n12848), .A2(n15101), .B1(n15078), .B2(n12847), .ZN(
        n12849) );
  NAND2_X1 U15143 ( .A1(n12850), .A2(n12849), .ZN(n12902) );
  MUX2_X1 U15144 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n12902), .S(n15157), .Z(
        P3_U3484) );
  NAND2_X1 U15145 ( .A1(n12851), .A2(n15078), .ZN(n12852) );
  OAI211_X1 U15146 ( .C1(n14458), .C2(n12854), .A(n12853), .B(n12852), .ZN(
        n12903) );
  MUX2_X1 U15147 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n12903), .S(n15157), .Z(
        P3_U3483) );
  INV_X1 U15148 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n15304) );
  AOI21_X1 U15149 ( .B1(n12856), .B2(n15101), .A(n12855), .ZN(n12904) );
  MUX2_X1 U15150 ( .A(n15304), .B(n12904), .S(n15157), .Z(n12857) );
  OAI21_X1 U15151 ( .B1(n12907), .B2(n12894), .A(n12857), .ZN(P3_U3482) );
  INV_X1 U15152 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12860) );
  AOI21_X1 U15153 ( .B1(n15101), .B2(n12859), .A(n12858), .ZN(n12908) );
  MUX2_X1 U15154 ( .A(n12860), .B(n12908), .S(n15157), .Z(n12861) );
  OAI21_X1 U15155 ( .B1(n12911), .B2(n12894), .A(n12861), .ZN(P3_U3481) );
  INV_X1 U15156 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12865) );
  INV_X1 U15157 ( .A(n12862), .ZN(n12863) );
  AOI21_X1 U15158 ( .B1(n15101), .B2(n12864), .A(n12863), .ZN(n12912) );
  MUX2_X1 U15159 ( .A(n12865), .B(n12912), .S(n15157), .Z(n12866) );
  OAI21_X1 U15160 ( .B1(n6818), .B2(n12894), .A(n12866), .ZN(P3_U3480) );
  INV_X1 U15161 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n15282) );
  AOI21_X1 U15162 ( .B1(n12868), .B2(n15101), .A(n12867), .ZN(n12915) );
  MUX2_X1 U15163 ( .A(n15282), .B(n12915), .S(n15157), .Z(n12869) );
  OAI21_X1 U15164 ( .B1(n12918), .B2(n12894), .A(n12869), .ZN(P3_U3479) );
  NAND2_X1 U15165 ( .A1(n12870), .A2(n15101), .ZN(n12871) );
  NAND2_X1 U15166 ( .A1(n12872), .A2(n12871), .ZN(n12919) );
  MUX2_X1 U15167 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n12919), .S(n15157), .Z(
        n12873) );
  INV_X1 U15168 ( .A(n12873), .ZN(n12874) );
  OAI21_X1 U15169 ( .B1(n12922), .B2(n12894), .A(n12874), .ZN(P3_U3478) );
  OR2_X1 U15170 ( .A1(n12875), .A2(n14458), .ZN(n12876) );
  NAND2_X1 U15171 ( .A1(n12877), .A2(n12876), .ZN(n12923) );
  MUX2_X1 U15172 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n12923), .S(n15157), .Z(
        n12878) );
  AOI21_X1 U15173 ( .B1(n12884), .B2(n12925), .A(n12878), .ZN(n12879) );
  INV_X1 U15174 ( .A(n12879), .ZN(P3_U3477) );
  NAND2_X1 U15175 ( .A1(n12880), .A2(n15101), .ZN(n12881) );
  NAND2_X1 U15176 ( .A1(n12882), .A2(n12881), .ZN(n12927) );
  MUX2_X1 U15177 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12927), .S(n15157), .Z(
        n12883) );
  AOI21_X1 U15178 ( .B1(n12884), .B2(n12929), .A(n12883), .ZN(n12885) );
  INV_X1 U15179 ( .A(n12885), .ZN(P3_U3476) );
  AOI21_X1 U15180 ( .B1(n12887), .B2(n15101), .A(n12886), .ZN(n12932) );
  MUX2_X1 U15181 ( .A(n12888), .B(n12932), .S(n15157), .Z(n12889) );
  OAI21_X1 U15182 ( .B1(n12935), .B2(n12894), .A(n12889), .ZN(P3_U3475) );
  INV_X1 U15183 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12892) );
  AOI21_X1 U15184 ( .B1(n12891), .B2(n15101), .A(n12890), .ZN(n12936) );
  MUX2_X1 U15185 ( .A(n12892), .B(n12936), .S(n15157), .Z(n12893) );
  OAI21_X1 U15186 ( .B1(n12940), .B2(n12894), .A(n12893), .ZN(P3_U3474) );
  INV_X1 U15187 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n12896) );
  MUX2_X1 U15188 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n12898), .S(n15141), .Z(
        P3_U3454) );
  INV_X1 U15189 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12900) );
  MUX2_X1 U15190 ( .A(n12900), .B(n12899), .S(n15141), .Z(n12901) );
  OAI21_X1 U15191 ( .B1(n7493), .B2(n12939), .A(n12901), .ZN(P3_U3453) );
  MUX2_X1 U15192 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n12902), .S(n15141), .Z(
        P3_U3452) );
  MUX2_X1 U15193 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n12903), .S(n15141), .Z(
        P3_U3451) );
  INV_X1 U15194 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12905) );
  MUX2_X1 U15195 ( .A(n12905), .B(n12904), .S(n15141), .Z(n12906) );
  OAI21_X1 U15196 ( .B1(n12907), .B2(n12939), .A(n12906), .ZN(P3_U3450) );
  INV_X1 U15197 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12909) );
  MUX2_X1 U15198 ( .A(n12909), .B(n12908), .S(n15141), .Z(n12910) );
  OAI21_X1 U15199 ( .B1(n12911), .B2(n12939), .A(n12910), .ZN(P3_U3449) );
  INV_X1 U15200 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12913) );
  MUX2_X1 U15201 ( .A(n12913), .B(n12912), .S(n15141), .Z(n12914) );
  OAI21_X1 U15202 ( .B1(n6818), .B2(n12939), .A(n12914), .ZN(P3_U3448) );
  INV_X1 U15203 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12916) );
  MUX2_X1 U15204 ( .A(n12916), .B(n12915), .S(n15141), .Z(n12917) );
  OAI21_X1 U15205 ( .B1(n12918), .B2(n12939), .A(n12917), .ZN(P3_U3447) );
  MUX2_X1 U15206 ( .A(n12919), .B(P3_REG0_REG_19__SCAN_IN), .S(n15142), .Z(
        n12920) );
  INV_X1 U15207 ( .A(n12920), .ZN(n12921) );
  OAI21_X1 U15208 ( .B1(n12922), .B2(n12939), .A(n12921), .ZN(P3_U3446) );
  INV_X1 U15209 ( .A(n12939), .ZN(n12930) );
  MUX2_X1 U15210 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n12923), .S(n15141), .Z(
        n12924) );
  AOI21_X1 U15211 ( .B1(n12930), .B2(n12925), .A(n12924), .ZN(n12926) );
  INV_X1 U15212 ( .A(n12926), .ZN(P3_U3444) );
  MUX2_X1 U15213 ( .A(n12927), .B(P3_REG0_REG_17__SCAN_IN), .S(n15142), .Z(
        n12928) );
  AOI21_X1 U15214 ( .B1(n12930), .B2(n12929), .A(n12928), .ZN(n12931) );
  INV_X1 U15215 ( .A(n12931), .ZN(P3_U3441) );
  INV_X1 U15216 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12933) );
  MUX2_X1 U15217 ( .A(n12933), .B(n12932), .S(n15141), .Z(n12934) );
  OAI21_X1 U15218 ( .B1(n12935), .B2(n12939), .A(n12934), .ZN(P3_U3438) );
  INV_X1 U15219 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12937) );
  MUX2_X1 U15220 ( .A(n12937), .B(n12936), .S(n15141), .Z(n12938) );
  OAI21_X1 U15221 ( .B1(n12940), .B2(n12939), .A(n12938), .ZN(P3_U3435) );
  MUX2_X1 U15222 ( .A(n12942), .B(P3_D_REG_0__SCAN_IN), .S(n12941), .Z(
        P3_U3376) );
  NAND2_X1 U15223 ( .A1(n12943), .A2(n14320), .ZN(n12946) );
  OR4_X1 U15224 ( .A1(n12944), .A2(P3_IR_REG_30__SCAN_IN), .A3(n9225), .A4(
        P3_U3151), .ZN(n12945) );
  OAI211_X1 U15225 ( .C1(n12962), .C2(n12947), .A(n12946), .B(n12945), .ZN(
        P3_U3264) );
  OAI222_X1 U15226 ( .A1(P3_U3151), .A2(n12950), .B1(n12960), .B2(n12949), 
        .C1(n12948), .C2(n12962), .ZN(P3_U3265) );
  INV_X1 U15227 ( .A(n12951), .ZN(n12953) );
  OAI222_X1 U15228 ( .A1(n12962), .A2(n12954), .B1(n12960), .B2(n12953), .C1(
        P3_U3151), .C2(n12952), .ZN(P3_U3266) );
  INV_X1 U15229 ( .A(n12955), .ZN(n12956) );
  OAI222_X1 U15230 ( .A1(n12962), .A2(n12957), .B1(P3_U3151), .B2(n9384), .C1(
        n12960), .C2(n12956), .ZN(P3_U3267) );
  INV_X1 U15231 ( .A(n12958), .ZN(n12959) );
  OAI222_X1 U15232 ( .A1(P3_U3151), .A2(n6679), .B1(n12962), .B2(n12961), .C1(
        n12960), .C2(n12959), .ZN(P3_U3269) );
  XOR2_X1 U15233 ( .A(n12965), .B(n12964), .Z(n12971) );
  AND2_X1 U15234 ( .A1(n13122), .A2(n13050), .ZN(n12966) );
  AOI21_X1 U15235 ( .B1(n13120), .B2(n13061), .A(n12966), .ZN(n13515) );
  INV_X1 U15236 ( .A(n12967), .ZN(n13344) );
  AOI22_X1 U15237 ( .A1(n13344), .A2(n13110), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12968) );
  OAI21_X1 U15238 ( .B1(n13515), .B2(n13108), .A(n12968), .ZN(n12969) );
  AOI21_X1 U15239 ( .B1(n13587), .B2(n13081), .A(n12969), .ZN(n12970) );
  OAI21_X1 U15240 ( .B1(n12971), .B2(n13070), .A(n12970), .ZN(P2_U3188) );
  NAND2_X1 U15241 ( .A1(n12972), .A2(n12973), .ZN(n13071) );
  XNOR2_X1 U15242 ( .A(n12975), .B(n12974), .ZN(n13072) );
  NOR2_X1 U15243 ( .A1(n13071), .A2(n13072), .ZN(n13069) );
  NOR2_X1 U15244 ( .A1(n13069), .A2(n12976), .ZN(n12980) );
  NAND2_X1 U15245 ( .A1(n12978), .A2(n12977), .ZN(n12979) );
  XNOR2_X1 U15246 ( .A(n12980), .B(n12979), .ZN(n12985) );
  AOI22_X1 U15247 ( .A1(n13124), .A2(n13061), .B1(n13050), .B2(n12981), .ZN(
        n13402) );
  NAND2_X1 U15248 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13252)
         );
  NAND2_X1 U15249 ( .A1(n13110), .A2(n13405), .ZN(n12982) );
  OAI211_X1 U15250 ( .C1(n13402), .C2(n13108), .A(n13252), .B(n12982), .ZN(
        n12983) );
  AOI21_X1 U15251 ( .B1(n13537), .B2(n13081), .A(n12983), .ZN(n12984) );
  OAI21_X1 U15252 ( .B1(n12985), .B2(n13070), .A(n12984), .ZN(P2_U3191) );
  INV_X1 U15253 ( .A(n12986), .ZN(n12987) );
  NAND2_X1 U15254 ( .A1(n13117), .A2(n13460), .ZN(n12989) );
  XOR2_X1 U15255 ( .A(n12990), .B(n12989), .Z(n12991) );
  XNOR2_X1 U15256 ( .A(n13489), .B(n12991), .ZN(n12992) );
  NAND2_X1 U15257 ( .A1(n13118), .A2(n13050), .ZN(n12995) );
  OR2_X1 U15258 ( .A1(n12993), .A2(n13094), .ZN(n12994) );
  AND2_X1 U15259 ( .A1(n12995), .A2(n12994), .ZN(n13268) );
  AOI22_X1 U15260 ( .A1(n13263), .A2(n13110), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12996) );
  OAI21_X1 U15261 ( .B1(n13268), .B2(n13108), .A(n12996), .ZN(n12997) );
  AOI21_X1 U15262 ( .B1(n13489), .B2(n13081), .A(n12997), .ZN(n12998) );
  AOI211_X1 U15263 ( .C1(n13001), .C2(n13000), .A(n13070), .B(n12999), .ZN(
        n13002) );
  INV_X1 U15264 ( .A(n13002), .ZN(n13006) );
  AOI22_X1 U15265 ( .A1(n13122), .A2(n13061), .B1(n13050), .B2(n13124), .ZN(
        n13380) );
  OAI22_X1 U15266 ( .A1(n13380), .A2(n13108), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13003), .ZN(n13004) );
  AOI21_X1 U15267 ( .B1(n13374), .B2(n13110), .A(n13004), .ZN(n13005) );
  OAI211_X1 U15268 ( .C1(n13376), .C2(n13114), .A(n13006), .B(n13005), .ZN(
        P2_U3195) );
  AND2_X1 U15269 ( .A1(n13120), .A2(n13050), .ZN(n13007) );
  AOI21_X1 U15270 ( .B1(n13119), .B2(n13061), .A(n13007), .ZN(n13313) );
  AOI22_X1 U15271 ( .A1(n13318), .A2(n13110), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13008) );
  OAI21_X1 U15272 ( .B1(n13313), .B2(n13108), .A(n13008), .ZN(n13013) );
  AOI211_X1 U15273 ( .C1(n13009), .C2(n13011), .A(n13070), .B(n13010), .ZN(
        n13012) );
  AOI21_X1 U15274 ( .B1(n13016), .B2(n13015), .A(n13014), .ZN(n13022) );
  NOR2_X1 U15275 ( .A1(n13097), .A2(n13456), .ZN(n13020) );
  AND2_X1 U15276 ( .A1(n13128), .A2(n13050), .ZN(n13017) );
  AOI21_X1 U15277 ( .B1(n13126), .B2(n13061), .A(n13017), .ZN(n13453) );
  OAI21_X1 U15278 ( .B1(n13108), .B2(n13453), .A(n13018), .ZN(n13019) );
  AOI211_X1 U15279 ( .C1(n13551), .C2(n13081), .A(n13020), .B(n13019), .ZN(
        n13021) );
  OAI21_X1 U15280 ( .B1(n13022), .B2(n13070), .A(n13021), .ZN(P2_U3198) );
  INV_X1 U15281 ( .A(n12972), .ZN(n13026) );
  NOR3_X1 U15282 ( .A1(n13014), .A2(n13024), .A3(n13023), .ZN(n13025) );
  OAI21_X1 U15283 ( .B1(n13026), .B2(n13025), .A(n9789), .ZN(n13034) );
  INV_X1 U15284 ( .A(n13438), .ZN(n13032) );
  OAI22_X1 U15285 ( .A1(n13028), .A2(n13094), .B1(n13027), .B2(n13092), .ZN(
        n13029) );
  INV_X1 U15286 ( .A(n13029), .ZN(n13433) );
  OAI22_X1 U15287 ( .A1(n13433), .A2(n13108), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13030), .ZN(n13031) );
  AOI21_X1 U15288 ( .B1(n13032), .B2(n13110), .A(n13031), .ZN(n13033) );
  OAI211_X1 U15289 ( .C1(n13035), .C2(n13114), .A(n13034), .B(n13033), .ZN(
        P2_U3200) );
  AOI211_X1 U15290 ( .C1(n13038), .C2(n13037), .A(n13070), .B(n13036), .ZN(
        n13039) );
  INV_X1 U15291 ( .A(n13039), .ZN(n13044) );
  OAI22_X1 U15292 ( .A1(n13093), .A2(n13094), .B1(n13040), .B2(n13092), .ZN(
        n13325) );
  OAI22_X1 U15293 ( .A1(n13332), .A2(n13097), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13041), .ZN(n13042) );
  AOI21_X1 U15294 ( .B1(n13325), .B2(n13099), .A(n13042), .ZN(n13043) );
  OAI211_X1 U15295 ( .C1(n13584), .C2(n13114), .A(n13044), .B(n13043), .ZN(
        P2_U3201) );
  INV_X1 U15296 ( .A(n13046), .ZN(n13047) );
  NOR2_X1 U15297 ( .A1(n13048), .A2(n13047), .ZN(n13049) );
  XNOR2_X1 U15298 ( .A(n13045), .B(n13049), .ZN(n13055) );
  AOI22_X1 U15299 ( .A1(n13123), .A2(n13061), .B1(n13050), .B2(n13125), .ZN(
        n13394) );
  INV_X1 U15300 ( .A(n13394), .ZN(n13051) );
  AOI22_X1 U15301 ( .A1(n13051), .A2(n13099), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13052) );
  OAI21_X1 U15302 ( .B1(n13389), .B2(n13097), .A(n13052), .ZN(n13053) );
  AOI21_X1 U15303 ( .B1(n13387), .B2(n13081), .A(n13053), .ZN(n13054) );
  OAI21_X1 U15304 ( .B1(n13055), .B2(n13070), .A(n13054), .ZN(P2_U3205) );
  OAI211_X1 U15305 ( .C1(n13058), .C2(n13057), .A(n13056), .B(n9789), .ZN(
        n13065) );
  NOR2_X1 U15306 ( .A1(n13361), .A2(n13097), .ZN(n13063) );
  NOR2_X1 U15307 ( .A1(n13059), .A2(n13092), .ZN(n13060) );
  AOI21_X1 U15308 ( .B1(n13121), .B2(n13061), .A(n13060), .ZN(n13366) );
  NOR2_X1 U15309 ( .A1(n13366), .A2(n13108), .ZN(n13062) );
  AOI211_X1 U15310 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(P2_U3088), .A(n13063), 
        .B(n13062), .ZN(n13064) );
  OAI211_X1 U15311 ( .C1(n13359), .C2(n13114), .A(n13065), .B(n13064), .ZN(
        P2_U3207) );
  OAI22_X1 U15312 ( .A1(n13067), .A2(n13094), .B1(n13066), .B2(n13092), .ZN(
        n13413) );
  AOI22_X1 U15313 ( .A1(n13413), .A2(n13099), .B1(P2_REG3_REG_18__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13068) );
  OAI21_X1 U15314 ( .B1(n13418), .B2(n13097), .A(n13068), .ZN(n13074) );
  AOI211_X1 U15315 ( .C1(n13072), .C2(n13071), .A(n13070), .B(n13069), .ZN(
        n13073) );
  AOI211_X1 U15316 ( .C1(n13541), .C2(n13081), .A(n13074), .B(n13073), .ZN(
        n13075) );
  INV_X1 U15317 ( .A(n13075), .ZN(P2_U3210) );
  XOR2_X1 U15318 ( .A(n13077), .B(n13076), .Z(n13078) );
  NAND2_X1 U15319 ( .A1(n13078), .A2(n9789), .ZN(n13087) );
  AND2_X1 U15320 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n13191) );
  AOI21_X1 U15321 ( .B1(n13099), .B2(n13079), .A(n13191), .ZN(n13086) );
  NAND2_X1 U15322 ( .A1(n13081), .A2(n13080), .ZN(n13085) );
  INV_X1 U15323 ( .A(n13082), .ZN(n13083) );
  NAND2_X1 U15324 ( .A1(n13110), .A2(n13083), .ZN(n13084) );
  NAND4_X1 U15325 ( .A1(n13087), .A2(n13086), .A3(n13085), .A4(n13084), .ZN(
        P2_U3211) );
  OAI21_X1 U15326 ( .B1(n13088), .B2(n13090), .A(n13089), .ZN(n13091) );
  NAND2_X1 U15327 ( .A1(n13091), .A2(n9789), .ZN(n13101) );
  OAI22_X1 U15328 ( .A1(n13095), .A2(n13094), .B1(n13093), .B2(n13092), .ZN(
        n13295) );
  OAI22_X1 U15329 ( .A1(n13301), .A2(n13097), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13096), .ZN(n13098) );
  AOI21_X1 U15330 ( .B1(n13295), .B2(n13099), .A(n13098), .ZN(n13100) );
  OAI211_X1 U15331 ( .C1(n13102), .C2(n13114), .A(n13101), .B(n13100), .ZN(
        P2_U3212) );
  OAI211_X1 U15332 ( .C1(n13105), .C2(n13104), .A(n13103), .B(n9789), .ZN(
        n13113) );
  OAI22_X1 U15333 ( .A1(n13108), .A2(n13107), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13106), .ZN(n13109) );
  AOI21_X1 U15334 ( .B1(n13111), .B2(n13110), .A(n13109), .ZN(n13112) );
  OAI211_X1 U15335 ( .C1(n13115), .C2(n13114), .A(n13113), .B(n13112), .ZN(
        P2_U3213) );
  MUX2_X1 U15336 ( .A(n13116), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13132), .Z(
        P2_U3561) );
  MUX2_X1 U15337 ( .A(n13117), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13132), .Z(
        P2_U3559) );
  MUX2_X1 U15338 ( .A(n13118), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13132), .Z(
        P2_U3558) );
  MUX2_X1 U15339 ( .A(n13119), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13132), .Z(
        P2_U3557) );
  MUX2_X1 U15340 ( .A(n13120), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13132), .Z(
        P2_U3555) );
  MUX2_X1 U15341 ( .A(n13121), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13132), .Z(
        P2_U3554) );
  MUX2_X1 U15342 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13122), .S(P2_U3947), .Z(
        P2_U3553) );
  MUX2_X1 U15343 ( .A(n13123), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13132), .Z(
        P2_U3552) );
  MUX2_X1 U15344 ( .A(n13124), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13132), .Z(
        P2_U3551) );
  MUX2_X1 U15345 ( .A(n13125), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13132), .Z(
        P2_U3550) );
  MUX2_X1 U15346 ( .A(n13126), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13132), .Z(
        P2_U3548) );
  MUX2_X1 U15347 ( .A(n13127), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13132), .Z(
        P2_U3547) );
  MUX2_X1 U15348 ( .A(n13128), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13132), .Z(
        P2_U3546) );
  MUX2_X1 U15349 ( .A(n13129), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13132), .Z(
        P2_U3545) );
  MUX2_X1 U15350 ( .A(n13130), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13132), .Z(
        P2_U3544) );
  MUX2_X1 U15351 ( .A(n13131), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13132), .Z(
        P2_U3543) );
  MUX2_X1 U15352 ( .A(n13133), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13132), .Z(
        P2_U3542) );
  MUX2_X1 U15353 ( .A(n13134), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13132), .Z(
        P2_U3541) );
  MUX2_X1 U15354 ( .A(n13135), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13132), .Z(
        P2_U3540) );
  MUX2_X1 U15355 ( .A(n13136), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13132), .Z(
        P2_U3539) );
  MUX2_X1 U15356 ( .A(n13137), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13132), .Z(
        P2_U3538) );
  MUX2_X1 U15357 ( .A(n13138), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13132), .Z(
        P2_U3537) );
  MUX2_X1 U15358 ( .A(n13139), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13132), .Z(
        P2_U3536) );
  MUX2_X1 U15359 ( .A(n13140), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13132), .Z(
        P2_U3535) );
  MUX2_X1 U15360 ( .A(n13141), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13132), .Z(
        P2_U3534) );
  MUX2_X1 U15361 ( .A(n13142), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13132), .Z(
        P2_U3533) );
  MUX2_X1 U15362 ( .A(n11872), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13132), .Z(
        P2_U3532) );
  MUX2_X1 U15363 ( .A(n13143), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13132), .Z(
        P2_U3531) );
  INV_X1 U15364 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n13145) );
  OAI22_X1 U15365 ( .A1(n14791), .A2(n13145), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13144), .ZN(n13146) );
  AOI21_X1 U15366 ( .B1(n13147), .B2(n14818), .A(n13146), .ZN(n13159) );
  MUX2_X1 U15367 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9939), .S(n13152), .Z(
        n13150) );
  NAND3_X1 U15368 ( .A1(n13150), .A2(n13149), .A3(n13148), .ZN(n13151) );
  NAND3_X1 U15369 ( .A1(n14814), .A2(n13164), .A3(n13151), .ZN(n13158) );
  MUX2_X1 U15370 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n7737), .S(n13152), .Z(
        n13155) );
  NAND3_X1 U15371 ( .A1(n13155), .A2(n13154), .A3(n13153), .ZN(n13156) );
  NAND3_X1 U15372 ( .A1(n14820), .A2(n13169), .A3(n13156), .ZN(n13157) );
  NAND3_X1 U15373 ( .A1(n13159), .A2(n13158), .A3(n13157), .ZN(P2_U3216) );
  NOR2_X1 U15374 ( .A1(n14769), .A2(n13166), .ZN(n13160) );
  AOI211_X1 U15375 ( .C1(n14812), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n13161), .B(
        n13160), .ZN(n13173) );
  MUX2_X1 U15376 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9942), .S(n13166), .Z(
        n13162) );
  NAND3_X1 U15377 ( .A1(n13164), .A2(n13163), .A3(n13162), .ZN(n13165) );
  NAND3_X1 U15378 ( .A1(n14814), .A2(n13178), .A3(n13165), .ZN(n13172) );
  MUX2_X1 U15379 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10642), .S(n13166), .Z(
        n13168) );
  NAND3_X1 U15380 ( .A1(n13169), .A2(n13168), .A3(n13167), .ZN(n13170) );
  NAND3_X1 U15381 ( .A1(n14820), .A2(n13184), .A3(n13170), .ZN(n13171) );
  NAND3_X1 U15382 ( .A1(n13173), .A2(n13172), .A3(n13171), .ZN(P2_U3217) );
  NOR2_X1 U15383 ( .A1(n14769), .A2(n13181), .ZN(n13174) );
  AOI211_X1 U15384 ( .C1(n14812), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n13175), .B(
        n13174), .ZN(n13189) );
  MUX2_X1 U15385 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9945), .S(n13181), .Z(
        n13176) );
  NAND3_X1 U15386 ( .A1(n13178), .A2(n13177), .A3(n13176), .ZN(n13179) );
  NAND3_X1 U15387 ( .A1(n14814), .A2(n13180), .A3(n13179), .ZN(n13188) );
  MUX2_X1 U15388 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10774), .S(n13181), .Z(
        n13182) );
  NAND3_X1 U15389 ( .A1(n13184), .A2(n13183), .A3(n13182), .ZN(n13185) );
  NAND3_X1 U15390 ( .A1(n14820), .A2(n13186), .A3(n13185), .ZN(n13187) );
  NAND3_X1 U15391 ( .A1(n13189), .A2(n13188), .A3(n13187), .ZN(P2_U3218) );
  NOR2_X1 U15392 ( .A1(n14769), .A2(n13196), .ZN(n13190) );
  AOI211_X1 U15393 ( .C1(n14812), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n13191), .B(
        n13190), .ZN(n13203) );
  MUX2_X1 U15394 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10067), .S(n13196), .Z(
        n13192) );
  NAND3_X1 U15395 ( .A1(n13194), .A2(n13193), .A3(n13192), .ZN(n13195) );
  NAND3_X1 U15396 ( .A1(n14814), .A2(n13208), .A3(n13195), .ZN(n13202) );
  MUX2_X1 U15397 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11035), .S(n13196), .Z(
        n13197) );
  NAND3_X1 U15398 ( .A1(n13199), .A2(n13198), .A3(n13197), .ZN(n13200) );
  NAND3_X1 U15399 ( .A1(n14820), .A2(n13213), .A3(n13200), .ZN(n13201) );
  NAND3_X1 U15400 ( .A1(n13203), .A2(n13202), .A3(n13201), .ZN(P2_U3220) );
  NOR2_X1 U15401 ( .A1(n14769), .A2(n13210), .ZN(n13204) );
  AOI211_X1 U15402 ( .C1(n14812), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n13205), .B(
        n13204), .ZN(n13217) );
  MUX2_X1 U15403 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10070), .S(n13210), .Z(
        n13206) );
  NAND3_X1 U15404 ( .A1(n13208), .A2(n13207), .A3(n13206), .ZN(n13209) );
  NAND3_X1 U15405 ( .A1(n14814), .A2(n13224), .A3(n13209), .ZN(n13216) );
  MUX2_X1 U15406 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10084), .S(n13210), .Z(
        n13211) );
  NAND3_X1 U15407 ( .A1(n13213), .A2(n13212), .A3(n13211), .ZN(n13214) );
  NAND3_X1 U15408 ( .A1(n14820), .A2(n13230), .A3(n13214), .ZN(n13215) );
  NAND3_X1 U15409 ( .A1(n13217), .A2(n13216), .A3(n13215), .ZN(P2_U3221) );
  INV_X1 U15410 ( .A(n13218), .ZN(n13220) );
  NOR2_X1 U15411 ( .A1(n14769), .A2(n13227), .ZN(n13219) );
  AOI211_X1 U15412 ( .C1(n14812), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n13220), .B(
        n13219), .ZN(n13235) );
  MUX2_X1 U15413 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n13221), .S(n13227), .Z(
        n13222) );
  NAND3_X1 U15414 ( .A1(n13224), .A2(n13223), .A3(n13222), .ZN(n13225) );
  NAND3_X1 U15415 ( .A1(n14814), .A2(n13226), .A3(n13225), .ZN(n13234) );
  MUX2_X1 U15416 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10991), .S(n13227), .Z(
        n13228) );
  NAND3_X1 U15417 ( .A1(n13230), .A2(n13229), .A3(n13228), .ZN(n13231) );
  NAND3_X1 U15418 ( .A1(n14820), .A2(n13232), .A3(n13231), .ZN(n13233) );
  NAND3_X1 U15419 ( .A1(n13235), .A2(n13234), .A3(n13233), .ZN(P2_U3222) );
  NOR2_X1 U15420 ( .A1(n13241), .A2(n13236), .ZN(n13237) );
  NOR2_X1 U15421 ( .A1(n13238), .A2(n13237), .ZN(n13239) );
  XOR2_X1 U15422 ( .A(n13239), .B(P2_REG2_REG_19__SCAN_IN), .Z(n13248) );
  INV_X1 U15423 ( .A(n13248), .ZN(n13246) );
  NAND2_X1 U15424 ( .A1(n13241), .A2(n13240), .ZN(n13242) );
  NAND2_X1 U15425 ( .A1(n13243), .A2(n13242), .ZN(n13244) );
  XOR2_X1 U15426 ( .A(n13244), .B(P2_REG1_REG_19__SCAN_IN), .Z(n13247) );
  NOR2_X1 U15427 ( .A1(n13247), .A2(n14750), .ZN(n13245) );
  AOI211_X1 U15428 ( .C1(n13246), .C2(n14820), .A(n14818), .B(n13245), .ZN(
        n13251) );
  AOI22_X1 U15429 ( .A1(n13248), .A2(n14820), .B1(n14814), .B2(n13247), .ZN(
        n13250) );
  MUX2_X1 U15430 ( .A(n13251), .B(n13250), .S(n13249), .Z(n13253) );
  OAI211_X1 U15431 ( .C1(n13254), .C2(n14791), .A(n13253), .B(n13252), .ZN(
        P2_U3233) );
  NAND2_X1 U15432 ( .A1(n13564), .A2(n13255), .ZN(n13256) );
  NAND3_X1 U15433 ( .A1(n13257), .A2(n13372), .A3(n13256), .ZN(n13485) );
  AOI21_X1 U15434 ( .B1(n13428), .B2(P2_REG2_REG_30__SCAN_IN), .A(n13258), 
        .ZN(n13260) );
  NAND2_X1 U15435 ( .A1(n13564), .A2(n13476), .ZN(n13259) );
  OAI211_X1 U15436 ( .C1(n13485), .C2(n13350), .A(n13260), .B(n13259), .ZN(
        P2_U3235) );
  XNOR2_X1 U15437 ( .A(n13262), .B(n13261), .ZN(n13272) );
  INV_X1 U15438 ( .A(n13272), .ZN(n13492) );
  INV_X1 U15439 ( .A(n13263), .ZN(n13273) );
  NAND2_X1 U15440 ( .A1(n13264), .A2(n13430), .ZN(n13270) );
  AOI211_X1 U15441 ( .C1(n13489), .C2(n13285), .A(n13460), .B(n6554), .ZN(
        n13488) );
  INV_X1 U15442 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13275) );
  OAI22_X1 U15443 ( .A1(n13276), .A2(n13463), .B1(n13275), .B2(n13468), .ZN(
        n13277) );
  AOI21_X1 U15444 ( .B1(n13488), .B2(n13478), .A(n13277), .ZN(n13278) );
  XNOR2_X1 U15445 ( .A(n13281), .B(n13280), .ZN(n13572) );
  INV_X1 U15446 ( .A(n13494), .ZN(n13292) );
  OAI211_X1 U15447 ( .C1(n13286), .C2(n13305), .A(n13372), .B(n13285), .ZN(
        n13493) );
  INV_X1 U15448 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13287) );
  OAI22_X1 U15449 ( .A1(n13288), .A2(n13472), .B1(n13287), .B2(n13468), .ZN(
        n13289) );
  AOI21_X1 U15450 ( .B1(n13569), .B2(n13476), .A(n13289), .ZN(n13290) );
  OAI21_X1 U15451 ( .B1(n13493), .B2(n13350), .A(n13290), .ZN(n13291) );
  AOI21_X1 U15452 ( .B1(n13292), .B2(n13468), .A(n13291), .ZN(n13293) );
  OAI21_X1 U15453 ( .B1(n13467), .B2(n13572), .A(n13293), .ZN(P2_U3238) );
  XNOR2_X1 U15454 ( .A(n13294), .B(n13299), .ZN(n13297) );
  INV_X1 U15455 ( .A(n13295), .ZN(n13296) );
  OAI21_X1 U15456 ( .B1(n13297), .B2(n13454), .A(n13296), .ZN(n13498) );
  XNOR2_X1 U15457 ( .A(n13299), .B(n13298), .ZN(n13576) );
  INV_X1 U15458 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n13300) );
  OAI22_X1 U15459 ( .A1(n13301), .A2(n13472), .B1(n13300), .B2(n13468), .ZN(
        n13302) );
  AOI21_X1 U15460 ( .B1(n13500), .B2(n13476), .A(n13302), .ZN(n13307) );
  NAND2_X1 U15461 ( .A1(n13500), .A2(n13315), .ZN(n13303) );
  NAND2_X1 U15462 ( .A1(n13303), .A2(n13372), .ZN(n13304) );
  NOR2_X1 U15463 ( .A1(n13305), .A2(n13304), .ZN(n13499) );
  NAND2_X1 U15464 ( .A1(n13499), .A2(n13478), .ZN(n13306) );
  OAI211_X1 U15465 ( .C1(n13576), .C2(n13467), .A(n13307), .B(n13306), .ZN(
        n13308) );
  AOI21_X1 U15466 ( .B1(n13498), .B2(n13468), .A(n13308), .ZN(n13309) );
  INV_X1 U15467 ( .A(n13309), .ZN(P2_U3239) );
  XOR2_X1 U15468 ( .A(n13310), .B(n13312), .Z(n13580) );
  XOR2_X1 U15469 ( .A(n13311), .B(n13312), .Z(n13314) );
  OAI21_X1 U15470 ( .B1(n13314), .B2(n13454), .A(n13313), .ZN(n13503) );
  NAND2_X1 U15471 ( .A1(n13503), .A2(n13468), .ZN(n13323) );
  INV_X1 U15472 ( .A(n13315), .ZN(n13316) );
  AOI211_X1 U15473 ( .C1(n13505), .C2(n13317), .A(n13460), .B(n13316), .ZN(
        n13504) );
  AOI22_X1 U15474 ( .A1(n13318), .A2(n13419), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n13428), .ZN(n13319) );
  OAI21_X1 U15475 ( .B1(n13320), .B2(n13463), .A(n13319), .ZN(n13321) );
  AOI21_X1 U15476 ( .B1(n13504), .B2(n13478), .A(n13321), .ZN(n13322) );
  OAI211_X1 U15477 ( .C1(n13467), .C2(n13580), .A(n13323), .B(n13322), .ZN(
        P2_U3240) );
  XNOR2_X1 U15478 ( .A(n13324), .B(n13329), .ZN(n13327) );
  INV_X1 U15479 ( .A(n13325), .ZN(n13326) );
  OAI21_X1 U15480 ( .B1(n13327), .B2(n13454), .A(n13326), .ZN(n13507) );
  INV_X1 U15481 ( .A(n13507), .ZN(n13338) );
  XNOR2_X1 U15482 ( .A(n13328), .B(n13329), .ZN(n13509) );
  AOI211_X1 U15483 ( .C1(n13331), .C2(n13347), .A(n13460), .B(n13330), .ZN(
        n13508) );
  NAND2_X1 U15484 ( .A1(n13508), .A2(n13478), .ZN(n13335) );
  INV_X1 U15485 ( .A(n13332), .ZN(n13333) );
  AOI22_X1 U15486 ( .A1(n13333), .A2(n13419), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n13428), .ZN(n13334) );
  OAI211_X1 U15487 ( .C1(n13584), .C2(n13463), .A(n13335), .B(n13334), .ZN(
        n13336) );
  AOI21_X1 U15488 ( .B1(n13470), .B2(n13509), .A(n13336), .ZN(n13337) );
  OAI21_X1 U15489 ( .B1(n13428), .B2(n13338), .A(n13337), .ZN(P2_U3241) );
  INV_X1 U15490 ( .A(n13515), .ZN(n13343) );
  INV_X1 U15491 ( .A(n13339), .ZN(n13346) );
  XNOR2_X1 U15492 ( .A(n13340), .B(n13346), .ZN(n13341) );
  NAND2_X1 U15493 ( .A1(n13341), .A2(n13430), .ZN(n13514) );
  INV_X1 U15494 ( .A(n13514), .ZN(n13342) );
  AOI211_X1 U15495 ( .C1(n13419), .C2(n13344), .A(n13343), .B(n13342), .ZN(
        n13353) );
  XNOR2_X1 U15496 ( .A(n13345), .B(n13346), .ZN(n13512) );
  OAI211_X1 U15497 ( .C1(n13348), .C2(n13358), .A(n13372), .B(n13347), .ZN(
        n13513) );
  AOI22_X1 U15498 ( .A1(n13587), .A2(n13476), .B1(n13428), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n13349) );
  OAI21_X1 U15499 ( .B1(n13513), .B2(n13350), .A(n13349), .ZN(n13351) );
  AOI21_X1 U15500 ( .B1(n13512), .B2(n13470), .A(n13351), .ZN(n13352) );
  OAI21_X1 U15501 ( .B1(n13353), .B2(n13428), .A(n13352), .ZN(P2_U3242) );
  INV_X1 U15502 ( .A(n13354), .ZN(n13357) );
  OAI21_X1 U15503 ( .B1(n13357), .B2(n13356), .A(n13355), .ZN(n13594) );
  AOI211_X1 U15504 ( .C1(n13591), .C2(n13371), .A(n13460), .B(n13358), .ZN(
        n13519) );
  NOR2_X1 U15505 ( .A1(n13359), .A2(n13463), .ZN(n13363) );
  OAI22_X1 U15506 ( .A1(n13361), .A2(n13472), .B1(n13360), .B2(n13468), .ZN(
        n13362) );
  AOI211_X1 U15507 ( .C1(n13519), .C2(n13478), .A(n13363), .B(n13362), .ZN(
        n13369) );
  XNOR2_X1 U15508 ( .A(n13364), .B(n13365), .ZN(n13367) );
  OAI21_X1 U15509 ( .B1(n13367), .B2(n13454), .A(n13366), .ZN(n13520) );
  NAND2_X1 U15510 ( .A1(n13520), .A2(n13468), .ZN(n13368) );
  OAI211_X1 U15511 ( .C1(n13467), .C2(n13594), .A(n13369), .B(n13368), .ZN(
        P2_U3243) );
  XOR2_X1 U15512 ( .A(n13378), .B(n13370), .Z(n13598) );
  OAI211_X1 U15513 ( .C1(n13376), .C2(n13385), .A(n13372), .B(n13371), .ZN(
        n13373) );
  INV_X1 U15514 ( .A(n13373), .ZN(n13525) );
  AOI22_X1 U15515 ( .A1(n13374), .A2(n13419), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n13428), .ZN(n13375) );
  OAI21_X1 U15516 ( .B1(n13376), .B2(n13463), .A(n13375), .ZN(n13377) );
  AOI21_X1 U15517 ( .B1(n13525), .B2(n13478), .A(n13377), .ZN(n13383) );
  XOR2_X1 U15518 ( .A(n13379), .B(n13378), .Z(n13381) );
  OAI21_X1 U15519 ( .B1(n13381), .B2(n13454), .A(n13380), .ZN(n13524) );
  NAND2_X1 U15520 ( .A1(n13524), .A2(n13468), .ZN(n13382) );
  OAI211_X1 U15521 ( .C1(n13598), .C2(n13467), .A(n13383), .B(n13382), .ZN(
        P2_U3244) );
  XOR2_X1 U15522 ( .A(n13384), .B(n13392), .Z(n13531) );
  INV_X1 U15523 ( .A(n13531), .ZN(n13398) );
  INV_X1 U15524 ( .A(n13404), .ZN(n13386) );
  AOI211_X1 U15525 ( .C1(n13387), .C2(n13386), .A(n13460), .B(n13385), .ZN(
        n13530) );
  NOR2_X1 U15526 ( .A1(n13603), .A2(n13463), .ZN(n13391) );
  OAI22_X1 U15527 ( .A1(n13389), .A2(n13472), .B1(n13388), .B2(n13468), .ZN(
        n13390) );
  AOI211_X1 U15528 ( .C1(n13530), .C2(n13478), .A(n13391), .B(n13390), .ZN(
        n13397) );
  XOR2_X1 U15529 ( .A(n13393), .B(n13392), .Z(n13395) );
  OAI21_X1 U15530 ( .B1(n13395), .B2(n13454), .A(n13394), .ZN(n13529) );
  NAND2_X1 U15531 ( .A1(n13529), .A2(n13468), .ZN(n13396) );
  OAI211_X1 U15532 ( .C1(n13398), .C2(n13467), .A(n13397), .B(n13396), .ZN(
        P2_U3245) );
  XNOR2_X1 U15533 ( .A(n13399), .B(n13401), .ZN(n13539) );
  XOR2_X1 U15534 ( .A(n13400), .B(n13401), .Z(n13403) );
  OAI21_X1 U15535 ( .B1(n13403), .B2(n13454), .A(n13402), .ZN(n13535) );
  NAND2_X1 U15536 ( .A1(n13535), .A2(n13468), .ZN(n13410) );
  AOI211_X1 U15537 ( .C1(n13537), .C2(n13415), .A(n13460), .B(n13404), .ZN(
        n13536) );
  INV_X1 U15538 ( .A(n13537), .ZN(n13407) );
  AOI22_X1 U15539 ( .A1(P2_REG2_REG_19__SCAN_IN), .A2(n13428), .B1(n13405), 
        .B2(n13419), .ZN(n13406) );
  OAI21_X1 U15540 ( .B1(n13407), .B2(n13463), .A(n13406), .ZN(n13408) );
  AOI21_X1 U15541 ( .B1(n13536), .B2(n13478), .A(n13408), .ZN(n13409) );
  OAI211_X1 U15542 ( .C1(n13467), .C2(n13539), .A(n13410), .B(n13409), .ZN(
        P2_U3246) );
  XNOR2_X1 U15543 ( .A(n13412), .B(n13411), .ZN(n13414) );
  AOI21_X1 U15544 ( .B1(n13414), .B2(n13430), .A(n13413), .ZN(n13543) );
  INV_X1 U15545 ( .A(n13443), .ZN(n13417) );
  INV_X1 U15546 ( .A(n13415), .ZN(n13416) );
  AOI211_X1 U15547 ( .C1(n13541), .C2(n13417), .A(n13460), .B(n13416), .ZN(
        n13540) );
  INV_X1 U15548 ( .A(n13418), .ZN(n13420) );
  AOI22_X1 U15549 ( .A1(n13428), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13420), 
        .B2(n13419), .ZN(n13421) );
  OAI21_X1 U15550 ( .B1(n13422), .B2(n13463), .A(n13421), .ZN(n13426) );
  AOI21_X1 U15551 ( .B1(n13424), .B2(n13423), .A(n6590), .ZN(n13544) );
  NOR2_X1 U15552 ( .A1(n13544), .A2(n13467), .ZN(n13425) );
  AOI211_X1 U15553 ( .C1(n13540), .C2(n13478), .A(n13426), .B(n13425), .ZN(
        n13427) );
  OAI21_X1 U15554 ( .B1(n13428), .B2(n13543), .A(n13427), .ZN(P2_U3247) );
  OAI211_X1 U15555 ( .C1(n13432), .C2(n13431), .A(n13430), .B(n13429), .ZN(
        n13434) );
  NAND2_X1 U15556 ( .A1(n13434), .A2(n13433), .ZN(n13545) );
  OAI21_X1 U15557 ( .B1(n13437), .B2(n13436), .A(n13435), .ZN(n13609) );
  OAI22_X1 U15558 ( .A1(n13468), .A2(n13439), .B1(n13438), .B2(n13472), .ZN(
        n13440) );
  AOI21_X1 U15559 ( .B1(n11978), .B2(n13476), .A(n13440), .ZN(n13445) );
  NAND2_X1 U15560 ( .A1(n11978), .A2(n13458), .ZN(n13441) );
  NAND2_X1 U15561 ( .A1(n13441), .A2(n13372), .ZN(n13442) );
  NOR2_X1 U15562 ( .A1(n13443), .A2(n13442), .ZN(n13546) );
  NAND2_X1 U15563 ( .A1(n13546), .A2(n13478), .ZN(n13444) );
  OAI211_X1 U15564 ( .C1(n13609), .C2(n13467), .A(n13445), .B(n13444), .ZN(
        n13446) );
  AOI21_X1 U15565 ( .B1(n13468), .B2(n13545), .A(n13446), .ZN(n13447) );
  INV_X1 U15566 ( .A(n13447), .ZN(P2_U3248) );
  NAND2_X1 U15567 ( .A1(n13448), .A2(n13452), .ZN(n13449) );
  NAND2_X1 U15568 ( .A1(n13450), .A2(n13449), .ZN(n13613) );
  XOR2_X1 U15569 ( .A(n13452), .B(n13451), .Z(n13455) );
  OAI21_X1 U15570 ( .B1(n13455), .B2(n13454), .A(n13453), .ZN(n13549) );
  NOR2_X1 U15571 ( .A1(n13472), .A2(n13456), .ZN(n13457) );
  OAI21_X1 U15572 ( .B1(n13549), .B2(n13457), .A(n13468), .ZN(n13466) );
  INV_X1 U15573 ( .A(n13458), .ZN(n13459) );
  AOI211_X1 U15574 ( .C1(n13551), .C2(n13461), .A(n13460), .B(n13459), .ZN(
        n13550) );
  OAI22_X1 U15575 ( .A1(n7107), .A2(n13463), .B1(n13462), .B2(n13468), .ZN(
        n13464) );
  AOI21_X1 U15576 ( .B1(n13550), .B2(n13478), .A(n13464), .ZN(n13465) );
  OAI211_X1 U15577 ( .C1(n13467), .C2(n13613), .A(n13466), .B(n13465), .ZN(
        P2_U3249) );
  NAND2_X1 U15578 ( .A1(n13469), .A2(n13468), .ZN(n13483) );
  NAND2_X1 U15579 ( .A1(n13471), .A2(n13470), .ZN(n13482) );
  OAI22_X1 U15580 ( .A1(n13468), .A2(n13474), .B1(n13473), .B2(n13472), .ZN(
        n13475) );
  AOI21_X1 U15581 ( .B1(n13477), .B2(n13476), .A(n13475), .ZN(n13481) );
  NAND2_X1 U15582 ( .A1(n13479), .A2(n13478), .ZN(n13480) );
  NAND4_X1 U15583 ( .A1(n13483), .A2(n13482), .A3(n13481), .A4(n13480), .ZN(
        P2_U3256) );
  NAND2_X1 U15584 ( .A1(n13485), .A2(n13484), .ZN(n13562) );
  MUX2_X1 U15585 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13562), .S(n14864), .Z(
        n13486) );
  AOI21_X1 U15586 ( .B1(n13558), .B2(n13564), .A(n13486), .ZN(n13487) );
  INV_X1 U15587 ( .A(n13487), .ZN(P2_U3529) );
  AOI21_X1 U15588 ( .B1(n14845), .B2(n13489), .A(n13488), .ZN(n13490) );
  MUX2_X1 U15589 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13566), .S(n14864), .Z(
        P2_U3527) );
  MUX2_X1 U15590 ( .A(n13495), .B(n13567), .S(n14864), .Z(n13497) );
  NAND2_X1 U15591 ( .A1(n13569), .A2(n13558), .ZN(n13496) );
  AOI211_X1 U15592 ( .C1(n14845), .C2(n13500), .A(n13499), .B(n13498), .ZN(
        n13573) );
  MUX2_X1 U15593 ( .A(n13501), .B(n13573), .S(n14864), .Z(n13502) );
  OAI21_X1 U15594 ( .B1(n13576), .B2(n13561), .A(n13502), .ZN(P2_U3525) );
  AOI211_X1 U15595 ( .C1(n14845), .C2(n13505), .A(n13504), .B(n13503), .ZN(
        n13577) );
  MUX2_X1 U15596 ( .A(n15194), .B(n13577), .S(n13552), .Z(n13506) );
  OAI21_X1 U15597 ( .B1(n13580), .B2(n13561), .A(n13506), .ZN(P2_U3524) );
  AOI211_X1 U15598 ( .C1(n14850), .C2(n13509), .A(n13508), .B(n13507), .ZN(
        n13581) );
  MUX2_X1 U15599 ( .A(n13510), .B(n13581), .S(n13552), .Z(n13511) );
  OAI21_X1 U15600 ( .B1(n13584), .B2(n13534), .A(n13511), .ZN(P2_U3523) );
  NAND2_X1 U15601 ( .A1(n13512), .A2(n14850), .ZN(n13516) );
  NAND4_X1 U15602 ( .A1(n13516), .A2(n13515), .A3(n13514), .A4(n13513), .ZN(
        n13585) );
  MUX2_X1 U15603 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13585), .S(n13552), .Z(
        n13517) );
  AOI21_X1 U15604 ( .B1(n13558), .B2(n13587), .A(n13517), .ZN(n13518) );
  INV_X1 U15605 ( .A(n13518), .ZN(P2_U3522) );
  INV_X1 U15606 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n13521) );
  NOR2_X1 U15607 ( .A1(n13520), .A2(n13519), .ZN(n13589) );
  MUX2_X1 U15608 ( .A(n13521), .B(n13589), .S(n14864), .Z(n13523) );
  NAND2_X1 U15609 ( .A1(n13591), .A2(n13558), .ZN(n13522) );
  OAI211_X1 U15610 ( .C1(n13561), .C2(n13594), .A(n13523), .B(n13522), .ZN(
        P2_U3521) );
  AOI211_X1 U15611 ( .C1(n14845), .C2(n13526), .A(n13525), .B(n13524), .ZN(
        n13595) );
  MUX2_X1 U15612 ( .A(n13527), .B(n13595), .S(n13552), .Z(n13528) );
  OAI21_X1 U15613 ( .B1(n13598), .B2(n13561), .A(n13528), .ZN(P2_U3520) );
  INV_X1 U15614 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n13532) );
  AOI211_X1 U15615 ( .C1(n13531), .C2(n14850), .A(n13530), .B(n13529), .ZN(
        n13599) );
  MUX2_X1 U15616 ( .A(n13532), .B(n13599), .S(n13552), .Z(n13533) );
  OAI21_X1 U15617 ( .B1(n13603), .B2(n13534), .A(n13533), .ZN(P2_U3519) );
  AOI211_X1 U15618 ( .C1(n14845), .C2(n13537), .A(n13536), .B(n13535), .ZN(
        n13538) );
  OAI21_X1 U15619 ( .B1(n14841), .B2(n13539), .A(n13538), .ZN(n13604) );
  MUX2_X1 U15620 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13604), .S(n14864), .Z(
        P2_U3518) );
  AOI21_X1 U15621 ( .B1(n14845), .B2(n13541), .A(n13540), .ZN(n13542) );
  OAI211_X1 U15622 ( .C1(n13544), .C2(n14841), .A(n13543), .B(n13542), .ZN(
        n13605) );
  MUX2_X1 U15623 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13605), .S(n13552), .Z(
        P2_U3517) );
  AOI211_X1 U15624 ( .C1(n14845), .C2(n11978), .A(n13546), .B(n13545), .ZN(
        n13606) );
  MUX2_X1 U15625 ( .A(n13547), .B(n13606), .S(n14864), .Z(n13548) );
  OAI21_X1 U15626 ( .B1(n13561), .B2(n13609), .A(n13548), .ZN(P2_U3516) );
  AOI211_X1 U15627 ( .C1(n14845), .C2(n13551), .A(n13550), .B(n13549), .ZN(
        n13610) );
  MUX2_X1 U15628 ( .A(n13553), .B(n13610), .S(n13552), .Z(n13554) );
  OAI21_X1 U15629 ( .B1(n13561), .B2(n13613), .A(n13554), .ZN(P2_U3515) );
  NOR2_X1 U15630 ( .A1(n13556), .A2(n13555), .ZN(n13614) );
  MUX2_X1 U15631 ( .A(n13557), .B(n13614), .S(n14864), .Z(n13560) );
  NAND2_X1 U15632 ( .A1(n13617), .A2(n13558), .ZN(n13559) );
  OAI211_X1 U15633 ( .C1(n13621), .C2(n13561), .A(n13560), .B(n13559), .ZN(
        P2_U3514) );
  MUX2_X1 U15634 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13562), .S(n14859), .Z(
        n13563) );
  AOI21_X1 U15635 ( .B1(n13616), .B2(n13564), .A(n13563), .ZN(n13565) );
  INV_X1 U15636 ( .A(n13565), .ZN(P2_U3497) );
  MUX2_X1 U15637 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13566), .S(n14859), .Z(
        P2_U3495) );
  INV_X1 U15638 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n13568) );
  NAND2_X1 U15639 ( .A1(n13569), .A2(n13616), .ZN(n13570) );
  INV_X1 U15640 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n13574) );
  MUX2_X1 U15641 ( .A(n13574), .B(n13573), .S(n14859), .Z(n13575) );
  OAI21_X1 U15642 ( .B1(n13576), .B2(n13620), .A(n13575), .ZN(P2_U3493) );
  INV_X1 U15643 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n13578) );
  MUX2_X1 U15644 ( .A(n13578), .B(n13577), .S(n14859), .Z(n13579) );
  OAI21_X1 U15645 ( .B1(n13580), .B2(n13620), .A(n13579), .ZN(P2_U3492) );
  INV_X1 U15646 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n13582) );
  MUX2_X1 U15647 ( .A(n13582), .B(n13581), .S(n14859), .Z(n13583) );
  OAI21_X1 U15648 ( .B1(n13584), .B2(n13602), .A(n13583), .ZN(P2_U3491) );
  MUX2_X1 U15649 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13585), .S(n14859), .Z(
        n13586) );
  AOI21_X1 U15650 ( .B1(n13616), .B2(n13587), .A(n13586), .ZN(n13588) );
  INV_X1 U15651 ( .A(n13588), .ZN(P2_U3490) );
  INV_X1 U15652 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n13590) );
  MUX2_X1 U15653 ( .A(n13590), .B(n13589), .S(n14859), .Z(n13593) );
  NAND2_X1 U15654 ( .A1(n13591), .A2(n13616), .ZN(n13592) );
  OAI211_X1 U15655 ( .C1(n13594), .C2(n13620), .A(n13593), .B(n13592), .ZN(
        P2_U3489) );
  INV_X1 U15656 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n13596) );
  MUX2_X1 U15657 ( .A(n13596), .B(n13595), .S(n14859), .Z(n13597) );
  OAI21_X1 U15658 ( .B1(n13598), .B2(n13620), .A(n13597), .ZN(P2_U3488) );
  INV_X1 U15659 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n13600) );
  MUX2_X1 U15660 ( .A(n13600), .B(n13599), .S(n14859), .Z(n13601) );
  OAI21_X1 U15661 ( .B1(n13603), .B2(n13602), .A(n13601), .ZN(P2_U3487) );
  MUX2_X1 U15662 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13604), .S(n14859), .Z(
        P2_U3486) );
  MUX2_X1 U15663 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13605), .S(n14859), .Z(
        P2_U3484) );
  INV_X1 U15664 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n13607) );
  MUX2_X1 U15665 ( .A(n13607), .B(n13606), .S(n14859), .Z(n13608) );
  OAI21_X1 U15666 ( .B1(n13609), .B2(n13620), .A(n13608), .ZN(P2_U3481) );
  INV_X1 U15667 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n13611) );
  MUX2_X1 U15668 ( .A(n13611), .B(n13610), .S(n14859), .Z(n13612) );
  OAI21_X1 U15669 ( .B1(n13613), .B2(n13620), .A(n13612), .ZN(P2_U3478) );
  MUX2_X1 U15670 ( .A(n13615), .B(n13614), .S(n14859), .Z(n13619) );
  NAND2_X1 U15671 ( .A1(n13617), .A2(n13616), .ZN(n13618) );
  OAI211_X1 U15672 ( .C1(n13621), .C2(n13620), .A(n13619), .B(n13618), .ZN(
        P2_U3475) );
  INV_X1 U15673 ( .A(n13622), .ZN(n14190) );
  NAND3_X1 U15674 ( .A1(n13623), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n13626) );
  OAI22_X1 U15675 ( .A1(n7191), .A2(n13626), .B1(n13625), .B2(n13624), .ZN(
        n13627) );
  INV_X1 U15676 ( .A(n13627), .ZN(n13628) );
  OAI21_X1 U15677 ( .B1(n14190), .B2(n13645), .A(n13628), .ZN(P2_U3296) );
  OAI222_X1 U15678 ( .A1(n13645), .A2(n13631), .B1(n13629), .B2(P2_U3088), 
        .C1(n13630), .C2(n13650), .ZN(P2_U3297) );
  INV_X1 U15679 ( .A(n13632), .ZN(n14191) );
  OAI222_X1 U15680 ( .A1(n13645), .A2(n14191), .B1(n13634), .B2(P2_U3088), 
        .C1(n13633), .C2(n13650), .ZN(P2_U3298) );
  NAND2_X1 U15681 ( .A1(n14193), .A2(n13635), .ZN(n13637) );
  OAI211_X1 U15682 ( .C1(n13650), .C2(n13638), .A(n13637), .B(n13636), .ZN(
        P2_U3299) );
  INV_X1 U15683 ( .A(n13639), .ZN(n14196) );
  OAI222_X1 U15684 ( .A1(n13650), .A2(n13641), .B1(n13651), .B2(n14196), .C1(
        P2_U3088), .C2(n13640), .ZN(P2_U3300) );
  INV_X1 U15685 ( .A(n13642), .ZN(n14198) );
  OAI222_X1 U15686 ( .A1(n13645), .A2(n14198), .B1(P2_U3088), .B2(n13644), 
        .C1(n13643), .C2(n13650), .ZN(P2_U3301) );
  OAI222_X1 U15687 ( .A1(n13650), .A2(n13648), .B1(n13651), .B2(n13647), .C1(
        n13646), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U15688 ( .A(n13649), .ZN(n14203) );
  OAI222_X1 U15689 ( .A1(P2_U3088), .A2(n13652), .B1(n13651), .B2(n14203), 
        .C1(n13650), .C2(n8952), .ZN(P2_U3303) );
  INV_X1 U15690 ( .A(n13653), .ZN(n13654) );
  MUX2_X1 U15691 ( .A(n13654), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI21_X1 U15692 ( .B1(n13657), .B2(n13656), .A(n13655), .ZN(n13658) );
  AOI22_X1 U15693 ( .A1(n14510), .A2(n13944), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13659) );
  OAI21_X1 U15694 ( .B1(n13660), .B2(n13791), .A(n13659), .ZN(n13661) );
  AOI21_X1 U15695 ( .B1(n13662), .B2(n13794), .A(n13661), .ZN(n13663) );
  INV_X1 U15696 ( .A(n13665), .ZN(n13760) );
  INV_X1 U15697 ( .A(n13666), .ZN(n13668) );
  NOR3_X1 U15698 ( .A1(n13760), .A2(n13668), .A3(n13667), .ZN(n13670) );
  INV_X1 U15699 ( .A(n13669), .ZN(n13730) );
  OAI21_X1 U15700 ( .B1(n13670), .B2(n13730), .A(n14580), .ZN(n13675) );
  NAND2_X1 U15701 ( .A1(n14004), .A2(n14339), .ZN(n13672) );
  NAND2_X1 U15702 ( .A1(n13943), .A2(n14050), .ZN(n13671) );
  AND2_X1 U15703 ( .A1(n13672), .A2(n13671), .ZN(n14110) );
  OAI22_X1 U15704 ( .A1(n14496), .A2(n14110), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15301), .ZN(n13673) );
  AOI21_X1 U15705 ( .B1(n13980), .B2(n13794), .A(n13673), .ZN(n13674) );
  OAI211_X1 U15706 ( .C1(n14112), .C2(n14577), .A(n13675), .B(n13674), .ZN(
        P1_U3216) );
  INV_X1 U15707 ( .A(n13676), .ZN(n13767) );
  OAI21_X1 U15708 ( .B1(n13767), .B2(n13678), .A(n13677), .ZN(n13680) );
  NAND3_X1 U15709 ( .A1(n13680), .A2(n14580), .A3(n13679), .ZN(n13685) );
  NOR2_X1 U15710 ( .A1(n14572), .A2(n14040), .ZN(n13683) );
  INV_X1 U15711 ( .A(n14510), .ZN(n13723) );
  NAND2_X1 U15712 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13891)
         );
  OAI21_X1 U15713 ( .B1(n13723), .B2(n13681), .A(n13891), .ZN(n13682) );
  AOI211_X1 U15714 ( .C1(n14512), .C2(n14039), .A(n13683), .B(n13682), .ZN(
        n13684) );
  OAI211_X1 U15715 ( .C1(n14136), .C2(n14577), .A(n13685), .B(n13684), .ZN(
        P1_U3219) );
  AOI21_X1 U15716 ( .B1(n13687), .B2(n13686), .A(n6468), .ZN(n13692) );
  AND2_X1 U15717 ( .A1(n14012), .A2(n14740), .ZN(n14124) );
  NOR2_X1 U15718 ( .A1(n14572), .A2(n14009), .ZN(n13690) );
  AOI22_X1 U15719 ( .A1(n14510), .A2(n14039), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13688) );
  OAI21_X1 U15720 ( .B1(n6899), .B2(n13791), .A(n13688), .ZN(n13689) );
  AOI211_X1 U15721 ( .C1(n14124), .C2(n14564), .A(n13690), .B(n13689), .ZN(
        n13691) );
  OAI21_X1 U15722 ( .B1(n13692), .B2(n14565), .A(n13691), .ZN(P1_U3223) );
  INV_X1 U15723 ( .A(n13693), .ZN(n13731) );
  INV_X1 U15724 ( .A(n13694), .ZN(n13696) );
  NOR3_X1 U15725 ( .A1(n13731), .A2(n13696), .A3(n13695), .ZN(n13699) );
  INV_X1 U15726 ( .A(n13697), .ZN(n13698) );
  OAI21_X1 U15727 ( .B1(n13699), .B2(n13698), .A(n14580), .ZN(n13704) );
  AOI22_X1 U15728 ( .A1(n14510), .A2(n13943), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13700) );
  OAI21_X1 U15729 ( .B1(n13701), .B2(n13791), .A(n13700), .ZN(n13702) );
  AOI21_X1 U15730 ( .B1(n13945), .B2(n13794), .A(n13702), .ZN(n13703) );
  OAI211_X1 U15731 ( .C1(n14100), .C2(n14577), .A(n13704), .B(n13703), .ZN(
        P1_U3225) );
  INV_X1 U15732 ( .A(n13705), .ZN(n13706) );
  AOI21_X1 U15733 ( .B1(n13708), .B2(n13707), .A(n13706), .ZN(n13714) );
  OAI22_X1 U15734 ( .A1(n14496), .A2(n14154), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13709), .ZN(n13711) );
  NOR2_X1 U15735 ( .A1(n14156), .A2(n14577), .ZN(n13710) );
  AOI211_X1 U15736 ( .C1(n13794), .C2(n13712), .A(n13711), .B(n13710), .ZN(
        n13713) );
  OAI21_X1 U15737 ( .B1(n13714), .B2(n14565), .A(n13713), .ZN(P1_U3226) );
  XNOR2_X1 U15738 ( .A(n13717), .B(n13716), .ZN(n13718) );
  XNOR2_X1 U15739 ( .A(n13715), .B(n13718), .ZN(n13726) );
  AOI21_X1 U15740 ( .B1(n14512), .B2(n14038), .A(n13719), .ZN(n13722) );
  NAND2_X1 U15741 ( .A1(n13794), .A2(n13720), .ZN(n13721) );
  OAI211_X1 U15742 ( .C1(n13792), .C2(n13723), .A(n13722), .B(n13721), .ZN(
        n13724) );
  AOI21_X1 U15743 ( .B1(n14150), .B2(n13739), .A(n13724), .ZN(n13725) );
  OAI21_X1 U15744 ( .B1(n13726), .B2(n14565), .A(n13725), .ZN(P1_U3228) );
  INV_X1 U15745 ( .A(n13727), .ZN(n13729) );
  NOR3_X1 U15746 ( .A1(n13730), .A2(n13729), .A3(n13728), .ZN(n13732) );
  OAI21_X1 U15747 ( .B1(n13732), .B2(n13731), .A(n14580), .ZN(n13736) );
  AOI22_X1 U15748 ( .A1(n14510), .A2(n13958), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13733) );
  OAI21_X1 U15749 ( .B1(n13779), .B2(n13791), .A(n13733), .ZN(n13734) );
  AOI21_X1 U15750 ( .B1(n13967), .B2(n13794), .A(n13734), .ZN(n13735) );
  OAI211_X1 U15751 ( .C1(n7220), .C2(n14577), .A(n13736), .B(n13735), .ZN(
        P1_U3229) );
  XOR2_X1 U15752 ( .A(n13737), .B(n13738), .Z(n13745) );
  NAND2_X1 U15753 ( .A1(n14130), .A2(n13739), .ZN(n13743) );
  NAND2_X1 U15754 ( .A1(n13802), .A2(n14050), .ZN(n13741) );
  NAND2_X1 U15755 ( .A1(n14051), .A2(n14339), .ZN(n13740) );
  NAND2_X1 U15756 ( .A1(n13741), .A2(n13740), .ZN(n14021) );
  AOI22_X1 U15757 ( .A1(n14584), .A2(n14021), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13742) );
  OAI211_X1 U15758 ( .C1(n14572), .C2(n14025), .A(n13743), .B(n13742), .ZN(
        n13744) );
  AOI21_X1 U15759 ( .B1(n13745), .B2(n14580), .A(n13744), .ZN(n13746) );
  INV_X1 U15760 ( .A(n13746), .ZN(P1_U3233) );
  OAI211_X1 U15761 ( .C1(n13749), .C2(n13748), .A(n13747), .B(n14580), .ZN(
        n13757) );
  NAND2_X1 U15762 ( .A1(n14510), .A2(n14511), .ZN(n13752) );
  INV_X1 U15763 ( .A(n13750), .ZN(n13751) );
  OAI211_X1 U15764 ( .C1(n13753), .C2(n13791), .A(n13752), .B(n13751), .ZN(
        n13755) );
  NOR2_X1 U15765 ( .A1(n14572), .A2(n14340), .ZN(n13754) );
  NOR2_X1 U15766 ( .A1(n13755), .A2(n13754), .ZN(n13756) );
  OAI211_X1 U15767 ( .C1(n14526), .C2(n14577), .A(n13757), .B(n13756), .ZN(
        P1_U3234) );
  NOR3_X1 U15768 ( .A1(n6468), .A2(n6660), .A3(n13759), .ZN(n13761) );
  OAI21_X1 U15769 ( .B1(n13761), .B2(n13760), .A(n14580), .ZN(n13765) );
  AND2_X1 U15770 ( .A1(n13958), .A2(n14050), .ZN(n13762) );
  AOI21_X1 U15771 ( .B1(n13802), .B2(n14339), .A(n13762), .ZN(n14117) );
  OAI22_X1 U15772 ( .A1(n14496), .A2(n14117), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15165), .ZN(n13763) );
  AOI21_X1 U15773 ( .B1(n13994), .B2(n13794), .A(n13763), .ZN(n13764) );
  OAI211_X1 U15774 ( .C1(n14577), .C2(n14119), .A(n13765), .B(n13764), .ZN(
        P1_U3235) );
  AOI21_X1 U15775 ( .B1(n13768), .B2(n13766), .A(n13767), .ZN(n13774) );
  NAND2_X1 U15776 ( .A1(n14510), .A2(n14052), .ZN(n13769) );
  NAND2_X1 U15777 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13857)
         );
  OAI211_X1 U15778 ( .C1(n13770), .C2(n13791), .A(n13769), .B(n13857), .ZN(
        n13772) );
  NOR2_X1 U15779 ( .A1(n14064), .A2(n14577), .ZN(n13771) );
  AOI211_X1 U15780 ( .C1(n13794), .C2(n14061), .A(n13772), .B(n13771), .ZN(
        n13773) );
  OAI21_X1 U15781 ( .B1(n13774), .B2(n14565), .A(n13773), .ZN(P1_U3238) );
  OAI21_X1 U15782 ( .B1(n13777), .B2(n13776), .A(n13775), .ZN(n13784) );
  NAND2_X1 U15783 ( .A1(n13921), .A2(n14740), .ZN(n14092) );
  NAND2_X1 U15784 ( .A1(n13801), .A2(n14050), .ZN(n13778) );
  OAI21_X1 U15785 ( .B1(n13779), .B2(n14622), .A(n13778), .ZN(n13930) );
  AOI22_X1 U15786 ( .A1(n14584), .A2(n13930), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13781) );
  NAND2_X1 U15787 ( .A1(n13794), .A2(n13924), .ZN(n13780) );
  OAI211_X1 U15788 ( .C1(n14092), .C2(n13782), .A(n13781), .B(n13780), .ZN(
        n13783) );
  AOI21_X1 U15789 ( .B1(n13784), .B2(n14580), .A(n13783), .ZN(n13785) );
  INV_X1 U15790 ( .A(n13785), .ZN(P1_U3240) );
  OAI211_X1 U15791 ( .C1(n13788), .C2(n13787), .A(n13786), .B(n14580), .ZN(
        n13797) );
  NAND2_X1 U15792 ( .A1(n14510), .A2(n14338), .ZN(n13790) );
  OAI211_X1 U15793 ( .C1(n13792), .C2(n13791), .A(n13790), .B(n13789), .ZN(
        n13793) );
  AOI21_X1 U15794 ( .B1(n13795), .B2(n13794), .A(n13793), .ZN(n13796) );
  OAI211_X1 U15795 ( .C1(n14162), .C2(n14577), .A(n13797), .B(n13796), .ZN(
        P1_U3241) );
  MUX2_X1 U15796 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13798), .S(n13812), .Z(
        P1_U3590) );
  MUX2_X1 U15797 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13799), .S(n13812), .Z(
        P1_U3589) );
  MUX2_X1 U15798 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13800), .S(n13812), .Z(
        P1_U3588) );
  MUX2_X1 U15799 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13801), .S(n13812), .Z(
        P1_U3587) );
  MUX2_X1 U15800 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13944), .S(n13812), .Z(
        P1_U3586) );
  MUX2_X1 U15801 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13959), .S(n13812), .Z(
        P1_U3585) );
  MUX2_X1 U15802 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13958), .S(n13812), .Z(
        P1_U3583) );
  MUX2_X1 U15803 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14004), .S(n13812), .Z(
        P1_U3582) );
  MUX2_X1 U15804 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13802), .S(n13812), .Z(
        P1_U3581) );
  MUX2_X1 U15805 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14052), .S(n13812), .Z(
        P1_U3577) );
  MUX2_X1 U15806 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13803), .S(n13812), .Z(
        P1_U3576) );
  MUX2_X1 U15807 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14484), .S(n13812), .Z(
        P1_U3575) );
  MUX2_X1 U15808 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14338), .S(n13812), .Z(
        P1_U3574) );
  MUX2_X1 U15809 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14483), .S(n13812), .Z(
        P1_U3573) );
  MUX2_X1 U15810 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14511), .S(n13812), .Z(
        P1_U3572) );
  MUX2_X1 U15811 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13804), .S(n13812), .Z(
        P1_U3571) );
  MUX2_X1 U15812 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14509), .S(n13812), .Z(
        P1_U3570) );
  MUX2_X1 U15813 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13805), .S(n13812), .Z(
        P1_U3569) );
  MUX2_X1 U15814 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13806), .S(n13812), .Z(
        P1_U3568) );
  MUX2_X1 U15815 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13807), .S(n13812), .Z(
        P1_U3567) );
  MUX2_X1 U15816 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13808), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15817 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13809), .S(n13812), .Z(
        P1_U3565) );
  MUX2_X1 U15818 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13810), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15819 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13811), .S(n13812), .Z(
        P1_U3563) );
  MUX2_X1 U15820 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n8828), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15821 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6863), .S(n13812), .Z(
        P1_U3561) );
  MUX2_X1 U15822 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13813), .S(P1_U4016), .Z(
        P1_U3560) );
  AND2_X1 U15823 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n13816) );
  NOR2_X1 U15824 ( .A1(n14601), .A2(n13814), .ZN(n13815) );
  AOI211_X1 U15825 ( .C1(n13852), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n13816), .B(
        n13815), .ZN(n13825) );
  OAI211_X1 U15826 ( .C1(n13819), .C2(n13818), .A(n14591), .B(n13817), .ZN(
        n13824) );
  AOI211_X1 U15827 ( .C1(n13821), .C2(n13820), .A(n13838), .B(n14596), .ZN(
        n13822) );
  INV_X1 U15828 ( .A(n13822), .ZN(n13823) );
  NAND3_X1 U15829 ( .A1(n13825), .A2(n13824), .A3(n13823), .ZN(P1_U3246) );
  NOR2_X1 U15830 ( .A1(n14601), .A2(n13826), .ZN(n13827) );
  AOI211_X1 U15831 ( .C1(n13852), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n13828), .B(
        n13827), .ZN(n13841) );
  OAI211_X1 U15832 ( .C1(n13831), .C2(n13830), .A(n14591), .B(n13829), .ZN(
        n13840) );
  MUX2_X1 U15833 ( .A(n10017), .B(P1_REG2_REG_4__SCAN_IN), .S(n13832), .Z(
        n13835) );
  INV_X1 U15834 ( .A(n13833), .ZN(n13834) );
  NAND2_X1 U15835 ( .A1(n13835), .A2(n13834), .ZN(n13837) );
  OAI211_X1 U15836 ( .C1(n13838), .C2(n13837), .A(n13887), .B(n13836), .ZN(
        n13839) );
  NAND4_X1 U15837 ( .A1(n13842), .A2(n13841), .A3(n13840), .A4(n13839), .ZN(
        P1_U3247) );
  OAI211_X1 U15838 ( .C1(n13845), .C2(n13844), .A(n13887), .B(n13843), .ZN(
        n13856) );
  NAND2_X1 U15839 ( .A1(n13860), .A2(n13846), .ZN(n13855) );
  OAI21_X1 U15840 ( .B1(n13849), .B2(n13848), .A(n13847), .ZN(n13850) );
  NAND2_X1 U15841 ( .A1(n14591), .A2(n13850), .ZN(n13854) );
  NAND2_X1 U15842 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14488)
         );
  INV_X1 U15843 ( .A(n14488), .ZN(n13851) );
  AOI21_X1 U15844 ( .B1(n13852), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n13851), 
        .ZN(n13853) );
  NAND4_X1 U15845 ( .A1(n13856), .A2(n13855), .A3(n13854), .A4(n13853), .ZN(
        P1_U3257) );
  INV_X1 U15846 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n13858) );
  OAI21_X1 U15847 ( .B1(n14605), .B2(n13858), .A(n13857), .ZN(n13859) );
  AOI21_X1 U15848 ( .B1(n13880), .B2(n13860), .A(n13859), .ZN(n13872) );
  XNOR2_X1 U15849 ( .A(n13873), .B(n13874), .ZN(n13863) );
  INV_X1 U15850 ( .A(n13863), .ZN(n13865) );
  INV_X1 U15851 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n15302) );
  NOR2_X1 U15852 ( .A1(n15302), .A2(n13863), .ZN(n13876) );
  INV_X1 U15853 ( .A(n13876), .ZN(n13864) );
  OAI211_X1 U15854 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n13865), .A(n14591), 
        .B(n13864), .ZN(n13871) );
  OAI21_X1 U15855 ( .B1(n13868), .B2(n13867), .A(n13866), .ZN(n13879) );
  XNOR2_X1 U15856 ( .A(n13873), .B(n13879), .ZN(n13869) );
  NAND2_X1 U15857 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n13869), .ZN(n13881) );
  OAI211_X1 U15858 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n13869), .A(n13887), 
        .B(n13881), .ZN(n13870) );
  NAND3_X1 U15859 ( .A1(n13872), .A2(n13871), .A3(n13870), .ZN(P1_U3261) );
  NOR2_X1 U15860 ( .A1(n13874), .A2(n13873), .ZN(n13875) );
  INV_X1 U15861 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13877) );
  XOR2_X1 U15862 ( .A(n13878), .B(n13877), .Z(n13888) );
  INV_X1 U15863 ( .A(n13888), .ZN(n13885) );
  NAND2_X1 U15864 ( .A1(n13880), .A2(n13879), .ZN(n13882) );
  NAND2_X1 U15865 ( .A1(n13882), .A2(n13881), .ZN(n13883) );
  XOR2_X1 U15866 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n13883), .Z(n13886) );
  OAI21_X1 U15867 ( .B1(n13886), .B2(n14596), .A(n14601), .ZN(n13884) );
  AOI21_X1 U15868 ( .B1(n13885), .B2(n14591), .A(n13884), .ZN(n13890) );
  AOI22_X1 U15869 ( .A1(n13888), .A2(n14591), .B1(n13887), .B2(n13886), .ZN(
        n13889) );
  OAI211_X1 U15870 ( .C1(n13893), .C2(n14605), .A(n13892), .B(n13891), .ZN(
        P1_U3262) );
  NAND2_X1 U15871 ( .A1(n14072), .A2(n13901), .ZN(n13894) );
  XNOR2_X1 U15872 ( .A(n14069), .B(n13894), .ZN(n13895) );
  NAND2_X1 U15873 ( .A1(n13895), .A2(n14637), .ZN(n14068) );
  NAND2_X1 U15874 ( .A1(n13897), .A2(n13896), .ZN(n14070) );
  NOR2_X1 U15875 ( .A1(n14646), .A2(n14070), .ZN(n13904) );
  NOR2_X1 U15876 ( .A1(n14069), .A2(n14640), .ZN(n13898) );
  AOI211_X1 U15877 ( .C1(n14646), .C2(P1_REG2_REG_31__SCAN_IN), .A(n13904), 
        .B(n13898), .ZN(n13899) );
  OAI21_X1 U15878 ( .B1(n14068), .B2(n14639), .A(n13899), .ZN(P1_U3263) );
  XNOR2_X1 U15879 ( .A(n13901), .B(n13900), .ZN(n13902) );
  NAND2_X1 U15880 ( .A1(n13902), .A2(n14637), .ZN(n14071) );
  NOR2_X1 U15881 ( .A1(n14072), .A2(n14640), .ZN(n13903) );
  AOI211_X1 U15882 ( .C1(n14646), .C2(P1_REG2_REG_30__SCAN_IN), .A(n13904), 
        .B(n13903), .ZN(n13905) );
  OAI21_X1 U15883 ( .B1(n14639), .B2(n14071), .A(n13905), .ZN(P1_U3264) );
  OAI21_X1 U15884 ( .B1(n13908), .B2(n13907), .A(n13906), .ZN(n14085) );
  AOI21_X1 U15885 ( .B1(n13909), .B2(n14082), .A(n14058), .ZN(n13911) );
  AOI22_X1 U15886 ( .A1(n14610), .A2(n14081), .B1(n13912), .B2(n14636), .ZN(
        n13914) );
  NAND2_X1 U15887 ( .A1(n14646), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n13913) );
  OAI211_X1 U15888 ( .C1(n6883), .C2(n14640), .A(n13914), .B(n13913), .ZN(
        n13915) );
  AOI21_X1 U15889 ( .B1(n14080), .B2(n13991), .A(n13915), .ZN(n13919) );
  XNOR2_X1 U15890 ( .A(n13917), .B(n13916), .ZN(n14083) );
  NAND2_X1 U15891 ( .A1(n14083), .A2(n14045), .ZN(n13918) );
  OAI211_X1 U15892 ( .C1(n14085), .C2(n14352), .A(n13919), .B(n13918), .ZN(
        P1_U3265) );
  XNOR2_X1 U15893 ( .A(n6555), .B(n13920), .ZN(n14096) );
  INV_X1 U15894 ( .A(n14096), .ZN(n13935) );
  AOI21_X1 U15895 ( .B1(n13942), .B2(n13921), .A(n14058), .ZN(n13923) );
  NAND2_X1 U15896 ( .A1(n13923), .A2(n13922), .ZN(n14091) );
  INV_X1 U15897 ( .A(n14091), .ZN(n13933) );
  AOI22_X1 U15898 ( .A1(n14646), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n13924), 
        .B2(n14636), .ZN(n13925) );
  OAI21_X1 U15899 ( .B1(n6903), .B2(n14640), .A(n13925), .ZN(n13932) );
  OAI21_X1 U15900 ( .B1(n13928), .B2(n13927), .A(n13926), .ZN(n13929) );
  NAND2_X1 U15901 ( .A1(n13929), .A2(n14138), .ZN(n14094) );
  INV_X1 U15902 ( .A(n13930), .ZN(n14093) );
  AOI21_X1 U15903 ( .B1(n14094), .B2(n14093), .A(n14646), .ZN(n13931) );
  AOI211_X1 U15904 ( .C1(n13933), .C2(n14060), .A(n13932), .B(n13931), .ZN(
        n13934) );
  OAI21_X1 U15905 ( .B1(n13935), .B2(n14352), .A(n13934), .ZN(P1_U3267) );
  XNOR2_X1 U15906 ( .A(n13939), .B(n13936), .ZN(n14104) );
  AOI21_X1 U15907 ( .B1(n13939), .B2(n13938), .A(n13937), .ZN(n14102) );
  AOI21_X1 U15908 ( .B1(n13940), .B2(n13965), .A(n14058), .ZN(n13941) );
  NAND2_X1 U15909 ( .A1(n13942), .A2(n13941), .ZN(n14099) );
  AOI22_X1 U15910 ( .A1(n13944), .A2(n14050), .B1(n14339), .B2(n13943), .ZN(
        n14098) );
  INV_X1 U15911 ( .A(n13945), .ZN(n13946) );
  OAI22_X1 U15912 ( .A1(n14646), .A2(n14098), .B1(n13946), .B2(n14608), .ZN(
        n13948) );
  NOR2_X1 U15913 ( .A1(n14100), .A2(n14640), .ZN(n13947) );
  AOI211_X1 U15914 ( .C1(n14646), .C2(P1_REG2_REG_25__SCAN_IN), .A(n13948), 
        .B(n13947), .ZN(n13949) );
  OAI21_X1 U15915 ( .B1(n14639), .B2(n14099), .A(n13949), .ZN(n13950) );
  AOI21_X1 U15916 ( .B1(n14102), .B2(n14618), .A(n13950), .ZN(n13951) );
  OAI21_X1 U15917 ( .B1(n14351), .B2(n14104), .A(n13951), .ZN(P1_U3268) );
  OAI21_X1 U15918 ( .B1(n13954), .B2(n13953), .A(n13952), .ZN(n14105) );
  NAND2_X1 U15919 ( .A1(n14105), .A2(n14056), .ZN(n13963) );
  OAI211_X1 U15920 ( .C1(n13957), .C2(n13956), .A(n13955), .B(n14138), .ZN(
        n13961) );
  AOI22_X1 U15921 ( .A1(n13959), .A2(n14050), .B1(n14339), .B2(n13958), .ZN(
        n13960) );
  AND2_X1 U15922 ( .A1(n13961), .A2(n13960), .ZN(n13962) );
  NAND2_X1 U15923 ( .A1(n13963), .A2(n13962), .ZN(n14108) );
  INV_X1 U15924 ( .A(n14108), .ZN(n13972) );
  AOI21_X1 U15925 ( .B1(n13964), .B2(n13978), .A(n14058), .ZN(n13966) );
  NAND2_X1 U15926 ( .A1(n13966), .A2(n13965), .ZN(n14106) );
  NOR2_X1 U15927 ( .A1(n14106), .A2(n14639), .ZN(n13970) );
  AOI22_X1 U15928 ( .A1(n14646), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n13967), 
        .B2(n14636), .ZN(n13968) );
  OAI21_X1 U15929 ( .B1(n7220), .B2(n14640), .A(n13968), .ZN(n13969) );
  AOI211_X1 U15930 ( .C1(n14105), .C2(n14066), .A(n13970), .B(n13969), .ZN(
        n13971) );
  OAI21_X1 U15931 ( .B1(n13972), .B2(n14646), .A(n13971), .ZN(P1_U3269) );
  OAI21_X1 U15932 ( .B1(n6568), .B2(n12356), .A(n13973), .ZN(n14116) );
  OAI21_X1 U15933 ( .B1(n13976), .B2(n13975), .A(n13974), .ZN(n14114) );
  INV_X1 U15934 ( .A(n13993), .ZN(n13977) );
  AOI21_X1 U15935 ( .B1(n13977), .B2(n8838), .A(n14058), .ZN(n13979) );
  NAND2_X1 U15936 ( .A1(n13979), .A2(n13978), .ZN(n14111) );
  INV_X1 U15937 ( .A(n13980), .ZN(n13981) );
  OAI22_X1 U15938 ( .A1(n14646), .A2(n14110), .B1(n13981), .B2(n14608), .ZN(
        n13983) );
  NOR2_X1 U15939 ( .A1(n14112), .A2(n14640), .ZN(n13982) );
  AOI211_X1 U15940 ( .C1(n14646), .C2(P1_REG2_REG_23__SCAN_IN), .A(n13983), 
        .B(n13982), .ZN(n13984) );
  OAI21_X1 U15941 ( .B1(n14639), .B2(n14111), .A(n13984), .ZN(n13985) );
  AOI21_X1 U15942 ( .B1(n14045), .B2(n14114), .A(n13985), .ZN(n13986) );
  OAI21_X1 U15943 ( .B1(n14352), .B2(n14116), .A(n13986), .ZN(P1_U3270) );
  XOR2_X1 U15944 ( .A(n13987), .B(n13989), .Z(n14123) );
  OAI21_X1 U15945 ( .B1(n13990), .B2(n13989), .A(n13988), .ZN(n14121) );
  INV_X1 U15946 ( .A(n13991), .ZN(n13999) );
  OAI21_X1 U15947 ( .B1(n14119), .B2(n14015), .A(n14637), .ZN(n13992) );
  OR2_X1 U15948 ( .A1(n13993), .A2(n13992), .ZN(n14118) );
  INV_X1 U15949 ( .A(n13994), .ZN(n13995) );
  OAI22_X1 U15950 ( .A1(n14646), .A2(n14117), .B1(n13995), .B2(n14608), .ZN(
        n13997) );
  NOR2_X1 U15951 ( .A1(n14119), .A2(n14640), .ZN(n13996) );
  AOI211_X1 U15952 ( .C1(n14646), .C2(P1_REG2_REG_22__SCAN_IN), .A(n13997), 
        .B(n13996), .ZN(n13998) );
  OAI21_X1 U15953 ( .B1(n13999), .B2(n14118), .A(n13998), .ZN(n14000) );
  AOI21_X1 U15954 ( .B1(n14618), .B2(n14121), .A(n14000), .ZN(n14001) );
  OAI21_X1 U15955 ( .B1(n14123), .B2(n14351), .A(n14001), .ZN(P1_U3271) );
  XOR2_X1 U15956 ( .A(n14002), .B(n14008), .Z(n14003) );
  AOI222_X1 U15957 ( .A1(n14039), .A2(n14339), .B1(n14004), .B2(n14050), .C1(
        n14138), .C2(n14003), .ZN(n14127) );
  INV_X1 U15958 ( .A(n14006), .ZN(n14007) );
  AOI21_X1 U15959 ( .B1(n14008), .B2(n14005), .A(n14007), .ZN(n14128) );
  INV_X1 U15960 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14010) );
  OAI22_X1 U15961 ( .A1(n14610), .A2(n14010), .B1(n14009), .B2(n14608), .ZN(
        n14011) );
  AOI21_X1 U15962 ( .B1(n14012), .B2(n14613), .A(n14011), .ZN(n14017) );
  NAND2_X1 U15963 ( .A1(n14012), .A2(n14028), .ZN(n14013) );
  NAND2_X1 U15964 ( .A1(n14013), .A2(n14637), .ZN(n14014) );
  NOR2_X1 U15965 ( .A1(n14015), .A2(n14014), .ZN(n14125) );
  NAND2_X1 U15966 ( .A1(n14125), .A2(n14060), .ZN(n14016) );
  OAI211_X1 U15967 ( .C1(n14128), .C2(n14352), .A(n14017), .B(n14016), .ZN(
        n14018) );
  INV_X1 U15968 ( .A(n14018), .ZN(n14019) );
  OAI21_X1 U15969 ( .B1(n14127), .B2(n14646), .A(n14019), .ZN(P1_U3272) );
  AOI21_X1 U15970 ( .B1(n14020), .B2(n12350), .A(n14621), .ZN(n14022) );
  AOI21_X1 U15971 ( .B1(n14023), .B2(n14022), .A(n14021), .ZN(n14132) );
  OAI21_X1 U15972 ( .B1(n7570), .B2(n12350), .A(n14024), .ZN(n14133) );
  INV_X1 U15973 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14026) );
  OAI22_X1 U15974 ( .A1(n14610), .A2(n14026), .B1(n14025), .B2(n14608), .ZN(
        n14027) );
  AOI21_X1 U15975 ( .B1(n14130), .B2(n14613), .A(n14027), .ZN(n14031) );
  AOI21_X1 U15976 ( .B1(n14130), .B2(n14037), .A(n14058), .ZN(n14029) );
  AND2_X1 U15977 ( .A1(n14029), .A2(n14028), .ZN(n14129) );
  NAND2_X1 U15978 ( .A1(n14129), .A2(n14060), .ZN(n14030) );
  OAI211_X1 U15979 ( .C1(n14133), .C2(n14352), .A(n14031), .B(n14030), .ZN(
        n14032) );
  INV_X1 U15980 ( .A(n14032), .ZN(n14033) );
  OAI21_X1 U15981 ( .B1(n14646), .B2(n14132), .A(n14033), .ZN(P1_U3273) );
  XNOR2_X1 U15982 ( .A(n14034), .B(n7266), .ZN(n14141) );
  OAI21_X1 U15983 ( .B1(n7574), .B2(n14036), .A(n14035), .ZN(n14139) );
  OAI211_X1 U15984 ( .C1(n14136), .C2(n14057), .A(n14637), .B(n14037), .ZN(
        n14135) );
  AOI22_X1 U15985 ( .A1(n14039), .A2(n14050), .B1(n14339), .B2(n14038), .ZN(
        n14134) );
  OAI22_X1 U15986 ( .A1(n14646), .A2(n14134), .B1(n14040), .B2(n14608), .ZN(
        n14042) );
  NOR2_X1 U15987 ( .A1(n14136), .A2(n14640), .ZN(n14041) );
  AOI211_X1 U15988 ( .C1(n14646), .C2(P1_REG2_REG_19__SCAN_IN), .A(n14042), 
        .B(n14041), .ZN(n14043) );
  OAI21_X1 U15989 ( .B1(n14639), .B2(n14135), .A(n14043), .ZN(n14044) );
  AOI21_X1 U15990 ( .B1(n14139), .B2(n14045), .A(n14044), .ZN(n14046) );
  OAI21_X1 U15991 ( .B1(n14141), .B2(n14352), .A(n14046), .ZN(P1_U3274) );
  XNOR2_X1 U15992 ( .A(n14047), .B(n14048), .ZN(n14142) );
  XNOR2_X1 U15993 ( .A(n14049), .B(n14048), .ZN(n14054) );
  AOI22_X1 U15994 ( .A1(n14339), .A2(n14052), .B1(n14051), .B2(n14050), .ZN(
        n14053) );
  OAI21_X1 U15995 ( .B1(n14054), .B2(n14621), .A(n14053), .ZN(n14055) );
  AOI21_X1 U15996 ( .B1(n14142), .B2(n14056), .A(n14055), .ZN(n14146) );
  AOI211_X1 U15997 ( .C1(n14144), .C2(n14059), .A(n14058), .B(n14057), .ZN(
        n14143) );
  NAND2_X1 U15998 ( .A1(n14143), .A2(n14060), .ZN(n14063) );
  AOI22_X1 U15999 ( .A1(n14646), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14061), 
        .B2(n14636), .ZN(n14062) );
  OAI211_X1 U16000 ( .C1(n14064), .C2(n14640), .A(n14063), .B(n14062), .ZN(
        n14065) );
  AOI21_X1 U16001 ( .B1(n14142), .B2(n14066), .A(n14065), .ZN(n14067) );
  OAI21_X1 U16002 ( .B1(n14146), .B2(n14646), .A(n14067), .ZN(P1_U3275) );
  OAI211_X1 U16003 ( .C1(n14069), .C2(n14711), .A(n14068), .B(n14070), .ZN(
        n14169) );
  MUX2_X1 U16004 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14169), .S(n14748), .Z(
        P1_U3559) );
  OAI211_X1 U16005 ( .C1(n14072), .C2(n14711), .A(n14071), .B(n14070), .ZN(
        n14170) );
  MUX2_X1 U16006 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14170), .S(n14748), .Z(
        P1_U3558) );
  OAI211_X1 U16007 ( .C1(n7229), .C2(n14711), .A(n14074), .B(n14073), .ZN(
        n14075) );
  MUX2_X1 U16008 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14171), .S(n14748), .Z(
        P1_U3557) );
  NAND2_X1 U16009 ( .A1(n14083), .A2(n14138), .ZN(n14084) );
  MUX2_X1 U16010 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14172), .S(n14748), .Z(
        P1_U3556) );
  AOI21_X1 U16011 ( .B1(n14740), .B2(n14087), .A(n14086), .ZN(n14088) );
  OAI211_X1 U16012 ( .C1(n14090), .C2(n14743), .A(n14089), .B(n14088), .ZN(
        n14173) );
  MUX2_X1 U16013 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14173), .S(n14748), .Z(
        P1_U3555) );
  NAND4_X1 U16014 ( .A1(n14094), .A2(n14093), .A3(n14092), .A4(n14091), .ZN(
        n14095) );
  AOI21_X1 U16015 ( .B1(n14096), .B2(n14729), .A(n14095), .ZN(n14097) );
  INV_X1 U16016 ( .A(n14097), .ZN(n14174) );
  MUX2_X1 U16017 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14174), .S(n14748), .Z(
        P1_U3554) );
  OAI211_X1 U16018 ( .C1(n14100), .C2(n14711), .A(n14099), .B(n14098), .ZN(
        n14101) );
  AOI21_X1 U16019 ( .B1(n14102), .B2(n14729), .A(n14101), .ZN(n14103) );
  OAI21_X1 U16020 ( .B1(n14621), .B2(n14104), .A(n14103), .ZN(n14175) );
  MUX2_X1 U16021 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14175), .S(n14748), .Z(
        P1_U3553) );
  INV_X1 U16022 ( .A(n14743), .ZN(n14687) );
  NAND2_X1 U16023 ( .A1(n14105), .A2(n14687), .ZN(n14107) );
  OAI211_X1 U16024 ( .C1(n7220), .C2(n14711), .A(n14107), .B(n14106), .ZN(
        n14109) );
  MUX2_X1 U16025 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14176), .S(n14748), .Z(
        P1_U3552) );
  OAI211_X1 U16026 ( .C1(n14112), .C2(n14711), .A(n14111), .B(n14110), .ZN(
        n14113) );
  AOI21_X1 U16027 ( .B1(n14114), .B2(n14138), .A(n14113), .ZN(n14115) );
  OAI21_X1 U16028 ( .B1(n14116), .B2(n14153), .A(n14115), .ZN(n14177) );
  MUX2_X1 U16029 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14177), .S(n14748), .Z(
        P1_U3551) );
  OAI211_X1 U16030 ( .C1(n14711), .C2(n14119), .A(n14118), .B(n14117), .ZN(
        n14120) );
  AOI21_X1 U16031 ( .B1(n14121), .B2(n14729), .A(n14120), .ZN(n14122) );
  OAI21_X1 U16032 ( .B1(n14621), .B2(n14123), .A(n14122), .ZN(n14178) );
  MUX2_X1 U16033 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14178), .S(n14748), .Z(
        P1_U3550) );
  NOR2_X1 U16034 ( .A1(n14125), .A2(n14124), .ZN(n14126) );
  OAI211_X1 U16035 ( .C1(n14153), .C2(n14128), .A(n14127), .B(n14126), .ZN(
        n14179) );
  MUX2_X1 U16036 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14179), .S(n14748), .Z(
        P1_U3549) );
  AOI21_X1 U16037 ( .B1(n14740), .B2(n14130), .A(n14129), .ZN(n14131) );
  OAI211_X1 U16038 ( .C1(n14133), .C2(n14153), .A(n14132), .B(n14131), .ZN(
        n14180) );
  MUX2_X1 U16039 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14180), .S(n14748), .Z(
        P1_U3548) );
  OAI211_X1 U16040 ( .C1(n14136), .C2(n14711), .A(n14135), .B(n14134), .ZN(
        n14137) );
  AOI21_X1 U16041 ( .B1(n14139), .B2(n14138), .A(n14137), .ZN(n14140) );
  OAI21_X1 U16042 ( .B1(n14141), .B2(n14153), .A(n14140), .ZN(n14181) );
  MUX2_X1 U16043 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14181), .S(n14748), .Z(
        P1_U3547) );
  INV_X1 U16044 ( .A(n14142), .ZN(n14147) );
  AOI21_X1 U16045 ( .B1(n14740), .B2(n14144), .A(n14143), .ZN(n14145) );
  OAI211_X1 U16046 ( .C1(n14147), .C2(n14743), .A(n14146), .B(n14145), .ZN(
        n14182) );
  MUX2_X1 U16047 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14182), .S(n14748), .Z(
        P1_U3546) );
  AOI211_X1 U16048 ( .C1(n14740), .C2(n14150), .A(n14149), .B(n14148), .ZN(
        n14151) );
  OAI21_X1 U16049 ( .B1(n14153), .B2(n14152), .A(n14151), .ZN(n14183) );
  MUX2_X1 U16050 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14183), .S(n14748), .Z(
        P1_U3545) );
  OAI211_X1 U16051 ( .C1(n14156), .C2(n14711), .A(n14155), .B(n14154), .ZN(
        n14157) );
  AOI21_X1 U16052 ( .B1(n14158), .B2(n14729), .A(n14157), .ZN(n14159) );
  OAI21_X1 U16053 ( .B1(n14160), .B2(n14621), .A(n14159), .ZN(n14184) );
  MUX2_X1 U16054 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14184), .S(n14748), .Z(
        P1_U3544) );
  OAI21_X1 U16055 ( .B1(n14162), .B2(n14711), .A(n14161), .ZN(n14163) );
  AOI211_X1 U16056 ( .C1(n14165), .C2(n14729), .A(n14164), .B(n14163), .ZN(
        n14166) );
  OAI21_X1 U16057 ( .B1(n14621), .B2(n14167), .A(n14166), .ZN(n14185) );
  MUX2_X1 U16058 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n14185), .S(n14748), .Z(
        P1_U3543) );
  MUX2_X1 U16059 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n14168), .S(n14748), .Z(
        P1_U3528) );
  MUX2_X1 U16060 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14169), .S(n15160), .Z(
        P1_U3527) );
  MUX2_X1 U16061 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14170), .S(n15160), .Z(
        P1_U3526) );
  MUX2_X1 U16062 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14173), .S(n15160), .Z(
        P1_U3523) );
  MUX2_X1 U16063 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14174), .S(n15160), .Z(
        P1_U3522) );
  MUX2_X1 U16064 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14175), .S(n15160), .Z(
        P1_U3521) );
  MUX2_X1 U16065 ( .A(n14176), .B(P1_REG0_REG_24__SCAN_IN), .S(n15158), .Z(
        P1_U3520) );
  MUX2_X1 U16066 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14177), .S(n15160), .Z(
        P1_U3519) );
  MUX2_X1 U16067 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14178), .S(n15160), .Z(
        P1_U3518) );
  MUX2_X1 U16068 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14179), .S(n15160), .Z(
        P1_U3517) );
  MUX2_X1 U16069 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14180), .S(n15160), .Z(
        P1_U3516) );
  MUX2_X1 U16070 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14181), .S(n15160), .Z(
        P1_U3515) );
  MUX2_X1 U16071 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14182), .S(n15160), .Z(
        P1_U3513) );
  MUX2_X1 U16072 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14183), .S(n15160), .Z(
        P1_U3510) );
  MUX2_X1 U16073 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14184), .S(n15160), .Z(
        P1_U3507) );
  MUX2_X1 U16074 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n14185), .S(n15160), .Z(
        P1_U3504) );
  NOR4_X1 U16075 ( .A1(n14186), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n8589), .ZN(n14187) );
  AOI21_X1 U16076 ( .B1(n14188), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14187), 
        .ZN(n14189) );
  OAI21_X1 U16077 ( .B1(n14190), .B2(n14204), .A(n14189), .ZN(P1_U3324) );
  OAI222_X1 U16078 ( .A1(n14192), .A2(P1_U3086), .B1(n14201), .B2(n7677), .C1(
        n14191), .C2(n14204), .ZN(P1_U3326) );
  INV_X1 U16079 ( .A(n14193), .ZN(n14195) );
  OAI222_X1 U16080 ( .A1(P1_U3086), .A2(n8882), .B1(n14204), .B2(n14195), .C1(
        n14194), .C2(n14201), .ZN(P1_U3327) );
  OAI222_X1 U16081 ( .A1(P1_U3086), .A2(n14197), .B1(n14204), .B2(n14196), 
        .C1(n15193), .C2(n14201), .ZN(P1_U3328) );
  OAI222_X1 U16082 ( .A1(n14201), .A2(n14200), .B1(P1_U3086), .B2(n14199), 
        .C1(n14198), .C2(n14204), .ZN(P1_U3329) );
  INV_X1 U16083 ( .A(n10222), .ZN(n14205) );
  OAI222_X1 U16084 ( .A1(P1_U3086), .A2(n14205), .B1(n14204), .B2(n14203), 
        .C1(n14202), .C2(n14201), .ZN(P1_U3331) );
  MUX2_X1 U16085 ( .A(n14206), .B(n8820), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U16086 ( .A(n14208), .B(n14207), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  INV_X1 U16087 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15298) );
  XOR2_X1 U16088 ( .A(n15298), .B(P1_ADDR_REG_18__SCAN_IN), .Z(n14362) );
  INV_X1 U16089 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14304) );
  NOR2_X1 U16090 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14304), .ZN(n14303) );
  INV_X1 U16091 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14300) );
  AND2_X1 U16092 ( .A1(n14300), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n14240) );
  INV_X1 U16093 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14239) );
  XOR2_X1 U16094 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n14247) );
  INV_X1 U16095 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14248) );
  INV_X1 U16096 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14235) );
  INV_X1 U16097 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14967) );
  INV_X1 U16098 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14231) );
  INV_X1 U16099 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14230) );
  INV_X1 U16100 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14228) );
  NAND2_X1 U16101 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(n14262), .ZN(n14261) );
  XOR2_X1 U16102 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), .Z(
        n14258) );
  NOR2_X1 U16103 ( .A1(n14259), .A2(n14258), .ZN(n14213) );
  XNOR2_X1 U16104 ( .A(n14215), .B(n14214), .ZN(n14257) );
  INV_X1 U16105 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14216) );
  NOR2_X1 U16106 ( .A1(n14217), .A2(n14216), .ZN(n14218) );
  NOR2_X1 U16107 ( .A1(n14221), .A2(n6849), .ZN(n14223) );
  NOR2_X1 U16108 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14225), .ZN(n14226) );
  XOR2_X1 U16109 ( .A(n14225), .B(P3_ADDR_REG_7__SCAN_IN), .Z(n14254) );
  XOR2_X1 U16110 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), .Z(
        n14283) );
  XOR2_X1 U16111 ( .A(n14230), .B(P1_ADDR_REG_9__SCAN_IN), .Z(n14288) );
  NAND2_X1 U16112 ( .A1(n14289), .A2(n14288), .ZN(n14229) );
  NAND2_X1 U16113 ( .A1(n14231), .A2(n14253), .ZN(n14233) );
  NOR2_X1 U16114 ( .A1(n14231), .A2(n14253), .ZN(n14232) );
  XNOR2_X1 U16115 ( .A(P1_ADDR_REG_11__SCAN_IN), .B(n14235), .ZN(n14294) );
  XOR2_X1 U16116 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(n14606), .Z(n14252) );
  AND2_X1 U16117 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14248), .ZN(n14237) );
  OAI22_X1 U16118 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14300), .B1(n14240), 
        .B2(n14302), .ZN(n14306) );
  NAND2_X1 U16119 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14304), .ZN(n14241) );
  OAI21_X1 U16120 ( .B1(n14303), .B2(n14306), .A(n14241), .ZN(n14242) );
  NOR2_X1 U16121 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14242), .ZN(n14244) );
  INV_X1 U16122 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14412) );
  XNOR2_X1 U16123 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14242), .ZN(n14245) );
  NOR2_X1 U16124 ( .A1(n14412), .A2(n14245), .ZN(n14243) );
  NOR2_X1 U16125 ( .A1(n14244), .A2(n14243), .ZN(n14361) );
  XNOR2_X1 U16126 ( .A(n14362), .B(n14361), .ZN(n14365) );
  XOR2_X1 U16127 ( .A(n14412), .B(n14245), .Z(n14358) );
  XNOR2_X1 U16128 ( .A(n14247), .B(n14246), .ZN(n14551) );
  XOR2_X1 U16129 ( .A(n14248), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n14250) );
  XNOR2_X1 U16130 ( .A(n14250), .B(n14249), .ZN(n14547) );
  XOR2_X1 U16131 ( .A(n14252), .B(n14251), .Z(n14295) );
  INV_X1 U16132 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14773) );
  XNOR2_X1 U16133 ( .A(n14254), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15327) );
  XNOR2_X1 U16134 ( .A(n14256), .B(n14255), .ZN(n14270) );
  INV_X1 U16135 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14268) );
  NAND2_X1 U16136 ( .A1(n14267), .A2(n14268), .ZN(n14269) );
  XOR2_X1 U16137 ( .A(n14257), .B(P1_ADDR_REG_3__SCAN_IN), .Z(n15330) );
  XOR2_X1 U16138 ( .A(n14259), .B(n14258), .Z(n14315) );
  XOR2_X1 U16139 ( .A(n14260), .B(n14261), .Z(n14263) );
  NOR2_X1 U16140 ( .A1(n14263), .A2(n9909), .ZN(n14264) );
  OAI21_X1 U16141 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n14262), .A(n14261), .ZN(
        n15324) );
  NAND2_X1 U16142 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15324), .ZN(n15334) );
  XOR2_X1 U16143 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n14263), .Z(n15333) );
  NOR2_X1 U16144 ( .A1(n15334), .A2(n15333), .ZN(n15332) );
  NOR2_X1 U16145 ( .A1(n14264), .A2(n15332), .ZN(n14314) );
  NOR2_X1 U16146 ( .A1(n14315), .A2(n14314), .ZN(n14265) );
  NAND2_X1 U16147 ( .A1(n14315), .A2(n14314), .ZN(n14313) );
  OAI21_X1 U16148 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n14265), .A(n14313), .ZN(
        n15329) );
  NAND2_X1 U16149 ( .A1(n15330), .A2(n15329), .ZN(n14266) );
  NOR2_X1 U16150 ( .A1(n15330), .A2(n15329), .ZN(n15328) );
  AOI21_X1 U16151 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n14266), .A(n15328), .ZN(
        n15320) );
  XOR2_X1 U16152 ( .A(n14268), .B(n14267), .Z(n15319) );
  NAND2_X1 U16153 ( .A1(n14270), .A2(n14272), .ZN(n14273) );
  INV_X1 U16154 ( .A(n14270), .ZN(n14271) );
  INV_X1 U16155 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15322) );
  XNOR2_X1 U16156 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n14274), .ZN(n14275) );
  XOR2_X1 U16157 ( .A(n14276), .B(n14275), .Z(n14325) );
  INV_X1 U16158 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n14277) );
  NOR2_X1 U16159 ( .A1(n14278), .A2(n14277), .ZN(n14279) );
  XNOR2_X1 U16160 ( .A(n14283), .B(n14282), .ZN(n14284) );
  NAND2_X1 U16161 ( .A1(n14286), .A2(n14284), .ZN(n14287) );
  INV_X1 U16162 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14328) );
  XOR2_X1 U16163 ( .A(n14289), .B(n14288), .Z(n14291) );
  NOR2_X1 U16164 ( .A1(n14291), .A2(n14290), .ZN(n14292) );
  XNOR2_X1 U16165 ( .A(n14294), .B(n14293), .ZN(n14541) );
  NAND2_X1 U16166 ( .A1(n14295), .A2(n14296), .ZN(n14297) );
  INV_X1 U16167 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14792) );
  INV_X1 U16168 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14299) );
  XNOR2_X1 U16169 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(n14300), .ZN(n14301) );
  INV_X1 U16170 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14557) );
  AOI21_X1 U16171 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(n14304), .A(n14303), 
        .ZN(n14305) );
  XOR2_X1 U16172 ( .A(n14306), .B(n14305), .Z(n14559) );
  NAND2_X1 U16173 ( .A1(n14358), .A2(n14359), .ZN(n14357) );
  OAI21_X1 U16174 ( .B1(n14365), .B2(n14364), .A(n14366), .ZN(n14310) );
  INV_X1 U16175 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n15255) );
  XOR2_X1 U16176 ( .A(n14310), .B(n15255), .Z(SUB_1596_U62) );
  AOI21_X1 U16177 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14311) );
  OAI21_X1 U16178 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14311), 
        .ZN(U28) );
  AOI21_X1 U16179 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14312) );
  OAI21_X1 U16180 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14312), 
        .ZN(U29) );
  OAI21_X1 U16181 ( .B1(n14315), .B2(n14314), .A(n14313), .ZN(n14316) );
  XNOR2_X1 U16182 ( .A(n14316), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI22_X1 U16183 ( .A1(n14317), .A2(n14320), .B1(SI_11_), .B2(n14319), .ZN(
        n14318) );
  OAI21_X1 U16184 ( .B1(P3_U3151), .B2(n14975), .A(n14318), .ZN(P3_U3284) );
  AOI22_X1 U16185 ( .A1(n14321), .A2(n14320), .B1(SI_12_), .B2(n14319), .ZN(
        n14322) );
  OAI21_X1 U16186 ( .B1(P3_U3151), .B2(n14323), .A(n14322), .ZN(P3_U3283) );
  AOI21_X1 U16187 ( .B1(n14326), .B2(n14325), .A(n14324), .ZN(SUB_1596_U57) );
  OAI21_X1 U16188 ( .B1(n14329), .B2(n14328), .A(n14327), .ZN(SUB_1596_U55) );
  AOI21_X1 U16189 ( .B1(n14773), .B2(n14331), .A(n14330), .ZN(SUB_1596_U54) );
  AOI21_X1 U16190 ( .B1(n14334), .B2(n14333), .A(n14332), .ZN(n14335) );
  XOR2_X1 U16191 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14335), .Z(SUB_1596_U70)
         );
  OAI211_X1 U16192 ( .C1(n14337), .C2(n14526), .A(n14637), .B(n14336), .ZN(
        n14525) );
  AOI22_X1 U16193 ( .A1(n14339), .A2(n14511), .B1(n14338), .B2(n14050), .ZN(
        n14524) );
  OAI21_X1 U16194 ( .B1(n14340), .B2(n14608), .A(n14524), .ZN(n14341) );
  AOI21_X1 U16195 ( .B1(n14343), .B2(n14342), .A(n14341), .ZN(n14344) );
  OAI21_X1 U16196 ( .B1(n14525), .B2(n14345), .A(n14344), .ZN(n14355) );
  OAI21_X1 U16197 ( .B1(n14348), .B2(n14347), .A(n14346), .ZN(n14530) );
  INV_X1 U16198 ( .A(n14530), .ZN(n14353) );
  XNOR2_X1 U16199 ( .A(n14350), .B(n14349), .ZN(n14527) );
  OAI22_X1 U16200 ( .A1(n14353), .A2(n14352), .B1(n14351), .B2(n14527), .ZN(
        n14354) );
  AOI221_X1 U16201 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n14646), .C1(n14355), 
        .C2(n14610), .A(n14354), .ZN(n14356) );
  INV_X1 U16202 ( .A(n14356), .ZN(P1_U3280) );
  OAI21_X1 U16203 ( .B1(n14359), .B2(n14358), .A(n14357), .ZN(n14360) );
  XNOR2_X1 U16204 ( .A(n14360), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  AND2_X1 U16205 ( .A1(n14362), .A2(n14361), .ZN(n14363) );
  AOI21_X1 U16206 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15298), .A(n14363), 
        .ZN(n14368) );
  AOI21_X1 U16207 ( .B1(n14371), .B2(n14370), .A(n14369), .ZN(n14385) );
  OAI21_X1 U16208 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n14373), .A(n14372), 
        .ZN(n14378) );
  AOI21_X1 U16209 ( .B1(n15030), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n14374), 
        .ZN(n14375) );
  OAI21_X1 U16210 ( .B1(n15033), .B2(n14376), .A(n14375), .ZN(n14377) );
  AOI21_X1 U16211 ( .B1(n14378), .B2(n15035), .A(n14377), .ZN(n14384) );
  AOI21_X1 U16212 ( .B1(n14381), .B2(n14380), .A(n14379), .ZN(n14382) );
  OR2_X1 U16213 ( .A1(n14382), .A2(n15018), .ZN(n14383) );
  OAI211_X1 U16214 ( .C1(n14385), .C2(n15043), .A(n14384), .B(n14383), .ZN(
        P3_U3197) );
  AOI21_X1 U16215 ( .B1(n14387), .B2(n14386), .A(n6580), .ZN(n14402) );
  OAI21_X1 U16216 ( .B1(n14390), .B2(n14389), .A(n14388), .ZN(n14395) );
  AOI21_X1 U16217 ( .B1(n15030), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n14391), 
        .ZN(n14392) );
  OAI21_X1 U16218 ( .B1(n15033), .B2(n14393), .A(n14392), .ZN(n14394) );
  AOI21_X1 U16219 ( .B1(n14395), .B2(n15035), .A(n14394), .ZN(n14401) );
  NOR2_X1 U16220 ( .A1(n6605), .A2(n14396), .ZN(n14398) );
  AOI21_X1 U16221 ( .B1(n14399), .B2(n14398), .A(n15018), .ZN(n14397) );
  OAI21_X1 U16222 ( .B1(n14399), .B2(n14398), .A(n14397), .ZN(n14400) );
  OAI211_X1 U16223 ( .C1(n14402), .C2(n15043), .A(n14401), .B(n14400), .ZN(
        P3_U3198) );
  AOI21_X1 U16224 ( .B1(n14405), .B2(n14404), .A(n14403), .ZN(n14419) );
  OAI21_X1 U16225 ( .B1(n14407), .B2(P3_REG1_REG_17__SCAN_IN), .A(n14406), 
        .ZN(n14408) );
  AND2_X1 U16226 ( .A1(n14408), .A2(n15035), .ZN(n14416) );
  AOI211_X1 U16227 ( .C1(n14411), .C2(n14410), .A(n15018), .B(n14409), .ZN(
        n14415) );
  OAI22_X1 U16228 ( .A1(n15033), .A2(n14413), .B1(n14412), .B2(n14996), .ZN(
        n14414) );
  NOR4_X1 U16229 ( .A1(n14417), .A2(n14416), .A3(n14415), .A4(n14414), .ZN(
        n14418) );
  OAI21_X1 U16230 ( .B1(n14419), .B2(n15043), .A(n14418), .ZN(P3_U3199) );
  AOI22_X1 U16231 ( .A1(n14992), .A2(n14420), .B1(n15030), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n14433) );
  OAI21_X1 U16232 ( .B1(n14423), .B2(n14422), .A(n14421), .ZN(n14428) );
  OAI21_X1 U16233 ( .B1(n14426), .B2(n14425), .A(n14424), .ZN(n14427) );
  AOI22_X1 U16234 ( .A1(n14428), .A2(n15035), .B1(n15037), .B2(n14427), .ZN(
        n14432) );
  XNOR2_X1 U16235 ( .A(n14434), .B(n14441), .ZN(n14439) );
  AOI222_X1 U16236 ( .A1(n15089), .A2(n14439), .B1(n14438), .B2(n14437), .C1(
        n14436), .C2(n14435), .ZN(n14463) );
  AOI22_X1 U16237 ( .A1(n15071), .A2(n14440), .B1(n15075), .B2(
        P3_REG2_REG_12__SCAN_IN), .ZN(n14447) );
  XNOR2_X1 U16238 ( .A(n14442), .B(n14441), .ZN(n14466) );
  INV_X1 U16239 ( .A(n14443), .ZN(n14444) );
  NOR2_X1 U16240 ( .A1(n14444), .A2(n15136), .ZN(n14465) );
  AOI22_X1 U16241 ( .A1(n14466), .A2(n14445), .B1(n15072), .B2(n14465), .ZN(
        n14446) );
  OAI211_X1 U16242 ( .C1(n15075), .C2(n14463), .A(n14447), .B(n14446), .ZN(
        P3_U3221) );
  INV_X1 U16243 ( .A(n9486), .ZN(n14449) );
  INV_X1 U16244 ( .A(n14448), .ZN(n14451) );
  AOI21_X1 U16245 ( .B1(n14449), .B2(n15078), .A(n14451), .ZN(n14468) );
  INV_X1 U16246 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n14450) );
  AOI22_X1 U16247 ( .A1(n15157), .A2(n14468), .B1(n14450), .B2(n15154), .ZN(
        P3_U3490) );
  AOI21_X1 U16248 ( .B1(n14452), .B2(n15078), .A(n14451), .ZN(n14470) );
  INV_X1 U16249 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n15217) );
  AOI22_X1 U16250 ( .A1(n15157), .A2(n14470), .B1(n15217), .B2(n15154), .ZN(
        P3_U3489) );
  NOR2_X1 U16251 ( .A1(n14453), .A2(n14458), .ZN(n14455) );
  AOI211_X1 U16252 ( .C1(n15078), .C2(n14456), .A(n14455), .B(n14454), .ZN(
        n14472) );
  AOI22_X1 U16253 ( .A1(n15157), .A2(n14472), .B1(n12615), .B2(n15154), .ZN(
        P3_U3473) );
  OAI22_X1 U16254 ( .A1(n14459), .A2(n14458), .B1(n15136), .B2(n14457), .ZN(
        n14460) );
  NOR2_X1 U16255 ( .A1(n14461), .A2(n14460), .ZN(n14474) );
  INV_X1 U16256 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14462) );
  AOI22_X1 U16257 ( .A1(n15157), .A2(n14474), .B1(n14462), .B2(n15154), .ZN(
        P3_U3472) );
  INV_X1 U16258 ( .A(n14463), .ZN(n14464) );
  AOI211_X1 U16259 ( .C1(n14466), .C2(n15101), .A(n14465), .B(n14464), .ZN(
        n14476) );
  AOI22_X1 U16260 ( .A1(n15157), .A2(n14476), .B1(n14467), .B2(n15154), .ZN(
        P3_U3471) );
  INV_X1 U16261 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14469) );
  AOI22_X1 U16262 ( .A1(n15142), .A2(n14469), .B1(n14468), .B2(n15141), .ZN(
        P3_U3458) );
  INV_X1 U16263 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14471) );
  AOI22_X1 U16264 ( .A1(n15142), .A2(n14471), .B1(n14470), .B2(n15141), .ZN(
        P3_U3457) );
  INV_X1 U16265 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n14473) );
  AOI22_X1 U16266 ( .A1(n15142), .A2(n14473), .B1(n14472), .B2(n15141), .ZN(
        P3_U3432) );
  INV_X1 U16267 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14475) );
  AOI22_X1 U16268 ( .A1(n15142), .A2(n14475), .B1(n14474), .B2(n15141), .ZN(
        P3_U3429) );
  INV_X1 U16269 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14477) );
  AOI22_X1 U16270 ( .A1(n15142), .A2(n14477), .B1(n14476), .B2(n15141), .ZN(
        P3_U3426) );
  INV_X1 U16271 ( .A(n13747), .ZN(n14480) );
  OAI21_X1 U16272 ( .B1(n14480), .B2(n14479), .A(n14478), .ZN(n14482) );
  AOI21_X1 U16273 ( .B1(n14482), .B2(n14481), .A(n14565), .ZN(n14487) );
  AOI22_X1 U16274 ( .A1(n14512), .A2(n14484), .B1(n14510), .B2(n14483), .ZN(
        n14485) );
  OAI21_X1 U16275 ( .B1(n14520), .B2(n14577), .A(n14485), .ZN(n14486) );
  NOR2_X1 U16276 ( .A1(n14487), .A2(n14486), .ZN(n14489) );
  OAI211_X1 U16277 ( .C1(n14490), .C2(n14572), .A(n14489), .B(n14488), .ZN(
        P1_U3215) );
  NAND2_X1 U16278 ( .A1(n14491), .A2(n14740), .ZN(n14724) );
  INV_X1 U16279 ( .A(n14724), .ZN(n14492) );
  AOI22_X1 U16280 ( .A1(n14492), .A2(n14564), .B1(P1_REG3_REG_10__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14502) );
  NAND2_X1 U16281 ( .A1(n14505), .A2(n14494), .ZN(n14495) );
  XNOR2_X1 U16282 ( .A(n14493), .B(n14495), .ZN(n14500) );
  AOI21_X1 U16283 ( .B1(n14498), .B2(n14497), .A(n14496), .ZN(n14499) );
  AOI21_X1 U16284 ( .B1(n14500), .B2(n14580), .A(n14499), .ZN(n14501) );
  OAI211_X1 U16285 ( .C1(n14572), .C2(n14503), .A(n14502), .B(n14501), .ZN(
        P1_U3217) );
  AOI21_X1 U16286 ( .B1(n14506), .B2(n14505), .A(n14504), .ZN(n14507) );
  OAI21_X1 U16287 ( .B1(n14508), .B2(n14507), .A(n14580), .ZN(n14514) );
  AOI22_X1 U16288 ( .A1(n14512), .A2(n14511), .B1(n14510), .B2(n14509), .ZN(
        n14513) );
  OAI211_X1 U16289 ( .C1(n14532), .C2(n14577), .A(n14514), .B(n14513), .ZN(
        n14515) );
  INV_X1 U16290 ( .A(n14515), .ZN(n14517) );
  OAI211_X1 U16291 ( .C1(n14518), .C2(n14572), .A(n14517), .B(n14516), .ZN(
        P1_U3236) );
  OAI21_X1 U16292 ( .B1(n14520), .B2(n14711), .A(n14519), .ZN(n14522) );
  AOI211_X1 U16293 ( .C1(n14523), .C2(n14729), .A(n14522), .B(n14521), .ZN(
        n14536) );
  AOI22_X1 U16294 ( .A1(n14748), .A2(n14536), .B1(n11267), .B2(n14746), .ZN(
        P1_U3542) );
  OAI211_X1 U16295 ( .C1(n14526), .C2(n14711), .A(n14525), .B(n14524), .ZN(
        n14529) );
  NOR2_X1 U16296 ( .A1(n14527), .A2(n14621), .ZN(n14528) );
  AOI211_X1 U16297 ( .C1(n14729), .C2(n14530), .A(n14529), .B(n14528), .ZN(
        n14537) );
  AOI22_X1 U16298 ( .A1(n14748), .A2(n14537), .B1(n10785), .B2(n14746), .ZN(
        P1_U3541) );
  OAI21_X1 U16299 ( .B1(n14532), .B2(n14711), .A(n14531), .ZN(n14534) );
  AOI211_X1 U16300 ( .C1(n14729), .C2(n14535), .A(n14534), .B(n14533), .ZN(
        n14538) );
  AOI22_X1 U16301 ( .A1(n14748), .A2(n14538), .B1(n10296), .B2(n14746), .ZN(
        P1_U3539) );
  AOI22_X1 U16302 ( .A1(n15160), .A2(n14536), .B1(n8555), .B2(n15158), .ZN(
        P1_U3501) );
  AOI22_X1 U16303 ( .A1(n15160), .A2(n14537), .B1(n8535), .B2(n15158), .ZN(
        P1_U3498) );
  AOI22_X1 U16304 ( .A1(n15160), .A2(n14538), .B1(n8506), .B2(n15158), .ZN(
        P1_U3492) );
  OAI21_X1 U16305 ( .B1(n14541), .B2(n14540), .A(n14539), .ZN(n14542) );
  XNOR2_X1 U16306 ( .A(n14542), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI21_X1 U16307 ( .B1(n14544), .B2(n14792), .A(n14543), .ZN(SUB_1596_U68) );
  OAI21_X1 U16308 ( .B1(n14547), .B2(n14546), .A(n14545), .ZN(n14548) );
  XNOR2_X1 U16309 ( .A(n14548), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  OAI21_X1 U16310 ( .B1(n14551), .B2(n14550), .A(n14549), .ZN(n14552) );
  XNOR2_X1 U16311 ( .A(n14552), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI222_X1 U16312 ( .A1(n14557), .A2(n14556), .B1(n14557), .B2(n14555), .C1(
        n14554), .C2(n14553), .ZN(SUB_1596_U65) );
  OAI21_X1 U16313 ( .B1(n14560), .B2(n14559), .A(n14558), .ZN(n14561) );
  XNOR2_X1 U16314 ( .A(n14561), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  NAND2_X1 U16315 ( .A1(n14562), .A2(n14740), .ZN(n14689) );
  INV_X1 U16316 ( .A(n14689), .ZN(n14563) );
  AOI22_X1 U16317 ( .A1(n14564), .A2(n14563), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14571) );
  AOI211_X1 U16318 ( .C1(n14567), .C2(n14566), .A(n14565), .B(n6606), .ZN(
        n14568) );
  AOI21_X1 U16319 ( .B1(n14584), .B2(n14569), .A(n14568), .ZN(n14570) );
  OAI211_X1 U16320 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n14572), .A(n14571), .B(
        n14570), .ZN(P1_U3218) );
  XNOR2_X1 U16321 ( .A(n14573), .B(n14574), .ZN(n14581) );
  NOR3_X1 U16322 ( .A1(n14576), .A2(n14627), .A3(n14575), .ZN(n14579) );
  NOR2_X1 U16323 ( .A1(n14577), .A2(n14676), .ZN(n14578) );
  AOI211_X1 U16324 ( .C1(n14581), .C2(n14580), .A(n14579), .B(n14578), .ZN(
        n14587) );
  INV_X1 U16325 ( .A(n14582), .ZN(n14585) );
  NOR2_X1 U16326 ( .A1(n8827), .A2(n14583), .ZN(n14633) );
  AOI22_X1 U16327 ( .A1(n14585), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n14584), 
        .B2(n14633), .ZN(n14586) );
  NAND2_X1 U16328 ( .A1(n14587), .A2(n14586), .ZN(P1_U3222) );
  OAI21_X1 U16329 ( .B1(n14590), .B2(n14589), .A(n14588), .ZN(n14592) );
  NAND2_X1 U16330 ( .A1(n14592), .A2(n14591), .ZN(n14599) );
  AOI21_X1 U16331 ( .B1(n14595), .B2(n14594), .A(n14593), .ZN(n14597) );
  OR2_X1 U16332 ( .A1(n14597), .A2(n14596), .ZN(n14598) );
  OAI211_X1 U16333 ( .C1(n14601), .C2(n14600), .A(n14599), .B(n14598), .ZN(
        n14602) );
  INV_X1 U16334 ( .A(n14602), .ZN(n14604) );
  OAI211_X1 U16335 ( .C1(n14606), .C2(n14605), .A(n14604), .B(n14603), .ZN(
        P1_U3255) );
  INV_X1 U16336 ( .A(n14607), .ZN(n14615) );
  OAI22_X1 U16337 ( .A1(n14610), .A2(n10047), .B1(n14609), .B2(n14608), .ZN(
        n14611) );
  AOI21_X1 U16338 ( .B1(n14613), .B2(n14612), .A(n14611), .ZN(n14614) );
  OAI21_X1 U16339 ( .B1(n14615), .B2(n14639), .A(n14614), .ZN(n14616) );
  AOI21_X1 U16340 ( .B1(n14618), .B2(n14617), .A(n14616), .ZN(n14619) );
  OAI21_X1 U16341 ( .B1(n14646), .B2(n14620), .A(n14619), .ZN(P1_U3287) );
  OAI21_X1 U16342 ( .B1(n14627), .B2(n14622), .A(n14621), .ZN(n14635) );
  NAND2_X1 U16343 ( .A1(n10686), .A2(n14622), .ZN(n14629) );
  AND2_X1 U16344 ( .A1(n14623), .A2(n10689), .ZN(n14624) );
  NOR2_X1 U16345 ( .A1(n14625), .A2(n14624), .ZN(n14638) );
  XNOR2_X1 U16346 ( .A(n14638), .B(n14626), .ZN(n14628) );
  MUX2_X1 U16347 ( .A(n14629), .B(n14628), .S(n14627), .Z(n14634) );
  XNOR2_X1 U16348 ( .A(n10686), .B(n14630), .ZN(n14674) );
  NOR2_X1 U16349 ( .A1(n14674), .A2(n14631), .ZN(n14632) );
  AOI211_X1 U16350 ( .C1(n14635), .C2(n14634), .A(n14633), .B(n14632), .ZN(
        n14677) );
  AOI22_X1 U16351 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(n14636), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(n14646), .ZN(n14645) );
  NAND2_X1 U16352 ( .A1(n14638), .A2(n14637), .ZN(n14675) );
  OAI22_X1 U16353 ( .A1(n14640), .A2(n14676), .B1(n14675), .B2(n14639), .ZN(
        n14643) );
  NOR2_X1 U16354 ( .A1(n14641), .A2(n14674), .ZN(n14642) );
  NOR2_X1 U16355 ( .A1(n14643), .A2(n14642), .ZN(n14644) );
  OAI211_X1 U16356 ( .C1(n14646), .C2(n14677), .A(n14645), .B(n14644), .ZN(
        P1_U3292) );
  INV_X1 U16357 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n14647) );
  NOR2_X1 U16358 ( .A1(n14673), .A2(n14647), .ZN(P1_U3294) );
  INV_X1 U16359 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n15260) );
  NOR2_X1 U16360 ( .A1(n14673), .A2(n15260), .ZN(P1_U3295) );
  INV_X1 U16361 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n15169) );
  NOR2_X1 U16362 ( .A1(n14673), .A2(n15169), .ZN(P1_U3296) );
  INV_X1 U16363 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n14648) );
  NOR2_X1 U16364 ( .A1(n14660), .A2(n14648), .ZN(P1_U3297) );
  INV_X1 U16365 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n14649) );
  NOR2_X1 U16366 ( .A1(n14660), .A2(n14649), .ZN(P1_U3298) );
  INV_X1 U16367 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n14650) );
  NOR2_X1 U16368 ( .A1(n14660), .A2(n14650), .ZN(P1_U3299) );
  INV_X1 U16369 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n14651) );
  NOR2_X1 U16370 ( .A1(n14660), .A2(n14651), .ZN(P1_U3300) );
  INV_X1 U16371 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n14652) );
  NOR2_X1 U16372 ( .A1(n14660), .A2(n14652), .ZN(P1_U3301) );
  INV_X1 U16373 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n14653) );
  NOR2_X1 U16374 ( .A1(n14660), .A2(n14653), .ZN(P1_U3302) );
  INV_X1 U16375 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n14654) );
  NOR2_X1 U16376 ( .A1(n14660), .A2(n14654), .ZN(P1_U3303) );
  INV_X1 U16377 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n14655) );
  NOR2_X1 U16378 ( .A1(n14660), .A2(n14655), .ZN(P1_U3304) );
  INV_X1 U16379 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n14656) );
  NOR2_X1 U16380 ( .A1(n14660), .A2(n14656), .ZN(P1_U3305) );
  INV_X1 U16381 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n14657) );
  NOR2_X1 U16382 ( .A1(n14660), .A2(n14657), .ZN(P1_U3306) );
  INV_X1 U16383 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n14658) );
  NOR2_X1 U16384 ( .A1(n14660), .A2(n14658), .ZN(P1_U3307) );
  INV_X1 U16385 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n14659) );
  NOR2_X1 U16386 ( .A1(n14660), .A2(n14659), .ZN(P1_U3308) );
  INV_X1 U16387 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n14661) );
  NOR2_X1 U16388 ( .A1(n14673), .A2(n14661), .ZN(P1_U3309) );
  INV_X1 U16389 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15247) );
  NOR2_X1 U16390 ( .A1(n14673), .A2(n15247), .ZN(P1_U3310) );
  INV_X1 U16391 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n14662) );
  NOR2_X1 U16392 ( .A1(n14673), .A2(n14662), .ZN(P1_U3311) );
  INV_X1 U16393 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n14663) );
  NOR2_X1 U16394 ( .A1(n14673), .A2(n14663), .ZN(P1_U3312) );
  INV_X1 U16395 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n14664) );
  NOR2_X1 U16396 ( .A1(n14673), .A2(n14664), .ZN(P1_U3313) );
  INV_X1 U16397 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n15241) );
  NOR2_X1 U16398 ( .A1(n14673), .A2(n15241), .ZN(P1_U3314) );
  INV_X1 U16399 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n14665) );
  NOR2_X1 U16400 ( .A1(n14673), .A2(n14665), .ZN(P1_U3315) );
  INV_X1 U16401 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n14666) );
  NOR2_X1 U16402 ( .A1(n14673), .A2(n14666), .ZN(P1_U3316) );
  INV_X1 U16403 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n14667) );
  NOR2_X1 U16404 ( .A1(n14673), .A2(n14667), .ZN(P1_U3317) );
  INV_X1 U16405 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n14668) );
  NOR2_X1 U16406 ( .A1(n14673), .A2(n14668), .ZN(P1_U3318) );
  INV_X1 U16407 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n14669) );
  NOR2_X1 U16408 ( .A1(n14673), .A2(n14669), .ZN(P1_U3319) );
  INV_X1 U16409 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n14670) );
  NOR2_X1 U16410 ( .A1(n14673), .A2(n14670), .ZN(P1_U3320) );
  INV_X1 U16411 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n14671) );
  NOR2_X1 U16412 ( .A1(n14673), .A2(n14671), .ZN(P1_U3321) );
  INV_X1 U16413 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n14672) );
  NOR2_X1 U16414 ( .A1(n14673), .A2(n14672), .ZN(P1_U3322) );
  INV_X1 U16415 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15246) );
  NOR2_X1 U16416 ( .A1(n14673), .A2(n15246), .ZN(P1_U3323) );
  INV_X1 U16417 ( .A(n14674), .ZN(n14680) );
  OAI21_X1 U16418 ( .B1(n14676), .B2(n14711), .A(n14675), .ZN(n14679) );
  INV_X1 U16419 ( .A(n14677), .ZN(n14678) );
  AOI211_X1 U16420 ( .C1(n14687), .C2(n14680), .A(n14679), .B(n14678), .ZN(
        n14730) );
  INV_X1 U16421 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14681) );
  AOI22_X1 U16422 ( .A1(n15160), .A2(n14730), .B1(n14681), .B2(n15158), .ZN(
        P1_U3462) );
  INV_X1 U16423 ( .A(n14682), .ZN(n14686) );
  OAI21_X1 U16424 ( .B1(n7038), .B2(n14711), .A(n14683), .ZN(n14685) );
  AOI211_X1 U16425 ( .C1(n14687), .C2(n14686), .A(n14685), .B(n14684), .ZN(
        n14731) );
  AOI22_X1 U16426 ( .A1(n15160), .A2(n14731), .B1(n8354), .B2(n15158), .ZN(
        P1_U3465) );
  INV_X1 U16427 ( .A(n14688), .ZN(n14694) );
  NAND4_X1 U16428 ( .A1(n14692), .A2(n14691), .A3(n14690), .A4(n14689), .ZN(
        n14693) );
  AOI21_X1 U16429 ( .B1(n14694), .B2(n14729), .A(n14693), .ZN(n14732) );
  INV_X1 U16430 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14695) );
  AOI22_X1 U16431 ( .A1(n15160), .A2(n14732), .B1(n14695), .B2(n15158), .ZN(
        P1_U3468) );
  OR4_X1 U16432 ( .A1(n14699), .A2(n14698), .A3(n14697), .A4(n14696), .ZN(
        n14700) );
  AOI21_X1 U16433 ( .B1(n14701), .B2(n14729), .A(n14700), .ZN(n14733) );
  INV_X1 U16434 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14702) );
  AOI22_X1 U16435 ( .A1(n15160), .A2(n14733), .B1(n14702), .B2(n15158), .ZN(
        P1_U3471) );
  INV_X1 U16436 ( .A(n14703), .ZN(n14709) );
  OR3_X1 U16437 ( .A1(n14706), .A2(n14705), .A3(n14704), .ZN(n14707) );
  AOI211_X1 U16438 ( .C1(n14709), .C2(n14729), .A(n14708), .B(n14707), .ZN(
        n14735) );
  AOI22_X1 U16439 ( .A1(n15160), .A2(n14735), .B1(n8403), .B2(n15158), .ZN(
        P1_U3474) );
  OAI21_X1 U16440 ( .B1(n14712), .B2(n14711), .A(n14710), .ZN(n14714) );
  AOI211_X1 U16441 ( .C1(n14729), .C2(n14715), .A(n14714), .B(n14713), .ZN(
        n14736) );
  INV_X1 U16442 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14716) );
  AOI22_X1 U16443 ( .A1(n15160), .A2(n14736), .B1(n14716), .B2(n15158), .ZN(
        P1_U3480) );
  AOI22_X1 U16444 ( .A1(n14718), .A2(n14729), .B1(n14740), .B2(n14717), .ZN(
        n14720) );
  NAND2_X1 U16445 ( .A1(n14720), .A2(n14719), .ZN(n14721) );
  NOR2_X1 U16446 ( .A1(n14722), .A2(n14721), .ZN(n14737) );
  INV_X1 U16447 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14723) );
  AOI22_X1 U16448 ( .A1(n15160), .A2(n14737), .B1(n14723), .B2(n15158), .ZN(
        P1_U3483) );
  NAND3_X1 U16449 ( .A1(n14726), .A2(n14725), .A3(n14724), .ZN(n14727) );
  AOI21_X1 U16450 ( .B1(n14729), .B2(n14728), .A(n14727), .ZN(n14747) );
  AOI22_X1 U16451 ( .A1(n15160), .A2(n14747), .B1(n8487), .B2(n15158), .ZN(
        P1_U3489) );
  AOI22_X1 U16452 ( .A1(n14748), .A2(n14730), .B1(n15162), .B2(n14746), .ZN(
        P1_U3529) );
  AOI22_X1 U16453 ( .A1(n14748), .A2(n14731), .B1(n10007), .B2(n14746), .ZN(
        P1_U3530) );
  AOI22_X1 U16454 ( .A1(n14748), .A2(n14732), .B1(n10008), .B2(n14746), .ZN(
        P1_U3531) );
  AOI22_X1 U16455 ( .A1(n14748), .A2(n14733), .B1(n15244), .B2(n14746), .ZN(
        P1_U3532) );
  INV_X1 U16456 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n14734) );
  AOI22_X1 U16457 ( .A1(n14748), .A2(n14735), .B1(n14734), .B2(n14746), .ZN(
        P1_U3533) );
  AOI22_X1 U16458 ( .A1(n14748), .A2(n14736), .B1(n10057), .B2(n14746), .ZN(
        P1_U3535) );
  AOI22_X1 U16459 ( .A1(n14748), .A2(n14737), .B1(n10058), .B2(n14746), .ZN(
        P1_U3536) );
  AOI21_X1 U16460 ( .B1(n14740), .B2(n14739), .A(n14738), .ZN(n14741) );
  OAI211_X1 U16461 ( .C1(n14744), .C2(n14743), .A(n14742), .B(n14741), .ZN(
        n15159) );
  OAI22_X1 U16462 ( .A1(n14746), .A2(n15159), .B1(P1_REG1_REG_9__SCAN_IN), 
        .B2(n14748), .ZN(n14745) );
  INV_X1 U16463 ( .A(n14745), .ZN(P1_U3537) );
  AOI22_X1 U16464 ( .A1(n14748), .A2(n14747), .B1(n10205), .B2(n14746), .ZN(
        P1_U3538) );
  NOR2_X1 U16465 ( .A1(n14812), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI21_X1 U16466 ( .B1(n14820), .B2(P2_REG2_REG_0__SCAN_IN), .A(n14749), .ZN(
        n14755) );
  AOI22_X1 U16467 ( .A1(n14812), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14754) );
  OAI22_X1 U16468 ( .A1(n14751), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n14750), .ZN(n14752) );
  OAI21_X1 U16469 ( .B1(n14818), .B2(n14752), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n14753) );
  OAI211_X1 U16470 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n14755), .A(n14754), .B(
        n14753), .ZN(P2_U3214) );
  NAND2_X1 U16471 ( .A1(n14757), .A2(n14756), .ZN(n14758) );
  NAND2_X1 U16472 ( .A1(n14759), .A2(n14758), .ZN(n14760) );
  NAND2_X1 U16473 ( .A1(n14814), .A2(n14760), .ZN(n14767) );
  NAND2_X1 U16474 ( .A1(n14762), .A2(n14761), .ZN(n14763) );
  NAND2_X1 U16475 ( .A1(n14764), .A2(n14763), .ZN(n14765) );
  NAND2_X1 U16476 ( .A1(n14820), .A2(n14765), .ZN(n14766) );
  OAI211_X1 U16477 ( .C1(n14769), .C2(n14768), .A(n14767), .B(n14766), .ZN(
        n14770) );
  INV_X1 U16478 ( .A(n14770), .ZN(n14772) );
  OAI211_X1 U16479 ( .C1(n14773), .C2(n14791), .A(n14772), .B(n14771), .ZN(
        P2_U3223) );
  AND2_X1 U16480 ( .A1(n14775), .A2(n14774), .ZN(n14778) );
  OAI21_X1 U16481 ( .B1(n14778), .B2(n14777), .A(n14776), .ZN(n14788) );
  INV_X1 U16482 ( .A(n14779), .ZN(n14787) );
  INV_X1 U16483 ( .A(n14780), .ZN(n14785) );
  NAND3_X1 U16484 ( .A1(n14783), .A2(n14782), .A3(n14781), .ZN(n14784) );
  NAND2_X1 U16485 ( .A1(n14785), .A2(n14784), .ZN(n14786) );
  AOI222_X1 U16486 ( .A1(n14788), .A2(n14814), .B1(n14787), .B2(n14818), .C1(
        n14786), .C2(n14820), .ZN(n14790) );
  NAND2_X1 U16487 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14789)
         );
  OAI211_X1 U16488 ( .C1(n14792), .C2(n14791), .A(n14790), .B(n14789), .ZN(
        P2_U3226) );
  AOI22_X1 U16489 ( .A1(n14812), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3088), .ZN(n14802) );
  NAND2_X1 U16490 ( .A1(n14818), .A2(n14793), .ZN(n14801) );
  OAI211_X1 U16491 ( .C1(n14795), .C2(P2_REG2_REG_14__SCAN_IN), .A(n14794), 
        .B(n14820), .ZN(n14800) );
  OAI211_X1 U16492 ( .C1(n14798), .C2(n14797), .A(n14796), .B(n14814), .ZN(
        n14799) );
  NAND4_X1 U16493 ( .A1(n14802), .A2(n14801), .A3(n14800), .A4(n14799), .ZN(
        P2_U3228) );
  AOI22_X1 U16494 ( .A1(n14812), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14811) );
  OAI211_X1 U16495 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n14804), .A(n14820), 
        .B(n14803), .ZN(n14810) );
  NAND2_X1 U16496 ( .A1(n14818), .A2(n14805), .ZN(n14809) );
  OAI211_X1 U16497 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n14807), .A(n14814), 
        .B(n14806), .ZN(n14808) );
  NAND4_X1 U16498 ( .A1(n14811), .A2(n14810), .A3(n14809), .A4(n14808), .ZN(
        P2_U3229) );
  AOI22_X1 U16499 ( .A1(n14812), .A2(P2_ADDR_REG_17__SCAN_IN), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3088), .ZN(n14826) );
  OAI211_X1 U16500 ( .C1(n14816), .C2(n14815), .A(n14814), .B(n14813), .ZN(
        n14825) );
  NAND2_X1 U16501 ( .A1(n14818), .A2(n14817), .ZN(n14824) );
  OAI211_X1 U16502 ( .C1(n14822), .C2(n14821), .A(n14820), .B(n14819), .ZN(
        n14823) );
  NAND4_X1 U16503 ( .A1(n14826), .A2(n14825), .A3(n14824), .A4(n14823), .ZN(
        P2_U3231) );
  INV_X1 U16504 ( .A(n14835), .ZN(n14832) );
  INV_X1 U16505 ( .A(n14828), .ZN(n14829) );
  AND2_X1 U16506 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14829), .ZN(P2_U3266) );
  AND2_X1 U16507 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14829), .ZN(P2_U3267) );
  AND2_X1 U16508 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14829), .ZN(P2_U3268) );
  AND2_X1 U16509 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14829), .ZN(P2_U3269) );
  AND2_X1 U16510 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14829), .ZN(P2_U3270) );
  AND2_X1 U16511 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14829), .ZN(P2_U3271) );
  AND2_X1 U16512 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14829), .ZN(P2_U3272) );
  AND2_X1 U16513 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14829), .ZN(P2_U3273) );
  AND2_X1 U16514 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14829), .ZN(P2_U3274) );
  AND2_X1 U16515 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14829), .ZN(P2_U3275) );
  AND2_X1 U16516 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14829), .ZN(P2_U3276) );
  AND2_X1 U16517 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14829), .ZN(P2_U3277) );
  AND2_X1 U16518 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14829), .ZN(P2_U3278) );
  AND2_X1 U16519 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14829), .ZN(P2_U3279) );
  AND2_X1 U16520 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14829), .ZN(P2_U3280) );
  AND2_X1 U16521 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14829), .ZN(P2_U3281) );
  AND2_X1 U16522 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14829), .ZN(P2_U3282) );
  AND2_X1 U16523 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14829), .ZN(P2_U3283) );
  INV_X1 U16524 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n15163) );
  NOR2_X1 U16525 ( .A1(n14828), .A2(n15163), .ZN(P2_U3284) );
  AND2_X1 U16526 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14829), .ZN(P2_U3285) );
  INV_X1 U16527 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n15175) );
  NOR2_X1 U16528 ( .A1(n14828), .A2(n15175), .ZN(P2_U3286) );
  AND2_X1 U16529 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14829), .ZN(P2_U3287) );
  AND2_X1 U16530 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14829), .ZN(P2_U3288) );
  AND2_X1 U16531 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14829), .ZN(P2_U3289) );
  AND2_X1 U16532 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14829), .ZN(P2_U3290) );
  AND2_X1 U16533 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14829), .ZN(P2_U3291) );
  AND2_X1 U16534 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14829), .ZN(P2_U3292) );
  INV_X1 U16535 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n15235) );
  NOR2_X1 U16536 ( .A1(n14828), .A2(n15235), .ZN(P2_U3293) );
  AND2_X1 U16537 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14829), .ZN(P2_U3294) );
  AND2_X1 U16538 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14829), .ZN(P2_U3295) );
  AOI22_X1 U16539 ( .A1(n14835), .A2(n14831), .B1(n14830), .B2(n14832), .ZN(
        P2_U3416) );
  AOI22_X1 U16540 ( .A1(n14835), .A2(n14834), .B1(n14833), .B2(n14832), .ZN(
        P2_U3417) );
  AOI21_X1 U16541 ( .B1(n14845), .B2(n14837), .A(n14836), .ZN(n14839) );
  OAI211_X1 U16542 ( .C1(n14841), .C2(n14840), .A(n14839), .B(n14838), .ZN(
        n14842) );
  INV_X1 U16543 ( .A(n14842), .ZN(n14860) );
  AOI22_X1 U16544 ( .A1(n14859), .A2(n14860), .B1(n7738), .B2(n14858), .ZN(
        P2_U3436) );
  AOI21_X1 U16545 ( .B1(n14845), .B2(n14844), .A(n14843), .ZN(n14846) );
  OAI211_X1 U16546 ( .C1(n14848), .C2(n11860), .A(n14847), .B(n14846), .ZN(
        n14849) );
  INV_X1 U16547 ( .A(n14849), .ZN(n14861) );
  AOI22_X1 U16548 ( .A1(n14859), .A2(n14861), .B1(n7772), .B2(n14858), .ZN(
        P2_U3442) );
  AND2_X1 U16549 ( .A1(n14851), .A2(n14850), .ZN(n14857) );
  OAI21_X1 U16550 ( .B1(n14854), .B2(n14853), .A(n14852), .ZN(n14855) );
  NOR3_X1 U16551 ( .A1(n14857), .A2(n14856), .A3(n14855), .ZN(n14863) );
  AOI22_X1 U16552 ( .A1(n14859), .A2(n14863), .B1(n7898), .B2(n14858), .ZN(
        P2_U3463) );
  AOI22_X1 U16553 ( .A1(n14864), .A2(n14860), .B1(n9939), .B2(n14862), .ZN(
        P2_U3501) );
  AOI22_X1 U16554 ( .A1(n14864), .A2(n14861), .B1(n9945), .B2(n14862), .ZN(
        P2_U3503) );
  AOI22_X1 U16555 ( .A1(n14864), .A2(n14863), .B1(n10124), .B2(n14862), .ZN(
        P2_U3510) );
  NOR2_X1 U16556 ( .A1(P3_U3897), .A2(n15030), .ZN(P3_U3150) );
  NOR3_X1 U16557 ( .A1(n15035), .A2(n14866), .A3(n15037), .ZN(n14876) );
  AOI22_X1 U16558 ( .A1(n15035), .A2(n14867), .B1(n14866), .B2(n14865), .ZN(
        n14874) );
  NAND2_X1 U16559 ( .A1(n15037), .A2(n14868), .ZN(n14869) );
  AOI22_X1 U16560 ( .A1(n15030), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n14871) );
  AND2_X1 U16561 ( .A1(n14872), .A2(n14871), .ZN(n14873) );
  OAI211_X1 U16562 ( .C1(n14876), .C2(n14875), .A(n14874), .B(n14873), .ZN(
        P3_U3182) );
  OR2_X1 U16563 ( .A1(n14877), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n14878) );
  AND2_X1 U16564 ( .A1(n14879), .A2(n14878), .ZN(n14894) );
  AND3_X1 U16565 ( .A1(n14882), .A2(n14881), .A3(n14880), .ZN(n14883) );
  OAI21_X1 U16566 ( .B1(n14884), .B2(n14883), .A(n15037), .ZN(n14887) );
  INV_X1 U16567 ( .A(n14885), .ZN(n14886) );
  OAI211_X1 U16568 ( .C1(n14996), .C2(n14214), .A(n14887), .B(n14886), .ZN(
        n14888) );
  AOI21_X1 U16569 ( .B1(n14889), .B2(n14992), .A(n14888), .ZN(n14893) );
  XNOR2_X1 U16570 ( .A(n14890), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n14891) );
  NAND2_X1 U16571 ( .A1(n15035), .A2(n14891), .ZN(n14892) );
  OAI211_X1 U16572 ( .C1(n14894), .C2(n15043), .A(n14893), .B(n14892), .ZN(
        P3_U3185) );
  NOR2_X1 U16573 ( .A1(n14896), .A2(n14895), .ZN(n14897) );
  NOR2_X1 U16574 ( .A1(n14898), .A2(n14897), .ZN(n14915) );
  INV_X1 U16575 ( .A(n14899), .ZN(n14900) );
  OAI21_X1 U16576 ( .B1(n14996), .B2(n14216), .A(n14900), .ZN(n14906) );
  AOI21_X1 U16577 ( .B1(n14903), .B2(n14902), .A(n14901), .ZN(n14904) );
  NOR2_X1 U16578 ( .A1(n14904), .A2(n15018), .ZN(n14905) );
  AOI211_X1 U16579 ( .C1(n14992), .C2(n14907), .A(n14906), .B(n14905), .ZN(
        n14914) );
  AOI21_X1 U16580 ( .B1(n14910), .B2(n14909), .A(n14908), .ZN(n14911) );
  OR2_X1 U16581 ( .A1(n14912), .A2(n14911), .ZN(n14913) );
  OAI211_X1 U16582 ( .C1(n14915), .C2(n15043), .A(n14914), .B(n14913), .ZN(
        P3_U3186) );
  AOI21_X1 U16583 ( .B1(n14918), .B2(n14917), .A(n14916), .ZN(n14931) );
  NOR2_X1 U16584 ( .A1(n14920), .A2(n14919), .ZN(n14921) );
  XNOR2_X1 U16585 ( .A(n6601), .B(n14921), .ZN(n14923) );
  OAI22_X1 U16586 ( .A1(n14923), .A2(n15018), .B1(n14922), .B2(n15033), .ZN(
        n14924) );
  AOI211_X1 U16587 ( .C1(P3_ADDR_REG_5__SCAN_IN), .C2(n15030), .A(n14925), .B(
        n14924), .ZN(n14930) );
  OAI21_X1 U16588 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n14927), .A(n14926), .ZN(
        n14928) );
  NAND2_X1 U16589 ( .A1(n15035), .A2(n14928), .ZN(n14929) );
  OAI211_X1 U16590 ( .C1(n14931), .C2(n15043), .A(n14930), .B(n14929), .ZN(
        P3_U3187) );
  AOI21_X1 U16591 ( .B1(n14934), .B2(n14933), .A(n14932), .ZN(n14949) );
  INV_X1 U16592 ( .A(n14935), .ZN(n14937) );
  NAND2_X1 U16593 ( .A1(n14937), .A2(n14936), .ZN(n14938) );
  XNOR2_X1 U16594 ( .A(n14939), .B(n14938), .ZN(n14941) );
  OAI22_X1 U16595 ( .A1(n14941), .A2(n15018), .B1(n14940), .B2(n15033), .ZN(
        n14942) );
  AOI211_X1 U16596 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15030), .A(n14943), .B(
        n14942), .ZN(n14948) );
  OAI21_X1 U16597 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n14945), .A(n14944), .ZN(
        n14946) );
  NAND2_X1 U16598 ( .A1(n14946), .A2(n15035), .ZN(n14947) );
  OAI211_X1 U16599 ( .C1(n14949), .C2(n15043), .A(n14948), .B(n14947), .ZN(
        P3_U3191) );
  OAI21_X1 U16600 ( .B1(n14952), .B2(n14951), .A(n14950), .ZN(n14954) );
  AOI21_X1 U16601 ( .B1(n14954), .B2(n15035), .A(n14953), .ZN(n14966) );
  AOI21_X1 U16602 ( .B1(n14957), .B2(n14956), .A(n14955), .ZN(n14962) );
  AOI21_X1 U16603 ( .B1(n14960), .B2(n14959), .A(n14958), .ZN(n14961) );
  OAI222_X1 U16604 ( .A1(n15033), .A2(n14963), .B1(n15018), .B2(n14962), .C1(
        n15043), .C2(n14961), .ZN(n14964) );
  INV_X1 U16605 ( .A(n14964), .ZN(n14965) );
  OAI211_X1 U16606 ( .C1(n14996), .C2(n14967), .A(n14966), .B(n14965), .ZN(
        P3_U3192) );
  AOI21_X1 U16607 ( .B1(n14970), .B2(n14969), .A(n14968), .ZN(n14984) );
  OAI21_X1 U16608 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n14972), .A(n14971), 
        .ZN(n14977) );
  AOI21_X1 U16609 ( .B1(n15030), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n14973), 
        .ZN(n14974) );
  OAI21_X1 U16610 ( .B1(n15033), .B2(n14975), .A(n14974), .ZN(n14976) );
  AOI21_X1 U16611 ( .B1(n14977), .B2(n15035), .A(n14976), .ZN(n14983) );
  NOR2_X1 U16612 ( .A1(n14979), .A2(n14978), .ZN(n14980) );
  OAI21_X1 U16613 ( .B1(n14981), .B2(n14980), .A(n15037), .ZN(n14982) );
  OAI211_X1 U16614 ( .C1(n14984), .C2(n15043), .A(n14983), .B(n14982), .ZN(
        P3_U3193) );
  AOI21_X1 U16615 ( .B1(n14987), .B2(n14986), .A(n14985), .ZN(n15005) );
  OAI21_X1 U16616 ( .B1(n14990), .B2(n14989), .A(n14988), .ZN(n14999) );
  INV_X1 U16617 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14997) );
  NAND2_X1 U16618 ( .A1(n14992), .A2(n14991), .ZN(n14995) );
  INV_X1 U16619 ( .A(n14993), .ZN(n14994) );
  OAI211_X1 U16620 ( .C1(n14997), .C2(n14996), .A(n14995), .B(n14994), .ZN(
        n14998) );
  AOI21_X1 U16621 ( .B1(n14999), .B2(n15035), .A(n14998), .ZN(n15004) );
  OAI211_X1 U16622 ( .C1(n15002), .C2(n15001), .A(n15037), .B(n15000), .ZN(
        n15003) );
  OAI211_X1 U16623 ( .C1(n15005), .C2(n15043), .A(n15004), .B(n15003), .ZN(
        P3_U3194) );
  AOI21_X1 U16624 ( .B1(n15242), .B2(n15007), .A(n15006), .ZN(n15022) );
  OAI21_X1 U16625 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n15009), .A(n15008), 
        .ZN(n15014) );
  AOI21_X1 U16626 ( .B1(n15030), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n15010), 
        .ZN(n15011) );
  OAI21_X1 U16627 ( .B1(n15033), .B2(n15012), .A(n15011), .ZN(n15013) );
  AOI21_X1 U16628 ( .B1(n15014), .B2(n15035), .A(n15013), .ZN(n15021) );
  AOI21_X1 U16629 ( .B1(n15017), .B2(n15016), .A(n15015), .ZN(n15019) );
  OR2_X1 U16630 ( .A1(n15019), .A2(n15018), .ZN(n15020) );
  OAI211_X1 U16631 ( .C1(n15022), .C2(n15043), .A(n15021), .B(n15020), .ZN(
        P3_U3195) );
  AOI21_X1 U16632 ( .B1(n15025), .B2(n15024), .A(n15023), .ZN(n15044) );
  OAI21_X1 U16633 ( .B1(n15028), .B2(n15027), .A(n15026), .ZN(n15036) );
  AOI21_X1 U16634 ( .B1(n15030), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n15029), 
        .ZN(n15031) );
  OAI21_X1 U16635 ( .B1(n15033), .B2(n15032), .A(n15031), .ZN(n15034) );
  AOI21_X1 U16636 ( .B1(n15036), .B2(n15035), .A(n15034), .ZN(n15042) );
  OAI211_X1 U16637 ( .C1(n15040), .C2(n15039), .A(n15038), .B(n15037), .ZN(
        n15041) );
  OAI211_X1 U16638 ( .C1(n15044), .C2(n15043), .A(n15042), .B(n15041), .ZN(
        P3_U3196) );
  XNOR2_X1 U16639 ( .A(n15045), .B(n15051), .ZN(n15124) );
  OAI22_X1 U16640 ( .A1(n15087), .A2(n15046), .B1(n15061), .B2(n15084), .ZN(
        n15053) );
  INV_X1 U16641 ( .A(n15047), .ZN(n15048) );
  AOI211_X1 U16642 ( .C1(n15051), .C2(n15050), .A(n15049), .B(n15048), .ZN(
        n15052) );
  AOI211_X1 U16643 ( .C1(n15124), .C2(n15054), .A(n15053), .B(n15052), .ZN(
        n15121) );
  AOI22_X1 U16644 ( .A1(n15071), .A2(n15055), .B1(n15075), .B2(
        P3_REG2_REG_6__SCAN_IN), .ZN(n15059) );
  NOR2_X1 U16645 ( .A1(n15056), .A2(n15136), .ZN(n15123) );
  AOI22_X1 U16646 ( .A1(n15124), .A2(n15057), .B1(n15072), .B2(n15123), .ZN(
        n15058) );
  OAI211_X1 U16647 ( .C1(n15075), .C2(n15121), .A(n15059), .B(n15058), .ZN(
        P3_U3227) );
  XNOR2_X1 U16648 ( .A(n15060), .B(n15064), .ZN(n15068) );
  INV_X1 U16649 ( .A(n15068), .ZN(n15115) );
  OAI22_X1 U16650 ( .A1(n15087), .A2(n15061), .B1(n15086), .B2(n15084), .ZN(
        n15062) );
  INV_X1 U16651 ( .A(n15062), .ZN(n15067) );
  OAI211_X1 U16652 ( .C1(n15065), .C2(n15064), .A(n15063), .B(n15089), .ZN(
        n15066) );
  OAI211_X1 U16653 ( .C1(n15068), .C2(n15093), .A(n15067), .B(n15066), .ZN(
        n15113) );
  AOI21_X1 U16654 ( .B1(n15095), .B2(n15115), .A(n15113), .ZN(n15074) );
  INV_X1 U16655 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n15300) );
  AND2_X1 U16656 ( .A1(n15078), .A2(n15069), .ZN(n15114) );
  AOI22_X1 U16657 ( .A1(n15072), .A2(n15114), .B1(n15071), .B2(n15070), .ZN(
        n15073) );
  OAI221_X1 U16658 ( .B1(n15075), .B2(n15074), .C1(n15096), .C2(n15300), .A(
        n15073), .ZN(P3_U3229) );
  XNOR2_X1 U16659 ( .A(n15082), .B(n15076), .ZN(n15092) );
  INV_X1 U16660 ( .A(n15092), .ZN(n15105) );
  AND2_X1 U16661 ( .A1(n15078), .A2(n15077), .ZN(n15104) );
  NAND2_X1 U16662 ( .A1(n15104), .A2(n15079), .ZN(n15080) );
  OAI21_X1 U16663 ( .B1(n15081), .B2(n15258), .A(n15080), .ZN(n15094) );
  XNOR2_X1 U16664 ( .A(n15083), .B(n15082), .ZN(n15090) );
  OAI22_X1 U16665 ( .A1(n15087), .A2(n15086), .B1(n15085), .B2(n15084), .ZN(
        n15088) );
  AOI21_X1 U16666 ( .B1(n15090), .B2(n15089), .A(n15088), .ZN(n15091) );
  OAI21_X1 U16667 ( .B1(n15093), .B2(n15092), .A(n15091), .ZN(n15103) );
  AOI211_X1 U16668 ( .C1(n15095), .C2(n15105), .A(n15094), .B(n15103), .ZN(
        n15097) );
  AOI22_X1 U16669 ( .A1(n15075), .A2(n10457), .B1(n15097), .B2(n15096), .ZN(
        P3_U3231) );
  INV_X1 U16670 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15102) );
  AOI211_X1 U16671 ( .C1(n15101), .C2(n15100), .A(n15099), .B(n15098), .ZN(
        n15143) );
  AOI22_X1 U16672 ( .A1(n15142), .A2(n15102), .B1(n15143), .B2(n15141), .ZN(
        P3_U3393) );
  INV_X1 U16673 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15106) );
  AOI211_X1 U16674 ( .C1(n15105), .C2(n15133), .A(n15104), .B(n15103), .ZN(
        n15144) );
  AOI22_X1 U16675 ( .A1(n15142), .A2(n15106), .B1(n15144), .B2(n15141), .ZN(
        P3_U3396) );
  INV_X1 U16676 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15112) );
  INV_X1 U16677 ( .A(n15107), .ZN(n15111) );
  NOR2_X1 U16678 ( .A1(n15108), .A2(n15136), .ZN(n15110) );
  AOI211_X1 U16679 ( .C1(n15111), .C2(n15133), .A(n15110), .B(n15109), .ZN(
        n15145) );
  AOI22_X1 U16680 ( .A1(n15142), .A2(n15112), .B1(n15145), .B2(n15141), .ZN(
        P3_U3399) );
  INV_X1 U16681 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15116) );
  AOI211_X1 U16682 ( .C1(n15115), .C2(n15133), .A(n15114), .B(n15113), .ZN(
        n15146) );
  AOI22_X1 U16683 ( .A1(n15142), .A2(n15116), .B1(n15146), .B2(n15141), .ZN(
        P3_U3402) );
  INV_X1 U16684 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15120) );
  AOI211_X1 U16685 ( .C1(n15119), .C2(n15133), .A(n15118), .B(n15117), .ZN(
        n15148) );
  AOI22_X1 U16686 ( .A1(n15142), .A2(n15120), .B1(n15148), .B2(n15141), .ZN(
        P3_U3405) );
  INV_X1 U16687 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15125) );
  INV_X1 U16688 ( .A(n15121), .ZN(n15122) );
  AOI211_X1 U16689 ( .C1(n15124), .C2(n15133), .A(n15123), .B(n15122), .ZN(
        n15150) );
  AOI22_X1 U16690 ( .A1(n15142), .A2(n15125), .B1(n15150), .B2(n15141), .ZN(
        P3_U3408) );
  INV_X1 U16691 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15129) );
  AOI211_X1 U16692 ( .C1(n15128), .C2(n15133), .A(n15127), .B(n15126), .ZN(
        n15152) );
  AOI22_X1 U16693 ( .A1(n15142), .A2(n15129), .B1(n15152), .B2(n15141), .ZN(
        P3_U3411) );
  INV_X1 U16694 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15134) );
  AOI211_X1 U16695 ( .C1(n15133), .C2(n15132), .A(n15131), .B(n15130), .ZN(
        n15153) );
  AOI22_X1 U16696 ( .A1(n15142), .A2(n15134), .B1(n15153), .B2(n15141), .ZN(
        P3_U3414) );
  INV_X1 U16697 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15281) );
  OAI22_X1 U16698 ( .A1(n15138), .A2(n15137), .B1(n15136), .B2(n15135), .ZN(
        n15139) );
  NOR2_X1 U16699 ( .A1(n15140), .A2(n15139), .ZN(n15156) );
  AOI22_X1 U16700 ( .A1(n15142), .A2(n15281), .B1(n15156), .B2(n15141), .ZN(
        P3_U3417) );
  AOI22_X1 U16701 ( .A1(n15157), .A2(n15143), .B1(n10408), .B2(n15154), .ZN(
        P3_U3460) );
  AOI22_X1 U16702 ( .A1(n15157), .A2(n15144), .B1(n10456), .B2(n15154), .ZN(
        P3_U3461) );
  AOI22_X1 U16703 ( .A1(n15157), .A2(n15145), .B1(n10462), .B2(n15154), .ZN(
        P3_U3462) );
  AOI22_X1 U16704 ( .A1(n15157), .A2(n15146), .B1(n10435), .B2(n15154), .ZN(
        P3_U3463) );
  INV_X1 U16705 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15147) );
  AOI22_X1 U16706 ( .A1(n15157), .A2(n15148), .B1(n15147), .B2(n15154), .ZN(
        P3_U3464) );
  AOI22_X1 U16707 ( .A1(n15157), .A2(n15150), .B1(n15149), .B2(n15154), .ZN(
        P3_U3465) );
  INV_X1 U16708 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15151) );
  AOI22_X1 U16709 ( .A1(n15157), .A2(n15152), .B1(n15151), .B2(n15154), .ZN(
        P3_U3466) );
  AOI22_X1 U16710 ( .A1(n15157), .A2(n15153), .B1(n10553), .B2(n15154), .ZN(
        P3_U3467) );
  AOI22_X1 U16711 ( .A1(n15157), .A2(n15156), .B1(n15155), .B2(n15154), .ZN(
        P3_U3468) );
  AOI22_X1 U16712 ( .A1(n15160), .A2(n15159), .B1(P1_REG0_REG_9__SCAN_IN), 
        .B2(n15158), .ZN(n15317) );
  AOI22_X1 U16713 ( .A1(n15163), .A2(keyinput60), .B1(n15162), .B2(keyinput10), 
        .ZN(n15161) );
  OAI221_X1 U16714 ( .B1(n15163), .B2(keyinput60), .C1(n15162), .C2(keyinput10), .A(n15161), .ZN(n15173) );
  AOI22_X1 U16715 ( .A1(n15165), .A2(keyinput8), .B1(n15299), .B2(keyinput63), 
        .ZN(n15164) );
  OAI221_X1 U16716 ( .B1(n15165), .B2(keyinput8), .C1(n15299), .C2(keyinput63), 
        .A(n15164), .ZN(n15172) );
  AOI22_X1 U16717 ( .A1(n15300), .A2(keyinput16), .B1(keyinput19), .B2(n15167), 
        .ZN(n15166) );
  OAI221_X1 U16718 ( .B1(n15300), .B2(keyinput16), .C1(n15167), .C2(keyinput19), .A(n15166), .ZN(n15171) );
  AOI22_X1 U16719 ( .A1(n15169), .A2(keyinput37), .B1(keyinput14), .B2(n15301), 
        .ZN(n15168) );
  OAI221_X1 U16720 ( .B1(n15169), .B2(keyinput37), .C1(n15301), .C2(keyinput14), .A(n15168), .ZN(n15170) );
  NOR4_X1 U16721 ( .A1(n15173), .A2(n15172), .A3(n15171), .A4(n15170), .ZN(
        n15214) );
  AOI22_X1 U16722 ( .A1(n15175), .A2(keyinput48), .B1(n15286), .B2(keyinput5), 
        .ZN(n15174) );
  OAI221_X1 U16723 ( .B1(n15175), .B2(keyinput48), .C1(n15286), .C2(keyinput5), 
        .A(n15174), .ZN(n15185) );
  AOI22_X1 U16724 ( .A1(n15178), .A2(keyinput17), .B1(keyinput11), .B2(n15177), 
        .ZN(n15176) );
  OAI221_X1 U16725 ( .B1(n15178), .B2(keyinput17), .C1(n15177), .C2(keyinput11), .A(n15176), .ZN(n15184) );
  INV_X1 U16726 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n15273) );
  AOI22_X1 U16727 ( .A1(n15273), .A2(keyinput47), .B1(n15298), .B2(keyinput4), 
        .ZN(n15179) );
  OAI221_X1 U16728 ( .B1(n15273), .B2(keyinput47), .C1(n15298), .C2(keyinput4), 
        .A(n15179), .ZN(n15183) );
  AOI22_X1 U16729 ( .A1(n15181), .A2(keyinput59), .B1(keyinput15), .B2(n13360), 
        .ZN(n15180) );
  OAI221_X1 U16730 ( .B1(n15181), .B2(keyinput59), .C1(n13360), .C2(keyinput15), .A(n15180), .ZN(n15182) );
  NOR4_X1 U16731 ( .A1(n15185), .A2(n15184), .A3(n15183), .A4(n15182), .ZN(
        n15213) );
  INV_X1 U16732 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n15188) );
  INV_X1 U16733 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n15187) );
  AOI22_X1 U16734 ( .A1(n15188), .A2(keyinput26), .B1(keyinput42), .B2(n15187), 
        .ZN(n15186) );
  OAI221_X1 U16735 ( .B1(n15188), .B2(keyinput26), .C1(n15187), .C2(keyinput42), .A(n15186), .ZN(n15200) );
  AOI22_X1 U16736 ( .A1(n15191), .A2(keyinput31), .B1(n15190), .B2(keyinput25), 
        .ZN(n15189) );
  OAI221_X1 U16737 ( .B1(n15191), .B2(keyinput31), .C1(n15190), .C2(keyinput25), .A(n15189), .ZN(n15199) );
  AOI22_X1 U16738 ( .A1(n15194), .A2(keyinput34), .B1(n15193), .B2(keyinput49), 
        .ZN(n15192) );
  OAI221_X1 U16739 ( .B1(n15194), .B2(keyinput34), .C1(n15193), .C2(keyinput49), .A(n15192), .ZN(n15198) );
  XNOR2_X1 U16740 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput50), .ZN(n15196) );
  XNOR2_X1 U16741 ( .A(P1_REG1_REG_19__SCAN_IN), .B(keyinput56), .ZN(n15195)
         );
  NAND2_X1 U16742 ( .A1(n15196), .A2(n15195), .ZN(n15197) );
  NOR4_X1 U16743 ( .A1(n15200), .A2(n15199), .A3(n15198), .A4(n15197), .ZN(
        n15212) );
  AOI22_X1 U16744 ( .A1(n15304), .A2(keyinput21), .B1(n15289), .B2(keyinput53), 
        .ZN(n15201) );
  OAI221_X1 U16745 ( .B1(n15304), .B2(keyinput21), .C1(n15289), .C2(keyinput53), .A(n15201), .ZN(n15210) );
  AOI22_X1 U16746 ( .A1(n15302), .A2(keyinput58), .B1(n15303), .B2(keyinput40), 
        .ZN(n15202) );
  OAI221_X1 U16747 ( .B1(n15302), .B2(keyinput58), .C1(n15303), .C2(keyinput40), .A(n15202), .ZN(n15209) );
  INV_X1 U16748 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n15203) );
  XOR2_X1 U16749 ( .A(n15203), .B(keyinput20), .Z(n15207) );
  XNOR2_X1 U16750 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput55), .ZN(n15206) );
  XNOR2_X1 U16751 ( .A(P3_REG3_REG_22__SCAN_IN), .B(keyinput1), .ZN(n15205) );
  XNOR2_X1 U16752 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput33), .ZN(n15204) );
  NAND4_X1 U16753 ( .A1(n15207), .A2(n15206), .A3(n15205), .A4(n15204), .ZN(
        n15208) );
  NOR3_X1 U16754 ( .A1(n15210), .A2(n15209), .A3(n15208), .ZN(n15211) );
  NAND4_X1 U16755 ( .A1(n15214), .A2(n15213), .A3(n15212), .A4(n15211), .ZN(
        n15272) );
  AOI22_X1 U16756 ( .A1(n15217), .A2(keyinput24), .B1(keyinput3), .B2(n15216), 
        .ZN(n15215) );
  OAI221_X1 U16757 ( .B1(n15217), .B2(keyinput24), .C1(n15216), .C2(keyinput3), 
        .A(n15215), .ZN(n15227) );
  AOI22_X1 U16758 ( .A1(n8677), .A2(keyinput18), .B1(n15219), .B2(keyinput22), 
        .ZN(n15218) );
  OAI221_X1 U16759 ( .B1(n8677), .B2(keyinput18), .C1(n15219), .C2(keyinput22), 
        .A(n15218), .ZN(n15226) );
  AOI22_X1 U16760 ( .A1(n15221), .A2(keyinput6), .B1(n7091), .B2(keyinput45), 
        .ZN(n15220) );
  OAI221_X1 U16761 ( .B1(n15221), .B2(keyinput6), .C1(n7091), .C2(keyinput45), 
        .A(n15220), .ZN(n15225) );
  XOR2_X1 U16762 ( .A(n14255), .B(keyinput13), .Z(n15223) );
  XNOR2_X1 U16763 ( .A(P3_IR_REG_2__SCAN_IN), .B(keyinput30), .ZN(n15222) );
  NAND2_X1 U16764 ( .A1(n15223), .A2(n15222), .ZN(n15224) );
  NOR4_X1 U16765 ( .A1(n15227), .A2(n15226), .A3(n15225), .A4(n15224), .ZN(
        n15270) );
  AOI22_X1 U16766 ( .A1(n15229), .A2(keyinput51), .B1(keyinput62), .B2(n15281), 
        .ZN(n15228) );
  OAI221_X1 U16767 ( .B1(n15229), .B2(keyinput51), .C1(n15281), .C2(keyinput62), .A(n15228), .ZN(n15239) );
  AOI22_X1 U16768 ( .A1(n15295), .A2(keyinput57), .B1(keyinput41), .B2(n15231), 
        .ZN(n15230) );
  OAI221_X1 U16769 ( .B1(n15295), .B2(keyinput57), .C1(n15231), .C2(keyinput41), .A(n15230), .ZN(n15238) );
  XOR2_X1 U16770 ( .A(n13144), .B(keyinput2), .Z(n15234) );
  XNOR2_X1 U16771 ( .A(P3_IR_REG_8__SCAN_IN), .B(keyinput61), .ZN(n15233) );
  XNOR2_X1 U16772 ( .A(P2_IR_REG_24__SCAN_IN), .B(keyinput0), .ZN(n15232) );
  NAND3_X1 U16773 ( .A1(n15234), .A2(n15233), .A3(n15232), .ZN(n15237) );
  XNOR2_X1 U16774 ( .A(n15235), .B(keyinput12), .ZN(n15236) );
  NOR4_X1 U16775 ( .A1(n15239), .A2(n15238), .A3(n15237), .A4(n15236), .ZN(
        n15269) );
  AOI22_X1 U16776 ( .A1(n15242), .A2(keyinput38), .B1(keyinput9), .B2(n15241), 
        .ZN(n15240) );
  OAI221_X1 U16777 ( .B1(n15242), .B2(keyinput38), .C1(n15241), .C2(keyinput9), 
        .A(n15240), .ZN(n15253) );
  AOI22_X1 U16778 ( .A1(n15276), .A2(keyinput27), .B1(keyinput32), .B2(n15244), 
        .ZN(n15243) );
  OAI221_X1 U16779 ( .B1(n15276), .B2(keyinput27), .C1(n15244), .C2(keyinput32), .A(n15243), .ZN(n15252) );
  INV_X1 U16780 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n15280) );
  AOI22_X1 U16781 ( .A1(n15280), .A2(keyinput28), .B1(n15246), .B2(keyinput35), 
        .ZN(n15245) );
  OAI221_X1 U16782 ( .B1(n15280), .B2(keyinput28), .C1(n15246), .C2(keyinput35), .A(n15245), .ZN(n15251) );
  XOR2_X1 U16783 ( .A(n15247), .B(keyinput39), .Z(n15249) );
  XNOR2_X1 U16784 ( .A(SI_3_), .B(keyinput52), .ZN(n15248) );
  NAND2_X1 U16785 ( .A1(n15249), .A2(n15248), .ZN(n15250) );
  NOR4_X1 U16786 ( .A1(n15253), .A2(n15252), .A3(n15251), .A4(n15250), .ZN(
        n15268) );
  AOI22_X1 U16787 ( .A1(n15255), .A2(keyinput7), .B1(n9423), .B2(keyinput43), 
        .ZN(n15254) );
  OAI221_X1 U16788 ( .B1(n15255), .B2(keyinput7), .C1(n9423), .C2(keyinput43), 
        .A(n15254), .ZN(n15266) );
  INV_X1 U16789 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15257) );
  AOI22_X1 U16790 ( .A1(n15258), .A2(keyinput36), .B1(keyinput23), .B2(n15257), 
        .ZN(n15256) );
  OAI221_X1 U16791 ( .B1(n15258), .B2(keyinput36), .C1(n15257), .C2(keyinput23), .A(n15256), .ZN(n15265) );
  AOI22_X1 U16792 ( .A1(n13388), .A2(keyinput44), .B1(n15260), .B2(keyinput54), 
        .ZN(n15259) );
  OAI221_X1 U16793 ( .B1(n13388), .B2(keyinput44), .C1(n15260), .C2(keyinput54), .A(n15259), .ZN(n15264) );
  XNOR2_X1 U16794 ( .A(P3_REG1_REG_20__SCAN_IN), .B(keyinput29), .ZN(n15262)
         );
  XNOR2_X1 U16795 ( .A(SI_6_), .B(keyinput46), .ZN(n15261) );
  NAND2_X1 U16796 ( .A1(n15262), .A2(n15261), .ZN(n15263) );
  NOR4_X1 U16797 ( .A1(n15266), .A2(n15265), .A3(n15264), .A4(n15263), .ZN(
        n15267) );
  NAND4_X1 U16798 ( .A1(n15270), .A2(n15269), .A3(n15268), .A4(n15267), .ZN(
        n15271) );
  NOR2_X1 U16799 ( .A1(n15272), .A2(n15271), .ZN(n15315) );
  NOR4_X1 U16800 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_ADDR_REG_5__SCAN_IN), .A4(n15273), .ZN(n15274) );
  NAND4_X1 U16801 ( .A1(n15275), .A2(P1_ADDR_REG_1__SCAN_IN), .A3(
        P2_ADDR_REG_3__SCAN_IN), .A4(n15274), .ZN(n15279) );
  NAND3_X1 U16802 ( .A1(P1_REG1_REG_4__SCAN_IN), .A2(P1_REG1_REG_1__SCAN_IN), 
        .A3(n15276), .ZN(n15277) );
  OR4_X1 U16803 ( .A1(SI_3_), .A2(n15169), .A3(SI_6_), .A4(n15277), .ZN(n15278) );
  NOR4_X1 U16804 ( .A1(n15279), .A2(P3_DATAO_REG_23__SCAN_IN), .A3(n15247), 
        .A4(n15278), .ZN(n15313) );
  NOR4_X1 U16805 ( .A1(P3_D_REG_1__SCAN_IN), .A2(P3_REG2_REG_13__SCAN_IN), 
        .A3(P2_REG2_REG_20__SCAN_IN), .A4(n15280), .ZN(n15312) );
  NAND4_X1 U16806 ( .A1(P3_REG1_REG_28__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), 
        .A3(P1_REG2_REG_22__SCAN_IN), .A4(n15281), .ZN(n15285) );
  NAND4_X1 U16807 ( .A1(P3_D_REG_9__SCAN_IN), .A2(SI_19_), .A3(
        P2_REG1_REG_13__SCAN_IN), .A4(P3_DATAO_REG_14__SCAN_IN), .ZN(n15284)
         );
  NAND3_X1 U16808 ( .A1(P3_REG3_REG_2__SCAN_IN), .A2(P3_REG1_REG_30__SCAN_IN), 
        .A3(n15282), .ZN(n15283) );
  NOR4_X1 U16809 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n15285), .A3(n15284), 
        .A4(n15283), .ZN(n15311) );
  NAND4_X1 U16810 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), 
        .A3(P2_D_REG_11__SCAN_IN), .A4(n15286), .ZN(n15294) );
  INV_X1 U16811 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n15288) );
  NOR4_X1 U16812 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P1_REG0_REG_21__SCAN_IN), 
        .A3(P2_REG0_REG_13__SCAN_IN), .A4(n13144), .ZN(n15287) );
  NAND4_X1 U16813 ( .A1(n15289), .A2(n15288), .A3(P1_REG1_REG_19__SCAN_IN), 
        .A4(n15287), .ZN(n15293) );
  NAND4_X1 U16814 ( .A1(n15290), .A2(P2_IR_REG_9__SCAN_IN), .A3(
        P2_REG1_REG_25__SCAN_IN), .A4(P2_DATAO_REG_27__SCAN_IN), .ZN(n15292)
         );
  NAND2_X1 U16815 ( .A1(P3_DATAO_REG_30__SCAN_IN), .A2(
        P3_DATAO_REG_24__SCAN_IN), .ZN(n15291) );
  NOR4_X1 U16816 ( .A1(n15294), .A2(n15293), .A3(n15292), .A4(n15291), .ZN(
        n15297) );
  NOR3_X1 U16817 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        n15295), .ZN(n15296) );
  NAND2_X1 U16818 ( .A1(n15297), .A2(n15296), .ZN(n15309) );
  NOR4_X1 U16819 ( .A1(P2_REG2_REG_22__SCAN_IN), .A2(P1_REG3_REG_22__SCAN_IN), 
        .A3(n15299), .A4(n15298), .ZN(n15307) );
  NOR3_X1 U16820 ( .A1(P2_REG0_REG_5__SCAN_IN), .A2(n15301), .A3(n15300), .ZN(
        n15306) );
  NOR4_X1 U16821 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n15304), .A3(n15303), 
        .A4(n15302), .ZN(n15305) );
  NAND4_X1 U16822 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15307), .A3(n15306), .A4(
        n15305), .ZN(n15308) );
  NOR2_X1 U16823 ( .A1(n15309), .A2(n15308), .ZN(n15310) );
  NAND4_X1 U16824 ( .A1(n15313), .A2(n15312), .A3(n15311), .A4(n15310), .ZN(
        n15314) );
  XNOR2_X1 U16825 ( .A(n15315), .B(n15314), .ZN(n15316) );
  XNOR2_X1 U16826 ( .A(n15317), .B(n15316), .ZN(P1_U3486) );
  OAI21_X1 U16827 ( .B1(n15320), .B2(n15319), .A(n15318), .ZN(SUB_1596_U59) );
  OAI21_X1 U16828 ( .B1(n15323), .B2(n15322), .A(n15321), .ZN(SUB_1596_U58) );
  XOR2_X1 U16829 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15324), .Z(SUB_1596_U53) );
  AOI21_X1 U16830 ( .B1(n15327), .B2(n15326), .A(n15325), .ZN(SUB_1596_U56) );
  AOI21_X1 U16831 ( .B1(n15330), .B2(n15329), .A(n15328), .ZN(n15331) );
  XOR2_X1 U16832 ( .A(n15331), .B(P2_ADDR_REG_3__SCAN_IN), .Z(SUB_1596_U60) );
  AOI21_X1 U16833 ( .B1(n15334), .B2(n15333), .A(n15332), .ZN(SUB_1596_U5) );
  CLKBUF_X1 U7191 ( .A(n8369), .Z(n8769) );
  NAND2_X1 U10211 ( .A1(n7804), .A2(n7803), .ZN(n13080) );
  AND2_X2 U7257 ( .A1(n9048), .A2(n9834), .ZN(n9059) );
  NAND2_X2 U9019 ( .A1(n7742), .A2(n9834), .ZN(n7724) );
  CLKBUF_X1 U7196 ( .A(n9676), .Z(n6840) );
  CLKBUF_X1 U7204 ( .A(n6436), .Z(n12628) );
  CLKBUF_X1 U7207 ( .A(n7788), .Z(n9918) );
  CLKBUF_X1 U7208 ( .A(n9059), .Z(n6437) );
  OR2_X1 U7219 ( .A1(n13448), .A2(n13452), .ZN(n13450) );
  NAND4_X2 U7237 ( .A1(n7721), .A2(n7720), .A3(n7719), .A4(n7718), .ZN(n11872)
         );
  AND3_X2 U7253 ( .A1(n6695), .A2(n6750), .A3(n6751), .ZN(n15339) );
endmodule

