

module b15_C_SARLock_k_64_4 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789;

  INV_X1 U3417 ( .A(n5946), .ZN(n5937) );
  INV_X1 U3418 ( .A(n4365), .ZN(n6042) );
  BUF_X2 U3419 ( .A(n3667), .Z(n5658) );
  NAND2_X2 U3420 ( .A1(n4266), .A2(n3402), .ZN(n3578) );
  CLKBUF_X2 U3421 ( .A(n3213), .Z(n4188) );
  CLKBUF_X2 U3422 ( .A(n4070), .Z(n4229) );
  OR2_X1 U3423 ( .A1(n3177), .A2(n3176), .ZN(n3633) );
  AND2_X1 U3424 ( .A1(n3056), .A2(n4538), .ZN(n3273) );
  AND2_X1 U3425 ( .A1(n3056), .A2(n4512), .ZN(n3292) );
  INV_X2 U3426 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3754) );
  INV_X4 U3427 ( .A(n3095), .ZN(n2971) );
  CLKBUF_X2 U3428 ( .A(n3204), .Z(n4240) );
  AOI22_X1 U3429 ( .A1(keyinput5), .A2(n6703), .B1(keyinput6), .B2(n6701), 
        .ZN(n6702) );
  AND3_X1 U3430 ( .A1(n3259), .A2(n3258), .A3(n3257), .ZN(n3325) );
  INV_X1 U3431 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3538) );
  NOR2_X1 U3432 ( .A1(n4268), .A2(n4271), .ZN(n4505) );
  OAI21_X1 U3433 ( .B1(n6703), .B2(keyinput5), .A(n6702), .ZN(n6715) );
  NAND2_X1 U3434 ( .A1(n3249), .A2(n3248), .ZN(n3327) );
  NAND4_X1 U3435 ( .A1(n3212), .A2(n3211), .A3(n3210), .A4(n3209), .ZN(n3255)
         );
  INV_X1 U3438 ( .A(n3255), .ZN(n3054) );
  NOR2_X1 U3439 ( .A1(n5934), .A2(n6513), .ZN(n4975) );
  OR2_X1 U3440 ( .A1(n5192), .A2(n5210), .ZN(n5241) );
  AND2_X1 U3441 ( .A1(n5741), .A2(n5333), .ZN(n5734) );
  INV_X1 U3442 ( .A(n5968), .ZN(n5993) );
  INV_X1 U3444 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6718) );
  NAND2_X2 U34450 ( .A1(n5523), .A2(n5525), .ZN(n5506) );
  NOR2_X2 U34460 ( .A1(n5805), .A2(n3533), .ZN(n5523) );
  NOR2_X4 U34470 ( .A1(n4650), .A2(n3050), .ZN(n5930) );
  NAND2_X2 U34480 ( .A1(n3664), .A2(n3663), .ZN(n4650) );
  CLKBUF_X1 U3449 ( .A(n4101), .Z(n2968) );
  OAI22_X2 U3450 ( .A1(n5553), .A2(n5540), .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5545), .ZN(n3021) );
  NAND2_X2 U34510 ( .A1(n3397), .A2(n3015), .ZN(n4425) );
  BUF_X2 U34520 ( .A(n3293), .Z(n2969) );
  BUF_X4 U34530 ( .A(n3293), .Z(n2970) );
  NOR2_X2 U3454 ( .A1(n6042), .A2(n4367), .ZN(n6598) );
  AND2_X1 U34550 ( .A1(n5417), .A2(n5753), .ZN(n5741) );
  NAND2_X1 U34560 ( .A1(n4988), .A2(n3515), .ZN(n5063) );
  AND2_X1 U3457 ( .A1(n3736), .A2(n5658), .ZN(n4296) );
  NAND2_X1 U3458 ( .A1(n5755), .A2(REIP_REG_20__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U34590 ( .A1(n5447), .A2(REIP_REG_17__SCAN_IN), .ZN(n5898) );
  NOR2_X1 U34600 ( .A1(n5918), .A2(n5899), .ZN(n5447) );
  NAND2_X1 U34610 ( .A1(n4975), .A2(REIP_REG_8__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U34620 ( .A1(n5936), .A2(REIP_REG_6__SCAN_IN), .ZN(n5934) );
  AND2_X1 U34630 ( .A1(n3509), .A2(n3508), .ZN(n2986) );
  CLKBUF_X2 U34640 ( .A(n6089), .Z(n6101) );
  CLKBUF_X2 U34650 ( .A(n2992), .Z(n3570) );
  AND2_X1 U3466 ( .A1(n3054), .A2(n2981), .ZN(n3334) );
  INV_X1 U3467 ( .A(n3667), .ZN(n3239) );
  NAND2_X1 U34680 ( .A1(n3753), .A2(n3229), .ZN(n3232) );
  INV_X2 U34700 ( .A(n3633), .ZN(n3611) );
  INV_X1 U34710 ( .A(n3253), .ZN(n4559) );
  NAND2_X1 U34720 ( .A1(n3346), .A2(n3255), .ZN(n3667) );
  BUF_X2 U34730 ( .A(n4143), .Z(n4238) );
  BUF_X2 U34740 ( .A(n3194), .Z(n4230) );
  BUF_X2 U3475 ( .A(n4164), .Z(n4231) );
  CLKBUF_X1 U3476 ( .A(n4101), .Z(n2980) );
  BUF_X2 U3477 ( .A(n3178), .Z(n4239) );
  BUF_X2 U3478 ( .A(n3199), .Z(n4232) );
  AND2_X1 U3479 ( .A1(n5805), .A2(n5524), .ZN(n5507) );
  NAND2_X1 U3480 ( .A1(n3093), .A2(n5568), .ZN(n5567) );
  AOI21_X1 U3481 ( .B1(n5356), .B2(n6133), .A(n4327), .ZN(n4328) );
  AND2_X1 U3482 ( .A1(n5381), .A2(n5367), .ZN(n5783) );
  CLKBUF_X1 U3483 ( .A(n5378), .Z(n5379) );
  NAND2_X1 U3484 ( .A1(n3070), .A2(n3069), .ZN(n5534) );
  NAND2_X1 U3485 ( .A1(n3020), .A2(n3061), .ZN(n5220) );
  AND2_X2 U3486 ( .A1(n5419), .A2(n5474), .ZN(n5405) );
  XNOR2_X1 U3487 ( .A(n4299), .B(n4298), .ZN(n5454) );
  AND2_X2 U3488 ( .A1(n5484), .A2(n3086), .ZN(n5419) );
  AND2_X2 U3489 ( .A1(n5312), .A2(n4010), .ZN(n5484) );
  NAND2_X1 U3490 ( .A1(n4990), .A2(n4989), .ZN(n4988) );
  NAND2_X1 U3491 ( .A1(n5203), .A2(n3085), .ZN(n5287) );
  AOI21_X1 U3492 ( .B1(n2985), .B2(n3067), .A(n2996), .ZN(n3061) );
  AND2_X1 U3493 ( .A1(n3064), .A2(n2990), .ZN(n2985) );
  AOI21_X1 U3494 ( .B1(n3066), .B2(n5061), .A(n3065), .ZN(n3064) );
  AOI211_X2 U3495 ( .C1(n6364), .C2(n5137), .A(n6362), .B(n4927), .ZN(n4969)
         );
  NAND2_X1 U3496 ( .A1(n3812), .A2(n3811), .ZN(n4916) );
  INV_X4 U3497 ( .A(n2986), .ZN(n5539) );
  AND3_X1 U3498 ( .A1(n4420), .A2(n4586), .A3(n4585), .ZN(n4584) );
  AOI21_X1 U3499 ( .B1(n3799), .B2(n3936), .A(n3798), .ZN(n4652) );
  NAND2_X1 U3500 ( .A1(n3483), .A2(n3482), .ZN(n3509) );
  NAND2_X1 U3501 ( .A1(n3778), .A2(n3777), .ZN(n4420) );
  OR2_X1 U3502 ( .A1(n5977), .A2(n4358), .ZN(n5953) );
  INV_X1 U3503 ( .A(n3485), .ZN(n3483) );
  NAND2_X1 U3504 ( .A1(n4334), .A2(n4333), .ZN(n5977) );
  XNOR2_X1 U3505 ( .A(n3460), .B(n3469), .ZN(n3799) );
  NOR2_X2 U3506 ( .A1(n5241), .A2(n5240), .ZN(n5274) );
  NAND2_X1 U3507 ( .A1(n4416), .A2(n3774), .ZN(n4571) );
  OAI21_X1 U3508 ( .B1(n3779), .B2(n3887), .A(n3785), .ZN(n4586) );
  AND3_X1 U3509 ( .A1(n6491), .A2(n6602), .A3(n5357), .ZN(n4332) );
  INV_X1 U3510 ( .A(n6598), .ZN(n5357) );
  OAI21_X1 U3511 ( .B1(n4429), .B2(n3887), .A(n3769), .ZN(n3770) );
  NAND2_X1 U3512 ( .A1(n3382), .A2(n3381), .ZN(n3388) );
  AND2_X1 U3513 ( .A1(n3414), .A2(n3413), .ZN(n4489) );
  CLKBUF_X1 U3514 ( .A(n3752), .Z(n5707) );
  NAND2_X1 U3515 ( .A1(n3681), .A2(n3680), .ZN(n5055) );
  INV_X1 U3516 ( .A(n4494), .ZN(n5028) );
  INV_X1 U3517 ( .A(n4593), .ZN(n3664) );
  NAND2_X1 U3518 ( .A1(n4570), .A2(n4421), .ZN(n4593) );
  CLKBUF_X1 U3519 ( .A(n3762), .Z(n3763) );
  NAND2_X1 U3520 ( .A1(n3401), .A2(n3400), .ZN(n4409) );
  AND2_X1 U3521 ( .A1(n4568), .A2(n4567), .ZN(n4570) );
  AOI21_X1 U3522 ( .B1(n3001), .B2(n2987), .A(n3000), .ZN(n3565) );
  AND2_X1 U3523 ( .A1(n3053), .A2(n3052), .ZN(n4568) );
  AND2_X1 U3524 ( .A1(n3325), .A2(n3630), .ZN(n3261) );
  OAI21_X1 U3525 ( .B1(n3342), .B2(n3079), .A(n3507), .ZN(n3078) );
  NOR2_X1 U3526 ( .A1(n3079), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3076) );
  NAND2_X1 U3527 ( .A1(n3002), .A2(n3004), .ZN(n3001) );
  INV_X1 U3528 ( .A(n3556), .ZN(n3000) );
  INV_X1 U3529 ( .A(n4592), .ZN(n3663) );
  INV_X1 U3530 ( .A(n3484), .ZN(n3482) );
  AND2_X1 U3531 ( .A1(n3057), .A2(n3260), .ZN(n3630) );
  NAND2_X1 U3532 ( .A1(n3586), .A2(n3054), .ZN(n3616) );
  OAI21_X1 U3533 ( .B1(n3654), .B2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n3653), 
        .ZN(n3657) );
  NAND2_X1 U3534 ( .A1(n3024), .A2(n3023), .ZN(n3653) );
  INV_X1 U3535 ( .A(n3286), .ZN(n3342) );
  AND3_X1 U3536 ( .A1(n3587), .A2(n5003), .A3(n3228), .ZN(n3241) );
  OR2_X1 U3537 ( .A1(n3725), .A2(EBX_REG_1__SCAN_IN), .ZN(n3024) );
  NOR2_X1 U3538 ( .A1(n5001), .A2(n3537), .ZN(n3563) );
  INV_X1 U3539 ( .A(n3624), .ZN(n3335) );
  INV_X2 U3540 ( .A(n4254), .ZN(n4313) );
  OR2_X1 U3541 ( .A1(n2981), .A2(n6603), .ZN(n3402) );
  INV_X1 U3542 ( .A(n4271), .ZN(n5001) );
  NOR2_X1 U3543 ( .A1(n3288), .A2(n6603), .ZN(n3291) );
  INV_X1 U3544 ( .A(n3287), .ZN(n2981) );
  NAND2_X1 U3545 ( .A1(n3611), .A2(n3346), .ZN(n3624) );
  CLKBUF_X1 U3546 ( .A(n3287), .Z(n4474) );
  INV_X1 U3547 ( .A(n3287), .ZN(n2982) );
  CLKBUF_X1 U3548 ( .A(n3229), .Z(n3230) );
  OR2_X1 U3549 ( .A1(n3284), .A2(n3283), .ZN(n3390) );
  OR2_X1 U3550 ( .A1(n3303), .A2(n3302), .ZN(n3389) );
  OR2_X1 U3551 ( .A1(n3272), .A2(n3271), .ZN(n3511) );
  OR2_X1 U3552 ( .A1(n3253), .A2(n6603), .ZN(n4266) );
  AND3_X2 U3553 ( .A1(n3225), .A2(n2994), .A3(n3006), .ZN(n3287) );
  AND2_X1 U3554 ( .A1(n3012), .A2(n3226), .ZN(n3006) );
  NAND2_X1 U3555 ( .A1(n3156), .A2(n3155), .ZN(n3167) );
  AND4_X1 U3556 ( .A1(n3193), .A2(n3192), .A3(n3191), .A4(n3190), .ZN(n3212)
         );
  AND4_X1 U3557 ( .A1(n3208), .A2(n3207), .A3(n3206), .A4(n3205), .ZN(n3209)
         );
  AND4_X1 U3558 ( .A1(n3103), .A2(n3102), .A3(n3101), .A4(n3100), .ZN(n3124)
         );
  AND4_X1 U3559 ( .A1(n3164), .A2(n3163), .A3(n3162), .A4(n3161), .ZN(n3165)
         );
  AND4_X1 U3560 ( .A1(n3154), .A2(n3153), .A3(n3152), .A4(n3151), .ZN(n3155)
         );
  AND4_X1 U3561 ( .A1(n3148), .A2(n3147), .A3(n3146), .A4(n3145), .ZN(n3156)
         );
  AND4_X1 U3562 ( .A1(n3217), .A2(n3216), .A3(n3215), .A4(n3214), .ZN(n3226)
         );
  AND4_X1 U3563 ( .A1(n3140), .A2(n3139), .A3(n3138), .A4(n3137), .ZN(n3141)
         );
  AND4_X1 U3564 ( .A1(n3198), .A2(n3197), .A3(n3196), .A4(n3195), .ZN(n3211)
         );
  AND2_X1 U3565 ( .A1(n3150), .A2(n3149), .ZN(n3152) );
  AND4_X1 U3566 ( .A1(n3128), .A2(n3127), .A3(n3126), .A4(n3125), .ZN(n3144)
         );
  AND4_X1 U3567 ( .A1(n3160), .A2(n3159), .A3(n3158), .A4(n3157), .ZN(n3166)
         );
  AND4_X1 U3568 ( .A1(n3203), .A2(n3202), .A3(n3201), .A4(n3200), .ZN(n3210)
         );
  AND4_X1 U3569 ( .A1(n3136), .A2(n3135), .A3(n3134), .A4(n3133), .ZN(n3142)
         );
  AND4_X1 U3570 ( .A1(n3114), .A2(n3113), .A3(n3112), .A4(n3111), .ZN(n3122)
         );
  AND4_X1 U3571 ( .A1(n3222), .A2(n3221), .A3(n3220), .A4(n3219), .ZN(n3225)
         );
  NOR2_X1 U3572 ( .A1(n6145), .A2(n6720), .ZN(n6402) );
  INV_X2 U3573 ( .A(n6145), .ZN(n6133) );
  AND4_X1 U3574 ( .A1(n3109), .A2(n3108), .A3(n3107), .A4(n3106), .ZN(n3123)
         );
  AND4_X1 U3575 ( .A1(n3120), .A2(n3119), .A3(n3118), .A4(n3117), .ZN(n3121)
         );
  BUF_X2 U3576 ( .A(n3273), .Z(n4237) );
  INV_X1 U3577 ( .A(n4317), .ZN(n3399) );
  OR2_X1 U3578 ( .A1(n6586), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4317) );
  INV_X2 U3579 ( .A(n6611), .ZN(n6597) );
  AND2_X2 U3580 ( .A1(n3116), .A2(n3056), .ZN(n4164) );
  AND2_X2 U3581 ( .A1(n3110), .A2(n4504), .ZN(n4101) );
  AND2_X1 U3582 ( .A1(n3104), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3115)
         );
  NAND2_X2 U3583 ( .A1(n6718), .A2(n6601), .ZN(n6364) );
  AND2_X2 U3584 ( .A1(n4512), .A2(n4504), .ZN(n3183) );
  AND2_X1 U3585 ( .A1(n3099), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3056)
         );
  INV_X1 U3586 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6634) );
  INV_X2 U3587 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6603) );
  AND2_X2 U3588 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4504) );
  NOR2_X2 U3589 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4519) );
  OR2_X1 U3590 ( .A1(n4911), .A2(n4854), .ZN(n2972) );
  OR2_X1 U3591 ( .A1(n4855), .A2(n4854), .ZN(n4853) );
  NOR2_X1 U3592 ( .A1(n5406), .A2(n5464), .ZN(n2973) );
  INV_X1 U3593 ( .A(n5207), .ZN(n2974) );
  INV_X1 U3594 ( .A(n5715), .ZN(n2975) );
  XNOR2_X1 U3595 ( .A(n4316), .B(n4315), .ZN(n2976) );
  OR2_X1 U3596 ( .A1(n3379), .A2(n3378), .ZN(n2977) );
  NAND2_X1 U3597 ( .A1(n2977), .A2(n3377), .ZN(n3383) );
  INV_X1 U3598 ( .A(n3595), .ZN(n2978) );
  NOR2_X1 U3599 ( .A1(n5406), .A2(n5464), .ZN(n5394) );
  AOI21_X1 U3600 ( .B1(n5187), .B2(n5204), .A(n5205), .ZN(n5203) );
  XNOR2_X1 U3601 ( .A(n3329), .B(n3328), .ZN(n4427) );
  XNOR2_X1 U3602 ( .A(n4316), .B(n4315), .ZN(n5356) );
  NAND2_X1 U3603 ( .A1(n3077), .A2(n3075), .ZN(n3379) );
  NAND2_X1 U3604 ( .A1(n3332), .A2(n3331), .ZN(n3377) );
  AND2_X1 U3605 ( .A1(n3383), .A2(n3380), .ZN(n3381) );
  NOR2_X1 U3606 ( .A1(n3312), .A2(n3092), .ZN(n3586) );
  OAI21_X1 U3607 ( .B1(n5672), .B2(n3531), .A(n3060), .ZN(n5807) );
  AND2_X1 U3608 ( .A1(n5672), .A2(n5535), .ZN(n3093) );
  NOR2_X1 U3609 ( .A1(n4652), .A2(n4667), .ZN(n3804) );
  AND2_X1 U3610 ( .A1(n3240), .A2(n4508), .ZN(n3258) );
  NAND2_X1 U3611 ( .A1(n5186), .A2(n5189), .ZN(n5187) );
  AND2_X2 U3612 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4512) );
  AND2_X1 U3613 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4511) );
  NAND2_X1 U3614 ( .A1(n6122), .A2(n6121), .ZN(n6120) );
  XNOR2_X1 U3615 ( .A(n3425), .B(n3424), .ZN(n6122) );
  INV_X1 U3616 ( .A(n3907), .ZN(n5068) );
  NAND2_X1 U3617 ( .A1(n4336), .A2(n3082), .ZN(n3907) );
  AND2_X2 U3618 ( .A1(n4512), .A2(n4504), .ZN(n2979) );
  AND2_X2 U3619 ( .A1(n3754), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3116)
         );
  NOR2_X1 U3620 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3105) );
  INV_X1 U3621 ( .A(n3468), .ZN(n3447) );
  NAND2_X2 U3622 ( .A1(n3468), .A2(n3418), .ZN(n3779) );
  OAI21_X2 U3623 ( .B1(n5220), .B2(n5223), .A(n5221), .ZN(n5246) );
  NAND2_X2 U3624 ( .A1(n3014), .A2(n3018), .ZN(n3397) );
  AND2_X2 U3625 ( .A1(n4584), .A2(n3804), .ZN(n4666) );
  AND4_X1 U3626 ( .A1(n3132), .A2(n3131), .A3(n3130), .A4(n3129), .ZN(n3143)
         );
  OAI22_X2 U3627 ( .A1(n4425), .A2(STATE2_REG_0__SCAN_IN), .B1(n3419), .B2(
        n4266), .ZN(n3385) );
  AND2_X1 U3628 ( .A1(n5370), .A2(n5369), .ZN(n5780) );
  XNOR2_X1 U3629 ( .A(n5370), .B(n2997), .ZN(n5327) );
  XNOR2_X2 U3630 ( .A(n3907), .B(n3908), .ZN(n5186) );
  AND2_X2 U3631 ( .A1(n3116), .A2(n3115), .ZN(n3213) );
  NOR2_X2 U3632 ( .A1(n3308), .A2(n3589), .ZN(n3608) );
  BUF_X4 U3633 ( .A(n3334), .Z(n2984) );
  NAND2_X2 U3634 ( .A1(n3388), .A2(n3417), .ZN(n4429) );
  NOR2_X1 U3635 ( .A1(n3088), .A2(n5434), .ZN(n3087) );
  INV_X1 U3636 ( .A(n5569), .ZN(n3088) );
  OR2_X1 U3637 ( .A1(n6431), .A2(n6603), .ZN(n4154) );
  NAND2_X1 U3638 ( .A1(n3755), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4254) );
  NAND2_X1 U3639 ( .A1(n5378), .A2(n3089), .ZN(n5370) );
  NOR2_X1 U3640 ( .A1(n5368), .A2(n3090), .ZN(n3089) );
  INV_X1 U3641 ( .A(n5380), .ZN(n3090) );
  NAND2_X1 U3642 ( .A1(n6468), .A2(n4273), .ZN(n6043) );
  INV_X1 U3643 ( .A(n4418), .ZN(n4297) );
  OR2_X1 U3644 ( .A1(n5539), .A2(n3524), .ZN(n3525) );
  OAI21_X1 U3645 ( .B1(n3522), .B2(n3072), .A(n3521), .ZN(n3071) );
  NAND2_X1 U3646 ( .A1(n5279), .A2(n5280), .ZN(n3072) );
  NAND2_X1 U3647 ( .A1(n5278), .A2(n3073), .ZN(n3070) );
  NOR2_X1 U3648 ( .A1(n3522), .A2(n3074), .ZN(n3073) );
  OR2_X1 U3649 ( .A1(n5539), .A2(n3517), .ZN(n3518) );
  INV_X1 U3650 ( .A(n5061), .ZN(n3067) );
  NAND2_X1 U3651 ( .A1(n3363), .A2(n3362), .ZN(n3018) );
  OR2_X1 U3652 ( .A1(n5408), .A2(n5465), .ZN(n5466) );
  NAND2_X1 U3653 ( .A1(n4341), .A2(n3095), .ZN(n5015) );
  NAND2_X1 U3654 ( .A1(n4664), .A2(n3051), .ZN(n3050) );
  INV_X1 U3655 ( .A(n4649), .ZN(n3051) );
  AND2_X1 U3656 ( .A1(n6601), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4312) );
  INV_X1 U3657 ( .A(n5397), .ZN(n4161) );
  AND2_X1 U3658 ( .A1(n4339), .A2(n5758), .ZN(n4024) );
  AND2_X1 U3659 ( .A1(n3975), .A2(n2998), .ZN(n3085) );
  INV_X1 U3660 ( .A(n5288), .ZN(n3975) );
  NOR2_X1 U3661 ( .A1(n3920), .A2(n3919), .ZN(n3924) );
  NAND2_X1 U3662 ( .A1(n6120), .A2(n3426), .ZN(n4583) );
  NOR2_X2 U3663 ( .A1(n5466), .A2(n5398), .ZN(n5605) );
  AND2_X1 U3664 ( .A1(n5539), .A2(n6674), .ZN(n3533) );
  NAND2_X1 U3665 ( .A1(n5560), .A2(n5551), .ZN(n5545) );
  AND2_X1 U3666 ( .A1(n5539), .A2(n5299), .ZN(n5280) );
  INV_X1 U3667 ( .A(n5107), .ZN(n3065) );
  INV_X1 U3668 ( .A(n5060), .ZN(n3066) );
  OR2_X1 U3669 ( .A1(n5063), .A2(n3067), .ZN(n3062) );
  OR2_X1 U3670 ( .A1(n5539), .A2(n3516), .ZN(n5128) );
  OR2_X1 U3671 ( .A1(n5702), .A2(n5255), .ZN(n5684) );
  NAND2_X1 U3672 ( .A1(n3615), .A2(n3614), .ZN(n3742) );
  OR2_X1 U3673 ( .A1(n6043), .A2(n3613), .ZN(n3614) );
  AND2_X1 U3674 ( .A1(n2978), .A2(n3227), .ZN(n6434) );
  OR2_X1 U3675 ( .A1(n3779), .A2(n4463), .ZN(n4622) );
  INV_X1 U3676 ( .A(n4429), .ZN(n4463) );
  CLKBUF_X1 U3677 ( .A(n4424), .Z(n4924) );
  AND2_X1 U3678 ( .A1(n3577), .A2(n3576), .ZN(n3602) );
  AND2_X1 U3679 ( .A1(n6459), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3574)
         );
  OAI22_X1 U3680 ( .A1(n3565), .A2(n3564), .B1(n3570), .B2(n3599), .ZN(n3572)
         );
  NAND2_X1 U3681 ( .A1(n3570), .A2(n3547), .ZN(n3582) );
  INV_X2 U3682 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6601) );
  NAND2_X1 U3683 ( .A1(n3005), .A2(n3618), .ZN(n4365) );
  INV_X1 U3684 ( .A(n6043), .ZN(n3005) );
  AND3_X1 U3685 ( .A1(n3736), .A2(n3047), .A3(n3046), .ZN(n3737) );
  INV_X1 U3686 ( .A(n5961), .ZN(n5982) );
  NAND2_X2 U3687 ( .A1(n4284), .A2(n4283), .ZN(n5997) );
  AND2_X1 U3688 ( .A1(n5200), .A2(n4278), .ZN(n6009) );
  AND2_X1 U3689 ( .A1(n5200), .A2(n4276), .ZN(n6006) );
  XNOR2_X1 U3690 ( .A(n4324), .B(n4323), .ZN(n4343) );
  OR2_X1 U3691 ( .A1(n4322), .A2(n5325), .ZN(n4324) );
  XNOR2_X1 U3692 ( .A(n4292), .B(n5349), .ZN(n4307) );
  NAND2_X1 U3693 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6468), .ZN(n6578) );
  OR2_X1 U3694 ( .A1(n4822), .A2(n4731), .ZN(n4754) );
  NAND2_X1 U3695 ( .A1(n4101), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3140)
         );
  NAND2_X1 U3696 ( .A1(n3232), .A2(n4559), .ZN(n3236) );
  NAND2_X1 U3697 ( .A1(n3447), .A2(n3097), .ZN(n3485) );
  AND2_X1 U3698 ( .A1(n3481), .A2(n3480), .ZN(n3484) );
  OR2_X1 U3699 ( .A1(n3436), .A2(n3435), .ZN(n3487) );
  OR2_X1 U3700 ( .A1(n3457), .A2(n3456), .ZN(n3486) );
  OR2_X1 U3701 ( .A1(n3374), .A2(n3373), .ZN(n3391) );
  NAND2_X1 U3702 ( .A1(n3253), .A2(n3091), .ZN(n3250) );
  OAI211_X1 U3703 ( .C1(n3254), .C2(n3253), .A(n4275), .B(n3232), .ZN(n3081)
         );
  AOI21_X1 U3704 ( .B1(n3199), .B2(INSTQUEUE_REG_0__0__SCAN_IN), .A(n3013), 
        .ZN(n3012) );
  NAND2_X1 U3705 ( .A1(n3223), .A2(n3224), .ZN(n3013) );
  NOR2_X1 U3706 ( .A1(n3009), .A2(n2991), .ZN(n3008) );
  AND2_X1 U3707 ( .A1(n3292), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3009) );
  NAND2_X1 U3708 ( .A1(n3178), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3007)
         );
  NAND2_X1 U3709 ( .A1(n3194), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3010) );
  NAND2_X1 U3710 ( .A1(n3204), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3011) );
  NAND2_X1 U3711 ( .A1(n3003), .A2(n3582), .ZN(n3002) );
  NOR2_X1 U3712 ( .A1(n5069), .A2(n3083), .ZN(n3082) );
  INV_X1 U3713 ( .A(n3084), .ZN(n3083) );
  AND2_X1 U3714 ( .A1(n4997), .A2(n4337), .ZN(n3084) );
  NAND2_X1 U3715 ( .A1(n3447), .A2(n3096), .ZN(n3460) );
  NOR2_X1 U3716 ( .A1(n3071), .A2(n2995), .ZN(n3069) );
  AND2_X1 U3717 ( .A1(n3673), .A2(n3672), .ZN(n4849) );
  NAND2_X1 U3718 ( .A1(n5658), .A2(EBX_REG_1__SCAN_IN), .ZN(n3023) );
  INV_X1 U3719 ( .A(n4308), .ZN(n3619) );
  OR2_X1 U3720 ( .A1(n3412), .A2(n3411), .ZN(n3439) );
  AND2_X1 U3721 ( .A1(n3398), .A2(n4726), .ZN(n4681) );
  AOI22_X1 U3722 ( .A1(n4143), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3154) );
  INV_X1 U3723 ( .A(n4683), .ZN(n4771) );
  XNOR2_X1 U3724 ( .A(n3397), .B(n4409), .ZN(n4424) );
  OAI21_X1 U3725 ( .B1(n6607), .B2(n6473), .A(n6578), .ZN(n4430) );
  INV_X1 U3726 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6442) );
  OR2_X1 U3727 ( .A1(n3575), .A2(n3576), .ZN(n3600) );
  NAND2_X1 U3728 ( .A1(n3238), .A2(n4559), .ZN(n4308) );
  CLKBUF_X1 U3729 ( .A(n3617), .Z(n3618) );
  OR2_X1 U3730 ( .A1(n3733), .A2(n5658), .ZN(n3047) );
  NAND2_X1 U3731 ( .A1(n3733), .A2(n3732), .ZN(n3736) );
  AND2_X2 U3732 ( .A1(n5382), .A2(n5383), .ZN(n3733) );
  NAND2_X1 U3733 ( .A1(n3227), .A2(n3287), .ZN(n5003) );
  AND2_X1 U3734 ( .A1(n4100), .A2(n4099), .ZN(n5474) );
  NAND2_X1 U3735 ( .A1(n3038), .A2(n3037), .ZN(n3692) );
  NAND2_X1 U3736 ( .A1(n5658), .A2(EBX_REG_16__SCAN_IN), .ZN(n3037) );
  NAND2_X1 U3737 ( .A1(n3036), .A2(n3035), .ZN(n3689) );
  NAND2_X1 U3738 ( .A1(n5658), .A2(EBX_REG_14__SCAN_IN), .ZN(n3035) );
  NAND2_X1 U3739 ( .A1(n3032), .A2(n3031), .ZN(n3670) );
  NAND2_X1 U3740 ( .A1(n5658), .A2(EBX_REG_8__SCAN_IN), .ZN(n3031) );
  NAND2_X1 U3741 ( .A1(n3030), .A2(n3029), .ZN(n3668) );
  NAND2_X1 U3742 ( .A1(n5658), .A2(EBX_REG_6__SCAN_IN), .ZN(n3029) );
  NAND2_X1 U3743 ( .A1(n3028), .A2(n3027), .ZN(n3662) );
  NAND2_X1 U3744 ( .A1(n5658), .A2(EBX_REG_4__SCAN_IN), .ZN(n3027) );
  INV_X1 U3745 ( .A(n5370), .ZN(n4311) );
  OR2_X1 U3746 ( .A1(n4227), .A2(n4226), .ZN(n5368) );
  AND2_X1 U3747 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n4182), .ZN(n4183)
         );
  NAND2_X1 U3748 ( .A1(n4183), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4223)
         );
  NAND2_X1 U3749 ( .A1(n4135), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4181)
         );
  NOR2_X1 U3750 ( .A1(n4095), .A2(n5554), .ZN(n4096) );
  AND2_X1 U3751 ( .A1(n4096), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4113)
         );
  AND2_X1 U3752 ( .A1(n3087), .A2(n4064), .ZN(n3086) );
  INV_X1 U3753 ( .A(n5418), .ZN(n4064) );
  AND2_X1 U3754 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n4042), .ZN(n4043)
         );
  INV_X1 U3755 ( .A(n4041), .ZN(n4042) );
  NAND2_X1 U3756 ( .A1(n4043), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4095)
         );
  NOR2_X1 U3757 ( .A1(n3993), .A2(n3992), .ZN(n3994) );
  NAND2_X1 U3758 ( .A1(n3994), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4041)
         );
  INV_X1 U3759 ( .A(n5312), .ZN(n5486) );
  AND2_X1 U3760 ( .A1(n3970), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3971)
         );
  NAND2_X1 U3761 ( .A1(n3971), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3993)
         );
  NOR2_X1 U3762 ( .A1(n3939), .A2(n5907), .ZN(n3970) );
  NAND2_X1 U3763 ( .A1(n3924), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3939)
         );
  AND2_X1 U3764 ( .A1(n2974), .A2(n5238), .ZN(n5237) );
  NAND2_X1 U3765 ( .A1(n5068), .A2(n3908), .ZN(n5204) );
  AND3_X1 U3766 ( .A1(n3923), .A2(n3922), .A3(n3921), .ZN(n5205) );
  NAND2_X1 U3767 ( .A1(n3891), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3920)
         );
  CLKBUF_X1 U3768 ( .A(n5187), .Z(n5188) );
  INV_X1 U3769 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6703) );
  NOR2_X1 U3770 ( .A1(n6703), .A2(n3857), .ZN(n3891) );
  NOR2_X1 U3771 ( .A1(n3842), .A2(n5101), .ZN(n3856) );
  OR2_X1 U3772 ( .A1(n3827), .A2(n4979), .ZN(n3842) );
  NOR2_X1 U3773 ( .A1(n3807), .A2(n3806), .ZN(n3808) );
  NAND2_X1 U3774 ( .A1(n3795), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3807)
         );
  NOR2_X1 U3775 ( .A1(n3790), .A2(n5964), .ZN(n3795) );
  INV_X1 U3776 ( .A(n3780), .ZN(n3781) );
  NAND2_X1 U3777 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3780) );
  NOR2_X1 U3778 ( .A1(n5506), .A2(n3748), .ZN(n4291) );
  INV_X1 U3779 ( .A(n3733), .ZN(n5385) );
  NAND2_X1 U3780 ( .A1(n3530), .A2(n5539), .ZN(n3060) );
  NAND2_X1 U3781 ( .A1(n3040), .A2(n3039), .ZN(n3711) );
  NAND2_X1 U3782 ( .A1(n5658), .A2(EBX_REG_23__SCAN_IN), .ZN(n3039) );
  OR2_X1 U3783 ( .A1(n5657), .A2(n3704), .ZN(n5438) );
  NAND2_X1 U3784 ( .A1(n5292), .A2(n3048), .ZN(n5657) );
  NOR2_X1 U3785 ( .A1(n5488), .A2(n3049), .ZN(n3048) );
  INV_X1 U3786 ( .A(n5291), .ZN(n3049) );
  NAND2_X1 U3787 ( .A1(n5671), .A2(n5679), .ZN(n5672) );
  INV_X1 U3788 ( .A(n3071), .ZN(n3068) );
  NAND2_X1 U3789 ( .A1(n3034), .A2(n3033), .ZN(n3685) );
  NAND2_X1 U3790 ( .A1(n5658), .A2(EBX_REG_12__SCAN_IN), .ZN(n3033) );
  NAND2_X1 U3791 ( .A1(n5063), .A2(n2985), .ZN(n3020) );
  INV_X1 U3792 ( .A(n5225), .ZN(n5656) );
  NOR2_X1 U3793 ( .A1(n4349), .A2(n4912), .ZN(n3680) );
  INV_X1 U3794 ( .A(n4348), .ZN(n3681) );
  AND2_X1 U3795 ( .A1(n3058), .A2(n3019), .ZN(n6121) );
  OR2_X1 U3796 ( .A1(n6131), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3019)
         );
  NAND2_X1 U3797 ( .A1(n3026), .A2(n3025), .ZN(n3658) );
  NAND2_X1 U3798 ( .A1(n5658), .A2(EBX_REG_2__SCAN_IN), .ZN(n3025) );
  NAND2_X1 U3799 ( .A1(n3017), .A2(n3016), .ZN(n3015) );
  OR2_X1 U3800 ( .A1(n4931), .A2(n5707), .ZN(n5029) );
  OR2_X1 U3801 ( .A1(n4429), .A2(n3415), .ZN(n6260) );
  INV_X1 U3802 ( .A(n4622), .ZN(n4628) );
  OAI21_X1 U3803 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6718), .A(n4771), 
        .ZN(n6362) );
  OR2_X1 U3804 ( .A1(n5707), .A2(n5028), .ZN(n6229) );
  OR2_X1 U3805 ( .A1(n4429), .A2(n4489), .ZN(n4822) );
  NOR2_X1 U3806 ( .A1(n4368), .A2(n6474), .ZN(n4367) );
  AND2_X1 U3807 ( .A1(n4357), .A2(n5357), .ZN(n5967) );
  AND2_X1 U3808 ( .A1(n4354), .A2(n4347), .ZN(n5961) );
  AND2_X1 U3809 ( .A1(n4343), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4344) );
  AND2_X1 U3810 ( .A1(n5015), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U3811 ( .A1(n4914), .A2(n4913), .ZN(n5244) );
  AOI21_X1 U3812 ( .B1(n4407), .B2(n4273), .A(n4272), .ZN(n4274) );
  INV_X1 U3813 ( .A(n5244), .ZN(n5201) );
  INV_X1 U3814 ( .A(n6006), .ZN(n5499) );
  OR3_X1 U3815 ( .A1(n6043), .A2(n4440), .A3(n6490), .ZN(n6038) );
  INV_X1 U3817 ( .A(n6038), .ZN(n6040) );
  NOR2_X1 U3818 ( .A1(n5379), .A2(n5519), .ZN(n5786) );
  NAND2_X1 U3819 ( .A1(n5484), .A2(n5569), .ZN(n5435) );
  NOR2_X1 U3820 ( .A1(n2989), .A2(n3042), .ZN(n3041) );
  INV_X1 U3821 ( .A(n5323), .ZN(n3042) );
  AND2_X1 U3822 ( .A1(n5827), .A2(n5619), .ZN(n5608) );
  OR2_X1 U3823 ( .A1(n5382), .A2(n5606), .ZN(n5774) );
  XNOR2_X1 U3824 ( .A(n3021), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5629)
         );
  OR2_X1 U3825 ( .A1(n5644), .A2(n3746), .ZN(n5631) );
  AND2_X1 U3826 ( .A1(n5833), .A2(n3745), .ZN(n5676) );
  AND2_X1 U3827 ( .A1(n5489), .A2(n5319), .ZN(n5895) );
  OAI21_X1 U3828 ( .B1(n5278), .B2(n5280), .A(n5279), .ZN(n5298) );
  NAND2_X1 U3829 ( .A1(n3062), .A2(n3064), .ZN(n5129) );
  NAND2_X1 U3830 ( .A1(n5063), .A2(n5060), .ZN(n3063) );
  NOR2_X1 U3831 ( .A1(n3646), .A2(n4481), .ZN(n6217) );
  INV_X1 U3832 ( .A(n6198), .ZN(n6218) );
  AND2_X1 U3833 ( .A1(n3742), .A2(n6434), .ZN(n5702) );
  INV_X1 U3834 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6356) );
  CLKBUF_X1 U3835 ( .A(n4425), .Z(n4426) );
  INV_X1 U3836 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6446) );
  INV_X1 U3837 ( .A(n5176), .ZN(n5182) );
  INV_X1 U3838 ( .A(n6265), .ZN(n6295) );
  OR2_X1 U3839 ( .A1(n6260), .A2(n4676), .ZN(n4719) );
  NOR2_X1 U3840 ( .A1(n4986), .A2(n4683), .ZN(n6286) );
  NOR2_X1 U3841 ( .A1(n6080), .A2(n4683), .ZN(n6350) );
  OAI211_X1 U3842 ( .C1(n4738), .C2(n6718), .A(n4737), .B(n4736), .ZN(n4764)
         );
  INV_X1 U3843 ( .A(n4754), .ZN(n6411) );
  OR2_X1 U3844 ( .A1(n4822), .A2(n6229), .ZN(n6777) );
  NOR2_X1 U3845 ( .A1(n6067), .A2(n4683), .ZN(n6421) );
  INV_X1 U3846 ( .A(n6423), .ZN(n4905) );
  OR2_X1 U3847 ( .A1(n4822), .A2(n4676), .ZN(n6423) );
  INV_X1 U3848 ( .A(n6350), .ZN(n6786) );
  OR2_X1 U3849 ( .A1(n3582), .A2(n3581), .ZN(n3583) );
  INV_X1 U3850 ( .A(n6553), .ZN(n6555) );
  NAND2_X1 U3851 ( .A1(n3045), .A2(n3044), .ZN(n4285) );
  OR2_X1 U3852 ( .A1(n5997), .A2(n5336), .ZN(n3044) );
  OAI21_X1 U3853 ( .B1(n4307), .B2(n6137), .A(n4328), .ZN(U2955) );
  NAND2_X1 U3854 ( .A1(n2974), .A2(n2998), .ZN(n5270) );
  NAND2_X1 U3855 ( .A1(n4336), .A2(n3084), .ZN(n4996) );
  OR2_X2 U3856 ( .A1(n3729), .A2(n2983), .ZN(n3654) );
  NAND2_X1 U3857 ( .A1(n3070), .A2(n3068), .ZN(n5573) );
  AND2_X2 U3858 ( .A1(n4538), .A2(n4504), .ZN(n3178) );
  AND2_X2 U3859 ( .A1(n3115), .A2(n4538), .ZN(n3194) );
  OR3_X1 U3860 ( .A1(n3551), .A2(n6603), .A3(n3550), .ZN(n2987) );
  NAND2_X1 U3861 ( .A1(n5484), .A2(n3087), .ZN(n2988) );
  NAND2_X1 U3862 ( .A1(n5507), .A2(n3532), .ZN(n4289) );
  INV_X1 U3863 ( .A(n3529), .ZN(n5671) );
  AND3_X1 U3864 ( .A1(n5608), .A2(n4300), .A3(n3535), .ZN(n2989) );
  NAND2_X1 U3865 ( .A1(n5539), .A2(n3517), .ZN(n2990) );
  AND2_X1 U3866 ( .A1(n3183), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n2991) );
  AND2_X1 U3867 ( .A1(n3253), .A2(n3055), .ZN(n2992) );
  NAND2_X1 U3868 ( .A1(n3254), .A2(n3253), .ZN(n2993) );
  AND4_X1 U3869 ( .A1(n3011), .A2(n3010), .A3(n3008), .A4(n3007), .ZN(n2994)
         );
  AND2_X1 U3870 ( .A1(n5539), .A2(n3523), .ZN(n2995) );
  NAND2_X1 U3871 ( .A1(n5128), .A2(n3518), .ZN(n2996) );
  NAND2_X1 U3872 ( .A1(n5409), .A2(n5410), .ZN(n5408) );
  AND2_X1 U3873 ( .A1(n5605), .A2(n5604), .ZN(n5382) );
  INV_X1 U3874 ( .A(n6097), .ZN(n6102) );
  BUF_X1 U3875 ( .A(n3167), .Z(n3753) );
  NAND2_X1 U3876 ( .A1(n5070), .A2(n5193), .ZN(n5192) );
  AND2_X1 U3877 ( .A1(n4336), .A2(n4337), .ZN(n4335) );
  NAND2_X1 U3878 ( .A1(n3063), .A2(n5061), .ZN(n5108) );
  INV_X1 U3879 ( .A(n5279), .ZN(n3074) );
  AND2_X1 U3880 ( .A1(n4608), .A2(n4275), .ZN(n3091) );
  NAND2_X1 U3881 ( .A1(n5292), .A2(n5291), .ZN(n5290) );
  AND2_X1 U3882 ( .A1(n4260), .A2(n4259), .ZN(n2997) );
  AND2_X1 U3883 ( .A1(n3238), .A2(n3227), .ZN(n3547) );
  INV_X1 U3884 ( .A(n3547), .ZN(n3561) );
  NAND2_X1 U3885 ( .A1(n5997), .A2(n3755), .ZN(n5773) );
  INV_X1 U3886 ( .A(n5773), .ZN(n5995) );
  NOR2_X1 U3887 ( .A1(n4650), .A2(n4649), .ZN(n4648) );
  AND2_X1 U3888 ( .A1(n5271), .A2(n5238), .ZN(n2998) );
  NAND2_X1 U3889 ( .A1(n5930), .A2(n3674), .ZN(n4348) );
  AND2_X1 U3890 ( .A1(n4505), .A2(n4277), .ZN(n3621) );
  INV_X1 U3891 ( .A(n4294), .ZN(n3046) );
  NOR2_X1 U3892 ( .A1(n4609), .A2(n3755), .ZN(n2999) );
  NAND2_X1 U3893 ( .A1(n6565), .A2(n4430), .ZN(n4609) );
  OR2_X1 U3894 ( .A1(n6482), .A2(n6364), .ZN(n6145) );
  OAI211_X1 U3895 ( .C1(n3549), .C2(n3597), .A(n3546), .B(n3545), .ZN(n3003)
         );
  NAND2_X1 U3896 ( .A1(n3548), .A2(n3597), .ZN(n3004) );
  NOR2_X2 U3897 ( .A1(n5898), .A2(n5766), .ZN(n5755) );
  NAND2_X2 U3898 ( .A1(n3584), .A2(n3583), .ZN(n6468) );
  NAND2_X1 U3899 ( .A1(n5339), .A2(n6542), .ZN(n5417) );
  NOR2_X2 U3900 ( .A1(n5190), .A2(n5191), .ZN(n5925) );
  INV_X2 U3901 ( .A(n3287), .ZN(n4441) );
  NAND2_X1 U3902 ( .A1(n3054), .A2(n3287), .ZN(n4271) );
  INV_X1 U3903 ( .A(n3018), .ZN(n3016) );
  INV_X1 U3904 ( .A(n3017), .ZN(n3014) );
  NAND2_X1 U3905 ( .A1(n3358), .A2(n3357), .ZN(n3017) );
  OAI21_X2 U3906 ( .B1(n3779), .B2(n3561), .A(n3423), .ZN(n3425) );
  NAND2_X2 U3907 ( .A1(n3022), .A2(n3520), .ZN(n5278) );
  NAND2_X1 U3908 ( .A1(n5246), .A2(n5247), .ZN(n3022) );
  AND2_X2 U3909 ( .A1(n4538), .A2(n4519), .ZN(n3199) );
  NOR2_X4 U3910 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4538) );
  NAND3_X1 U3911 ( .A1(n3241), .A2(n3258), .A3(n3057), .ZN(n3080) );
  NAND2_X1 U3912 ( .A1(n5001), .A2(n3312), .ZN(n3057) );
  OR2_X1 U3913 ( .A1(n3725), .A2(EBX_REG_2__SCAN_IN), .ZN(n3026) );
  OR2_X1 U3914 ( .A1(n3725), .A2(EBX_REG_4__SCAN_IN), .ZN(n3028) );
  OR2_X1 U3915 ( .A1(n3725), .A2(EBX_REG_6__SCAN_IN), .ZN(n3030) );
  OR2_X1 U3916 ( .A1(n3725), .A2(EBX_REG_8__SCAN_IN), .ZN(n3032) );
  OR2_X1 U3917 ( .A1(n3725), .A2(EBX_REG_12__SCAN_IN), .ZN(n3034) );
  OR2_X1 U3918 ( .A1(n3725), .A2(EBX_REG_14__SCAN_IN), .ZN(n3036) );
  OR2_X1 U3919 ( .A1(n3725), .A2(EBX_REG_16__SCAN_IN), .ZN(n3038) );
  OR2_X1 U3920 ( .A1(n3725), .A2(EBX_REG_23__SCAN_IN), .ZN(n3040) );
  AND2_X2 U3921 ( .A1(n4418), .A2(n5658), .ZN(n3725) );
  NAND2_X1 U3922 ( .A1(n3043), .A2(n3041), .ZN(n3749) );
  NAND2_X1 U3923 ( .A1(n5346), .A2(n4302), .ZN(n3043) );
  NAND2_X1 U3924 ( .A1(n5346), .A2(n5995), .ZN(n3045) );
  INV_X1 U3925 ( .A(n3657), .ZN(n3052) );
  NAND2_X1 U3926 ( .A1(n4417), .A2(n4418), .ZN(n3053) );
  AND2_X2 U3927 ( .A1(n5477), .A2(n5476), .ZN(n5409) );
  AND2_X2 U3928 ( .A1(n5426), .A2(n5425), .ZN(n5477) );
  AND2_X2 U3929 ( .A1(n5053), .A2(n3686), .ZN(n5070) );
  NOR2_X2 U3930 ( .A1(n5055), .A2(n5054), .ZN(n5053) );
  AND2_X1 U3931 ( .A1(n2982), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3055) );
  AND2_X1 U3932 ( .A1(n3309), .A2(n4441), .ZN(n3729) );
  AND2_X2 U3933 ( .A1(n4519), .A2(n4512), .ZN(n3204) );
  AND2_X2 U3934 ( .A1(n3110), .A2(n4519), .ZN(n4143) );
  AND2_X2 U3935 ( .A1(n3116), .A2(n4519), .ZN(n4070) );
  NAND2_X1 U3936 ( .A1(n3059), .A2(n6129), .ZN(n3058) );
  NAND2_X1 U3937 ( .A1(n6131), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3059)
         );
  AND2_X2 U3938 ( .A1(n5807), .A2(n5808), .ZN(n5805) );
  NAND2_X1 U3939 ( .A1(n3762), .A2(n3076), .ZN(n3075) );
  INV_X1 U3940 ( .A(n3078), .ZN(n3077) );
  NAND2_X1 U3941 ( .A1(n3762), .A2(n6603), .ZN(n3340) );
  INV_X1 U3942 ( .A(n3343), .ZN(n3079) );
  NAND2_X1 U3943 ( .A1(n3080), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3315) );
  NAND2_X1 U3944 ( .A1(n3080), .A2(n3242), .ZN(n3249) );
  NOR2_X2 U3945 ( .A1(n3081), .A2(n3624), .ZN(n3587) );
  OAI22_X1 U3946 ( .A1(n3256), .A2(n3081), .B1(n3729), .B2(n3227), .ZN(n3257)
         );
  AOI21_X1 U3947 ( .B1(n2983), .B2(n3081), .A(n3625), .ZN(n3626) );
  NAND2_X1 U3948 ( .A1(n5378), .A2(n5380), .ZN(n5367) );
  NAND2_X1 U3949 ( .A1(n3386), .A2(n3387), .ZN(n3417) );
  NAND2_X1 U3950 ( .A1(n6108), .A2(n6107), .ZN(n6106) );
  NAND2_X1 U3951 ( .A1(n3339), .A2(n3338), .ZN(n4479) );
  AOI21_X1 U3952 ( .B1(n5500), .B2(n5586), .A(n4291), .ZN(n3536) );
  AOI21_X1 U3953 ( .B1(n5587), .B2(n5516), .A(n5500), .ZN(n5501) );
  NAND2_X1 U3954 ( .A1(n5567), .A2(n5537), .ZN(n5561) );
  AOI22_X1 U3955 ( .A1(n3204), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3184) );
  XNOR2_X1 U3956 ( .A(n3333), .B(n3377), .ZN(n3752) );
  XNOR2_X1 U3957 ( .A(n3379), .B(n3378), .ZN(n3333) );
  CLKBUF_X1 U3958 ( .A(n4584), .Z(n4670) );
  OAI21_X1 U3959 ( .B1(n4429), .B2(n3561), .A(n3395), .ZN(n3396) );
  XNOR2_X1 U3960 ( .A(n3536), .B(n3535), .ZN(n5329) );
  AND2_X1 U3961 ( .A1(n4441), .A2(n4332), .ZN(n4333) );
  AND2_X2 U3962 ( .A1(n4441), .A2(n3227), .ZN(n4418) );
  AND2_X1 U3963 ( .A1(n3608), .A2(n4441), .ZN(n3617) );
  NAND2_X1 U3964 ( .A1(n3238), .A2(n4608), .ZN(n3254) );
  NOR2_X2 U3965 ( .A1(n5287), .A2(n5313), .ZN(n5312) );
  NAND2_X2 U3966 ( .A1(n3416), .A2(n3415), .ZN(n3468) );
  CLKBUF_X1 U3967 ( .A(n2969), .Z(n4165) );
  INV_X1 U3968 ( .A(n3167), .ZN(n4608) );
  INV_X1 U3969 ( .A(n3417), .ZN(n3416) );
  AOI21_X1 U3970 ( .B1(n5327), .B2(n6133), .A(n5326), .ZN(n5328) );
  NOR2_X2 U3971 ( .A1(n5561), .A2(n5562), .ZN(n5560) );
  AND2_X1 U3972 ( .A1(n3753), .A2(n4275), .ZN(n3310) );
  NAND2_X1 U3973 ( .A1(n5997), .A2(n4275), .ZN(n5480) );
  INV_X1 U3974 ( .A(n5480), .ZN(n4286) );
  INV_X1 U3975 ( .A(n4202), .ZN(n4251) );
  INV_X1 U3976 ( .A(n4251), .ZN(n4339) );
  OR2_X1 U3977 ( .A1(n4308), .A2(n4441), .ZN(n3092) );
  INV_X1 U3978 ( .A(n3250), .ZN(n3585) );
  INV_X1 U3979 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3806) );
  NOR2_X2 U3980 ( .A1(n3753), .A2(n6601), .ZN(n3936) );
  INV_X1 U3981 ( .A(n6137), .ZN(n4310) );
  INV_X1 U3982 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3771) );
  AND2_X1 U3983 ( .A1(n4280), .A2(n4279), .ZN(n3094) );
  NAND2_X1 U3984 ( .A1(n4384), .A2(n6603), .ZN(n3095) );
  NAND2_X1 U3985 ( .A1(n3438), .A2(n3437), .ZN(n3096) );
  AND2_X1 U3986 ( .A1(n3096), .A2(n3469), .ZN(n3097) );
  AND4_X1 U3987 ( .A1(n5608), .A2(n4300), .A3(INSTADDRPOINTER_REG_30__SCAN_IN), 
        .A4(n5349), .ZN(n3098) );
  NOR2_X1 U3988 ( .A1(n5684), .A2(n3639), .ZN(n5686) );
  INV_X1 U3989 ( .A(n3396), .ZN(n6129) );
  NAND2_X1 U3990 ( .A1(n2993), .A2(n3239), .ZN(n3256) );
  OR2_X1 U3991 ( .A1(n3244), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3243)
         );
  INV_X1 U3992 ( .A(n3364), .ZN(n4189) );
  INV_X1 U3993 ( .A(n3391), .ZN(n3419) );
  INV_X1 U3994 ( .A(n3394), .ZN(n3395) );
  AND2_X1 U3995 ( .A1(n6356), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3540)
         );
  OR2_X1 U3996 ( .A1(n3247), .A2(n3246), .ZN(n3248) );
  NAND2_X1 U3997 ( .A1(n3327), .A2(n3326), .ZN(n3356) );
  NAND2_X1 U3998 ( .A1(n3204), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3132) );
  AOI22_X1 U3999 ( .A1(n4164), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3147) );
  INV_X1 U4000 ( .A(n5485), .ZN(n4010) );
  OR2_X1 U4001 ( .A1(n3479), .A2(n3478), .ZN(n3500) );
  INV_X1 U4002 ( .A(n3356), .ZN(n3328) );
  OAI21_X1 U4003 ( .B1(n3236), .B2(n3091), .A(n3633), .ZN(n3234) );
  OR2_X1 U4004 ( .A1(n3575), .A2(n3574), .ZN(n3577) );
  INV_X1 U4005 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4521) );
  NOR2_X1 U4006 ( .A1(n4223), .A2(n5513), .ZN(n4224) );
  INV_X1 U4007 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3919) );
  AND2_X1 U4008 ( .A1(n3684), .A2(n3683), .ZN(n5054) );
  INV_X1 U4009 ( .A(n3729), .ZN(n3724) );
  NAND2_X1 U4010 ( .A1(n4224), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4322)
         );
  OR2_X1 U4011 ( .A1(n4185), .A2(n4184), .ZN(n5518) );
  NAND2_X1 U4012 ( .A1(n3856), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3857)
         );
  OR3_X1 U4013 ( .A1(n4408), .A2(n4407), .A3(n4406), .ZN(n4534) );
  OR2_X1 U4014 ( .A1(n5707), .A2(n6602), .ZN(n4621) );
  INV_X1 U4015 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5101) );
  INV_X1 U4016 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4979) );
  AND2_X1 U4017 ( .A1(n4113), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4135)
         );
  AOI21_X1 U4018 ( .B1(n5097), .B2(n4202), .A(n3841), .ZN(n4911) );
  INV_X1 U4019 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5964) );
  INV_X1 U4020 ( .A(n6474), .ZN(n4273) );
  INV_X1 U4021 ( .A(n4289), .ZN(n5500) );
  OR2_X1 U4022 ( .A1(n5539), .A2(n5299), .ZN(n5279) );
  AND2_X1 U4023 ( .A1(n3742), .A2(n3636), .ZN(n5255) );
  NAND2_X1 U4024 ( .A1(n3742), .A2(n3741), .ZN(n6213) );
  INV_X1 U4025 ( .A(n4534), .ZN(n6436) );
  OR2_X1 U4026 ( .A1(n4931), .A2(n4676), .ZN(n4964) );
  OR2_X1 U4027 ( .A1(n6260), .A2(n4731), .ZN(n6234) );
  INV_X1 U4028 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4863) );
  OR2_X1 U4029 ( .A1(n5707), .A2(n4494), .ZN(n4731) );
  INV_X1 U4030 ( .A(n3618), .ZN(n4373) );
  OR2_X1 U4031 ( .A1(n4265), .A2(n6603), .ZN(n6474) );
  INV_X1 U4032 ( .A(n5742), .ZN(n5393) );
  AND2_X1 U4033 ( .A1(n5015), .A2(n4344), .ZN(n5968) );
  AND2_X1 U4034 ( .A1(n5200), .A2(n3755), .ZN(n4329) );
  AND2_X1 U4035 ( .A1(n5200), .A2(n4277), .ZN(n6005) );
  INV_X1 U4036 ( .A(n5200), .ZN(n6008) );
  INV_X1 U4037 ( .A(n6600), .ZN(n6030) );
  INV_X1 U4038 ( .A(n6104), .ZN(n6094) );
  AND2_X1 U4039 ( .A1(n2988), .A2(n5436), .ZN(n5797) );
  NAND2_X1 U4040 ( .A1(n3808), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3827)
         );
  INV_X1 U4041 ( .A(n6139), .ZN(n5821) );
  NAND2_X1 U4042 ( .A1(n3781), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3790)
         );
  INV_X1 U4043 ( .A(n5824), .ZN(n6142) );
  INV_X1 U4044 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3535) );
  OR2_X1 U4045 ( .A1(n5634), .A2(n3649), .ZN(n5826) );
  NAND2_X1 U4046 ( .A1(n3742), .A2(n4375), .ZN(n6209) );
  AND2_X1 U4047 ( .A1(n3352), .A2(n3353), .ZN(n4480) );
  NAND2_X1 U4048 ( .A1(n6603), .A2(n4430), .ZN(n4683) );
  INV_X1 U4049 ( .A(n4964), .ZN(n4660) );
  INV_X1 U4050 ( .A(n6234), .ZN(n6254) );
  INV_X1 U4051 ( .A(n6300), .ZN(n6330) );
  INV_X1 U4052 ( .A(n4719), .ZN(n6328) );
  INV_X1 U4053 ( .A(n4772), .ZN(n4812) );
  AND2_X1 U4054 ( .A1(n5707), .A2(n5028), .ZN(n4932) );
  INV_X1 U4055 ( .A(n6777), .ZN(n6408) );
  INV_X1 U4056 ( .A(n6424), .ZN(n6782) );
  INV_X1 U4057 ( .A(n5967), .ZN(n5981) );
  NAND4_X1 U4058 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_12__SCAN_IN), .A4(n5925), .ZN(n5918) );
  NAND2_X1 U4059 ( .A1(n5015), .A2(n4342), .ZN(n5946) );
  INV_X1 U4060 ( .A(n5987), .ZN(n5963) );
  NAND2_X1 U4061 ( .A1(n6097), .A2(n4274), .ZN(n5200) );
  OR2_X1 U4062 ( .A1(n6043), .A2(n6463), .ZN(n6104) );
  NAND2_X1 U4063 ( .A1(n6137), .A2(n4319), .ZN(n5824) );
  NAND2_X1 U4064 ( .A1(n5824), .A2(n4388), .ZN(n6139) );
  NOR2_X1 U4065 ( .A1(n3743), .A2(n5656), .ZN(n6151) );
  NAND2_X1 U4066 ( .A1(n3742), .A2(n3623), .ZN(n6198) );
  INV_X1 U4067 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6459) );
  NAND2_X1 U4068 ( .A1(n4866), .A2(n5028), .ZN(n5051) );
  OR2_X1 U4069 ( .A1(n6261), .A2(n6260), .ZN(n6300) );
  NOR2_X1 U4070 ( .A1(n4686), .A2(n4685), .ZN(n4724) );
  NAND2_X1 U4071 ( .A1(n4628), .A2(n4620), .ZN(n4708) );
  INV_X1 U4072 ( .A(n4779), .ZN(n4818) );
  NAND2_X1 U4073 ( .A1(n4628), .A2(n4932), .ZN(n6354) );
  INV_X1 U4074 ( .A(n6359), .ZN(n6416) );
  INV_X1 U4075 ( .A(n6286), .ZN(n6401) );
  OR2_X1 U4076 ( .A1(n6261), .A2(n4822), .ZN(n6424) );
  INV_X1 U4077 ( .A(n6564), .ZN(n6560) );
  INV_X1 U4078 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6708) );
  OAI21_X1 U4079 ( .B1(n5329), .B2(n6198), .A(n3751), .ZN(U2988) );
  AND2_X2 U4080 ( .A1(n3538), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3110)
         );
  NAND2_X1 U4081 ( .A1(n4101), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3103)
         );
  INV_X1 U4082 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3099) );
  NAND2_X1 U4083 ( .A1(n3292), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3102) );
  NAND2_X1 U4084 ( .A1(n2979), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3101)
         );
  NAND2_X1 U4085 ( .A1(n3204), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3100) );
  INV_X1 U4086 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3104) );
  NAND2_X1 U4087 ( .A1(n3213), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3109) );
  NAND2_X1 U4088 ( .A1(n4143), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3108) );
  NAND2_X1 U4089 ( .A1(n4070), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3107) );
  AND2_X2 U4090 ( .A1(n4511), .A2(n3105), .ZN(n3895) );
  NAND2_X1 U4091 ( .A1(n3895), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3106) );
  AND2_X2 U4092 ( .A1(n3110), .A2(n3115), .ZN(n3293) );
  NAND2_X1 U4093 ( .A1(n2970), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3114)
         );
  NAND2_X1 U4094 ( .A1(n4164), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3113) );
  NAND2_X1 U4095 ( .A1(n3273), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3112) );
  NAND2_X1 U4096 ( .A1(n3194), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3111) );
  AND2_X2 U4097 ( .A1(n3115), .A2(n4512), .ZN(n3266) );
  NAND2_X1 U4098 ( .A1(n3266), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3120)
         );
  AND2_X4 U4099 ( .A1(n3116), .A2(n4504), .ZN(n3218) );
  NAND2_X1 U4100 ( .A1(n3218), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3119)
         );
  NAND2_X1 U4101 ( .A1(n3199), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3118) );
  NAND2_X1 U4102 ( .A1(n3178), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3117)
         );
  NAND4_X2 U4103 ( .A1(n3124), .A2(n3123), .A3(n3122), .A4(n3121), .ZN(n3253)
         );
  NAND2_X1 U4104 ( .A1(n4143), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3128) );
  NAND2_X1 U4105 ( .A1(n3194), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3127) );
  NAND2_X1 U4106 ( .A1(n3218), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3126)
         );
  NAND2_X1 U4107 ( .A1(n3199), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3125) );
  NAND2_X1 U4108 ( .A1(n4164), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3131) );
  NAND2_X1 U4109 ( .A1(n3266), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3130)
         );
  NAND2_X1 U4110 ( .A1(n3183), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3129)
         );
  NAND2_X1 U4111 ( .A1(n3213), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3136) );
  NAND2_X1 U4112 ( .A1(n4070), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3135) );
  NAND2_X1 U4113 ( .A1(n3895), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3134) );
  NAND2_X1 U4114 ( .A1(n3178), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3133)
         );
  NAND2_X1 U4115 ( .A1(n3273), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3139) );
  NAND2_X1 U4116 ( .A1(n3292), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3138) );
  NAND2_X1 U4117 ( .A1(n2970), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3137)
         );
  NAND4_X4 U4118 ( .A1(n3144), .A2(n3143), .A3(n3142), .A4(n3141), .ZN(n3238)
         );
  AOI22_X1 U4119 ( .A1(n4101), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3292), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3148) );
  AOI22_X1 U4120 ( .A1(n2969), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3146) );
  AOI22_X1 U4121 ( .A1(n3204), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3145) );
  AOI22_X1 U4122 ( .A1(n3266), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3153) );
  NAND2_X1 U4123 ( .A1(n3178), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3150)
         );
  NAND2_X1 U4124 ( .A1(n3218), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3149)
         );
  AOI22_X1 U4125 ( .A1(n4070), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3151) );
  AOI22_X1 U4126 ( .A1(n3266), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3160) );
  AOI22_X1 U4127 ( .A1(n4143), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3159) );
  AOI22_X1 U4128 ( .A1(n3218), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3178), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3158) );
  AOI22_X1 U4129 ( .A1(n4070), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3157) );
  AOI22_X1 U4130 ( .A1(n4101), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3292), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3164) );
  AOI22_X1 U4131 ( .A1(n4164), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3163) );
  AOI22_X1 U4132 ( .A1(n2969), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3162) );
  AOI22_X1 U4133 ( .A1(n3204), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3161) );
  NAND2_X2 U4134 ( .A1(n3166), .A2(n3165), .ZN(n4275) );
  INV_X1 U4135 ( .A(n3238), .ZN(n3229) );
  AOI22_X1 U4136 ( .A1(n4101), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3171) );
  AOI22_X1 U4137 ( .A1(n4070), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3170) );
  AOI22_X1 U4138 ( .A1(n2970), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3178), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3169) );
  AOI22_X1 U4139 ( .A1(n4164), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3168) );
  NAND4_X1 U4140 ( .A1(n3171), .A2(n3170), .A3(n3169), .A4(n3168), .ZN(n3177)
         );
  AOI22_X1 U4141 ( .A1(n3194), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3175) );
  AOI22_X1 U4142 ( .A1(n3273), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3174) );
  AOI22_X1 U4143 ( .A1(n3292), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3173) );
  AOI22_X1 U4144 ( .A1(n3266), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3218), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3172) );
  NAND4_X1 U4145 ( .A1(n3175), .A2(n3174), .A3(n3173), .A4(n3172), .ZN(n3176)
         );
  AOI22_X1 U4146 ( .A1(n4143), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3182) );
  AOI22_X1 U4147 ( .A1(n3266), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3181) );
  AOI22_X1 U4148 ( .A1(n3218), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3178), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3180) );
  AOI22_X1 U4149 ( .A1(n4070), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3179) );
  NAND4_X1 U4150 ( .A1(n3182), .A2(n3181), .A3(n3180), .A4(n3179), .ZN(n3189)
         );
  AOI22_X1 U4151 ( .A1(n4101), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3292), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3187) );
  AOI22_X1 U4152 ( .A1(n4164), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3186) );
  AOI22_X1 U4153 ( .A1(n2970), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3185) );
  NAND4_X1 U4154 ( .A1(n3187), .A2(n3186), .A3(n3185), .A4(n3184), .ZN(n3188)
         );
  OR2_X2 U4155 ( .A1(n3189), .A2(n3188), .ZN(n3346) );
  NAND2_X1 U4156 ( .A1(n3213), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3193) );
  NAND2_X1 U4157 ( .A1(n4143), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3192) );
  NAND2_X1 U4158 ( .A1(n4070), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3191) );
  NAND2_X1 U4159 ( .A1(n3895), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3190) );
  NAND2_X1 U4160 ( .A1(n2970), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3198)
         );
  NAND2_X1 U4161 ( .A1(n4164), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3197) );
  NAND2_X1 U4162 ( .A1(n3273), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3196) );
  NAND2_X1 U4163 ( .A1(n3194), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3195) );
  NAND2_X1 U4164 ( .A1(n3266), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3203)
         );
  NAND2_X1 U4165 ( .A1(n3218), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3202)
         );
  NAND2_X1 U4166 ( .A1(n3199), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3201) );
  NAND2_X1 U4167 ( .A1(n3178), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3200)
         );
  NAND2_X1 U4168 ( .A1(n3292), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3208) );
  NAND2_X1 U4169 ( .A1(n4101), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3207)
         );
  NAND2_X1 U4170 ( .A1(n3183), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3206)
         );
  NAND2_X1 U4171 ( .A1(n3204), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3205) );
  NAND2_X1 U4172 ( .A1(n3273), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3217) );
  NAND2_X1 U4173 ( .A1(n4143), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3216) );
  NAND2_X1 U4174 ( .A1(n4101), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3215)
         );
  NAND2_X1 U4175 ( .A1(n3213), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3214) );
  NAND2_X1 U4176 ( .A1(n3266), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3222)
         );
  NAND2_X1 U4177 ( .A1(n4070), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3221) );
  NAND2_X1 U4178 ( .A1(n3218), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3220)
         );
  NAND2_X1 U4179 ( .A1(n3895), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3219) );
  NAND2_X1 U4180 ( .A1(n3293), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3224)
         );
  NAND2_X1 U4181 ( .A1(n4164), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3223) );
  NAND2_X1 U4182 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6499) );
  OAI21_X1 U4183 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6499), .ZN(n3596) );
  NAND2_X1 U4184 ( .A1(n3054), .A2(n3596), .ZN(n3311) );
  BUF_X1 U4185 ( .A(n3229), .Z(n4575) );
  NAND2_X1 U4186 ( .A1(n3311), .A2(n4575), .ZN(n3228) );
  AOI22_X1 U4187 ( .A1(n3310), .A2(n3230), .B1(n3633), .B2(n4275), .ZN(n3231)
         );
  NAND2_X1 U4188 ( .A1(n3250), .A2(n3231), .ZN(n3235) );
  NAND2_X1 U4189 ( .A1(n3254), .A2(n3346), .ZN(n3233) );
  NAND3_X1 U4190 ( .A1(n3235), .A2(n3234), .A3(n3233), .ZN(n3312) );
  INV_X1 U4191 ( .A(n3236), .ZN(n3237) );
  INV_X1 U4192 ( .A(n4275), .ZN(n3755) );
  NAND2_X1 U4193 ( .A1(n3237), .A2(n4275), .ZN(n3589) );
  NAND2_X1 U4194 ( .A1(n3589), .A2(n3334), .ZN(n3240) );
  NAND2_X1 U4195 ( .A1(n3239), .A2(n3619), .ZN(n4508) );
  NAND2_X1 U4196 ( .A1(n6634), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4265) );
  NAND2_X1 U4197 ( .A1(n6634), .A2(n6718), .ZN(n6586) );
  MUX2_X1 U4198 ( .A(n4265), .B(n3399), .S(n6356), .Z(n3244) );
  AND2_X1 U4199 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n3243), .ZN(n3242) );
  INV_X1 U4200 ( .A(n3243), .ZN(n3247) );
  NAND2_X1 U4201 ( .A1(n2992), .A2(n3254), .ZN(n3314) );
  INV_X1 U4202 ( .A(n3244), .ZN(n3245) );
  AND2_X1 U4203 ( .A1(n3314), .A2(n3245), .ZN(n3246) );
  INV_X1 U4204 ( .A(n3254), .ZN(n3590) );
  OR2_X1 U4205 ( .A1(n6586), .A2(n6603), .ZN(n6475) );
  AOI21_X1 U4206 ( .B1(n3590), .B2(n2984), .A(n6475), .ZN(n3252) );
  NAND2_X1 U4208 ( .A1(n3585), .A2(n3309), .ZN(n3251) );
  AND2_X1 U4209 ( .A1(n3252), .A2(n3251), .ZN(n3259) );
  INV_X1 U4210 ( .A(n5003), .ZN(n4371) );
  AOI22_X1 U4211 ( .A1(n4371), .A2(n4308), .B1(n4441), .B2(n3633), .ZN(n3260)
         );
  XNOR2_X2 U4212 ( .A(n3327), .B(n3261), .ZN(n3762) );
  AOI22_X1 U4213 ( .A1(n4238), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4229), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3265) );
  AOI22_X1 U4214 ( .A1(n4231), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3264) );
  AOI22_X1 U4215 ( .A1(n2968), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3263) );
  AOI22_X1 U4216 ( .A1(n2970), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4240), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3262) );
  NAND4_X1 U4217 ( .A1(n3265), .A2(n3264), .A3(n3263), .A4(n3262), .ZN(n3272)
         );
  AOI22_X1 U4218 ( .A1(n3213), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4228), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3270) );
  INV_X1 U4219 ( .A(n3364), .ZN(n3278) );
  AOI22_X1 U4220 ( .A1(n3278), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3269) );
  AOI22_X1 U4222 ( .A1(n4069), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3268) );
  AOI22_X1 U4223 ( .A1(n4237), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3267) );
  NAND4_X1 U4224 ( .A1(n3270), .A2(n3269), .A3(n3268), .A4(n3267), .ZN(n3271)
         );
  NOR2_X1 U4225 ( .A1(n4266), .A2(n3511), .ZN(n3304) );
  NAND2_X1 U4226 ( .A1(n4559), .A2(n3511), .ZN(n3288) );
  AOI22_X1 U4227 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n4238), .B1(n4237), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3277) );
  AOI22_X1 U4228 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n2969), .B1(n2980), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3276) );
  AOI22_X1 U4229 ( .A1(n4229), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3275) );
  AOI22_X1 U4230 ( .A1(n3218), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3274) );
  NAND4_X1 U4231 ( .A1(n3277), .A2(n3276), .A3(n3275), .A4(n3274), .ZN(n3284)
         );
  AOI22_X1 U4232 ( .A1(n3278), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3282) );
  AOI22_X1 U4233 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n3213), .B1(n4240), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3281) );
  AOI22_X1 U4234 ( .A1(n4069), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3280) );
  AOI22_X1 U4235 ( .A1(n4231), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3279) );
  NAND4_X1 U4236 ( .A1(n3282), .A2(n3281), .A3(n3280), .A4(n3279), .ZN(n3283)
         );
  INV_X1 U4237 ( .A(n3390), .ZN(n3285) );
  MUX2_X1 U4238 ( .A(n3304), .B(n3291), .S(n3285), .Z(n3286) );
  INV_X1 U4239 ( .A(n3570), .ZN(n3555) );
  INV_X1 U4240 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3290) );
  AOI21_X1 U4241 ( .B1(n4474), .B2(n3390), .A(n6603), .ZN(n3289) );
  OAI211_X1 U4242 ( .C1(n3555), .C2(n3290), .A(n3289), .B(n3288), .ZN(n3343)
         );
  INV_X1 U4243 ( .A(n3291), .ZN(n3507) );
  AOI22_X1 U4244 ( .A1(n4231), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3297) );
  INV_X1 U4245 ( .A(n3292), .ZN(n3364) );
  AOI22_X1 U4246 ( .A1(n4189), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4247 ( .A1(n2970), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3295) );
  AOI22_X1 U4248 ( .A1(n3218), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3294) );
  NAND4_X1 U4249 ( .A1(n3297), .A2(n3296), .A3(n3295), .A4(n3294), .ZN(n3303)
         );
  AOI22_X1 U4250 ( .A1(n2980), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4251 ( .A1(n4229), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4252 ( .A1(n4238), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4240), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3299) );
  BUF_X2 U4253 ( .A(n3266), .Z(n4069) );
  AOI22_X1 U4254 ( .A1(n4069), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3298) );
  NAND4_X1 U4255 ( .A1(n3301), .A2(n3300), .A3(n3299), .A4(n3298), .ZN(n3302)
         );
  INV_X1 U4256 ( .A(n3389), .ZN(n3307) );
  INV_X1 U4257 ( .A(n3304), .ZN(n3306) );
  NAND2_X1 U4258 ( .A1(n3570), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3305) );
  OAI211_X1 U4259 ( .C1(n3307), .C2(n3402), .A(n3306), .B(n3305), .ZN(n3378)
         );
  NAND2_X1 U4260 ( .A1(n3335), .A2(n4575), .ZN(n3308) );
  NAND3_X1 U4261 ( .A1(n3309), .A2(n3611), .A3(n4575), .ZN(n4268) );
  AOI21_X1 U4262 ( .B1(n3617), .B2(n3311), .A(n3621), .ZN(n3313) );
  NAND2_X1 U4263 ( .A1(n3313), .A2(n3616), .ZN(n3324) );
  NAND2_X1 U4264 ( .A1(n3324), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3320) );
  NAND2_X1 U4265 ( .A1(n3315), .A2(n3314), .ZN(n3359) );
  NAND2_X1 U4266 ( .A1(n3359), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3319) );
  XNOR2_X1 U4267 ( .A(n4863), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5144)
         );
  NAND2_X1 U4268 ( .A1(n3399), .A2(n5144), .ZN(n3317) );
  NAND2_X1 U4269 ( .A1(n4265), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3316) );
  NAND2_X1 U4270 ( .A1(n3317), .A2(n3316), .ZN(n3321) );
  INV_X1 U4271 ( .A(n3321), .ZN(n3318) );
  NAND3_X1 U4272 ( .A1(n3320), .A2(n3319), .A3(n3318), .ZN(n3357) );
  OR2_X1 U4273 ( .A1(n3321), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3322)
         );
  AND2_X1 U4274 ( .A1(n3322), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3323) );
  NAND2_X1 U4275 ( .A1(n3324), .A2(n3323), .ZN(n3355) );
  NAND2_X1 U4276 ( .A1(n3357), .A2(n3355), .ZN(n3329) );
  NAND2_X1 U4277 ( .A1(n3630), .A2(n3325), .ZN(n3326) );
  NAND2_X1 U4278 ( .A1(n4427), .A2(n6603), .ZN(n3332) );
  INV_X1 U4279 ( .A(n4266), .ZN(n3330) );
  NAND2_X1 U4280 ( .A1(n3330), .A2(n3389), .ZN(n3331) );
  NAND2_X1 U4281 ( .A1(n3752), .A2(n3547), .ZN(n3339) );
  XNOR2_X1 U4282 ( .A(n3390), .B(n3389), .ZN(n3336) );
  INV_X1 U4283 ( .A(n2984), .ZN(n3591) );
  OAI211_X1 U4284 ( .C1(n3336), .C2(n3591), .A(n3335), .B(n3238), .ZN(n3337)
         );
  INV_X1 U4285 ( .A(n3337), .ZN(n3338) );
  NAND2_X1 U4286 ( .A1(n3340), .A2(n3343), .ZN(n3341) );
  NAND2_X1 U4287 ( .A1(n3341), .A2(n3342), .ZN(n3345) );
  NAND2_X1 U4288 ( .A1(n3286), .A2(n3343), .ZN(n3344) );
  AND2_X2 U4289 ( .A1(n3345), .A2(n3344), .ZN(n4494) );
  NAND2_X1 U4290 ( .A1(n4494), .A2(n3547), .ZN(n3349) );
  NAND2_X1 U4291 ( .A1(n4474), .A2(n3346), .ZN(n3392) );
  OAI21_X1 U4292 ( .B1(n3591), .B2(n3390), .A(n3392), .ZN(n3347) );
  INV_X1 U4293 ( .A(n3347), .ZN(n3348) );
  NAND2_X1 U4294 ( .A1(n3349), .A2(n3348), .ZN(n4387) );
  NAND2_X1 U4295 ( .A1(n4387), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3350)
         );
  INV_X1 U4296 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U4297 ( .A1(n3350), .A2(n6215), .ZN(n3352) );
  AND2_X1 U4298 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3351) );
  NAND2_X1 U4299 ( .A1(n4387), .A2(n3351), .ZN(n3353) );
  NAND2_X1 U4300 ( .A1(n4479), .A2(n4480), .ZN(n3354) );
  NAND2_X1 U4301 ( .A1(n3354), .A2(n3353), .ZN(n6131) );
  NAND2_X1 U4302 ( .A1(n3356), .A2(n3355), .ZN(n3358) );
  NAND2_X1 U4303 ( .A1(n3359), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3363) );
  NAND2_X1 U4304 ( .A1(n6442), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4919) );
  MUX2_X1 U4305 ( .A(n4919), .B(n6442), .S(n6356), .Z(n3361) );
  AND2_X1 U4306 ( .A1(n4863), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4730)
         );
  INV_X1 U4307 ( .A(n4730), .ZN(n3360) );
  NAND2_X1 U4308 ( .A1(n3361), .A2(n3360), .ZN(n4488) );
  AOI22_X1 U4309 ( .A1(n4488), .A2(n3399), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n4265), .ZN(n3362) );
  AOI22_X1 U4310 ( .A1(n2980), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4189), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4311 ( .A1(n4231), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4312 ( .A1(n4165), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4313 ( .A1(n4240), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3365) );
  NAND4_X1 U4314 ( .A1(n3368), .A2(n3367), .A3(n3366), .A4(n3365), .ZN(n3374)
         );
  AOI22_X1 U4315 ( .A1(n4238), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4316 ( .A1(n4069), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3371) );
  AOI22_X1 U4317 ( .A1(n3218), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4318 ( .A1(n4229), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3369) );
  NAND4_X1 U4319 ( .A1(n3372), .A2(n3371), .A3(n3370), .A4(n3369), .ZN(n3373)
         );
  INV_X1 U4320 ( .A(n3402), .ZN(n3375) );
  AOI22_X1 U4321 ( .A1(n3570), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3375), 
        .B2(n3391), .ZN(n3384) );
  INV_X1 U4322 ( .A(n3384), .ZN(n3376) );
  XNOR2_X1 U4323 ( .A(n3385), .B(n3376), .ZN(n3382) );
  NAND2_X1 U4324 ( .A1(n3379), .A2(n3378), .ZN(n3380) );
  INV_X1 U4325 ( .A(n3383), .ZN(n3387) );
  XNOR2_X1 U4326 ( .A(n3385), .B(n3384), .ZN(n3386) );
  NAND2_X1 U4327 ( .A1(n3390), .A2(n3389), .ZN(n3420) );
  XNOR2_X1 U4328 ( .A(n3420), .B(n3391), .ZN(n3393) );
  OAI21_X1 U4329 ( .B1(n3393), .B2(n3591), .A(n3392), .ZN(n3394) );
  NAND2_X1 U4330 ( .A1(n3359), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3401) );
  NOR3_X1 U4331 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6442), .A3(n4863), 
        .ZN(n6313) );
  NAND2_X1 U4332 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6313), .ZN(n6306) );
  NAND2_X1 U4333 ( .A1(n6446), .A2(n6306), .ZN(n3398) );
  NOR3_X1 U4334 ( .A1(n6446), .A2(n6442), .A3(n4863), .ZN(n4436) );
  NAND2_X1 U4335 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4436), .ZN(n4726) );
  AOI22_X1 U4336 ( .A1(n3399), .A2(n4681), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n4265), .ZN(n3400) );
  NAND2_X1 U4337 ( .A1(n4424), .A2(n6603), .ZN(n3414) );
  AOI22_X1 U4338 ( .A1(n4237), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n2980), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3406) );
  AOI22_X1 U4339 ( .A1(n4165), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3405) );
  INV_X1 U4340 ( .A(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n6617) );
  AOI22_X1 U4341 ( .A1(n4231), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3404) );
  BUF_X2 U4342 ( .A(n3218), .Z(n4228) );
  AOI22_X1 U4343 ( .A1(n4228), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3403) );
  NAND4_X1 U4344 ( .A1(n3406), .A2(n3405), .A3(n3404), .A4(n3403), .ZN(n3412)
         );
  AOI22_X1 U4345 ( .A1(n4238), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4229), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3410) );
  AOI22_X1 U4346 ( .A1(n4069), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3409) );
  AOI22_X1 U4347 ( .A1(n4189), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3408) );
  AOI22_X1 U4348 ( .A1(n4240), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3407) );
  NAND4_X1 U4349 ( .A1(n3410), .A2(n3409), .A3(n3408), .A4(n3407), .ZN(n3411)
         );
  AOI22_X1 U4350 ( .A1(n3578), .A2(n3439), .B1(n3570), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3413) );
  INV_X1 U4351 ( .A(n4489), .ZN(n3415) );
  NAND2_X1 U4352 ( .A1(n3417), .A2(n4489), .ZN(n3418) );
  NAND2_X1 U4353 ( .A1(n3420), .A2(n3419), .ZN(n3440) );
  INV_X1 U4354 ( .A(n3439), .ZN(n3421) );
  XNOR2_X1 U4355 ( .A(n3440), .B(n3421), .ZN(n3422) );
  NAND2_X1 U4356 ( .A1(n3422), .A2(n2984), .ZN(n3423) );
  INV_X1 U4357 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3424) );
  NAND2_X1 U4358 ( .A1(n3425), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3426)
         );
  AOI22_X1 U4359 ( .A1(n4237), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4360 ( .A1(n4188), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4228), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4361 ( .A1(n4165), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4362 ( .A1(n2980), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4240), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3427) );
  NAND4_X1 U4363 ( .A1(n3430), .A2(n3429), .A3(n3428), .A4(n3427), .ZN(n3436)
         );
  AOI22_X1 U4364 ( .A1(n4231), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4189), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3434) );
  AOI22_X1 U4365 ( .A1(n4069), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3433) );
  AOI22_X1 U4366 ( .A1(n4238), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3432) );
  AOI22_X1 U4367 ( .A1(n4239), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3431) );
  NAND4_X1 U4368 ( .A1(n3434), .A2(n3433), .A3(n3432), .A4(n3431), .ZN(n3435)
         );
  NAND2_X1 U4369 ( .A1(n3578), .A2(n3487), .ZN(n3438) );
  NAND2_X1 U4370 ( .A1(n3570), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3437) );
  XNOR2_X1 U4371 ( .A(n3468), .B(n3096), .ZN(n3786) );
  NAND2_X1 U4372 ( .A1(n3786), .A2(n3547), .ZN(n3443) );
  NAND2_X1 U4373 ( .A1(n3440), .A2(n3439), .ZN(n3489) );
  XNOR2_X1 U4374 ( .A(n3489), .B(n3487), .ZN(n3441) );
  NAND2_X1 U4375 ( .A1(n3441), .A2(n2984), .ZN(n3442) );
  NAND2_X1 U4376 ( .A1(n3443), .A2(n3442), .ZN(n3445) );
  INV_X1 U4377 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3444) );
  XNOR2_X1 U4378 ( .A(n3445), .B(n3444), .ZN(n4582) );
  NAND2_X1 U4379 ( .A1(n4583), .A2(n4582), .ZN(n4581) );
  NAND2_X1 U4380 ( .A1(n3445), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3446)
         );
  NAND2_X1 U4381 ( .A1(n4581), .A2(n3446), .ZN(n5693) );
  AOI22_X1 U4382 ( .A1(n2980), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4189), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4383 ( .A1(n4231), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4384 ( .A1(n4165), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4385 ( .A1(n4240), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3448) );
  NAND4_X1 U4386 ( .A1(n3451), .A2(n3450), .A3(n3449), .A4(n3448), .ZN(n3457)
         );
  AOI22_X1 U4387 ( .A1(n4238), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4388 ( .A1(n4069), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4389 ( .A1(n4228), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3453) );
  INV_X1 U4390 ( .A(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n6696) );
  AOI22_X1 U4391 ( .A1(n4229), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3452) );
  NAND4_X1 U4392 ( .A1(n3455), .A2(n3454), .A3(n3453), .A4(n3452), .ZN(n3456)
         );
  NAND2_X1 U4393 ( .A1(n3578), .A2(n3486), .ZN(n3459) );
  NAND2_X1 U4394 ( .A1(n3570), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3458) );
  NAND2_X1 U4395 ( .A1(n3459), .A2(n3458), .ZN(n3469) );
  NAND2_X1 U4396 ( .A1(n3799), .A2(n3547), .ZN(n3465) );
  INV_X1 U4397 ( .A(n3487), .ZN(n3461) );
  OR2_X1 U4398 ( .A1(n3489), .A2(n3461), .ZN(n3462) );
  XNOR2_X1 U4399 ( .A(n3462), .B(n3486), .ZN(n3463) );
  NAND2_X1 U4400 ( .A1(n3463), .A2(n2984), .ZN(n3464) );
  NAND2_X1 U4401 ( .A1(n3465), .A2(n3464), .ZN(n3466) );
  INV_X1 U4402 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5688) );
  XNOR2_X1 U4403 ( .A(n3466), .B(n5688), .ZN(n5692) );
  NAND2_X1 U4404 ( .A1(n5693), .A2(n5692), .ZN(n5691) );
  NAND2_X1 U4405 ( .A1(n3466), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3467)
         );
  NAND2_X1 U4406 ( .A1(n5691), .A2(n3467), .ZN(n4859) );
  AOI22_X1 U4407 ( .A1(n2980), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4189), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3473) );
  AOI22_X1 U4408 ( .A1(n4231), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3472) );
  AOI22_X1 U4409 ( .A1(n4165), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4410 ( .A1(n4240), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3470) );
  NAND4_X1 U4411 ( .A1(n3473), .A2(n3472), .A3(n3471), .A4(n3470), .ZN(n3479)
         );
  AOI22_X1 U4412 ( .A1(n4238), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3477) );
  AOI22_X1 U4413 ( .A1(n4069), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3476) );
  AOI22_X1 U4414 ( .A1(n4228), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3475) );
  AOI22_X1 U4415 ( .A1(n4229), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3474) );
  NAND4_X1 U4416 ( .A1(n3477), .A2(n3476), .A3(n3475), .A4(n3474), .ZN(n3478)
         );
  NAND2_X1 U4417 ( .A1(n3578), .A2(n3500), .ZN(n3481) );
  NAND2_X1 U4418 ( .A1(n3570), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3480) );
  NAND2_X1 U4419 ( .A1(n3485), .A2(n3484), .ZN(n3803) );
  NAND3_X1 U4420 ( .A1(n3509), .A2(n3547), .A3(n3803), .ZN(n3492) );
  NAND2_X1 U4421 ( .A1(n3487), .A2(n3486), .ZN(n3488) );
  OR2_X1 U4422 ( .A1(n3489), .A2(n3488), .ZN(n3499) );
  XNOR2_X1 U4423 ( .A(n3499), .B(n3500), .ZN(n3490) );
  NAND2_X1 U4424 ( .A1(n3490), .A2(n2984), .ZN(n3491) );
  NAND2_X1 U4425 ( .A1(n3492), .A2(n3491), .ZN(n3493) );
  INV_X1 U4426 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5120) );
  XNOR2_X1 U4427 ( .A(n3493), .B(n5120), .ZN(n4858) );
  NAND2_X1 U4428 ( .A1(n4859), .A2(n4858), .ZN(n4857) );
  NAND2_X1 U4429 ( .A1(n3493), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3494)
         );
  NAND2_X1 U4430 ( .A1(n4857), .A2(n3494), .ZN(n6108) );
  INV_X1 U4431 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3496) );
  NAND2_X1 U4432 ( .A1(n3578), .A2(n3511), .ZN(n3495) );
  OAI21_X1 U4433 ( .B1(n3496), .B2(n3555), .A(n3495), .ZN(n3497) );
  XNOR2_X1 U4434 ( .A(n3509), .B(n3497), .ZN(n3805) );
  INV_X1 U4435 ( .A(n3805), .ZN(n3498) );
  OR2_X1 U4436 ( .A1(n3498), .A2(n3561), .ZN(n3504) );
  INV_X1 U4437 ( .A(n3499), .ZN(n3501) );
  NAND2_X1 U4438 ( .A1(n3501), .A2(n3500), .ZN(n3510) );
  XNOR2_X1 U4439 ( .A(n3510), .B(n3511), .ZN(n3502) );
  NAND2_X1 U4440 ( .A1(n3502), .A2(n2984), .ZN(n3503) );
  NAND2_X1 U4441 ( .A1(n3504), .A2(n3503), .ZN(n3505) );
  INV_X1 U4442 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6175) );
  XNOR2_X1 U4443 ( .A(n3505), .B(n6175), .ZN(n6107) );
  NAND2_X1 U4444 ( .A1(n3505), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3506)
         );
  NAND2_X1 U4445 ( .A1(n6106), .A2(n3506), .ZN(n4990) );
  NOR2_X1 U4446 ( .A1(n3507), .A2(n3561), .ZN(n3508) );
  INV_X1 U4447 ( .A(n3510), .ZN(n3512) );
  NAND3_X1 U4448 ( .A1(n3512), .A2(n2984), .A3(n3511), .ZN(n3513) );
  NAND2_X1 U4449 ( .A1(n5539), .A2(n3513), .ZN(n3514) );
  INV_X1 U4450 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6169) );
  XNOR2_X1 U4451 ( .A(n3514), .B(n6169), .ZN(n4989) );
  NAND2_X1 U4452 ( .A1(n3514), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3515)
         );
  INV_X1 U4453 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5121) );
  NAND2_X1 U4454 ( .A1(n5539), .A2(n5121), .ZN(n5060) );
  OR2_X1 U4455 ( .A1(n5539), .A2(n5121), .ZN(n5061) );
  INV_X1 U4456 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3516) );
  NAND2_X1 U4457 ( .A1(n5539), .A2(n3516), .ZN(n5107) );
  INV_X1 U4458 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3517) );
  INV_X1 U4459 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5226) );
  NOR2_X1 U4460 ( .A1(n5539), .A2(n5226), .ZN(n5223) );
  NAND2_X1 U4461 ( .A1(n5539), .A2(n5226), .ZN(n5221) );
  XNOR2_X1 U4462 ( .A(n5539), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5247)
         );
  INV_X1 U4463 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3519) );
  NAND2_X1 U4464 ( .A1(n5539), .A2(n3519), .ZN(n3520) );
  INV_X1 U4465 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5299) );
  INV_X1 U4466 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5849) );
  NOR2_X1 U4467 ( .A1(n5539), .A2(n5849), .ZN(n3522) );
  NAND2_X1 U4468 ( .A1(n5539), .A2(n5849), .ZN(n3521) );
  AND2_X1 U4469 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3745) );
  NAND2_X1 U4470 ( .A1(n3745), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3523) );
  INV_X1 U4471 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5857) );
  INV_X1 U4472 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5834) );
  INV_X1 U4473 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6737) );
  AND3_X1 U4474 ( .A1(n5857), .A2(n5834), .A3(n6737), .ZN(n3524) );
  NAND2_X1 U4475 ( .A1(n5534), .A2(n3525), .ZN(n3529) );
  INV_X1 U4476 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5679) );
  NOR2_X1 U4477 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3527) );
  INV_X1 U4478 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5623) );
  INV_X1 U4479 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6633) );
  INV_X1 U4480 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3526) );
  NAND4_X1 U4481 ( .A1(n3527), .A2(n5623), .A3(n6633), .A4(n3526), .ZN(n3531)
         );
  AND2_X1 U4482 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5663) );
  AND2_X1 U4483 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3644) );
  NAND2_X1 U4484 ( .A1(n5663), .A2(n3644), .ZN(n5546) );
  NAND2_X1 U4485 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3747) );
  NOR2_X1 U4486 ( .A1(n5546), .A2(n3747), .ZN(n3528) );
  NAND2_X1 U4487 ( .A1(n3529), .A2(n3528), .ZN(n3530) );
  XNOR2_X1 U4488 ( .A(n5539), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5808)
         );
  NOR2_X1 U4489 ( .A1(n5539), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5524)
         );
  NOR2_X1 U4490 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3532) );
  INV_X1 U4491 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5586) );
  INV_X1 U4492 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6674) );
  INV_X1 U4493 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3534) );
  NOR2_X1 U4494 ( .A1(n2986), .A2(n3534), .ZN(n5525) );
  AND2_X1 U4495 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U4496 ( .A1(n5587), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3748) );
  AND2_X1 U4497 ( .A1(n3054), .A2(n3238), .ZN(n3537) );
  XNOR2_X1 U4498 ( .A(n3538), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3543)
         );
  OAI21_X1 U4499 ( .B1(n3619), .B2(n3543), .A(n4441), .ZN(n3539) );
  NAND2_X1 U4500 ( .A1(n3563), .A2(n3539), .ZN(n3545) );
  INV_X1 U4501 ( .A(n3545), .ZN(n3548) );
  XNOR2_X1 U4502 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3541) );
  NAND2_X1 U4503 ( .A1(n3540), .A2(n3541), .ZN(n3553) );
  OAI21_X1 U4504 ( .B1(n3541), .B2(n3540), .A(n3553), .ZN(n3550) );
  INV_X1 U4505 ( .A(n3550), .ZN(n3597) );
  NAND2_X1 U4506 ( .A1(n3578), .A2(n3227), .ZN(n3542) );
  NAND2_X1 U4507 ( .A1(n3542), .A2(n3238), .ZN(n3549) );
  INV_X1 U4508 ( .A(n3578), .ZN(n3544) );
  NOR2_X1 U4509 ( .A1(n3544), .A2(n3543), .ZN(n3546) );
  INV_X1 U4510 ( .A(n3549), .ZN(n3551) );
  NAND2_X1 U4511 ( .A1(n4863), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3552) );
  NAND2_X1 U4512 ( .A1(n3553), .A2(n3552), .ZN(n3558) );
  XNOR2_X1 U4513 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3557) );
  INV_X1 U4514 ( .A(n3557), .ZN(n3554) );
  XNOR2_X1 U4515 ( .A(n3558), .B(n3554), .ZN(n3598) );
  NAND2_X1 U4516 ( .A1(n3578), .A2(n3598), .ZN(n3562) );
  OAI211_X1 U4517 ( .C1(n3598), .C2(n3555), .A(n3563), .B(n3562), .ZN(n3556)
         );
  XNOR2_X1 U4518 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3566) );
  NAND2_X1 U4519 ( .A1(n3558), .A2(n3557), .ZN(n3560) );
  NAND2_X1 U4520 ( .A1(n6442), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3559) );
  NAND2_X1 U4521 ( .A1(n3560), .A2(n3559), .ZN(n3567) );
  XOR2_X1 U4522 ( .A(n3566), .B(n3567), .Z(n3599) );
  OAI22_X1 U4523 ( .A1(n3563), .A2(n3562), .B1(n3599), .B2(n3561), .ZN(n3564)
         );
  NAND2_X1 U4524 ( .A1(n3567), .A2(n3566), .ZN(n3569) );
  NAND2_X1 U4525 ( .A1(n6446), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3568) );
  NAND2_X1 U4526 ( .A1(n3569), .A2(n3568), .ZN(n3575) );
  NAND2_X1 U4527 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6613), .ZN(n3576) );
  NOR2_X1 U4528 ( .A1(n3570), .A2(n3600), .ZN(n3571) );
  OAI22_X1 U4529 ( .A1(n3572), .A2(n3571), .B1(n3582), .B2(n3600), .ZN(n3573)
         );
  AOI21_X1 U4530 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6603), .A(n3573), 
        .ZN(n3580) );
  NAND2_X1 U4531 ( .A1(n3578), .A2(n3602), .ZN(n3579) );
  NAND2_X1 U4532 ( .A1(n3580), .A2(n3579), .ZN(n3584) );
  INV_X1 U4533 ( .A(n3602), .ZN(n3581) );
  NAND2_X1 U4534 ( .A1(n3585), .A2(n3238), .ZN(n6431) );
  NOR2_X1 U4535 ( .A1(n6431), .A2(n3054), .ZN(n3637) );
  INV_X1 U4536 ( .A(n3637), .ZN(n3606) );
  INV_X1 U4537 ( .A(n3586), .ZN(n3595) );
  NAND2_X1 U4538 ( .A1(n6431), .A2(n4474), .ZN(n3588) );
  NAND2_X1 U4539 ( .A1(n3587), .A2(n3588), .ZN(n4309) );
  INV_X1 U4540 ( .A(n4309), .ZN(n3593) );
  NAND2_X1 U4541 ( .A1(n3589), .A2(n2981), .ZN(n3592) );
  MUX2_X1 U4542 ( .A(n3592), .B(n3591), .S(n3590), .Z(n3628) );
  NAND2_X1 U4543 ( .A1(n3593), .A2(n3628), .ZN(n3594) );
  NAND2_X1 U4544 ( .A1(n3595), .A2(n3594), .ZN(n4404) );
  OR2_X1 U4545 ( .A1(n3596), .A2(STATE_REG_0__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U4546 ( .A1(n3227), .A2(n6490), .ZN(n3604) );
  AND3_X1 U4547 ( .A1(n3599), .A2(n3598), .A3(n3597), .ZN(n3601) );
  OAI21_X1 U4548 ( .B1(n3602), .B2(n3601), .A(n3600), .ZN(n4376) );
  INV_X1 U4549 ( .A(READY_N), .ZN(n6491) );
  NAND2_X1 U4550 ( .A1(n4376), .A2(n6491), .ZN(n4262) );
  INV_X1 U4551 ( .A(n4262), .ZN(n3603) );
  NAND3_X1 U4552 ( .A1(n3604), .A2(n3633), .A3(n3603), .ZN(n3605) );
  OAI211_X1 U4553 ( .C1(n6468), .C2(n3606), .A(n4404), .B(n3605), .ZN(n3607)
         );
  NAND2_X1 U4554 ( .A1(n3607), .A2(n4273), .ZN(n3615) );
  NAND2_X1 U4555 ( .A1(n3054), .A2(n6490), .ZN(n4334) );
  NAND3_X1 U4556 ( .A1(n3608), .A2(n4334), .A3(n6491), .ZN(n3610) );
  INV_X1 U4557 ( .A(n4277), .ZN(n3609) );
  NAND3_X1 U4558 ( .A1(n3610), .A2(n2982), .A3(n3609), .ZN(n3612) );
  NAND2_X1 U4559 ( .A1(n3612), .A2(n3611), .ZN(n3613) );
  NAND2_X1 U4560 ( .A1(n3618), .A2(n3227), .ZN(n4400) );
  NOR2_X1 U4561 ( .A1(n3619), .A2(n5001), .ZN(n3620) );
  OR2_X1 U4562 ( .A1(n4309), .A2(n3620), .ZN(n4372) );
  NAND2_X1 U4563 ( .A1(n3621), .A2(n3253), .ZN(n3622) );
  NAND4_X1 U4564 ( .A1(n3616), .A2(n4400), .A3(n4372), .A4(n3622), .ZN(n3623)
         );
  NOR2_X1 U4565 ( .A1(n5003), .A2(n3633), .ZN(n4402) );
  OAI21_X1 U4566 ( .B1(n4402), .B2(n3654), .A(n3624), .ZN(n3627) );
  NOR2_X1 U4567 ( .A1(n4277), .A2(n3611), .ZN(n3625) );
  AND2_X1 U4568 ( .A1(n3627), .A2(n3626), .ZN(n3629) );
  NAND3_X1 U4569 ( .A1(n3630), .A2(n3629), .A3(n3628), .ZN(n4509) );
  INV_X1 U4570 ( .A(n4508), .ZN(n3631) );
  AOI22_X1 U4571 ( .A1(n4505), .A2(n3091), .B1(n3631), .B2(n4474), .ZN(n3634)
         );
  NAND2_X1 U4572 ( .A1(n3309), .A2(n4474), .ZN(n3632) );
  OR3_X1 U4573 ( .A1(n6431), .A2(n3633), .A3(n3632), .ZN(n4528) );
  NAND2_X1 U4574 ( .A1(n3634), .A2(n4528), .ZN(n3635) );
  NOR2_X1 U4575 ( .A1(n4509), .A2(n3635), .ZN(n3638) );
  INV_X1 U4576 ( .A(n3638), .ZN(n3636) );
  NAND2_X1 U4577 ( .A1(n3638), .A2(n3637), .ZN(n4518) );
  INV_X1 U4578 ( .A(n4518), .ZN(n4375) );
  INV_X1 U4579 ( .A(n6209), .ZN(n3639) );
  INV_X1 U4580 ( .A(n5686), .ZN(n5303) );
  NAND2_X1 U4581 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U4582 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6188) );
  NOR2_X1 U4583 ( .A1(n5683), .A2(n6188), .ZN(n5689) );
  NAND3_X1 U4584 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n5689), .ZN(n5117) );
  NOR2_X1 U4585 ( .A1(n6175), .A2(n6169), .ZN(n6164) );
  NAND3_X1 U4586 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6164), .ZN(n3640) );
  NOR2_X1 U4587 ( .A1(n5117), .A2(n3640), .ZN(n5254) );
  INV_X1 U4588 ( .A(n5254), .ZN(n5263) );
  NOR2_X1 U4589 ( .A1(n6364), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4384) );
  NOR2_X1 U4590 ( .A1(n3742), .A2(n2971), .ZN(n5703) );
  NOR2_X1 U4591 ( .A1(n5255), .A2(n3639), .ZN(n5260) );
  NOR2_X1 U4592 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5260), .ZN(n5698)
         );
  NOR2_X1 U4593 ( .A1(n5703), .A2(n5698), .ZN(n5681) );
  NAND2_X1 U4594 ( .A1(n6209), .A2(n5681), .ZN(n5655) );
  INV_X1 U4595 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6758) );
  NAND2_X1 U4596 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U4597 ( .A1(n6758), .A2(n6205), .ZN(n6206) );
  NAND3_X1 U4598 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n6206), .ZN(n5119) );
  NOR2_X1 U4599 ( .A1(n6209), .A2(n5119), .ZN(n5687) );
  NAND3_X1 U4600 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n5687), .ZN(n5116) );
  NOR2_X1 U4601 ( .A1(n3640), .A2(n5116), .ZN(n3743) );
  INV_X1 U4602 ( .A(n3743), .ZN(n5257) );
  AOI22_X1 U4603 ( .A1(n5684), .A2(n5263), .B1(n5655), .B2(n5257), .ZN(n6150)
         );
  NOR2_X1 U4604 ( .A1(n3517), .A2(n5226), .ZN(n5259) );
  NAND2_X1 U4605 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5259), .ZN(n5859) );
  NOR2_X1 U4606 ( .A1(n5299), .A2(n5859), .ZN(n5300) );
  NAND3_X1 U4607 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5300), .ZN(n3744) );
  NAND2_X1 U4608 ( .A1(n5303), .A2(n3744), .ZN(n3641) );
  NAND2_X1 U4609 ( .A1(n6150), .A2(n3641), .ZN(n5845) );
  NAND2_X1 U4610 ( .A1(n5663), .A2(n3745), .ZN(n3642) );
  AND2_X1 U4611 ( .A1(n5303), .A2(n3642), .ZN(n3643) );
  NOR2_X1 U4612 ( .A1(n5845), .A2(n3643), .ZN(n5643) );
  INV_X1 U4613 ( .A(n3644), .ZN(n3746) );
  NAND2_X1 U4614 ( .A1(n5303), .A2(n3746), .ZN(n3645) );
  NAND2_X1 U4615 ( .A1(n5643), .A2(n3645), .ZN(n5634) );
  INV_X1 U4616 ( .A(n5684), .ZN(n3646) );
  NOR2_X1 U4617 ( .A1(n5702), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4481)
         );
  INV_X1 U4618 ( .A(n6217), .ZN(n3647) );
  AND2_X1 U4619 ( .A1(n6209), .A2(n3647), .ZN(n5118) );
  INV_X1 U4620 ( .A(n3747), .ZN(n3648) );
  NOR2_X1 U4621 ( .A1(n5118), .A2(n3648), .ZN(n3649) );
  AND2_X1 U4622 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5619) );
  NOR2_X1 U4623 ( .A1(n5686), .A2(n5619), .ZN(n3650) );
  NOR2_X1 U4624 ( .A1(n5826), .A2(n3650), .ZN(n5595) );
  INV_X1 U4625 ( .A(n5587), .ZN(n3651) );
  NAND2_X1 U4626 ( .A1(n5303), .A2(n3651), .ZN(n3652) );
  NAND2_X1 U4627 ( .A1(n5595), .A2(n3652), .ZN(n5592) );
  AOI21_X1 U4628 ( .B1(n5586), .B2(n5303), .A(n5592), .ZN(n4303) );
  INV_X1 U4629 ( .A(n4303), .ZN(n3750) );
  NAND2_X1 U4630 ( .A1(n3729), .A2(EBX_REG_0__SCAN_IN), .ZN(n3656) );
  INV_X1 U4631 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4399) );
  NAND2_X1 U4632 ( .A1(n2983), .A2(n4399), .ZN(n3655) );
  NAND2_X1 U4633 ( .A1(n3656), .A2(n3655), .ZN(n4397) );
  XNOR2_X1 U4634 ( .A(n3657), .B(n4397), .ZN(n4417) );
  OAI21_X1 U4635 ( .B1(n3654), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .A(n3658), 
        .ZN(n3659) );
  INV_X1 U4636 ( .A(n3659), .ZN(n4567) );
  MUX2_X1 U4637 ( .A(n5658), .B(n3724), .S(EBX_REG_3__SCAN_IN), .Z(n3661) );
  NAND2_X1 U4638 ( .A1(n4297), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3660)
         );
  NAND2_X1 U4639 ( .A1(n3661), .A2(n3660), .ZN(n4421) );
  OAI21_X1 U4640 ( .B1(n3654), .B2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n3662), 
        .ZN(n4592) );
  MUX2_X1 U4641 ( .A(n2983), .B(n3729), .S(EBX_REG_5__SCAN_IN), .Z(n3666) );
  AND2_X1 U4642 ( .A1(n4297), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3665)
         );
  NOR2_X1 U4643 ( .A1(n3666), .A2(n3665), .ZN(n4649) );
  OAI21_X1 U4644 ( .B1(n3654), .B2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n3668), 
        .ZN(n3669) );
  INV_X1 U4645 ( .A(n3669), .ZN(n4664) );
  OAI21_X1 U4646 ( .B1(n3654), .B2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n3670), 
        .ZN(n4850) );
  INV_X1 U4647 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U4648 ( .A1(n4418), .A2(n5998), .ZN(n3671) );
  OAI211_X1 U4649 ( .C1(n3729), .C2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n5658), 
        .B(n3671), .ZN(n3673) );
  NAND2_X1 U4650 ( .A1(n2983), .A2(n5998), .ZN(n3672) );
  NOR2_X1 U4651 ( .A1(n4850), .A2(n4849), .ZN(n3674) );
  INV_X1 U4652 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4999) );
  NAND2_X1 U4653 ( .A1(n4418), .A2(n4999), .ZN(n3675) );
  OAI211_X1 U4654 ( .C1(n2983), .C2(n3516), .A(n3724), .B(n3675), .ZN(n3677)
         );
  NAND2_X1 U4655 ( .A1(n3725), .A2(n4999), .ZN(n3676) );
  NAND2_X1 U4656 ( .A1(n3677), .A2(n3676), .ZN(n4349) );
  MUX2_X1 U4657 ( .A(n2983), .B(n3729), .S(EBX_REG_9__SCAN_IN), .Z(n3679) );
  AND2_X1 U4658 ( .A1(n4297), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3678)
         );
  NOR2_X1 U4659 ( .A1(n3679), .A2(n3678), .ZN(n4912) );
  INV_X1 U4660 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5057) );
  NAND2_X1 U4661 ( .A1(n4418), .A2(n5057), .ZN(n3682) );
  OAI211_X1 U4662 ( .C1(n3729), .C2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n5658), .B(n3682), .ZN(n3684) );
  NAND2_X1 U4663 ( .A1(n2983), .A2(n5057), .ZN(n3683) );
  OAI21_X1 U4664 ( .B1(n3654), .B2(INSTADDRPOINTER_REG_12__SCAN_IN), .A(n3685), 
        .ZN(n5072) );
  INV_X1 U4665 ( .A(n5072), .ZN(n3686) );
  MUX2_X1 U4666 ( .A(n5658), .B(n3724), .S(EBX_REG_13__SCAN_IN), .Z(n3688) );
  NAND2_X1 U4667 ( .A1(n4297), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3687) );
  NAND2_X1 U4668 ( .A1(n3688), .A2(n3687), .ZN(n5193) );
  OAI21_X1 U4669 ( .B1(n3654), .B2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n3689), 
        .ZN(n5210) );
  MUX2_X1 U4670 ( .A(n2983), .B(n3729), .S(EBX_REG_15__SCAN_IN), .Z(n3691) );
  AND2_X1 U4671 ( .A1(n4297), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3690)
         );
  NOR2_X1 U4672 ( .A1(n3691), .A2(n3690), .ZN(n5240) );
  OAI21_X1 U4673 ( .B1(n3654), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n3692), 
        .ZN(n3693) );
  INV_X1 U4674 ( .A(n3693), .ZN(n5273) );
  AND2_X2 U4675 ( .A1(n5274), .A2(n5273), .ZN(n5292) );
  INV_X1 U4676 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U4677 ( .A1(n4418), .A2(n5294), .ZN(n3694) );
  OAI211_X1 U4678 ( .C1(n3729), .C2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5658), .B(n3694), .ZN(n3696) );
  NAND2_X1 U4679 ( .A1(n2983), .A2(n5294), .ZN(n3695) );
  NAND2_X1 U4680 ( .A1(n3696), .A2(n3695), .ZN(n5291) );
  INV_X1 U4681 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U4682 ( .A1(n4418), .A2(n5772), .ZN(n3698) );
  NAND2_X1 U4683 ( .A1(n5658), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3697) );
  NAND3_X1 U4684 ( .A1(n3724), .A2(n3698), .A3(n3697), .ZN(n3700) );
  NAND2_X1 U4685 ( .A1(n3725), .A2(n5772), .ZN(n3699) );
  NAND2_X1 U4686 ( .A1(n3700), .A2(n3699), .ZN(n5488) );
  OAI22_X1 U4687 ( .A1(n3654), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n4297), .ZN(n5660) );
  INV_X1 U4688 ( .A(n3654), .ZN(n3701) );
  INV_X1 U4689 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5321) );
  AND2_X1 U4690 ( .A1(n4418), .A2(n5321), .ZN(n5315) );
  AOI21_X1 U4691 ( .B1(n3701), .B2(n6737), .A(n5315), .ZN(n5316) );
  NAND2_X1 U4692 ( .A1(n5316), .A2(n5660), .ZN(n3703) );
  INV_X1 U4693 ( .A(n5316), .ZN(n5659) );
  NAND2_X1 U4694 ( .A1(n5659), .A2(n5658), .ZN(n3702) );
  OAI211_X1 U4695 ( .C1(n5658), .C2(n5660), .A(n3703), .B(n3702), .ZN(n3704)
         );
  INV_X1 U4696 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5481) );
  NAND2_X1 U4697 ( .A1(n4418), .A2(n5481), .ZN(n3706) );
  NAND2_X1 U4698 ( .A1(n5658), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3705) );
  NAND3_X1 U4699 ( .A1(n3724), .A2(n3706), .A3(n3705), .ZN(n3708) );
  NAND2_X1 U4700 ( .A1(n3725), .A2(n5481), .ZN(n3707) );
  NAND2_X1 U4701 ( .A1(n3708), .A2(n3707), .ZN(n5437) );
  NOR2_X2 U4702 ( .A1(n5438), .A2(n5437), .ZN(n5426) );
  MUX2_X1 U4703 ( .A(n5658), .B(n3724), .S(EBX_REG_22__SCAN_IN), .Z(n3710) );
  NAND2_X1 U4704 ( .A1(n4297), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3709) );
  NAND2_X1 U4705 ( .A1(n3710), .A2(n3709), .ZN(n5425) );
  OAI21_X1 U4706 ( .B1(n3654), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n3711), 
        .ZN(n3712) );
  INV_X1 U4707 ( .A(n3712), .ZN(n5476) );
  INV_X1 U4708 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6750) );
  NAND2_X1 U4709 ( .A1(n4418), .A2(n6750), .ZN(n3713) );
  OAI211_X1 U4710 ( .C1(n3729), .C2(INSTADDRPOINTER_REG_24__SCAN_IN), .A(n5658), .B(n3713), .ZN(n3715) );
  NAND2_X1 U4711 ( .A1(n2983), .A2(n6750), .ZN(n3714) );
  NAND2_X1 U4712 ( .A1(n3715), .A2(n3714), .ZN(n5410) );
  INV_X1 U4713 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U4714 ( .A1(n4418), .A2(n5735), .ZN(n3717) );
  NAND2_X1 U4715 ( .A1(n5658), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3716) );
  NAND3_X1 U4716 ( .A1(n3724), .A2(n3717), .A3(n3716), .ZN(n3719) );
  NAND2_X1 U4717 ( .A1(n3725), .A2(n5735), .ZN(n3718) );
  NAND2_X1 U4718 ( .A1(n3719), .A2(n3718), .ZN(n5465) );
  MUX2_X1 U4719 ( .A(n2983), .B(n3729), .S(EBX_REG_26__SCAN_IN), .Z(n3721) );
  AND2_X1 U4720 ( .A1(n4297), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3720)
         );
  NOR2_X1 U4721 ( .A1(n3721), .A2(n3720), .ZN(n5398) );
  INV_X1 U4722 ( .A(EBX_REG_27__SCAN_IN), .ZN(n6690) );
  NAND2_X1 U4723 ( .A1(n4418), .A2(n6690), .ZN(n3723) );
  NAND2_X1 U4724 ( .A1(n5658), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3722) );
  NAND3_X1 U4725 ( .A1(n3724), .A2(n3723), .A3(n3722), .ZN(n3727) );
  NAND2_X1 U4726 ( .A1(n3725), .A2(n6690), .ZN(n3726) );
  AND2_X1 U4727 ( .A1(n3727), .A2(n3726), .ZN(n5604) );
  INV_X1 U4728 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U4729 ( .A1(n4418), .A2(n5459), .ZN(n3728) );
  OAI211_X1 U4730 ( .C1(n3729), .C2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n3728), .B(n5658), .ZN(n3731) );
  NAND2_X1 U4731 ( .A1(n2983), .A2(n5459), .ZN(n3730) );
  NAND2_X1 U4732 ( .A1(n3731), .A2(n3730), .ZN(n5383) );
  OAI22_X1 U4733 ( .A1(n3654), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n4297), .ZN(n4293) );
  INV_X1 U4734 ( .A(n4293), .ZN(n3732) );
  INV_X1 U4735 ( .A(n4296), .ZN(n3739) );
  NAND2_X1 U4736 ( .A1(n3654), .A2(EBX_REG_30__SCAN_IN), .ZN(n3735) );
  NAND2_X1 U4737 ( .A1(n4297), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3734) );
  NAND2_X1 U4738 ( .A1(n3735), .A2(n3734), .ZN(n4294) );
  AOI21_X1 U4739 ( .B1(n3736), .B2(n3733), .A(n3046), .ZN(n3738) );
  AOI21_X1 U4740 ( .B1(n3739), .B2(n3738), .A(n3737), .ZN(n5346) );
  NAND2_X1 U4741 ( .A1(n3608), .A2(n2984), .ZN(n6463) );
  NAND2_X1 U4742 ( .A1(n3621), .A2(n4559), .ZN(n3740) );
  NAND2_X1 U4743 ( .A1(n6463), .A2(n3740), .ZN(n3741) );
  NAND2_X1 U4744 ( .A1(n2971), .A2(REIP_REG_30__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U4745 ( .A1(n5254), .A2(n6217), .ZN(n5225) );
  NOR2_X1 U4746 ( .A1(n3744), .A2(n6151), .ZN(n5833) );
  NAND2_X1 U4747 ( .A1(n5676), .A2(n5663), .ZN(n5644) );
  NOR2_X1 U4748 ( .A1(n5631), .A2(n3747), .ZN(n5827) );
  INV_X1 U4749 ( .A(n3748), .ZN(n4300) );
  AOI21_X1 U4750 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n3750), .A(n3749), 
        .ZN(n3751) );
  NAND2_X1 U4751 ( .A1(n3752), .A2(n3936), .ZN(n3760) );
  NAND2_X1 U4752 ( .A1(n4277), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3789) );
  NAND2_X1 U4753 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n6601), .ZN(n3757)
         );
  NAND2_X1 U4754 ( .A1(n4313), .A2(EAX_REG_1__SCAN_IN), .ZN(n3756) );
  OAI211_X1 U4755 ( .C1(n3789), .C2(n3754), .A(n3757), .B(n3756), .ZN(n3758)
         );
  INV_X1 U4756 ( .A(n3758), .ZN(n3759) );
  NAND2_X1 U4757 ( .A1(n3760), .A2(n3759), .ZN(n4414) );
  NAND2_X1 U4758 ( .A1(n5028), .A2(n3091), .ZN(n3761) );
  NAND2_X1 U4759 ( .A1(n3761), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4389) );
  NAND2_X1 U4760 ( .A1(n4313), .A2(EAX_REG_0__SCAN_IN), .ZN(n3765) );
  NAND2_X1 U4761 ( .A1(n6601), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3764)
         );
  OAI211_X1 U4762 ( .C1(n3789), .C2(n3538), .A(n3765), .B(n3764), .ZN(n3766)
         );
  AOI21_X1 U4763 ( .B1(n3763), .B2(n3936), .A(n3766), .ZN(n3767) );
  OR2_X1 U4764 ( .A1(n4389), .A2(n3767), .ZN(n4390) );
  INV_X1 U4765 ( .A(n3767), .ZN(n4391) );
  NOR2_X1 U4766 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4202) );
  OR2_X1 U4767 ( .A1(n4391), .A2(n4251), .ZN(n3768) );
  NAND2_X1 U4768 ( .A1(n4390), .A2(n3768), .ZN(n4413) );
  NAND2_X1 U4769 ( .A1(n4414), .A2(n4413), .ZN(n4416) );
  INV_X1 U4770 ( .A(n3936), .ZN(n3887) );
  INV_X1 U4771 ( .A(n4312), .ZN(n3769) );
  INV_X1 U4772 ( .A(n3770), .ZN(n3774) );
  OAI21_X1 U4773 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3780), .ZN(n6136) );
  AOI22_X1 U4774 ( .A1(n4339), .A2(n6136), .B1(n4312), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3773) );
  NAND2_X1 U4775 ( .A1(n4313), .A2(EAX_REG_2__SCAN_IN), .ZN(n3772) );
  OAI211_X1 U4776 ( .C1(n3789), .C2(n3771), .A(n3773), .B(n3772), .ZN(n4572)
         );
  NAND2_X1 U4777 ( .A1(n4571), .A2(n4572), .ZN(n3778) );
  INV_X1 U4778 ( .A(n4416), .ZN(n3776) );
  INV_X1 U4779 ( .A(n3774), .ZN(n3775) );
  NAND2_X1 U4780 ( .A1(n3776), .A2(n3775), .ZN(n3777) );
  OAI21_X1 U4781 ( .B1(n3781), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n3790), 
        .ZN(n6128) );
  AOI22_X1 U4782 ( .A1(n6128), .A2(n4339), .B1(n4312), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3783) );
  NAND2_X1 U4783 ( .A1(n4313), .A2(EAX_REG_3__SCAN_IN), .ZN(n3782) );
  OAI211_X1 U4784 ( .C1(n3789), .C2(n4521), .A(n3783), .B(n3782), .ZN(n3784)
         );
  INV_X1 U4785 ( .A(n3784), .ZN(n3785) );
  NAND2_X1 U4786 ( .A1(n3786), .A2(n3936), .ZN(n3794) );
  INV_X1 U4787 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6602) );
  OAI21_X1 U4788 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6602), .A(n6601), 
        .ZN(n3788) );
  NAND2_X1 U4789 ( .A1(n4313), .A2(EAX_REG_4__SCAN_IN), .ZN(n3787) );
  OAI211_X1 U4790 ( .C1(n3789), .C2(n6613), .A(n3788), .B(n3787), .ZN(n3792)
         );
  AOI21_X1 U4791 ( .B1(n3790), .B2(n5964), .A(n3795), .ZN(n5969) );
  NAND2_X1 U4792 ( .A1(n5969), .A2(n4339), .ZN(n3791) );
  NAND2_X1 U4793 ( .A1(n3792), .A2(n3791), .ZN(n3793) );
  NAND2_X1 U4794 ( .A1(n3794), .A2(n3793), .ZN(n4585) );
  INV_X1 U4795 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4987) );
  NAND2_X1 U4796 ( .A1(n4312), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3797)
         );
  OAI21_X1 U4797 ( .B1(n3795), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3807), 
        .ZN(n6119) );
  NAND2_X1 U4798 ( .A1(n6119), .A2(n4339), .ZN(n3796) );
  OAI211_X1 U4799 ( .C1(n4254), .C2(n4987), .A(n3797), .B(n3796), .ZN(n3798)
         );
  NAND2_X1 U4800 ( .A1(n4313), .A2(EAX_REG_6__SCAN_IN), .ZN(n3801) );
  OAI21_X1 U4801 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6602), .A(n6601), 
        .ZN(n3800) );
  XNOR2_X1 U4802 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n3807), .ZN(n5949) );
  AOI22_X1 U4803 ( .A1(n3801), .A2(n3800), .B1(n4339), .B2(n5949), .ZN(n3802)
         );
  AOI21_X1 U4804 ( .B1(n3803), .B2(n3936), .A(n3802), .ZN(n4667) );
  NAND2_X1 U4805 ( .A1(n3805), .A2(n3936), .ZN(n3812) );
  OAI21_X1 U4806 ( .B1(n3808), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3827), 
        .ZN(n6113) );
  NAND2_X1 U4807 ( .A1(n6113), .A2(n4339), .ZN(n3810) );
  AOI22_X1 U4808 ( .A1(n4313), .A2(EAX_REG_7__SCAN_IN), .B1(n4312), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3809) );
  AND2_X1 U4809 ( .A1(n3810), .A2(n3809), .ZN(n3811) );
  NAND2_X1 U4810 ( .A1(n4666), .A2(n4916), .ZN(n4855) );
  XNOR2_X1 U4811 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3827), .ZN(n4981) );
  INV_X1 U4812 ( .A(n4981), .ZN(n4992) );
  AOI22_X1 U4813 ( .A1(n2980), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4814 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n4165), .B1(n4228), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4815 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4189), .B1(n4232), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4816 ( .A1(n4238), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3813) );
  NAND4_X1 U4817 ( .A1(n3816), .A2(n3815), .A3(n3814), .A4(n3813), .ZN(n3822)
         );
  AOI22_X1 U4818 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n4237), .B1(n4231), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4819 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n4188), .B1(n4239), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4820 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n4230), .B1(n4240), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4821 ( .A1(n4229), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3817) );
  NAND4_X1 U4822 ( .A1(n3820), .A2(n3819), .A3(n3818), .A4(n3817), .ZN(n3821)
         );
  OAI21_X1 U4823 ( .B1(n3822), .B2(n3821), .A(n3936), .ZN(n3825) );
  NAND2_X1 U4824 ( .A1(n4313), .A2(EAX_REG_8__SCAN_IN), .ZN(n3824) );
  NAND2_X1 U4825 ( .A1(n4312), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3823)
         );
  NAND3_X1 U4826 ( .A1(n3825), .A2(n3824), .A3(n3823), .ZN(n3826) );
  AOI21_X1 U4827 ( .B1(n4992), .B2(n4339), .A(n3826), .ZN(n4854) );
  XNOR2_X1 U4828 ( .A(n3842), .B(n5101), .ZN(n5097) );
  AOI22_X1 U4829 ( .A1(n4238), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4189), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4830 ( .A1(n4188), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3830) );
  AOI22_X1 U4831 ( .A1(n4229), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4832 ( .A1(n2968), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3828) );
  NAND4_X1 U4833 ( .A1(n3831), .A2(n3830), .A3(n3829), .A4(n3828), .ZN(n3837)
         );
  AOI22_X1 U4834 ( .A1(n4231), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4835 ( .A1(n4165), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4836 ( .A1(n4069), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4837 ( .A1(n4228), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4240), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3832) );
  NAND4_X1 U4838 ( .A1(n3835), .A2(n3834), .A3(n3833), .A4(n3832), .ZN(n3836)
         );
  OAI21_X1 U4839 ( .B1(n3837), .B2(n3836), .A(n3936), .ZN(n3840) );
  NAND2_X1 U4840 ( .A1(n4313), .A2(EAX_REG_9__SCAN_IN), .ZN(n3839) );
  NAND2_X1 U4841 ( .A1(n4312), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3838)
         );
  NAND3_X1 U4842 ( .A1(n3840), .A2(n3839), .A3(n3838), .ZN(n3841) );
  NOR2_X2 U4843 ( .A1(n2972), .A2(n4855), .ZN(n4336) );
  INV_X1 U4844 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4352) );
  XNOR2_X1 U4845 ( .A(n4352), .B(n3856), .ZN(n5111) );
  AOI22_X1 U4846 ( .A1(n2968), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4189), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4847 ( .A1(n4231), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4848 ( .A1(n4188), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4228), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4849 ( .A1(n4229), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3843) );
  NAND4_X1 U4850 ( .A1(n3846), .A2(n3845), .A3(n3844), .A4(n3843), .ZN(n3852)
         );
  AOI22_X1 U4851 ( .A1(n4238), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4852 ( .A1(n4165), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4853 ( .A1(n4232), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4854 ( .A1(n4240), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3847) );
  NAND4_X1 U4855 ( .A1(n3850), .A2(n3849), .A3(n3848), .A4(n3847), .ZN(n3851)
         );
  OR2_X1 U4856 ( .A1(n3852), .A2(n3851), .ZN(n3853) );
  AOI22_X1 U4857 ( .A1(n3936), .A2(n3853), .B1(n4312), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3855) );
  NAND2_X1 U4858 ( .A1(n4313), .A2(EAX_REG_10__SCAN_IN), .ZN(n3854) );
  OAI211_X1 U4859 ( .C1(n5111), .C2(n4251), .A(n3855), .B(n3854), .ZN(n4337)
         );
  NAND2_X1 U4860 ( .A1(n3857), .A2(n6703), .ZN(n3859) );
  INV_X1 U4861 ( .A(n3891), .ZN(n3858) );
  NAND2_X1 U4862 ( .A1(n3859), .A2(n3858), .ZN(n5133) );
  NAND2_X1 U4863 ( .A1(n5133), .A2(n4339), .ZN(n3874) );
  AOI22_X1 U4864 ( .A1(n4238), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n2980), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4865 ( .A1(n4228), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4866 ( .A1(n4188), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4867 ( .A1(n4069), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3860) );
  NAND4_X1 U4868 ( .A1(n3863), .A2(n3862), .A3(n3861), .A4(n3860), .ZN(n3869)
         );
  AOI22_X1 U4869 ( .A1(n4189), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4870 ( .A1(n4231), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4871 ( .A1(n4165), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4872 ( .A1(n4240), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3864) );
  NAND4_X1 U4873 ( .A1(n3867), .A2(n3866), .A3(n3865), .A4(n3864), .ZN(n3868)
         );
  OAI21_X1 U4874 ( .B1(n3869), .B2(n3868), .A(n3936), .ZN(n3872) );
  NAND2_X1 U4875 ( .A1(n4313), .A2(EAX_REG_11__SCAN_IN), .ZN(n3871) );
  NAND2_X1 U4876 ( .A1(n4312), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3870)
         );
  AND3_X1 U4877 ( .A1(n3872), .A2(n3871), .A3(n3870), .ZN(n3873) );
  NAND2_X1 U4878 ( .A1(n3874), .A2(n3873), .ZN(n4997) );
  INV_X1 U4879 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5923) );
  XNOR2_X1 U4880 ( .A(n5923), .B(n3891), .ZN(n5919) );
  NAND2_X1 U4881 ( .A1(n5919), .A2(n4339), .ZN(n3890) );
  INV_X1 U4882 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5074) );
  OAI21_X1 U4883 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6602), .A(n6601), 
        .ZN(n3875) );
  OAI21_X1 U4884 ( .B1(n4254), .B2(n5074), .A(n3875), .ZN(n3889) );
  AOI22_X1 U4885 ( .A1(n4165), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n2980), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4886 ( .A1(n4231), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4887 ( .A1(n3199), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4888 ( .A1(n4189), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3876) );
  NAND4_X1 U4889 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3885)
         );
  AOI22_X1 U4890 ( .A1(n4238), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4891 ( .A1(n4228), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4892 ( .A1(n4229), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4893 ( .A1(n4069), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4240), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3880) );
  NAND4_X1 U4894 ( .A1(n3883), .A2(n3882), .A3(n3881), .A4(n3880), .ZN(n3884)
         );
  NOR2_X1 U4895 ( .A1(n3885), .A2(n3884), .ZN(n3886) );
  NOR2_X1 U4896 ( .A1(n3887), .A2(n3886), .ZN(n3888) );
  AOI21_X1 U4897 ( .B1(n3890), .B2(n3889), .A(n3888), .ZN(n5069) );
  NAND2_X1 U4898 ( .A1(n4313), .A2(EAX_REG_13__SCAN_IN), .ZN(n3894) );
  INV_X1 U4899 ( .A(n3920), .ZN(n3892) );
  XNOR2_X1 U4900 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n3892), .ZN(n5250)
         );
  AOI22_X1 U4901 ( .A1(n4202), .A2(n5250), .B1(n4312), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3893) );
  NAND2_X1 U4902 ( .A1(n3894), .A2(n3893), .ZN(n3908) );
  AOI22_X1 U4903 ( .A1(n4069), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4904 ( .A1(n2980), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4905 ( .A1(n4231), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4070), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4906 ( .A1(n4237), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3896) );
  NAND4_X1 U4907 ( .A1(n3899), .A2(n3898), .A3(n3897), .A4(n3896), .ZN(n3905)
         );
  AOI22_X1 U4908 ( .A1(n4228), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4240), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4909 ( .A1(n4165), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4910 ( .A1(n4238), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4911 ( .A1(n4189), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3900) );
  NAND4_X1 U4912 ( .A1(n3903), .A2(n3902), .A3(n3901), .A4(n3900), .ZN(n3904)
         );
  OR2_X1 U4913 ( .A1(n3905), .A2(n3904), .ZN(n3906) );
  AND2_X1 U4914 ( .A1(n3936), .A2(n3906), .ZN(n5189) );
  AOI22_X1 U4915 ( .A1(n4229), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4228), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4916 ( .A1(n4231), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4917 ( .A1(n4069), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4918 ( .A1(n4238), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3909) );
  NAND4_X1 U4919 ( .A1(n3912), .A2(n3911), .A3(n3910), .A4(n3909), .ZN(n3918)
         );
  AOI22_X1 U4920 ( .A1(n4165), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4921 ( .A1(n4188), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4922 ( .A1(n2968), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4923 ( .A1(n4189), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4240), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3913) );
  NAND4_X1 U4924 ( .A1(n3916), .A2(n3915), .A3(n3914), .A4(n3913), .ZN(n3917)
         );
  OAI21_X1 U4925 ( .B1(n3918), .B2(n3917), .A(n3936), .ZN(n3923) );
  XNOR2_X1 U4926 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3924), .ZN(n5282)
         );
  AOI22_X1 U4927 ( .A1(n4202), .A2(n5282), .B1(n4312), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3922) );
  NAND2_X1 U4928 ( .A1(n4313), .A2(EAX_REG_14__SCAN_IN), .ZN(n3921) );
  XNOR2_X1 U4929 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3939), .ZN(n5914)
         );
  AOI22_X1 U4930 ( .A1(n4238), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4931 ( .A1(n2968), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4932 ( .A1(n4230), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4933 ( .A1(n4229), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3925) );
  NAND4_X1 U4934 ( .A1(n3928), .A2(n3927), .A3(n3926), .A4(n3925), .ZN(n3934)
         );
  AOI22_X1 U4935 ( .A1(n4231), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4936 ( .A1(n4189), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4937 ( .A1(n4165), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4240), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4938 ( .A1(n4228), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3929) );
  NAND4_X1 U4939 ( .A1(n3932), .A2(n3931), .A3(n3930), .A4(n3929), .ZN(n3933)
         );
  OR2_X1 U4940 ( .A1(n3934), .A2(n3933), .ZN(n3935) );
  AOI22_X1 U4941 ( .A1(n3936), .A2(n3935), .B1(n4312), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3938) );
  NAND2_X1 U4942 ( .A1(n4313), .A2(EAX_REG_15__SCAN_IN), .ZN(n3937) );
  OAI211_X1 U4943 ( .C1(n5914), .C2(n4251), .A(n3938), .B(n3937), .ZN(n5238)
         );
  INV_X1 U4944 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5907) );
  INV_X1 U4945 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3940) );
  XNOR2_X1 U4946 ( .A(n3970), .B(n3940), .ZN(n5900) );
  OR2_X1 U4947 ( .A1(n5900), .A2(n4251), .ZN(n3955) );
  AOI22_X1 U4948 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n4188), .B1(n4228), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4949 ( .A1(n4237), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4950 ( .A1(n4069), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4951 ( .A1(n2980), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3941) );
  NAND4_X1 U4952 ( .A1(n3944), .A2(n3943), .A3(n3942), .A4(n3941), .ZN(n3950)
         );
  AOI22_X1 U4953 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4165), .B1(n4231), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4954 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n4238), .B1(n4229), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4955 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n4232), .B1(n4239), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4956 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n4189), .B1(n4240), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3945) );
  NAND4_X1 U4957 ( .A1(n3948), .A2(n3947), .A3(n3946), .A4(n3945), .ZN(n3949)
         );
  NOR2_X1 U4958 ( .A1(n3950), .A2(n3949), .ZN(n3952) );
  AOI22_X1 U4959 ( .A1(n4313), .A2(EAX_REG_16__SCAN_IN), .B1(n4312), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3951) );
  OAI21_X1 U4960 ( .B1(n4154), .B2(n3952), .A(n3951), .ZN(n3953) );
  INV_X1 U4961 ( .A(n3953), .ZN(n3954) );
  NAND2_X1 U4962 ( .A1(n3955), .A2(n3954), .ZN(n5271) );
  AOI22_X1 U4963 ( .A1(n4189), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3266), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4964 ( .A1(n4237), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4965 ( .A1(n4239), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4966 ( .A1(n2968), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3956) );
  NAND4_X1 U4967 ( .A1(n3959), .A2(n3958), .A3(n3957), .A4(n3956), .ZN(n3965)
         );
  AOI22_X1 U4968 ( .A1(n4165), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4231), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4969 ( .A1(n4188), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4229), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4970 ( .A1(n4238), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4971 ( .A1(n4228), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4240), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3960) );
  NAND4_X1 U4972 ( .A1(n3963), .A2(n3962), .A3(n3961), .A4(n3960), .ZN(n3964)
         );
  NOR2_X1 U4973 ( .A1(n3965), .A2(n3964), .ZN(n3969) );
  OAI21_X1 U4974 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6602), .A(n6601), 
        .ZN(n3966) );
  INV_X1 U4975 ( .A(n3966), .ZN(n3967) );
  AOI21_X1 U4976 ( .B1(n4313), .B2(EAX_REG_17__SCAN_IN), .A(n3967), .ZN(n3968)
         );
  OAI21_X1 U4977 ( .B1(n4154), .B2(n3969), .A(n3968), .ZN(n3974) );
  OAI21_X1 U4978 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3971), .A(n3993), 
        .ZN(n3972) );
  INV_X1 U4979 ( .A(n3972), .ZN(n5822) );
  NAND2_X1 U4980 ( .A1(n5822), .A2(n4339), .ZN(n3973) );
  NAND2_X1 U4981 ( .A1(n3974), .A2(n3973), .ZN(n5288) );
  AOI22_X1 U4982 ( .A1(n4188), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4983 ( .A1(n2968), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4228), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4984 ( .A1(n4231), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4985 ( .A1(n4238), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3976) );
  NAND4_X1 U4986 ( .A1(n3979), .A2(n3978), .A3(n3977), .A4(n3976), .ZN(n3987)
         );
  AOI22_X1 U4987 ( .A1(n4165), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3278), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4988 ( .A1(n4229), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4240), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4989 ( .A1(n4230), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3983) );
  AOI21_X1 U4990 ( .B1(n4081), .B2(INSTQUEUE_REG_9__2__SCAN_IN), .A(n4202), 
        .ZN(n3981) );
  NAND2_X1 U4991 ( .A1(n4237), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3980) );
  AND2_X1 U4992 ( .A1(n3981), .A2(n3980), .ZN(n3982) );
  NAND4_X1 U4993 ( .A1(n3985), .A2(n3984), .A3(n3983), .A4(n3982), .ZN(n3986)
         );
  NAND2_X1 U4994 ( .A1(n4154), .A2(n4251), .ZN(n4056) );
  OAI21_X1 U4995 ( .B1(n3987), .B2(n3986), .A(n4056), .ZN(n3989) );
  AOI22_X1 U4996 ( .A1(n4313), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6601), .ZN(n3988) );
  NAND2_X1 U4997 ( .A1(n3989), .A2(n3988), .ZN(n3991) );
  XNOR2_X1 U4998 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3993), .ZN(n5891)
         );
  NAND2_X1 U4999 ( .A1(n4202), .A2(n5891), .ZN(n3990) );
  NAND2_X1 U5000 ( .A1(n3991), .A2(n3990), .ZN(n5313) );
  INV_X1 U5001 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3992) );
  OR2_X1 U5002 ( .A1(n3994), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3995)
         );
  NAND2_X1 U5003 ( .A1(n3995), .A2(n4041), .ZN(n5817) );
  AOI22_X1 U5004 ( .A1(n4231), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n2980), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U5005 ( .A1(n4229), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U5006 ( .A1(n4188), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U5007 ( .A1(n4189), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3996) );
  NAND4_X1 U5008 ( .A1(n3999), .A2(n3998), .A3(n3997), .A4(n3996), .ZN(n4005)
         );
  AOI22_X1 U5009 ( .A1(n4165), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4228), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U5010 ( .A1(n4069), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4240), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U5011 ( .A1(n4238), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U5012 ( .A1(n4237), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4000) );
  NAND4_X1 U5013 ( .A1(n4003), .A2(n4002), .A3(n4001), .A4(n4000), .ZN(n4004)
         );
  NOR2_X1 U5014 ( .A1(n4005), .A2(n4004), .ZN(n4008) );
  OAI21_X1 U5015 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6602), .A(n6601), 
        .ZN(n4007) );
  NAND2_X1 U5016 ( .A1(n4313), .A2(EAX_REG_19__SCAN_IN), .ZN(n4006) );
  OAI211_X1 U5017 ( .C1(n4154), .C2(n4008), .A(n4007), .B(n4006), .ZN(n4009)
         );
  OAI21_X1 U5018 ( .B1(n5817), .B2(n4251), .A(n4009), .ZN(n5485) );
  AOI22_X1 U5019 ( .A1(n2968), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U5020 ( .A1(n3199), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4240), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4015) );
  AOI21_X1 U5021 ( .B1(n4081), .B2(INSTQUEUE_REG_9__4__SCAN_IN), .A(n4202), 
        .ZN(n4012) );
  NAND2_X1 U5022 ( .A1(n4165), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4011)
         );
  AND2_X1 U5023 ( .A1(n4012), .A2(n4011), .ZN(n4014) );
  AOI22_X1 U5024 ( .A1(n3278), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4013) );
  NAND4_X1 U5025 ( .A1(n4016), .A2(n4015), .A3(n4014), .A4(n4013), .ZN(n4022)
         );
  AOI22_X1 U5026 ( .A1(n4188), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4229), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U5027 ( .A1(n4237), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U5028 ( .A1(n4231), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U5029 ( .A1(n4228), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4017) );
  NAND4_X1 U5030 ( .A1(n4020), .A2(n4019), .A3(n4018), .A4(n4017), .ZN(n4021)
         );
  OR2_X1 U5031 ( .A1(n4022), .A2(n4021), .ZN(n4023) );
  NAND2_X1 U5032 ( .A1(n4056), .A2(n4023), .ZN(n4026) );
  AOI22_X1 U5033 ( .A1(n4313), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6601), .ZN(n4025) );
  XNOR2_X1 U5034 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n4041), .ZN(n5758)
         );
  AOI21_X1 U5035 ( .B1(n4026), .B2(n4025), .A(n4024), .ZN(n5569) );
  AOI22_X1 U5036 ( .A1(n2968), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U5037 ( .A1(n4231), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4029) );
  AOI22_X1 U5038 ( .A1(n4165), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4069), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U5039 ( .A1(n4229), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4027) );
  NAND4_X1 U5040 ( .A1(n4030), .A2(n4029), .A3(n4028), .A4(n4027), .ZN(n4036)
         );
  AOI22_X1 U5041 ( .A1(n4238), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U5042 ( .A1(n4228), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U5043 ( .A1(n4189), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4240), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U5044 ( .A1(n4230), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4031) );
  NAND4_X1 U5045 ( .A1(n4034), .A2(n4033), .A3(n4032), .A4(n4031), .ZN(n4035)
         );
  NOR2_X1 U5046 ( .A1(n4036), .A2(n4035), .ZN(n4040) );
  NAND2_X1 U5047 ( .A1(n6601), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4037)
         );
  NAND2_X1 U5048 ( .A1(n4251), .A2(n4037), .ZN(n4038) );
  AOI21_X1 U5049 ( .B1(n4313), .B2(EAX_REG_21__SCAN_IN), .A(n4038), .ZN(n4039)
         );
  OAI21_X1 U5050 ( .B1(n4154), .B2(n4040), .A(n4039), .ZN(n4045) );
  OAI21_X1 U5051 ( .B1(n4043), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n4095), 
        .ZN(n5564) );
  OR2_X1 U5052 ( .A1(n5564), .A2(n4251), .ZN(n4044) );
  NAND2_X1 U5053 ( .A1(n4045), .A2(n4044), .ZN(n5434) );
  AOI22_X1 U5054 ( .A1(n2980), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3278), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U5055 ( .A1(n4165), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U5056 ( .A1(n4069), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U5057 ( .A1(n4229), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4046) );
  NAND4_X1 U5058 ( .A1(n4049), .A2(n4048), .A3(n4047), .A4(n4046), .ZN(n4058)
         );
  AOI22_X1 U5059 ( .A1(n4188), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U5060 ( .A1(n4238), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4240), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4054) );
  AOI21_X1 U5061 ( .B1(n4081), .B2(INSTQUEUE_REG_9__6__SCAN_IN), .A(n4202), 
        .ZN(n4051) );
  NAND2_X1 U5062 ( .A1(n4164), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4050) );
  AND2_X1 U5063 ( .A1(n4051), .A2(n4050), .ZN(n4053) );
  AOI22_X1 U5064 ( .A1(n4228), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4052) );
  NAND4_X1 U5065 ( .A1(n4055), .A2(n4054), .A3(n4053), .A4(n4052), .ZN(n4057)
         );
  OAI21_X1 U5066 ( .B1(n4058), .B2(n4057), .A(n4056), .ZN(n4061) );
  INV_X1 U5067 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5554) );
  NOR2_X1 U5068 ( .A1(n5554), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4059) );
  AOI21_X1 U5069 ( .B1(n4313), .B2(EAX_REG_22__SCAN_IN), .A(n4059), .ZN(n4060)
         );
  NAND2_X1 U5070 ( .A1(n4061), .A2(n4060), .ZN(n4063) );
  XNOR2_X1 U5071 ( .A(n4095), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5558)
         );
  NAND2_X1 U5072 ( .A1(n5558), .A2(n4339), .ZN(n4062) );
  NAND2_X1 U5073 ( .A1(n4063), .A2(n4062), .ZN(n5418) );
  AOI22_X1 U5074 ( .A1(n2968), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4189), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U5075 ( .A1(n4164), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U5076 ( .A1(n4165), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U5077 ( .A1(n4240), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4065) );
  NAND4_X1 U5078 ( .A1(n4068), .A2(n4067), .A3(n4066), .A4(n4065), .ZN(n4076)
         );
  AOI22_X1 U5079 ( .A1(n4238), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4074) );
  AOI22_X1 U5080 ( .A1(n4069), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U5081 ( .A1(n4228), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U5082 ( .A1(n4070), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4071) );
  NAND4_X1 U5083 ( .A1(n4074), .A2(n4073), .A3(n4072), .A4(n4071), .ZN(n4075)
         );
  OR2_X1 U5084 ( .A1(n4076), .A2(n4075), .ZN(n4090) );
  AOI22_X1 U5085 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n4189), .B1(n2980), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4080) );
  AOI22_X1 U5086 ( .A1(n4164), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4079) );
  AOI22_X1 U5087 ( .A1(n4165), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U5088 ( .A1(n4240), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4077) );
  NAND4_X1 U5089 ( .A1(n4080), .A2(n4079), .A3(n4078), .A4(n4077), .ZN(n4087)
         );
  AOI22_X1 U5090 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n4238), .B1(n4188), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4085) );
  INV_X1 U5091 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n6739) );
  AOI22_X1 U5092 ( .A1(n3266), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U5093 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4228), .B1(n4239), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U5094 ( .A1(n4229), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4082) );
  NAND4_X1 U5095 ( .A1(n4085), .A2(n4084), .A3(n4083), .A4(n4082), .ZN(n4086)
         );
  OR2_X1 U5096 ( .A1(n4087), .A2(n4086), .ZN(n4089) );
  AND2_X1 U5097 ( .A1(n4089), .A2(n4090), .ZN(n4128) );
  INV_X1 U5098 ( .A(n4128), .ZN(n4088) );
  OAI21_X1 U5099 ( .B1(n4090), .B2(n4089), .A(n4088), .ZN(n4094) );
  NAND2_X1 U5100 ( .A1(n6601), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4091)
         );
  NAND2_X1 U5101 ( .A1(n4251), .A2(n4091), .ZN(n4092) );
  AOI21_X1 U5102 ( .B1(n4313), .B2(EAX_REG_23__SCAN_IN), .A(n4092), .ZN(n4093)
         );
  OAI21_X1 U5103 ( .B1(n4154), .B2(n4094), .A(n4093), .ZN(n4100) );
  NOR2_X1 U5104 ( .A1(n4096), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4097)
         );
  OR2_X1 U5105 ( .A1(n4113), .A2(n4097), .ZN(n5745) );
  INV_X1 U5106 ( .A(n5745), .ZN(n4098) );
  NAND2_X1 U5107 ( .A1(n4098), .A2(n4339), .ZN(n4099) );
  INV_X1 U5108 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4117) );
  AOI22_X1 U5109 ( .A1(n2980), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4189), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U5110 ( .A1(n4164), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5111 ( .A1(n2970), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U5112 ( .A1(n4240), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4102) );
  NAND4_X1 U5113 ( .A1(n4105), .A2(n4104), .A3(n4103), .A4(n4102), .ZN(n4111)
         );
  AOI22_X1 U5114 ( .A1(n4238), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U5115 ( .A1(n3266), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3199), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U5116 ( .A1(n4228), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U5117 ( .A1(n4229), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4106) );
  NAND4_X1 U5118 ( .A1(n4109), .A2(n4108), .A3(n4107), .A4(n4106), .ZN(n4110)
         );
  OR2_X1 U5119 ( .A1(n4111), .A2(n4110), .ZN(n4129) );
  XNOR2_X1 U5120 ( .A(n4128), .B(n4129), .ZN(n4112) );
  OR2_X1 U5121 ( .A1(n4154), .A2(n4112), .ZN(n4116) );
  NOR2_X1 U5122 ( .A1(n4113), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4114)
         );
  OR2_X1 U5123 ( .A1(n4135), .A2(n4114), .ZN(n5542) );
  AOI22_X1 U5124 ( .A1(n5542), .A2(n4202), .B1(n4312), .B2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4115) );
  OAI211_X1 U5125 ( .C1(n4254), .C2(n4117), .A(n4116), .B(n4115), .ZN(n5407)
         );
  NAND2_X1 U5126 ( .A1(n5405), .A2(n5407), .ZN(n5406) );
  AOI22_X1 U5127 ( .A1(n2969), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n2968), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4121) );
  AOI22_X1 U5128 ( .A1(n3266), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4229), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U5129 ( .A1(n4189), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4119) );
  AOI22_X1 U5130 ( .A1(n4228), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4118) );
  NAND4_X1 U5131 ( .A1(n4121), .A2(n4120), .A3(n4119), .A4(n4118), .ZN(n4127)
         );
  AOI22_X1 U5132 ( .A1(n4143), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5133 ( .A1(n4237), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5134 ( .A1(n4231), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4240), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U5135 ( .A1(n4230), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4122) );
  NAND4_X1 U5136 ( .A1(n4125), .A2(n4124), .A3(n4123), .A4(n4122), .ZN(n4126)
         );
  OR2_X1 U5137 ( .A1(n4127), .A2(n4126), .ZN(n4140) );
  NAND2_X1 U5138 ( .A1(n4129), .A2(n4128), .ZN(n4142) );
  INV_X1 U5139 ( .A(n4142), .ZN(n4130) );
  XNOR2_X1 U5140 ( .A(n4140), .B(n4130), .ZN(n4134) );
  INV_X1 U5141 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4131) );
  AOI21_X1 U5142 ( .B1(n4131), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4132) );
  AOI21_X1 U5143 ( .B1(n4313), .B2(EAX_REG_25__SCAN_IN), .A(n4132), .ZN(n4133)
         );
  OAI21_X1 U5144 ( .B1(n4154), .B2(n4134), .A(n4133), .ZN(n4139) );
  OR2_X1 U5145 ( .A1(n4135), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4136)
         );
  NAND2_X1 U5146 ( .A1(n4136), .A2(n4181), .ZN(n5812) );
  INV_X1 U5147 ( .A(n5812), .ZN(n4137) );
  NAND2_X1 U5148 ( .A1(n4137), .A2(n4339), .ZN(n4138) );
  NAND2_X1 U5149 ( .A1(n4139), .A2(n4138), .ZN(n5464) );
  INV_X1 U5150 ( .A(n4140), .ZN(n4141) );
  OR2_X1 U5151 ( .A1(n4142), .A2(n4141), .ZN(n4162) );
  AOI22_X1 U5152 ( .A1(n4143), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3278), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4147) );
  AOI22_X1 U5153 ( .A1(n2970), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4146) );
  AOI22_X1 U5154 ( .A1(n3266), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4145) );
  AOI22_X1 U5155 ( .A1(n4229), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4144) );
  NAND4_X1 U5156 ( .A1(n4147), .A2(n4146), .A3(n4145), .A4(n4144), .ZN(n4153)
         );
  AOI22_X1 U5157 ( .A1(n2980), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4228), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4151) );
  AOI22_X1 U5158 ( .A1(n4164), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U5159 ( .A1(n4188), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U5160 ( .A1(n4240), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4148) );
  NAND4_X1 U5161 ( .A1(n4151), .A2(n4150), .A3(n4149), .A4(n4148), .ZN(n4152)
         );
  NOR2_X1 U5162 ( .A1(n4153), .A2(n4152), .ZN(n4163) );
  XOR2_X1 U5163 ( .A(n4162), .B(n4163), .Z(n4155) );
  INV_X1 U5164 ( .A(n4154), .ZN(n4256) );
  NAND2_X1 U5165 ( .A1(n4155), .A2(n4256), .ZN(n4158) );
  INV_X1 U5166 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5530) );
  OAI21_X1 U5167 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5530), .A(n4251), .ZN(
        n4156) );
  AOI21_X1 U5168 ( .B1(n4313), .B2(EAX_REG_26__SCAN_IN), .A(n4156), .ZN(n4157)
         );
  NAND2_X1 U5169 ( .A1(n4158), .A2(n4157), .ZN(n4160) );
  XNOR2_X1 U5170 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .B(n4181), .ZN(n5528)
         );
  NAND2_X1 U5171 ( .A1(n4339), .A2(n5528), .ZN(n4159) );
  NAND2_X1 U5172 ( .A1(n4160), .A2(n4159), .ZN(n5397) );
  NAND2_X1 U5173 ( .A1(n5394), .A2(n4161), .ZN(n5395) );
  NOR2_X1 U5174 ( .A1(n4163), .A2(n4162), .ZN(n4187) );
  AOI22_X1 U5175 ( .A1(n2968), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4189), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U5176 ( .A1(n4164), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U5177 ( .A1(n4165), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4167) );
  AOI22_X1 U5178 ( .A1(n4240), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4166) );
  NAND4_X1 U5179 ( .A1(n4169), .A2(n4168), .A3(n4167), .A4(n4166), .ZN(n4175)
         );
  AOI22_X1 U5180 ( .A1(n4238), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4173) );
  AOI22_X1 U5181 ( .A1(n4069), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4172) );
  AOI22_X1 U5182 ( .A1(n4228), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4171) );
  AOI22_X1 U5183 ( .A1(n4229), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4170) );
  NAND4_X1 U5184 ( .A1(n4173), .A2(n4172), .A3(n4171), .A4(n4170), .ZN(n4174)
         );
  OR2_X1 U5185 ( .A1(n4175), .A2(n4174), .ZN(n4186) );
  INV_X1 U5186 ( .A(n4186), .ZN(n4176) );
  XNOR2_X1 U5187 ( .A(n4187), .B(n4176), .ZN(n4180) );
  INV_X1 U5188 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4178) );
  NAND2_X1 U5189 ( .A1(n6601), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4177)
         );
  OAI211_X1 U5190 ( .C1(n4254), .C2(n4178), .A(n4251), .B(n4177), .ZN(n4179)
         );
  AOI21_X1 U5191 ( .B1(n4180), .B2(n4256), .A(n4179), .ZN(n4185) );
  INV_X1 U5192 ( .A(n4181), .ZN(n4182) );
  OAI21_X1 U5193 ( .B1(n4183), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n4223), 
        .ZN(n5725) );
  NOR2_X1 U5194 ( .A1(n5725), .A2(n4251), .ZN(n4184) );
  NOR2_X2 U5195 ( .A1(n5395), .A2(n5518), .ZN(n5378) );
  NAND2_X1 U5196 ( .A1(n4187), .A2(n4186), .ZN(n4206) );
  AOI22_X1 U5197 ( .A1(n4189), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4193) );
  AOI22_X1 U5198 ( .A1(n4237), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4192) );
  AOI22_X1 U5199 ( .A1(n2969), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4191) );
  AOI22_X1 U5200 ( .A1(n4069), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4190) );
  NAND4_X1 U5201 ( .A1(n4193), .A2(n4192), .A3(n4191), .A4(n4190), .ZN(n4199)
         );
  AOI22_X1 U5202 ( .A1(n4238), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4229), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4197) );
  AOI22_X1 U5203 ( .A1(n2980), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4196) );
  AOI22_X1 U5204 ( .A1(n4228), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4240), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4195) );
  AOI22_X1 U5205 ( .A1(n4231), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4194) );
  NAND4_X1 U5206 ( .A1(n4197), .A2(n4196), .A3(n4195), .A4(n4194), .ZN(n4198)
         );
  NOR2_X1 U5207 ( .A1(n4199), .A2(n4198), .ZN(n4207) );
  XOR2_X1 U5208 ( .A(n4206), .B(n4207), .Z(n4200) );
  NAND2_X1 U5209 ( .A1(n4200), .A2(n4256), .ZN(n4205) );
  INV_X1 U5210 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5513) );
  OAI21_X1 U5211 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5513), .A(n4251), .ZN(
        n4201) );
  AOI21_X1 U5212 ( .B1(n4313), .B2(EAX_REG_28__SCAN_IN), .A(n4201), .ZN(n4204)
         );
  XNOR2_X1 U5213 ( .A(n4223), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5511)
         );
  AND2_X1 U5214 ( .A1(n5511), .A2(n4202), .ZN(n4203) );
  AOI21_X1 U5215 ( .B1(n4205), .B2(n4204), .A(n4203), .ZN(n5380) );
  NOR2_X1 U5216 ( .A1(n4207), .A2(n4206), .ZN(n4248) );
  AOI22_X1 U5217 ( .A1(n2980), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3278), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4211) );
  AOI22_X1 U5218 ( .A1(n4231), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4210) );
  AOI22_X1 U5219 ( .A1(n2970), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4209) );
  AOI22_X1 U5220 ( .A1(n4240), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3183), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4208) );
  NAND4_X1 U5221 ( .A1(n4211), .A2(n4210), .A3(n4209), .A4(n4208), .ZN(n4217)
         );
  AOI22_X1 U5222 ( .A1(n4238), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4215) );
  AOI22_X1 U5223 ( .A1(n4069), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4214) );
  AOI22_X1 U5224 ( .A1(n3218), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4213) );
  AOI22_X1 U5225 ( .A1(n4229), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4212) );
  NAND4_X1 U5226 ( .A1(n4215), .A2(n4214), .A3(n4213), .A4(n4212), .ZN(n4216)
         );
  OR2_X1 U5227 ( .A1(n4217), .A2(n4216), .ZN(n4247) );
  INV_X1 U5228 ( .A(n4247), .ZN(n4218) );
  XNOR2_X1 U5229 ( .A(n4248), .B(n4218), .ZN(n4222) );
  INV_X1 U5230 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4220) );
  NAND2_X1 U5231 ( .A1(n6601), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4219)
         );
  OAI211_X1 U5232 ( .C1(n4254), .C2(n4220), .A(n4251), .B(n4219), .ZN(n4221)
         );
  AOI21_X1 U5233 ( .B1(n4222), .B2(n4256), .A(n4221), .ZN(n4227) );
  OR2_X1 U5234 ( .A1(n4224), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4225)
         );
  NAND2_X1 U5235 ( .A1(n4322), .A2(n4225), .ZN(n5503) );
  NOR2_X1 U5236 ( .A1(n5503), .A2(n4251), .ZN(n4226) );
  AOI22_X1 U5237 ( .A1(n4229), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4228), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4236) );
  AOI22_X1 U5238 ( .A1(n4231), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4230), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4235) );
  AOI22_X1 U5239 ( .A1(n3278), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4232), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4234) );
  AOI22_X1 U5240 ( .A1(n4069), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3895), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4233) );
  NAND4_X1 U5241 ( .A1(n4236), .A2(n4235), .A3(n4234), .A4(n4233), .ZN(n4246)
         );
  AOI22_X1 U5242 ( .A1(n2969), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4244) );
  AOI22_X1 U5243 ( .A1(n4238), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4188), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4243) );
  AOI22_X1 U5244 ( .A1(n2968), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4242) );
  AOI22_X1 U5245 ( .A1(n4240), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n2979), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4241) );
  NAND4_X1 U5246 ( .A1(n4244), .A2(n4243), .A3(n4242), .A4(n4241), .ZN(n4245)
         );
  NOR2_X1 U5247 ( .A1(n4246), .A2(n4245), .ZN(n4250) );
  NAND2_X1 U5248 ( .A1(n4248), .A2(n4247), .ZN(n4249) );
  XOR2_X1 U5249 ( .A(n4250), .B(n4249), .Z(n4257) );
  INV_X1 U5250 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4253) );
  NAND2_X1 U5251 ( .A1(n6601), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4252)
         );
  OAI211_X1 U5252 ( .C1(n4254), .C2(n4253), .A(n4252), .B(n4251), .ZN(n4255)
         );
  AOI21_X1 U5253 ( .B1(n4257), .B2(n4256), .A(n4255), .ZN(n4258) );
  INV_X1 U5254 ( .A(n4258), .ZN(n4260) );
  XNOR2_X1 U5255 ( .A(n4322), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5341)
         );
  NAND2_X1 U5256 ( .A1(n5341), .A2(n4339), .ZN(n4259) );
  INV_X1 U5257 ( .A(n5327), .ZN(n5348) );
  NAND2_X1 U5258 ( .A1(n3227), .A2(n6491), .ZN(n4261) );
  OR2_X2 U5259 ( .A1(n4365), .A2(n4261), .ZN(n6097) );
  NOR2_X1 U5260 ( .A1(n4309), .A2(n4271), .ZN(n4516) );
  NAND2_X1 U5261 ( .A1(n6468), .A2(n4516), .ZN(n4264) );
  OR2_X1 U5262 ( .A1(n3616), .A2(n4262), .ZN(n4263) );
  NAND2_X1 U5263 ( .A1(n4264), .A2(n4263), .ZN(n4407) );
  INV_X1 U5264 ( .A(n4265), .ZN(n6467) );
  NAND3_X1 U5265 ( .A1(n3755), .A2(n6467), .A3(n3167), .ZN(n4267) );
  NOR2_X1 U5266 ( .A1(n4267), .A2(n4266), .ZN(n4270) );
  INV_X1 U5267 ( .A(n4268), .ZN(n4269) );
  NAND2_X1 U5268 ( .A1(n4270), .A2(n4269), .ZN(n4282) );
  NOR2_X1 U5269 ( .A1(n4282), .A2(n4271), .ZN(n4272) );
  AND2_X1 U5270 ( .A1(n4575), .A2(n4275), .ZN(n4278) );
  NOR2_X1 U5271 ( .A1(n4278), .A2(n4277), .ZN(n4276) );
  AOI22_X1 U5272 ( .A1(n6005), .A2(DATAI_30_), .B1(n6008), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n4280) );
  NAND2_X1 U5273 ( .A1(n6009), .A2(DATAI_14_), .ZN(n4279) );
  OAI21_X1 U5274 ( .B1(n5348), .B2(n5499), .A(n3094), .ZN(U2861) );
  OR2_X1 U5275 ( .A1(n4518), .A2(n6474), .ZN(n4281) );
  OR2_X1 U5276 ( .A1(n6468), .A2(n4281), .ZN(n4284) );
  OR2_X1 U5277 ( .A1(n4282), .A2(n4297), .ZN(n4283) );
  INV_X1 U5278 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5336) );
  AOI21_X1 U5279 ( .B1(n5327), .B2(n4286), .A(n4285), .ZN(n4287) );
  INV_X1 U5280 ( .A(n4287), .ZN(U2829) );
  NAND2_X1 U5281 ( .A1(n3535), .A2(n5586), .ZN(n4288) );
  NOR2_X1 U5282 ( .A1(n4289), .A2(n4288), .ZN(n4290) );
  AOI21_X1 U5283 ( .B1(n4291), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n4290), 
        .ZN(n4292) );
  INV_X1 U5284 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5349) );
  MUX2_X1 U5285 ( .A(n4293), .B(EBX_REG_29__SCAN_IN), .S(n2983), .Z(n5371) );
  NOR3_X1 U5286 ( .A1(n5385), .A2(n5371), .A3(n4294), .ZN(n4295) );
  NOR2_X1 U5287 ( .A1(n4296), .A2(n4295), .ZN(n4299) );
  OAI22_X1 U5288 ( .A1(n3654), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4297), .ZN(n4298) );
  INV_X1 U5289 ( .A(n6213), .ZN(n4302) );
  NAND2_X1 U5290 ( .A1(n2971), .A2(REIP_REG_31__SCAN_IN), .ZN(n4326) );
  INV_X1 U5291 ( .A(n4326), .ZN(n4301) );
  AOI211_X2 U5292 ( .C1(n5454), .C2(n4302), .A(n4301), .B(n3098), .ZN(n4306)
         );
  OAI21_X1 U5293 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5686), .A(n4303), 
        .ZN(n4304) );
  NAND2_X1 U5294 ( .A1(n4304), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4305) );
  OAI211_X1 U5295 ( .C1(n4307), .C2(n6198), .A(n4306), .B(n4305), .ZN(U2987)
         );
  OR2_X1 U5296 ( .A1(n4309), .A2(n4308), .ZN(n6454) );
  OR2_X2 U5297 ( .A1(n6043), .A2(n6454), .ZN(n6137) );
  NAND2_X1 U5298 ( .A1(n4311), .A2(n2997), .ZN(n4316) );
  AOI22_X1 U5299 ( .A1(n4313), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n4312), .ZN(n4314) );
  INV_X1 U5300 ( .A(n4314), .ZN(n4315) );
  NAND3_X1 U5301 ( .A1(n6603), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6482) );
  AND2_X1 U5302 ( .A1(n4317), .A2(n6364), .ZN(n6599) );
  INV_X1 U5303 ( .A(n6599), .ZN(n4318) );
  NAND2_X1 U5304 ( .A1(n4318), .A2(n6603), .ZN(n4319) );
  NAND2_X1 U5305 ( .A1(n6603), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4321) );
  NAND2_X1 U5306 ( .A1(n6602), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4320) );
  NAND2_X1 U5307 ( .A1(n4321), .A2(n4320), .ZN(n4388) );
  INV_X1 U5308 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5325) );
  INV_X1 U5309 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4323) );
  NAND2_X1 U5310 ( .A1(n6142), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4325)
         );
  OAI211_X1 U5311 ( .C1(n6139), .C2(n4343), .A(n4326), .B(n4325), .ZN(n4327)
         );
  NAND2_X1 U5312 ( .A1(n2976), .A2(n4329), .ZN(n4331) );
  AOI22_X1 U5313 ( .A1(n6005), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6008), .ZN(n4330) );
  NAND2_X1 U5314 ( .A1(n4331), .A2(n4330), .ZN(U2860) );
  INV_X1 U5315 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6721) );
  INV_X1 U5316 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U5317 ( .A1(n2978), .A2(n4376), .ZN(n4368) );
  INV_X1 U5318 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6587) );
  INV_X1 U5319 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6505) );
  INV_X1 U5320 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6503) );
  NOR3_X1 U5321 ( .A1(n6587), .A2(n6505), .A3(n6503), .ZN(n5971) );
  NAND2_X1 U5322 ( .A1(REIP_REG_4__SCAN_IN), .A2(n5971), .ZN(n4358) );
  NOR2_X2 U5323 ( .A1(n6509), .A2(n5953), .ZN(n5936) );
  INV_X1 U5324 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6513) );
  NOR3_X1 U5325 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6721), .A3(n5190), .ZN(n4363) );
  NOR2_X1 U5326 ( .A1(n4336), .A2(n4337), .ZN(n4338) );
  OR2_X1 U5327 ( .A1(n4335), .A2(n4338), .ZN(n5112) );
  NOR2_X1 U5328 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6607) );
  NAND2_X1 U5329 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6607), .ZN(n6471) );
  NAND3_X1 U5330 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n4339), .A3(n6603), .ZN(
        n6478) );
  OAI211_X1 U5331 ( .C1(n6603), .C2(n6471), .A(n6598), .B(n6478), .ZN(n4340)
         );
  INV_X1 U5332 ( .A(n4340), .ZN(n4341) );
  NOR2_X1 U5333 ( .A1(n4343), .A2(n6634), .ZN(n4342) );
  NOR2_X1 U5334 ( .A1(n5112), .A2(n5946), .ZN(n4362) );
  NAND2_X1 U5335 ( .A1(n6491), .A2(n6602), .ZN(n4345) );
  AND2_X1 U5336 ( .A1(n2981), .A2(n4345), .ZN(n4354) );
  AND2_X1 U5337 ( .A1(EBX_REG_31__SCAN_IN), .A2(n5357), .ZN(n4346) );
  AND2_X1 U5338 ( .A1(n3227), .A2(n4346), .ZN(n4347) );
  OAI21_X1 U5339 ( .B1(n4348), .B2(n4912), .A(n4349), .ZN(n4350) );
  AND2_X1 U5340 ( .A1(n4350), .A2(n5055), .ZN(n5124) );
  AOI22_X1 U5341 ( .A1(n5968), .A2(n5111), .B1(n5961), .B2(n5124), .ZN(n4351)
         );
  OAI211_X1 U5342 ( .C1(n5963), .C2(n4352), .A(n4351), .B(n3095), .ZN(n4361)
         );
  INV_X1 U5343 ( .A(n6490), .ZN(n4353) );
  NAND3_X1 U5344 ( .A1(n6491), .A2(n6602), .A3(n4353), .ZN(n6464) );
  NAND2_X1 U5345 ( .A1(n2984), .A2(n6464), .ZN(n4356) );
  INV_X1 U5346 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U5347 ( .A1(n4354), .A2(n5455), .ZN(n4355) );
  NAND2_X1 U5348 ( .A1(n4356), .A2(n4355), .ZN(n4357) );
  NAND2_X1 U5349 ( .A1(n5015), .A2(n5977), .ZN(n5423) );
  INV_X1 U5350 ( .A(n5015), .ZN(n5090) );
  NOR3_X1 U5351 ( .A1(n5090), .A2(n6509), .A3(n4358), .ZN(n5941) );
  NAND4_X1 U5352 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .A4(n5941), .ZN(n5076) );
  AND2_X1 U5353 ( .A1(n5423), .A2(n5076), .ZN(n5099) );
  NOR2_X1 U5354 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5190), .ZN(n5095) );
  OAI21_X1 U5355 ( .B1(n5099), .B2(n5095), .A(REIP_REG_10__SCAN_IN), .ZN(n4359) );
  OAI21_X1 U5356 ( .B1(n5981), .B2(n4999), .A(n4359), .ZN(n4360) );
  OR4_X1 U5357 ( .A1(n4363), .A2(n4362), .A3(n4361), .A4(n4360), .ZN(U2817) );
  INV_X1 U5358 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n4366) );
  INV_X1 U5359 ( .A(n4384), .ZN(n4364) );
  OAI211_X1 U5360 ( .C1(n4367), .C2(n4366), .A(n4365), .B(n4364), .ZN(U2788)
         );
  OR2_X1 U5361 ( .A1(n6468), .A2(n5001), .ZN(n4370) );
  NAND2_X1 U5362 ( .A1(n4368), .A2(n4373), .ZN(n4369) );
  NAND2_X1 U5363 ( .A1(n4370), .A2(n4369), .ZN(n5869) );
  OR2_X1 U5364 ( .A1(n2984), .A2(n4371), .ZN(n4386) );
  AOI21_X1 U5365 ( .B1(n4386), .B2(n6490), .A(READY_N), .ZN(n6605) );
  NOR2_X1 U5366 ( .A1(n5869), .A2(n6605), .ZN(n6452) );
  OR2_X1 U5367 ( .A1(n6452), .A2(n6474), .ZN(n4381) );
  INV_X1 U5368 ( .A(n4381), .ZN(n5875) );
  INV_X1 U5369 ( .A(MORE_REG_SCAN_IN), .ZN(n4383) );
  AND2_X1 U5370 ( .A1(n4373), .A2(n4372), .ZN(n4374) );
  OR2_X1 U5371 ( .A1(n6468), .A2(n4374), .ZN(n4380) );
  NAND2_X1 U5372 ( .A1(n6468), .A2(n4375), .ZN(n4379) );
  INV_X1 U5373 ( .A(n4376), .ZN(n4377) );
  NAND2_X1 U5374 ( .A1(n2978), .A2(n4377), .ZN(n4378) );
  AND3_X1 U5375 ( .A1(n4380), .A2(n4379), .A3(n4378), .ZN(n6455) );
  OR2_X1 U5376 ( .A1(n4381), .A2(n6455), .ZN(n4382) );
  OAI21_X1 U5377 ( .B1(n5875), .B2(n4383), .A(n4382), .ZN(U3471) );
  OAI21_X1 U5378 ( .B1(n4384), .B2(READREQUEST_REG_SCAN_IN), .A(n6598), .ZN(
        n4385) );
  OAI21_X1 U5379 ( .B1(n6598), .B2(n4386), .A(n4385), .ZN(U3474) );
  XOR2_X1 U5380 ( .A(n4387), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n5701) );
  INV_X1 U5381 ( .A(n5701), .ZN(n4396) );
  OAI21_X1 U5382 ( .B1(n6142), .B2(n4388), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4395) );
  INV_X1 U5383 ( .A(n4389), .ZN(n4392) );
  OAI21_X1 U5384 ( .B1(n4392), .B2(n4391), .A(n4390), .ZN(n5008) );
  INV_X1 U5385 ( .A(n5008), .ZN(n4393) );
  AOI22_X1 U5386 ( .A1(n4393), .A2(n6133), .B1(n2971), .B2(REIP_REG_0__SCAN_IN), .ZN(n4394) );
  OAI211_X1 U5387 ( .C1(n4396), .C2(n6137), .A(n4395), .B(n4394), .ZN(U2986)
         );
  INV_X1 U5388 ( .A(n4397), .ZN(n4398) );
  OAI21_X1 U5389 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n3654), .A(n4398), 
        .ZN(n5699) );
  OAI222_X1 U5390 ( .A1(n5008), .A2(n5480), .B1(n5997), .B2(n4399), .C1(n5699), 
        .C2(n5773), .ZN(U2859) );
  NOR2_X1 U5391 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6718), .ZN(n6565) );
  AOI21_X1 U5392 ( .B1(n4400), .B2(n6490), .A(READY_N), .ZN(n4401) );
  OAI211_X1 U5393 ( .C1(n3608), .C2(n6434), .A(n6468), .B(n4401), .ZN(n4405)
         );
  INV_X1 U5394 ( .A(n4402), .ZN(n4403) );
  NAND3_X1 U5395 ( .A1(n4405), .A2(n4404), .A3(n4403), .ZN(n4408) );
  NOR2_X1 U5396 ( .A1(n6468), .A2(n4518), .ZN(n4406) );
  INV_X1 U5397 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5874) );
  NOR2_X1 U5398 ( .A1(n6634), .A2(n6601), .ZN(n6473) );
  NAND2_X1 U5399 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6473), .ZN(n6566) );
  OAI22_X1 U5400 ( .A1(n6436), .A2(n6474), .B1(n5874), .B2(n6566), .ZN(n4411)
         );
  NOR2_X1 U5401 ( .A1(n6565), .A2(n4411), .ZN(n6583) );
  INV_X1 U5402 ( .A(n6583), .ZN(n6581) );
  INV_X1 U5403 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6613) );
  INV_X1 U5404 ( .A(n4409), .ZN(n4733) );
  OR2_X1 U5405 ( .A1(n3397), .A2(n4733), .ZN(n4410) );
  XNOR2_X1 U5406 ( .A(n4410), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5962)
         );
  INV_X1 U5407 ( .A(n6586), .ZN(n6571) );
  INV_X1 U5408 ( .A(n3616), .ZN(n4539) );
  NAND4_X1 U5409 ( .A1(n5962), .A2(n6571), .A3(n4539), .A4(n4411), .ZN(n4412)
         );
  OAI21_X1 U5410 ( .B1(n6581), .B2(n6613), .A(n4412), .ZN(U3455) );
  OR2_X1 U5411 ( .A1(n4414), .A2(n4413), .ZN(n4415) );
  NAND2_X1 U5412 ( .A1(n4416), .A2(n4415), .ZN(n6144) );
  XNOR2_X1 U5413 ( .A(n4417), .B(n4418), .ZN(n4483) );
  INV_X1 U5414 ( .A(n5997), .ZN(n5490) );
  AOI22_X1 U5415 ( .A1(n5995), .A2(n4483), .B1(n5490), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4419) );
  OAI21_X1 U5416 ( .B1(n5480), .B2(n6144), .A(n4419), .ZN(U2858) );
  XNOR2_X1 U5417 ( .A(n4586), .B(n4420), .ZN(n6123) );
  OR2_X1 U5418 ( .A1(n4570), .A2(n4421), .ZN(n4422) );
  AND2_X1 U5419 ( .A1(n4593), .A2(n4422), .ZN(n6197) );
  AOI22_X1 U5420 ( .A1(n5995), .A2(n6197), .B1(n5490), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4423) );
  OAI21_X1 U5421 ( .B1(n6123), .B2(n5480), .A(n4423), .ZN(U2856) );
  AND2_X1 U5422 ( .A1(n4924), .A2(n3763), .ZN(n6358) );
  INV_X1 U5423 ( .A(n4427), .ZN(n5715) );
  OR2_X1 U5424 ( .A1(n4426), .A2(n5715), .ZN(n4824) );
  INV_X1 U5425 ( .A(n4824), .ZN(n6303) );
  INV_X1 U5426 ( .A(n4726), .ZN(n6419) );
  AOI21_X1 U5427 ( .B1(n6358), .B2(n6303), .A(n6419), .ZN(n4433) );
  INV_X1 U5428 ( .A(n4436), .ZN(n4821) );
  OAI22_X1 U5429 ( .A1(n4433), .A2(n6364), .B1(n6601), .B2(n4821), .ZN(n6420)
         );
  INV_X1 U5430 ( .A(n6420), .ZN(n4725) );
  INV_X1 U5431 ( .A(DATAI_7_), .ZN(n6080) );
  INV_X1 U5432 ( .A(DATAI_31_), .ZN(n4428) );
  NOR2_X1 U5433 ( .A1(n6145), .A2(n4428), .ZN(n6412) );
  INV_X1 U5434 ( .A(n4932), .ZN(n6261) );
  NOR2_X1 U5435 ( .A1(n4609), .A2(n3755), .ZN(n6410) );
  INV_X1 U5436 ( .A(n6410), .ZN(n6780) );
  NAND2_X1 U5437 ( .A1(n6133), .A2(DATAI_23_), .ZN(n6301) );
  NAND2_X1 U5438 ( .A1(n5707), .A2(n4494), .ZN(n4676) );
  OAI22_X1 U5439 ( .A1(n6780), .A2(n4726), .B1(n6301), .B2(n6423), .ZN(n4431)
         );
  AOI21_X1 U5440 ( .B1(n6412), .B2(n6782), .A(n4431), .ZN(n4438) );
  INV_X1 U5441 ( .A(n6364), .ZN(n6312) );
  INV_X1 U5442 ( .A(n4822), .ZN(n4432) );
  AOI21_X1 U5443 ( .B1(n4432), .B2(n5707), .A(n6145), .ZN(n4434) );
  OR2_X1 U5444 ( .A1(n6364), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5138) );
  INV_X1 U5445 ( .A(n5138), .ZN(n4868) );
  OAI21_X1 U5446 ( .B1(n4434), .B2(n4868), .A(n4433), .ZN(n4435) );
  INV_X1 U5447 ( .A(n6362), .ZN(n6310) );
  OAI211_X1 U5448 ( .C1(n4436), .C2(n6312), .A(n4435), .B(n6310), .ZN(n6417)
         );
  NAND2_X1 U5449 ( .A1(n6417), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4437)
         );
  OAI211_X1 U5450 ( .C1(n4725), .C2(n6786), .A(n4438), .B(n4437), .ZN(U3147)
         );
  INV_X1 U5451 ( .A(n6463), .ZN(n4439) );
  NOR2_X1 U5452 ( .A1(n6434), .A2(n4439), .ZN(n4440) );
  NAND2_X1 U5453 ( .A1(n6040), .A2(n2982), .ZN(n6012) );
  NAND2_X1 U5454 ( .A1(n6473), .A2(n6603), .ZN(n6600) );
  NOR2_X4 U5455 ( .A1(n6040), .A2(n6036), .ZN(n6032) );
  AOI22_X1 U5456 ( .A1(n6036), .A2(UWORD_REG_14__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4442) );
  OAI21_X1 U5457 ( .B1(n4253), .B2(n6012), .A(n4442), .ZN(U2893) );
  AOI22_X1 U5458 ( .A1(n6036), .A2(UWORD_REG_11__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4443) );
  OAI21_X1 U5459 ( .B1(n4178), .B2(n6012), .A(n4443), .ZN(U2896) );
  INV_X1 U5460 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4445) );
  AOI22_X1 U5461 ( .A1(n6036), .A2(UWORD_REG_1__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4444) );
  OAI21_X1 U5462 ( .B1(n4445), .B2(n6012), .A(n4444), .ZN(U2906) );
  INV_X1 U5463 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6710) );
  AOI22_X1 U5464 ( .A1(n6036), .A2(UWORD_REG_2__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4446) );
  OAI21_X1 U5465 ( .B1(n6710), .B2(n6012), .A(n4446), .ZN(U2905) );
  INV_X1 U5466 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4448) );
  AOI22_X1 U5467 ( .A1(n6036), .A2(UWORD_REG_3__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4447) );
  OAI21_X1 U5468 ( .B1(n4448), .B2(n6012), .A(n4447), .ZN(U2904) );
  INV_X1 U5469 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4450) );
  AOI22_X1 U5470 ( .A1(n6036), .A2(UWORD_REG_5__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4449) );
  OAI21_X1 U5471 ( .B1(n4450), .B2(n6012), .A(n4449), .ZN(U2902) );
  INV_X1 U5472 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4452) );
  AOI22_X1 U5473 ( .A1(n6036), .A2(UWORD_REG_6__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4451) );
  OAI21_X1 U5474 ( .B1(n4452), .B2(n6012), .A(n4451), .ZN(U2901) );
  INV_X1 U5475 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4454) );
  AOI22_X1 U5476 ( .A1(n6036), .A2(UWORD_REG_7__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4453) );
  OAI21_X1 U5477 ( .B1(n4454), .B2(n6012), .A(n4453), .ZN(U2900) );
  AOI22_X1 U5478 ( .A1(n6036), .A2(UWORD_REG_8__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4455) );
  OAI21_X1 U5479 ( .B1(n4117), .B2(n6012), .A(n4455), .ZN(U2899) );
  AOI22_X1 U5480 ( .A1(n6036), .A2(UWORD_REG_13__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4456) );
  OAI21_X1 U5481 ( .B1(n4220), .B2(n6012), .A(n4456), .ZN(U2894) );
  INV_X1 U5482 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6057) );
  AOI22_X1 U5483 ( .A1(n6036), .A2(UWORD_REG_10__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4457) );
  OAI21_X1 U5484 ( .B1(n6057), .B2(n6012), .A(n4457), .ZN(U2897) );
  INV_X1 U5485 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6062) );
  AOI22_X1 U5486 ( .A1(n6036), .A2(UWORD_REG_12__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4458) );
  OAI21_X1 U5487 ( .B1(n6062), .B2(n6012), .A(n4458), .ZN(U2895) );
  INV_X1 U5488 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4460) );
  AOI22_X1 U5489 ( .A1(n6036), .A2(UWORD_REG_0__SCAN_IN), .B1(
        DATAO_REG_16__SCAN_IN), .B2(n6032), .ZN(n4459) );
  OAI21_X1 U5490 ( .B1(n4460), .B2(n6012), .A(n4459), .ZN(U2907) );
  INV_X1 U5491 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4462) );
  AOI22_X1 U5492 ( .A1(n6036), .A2(UWORD_REG_9__SCAN_IN), .B1(
        DATAO_REG_25__SCAN_IN), .B2(n6032), .ZN(n4461) );
  OAI21_X1 U5493 ( .B1(n4462), .B2(n6012), .A(n4461), .ZN(U2898) );
  NAND2_X1 U5494 ( .A1(n5707), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5710) );
  OAI21_X1 U5495 ( .B1(n4622), .B2(n5710), .A(n6312), .ZN(n4469) );
  AND2_X1 U5496 ( .A1(n2975), .A2(n4426), .ZN(n4923) );
  NAND2_X1 U5497 ( .A1(n4923), .A2(n4924), .ZN(n4781) );
  INV_X1 U5498 ( .A(n3763), .ZN(n6224) );
  OR2_X1 U5499 ( .A1(n4781), .A2(n6224), .ZN(n4465) );
  OR2_X1 U5500 ( .A1(n4919), .A2(n6446), .ZN(n4775) );
  NOR2_X1 U5501 ( .A1(n6356), .A2(n4775), .ZN(n6348) );
  INV_X1 U5502 ( .A(n6348), .ZN(n4464) );
  NAND2_X1 U5503 ( .A1(n4465), .A2(n4464), .ZN(n4467) );
  NAND2_X1 U5504 ( .A1(n4775), .A2(n6364), .ZN(n4466) );
  OAI211_X1 U5505 ( .C1(n4469), .C2(n4467), .A(n6310), .B(n4466), .ZN(n6351)
         );
  INV_X1 U5506 ( .A(n6351), .ZN(n4580) );
  INV_X1 U5507 ( .A(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4478) );
  INV_X1 U5508 ( .A(DATAI_0_), .ZN(n6067) );
  INV_X1 U5509 ( .A(n4467), .ZN(n4468) );
  OR2_X1 U5510 ( .A1(n4469), .A2(n4468), .ZN(n4472) );
  INV_X1 U5511 ( .A(n4775), .ZN(n4470) );
  NAND2_X1 U5512 ( .A1(n4470), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4471) );
  NAND2_X1 U5513 ( .A1(n4472), .A2(n4471), .ZN(n6349) );
  INV_X1 U5514 ( .A(DATAI_24_), .ZN(n4473) );
  NOR2_X1 U5515 ( .A1(n6145), .A2(n4473), .ZN(n6368) );
  INV_X1 U5516 ( .A(n6368), .ZN(n6425) );
  NOR2_X2 U5517 ( .A1(n4609), .A2(n4474), .ZN(n6418) );
  NOR2_X2 U5518 ( .A1(n4622), .A2(n4676), .ZN(n6347) );
  NAND2_X1 U5519 ( .A1(n6133), .A2(DATAI_16_), .ZN(n6422) );
  INV_X1 U5520 ( .A(n6422), .ZN(n6360) );
  AOI22_X1 U5521 ( .A1(n6418), .A2(n6348), .B1(n6347), .B2(n6360), .ZN(n4475)
         );
  OAI21_X1 U5522 ( .B1(n6354), .B2(n6425), .A(n4475), .ZN(n4476) );
  AOI21_X1 U5523 ( .B1(n6421), .B2(n6349), .A(n4476), .ZN(n4477) );
  OAI21_X1 U5524 ( .B1(n4580), .B2(n4478), .A(n4477), .ZN(U3108) );
  XNOR2_X1 U5525 ( .A(n4480), .B(n4479), .ZN(n6138) );
  OR3_X1 U5526 ( .A1(n5686), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4481), 
        .ZN(n4485) );
  NOR2_X1 U5527 ( .A1(n6215), .A2(n5681), .ZN(n4482) );
  NOR2_X1 U5528 ( .A1(n3095), .A2(n6587), .ZN(n6141) );
  AOI211_X1 U5529 ( .C1(n4302), .C2(n4483), .A(n4482), .B(n6141), .ZN(n4484)
         );
  OAI211_X1 U5530 ( .C1(n6138), .C2(n6198), .A(n4485), .B(n4484), .ZN(U3017)
         );
  NOR2_X1 U5531 ( .A1(n4426), .A2(n2975), .ZN(n6357) );
  INV_X1 U5532 ( .A(n6357), .ZN(n4732) );
  NOR2_X1 U5533 ( .A1(n4732), .A2(n6364), .ZN(n4741) );
  INV_X1 U5534 ( .A(n4924), .ZN(n6304) );
  NAND2_X1 U5535 ( .A1(n4741), .A2(n6304), .ZN(n4487) );
  AND2_X1 U5536 ( .A1(n4488), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6262) );
  NOR2_X1 U5537 ( .A1(n5144), .A2(n4681), .ZN(n4872) );
  NAND2_X1 U5538 ( .A1(n6262), .A2(n4872), .ZN(n4486) );
  NAND2_X1 U5539 ( .A1(n4487), .A2(n4486), .ZN(n4610) );
  INV_X1 U5540 ( .A(n4610), .ZN(n4663) );
  NAND2_X1 U5541 ( .A1(n4730), .A2(n6446), .ZN(n6231) );
  NOR2_X1 U5542 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6231), .ZN(n4611)
         );
  INV_X1 U5543 ( .A(n4611), .ZN(n4658) );
  NOR2_X1 U5544 ( .A1(n4488), .A2(n6601), .ZN(n6267) );
  OAI21_X1 U5545 ( .B1(n4872), .B2(n6601), .A(n4771), .ZN(n4864) );
  AOI211_X1 U5546 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4658), .A(n6267), .B(
        n4864), .ZN(n4493) );
  NAND2_X1 U5547 ( .A1(n3779), .A2(n4429), .ZN(n4931) );
  INV_X1 U5548 ( .A(n6260), .ZN(n4491) );
  INV_X1 U5549 ( .A(n4621), .ZN(n4490) );
  AOI21_X1 U5550 ( .B1(n4491), .B2(n4490), .A(n6364), .ZN(n6230) );
  NAND2_X1 U5551 ( .A1(n6357), .A2(n4733), .ZN(n6225) );
  OAI211_X1 U5552 ( .C1(n4868), .C2(n4964), .A(n6230), .B(n6225), .ZN(n4492)
         );
  NAND2_X1 U5553 ( .A1(n4493), .A2(n4492), .ZN(n4657) );
  NAND2_X1 U5554 ( .A1(n4657), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4497) );
  OAI22_X1 U5555 ( .A1(n6780), .A2(n4658), .B1(n6301), .B2(n6234), .ZN(n4495)
         );
  AOI21_X1 U5556 ( .B1(n6412), .B2(n4660), .A(n4495), .ZN(n4496) );
  OAI211_X1 U5557 ( .C1(n4663), .C2(n6786), .A(n4497), .B(n4496), .ZN(U3059)
         );
  INV_X1 U5558 ( .A(n6421), .ZN(n6371) );
  NAND2_X1 U5559 ( .A1(n4657), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4500) );
  INV_X1 U5560 ( .A(n6418), .ZN(n5179) );
  OAI22_X1 U5561 ( .A1(n5179), .A2(n4658), .B1(n6422), .B2(n6234), .ZN(n4498)
         );
  AOI21_X1 U5562 ( .B1(n6368), .B2(n4660), .A(n4498), .ZN(n4499) );
  OAI211_X1 U5563 ( .C1(n4663), .C2(n6371), .A(n4500), .B(n4499), .ZN(U3052)
         );
  NAND2_X1 U5564 ( .A1(n6133), .A2(DATAI_26_), .ZN(n6342) );
  NAND2_X1 U5565 ( .A1(n6133), .A2(DATAI_18_), .ZN(n6278) );
  INV_X1 U5566 ( .A(n6278), .ZN(n6378) );
  NOR2_X2 U5567 ( .A1(n4609), .A2(n3611), .ZN(n6379) );
  INV_X1 U5568 ( .A(n6379), .ZN(n5162) );
  INV_X1 U5569 ( .A(DATAI_2_), .ZN(n6071) );
  NOR2_X1 U5570 ( .A1(n6071), .A2(n4683), .ZN(n6339) );
  INV_X1 U5571 ( .A(n6339), .ZN(n6383) );
  OAI22_X1 U5572 ( .A1(n5162), .A2(n4726), .B1(n4725), .B2(n6383), .ZN(n4501)
         );
  AOI21_X1 U5573 ( .B1(n6378), .B2(n4905), .A(n4501), .ZN(n4503) );
  NAND2_X1 U5574 ( .A1(n6417), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4502)
         );
  OAI211_X1 U5575 ( .C1(n6424), .C2(n6342), .A(n4503), .B(n4502), .ZN(U3142)
         );
  NAND2_X1 U5576 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5874), .ZN(n4537) );
  INV_X1 U5577 ( .A(n4504), .ZN(n4536) );
  INV_X1 U5578 ( .A(n3608), .ZN(n4507) );
  INV_X1 U5579 ( .A(n4505), .ZN(n4506) );
  NAND4_X1 U5580 ( .A1(n4508), .A2(n3616), .A3(n4507), .A4(n4506), .ZN(n4510)
         );
  NOR2_X1 U5581 ( .A1(n4510), .A2(n4509), .ZN(n6430) );
  XNOR2_X1 U5582 ( .A(n4511), .B(n4521), .ZN(n4515) );
  INV_X1 U5583 ( .A(n4528), .ZN(n4514) );
  INV_X1 U5584 ( .A(n4512), .ZN(n4520) );
  OAI21_X1 U5585 ( .B1(n4520), .B2(n3771), .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .ZN(n4513) );
  NAND2_X1 U5586 ( .A1(n3364), .A2(n4513), .ZN(n6570) );
  AOI22_X1 U5587 ( .A1(n6434), .A2(n4515), .B1(n4514), .B2(n6570), .ZN(n4525)
         );
  INV_X1 U5588 ( .A(n4516), .ZN(n4517) );
  NAND2_X1 U5589 ( .A1(n4518), .A2(n4517), .ZN(n4531) );
  INV_X1 U5590 ( .A(n4519), .ZN(n4522) );
  INV_X1 U5591 ( .A(n4520), .ZN(n5714) );
  MUX2_X1 U5592 ( .A(n4522), .B(n4521), .S(n5714), .Z(n4523) );
  NAND3_X1 U5593 ( .A1(n4531), .A2(n4536), .A3(n4523), .ZN(n4524) );
  OAI211_X1 U5594 ( .C1(n6304), .C2(n6430), .A(n4525), .B(n4524), .ZN(n6572)
         );
  MUX2_X1 U5595 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6572), .S(n4534), 
        .Z(n6447) );
  OR2_X1 U5596 ( .A1(n4426), .A2(n6430), .ZN(n4533) );
  XNOR2_X1 U5597 ( .A(n5714), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4530)
         );
  XNOR2_X1 U5598 ( .A(n3771), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4526)
         );
  NAND2_X1 U5599 ( .A1(n6434), .A2(n4526), .ZN(n4527) );
  OAI21_X1 U5600 ( .B1(n4530), .B2(n4528), .A(n4527), .ZN(n4529) );
  AOI21_X1 U5601 ( .B1(n4531), .B2(n4530), .A(n4529), .ZN(n4532) );
  NAND2_X1 U5602 ( .A1(n4533), .A2(n4532), .ZN(n5353) );
  MUX2_X1 U5603 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n5353), .S(n4534), 
        .Z(n6441) );
  NAND3_X1 U5604 ( .A1(n6447), .A2(n6441), .A3(n6634), .ZN(n4535) );
  OAI21_X1 U5605 ( .B1(n4537), .B2(n4536), .A(n4535), .ZN(n6458) );
  INV_X1 U5606 ( .A(n4538), .ZN(n5719) );
  NAND2_X1 U5607 ( .A1(n6458), .A2(n5719), .ZN(n4543) );
  MUX2_X1 U5608 ( .A(n6436), .B(n5874), .S(STATE2_REG_1__SCAN_IN), .Z(n4541)
         );
  AND3_X1 U5609 ( .A1(n5962), .A2(n4539), .A3(n6634), .ZN(n4540) );
  AOI21_X1 U5610 ( .B1(n4541), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n4540), 
        .ZN(n6456) );
  AND3_X1 U5611 ( .A1(n4543), .A2(n5874), .A3(n6456), .ZN(n4542) );
  OAI21_X1 U5612 ( .B1(n4542), .B2(n6566), .A(n4683), .ZN(n6223) );
  AND3_X1 U5613 ( .A1(n4543), .A2(n6456), .A3(n6473), .ZN(n6465) );
  AND2_X1 U5614 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6718), .ZN(n5711) );
  OAI22_X1 U5615 ( .A1(n5028), .A2(n6364), .B1(n6224), .B2(n5711), .ZN(n4544)
         );
  OAI21_X1 U5616 ( .B1(n6465), .B2(n4544), .A(n6223), .ZN(n4545) );
  OAI21_X1 U5617 ( .B1(n6223), .B2(n6356), .A(n4545), .ZN(U3465) );
  NOR2_X1 U5618 ( .A1(n4822), .A2(n4621), .ZN(n6355) );
  INV_X1 U5619 ( .A(n6355), .ZN(n4547) );
  OR2_X1 U5620 ( .A1(n6260), .A2(n5710), .ZN(n6302) );
  AND2_X1 U5621 ( .A1(n4622), .A2(n6302), .ZN(n4546) );
  AOI21_X1 U5622 ( .B1(n4547), .B2(n4546), .A(n6364), .ZN(n4922) );
  OAI22_X1 U5623 ( .A1(n3779), .A2(n5138), .B1(n6304), .B2(n5711), .ZN(n4548)
         );
  OAI21_X1 U5624 ( .B1(n4922), .B2(n4548), .A(n6223), .ZN(n4549) );
  OAI21_X1 U5625 ( .B1(n6223), .B2(n6446), .A(n4549), .ZN(U3462) );
  AOI22_X1 U5626 ( .A1(n6379), .A2(n4611), .B1(n6339), .B2(n4610), .ZN(n4551)
         );
  INV_X1 U5627 ( .A(n6342), .ZN(n6380) );
  NAND2_X1 U5628 ( .A1(n4660), .A2(n6380), .ZN(n4550) );
  OAI211_X1 U5629 ( .C1(n6234), .C2(n6278), .A(n4551), .B(n4550), .ZN(n4552)
         );
  AOI21_X1 U5630 ( .B1(n4657), .B2(INSTQUEUE_REG_4__2__SCAN_IN), .A(n4552), 
        .ZN(n4553) );
  INV_X1 U5631 ( .A(n4553), .ZN(U3054) );
  NAND2_X1 U5632 ( .A1(n6133), .A2(DATAI_19_), .ZN(n6282) );
  NOR2_X2 U5633 ( .A1(n4609), .A2(n3309), .ZN(n6385) );
  INV_X1 U5634 ( .A(DATAI_3_), .ZN(n6073) );
  NOR2_X1 U5635 ( .A1(n6073), .A2(n4683), .ZN(n6279) );
  AOI22_X1 U5636 ( .A1(n6385), .A2(n4611), .B1(n6279), .B2(n4610), .ZN(n4556)
         );
  INV_X1 U5637 ( .A(DATAI_27_), .ZN(n4554) );
  NOR2_X1 U5638 ( .A1(n6145), .A2(n4554), .ZN(n6384) );
  NAND2_X1 U5639 ( .A1(n4660), .A2(n6384), .ZN(n4555) );
  OAI211_X1 U5640 ( .C1(n6234), .C2(n6282), .A(n4556), .B(n4555), .ZN(n4557)
         );
  AOI21_X1 U5641 ( .B1(n4657), .B2(INSTQUEUE_REG_4__3__SCAN_IN), .A(n4557), 
        .ZN(n4558) );
  INV_X1 U5642 ( .A(n4558), .ZN(U3055) );
  NAND2_X1 U5643 ( .A1(n6133), .A2(DATAI_20_), .ZN(n6285) );
  NOR2_X2 U5644 ( .A1(n4609), .A2(n4559), .ZN(n6391) );
  INV_X1 U5645 ( .A(DATAI_4_), .ZN(n6075) );
  NOR2_X1 U5646 ( .A1(n6075), .A2(n4683), .ZN(n6343) );
  AOI22_X1 U5647 ( .A1(n6391), .A2(n4611), .B1(n6343), .B2(n4610), .ZN(n4561)
         );
  NAND2_X1 U5648 ( .A1(n6133), .A2(DATAI_28_), .ZN(n6346) );
  INV_X1 U5649 ( .A(n6346), .ZN(n6390) );
  NAND2_X1 U5650 ( .A1(n4660), .A2(n6390), .ZN(n4560) );
  OAI211_X1 U5651 ( .C1(n6234), .C2(n6285), .A(n4561), .B(n4560), .ZN(n4562)
         );
  AOI21_X1 U5652 ( .B1(n4657), .B2(INSTQUEUE_REG_4__4__SCAN_IN), .A(n4562), 
        .ZN(n4563) );
  INV_X1 U5653 ( .A(n4563), .ZN(U3056) );
  INV_X1 U5654 ( .A(n6285), .ZN(n6392) );
  INV_X1 U5655 ( .A(n6391), .ZN(n5155) );
  INV_X1 U5656 ( .A(n6343), .ZN(n6395) );
  OAI22_X1 U5657 ( .A1(n5155), .A2(n4726), .B1(n4725), .B2(n6395), .ZN(n4564)
         );
  AOI21_X1 U5658 ( .B1(n6392), .B2(n4905), .A(n4564), .ZN(n4566) );
  NAND2_X1 U5659 ( .A1(n6417), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4565)
         );
  OAI211_X1 U5660 ( .C1(n6424), .C2(n6346), .A(n4566), .B(n4565), .ZN(U3144)
         );
  NOR2_X1 U5661 ( .A1(n4568), .A2(n4567), .ZN(n4569) );
  OR2_X1 U5662 ( .A1(n4570), .A2(n4569), .ZN(n6212) );
  INV_X1 U5663 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5980) );
  NOR2_X1 U5664 ( .A1(n4571), .A2(n4572), .ZN(n4573) );
  NOR2_X1 U5665 ( .A1(n4420), .A2(n4573), .ZN(n6132) );
  INV_X1 U5666 ( .A(n6132), .ZN(n4973) );
  OAI222_X1 U5667 ( .A1(n6212), .A2(n5773), .B1(n5980), .B2(n5997), .C1(n5480), 
        .C2(n4973), .ZN(U2857) );
  INV_X1 U5668 ( .A(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4579) );
  INV_X1 U5669 ( .A(DATAI_29_), .ZN(n4574) );
  NOR2_X1 U5670 ( .A1(n6145), .A2(n4574), .ZN(n6398) );
  INV_X1 U5671 ( .A(n6398), .ZN(n5167) );
  NOR2_X1 U5672 ( .A1(n4609), .A2(n4575), .ZN(n6397) );
  NAND2_X1 U5673 ( .A1(n6133), .A2(DATAI_21_), .ZN(n6289) );
  INV_X1 U5674 ( .A(n6289), .ZN(n6396) );
  AOI22_X1 U5675 ( .A1(n6397), .A2(n6348), .B1(n6347), .B2(n6396), .ZN(n4576)
         );
  OAI21_X1 U5676 ( .B1(n6354), .B2(n5167), .A(n4576), .ZN(n4577) );
  AOI21_X1 U5677 ( .B1(n6286), .B2(n6349), .A(n4577), .ZN(n4578) );
  OAI21_X1 U5678 ( .B1(n4580), .B2(n4579), .A(n4578), .ZN(U3113) );
  OAI21_X1 U5679 ( .B1(n4583), .B2(n4582), .A(n4581), .ZN(n6192) );
  AOI21_X1 U5680 ( .B1(n4420), .B2(n4586), .A(n4585), .ZN(n4587) );
  NOR2_X1 U5681 ( .A1(n4670), .A2(n4587), .ZN(n5970) );
  INV_X1 U5682 ( .A(n5969), .ZN(n4589) );
  NAND2_X1 U5683 ( .A1(n2971), .A2(REIP_REG_4__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U5684 ( .A1(n6142), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4588)
         );
  OAI211_X1 U5685 ( .C1(n6139), .C2(n4589), .A(n6189), .B(n4588), .ZN(n4590)
         );
  AOI21_X1 U5686 ( .B1(n5970), .B2(n6133), .A(n4590), .ZN(n4591) );
  OAI21_X1 U5687 ( .B1(n6137), .B2(n6192), .A(n4591), .ZN(U2982) );
  INV_X1 U5688 ( .A(n5970), .ZN(n4971) );
  INV_X1 U5689 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4595) );
  NAND2_X1 U5690 ( .A1(n4593), .A2(n4592), .ZN(n4594) );
  NAND2_X1 U5691 ( .A1(n4650), .A2(n4594), .ZN(n5960) );
  OAI222_X1 U5692 ( .A1(n4971), .A2(n5480), .B1(n5997), .B2(n4595), .C1(n5773), 
        .C2(n5960), .ZN(U2855) );
  NAND2_X1 U5693 ( .A1(n6133), .A2(DATAI_17_), .ZN(n6275) );
  NOR2_X2 U5694 ( .A1(n4609), .A2(n3054), .ZN(n6373) );
  INV_X1 U5695 ( .A(DATAI_1_), .ZN(n6069) );
  NOR2_X1 U5696 ( .A1(n6069), .A2(n4683), .ZN(n6335) );
  AOI22_X1 U5697 ( .A1(n6373), .A2(n4611), .B1(n6335), .B2(n4610), .ZN(n4598)
         );
  INV_X1 U5698 ( .A(DATAI_25_), .ZN(n4596) );
  NOR2_X1 U5699 ( .A1(n6145), .A2(n4596), .ZN(n6374) );
  NAND2_X1 U5700 ( .A1(n4660), .A2(n6374), .ZN(n4597) );
  OAI211_X1 U5701 ( .C1(n6234), .C2(n6275), .A(n4598), .B(n4597), .ZN(n4599)
         );
  AOI21_X1 U5702 ( .B1(n4657), .B2(INSTQUEUE_REG_4__1__SCAN_IN), .A(n4599), 
        .ZN(n4600) );
  INV_X1 U5703 ( .A(n4600), .ZN(U3053) );
  INV_X1 U5704 ( .A(n6384), .ZN(n5041) );
  NAND2_X1 U5705 ( .A1(n6349), .A2(n6279), .ZN(n4602) );
  INV_X1 U5706 ( .A(n6282), .ZN(n6386) );
  AOI22_X1 U5707 ( .A1(n6385), .A2(n6348), .B1(n6347), .B2(n6386), .ZN(n4601)
         );
  OAI211_X1 U5708 ( .C1(n5041), .C2(n6354), .A(n4602), .B(n4601), .ZN(n4603)
         );
  AOI21_X1 U5709 ( .B1(n6351), .B2(INSTQUEUE_REG_11__3__SCAN_IN), .A(n4603), 
        .ZN(n4604) );
  INV_X1 U5710 ( .A(n4604), .ZN(U3111) );
  INV_X1 U5711 ( .A(n6385), .ZN(n5147) );
  INV_X1 U5712 ( .A(n6279), .ZN(n6389) );
  OAI22_X1 U5713 ( .A1(n5147), .A2(n4726), .B1(n4725), .B2(n6389), .ZN(n4605)
         );
  AOI21_X1 U5714 ( .B1(n6386), .B2(n4905), .A(n4605), .ZN(n4607) );
  NAND2_X1 U5715 ( .A1(n6417), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4606)
         );
  OAI211_X1 U5716 ( .C1(n6424), .C2(n5041), .A(n4607), .B(n4606), .ZN(U3143)
         );
  NAND2_X1 U5717 ( .A1(n6133), .A2(DATAI_22_), .ZN(n6293) );
  NOR2_X2 U5718 ( .A1(n4609), .A2(n4608), .ZN(n6403) );
  INV_X1 U5719 ( .A(DATAI_6_), .ZN(n6078) );
  NOR2_X1 U5720 ( .A1(n6078), .A2(n4683), .ZN(n6290) );
  AOI22_X1 U5721 ( .A1(n6403), .A2(n4611), .B1(n6290), .B2(n4610), .ZN(n4613)
         );
  NAND2_X1 U5722 ( .A1(n4660), .A2(n6402), .ZN(n4612) );
  OAI211_X1 U5723 ( .C1(n6234), .C2(n6293), .A(n4613), .B(n4612), .ZN(n4614)
         );
  AOI21_X1 U5724 ( .B1(n4657), .B2(INSTQUEUE_REG_4__6__SCAN_IN), .A(n4614), 
        .ZN(n4615) );
  INV_X1 U5725 ( .A(n4615), .ZN(U3058) );
  INV_X1 U5726 ( .A(n6402), .ZN(n5036) );
  NAND2_X1 U5727 ( .A1(n6349), .A2(n6290), .ZN(n4617) );
  INV_X1 U5728 ( .A(n6293), .ZN(n6404) );
  AOI22_X1 U5729 ( .A1(n6403), .A2(n6348), .B1(n6347), .B2(n6404), .ZN(n4616)
         );
  OAI211_X1 U5730 ( .C1(n5036), .C2(n6354), .A(n4617), .B(n4616), .ZN(n4618)
         );
  AOI21_X1 U5731 ( .B1(n6351), .B2(INSTQUEUE_REG_11__6__SCAN_IN), .A(n4618), 
        .ZN(n4619) );
  INV_X1 U5732 ( .A(n4619), .ZN(U3114) );
  INV_X1 U5733 ( .A(n6412), .ZN(n6778) );
  INV_X1 U5734 ( .A(n4731), .ZN(n4620) );
  NAND2_X1 U5735 ( .A1(n5715), .A2(n4426), .ZN(n4867) );
  INV_X1 U5736 ( .A(n4867), .ZN(n4677) );
  NAND3_X1 U5737 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6442), .A3(n4863), .ZN(n4680) );
  NOR2_X1 U5738 ( .A1(n6356), .A2(n4680), .ZN(n4645) );
  AOI21_X1 U5739 ( .B1(n6358), .B2(n4677), .A(n4645), .ZN(n4626) );
  INV_X1 U5740 ( .A(n4626), .ZN(n4624) );
  OAI21_X1 U5741 ( .B1(n4622), .B2(n4621), .A(n6312), .ZN(n4625) );
  AOI21_X1 U5742 ( .B1(n6364), .B2(n4680), .A(n6362), .ZN(n4623) );
  OAI21_X1 U5743 ( .B1(n4624), .B2(n4625), .A(n4623), .ZN(n4644) );
  OAI22_X1 U5744 ( .A1(n4626), .A2(n4625), .B1(n6601), .B2(n4680), .ZN(n4643)
         );
  AOI22_X1 U5745 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4644), .B1(n6350), 
        .B2(n4643), .ZN(n4630) );
  INV_X1 U5746 ( .A(n6229), .ZN(n4627) );
  NAND2_X1 U5747 ( .A1(n4628), .A2(n4627), .ZN(n4772) );
  INV_X1 U5748 ( .A(n6301), .ZN(n6783) );
  AOI22_X1 U5749 ( .A1(n4812), .A2(n6783), .B1(n2999), .B2(n4645), .ZN(n4629)
         );
  OAI211_X1 U5750 ( .C1(n6778), .C2(n4708), .A(n4630), .B(n4629), .ZN(U3099)
         );
  AOI22_X1 U5751 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4644), .B1(n6343), 
        .B2(n4643), .ZN(n4632) );
  AOI22_X1 U5752 ( .A1(n4812), .A2(n6392), .B1(n6391), .B2(n4645), .ZN(n4631)
         );
  OAI211_X1 U5753 ( .C1(n6346), .C2(n4708), .A(n4632), .B(n4631), .ZN(U3096)
         );
  AOI22_X1 U5754 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4644), .B1(n6339), 
        .B2(n4643), .ZN(n4634) );
  AOI22_X1 U5755 ( .A1(n4812), .A2(n6378), .B1(n6379), .B2(n4645), .ZN(n4633)
         );
  OAI211_X1 U5756 ( .C1(n6342), .C2(n4708), .A(n4634), .B(n4633), .ZN(U3094)
         );
  AOI22_X1 U5757 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4644), .B1(n6286), 
        .B2(n4643), .ZN(n4636) );
  AOI22_X1 U5758 ( .A1(n4812), .A2(n6396), .B1(n6397), .B2(n4645), .ZN(n4635)
         );
  OAI211_X1 U5759 ( .C1(n5167), .C2(n4708), .A(n4636), .B(n4635), .ZN(U3097)
         );
  INV_X1 U5760 ( .A(n6374), .ZN(n6338) );
  AOI22_X1 U5761 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4644), .B1(n6335), 
        .B2(n4643), .ZN(n4638) );
  INV_X1 U5762 ( .A(n6275), .ZN(n6372) );
  AOI22_X1 U5763 ( .A1(n4812), .A2(n6372), .B1(n6373), .B2(n4645), .ZN(n4637)
         );
  OAI211_X1 U5764 ( .C1(n6338), .C2(n4708), .A(n4638), .B(n4637), .ZN(U3093)
         );
  AOI22_X1 U5765 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4644), .B1(n6290), 
        .B2(n4643), .ZN(n4640) );
  AOI22_X1 U5766 ( .A1(n4812), .A2(n6404), .B1(n6403), .B2(n4645), .ZN(n4639)
         );
  OAI211_X1 U5767 ( .C1(n5036), .C2(n4708), .A(n4640), .B(n4639), .ZN(U3098)
         );
  AOI22_X1 U5768 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4644), .B1(n6279), 
        .B2(n4643), .ZN(n4642) );
  AOI22_X1 U5769 ( .A1(n4812), .A2(n6386), .B1(n6385), .B2(n4645), .ZN(n4641)
         );
  OAI211_X1 U5770 ( .C1(n5041), .C2(n4708), .A(n4642), .B(n4641), .ZN(U3095)
         );
  AOI22_X1 U5771 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4644), .B1(n6421), 
        .B2(n4643), .ZN(n4647) );
  AOI22_X1 U5772 ( .A1(n4812), .A2(n6360), .B1(n6418), .B2(n4645), .ZN(n4646)
         );
  OAI211_X1 U5773 ( .C1(n6425), .C2(n4708), .A(n4647), .B(n4646), .ZN(U3092)
         );
  AND2_X1 U5774 ( .A1(n4650), .A2(n4649), .ZN(n4651) );
  NOR2_X1 U5775 ( .A1(n4648), .A2(n4651), .ZN(n5690) );
  INV_X1 U5776 ( .A(n5690), .ZN(n5957) );
  XNOR2_X1 U5777 ( .A(n4670), .B(n4652), .ZN(n6115) );
  INV_X1 U5778 ( .A(n6115), .ZN(n4985) );
  INV_X1 U5779 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4653) );
  OAI222_X1 U5780 ( .A1(n5957), .A2(n5773), .B1(n5480), .B2(n4985), .C1(n5997), 
        .C2(n4653), .ZN(U2854) );
  INV_X1 U5781 ( .A(n6397), .ZN(n5166) );
  OAI22_X1 U5782 ( .A1(n5166), .A2(n4726), .B1(n6289), .B2(n6423), .ZN(n4654)
         );
  AOI21_X1 U5783 ( .B1(n6398), .B2(n6782), .A(n4654), .ZN(n4656) );
  NAND2_X1 U5784 ( .A1(n6417), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4655)
         );
  OAI211_X1 U5785 ( .C1(n4725), .C2(n6401), .A(n4656), .B(n4655), .ZN(U3145)
         );
  NAND2_X1 U5786 ( .A1(n4657), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4662) );
  OAI22_X1 U5787 ( .A1(n5166), .A2(n4658), .B1(n6289), .B2(n6234), .ZN(n4659)
         );
  AOI21_X1 U5788 ( .B1(n6398), .B2(n4660), .A(n4659), .ZN(n4661) );
  OAI211_X1 U5789 ( .C1(n4663), .C2(n6401), .A(n4662), .B(n4661), .ZN(U3057)
         );
  NOR2_X1 U5790 ( .A1(n4648), .A2(n4664), .ZN(n4665) );
  OR2_X1 U5791 ( .A1(n5930), .A2(n4665), .ZN(n6177) );
  INV_X1 U5792 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4672) );
  INV_X1 U5793 ( .A(n4652), .ZN(n4669) );
  INV_X1 U5794 ( .A(n4667), .ZN(n4668) );
  AOI21_X1 U5795 ( .B1(n4670), .B2(n4669), .A(n4668), .ZN(n4671) );
  OR2_X1 U5796 ( .A1(n4666), .A2(n4671), .ZN(n5947) );
  OAI222_X1 U5797 ( .A1(n6177), .A2(n5773), .B1(n4672), .B2(n5997), .C1(n5947), 
        .C2(n5480), .ZN(U2853) );
  INV_X1 U5798 ( .A(n6373), .ZN(n5151) );
  INV_X1 U5799 ( .A(n6335), .ZN(n6377) );
  OAI22_X1 U5800 ( .A1(n5151), .A2(n4726), .B1(n4725), .B2(n6377), .ZN(n4673)
         );
  AOI21_X1 U5801 ( .B1(n6372), .B2(n4905), .A(n4673), .ZN(n4675) );
  NAND2_X1 U5802 ( .A1(n6417), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4674)
         );
  OAI211_X1 U5803 ( .C1(n6424), .C2(n6338), .A(n4675), .B(n4674), .ZN(U3141)
         );
  NAND3_X1 U5804 ( .A1(n4708), .A2(n6312), .A3(n4719), .ZN(n4679) );
  NAND2_X1 U5805 ( .A1(n4677), .A2(n4924), .ZN(n4687) );
  INV_X1 U5806 ( .A(n4687), .ZN(n4678) );
  AOI21_X1 U5807 ( .B1(n4679), .B2(n5138), .A(n4678), .ZN(n4686) );
  NOR2_X1 U5808 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4680), .ZN(n4716)
         );
  INV_X1 U5809 ( .A(n6262), .ZN(n4684) );
  INV_X1 U5810 ( .A(n4681), .ZN(n4682) );
  OR2_X1 U5811 ( .A1(n4682), .A2(n5144), .ZN(n4739) );
  AOI21_X1 U5812 ( .B1(n4739), .B2(STATE2_REG_2__SCAN_IN), .A(n4683), .ZN(
        n4735) );
  OAI211_X1 U5813 ( .C1(n6718), .C2(n4716), .A(n4684), .B(n4735), .ZN(n4685)
         );
  INV_X1 U5814 ( .A(n6267), .ZN(n4780) );
  OAI22_X1 U5815 ( .A1(n4687), .A2(n6364), .B1(n4780), .B2(n4739), .ZN(n4721)
         );
  INV_X1 U5816 ( .A(n4708), .ZN(n4717) );
  AOI22_X1 U5817 ( .A1(n6783), .A2(n4717), .B1(n6410), .B2(n4716), .ZN(n4688)
         );
  OAI21_X1 U5818 ( .B1(n6778), .B2(n4719), .A(n4688), .ZN(n4689) );
  AOI21_X1 U5819 ( .B1(n6350), .B2(n4721), .A(n4689), .ZN(n4690) );
  OAI21_X1 U5820 ( .B1(n4724), .B2(n6693), .A(n4690), .ZN(U3091) );
  INV_X1 U5821 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4694) );
  AOI22_X1 U5822 ( .A1(n6403), .A2(n4716), .B1(n6290), .B2(n4721), .ZN(n4691)
         );
  OAI21_X1 U5823 ( .B1(n6293), .B2(n4708), .A(n4691), .ZN(n4692) );
  AOI21_X1 U5824 ( .B1(n6402), .B2(n6328), .A(n4692), .ZN(n4693) );
  OAI21_X1 U5825 ( .B1(n4724), .B2(n4694), .A(n4693), .ZN(U3090) );
  INV_X1 U5826 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4698) );
  AOI22_X1 U5827 ( .A1(n6385), .A2(n4716), .B1(n6279), .B2(n4721), .ZN(n4695)
         );
  OAI21_X1 U5828 ( .B1(n6282), .B2(n4708), .A(n4695), .ZN(n4696) );
  AOI21_X1 U5829 ( .B1(n6384), .B2(n6328), .A(n4696), .ZN(n4697) );
  OAI21_X1 U5830 ( .B1(n4724), .B2(n4698), .A(n4697), .ZN(U3087) );
  INV_X1 U5831 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4702) );
  AOI22_X1 U5832 ( .A1(n6391), .A2(n4716), .B1(n6343), .B2(n4721), .ZN(n4699)
         );
  OAI21_X1 U5833 ( .B1(n6285), .B2(n4708), .A(n4699), .ZN(n4700) );
  AOI21_X1 U5834 ( .B1(n6390), .B2(n6328), .A(n4700), .ZN(n4701) );
  OAI21_X1 U5835 ( .B1(n4724), .B2(n4702), .A(n4701), .ZN(U3088) );
  INV_X1 U5836 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4706) );
  AOI22_X1 U5837 ( .A1(n6379), .A2(n4716), .B1(n6339), .B2(n4721), .ZN(n4703)
         );
  OAI21_X1 U5838 ( .B1(n6278), .B2(n4708), .A(n4703), .ZN(n4704) );
  AOI21_X1 U5839 ( .B1(n6380), .B2(n6328), .A(n4704), .ZN(n4705) );
  OAI21_X1 U5840 ( .B1(n4724), .B2(n4706), .A(n4705), .ZN(U3086) );
  INV_X1 U5841 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4711) );
  AOI22_X1 U5842 ( .A1(n6373), .A2(n4716), .B1(n6335), .B2(n4721), .ZN(n4707)
         );
  OAI21_X1 U5843 ( .B1(n6275), .B2(n4708), .A(n4707), .ZN(n4709) );
  AOI21_X1 U5844 ( .B1(n6374), .B2(n6328), .A(n4709), .ZN(n4710) );
  OAI21_X1 U5845 ( .B1(n4724), .B2(n4711), .A(n4710), .ZN(U3085) );
  INV_X1 U5846 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4715) );
  AOI22_X1 U5847 ( .A1(n6396), .A2(n4717), .B1(n6397), .B2(n4716), .ZN(n4712)
         );
  OAI21_X1 U5848 ( .B1(n5167), .B2(n4719), .A(n4712), .ZN(n4713) );
  AOI21_X1 U5849 ( .B1(n6286), .B2(n4721), .A(n4713), .ZN(n4714) );
  OAI21_X1 U5850 ( .B1(n4724), .B2(n4715), .A(n4714), .ZN(U3089) );
  INV_X1 U5851 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4723) );
  AOI22_X1 U5852 ( .A1(n6360), .A2(n4717), .B1(n6418), .B2(n4716), .ZN(n4718)
         );
  OAI21_X1 U5853 ( .B1(n6425), .B2(n4719), .A(n4718), .ZN(n4720) );
  AOI21_X1 U5854 ( .B1(n6421), .B2(n4721), .A(n4720), .ZN(n4722) );
  OAI21_X1 U5855 ( .B1(n4724), .B2(n4723), .A(n4722), .ZN(U3084) );
  INV_X1 U5856 ( .A(n6403), .ZN(n5171) );
  INV_X1 U5857 ( .A(n6290), .ZN(n6407) );
  OAI22_X1 U5858 ( .A1(n5171), .A2(n4726), .B1(n4725), .B2(n6407), .ZN(n4727)
         );
  AOI21_X1 U5859 ( .B1(n6404), .B2(n4905), .A(n4727), .ZN(n4729) );
  NAND2_X1 U5860 ( .A1(n6417), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4728)
         );
  OAI211_X1 U5861 ( .C1(n6424), .C2(n5036), .A(n4729), .B(n4728), .ZN(U3146)
         );
  INV_X1 U5862 ( .A(n6347), .ZN(n4770) );
  NAND2_X1 U5863 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4730), .ZN(n6363) );
  NOR2_X1 U5864 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6363), .ZN(n4738)
         );
  NOR3_X1 U5865 ( .A1(n6347), .A2(n6411), .A3(n6364), .ZN(n4734) );
  OAI22_X1 U5866 ( .A1(n4734), .A2(n4868), .B1(n4733), .B2(n4732), .ZN(n4737)
         );
  AND2_X1 U5867 ( .A1(n4780), .A2(n4735), .ZN(n4736) );
  NAND2_X1 U5868 ( .A1(n4764), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4744)
         );
  INV_X1 U5869 ( .A(n4738), .ZN(n4766) );
  INV_X1 U5870 ( .A(n4739), .ZN(n4740) );
  AOI22_X1 U5871 ( .A1(n4741), .A2(n4924), .B1(n4740), .B2(n6262), .ZN(n4765)
         );
  OAI22_X1 U5872 ( .A1(n5162), .A2(n4766), .B1(n4765), .B2(n6383), .ZN(n4742)
         );
  AOI21_X1 U5873 ( .B1(n6378), .B2(n6411), .A(n4742), .ZN(n4743) );
  OAI211_X1 U5874 ( .C1(n4770), .C2(n6342), .A(n4744), .B(n4743), .ZN(U3118)
         );
  NAND2_X1 U5875 ( .A1(n4764), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4747)
         );
  OAI22_X1 U5876 ( .A1(n6780), .A2(n4766), .B1(n6301), .B2(n4754), .ZN(n4745)
         );
  AOI21_X1 U5877 ( .B1(n6412), .B2(n6347), .A(n4745), .ZN(n4746) );
  OAI211_X1 U5878 ( .C1(n4765), .C2(n6786), .A(n4747), .B(n4746), .ZN(U3123)
         );
  NAND2_X1 U5879 ( .A1(n4764), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4750)
         );
  OAI22_X1 U5880 ( .A1(n5151), .A2(n4766), .B1(n4765), .B2(n6377), .ZN(n4748)
         );
  AOI21_X1 U5881 ( .B1(n6372), .B2(n6411), .A(n4748), .ZN(n4749) );
  OAI211_X1 U5882 ( .C1(n4770), .C2(n6338), .A(n4750), .B(n4749), .ZN(U3117)
         );
  NAND2_X1 U5883 ( .A1(n4764), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4753)
         );
  OAI22_X1 U5884 ( .A1(n5179), .A2(n4766), .B1(n6422), .B2(n4754), .ZN(n4751)
         );
  AOI21_X1 U5885 ( .B1(n6368), .B2(n6347), .A(n4751), .ZN(n4752) );
  OAI211_X1 U5886 ( .C1(n4765), .C2(n6371), .A(n4753), .B(n4752), .ZN(U3116)
         );
  NAND2_X1 U5887 ( .A1(n4764), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4757)
         );
  OAI22_X1 U5888 ( .A1(n5166), .A2(n4766), .B1(n6289), .B2(n4754), .ZN(n4755)
         );
  AOI21_X1 U5889 ( .B1(n6398), .B2(n6347), .A(n4755), .ZN(n4756) );
  OAI211_X1 U5890 ( .C1(n4765), .C2(n6401), .A(n4757), .B(n4756), .ZN(U3121)
         );
  NAND2_X1 U5891 ( .A1(n4764), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4760)
         );
  OAI22_X1 U5892 ( .A1(n5171), .A2(n4766), .B1(n4765), .B2(n6407), .ZN(n4758)
         );
  AOI21_X1 U5893 ( .B1(n6404), .B2(n6411), .A(n4758), .ZN(n4759) );
  OAI211_X1 U5894 ( .C1(n4770), .C2(n5036), .A(n4760), .B(n4759), .ZN(U3122)
         );
  NAND2_X1 U5895 ( .A1(n4764), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4763)
         );
  OAI22_X1 U5896 ( .A1(n5147), .A2(n4766), .B1(n4765), .B2(n6389), .ZN(n4761)
         );
  AOI21_X1 U5897 ( .B1(n6386), .B2(n6411), .A(n4761), .ZN(n4762) );
  OAI211_X1 U5898 ( .C1(n4770), .C2(n5041), .A(n4763), .B(n4762), .ZN(U3119)
         );
  NAND2_X1 U5899 ( .A1(n4764), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4769)
         );
  OAI22_X1 U5900 ( .A1(n5155), .A2(n4766), .B1(n4765), .B2(n6395), .ZN(n4767)
         );
  AOI21_X1 U5901 ( .B1(n6392), .B2(n6411), .A(n4767), .ZN(n4768) );
  OAI211_X1 U5902 ( .C1(n4770), .C2(n6346), .A(n4769), .B(n4768), .ZN(U3120)
         );
  OAI21_X1 U5903 ( .B1(n5144), .B2(n6601), .A(n4771), .ZN(n6266) );
  NOR2_X1 U5904 ( .A1(n6262), .A2(n6266), .ZN(n5141) );
  NAND2_X1 U5905 ( .A1(n6354), .A2(n4772), .ZN(n4773) );
  NAND2_X1 U5906 ( .A1(n4773), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4774) );
  NAND2_X1 U5907 ( .A1(n4774), .A2(n6312), .ZN(n4782) );
  INV_X1 U5908 ( .A(n4781), .ZN(n4776) );
  NOR2_X1 U5909 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4775), .ZN(n4811)
         );
  OAI22_X1 U5910 ( .A1(n4782), .A2(n4776), .B1(n4811), .B2(n6718), .ZN(n4777)
         );
  INV_X1 U5911 ( .A(n4777), .ZN(n4778) );
  OAI211_X1 U5912 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6601), .A(n5141), .B(n4778), .ZN(n4779) );
  INV_X1 U5913 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4786) );
  NAND2_X1 U5914 ( .A1(n5144), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4819) );
  OAI22_X1 U5915 ( .A1(n4782), .A2(n4781), .B1(n4780), .B2(n4819), .ZN(n4815)
         );
  AOI22_X1 U5916 ( .A1(n4812), .A2(n6368), .B1(n6418), .B2(n4811), .ZN(n4783)
         );
  OAI21_X1 U5917 ( .B1(n6354), .B2(n6422), .A(n4783), .ZN(n4784) );
  AOI21_X1 U5918 ( .B1(n4815), .B2(n6421), .A(n4784), .ZN(n4785) );
  OAI21_X1 U5919 ( .B1(n4818), .B2(n4786), .A(n4785), .ZN(U3100) );
  INV_X1 U5920 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4790) );
  AOI22_X1 U5921 ( .A1(n4812), .A2(n6380), .B1(n6379), .B2(n4811), .ZN(n4787)
         );
  OAI21_X1 U5922 ( .B1(n6354), .B2(n6278), .A(n4787), .ZN(n4788) );
  AOI21_X1 U5923 ( .B1(n4815), .B2(n6339), .A(n4788), .ZN(n4789) );
  OAI21_X1 U5924 ( .B1(n4818), .B2(n4790), .A(n4789), .ZN(U3102) );
  INV_X1 U5925 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4794) );
  AOI22_X1 U5926 ( .A1(n6373), .A2(n4811), .B1(n4812), .B2(n6374), .ZN(n4791)
         );
  OAI21_X1 U5927 ( .B1(n6354), .B2(n6275), .A(n4791), .ZN(n4792) );
  AOI21_X1 U5928 ( .B1(n4815), .B2(n6335), .A(n4792), .ZN(n4793) );
  OAI21_X1 U5929 ( .B1(n4818), .B2(n4794), .A(n4793), .ZN(U3101) );
  INV_X1 U5930 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4798) );
  AOI22_X1 U5931 ( .A1(n4812), .A2(n6390), .B1(n6391), .B2(n4811), .ZN(n4795)
         );
  OAI21_X1 U5932 ( .B1(n6354), .B2(n6285), .A(n4795), .ZN(n4796) );
  AOI21_X1 U5933 ( .B1(n4815), .B2(n6343), .A(n4796), .ZN(n4797) );
  OAI21_X1 U5934 ( .B1(n4818), .B2(n4798), .A(n4797), .ZN(U3104) );
  INV_X1 U5935 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4802) );
  AOI22_X1 U5936 ( .A1(n4812), .A2(n6412), .B1(n6410), .B2(n4811), .ZN(n4799)
         );
  OAI21_X1 U5937 ( .B1(n6354), .B2(n6301), .A(n4799), .ZN(n4800) );
  AOI21_X1 U5938 ( .B1(n4815), .B2(n6350), .A(n4800), .ZN(n4801) );
  OAI21_X1 U5939 ( .B1(n4818), .B2(n4802), .A(n4801), .ZN(U3107) );
  INV_X1 U5940 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4806) );
  AOI22_X1 U5941 ( .A1(n4812), .A2(n6402), .B1(n6403), .B2(n4811), .ZN(n4803)
         );
  OAI21_X1 U5942 ( .B1(n6354), .B2(n6293), .A(n4803), .ZN(n4804) );
  AOI21_X1 U5943 ( .B1(n4815), .B2(n6290), .A(n4804), .ZN(n4805) );
  OAI21_X1 U5944 ( .B1(n4818), .B2(n4806), .A(n4805), .ZN(U3106) );
  INV_X1 U5945 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4810) );
  AOI22_X1 U5946 ( .A1(n4812), .A2(n6398), .B1(n6397), .B2(n4811), .ZN(n4807)
         );
  OAI21_X1 U5947 ( .B1(n6354), .B2(n6289), .A(n4807), .ZN(n4808) );
  AOI21_X1 U5948 ( .B1(n4815), .B2(n6286), .A(n4808), .ZN(n4809) );
  OAI21_X1 U5949 ( .B1(n4818), .B2(n4810), .A(n4809), .ZN(U3105) );
  INV_X1 U5950 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4817) );
  AOI22_X1 U5951 ( .A1(n4812), .A2(n6384), .B1(n6385), .B2(n4811), .ZN(n4813)
         );
  OAI21_X1 U5952 ( .B1(n6354), .B2(n6282), .A(n4813), .ZN(n4814) );
  AOI21_X1 U5953 ( .B1(n4815), .B2(n6279), .A(n4814), .ZN(n4816) );
  OAI21_X1 U5954 ( .B1(n4818), .B2(n4817), .A(n4816), .ZN(U3103) );
  NOR2_X1 U5955 ( .A1(n4824), .A2(n6364), .ZN(n6264) );
  INV_X1 U5956 ( .A(n4819), .ZN(n4820) );
  AOI22_X1 U5957 ( .A1(n6264), .A2(n4924), .B1(n6262), .B2(n4820), .ZN(n6787)
         );
  NOR2_X1 U5958 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4821), .ZN(n4827)
         );
  NOR3_X1 U5959 ( .A1(n6266), .A2(n6446), .A3(n6267), .ZN(n4826) );
  OAI21_X1 U5960 ( .B1(n6782), .B2(n6408), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4823) );
  NAND3_X1 U5961 ( .A1(n4824), .A2(n6312), .A3(n4823), .ZN(n4825) );
  OAI211_X1 U5962 ( .C1(n4827), .C2(n6718), .A(n4826), .B(n4825), .ZN(n6776)
         );
  NAND2_X1 U5963 ( .A1(n6776), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4830)
         );
  INV_X1 U5964 ( .A(n4827), .ZN(n6779) );
  OAI22_X1 U5965 ( .A1(n5166), .A2(n6779), .B1(n5167), .B2(n6777), .ZN(n4828)
         );
  AOI21_X1 U5966 ( .B1(n6396), .B2(n6782), .A(n4828), .ZN(n4829) );
  OAI211_X1 U5967 ( .C1(n6787), .C2(n6401), .A(n4830), .B(n4829), .ZN(U3137)
         );
  NAND2_X1 U5968 ( .A1(n6776), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4833)
         );
  OAI22_X1 U5969 ( .A1(n5179), .A2(n6779), .B1(n6425), .B2(n6777), .ZN(n4831)
         );
  AOI21_X1 U5970 ( .B1(n6360), .B2(n6782), .A(n4831), .ZN(n4832) );
  OAI211_X1 U5971 ( .C1(n6787), .C2(n6371), .A(n4833), .B(n4832), .ZN(U3132)
         );
  NAND2_X1 U5972 ( .A1(n6776), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4836)
         );
  OAI22_X1 U5973 ( .A1(n5151), .A2(n6779), .B1(n6787), .B2(n6377), .ZN(n4834)
         );
  AOI21_X1 U5974 ( .B1(n6374), .B2(n6408), .A(n4834), .ZN(n4835) );
  OAI211_X1 U5975 ( .C1(n6424), .C2(n6275), .A(n4836), .B(n4835), .ZN(U3133)
         );
  NAND2_X1 U5976 ( .A1(n6776), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4839)
         );
  OAI22_X1 U5977 ( .A1(n5171), .A2(n6779), .B1(n6787), .B2(n6407), .ZN(n4837)
         );
  AOI21_X1 U5978 ( .B1(n6402), .B2(n6408), .A(n4837), .ZN(n4838) );
  OAI211_X1 U5979 ( .C1(n6424), .C2(n6293), .A(n4839), .B(n4838), .ZN(U3138)
         );
  NAND2_X1 U5980 ( .A1(n6776), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4842)
         );
  OAI22_X1 U5981 ( .A1(n5155), .A2(n6779), .B1(n6787), .B2(n6395), .ZN(n4840)
         );
  AOI21_X1 U5982 ( .B1(n6390), .B2(n6408), .A(n4840), .ZN(n4841) );
  OAI211_X1 U5983 ( .C1(n6424), .C2(n6285), .A(n4842), .B(n4841), .ZN(U3136)
         );
  NAND2_X1 U5984 ( .A1(n6776), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4845)
         );
  OAI22_X1 U5985 ( .A1(n5147), .A2(n6779), .B1(n6787), .B2(n6389), .ZN(n4843)
         );
  AOI21_X1 U5986 ( .B1(n6384), .B2(n6408), .A(n4843), .ZN(n4844) );
  OAI211_X1 U5987 ( .C1(n6424), .C2(n6282), .A(n4845), .B(n4844), .ZN(U3135)
         );
  NAND2_X1 U5988 ( .A1(n6776), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4848)
         );
  OAI22_X1 U5989 ( .A1(n5162), .A2(n6779), .B1(n6787), .B2(n6383), .ZN(n4846)
         );
  AOI21_X1 U5990 ( .B1(n6380), .B2(n6408), .A(n4846), .ZN(n4847) );
  OAI211_X1 U5991 ( .C1(n6424), .C2(n6278), .A(n4848), .B(n4847), .ZN(U3134)
         );
  INV_X1 U5992 ( .A(n4849), .ZN(n5929) );
  NAND2_X1 U5993 ( .A1(n5930), .A2(n5929), .ZN(n4851) );
  NAND2_X1 U5994 ( .A1(n4851), .A2(n4850), .ZN(n4852) );
  NAND2_X1 U5995 ( .A1(n4852), .A2(n4348), .ZN(n6159) );
  INV_X1 U5996 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U5997 ( .A1(n4855), .A2(n4854), .ZN(n4856) );
  AND2_X1 U5998 ( .A1(n4853), .A2(n4856), .ZN(n4994) );
  INV_X1 U5999 ( .A(n4994), .ZN(n4984) );
  OAI222_X1 U6000 ( .A1(n6159), .A2(n5773), .B1(n4976), .B2(n5997), .C1(n5480), 
        .C2(n4984), .ZN(U2851) );
  OAI21_X1 U6001 ( .B1(n4859), .B2(n4858), .A(n4857), .ZN(n6181) );
  NAND2_X1 U6002 ( .A1(n2971), .A2(REIP_REG_6__SCAN_IN), .ZN(n6178) );
  OAI21_X1 U6003 ( .B1(n5824), .B2(n3806), .A(n6178), .ZN(n4861) );
  NOR2_X1 U6004 ( .A1(n5947), .A2(n6145), .ZN(n4860) );
  AOI211_X1 U6005 ( .C1(n5821), .C2(n5949), .A(n4861), .B(n4860), .ZN(n4862)
         );
  OAI21_X1 U6006 ( .B1(n6137), .B2(n6181), .A(n4862), .ZN(U2980) );
  NAND3_X1 U6007 ( .A1(n6446), .A2(n6442), .A3(n4863), .ZN(n5025) );
  NOR2_X1 U6008 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5025), .ZN(n4904)
         );
  INV_X1 U6009 ( .A(n4904), .ZN(n4865) );
  AOI211_X1 U6010 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4865), .A(n6262), .B(
        n4864), .ZN(n4871) );
  INV_X1 U6011 ( .A(n5029), .ZN(n4866) );
  INV_X1 U6012 ( .A(n5051), .ZN(n4882) );
  NOR3_X1 U6013 ( .A1(n4882), .A2(n4905), .A3(n6364), .ZN(n4869) );
  OR2_X1 U6014 ( .A1(n4924), .A2(n4867), .ZN(n5021) );
  OAI21_X1 U6015 ( .B1(n4869), .B2(n4868), .A(n5021), .ZN(n4870) );
  NAND2_X1 U6016 ( .A1(n4871), .A2(n4870), .ZN(n4909) );
  AOI22_X1 U6017 ( .A1(n4882), .A2(n6783), .B1(n2999), .B2(n4904), .ZN(n4875)
         );
  NAND2_X1 U6018 ( .A1(n6267), .A2(n4872), .ZN(n4873) );
  OAI21_X1 U6019 ( .B1(n5021), .B2(n6364), .A(n4873), .ZN(n4903) );
  NAND2_X1 U6020 ( .A1(n6350), .A2(n4903), .ZN(n4874) );
  OAI211_X1 U6021 ( .C1(n6423), .C2(n6778), .A(n4875), .B(n4874), .ZN(n4876)
         );
  AOI21_X1 U6022 ( .B1(n4909), .B2(INSTQUEUE_REG_0__7__SCAN_IN), .A(n4876), 
        .ZN(n4877) );
  INV_X1 U6023 ( .A(n4877), .ZN(U3027) );
  AOI22_X1 U6024 ( .A1(n4882), .A2(n6396), .B1(n6397), .B2(n4904), .ZN(n4879)
         );
  NAND2_X1 U6025 ( .A1(n6286), .A2(n4903), .ZN(n4878) );
  OAI211_X1 U6026 ( .C1(n6423), .C2(n5167), .A(n4879), .B(n4878), .ZN(n4880)
         );
  AOI21_X1 U6027 ( .B1(n4909), .B2(INSTQUEUE_REG_0__5__SCAN_IN), .A(n4880), 
        .ZN(n4881) );
  INV_X1 U6028 ( .A(n4881), .ZN(U3025) );
  AOI22_X1 U6029 ( .A1(n4882), .A2(n6360), .B1(n6418), .B2(n4904), .ZN(n4884)
         );
  NAND2_X1 U6030 ( .A1(n6421), .A2(n4903), .ZN(n4883) );
  OAI211_X1 U6031 ( .C1(n6423), .C2(n6425), .A(n4884), .B(n4883), .ZN(n4885)
         );
  AOI21_X1 U6032 ( .B1(n4909), .B2(INSTQUEUE_REG_0__0__SCAN_IN), .A(n4885), 
        .ZN(n4886) );
  INV_X1 U6033 ( .A(n4886), .ZN(U3020) );
  AOI22_X1 U6034 ( .A1(n6379), .A2(n4904), .B1(n6339), .B2(n4903), .ZN(n4888)
         );
  NAND2_X1 U6035 ( .A1(n4905), .A2(n6380), .ZN(n4887) );
  OAI211_X1 U6036 ( .C1(n5051), .C2(n6278), .A(n4888), .B(n4887), .ZN(n4889)
         );
  AOI21_X1 U6037 ( .B1(n4909), .B2(INSTQUEUE_REG_0__2__SCAN_IN), .A(n4889), 
        .ZN(n4890) );
  INV_X1 U6038 ( .A(n4890), .ZN(U3022) );
  AOI22_X1 U6039 ( .A1(n6385), .A2(n4904), .B1(n6279), .B2(n4903), .ZN(n4892)
         );
  NAND2_X1 U6040 ( .A1(n4905), .A2(n6384), .ZN(n4891) );
  OAI211_X1 U6041 ( .C1(n5051), .C2(n6282), .A(n4892), .B(n4891), .ZN(n4893)
         );
  AOI21_X1 U6042 ( .B1(n4909), .B2(INSTQUEUE_REG_0__3__SCAN_IN), .A(n4893), 
        .ZN(n4894) );
  INV_X1 U6043 ( .A(n4894), .ZN(U3023) );
  AOI22_X1 U6044 ( .A1(n6373), .A2(n4904), .B1(n6335), .B2(n4903), .ZN(n4896)
         );
  NAND2_X1 U6045 ( .A1(n4905), .A2(n6374), .ZN(n4895) );
  OAI211_X1 U6046 ( .C1(n5051), .C2(n6275), .A(n4896), .B(n4895), .ZN(n4897)
         );
  AOI21_X1 U6047 ( .B1(n4909), .B2(INSTQUEUE_REG_0__1__SCAN_IN), .A(n4897), 
        .ZN(n4898) );
  INV_X1 U6048 ( .A(n4898), .ZN(U3021) );
  AOI22_X1 U6049 ( .A1(n6403), .A2(n4904), .B1(n6290), .B2(n4903), .ZN(n4900)
         );
  NAND2_X1 U6050 ( .A1(n4905), .A2(n6402), .ZN(n4899) );
  OAI211_X1 U6051 ( .C1(n5051), .C2(n6293), .A(n4900), .B(n4899), .ZN(n4901)
         );
  AOI21_X1 U6052 ( .B1(n4909), .B2(INSTQUEUE_REG_0__6__SCAN_IN), .A(n4901), 
        .ZN(n4902) );
  INV_X1 U6053 ( .A(n4902), .ZN(U3026) );
  AOI22_X1 U6054 ( .A1(n6391), .A2(n4904), .B1(n6343), .B2(n4903), .ZN(n4907)
         );
  NAND2_X1 U6055 ( .A1(n4905), .A2(n6390), .ZN(n4906) );
  OAI211_X1 U6056 ( .C1(n5051), .C2(n6285), .A(n4907), .B(n4906), .ZN(n4908)
         );
  AOI21_X1 U6057 ( .B1(n4909), .B2(INSTQUEUE_REG_0__4__SCAN_IN), .A(n4908), 
        .ZN(n4910) );
  INV_X1 U6058 ( .A(n4910), .ZN(U3024) );
  AOI21_X1 U6059 ( .B1(n4911), .B2(n4853), .A(n4336), .ZN(n5104) );
  INV_X1 U6060 ( .A(n5104), .ZN(n5067) );
  XNOR2_X1 U6061 ( .A(n4348), .B(n4912), .ZN(n5098) );
  INV_X1 U6062 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5096) );
  OAI222_X1 U6063 ( .A1(n5067), .A2(n5480), .B1(n5773), .B2(n5098), .C1(n5997), 
        .C2(n5096), .ZN(U2850) );
  INV_X1 U6064 ( .A(n6005), .ZN(n4914) );
  INV_X1 U6065 ( .A(n6009), .ZN(n4913) );
  AOI22_X1 U6066 ( .A1(n5244), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n6008), .ZN(n4915) );
  OAI21_X1 U6067 ( .B1(n4984), .B2(n5499), .A(n4915), .ZN(U2883) );
  XOR2_X1 U6068 ( .A(n4916), .B(n4666), .Z(n6110) );
  INV_X1 U6069 ( .A(n6110), .ZN(n4918) );
  AOI22_X1 U6070 ( .A1(n5244), .A2(DATAI_7_), .B1(EAX_REG_7__SCAN_IN), .B2(
        n6008), .ZN(n4917) );
  OAI21_X1 U6071 ( .B1(n4918), .B2(n5499), .A(n4917), .ZN(U2884) );
  OR2_X1 U6072 ( .A1(n4919), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5137)
         );
  INV_X1 U6073 ( .A(n5710), .ZN(n4920) );
  AOI21_X1 U6074 ( .B1(n4920), .B2(n4429), .A(n6364), .ZN(n4921) );
  NOR2_X1 U6075 ( .A1(n4922), .A2(n4921), .ZN(n4930) );
  INV_X1 U6076 ( .A(n4923), .ZN(n4925) );
  NOR2_X1 U6077 ( .A1(n4925), .A2(n4924), .ZN(n5146) );
  INV_X1 U6078 ( .A(n5146), .ZN(n5139) );
  NOR2_X1 U6079 ( .A1(n6356), .A2(n5137), .ZN(n4962) );
  INV_X1 U6080 ( .A(n4962), .ZN(n4926) );
  OAI21_X1 U6081 ( .B1(n5139), .B2(n6224), .A(n4926), .ZN(n4928) );
  NOR2_X1 U6082 ( .A1(n4930), .A2(n4928), .ZN(n4927) );
  INV_X1 U6083 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4937) );
  INV_X1 U6084 ( .A(n4928), .ZN(n4929) );
  OAI22_X1 U6085 ( .A1(n4930), .A2(n4929), .B1(n6601), .B2(n5137), .ZN(n4966)
         );
  INV_X1 U6086 ( .A(n4931), .ZN(n4933) );
  NAND2_X1 U6087 ( .A1(n4933), .A2(n4932), .ZN(n5176) );
  AOI22_X1 U6088 ( .A1(n2999), .A2(n4962), .B1(n5182), .B2(n6412), .ZN(n4934)
         );
  OAI21_X1 U6089 ( .B1(n6301), .B2(n4964), .A(n4934), .ZN(n4935) );
  AOI21_X1 U6090 ( .B1(n4966), .B2(n6350), .A(n4935), .ZN(n4936) );
  OAI21_X1 U6091 ( .B1(n4969), .B2(n4937), .A(n4936), .ZN(U3051) );
  INV_X1 U6092 ( .A(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4941) );
  AOI22_X1 U6093 ( .A1(n6403), .A2(n4962), .B1(n5182), .B2(n6402), .ZN(n4938)
         );
  OAI21_X1 U6094 ( .B1(n6293), .B2(n4964), .A(n4938), .ZN(n4939) );
  AOI21_X1 U6095 ( .B1(n4966), .B2(n6290), .A(n4939), .ZN(n4940) );
  OAI21_X1 U6096 ( .B1(n4969), .B2(n4941), .A(n4940), .ZN(U3050) );
  INV_X1 U6097 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4945) );
  AOI22_X1 U6098 ( .A1(n6397), .A2(n4962), .B1(n5182), .B2(n6398), .ZN(n4942)
         );
  OAI21_X1 U6099 ( .B1(n6289), .B2(n4964), .A(n4942), .ZN(n4943) );
  AOI21_X1 U6100 ( .B1(n4966), .B2(n6286), .A(n4943), .ZN(n4944) );
  OAI21_X1 U6101 ( .B1(n4969), .B2(n4945), .A(n4944), .ZN(U3049) );
  INV_X1 U6102 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4949) );
  AOI22_X1 U6103 ( .A1(n6391), .A2(n4962), .B1(n5182), .B2(n6390), .ZN(n4946)
         );
  OAI21_X1 U6104 ( .B1(n6285), .B2(n4964), .A(n4946), .ZN(n4947) );
  AOI21_X1 U6105 ( .B1(n4966), .B2(n6343), .A(n4947), .ZN(n4948) );
  OAI21_X1 U6106 ( .B1(n4969), .B2(n4949), .A(n4948), .ZN(U3048) );
  INV_X1 U6107 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4953) );
  AOI22_X1 U6108 ( .A1(n6385), .A2(n4962), .B1(n5182), .B2(n6384), .ZN(n4950)
         );
  OAI21_X1 U6109 ( .B1(n6282), .B2(n4964), .A(n4950), .ZN(n4951) );
  AOI21_X1 U6110 ( .B1(n4966), .B2(n6279), .A(n4951), .ZN(n4952) );
  OAI21_X1 U6111 ( .B1(n4969), .B2(n4953), .A(n4952), .ZN(U3047) );
  INV_X1 U6112 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4957) );
  AOI22_X1 U6113 ( .A1(n6418), .A2(n4962), .B1(n5182), .B2(n6368), .ZN(n4954)
         );
  OAI21_X1 U6114 ( .B1(n6422), .B2(n4964), .A(n4954), .ZN(n4955) );
  AOI21_X1 U6115 ( .B1(n4966), .B2(n6421), .A(n4955), .ZN(n4956) );
  OAI21_X1 U6116 ( .B1(n4969), .B2(n4957), .A(n4956), .ZN(U3044) );
  INV_X1 U6117 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4961) );
  AOI22_X1 U6118 ( .A1(n6379), .A2(n4962), .B1(n5182), .B2(n6380), .ZN(n4958)
         );
  OAI21_X1 U6119 ( .B1(n6278), .B2(n4964), .A(n4958), .ZN(n4959) );
  AOI21_X1 U6120 ( .B1(n4966), .B2(n6339), .A(n4959), .ZN(n4960) );
  OAI21_X1 U6121 ( .B1(n4969), .B2(n4961), .A(n4960), .ZN(U3046) );
  INV_X1 U6122 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4968) );
  AOI22_X1 U6123 ( .A1(n6373), .A2(n4962), .B1(n5182), .B2(n6374), .ZN(n4963)
         );
  OAI21_X1 U6124 ( .B1(n6275), .B2(n4964), .A(n4963), .ZN(n4965) );
  AOI21_X1 U6125 ( .B1(n4966), .B2(n6335), .A(n4965), .ZN(n4967) );
  OAI21_X1 U6126 ( .B1(n4969), .B2(n4968), .A(n4967), .ZN(U3045) );
  AOI22_X1 U6127 ( .A1(n5244), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n6008), .ZN(n4970) );
  OAI21_X1 U6128 ( .B1(n5112), .B2(n5499), .A(n4970), .ZN(U2881) );
  INV_X1 U6129 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6616) );
  OAI222_X1 U6130 ( .A1(n4971), .A2(n5499), .B1(n5201), .B2(n6075), .C1(n5200), 
        .C2(n6616), .ZN(U2887) );
  INV_X1 U6131 ( .A(EAX_REG_3__SCAN_IN), .ZN(n4972) );
  OAI222_X1 U6132 ( .A1(n6123), .A2(n5499), .B1(n5201), .B2(n6073), .C1(n5200), 
        .C2(n4972), .ZN(U2888) );
  INV_X1 U6133 ( .A(DATAI_9_), .ZN(n6740) );
  INV_X1 U6134 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6023) );
  OAI222_X1 U6135 ( .A1(n5067), .A2(n5499), .B1(n5201), .B2(n6740), .C1(n5200), 
        .C2(n6023), .ZN(U2882) );
  INV_X1 U6136 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6028) );
  OAI222_X1 U6137 ( .A1(n5947), .A2(n5499), .B1(n5201), .B2(n6078), .C1(n5200), 
        .C2(n6028), .ZN(U2885) );
  INV_X1 U6138 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6039) );
  OAI222_X1 U6139 ( .A1(n6144), .A2(n5499), .B1(n5201), .B2(n6069), .C1(n5200), 
        .C2(n6039), .ZN(U2890) );
  INV_X1 U6140 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6035) );
  OAI222_X1 U6141 ( .A1(n4973), .A2(n5499), .B1(n5201), .B2(n6071), .C1(n5200), 
        .C2(n6035), .ZN(U2889) );
  INV_X1 U6142 ( .A(EAX_REG_0__SCAN_IN), .ZN(n4974) );
  OAI222_X1 U6143 ( .A1(n5008), .A2(n5499), .B1(n6067), .B2(n5201), .C1(n4974), 
        .C2(n5200), .ZN(U2891) );
  OAI21_X1 U6144 ( .B1(REIP_REG_8__SCAN_IN), .B2(n4975), .A(n5099), .ZN(n4983)
         );
  OAI22_X1 U6145 ( .A1(n6159), .A2(n5982), .B1(n5981), .B2(n4976), .ZN(n4977)
         );
  INV_X1 U6146 ( .A(n4977), .ZN(n4978) );
  OAI211_X1 U6147 ( .C1(n5963), .C2(n4979), .A(n4978), .B(n3095), .ZN(n4980)
         );
  AOI21_X1 U6148 ( .B1(n4981), .B2(n5968), .A(n4980), .ZN(n4982) );
  OAI211_X1 U6149 ( .C1(n5946), .C2(n4984), .A(n4983), .B(n4982), .ZN(U2819)
         );
  INV_X1 U6150 ( .A(DATAI_5_), .ZN(n4986) );
  OAI222_X1 U6151 ( .A1(n5200), .A2(n4987), .B1(n4986), .B2(n5201), .C1(n5499), 
        .C2(n4985), .ZN(U2886) );
  OAI21_X1 U6152 ( .B1(n4990), .B2(n4989), .A(n4988), .ZN(n6163) );
  NAND2_X1 U6153 ( .A1(n2971), .A2(REIP_REG_8__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U6154 ( .A1(n6142), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4991)
         );
  OAI211_X1 U6155 ( .C1(n6139), .C2(n4992), .A(n6160), .B(n4991), .ZN(n4993)
         );
  AOI21_X1 U6156 ( .B1(n4994), .B2(n6133), .A(n4993), .ZN(n4995) );
  OAI21_X1 U6157 ( .B1(n6163), .B2(n6137), .A(n4995), .ZN(U2978) );
  OAI21_X1 U6158 ( .B1(n4335), .B2(n4997), .A(n4996), .ZN(n5052) );
  AOI22_X1 U6159 ( .A1(n5244), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n6008), .ZN(n4998) );
  OAI21_X1 U6160 ( .B1(n5052), .B2(n5499), .A(n4998), .ZN(U2880) );
  INV_X1 U6161 ( .A(n5124), .ZN(n5000) );
  OAI222_X1 U6162 ( .A1(n5000), .A2(n5773), .B1(n4999), .B2(n5997), .C1(n5112), 
        .C2(n5480), .ZN(U2849) );
  NAND2_X1 U6163 ( .A1(n5001), .A2(n5357), .ZN(n5002) );
  NAND2_X1 U6164 ( .A1(n5946), .A2(n5002), .ZN(n5986) );
  INV_X1 U6165 ( .A(n5986), .ZN(n5020) );
  NOR2_X1 U6166 ( .A1(n5003), .A2(n6598), .ZN(n5984) );
  OAI22_X1 U6167 ( .A1(n4399), .A2(n5981), .B1(n5699), .B2(n5982), .ZN(n5005)
         );
  INV_X1 U6168 ( .A(n5423), .ZN(n5942) );
  INV_X1 U6169 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6593) );
  NOR2_X1 U6170 ( .A1(n5942), .A2(n6593), .ZN(n5004) );
  AOI211_X1 U6171 ( .C1(n5984), .C2(n3763), .A(n5005), .B(n5004), .ZN(n5007)
         );
  OAI21_X1 U6172 ( .B1(n5987), .B2(n5968), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5006) );
  OAI211_X1 U6173 ( .C1(n5020), .C2(n5008), .A(n5007), .B(n5006), .ZN(U2827)
         );
  INV_X1 U6174 ( .A(n6128), .ZN(n5014) );
  INV_X1 U6175 ( .A(n5984), .ZN(n5087) );
  NAND2_X1 U6176 ( .A1(n5987), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5010)
         );
  AOI22_X1 U6177 ( .A1(n6197), .A2(n5961), .B1(n5967), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n5009) );
  OAI211_X1 U6178 ( .C1(n6304), .C2(n5087), .A(n5010), .B(n5009), .ZN(n5013)
         );
  INV_X1 U6179 ( .A(n5971), .ZN(n5011) );
  OAI21_X1 U6180 ( .B1(n5090), .B2(n5011), .A(n5423), .ZN(n5965) );
  NOR2_X1 U6181 ( .A1(n5965), .A2(n6505), .ZN(n5012) );
  AOI211_X1 U6182 ( .C1(n5968), .C2(n5014), .A(n5013), .B(n5012), .ZN(n5019)
         );
  NAND2_X1 U6183 ( .A1(n5015), .A2(REIP_REG_1__SCAN_IN), .ZN(n5016) );
  NAND2_X1 U6184 ( .A1(n5423), .A2(n5016), .ZN(n5017) );
  NAND2_X1 U6185 ( .A1(n5017), .A2(REIP_REG_2__SCAN_IN), .ZN(n5979) );
  OR3_X1 U6186 ( .A1(n5979), .A2(n5971), .A3(n5977), .ZN(n5018) );
  OAI211_X1 U6187 ( .C1(n5020), .C2(n6123), .A(n5019), .B(n5018), .ZN(U2824)
         );
  OAI21_X1 U6188 ( .B1(n5029), .B2(n6602), .A(n6312), .ZN(n5027) );
  INV_X1 U6189 ( .A(n5021), .ZN(n5022) );
  NOR2_X1 U6190 ( .A1(n6356), .A2(n5025), .ZN(n5048) );
  AOI21_X1 U6191 ( .B1(n5022), .B2(n3763), .A(n5048), .ZN(n5026) );
  INV_X1 U6192 ( .A(n5026), .ZN(n5024) );
  AOI21_X1 U6193 ( .B1(n6364), .B2(n5025), .A(n6362), .ZN(n5023) );
  OAI21_X1 U6194 ( .B1(n5027), .B2(n5024), .A(n5023), .ZN(n5047) );
  OAI22_X1 U6195 ( .A1(n5027), .A2(n5026), .B1(n6601), .B2(n5025), .ZN(n5046)
         );
  AOI22_X1 U6196 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5047), .B1(n6421), 
        .B2(n5046), .ZN(n5031) );
  NOR2_X2 U6197 ( .A1(n5029), .A2(n5028), .ZN(n5173) );
  AOI22_X1 U6198 ( .A1(n5173), .A2(n6360), .B1(n6418), .B2(n5048), .ZN(n5030)
         );
  OAI211_X1 U6199 ( .C1(n6425), .C2(n5051), .A(n5031), .B(n5030), .ZN(U3028)
         );
  AOI22_X1 U6200 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n5047), .B1(n6286), 
        .B2(n5046), .ZN(n5033) );
  AOI22_X1 U6201 ( .A1(n5173), .A2(n6396), .B1(n6397), .B2(n5048), .ZN(n5032)
         );
  OAI211_X1 U6202 ( .C1(n5167), .C2(n5051), .A(n5033), .B(n5032), .ZN(U3033)
         );
  AOI22_X1 U6203 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n5047), .B1(n6290), 
        .B2(n5046), .ZN(n5035) );
  AOI22_X1 U6204 ( .A1(n5173), .A2(n6404), .B1(n6403), .B2(n5048), .ZN(n5034)
         );
  OAI211_X1 U6205 ( .C1(n5036), .C2(n5051), .A(n5035), .B(n5034), .ZN(U3034)
         );
  AOI22_X1 U6206 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5047), .B1(n6339), 
        .B2(n5046), .ZN(n5038) );
  AOI22_X1 U6207 ( .A1(n5173), .A2(n6378), .B1(n6379), .B2(n5048), .ZN(n5037)
         );
  OAI211_X1 U6208 ( .C1(n6342), .C2(n5051), .A(n5038), .B(n5037), .ZN(U3030)
         );
  AOI22_X1 U6209 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5047), .B1(n6279), 
        .B2(n5046), .ZN(n5040) );
  AOI22_X1 U6210 ( .A1(n5173), .A2(n6386), .B1(n6385), .B2(n5048), .ZN(n5039)
         );
  OAI211_X1 U6211 ( .C1(n5041), .C2(n5051), .A(n5040), .B(n5039), .ZN(U3031)
         );
  AOI22_X1 U6212 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5047), .B1(n6335), 
        .B2(n5046), .ZN(n5043) );
  AOI22_X1 U6213 ( .A1(n5173), .A2(n6372), .B1(n6373), .B2(n5048), .ZN(n5042)
         );
  OAI211_X1 U6214 ( .C1(n6338), .C2(n5051), .A(n5043), .B(n5042), .ZN(U3029)
         );
  AOI22_X1 U6215 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n5047), .B1(n6350), 
        .B2(n5046), .ZN(n5045) );
  AOI22_X1 U6216 ( .A1(n5173), .A2(n6783), .B1(n2999), .B2(n5048), .ZN(n5044)
         );
  OAI211_X1 U6217 ( .C1(n6778), .C2(n5051), .A(n5045), .B(n5044), .ZN(U3035)
         );
  AOI22_X1 U6218 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5047), .B1(n6343), 
        .B2(n5046), .ZN(n5050) );
  AOI22_X1 U6219 ( .A1(n5173), .A2(n6392), .B1(n6391), .B2(n5048), .ZN(n5049)
         );
  OAI211_X1 U6220 ( .C1(n6346), .C2(n5051), .A(n5050), .B(n5049), .ZN(U3032)
         );
  INV_X1 U6221 ( .A(n5052), .ZN(n5135) );
  INV_X1 U6222 ( .A(n5053), .ZN(n5071) );
  NAND2_X1 U6223 ( .A1(n5055), .A2(n5054), .ZN(n5056) );
  NAND2_X1 U6224 ( .A1(n5071), .A2(n5056), .ZN(n6147) );
  OAI22_X1 U6225 ( .A1(n5773), .A2(n6147), .B1(n5057), .B2(n5997), .ZN(n5058)
         );
  AOI21_X1 U6226 ( .B1(n5135), .B2(n4286), .A(n5058), .ZN(n5059) );
  INV_X1 U6227 ( .A(n5059), .ZN(U2848) );
  NAND2_X1 U6228 ( .A1(n5061), .A2(n5060), .ZN(n5062) );
  XNOR2_X1 U6229 ( .A(n5063), .B(n5062), .ZN(n6155) );
  NAND2_X1 U6230 ( .A1(n6155), .A2(n4310), .ZN(n5066) );
  AND2_X1 U6231 ( .A1(n2971), .A2(REIP_REG_9__SCAN_IN), .ZN(n6152) );
  NOR2_X1 U6232 ( .A1(n6139), .A2(n5097), .ZN(n5064) );
  AOI211_X1 U6233 ( .C1(n6142), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6152), 
        .B(n5064), .ZN(n5065) );
  OAI211_X1 U6234 ( .C1(n6145), .C2(n5067), .A(n5066), .B(n5065), .ZN(U2977)
         );
  AOI21_X1 U6235 ( .B1(n5069), .B2(n4996), .A(n5068), .ZN(n5920) );
  INV_X1 U6236 ( .A(n5920), .ZN(n5075) );
  AOI21_X1 U6237 ( .B1(n5072), .B2(n5071), .A(n5070), .ZN(n5921) );
  AOI22_X1 U6238 ( .A1(n5921), .A2(n5995), .B1(n5490), .B2(EBX_REG_12__SCAN_IN), .ZN(n5073) );
  OAI21_X1 U6239 ( .B1(n5075), .B2(n5480), .A(n5073), .ZN(U2847) );
  INV_X1 U6240 ( .A(DATAI_12_), .ZN(n6060) );
  OAI222_X1 U6241 ( .A1(n5075), .A2(n5499), .B1(n6060), .B2(n5201), .C1(n5074), 
        .C2(n5200), .ZN(U2879) );
  NAND3_X1 U6242 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .A3(
        REIP_REG_10__SCAN_IN), .ZN(n5191) );
  NOR2_X1 U6243 ( .A1(n5076), .A2(n5191), .ZN(n5209) );
  NOR2_X1 U6244 ( .A1(n5942), .A2(n5209), .ZN(n5926) );
  NAND2_X1 U6245 ( .A1(n5926), .A2(REIP_REG_11__SCAN_IN), .ZN(n5080) );
  AOI21_X1 U6246 ( .B1(n5967), .B2(EBX_REG_11__SCAN_IN), .A(n2971), .ZN(n5077)
         );
  OAI21_X1 U6247 ( .B1(n6147), .B2(n5982), .A(n5077), .ZN(n5078) );
  AOI21_X1 U6248 ( .B1(n5987), .B2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n5078), 
        .ZN(n5079) );
  OAI211_X1 U6249 ( .C1(n5993), .C2(n5133), .A(n5080), .B(n5079), .ZN(n5083)
         );
  NAND2_X1 U6250 ( .A1(REIP_REG_9__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .ZN(
        n5081) );
  NOR3_X1 U6251 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5081), .A3(n5190), .ZN(n5082) );
  AOI211_X1 U6252 ( .C1(n5135), .C2(n5937), .A(n5083), .B(n5082), .ZN(n5084)
         );
  INV_X1 U6253 ( .A(n5084), .ZN(U2816) );
  INV_X1 U6254 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5094) );
  INV_X1 U6255 ( .A(n5977), .ZN(n5972) );
  AOI22_X1 U6256 ( .A1(n5967), .A2(EBX_REG_1__SCAN_IN), .B1(n5972), .B2(n6587), 
        .ZN(n5086) );
  NAND2_X1 U6257 ( .A1(n4417), .A2(n5961), .ZN(n5085) );
  OAI211_X1 U6258 ( .C1(n5715), .C2(n5087), .A(n5086), .B(n5085), .ZN(n5089)
         );
  NOR2_X1 U6259 ( .A1(n5993), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5088)
         );
  AOI211_X1 U6260 ( .C1(n5090), .C2(REIP_REG_1__SCAN_IN), .A(n5089), .B(n5088), 
        .ZN(n5093) );
  INV_X1 U6261 ( .A(n6144), .ZN(n5091) );
  NAND2_X1 U6262 ( .A1(n5986), .A2(n5091), .ZN(n5092) );
  OAI211_X1 U6263 ( .C1(n5094), .C2(n5963), .A(n5093), .B(n5092), .ZN(U2826)
         );
  INV_X1 U6264 ( .A(n5095), .ZN(n5106) );
  OAI22_X1 U6265 ( .A1(n5993), .A2(n5097), .B1(n5096), .B2(n5981), .ZN(n5103)
         );
  INV_X1 U6266 ( .A(n5098), .ZN(n6153) );
  AOI22_X1 U6267 ( .A1(n5099), .A2(REIP_REG_9__SCAN_IN), .B1(n5961), .B2(n6153), .ZN(n5100) );
  OAI211_X1 U6268 ( .C1(n5963), .C2(n5101), .A(n5100), .B(n3095), .ZN(n5102)
         );
  AOI211_X1 U6269 ( .C1(n5104), .C2(n5937), .A(n5103), .B(n5102), .ZN(n5105)
         );
  NAND2_X1 U6270 ( .A1(n5106), .A2(n5105), .ZN(U2818) );
  NAND2_X1 U6271 ( .A1(n5128), .A2(n5107), .ZN(n5109) );
  XOR2_X1 U6272 ( .A(n5109), .B(n5108), .Z(n5127) );
  AND2_X1 U6273 ( .A1(n2971), .A2(REIP_REG_10__SCAN_IN), .ZN(n5123) );
  AND2_X1 U6274 ( .A1(n6142), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5110)
         );
  AOI211_X1 U6275 ( .C1(n5821), .C2(n5111), .A(n5123), .B(n5110), .ZN(n5115)
         );
  INV_X1 U6276 ( .A(n5112), .ZN(n5113) );
  NAND2_X1 U6277 ( .A1(n5113), .A2(n6133), .ZN(n5114) );
  OAI211_X1 U6278 ( .C1(n5127), .C2(n6137), .A(n5115), .B(n5114), .ZN(U2976)
         );
  AOI22_X1 U6279 ( .A1(n5684), .A2(n5117), .B1(n5655), .B2(n5116), .ZN(n6176)
         );
  OAI21_X1 U6280 ( .B1(n5686), .B2(n6164), .A(n6176), .ZN(n6154) );
  AOI21_X1 U6281 ( .B1(n5683), .B2(n6209), .A(n5118), .ZN(n6187) );
  NOR2_X1 U6282 ( .A1(n5688), .A2(n5119), .ZN(n5685) );
  NAND2_X1 U6283 ( .A1(n6187), .A2(n5685), .ZN(n6186) );
  NOR2_X1 U6284 ( .A1(n5120), .A2(n6186), .ZN(n6172) );
  NAND2_X1 U6285 ( .A1(n6164), .A2(n6172), .ZN(n6158) );
  AOI221_X1 U6286 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n5121), .C2(n3516), .A(n6158), 
        .ZN(n5122) );
  AOI21_X1 U6287 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6154), .A(n5122), 
        .ZN(n5126) );
  AOI21_X1 U6288 ( .B1(n4302), .B2(n5124), .A(n5123), .ZN(n5125) );
  OAI211_X1 U6289 ( .C1(n5127), .C2(n6198), .A(n5126), .B(n5125), .ZN(U3008)
         );
  NAND2_X1 U6290 ( .A1(n5129), .A2(n5128), .ZN(n5131) );
  XNOR2_X1 U6291 ( .A(n5539), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5130)
         );
  XNOR2_X1 U6292 ( .A(n5131), .B(n5130), .ZN(n6146) );
  AOI22_X1 U6293 ( .A1(n6142), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .B1(n2971), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n5132) );
  OAI21_X1 U6294 ( .B1(n5133), .B2(n6139), .A(n5132), .ZN(n5134) );
  AOI21_X1 U6295 ( .B1(n5135), .B2(n6133), .A(n5134), .ZN(n5136) );
  OAI21_X1 U6296 ( .B1(n6146), .B2(n6137), .A(n5136), .ZN(U2975) );
  NOR2_X1 U6297 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5137), .ZN(n5143)
         );
  OAI21_X1 U6298 ( .B1(n5173), .B2(n5182), .A(n5138), .ZN(n5140) );
  NAND2_X1 U6299 ( .A1(n5140), .A2(n5139), .ZN(n5142) );
  OAI221_X1 U6300 ( .B1(n5143), .B2(n6718), .C1(n5143), .C2(n5142), .A(n5141), 
        .ZN(n5177) );
  NAND2_X1 U6301 ( .A1(n5177), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5150) );
  INV_X1 U6302 ( .A(n5143), .ZN(n5178) );
  INV_X1 U6303 ( .A(n5144), .ZN(n5145) );
  NOR2_X1 U6304 ( .A1(n5145), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6263)
         );
  AOI22_X1 U6305 ( .A1(n5146), .A2(n6312), .B1(n6267), .B2(n6263), .ZN(n5185)
         );
  OAI22_X1 U6306 ( .A1(n5147), .A2(n5178), .B1(n5185), .B2(n6389), .ZN(n5148)
         );
  AOI21_X1 U6307 ( .B1(n6384), .B2(n5173), .A(n5148), .ZN(n5149) );
  OAI211_X1 U6308 ( .C1(n5176), .C2(n6282), .A(n5150), .B(n5149), .ZN(U3039)
         );
  NAND2_X1 U6309 ( .A1(n5177), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5154) );
  OAI22_X1 U6310 ( .A1(n5151), .A2(n5178), .B1(n5185), .B2(n6377), .ZN(n5152)
         );
  AOI21_X1 U6311 ( .B1(n6374), .B2(n5173), .A(n5152), .ZN(n5153) );
  OAI211_X1 U6312 ( .C1(n6275), .C2(n5176), .A(n5154), .B(n5153), .ZN(U3037)
         );
  NAND2_X1 U6313 ( .A1(n5177), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5158) );
  OAI22_X1 U6314 ( .A1(n5155), .A2(n5178), .B1(n5185), .B2(n6395), .ZN(n5156)
         );
  AOI21_X1 U6315 ( .B1(n6390), .B2(n5173), .A(n5156), .ZN(n5157) );
  OAI211_X1 U6316 ( .C1(n5176), .C2(n6285), .A(n5158), .B(n5157), .ZN(U3040)
         );
  NAND2_X1 U6317 ( .A1(n5177), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5161) );
  INV_X1 U6318 ( .A(n5173), .ZN(n5180) );
  OAI22_X1 U6319 ( .A1(n6778), .A2(n5180), .B1(n6780), .B2(n5178), .ZN(n5159)
         );
  AOI21_X1 U6320 ( .B1(n6783), .B2(n5182), .A(n5159), .ZN(n5160) );
  OAI211_X1 U6321 ( .C1(n5185), .C2(n6786), .A(n5161), .B(n5160), .ZN(U3043)
         );
  NAND2_X1 U6322 ( .A1(n5177), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5165) );
  OAI22_X1 U6323 ( .A1(n5162), .A2(n5178), .B1(n5185), .B2(n6383), .ZN(n5163)
         );
  AOI21_X1 U6324 ( .B1(n6380), .B2(n5173), .A(n5163), .ZN(n5164) );
  OAI211_X1 U6325 ( .C1(n5176), .C2(n6278), .A(n5165), .B(n5164), .ZN(U3038)
         );
  NAND2_X1 U6326 ( .A1(n5177), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5170) );
  OAI22_X1 U6327 ( .A1(n5167), .A2(n5180), .B1(n5166), .B2(n5178), .ZN(n5168)
         );
  AOI21_X1 U6328 ( .B1(n6396), .B2(n5182), .A(n5168), .ZN(n5169) );
  OAI211_X1 U6329 ( .C1(n5185), .C2(n6401), .A(n5170), .B(n5169), .ZN(U3041)
         );
  NAND2_X1 U6330 ( .A1(n5177), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5175) );
  OAI22_X1 U6331 ( .A1(n5171), .A2(n5178), .B1(n5185), .B2(n6407), .ZN(n5172)
         );
  AOI21_X1 U6332 ( .B1(n6402), .B2(n5173), .A(n5172), .ZN(n5174) );
  OAI211_X1 U6333 ( .C1(n5176), .C2(n6293), .A(n5175), .B(n5174), .ZN(U3042)
         );
  NAND2_X1 U6334 ( .A1(n5177), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5184) );
  OAI22_X1 U6335 ( .A1(n6425), .A2(n5180), .B1(n5179), .B2(n5178), .ZN(n5181)
         );
  AOI21_X1 U6336 ( .B1(n6360), .B2(n5182), .A(n5181), .ZN(n5183) );
  OAI211_X1 U6337 ( .C1(n5185), .C2(n6371), .A(n5184), .B(n5183), .ZN(U3036)
         );
  OAI21_X1 U6338 ( .B1(n5186), .B2(n5189), .A(n5188), .ZN(n5248) );
  NAND2_X1 U6339 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n5208) );
  OAI211_X1 U6340 ( .C1(REIP_REG_13__SCAN_IN), .C2(REIP_REG_12__SCAN_IN), .A(
        n5925), .B(n5208), .ZN(n5199) );
  OAI21_X1 U6341 ( .B1(n5070), .B2(n5193), .A(n5192), .ZN(n5264) );
  NOR2_X1 U6342 ( .A1(n5264), .A2(n5982), .ZN(n5194) );
  AOI211_X1 U6343 ( .C1(n5967), .C2(EBX_REG_13__SCAN_IN), .A(n2971), .B(n5194), 
        .ZN(n5196) );
  NAND2_X1 U6344 ( .A1(n5987), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5195)
         );
  OAI211_X1 U6345 ( .C1(n5993), .C2(n5250), .A(n5196), .B(n5195), .ZN(n5197)
         );
  AOI21_X1 U6346 ( .B1(n5926), .B2(REIP_REG_13__SCAN_IN), .A(n5197), .ZN(n5198) );
  OAI211_X1 U6347 ( .C1(n5248), .C2(n5946), .A(n5199), .B(n5198), .ZN(U2814)
         );
  INV_X1 U6348 ( .A(DATAI_13_), .ZN(n6096) );
  INV_X1 U6349 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6018) );
  OAI222_X1 U6350 ( .A1(n5248), .A2(n5499), .B1(n5201), .B2(n6096), .C1(n6018), 
        .C2(n5200), .ZN(U2878) );
  INV_X1 U6351 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5202) );
  OAI222_X1 U6352 ( .A1(n5264), .A2(n5773), .B1(n5997), .B2(n5202), .C1(n5480), 
        .C2(n5248), .ZN(U2846) );
  INV_X1 U6353 ( .A(n5203), .ZN(n5207) );
  NAND3_X1 U6354 ( .A1(n5188), .A2(n5205), .A3(n5204), .ZN(n5206) );
  NAND2_X1 U6355 ( .A1(n5207), .A2(n5206), .ZN(n5286) );
  NOR2_X1 U6356 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5208), .ZN(n5217) );
  INV_X1 U6357 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6525) );
  NAND4_X1 U6358 ( .A1(n5209), .A2(REIP_REG_14__SCAN_IN), .A3(
        REIP_REG_13__SCAN_IN), .A4(REIP_REG_12__SCAN_IN), .ZN(n5331) );
  NAND2_X1 U6359 ( .A1(n5331), .A2(n5423), .ZN(n5910) );
  NAND2_X1 U6360 ( .A1(n5192), .A2(n5210), .ZN(n5211) );
  NAND2_X1 U6361 ( .A1(n5241), .A2(n5211), .ZN(n5860) );
  INV_X1 U6362 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5236) );
  OAI22_X1 U6363 ( .A1(n5860), .A2(n5982), .B1(n5981), .B2(n5236), .ZN(n5212)
         );
  INV_X1 U6364 ( .A(n5212), .ZN(n5213) );
  OAI21_X1 U6365 ( .B1(n6525), .B2(n5910), .A(n5213), .ZN(n5216) );
  AOI21_X1 U6366 ( .B1(n5987), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n2971), 
        .ZN(n5214) );
  OAI21_X1 U6367 ( .B1(n5993), .B2(n5282), .A(n5214), .ZN(n5215) );
  AOI211_X1 U6368 ( .C1(n5925), .C2(n5217), .A(n5216), .B(n5215), .ZN(n5218)
         );
  OAI21_X1 U6369 ( .B1(n5286), .B2(n5946), .A(n5218), .ZN(U2813) );
  AOI22_X1 U6370 ( .A1(n5244), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n6008), .ZN(n5219) );
  OAI21_X1 U6371 ( .B1(n5286), .B2(n5499), .A(n5219), .ZN(U2877) );
  INV_X1 U6372 ( .A(n5221), .ZN(n5222) );
  NOR2_X1 U6373 ( .A1(n5223), .A2(n5222), .ZN(n5224) );
  XNOR2_X1 U6374 ( .A(n5220), .B(n5224), .ZN(n5235) );
  AND2_X1 U6375 ( .A1(n2971), .A2(REIP_REG_12__SCAN_IN), .ZN(n5232) );
  AOI21_X1 U6376 ( .B1(n4302), .B2(n5921), .A(n5232), .ZN(n5230) );
  INV_X1 U6377 ( .A(n6150), .ZN(n5301) );
  AOI21_X1 U6378 ( .B1(n5225), .B2(n6209), .A(n5259), .ZN(n5228) );
  OAI21_X1 U6379 ( .B1(n6151), .B2(n3517), .A(n5226), .ZN(n5227) );
  OAI21_X1 U6380 ( .B1(n5301), .B2(n5228), .A(n5227), .ZN(n5229) );
  OAI211_X1 U6381 ( .C1(n5235), .C2(n6198), .A(n5230), .B(n5229), .ZN(U3006)
         );
  NOR2_X1 U6382 ( .A1(n5824), .A2(n5923), .ZN(n5231) );
  AOI211_X1 U6383 ( .C1(n5821), .C2(n5919), .A(n5232), .B(n5231), .ZN(n5234)
         );
  NAND2_X1 U6384 ( .A1(n5920), .A2(n6133), .ZN(n5233) );
  OAI211_X1 U6385 ( .C1(n5235), .C2(n6137), .A(n5234), .B(n5233), .ZN(U2974)
         );
  OAI222_X1 U6386 ( .A1(n5860), .A2(n5773), .B1(n5236), .B2(n5997), .C1(n5480), 
        .C2(n5286), .ZN(U2845) );
  NOR2_X1 U6387 ( .A1(n2974), .A2(n5238), .ZN(n5239) );
  OR2_X1 U6388 ( .A1(n5237), .A2(n5239), .ZN(n5913) );
  AND2_X1 U6389 ( .A1(n5241), .A2(n5240), .ZN(n5242) );
  NOR2_X1 U6390 ( .A1(n5274), .A2(n5242), .ZN(n5908) );
  AOI22_X1 U6391 ( .A1(n5908), .A2(n5995), .B1(EBX_REG_15__SCAN_IN), .B2(n5490), .ZN(n5243) );
  OAI21_X1 U6392 ( .B1(n5913), .B2(n5480), .A(n5243), .ZN(U2844) );
  AOI22_X1 U6393 ( .A1(n5244), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6008), .ZN(n5245) );
  OAI21_X1 U6394 ( .B1(n5913), .B2(n5499), .A(n5245), .ZN(U2876) );
  XOR2_X1 U6395 ( .A(n5246), .B(n5247), .Z(n5269) );
  INV_X1 U6396 ( .A(n5248), .ZN(n5252) );
  AOI22_X1 U6397 ( .A1(n6142), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .B1(n2971), 
        .B2(REIP_REG_13__SCAN_IN), .ZN(n5249) );
  OAI21_X1 U6398 ( .B1(n5250), .B2(n6139), .A(n5249), .ZN(n5251) );
  AOI21_X1 U6399 ( .B1(n5252), .B2(n6133), .A(n5251), .ZN(n5253) );
  OAI21_X1 U6400 ( .B1(n5269), .B2(n6137), .A(n5253), .ZN(U2973) );
  NAND3_X1 U6401 ( .A1(n5255), .A2(n5254), .A3(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5256) );
  INV_X1 U6402 ( .A(n5259), .ZN(n5262) );
  AOI211_X1 U6403 ( .C1(n5257), .C2(n5256), .A(INSTADDRPOINTER_REG_13__SCAN_IN), .B(n5262), .ZN(n5261) );
  AOI211_X1 U6404 ( .C1(n5702), .C2(n5859), .A(n5261), .B(n5301), .ZN(n5258)
         );
  OAI21_X1 U6405 ( .B1(n5260), .B2(n5259), .A(n5258), .ZN(n5863) );
  OAI21_X1 U6406 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5261), .A(n5863), 
        .ZN(n5268) );
  NOR3_X1 U6407 ( .A1(n5263), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n5262), 
        .ZN(n5266) );
  INV_X1 U6408 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6523) );
  OAI22_X1 U6409 ( .A1(n6213), .A2(n5264), .B1(n6523), .B2(n3095), .ZN(n5265)
         );
  AOI21_X1 U6410 ( .B1(n5702), .B2(n5266), .A(n5265), .ZN(n5267) );
  OAI211_X1 U6411 ( .C1(n5269), .C2(n6198), .A(n5268), .B(n5267), .ZN(U3005)
         );
  OR2_X1 U6412 ( .A1(n5237), .A2(n5271), .ZN(n5272) );
  AND2_X1 U6413 ( .A1(n5270), .A2(n5272), .ZN(n6007) );
  INV_X1 U6414 ( .A(n6007), .ZN(n5277) );
  INV_X1 U6415 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5276) );
  NOR2_X1 U6416 ( .A1(n5274), .A2(n5273), .ZN(n5275) );
  OR2_X1 U6417 ( .A1(n5292), .A2(n5275), .ZN(n5853) );
  OAI222_X1 U6418 ( .A1(n5277), .A2(n5480), .B1(n5997), .B2(n5276), .C1(n5853), 
        .C2(n5773), .ZN(U2843) );
  NOR2_X1 U6419 ( .A1(n3074), .A2(n5280), .ZN(n5281) );
  XNOR2_X1 U6420 ( .A(n5278), .B(n5281), .ZN(n5864) );
  NAND2_X1 U6421 ( .A1(n5864), .A2(n4310), .ZN(n5285) );
  AND2_X1 U6422 ( .A1(n2971), .A2(REIP_REG_14__SCAN_IN), .ZN(n5861) );
  NOR2_X1 U6423 ( .A1(n6139), .A2(n5282), .ZN(n5283) );
  AOI211_X1 U6424 ( .C1(n6142), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5861), 
        .B(n5283), .ZN(n5284) );
  OAI211_X1 U6425 ( .C1(n6145), .C2(n5286), .A(n5285), .B(n5284), .ZN(U2972)
         );
  NAND2_X1 U6426 ( .A1(n5270), .A2(n5288), .ZN(n5289) );
  AND2_X1 U6427 ( .A1(n5287), .A2(n5289), .ZN(n6002) );
  OR2_X1 U6428 ( .A1(n5292), .A2(n5291), .ZN(n5293) );
  NAND2_X1 U6429 ( .A1(n5290), .A2(n5293), .ZN(n5842) );
  OAI22_X1 U6430 ( .A1(n5842), .A2(n5773), .B1(n5294), .B2(n5997), .ZN(n5295)
         );
  AOI21_X1 U6431 ( .B1(n6002), .B2(n4286), .A(n5295), .ZN(n5296) );
  INV_X1 U6432 ( .A(n5296), .ZN(U2842) );
  XNOR2_X1 U6433 ( .A(n5539), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5297)
         );
  XNOR2_X1 U6434 ( .A(n5298), .B(n5297), .ZN(n5311) );
  NOR3_X1 U6435 ( .A1(n6151), .A2(n5859), .A3(n5299), .ZN(n5851) );
  INV_X1 U6436 ( .A(n5300), .ZN(n5302) );
  AOI21_X1 U6437 ( .B1(n5303), .B2(n5302), .A(n5301), .ZN(n5858) );
  NAND2_X1 U6438 ( .A1(n2971), .A2(REIP_REG_15__SCAN_IN), .ZN(n5307) );
  NAND2_X1 U6439 ( .A1(n5908), .A2(n4302), .ZN(n5304) );
  OAI211_X1 U6440 ( .C1(n5858), .C2(n5849), .A(n5307), .B(n5304), .ZN(n5305)
         );
  AOI21_X1 U6441 ( .B1(n5851), .B2(n5849), .A(n5305), .ZN(n5306) );
  OAI21_X1 U6442 ( .B1(n5311), .B2(n6198), .A(n5306), .ZN(U3003) );
  OAI21_X1 U6443 ( .B1(n5824), .B2(n5907), .A(n5307), .ZN(n5308) );
  AOI21_X1 U6444 ( .B1(n5821), .B2(n5914), .A(n5308), .ZN(n5310) );
  OR2_X1 U6445 ( .A1(n5913), .A2(n6145), .ZN(n5309) );
  OAI211_X1 U6446 ( .C1(n5311), .C2(n6137), .A(n5310), .B(n5309), .ZN(U2971)
         );
  NAND2_X1 U6447 ( .A1(n5287), .A2(n5313), .ZN(n5314) );
  AND2_X1 U6448 ( .A1(n5486), .A2(n5314), .ZN(n5999) );
  INV_X1 U6449 ( .A(n5999), .ZN(n5322) );
  MUX2_X1 U6450 ( .A(n5316), .B(n5315), .S(n2983), .Z(n5317) );
  INV_X1 U6451 ( .A(n5317), .ZN(n5318) );
  OR2_X1 U6452 ( .A1(n5290), .A2(n5318), .ZN(n5489) );
  NAND2_X1 U6453 ( .A1(n5290), .A2(n5318), .ZN(n5319) );
  INV_X1 U6454 ( .A(n5895), .ZN(n5320) );
  OAI222_X1 U6455 ( .A1(n5322), .A2(n5480), .B1(n5997), .B2(n5321), .C1(n5320), 
        .C2(n5773), .ZN(U2841) );
  NAND2_X1 U6456 ( .A1(n5821), .A2(n5341), .ZN(n5324) );
  OAI211_X1 U6457 ( .C1(n5824), .C2(n5325), .A(n5324), .B(n5323), .ZN(n5326)
         );
  OAI21_X1 U6458 ( .B1(n5329), .B2(n6137), .A(n5328), .ZN(U2956) );
  AND2_X1 U6459 ( .A1(REIP_REG_26__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5330) );
  OR2_X1 U6460 ( .A1(n5977), .A2(n5330), .ZN(n5333) );
  INV_X1 U6461 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6531) );
  NAND2_X1 U6462 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n5899) );
  NOR3_X1 U6463 ( .A1(n6531), .A2(n5331), .A3(n5899), .ZN(n5446) );
  NAND4_X1 U6464 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5446), .A3(
        REIP_REG_19__SCAN_IN), .A4(REIP_REG_18__SCAN_IN), .ZN(n5422) );
  NAND3_X1 U6465 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5332) );
  OAI21_X1 U6466 ( .B1(n5422), .B2(n5332), .A(n5423), .ZN(n5753) );
  NAND2_X1 U6467 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5766) );
  NOR2_X2 U6468 ( .A1(n5332), .A2(n5441), .ZN(n5339) );
  INV_X1 U6469 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U6470 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5340) );
  INV_X1 U6471 ( .A(n5340), .ZN(n5334) );
  OR2_X1 U6472 ( .A1(n5977), .A2(n5334), .ZN(n5335) );
  NAND2_X1 U6473 ( .A1(n5734), .A2(n5335), .ZN(n5387) );
  INV_X1 U6474 ( .A(n5387), .ZN(n5338) );
  INV_X1 U6475 ( .A(REIP_REG_30__SCAN_IN), .ZN(n5337) );
  OAI22_X1 U6476 ( .A1(n5338), .A2(n5337), .B1(n5981), .B2(n5336), .ZN(n5345)
         );
  NAND2_X1 U6477 ( .A1(n5339), .A2(REIP_REG_24__SCAN_IN), .ZN(n5742) );
  NAND3_X1 U6478 ( .A1(REIP_REG_26__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .A3(
        n5393), .ZN(n5724) );
  NOR2_X2 U6479 ( .A1(n5724), .A2(n5340), .ZN(n5376) );
  NAND2_X1 U6480 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .ZN(
        n5361) );
  OAI211_X1 U6481 ( .C1(REIP_REG_30__SCAN_IN), .C2(REIP_REG_29__SCAN_IN), .A(
        n5376), .B(n5361), .ZN(n5343) );
  AOI22_X1 U6482 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n5987), .B1(n5341), 
        .B2(n5968), .ZN(n5342) );
  NAND2_X1 U6483 ( .A1(n5343), .A2(n5342), .ZN(n5344) );
  AOI211_X1 U6484 ( .C1(n5961), .C2(n5346), .A(n5345), .B(n5344), .ZN(n5347)
         );
  OAI21_X1 U6485 ( .B1(n5348), .B2(n5946), .A(n5347), .ZN(U2797) );
  NAND2_X1 U6486 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5718) );
  AOI22_X1 U6487 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5349), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6215), .ZN(n5721) );
  OR2_X1 U6488 ( .A1(n5718), .A2(n5721), .ZN(n5351) );
  INV_X1 U6489 ( .A(n6578), .ZN(n6569) );
  NAND3_X1 U6490 ( .A1(n5714), .A2(n3771), .A3(n6569), .ZN(n5350) );
  NAND2_X1 U6491 ( .A1(n5351), .A2(n5350), .ZN(n5352) );
  AOI21_X1 U6492 ( .B1(n5353), .B2(n6571), .A(n5352), .ZN(n5355) );
  NOR2_X1 U6493 ( .A1(n5714), .A2(n6578), .ZN(n5720) );
  OAI21_X1 U6494 ( .B1(n6583), .B2(n5720), .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .ZN(n5354) );
  OAI21_X1 U6495 ( .B1(n6583), .B2(n5355), .A(n5354), .ZN(U3459) );
  INV_X1 U6496 ( .A(n2976), .ZN(n5366) );
  AOI21_X1 U6497 ( .B1(n5972), .B2(n5361), .A(n5387), .ZN(n5360) );
  INV_X1 U6498 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6558) );
  NAND2_X1 U6499 ( .A1(n5987), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5359)
         );
  NAND4_X1 U6500 ( .A1(n2984), .A2(EBX_REG_31__SCAN_IN), .A3(n6464), .A4(n5357), .ZN(n5358) );
  OAI211_X1 U6501 ( .C1(n5360), .C2(n6558), .A(n5359), .B(n5358), .ZN(n5364)
         );
  INV_X1 U6502 ( .A(n5376), .ZN(n5362) );
  NOR3_X1 U6503 ( .A1(n5362), .A2(REIP_REG_31__SCAN_IN), .A3(n5361), .ZN(n5363) );
  AOI211_X1 U6504 ( .C1(n5454), .C2(n5961), .A(n5364), .B(n5363), .ZN(n5365)
         );
  OAI21_X1 U6505 ( .B1(n5366), .B2(n5946), .A(n5365), .ZN(U2796) );
  NAND2_X1 U6506 ( .A1(n5367), .A2(n5368), .ZN(n5369) );
  INV_X1 U6507 ( .A(n5780), .ZN(n5458) );
  INV_X1 U6508 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6554) );
  XNOR2_X1 U6509 ( .A(n5385), .B(n5371), .ZN(n5590) );
  AOI22_X1 U6510 ( .A1(EBX_REG_29__SCAN_IN), .A2(n5967), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n5987), .ZN(n5372) );
  OAI21_X1 U6511 ( .B1(n5503), .B2(n5993), .A(n5372), .ZN(n5373) );
  AOI21_X1 U6512 ( .B1(REIP_REG_29__SCAN_IN), .B2(n5387), .A(n5373), .ZN(n5374) );
  OAI21_X1 U6513 ( .B1(n5590), .B2(n5982), .A(n5374), .ZN(n5375) );
  AOI21_X1 U6514 ( .B1(n5376), .B2(n6554), .A(n5375), .ZN(n5377) );
  OAI21_X1 U6515 ( .B1(n5458), .B2(n5946), .A(n5377), .ZN(U2798) );
  OR2_X1 U6516 ( .A1(n5379), .A2(n5380), .ZN(n5381) );
  INV_X1 U6517 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6547) );
  NOR3_X1 U6518 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6547), .A3(n5724), .ZN(n5391) );
  OR2_X1 U6519 ( .A1(n5382), .A2(n5383), .ZN(n5384) );
  NAND2_X1 U6520 ( .A1(n5385), .A2(n5384), .ZN(n5600) );
  OAI22_X1 U6521 ( .A1(n5459), .A2(n5981), .B1(n5513), .B2(n5963), .ZN(n5386)
         );
  AOI21_X1 U6522 ( .B1(n5387), .B2(REIP_REG_28__SCAN_IN), .A(n5386), .ZN(n5389) );
  NAND2_X1 U6523 ( .A1(n5968), .A2(n5511), .ZN(n5388) );
  OAI211_X1 U6524 ( .C1(n5600), .C2(n5982), .A(n5389), .B(n5388), .ZN(n5390)
         );
  AOI211_X1 U6525 ( .C1(n5783), .C2(n5937), .A(n5391), .B(n5390), .ZN(n5392)
         );
  INV_X1 U6526 ( .A(n5392), .ZN(U2799) );
  AOI21_X1 U6527 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5393), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5404) );
  INV_X1 U6528 ( .A(n2973), .ZN(n5463) );
  INV_X1 U6529 ( .A(n5395), .ZN(n5396) );
  AOI21_X1 U6530 ( .B1(n5397), .B2(n5463), .A(n5396), .ZN(n5532) );
  NAND2_X1 U6531 ( .A1(n5532), .A2(n5937), .ZN(n5403) );
  INV_X1 U6532 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6625) );
  OAI22_X1 U6533 ( .A1(n6625), .A2(n5981), .B1(n5530), .B2(n5963), .ZN(n5401)
         );
  AND2_X1 U6534 ( .A1(n5466), .A2(n5398), .ZN(n5399) );
  NOR2_X1 U6535 ( .A1(n5605), .A2(n5399), .ZN(n5615) );
  INV_X1 U6536 ( .A(n5615), .ZN(n5462) );
  NOR2_X1 U6537 ( .A1(n5462), .A2(n5982), .ZN(n5400) );
  AOI211_X1 U6538 ( .C1(n5968), .C2(n5528), .A(n5401), .B(n5400), .ZN(n5402)
         );
  OAI211_X1 U6539 ( .C1(n5734), .C2(n5404), .A(n5403), .B(n5402), .ZN(U2801)
         );
  OAI21_X1 U6540 ( .B1(n5405), .B2(n5407), .A(n5406), .ZN(n5471) );
  OR2_X1 U6541 ( .A1(n5409), .A2(n5410), .ZN(n5411) );
  NAND2_X1 U6542 ( .A1(n5408), .A2(n5411), .ZN(n5625) );
  INV_X1 U6543 ( .A(n5625), .ZN(n5415) );
  AOI22_X1 U6544 ( .A1(n5987), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .B1(n5967), 
        .B2(EBX_REG_24__SCAN_IN), .ZN(n5412) );
  OAI21_X1 U6545 ( .B1(n5993), .B2(n5542), .A(n5412), .ZN(n5414) );
  NOR2_X1 U6546 ( .A1(n5753), .A2(n6542), .ZN(n5413) );
  AOI211_X1 U6547 ( .C1(n5961), .C2(n5415), .A(n5414), .B(n5413), .ZN(n5416)
         );
  OAI211_X1 U6548 ( .C1(n5471), .C2(n5946), .A(n5417), .B(n5416), .ZN(U2803)
         );
  INV_X1 U6549 ( .A(n5441), .ZN(n5743) );
  OAI21_X1 U6550 ( .B1(REIP_REG_22__SCAN_IN), .B2(REIP_REG_21__SCAN_IN), .A(
        n5743), .ZN(n5433) );
  INV_X1 U6551 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6540) );
  INV_X1 U6552 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6537) );
  NOR2_X1 U6553 ( .A1(n6540), .A2(n6537), .ZN(n5744) );
  AND2_X1 U6554 ( .A1(n2988), .A2(n5418), .ZN(n5420) );
  OR2_X1 U6555 ( .A1(n5420), .A2(n5419), .ZN(n5555) );
  INV_X1 U6556 ( .A(n5555), .ZN(n5421) );
  NAND2_X1 U6557 ( .A1(n5421), .A2(n5937), .ZN(n5432) );
  NAND2_X1 U6558 ( .A1(n5423), .A2(n5422), .ZN(n5762) );
  AOI22_X1 U6559 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n5987), .B1(n5558), 
        .B2(n5968), .ZN(n5424) );
  OAI21_X1 U6560 ( .B1(n6540), .B2(n5762), .A(n5424), .ZN(n5430) );
  NOR2_X1 U6561 ( .A1(n5426), .A2(n5425), .ZN(n5427) );
  OR2_X1 U6562 ( .A1(n5477), .A2(n5427), .ZN(n5637) );
  INV_X1 U6563 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5428) );
  OAI22_X1 U6564 ( .A1(n5637), .A2(n5982), .B1(n5428), .B2(n5981), .ZN(n5429)
         );
  NOR2_X1 U6565 ( .A1(n5430), .A2(n5429), .ZN(n5431) );
  OAI211_X1 U6566 ( .C1(n5433), .C2(n5744), .A(n5432), .B(n5431), .ZN(U2805)
         );
  NAND2_X1 U6567 ( .A1(n5435), .A2(n5434), .ZN(n5436) );
  INV_X1 U6568 ( .A(n5797), .ZN(n5445) );
  XNOR2_X1 U6569 ( .A(n5438), .B(n5437), .ZN(n5649) );
  INV_X1 U6570 ( .A(n5649), .ZN(n5443) );
  OAI22_X1 U6571 ( .A1(n5481), .A2(n5981), .B1(n5564), .B2(n5993), .ZN(n5439)
         );
  AOI21_X1 U6572 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n5987), .A(n5439), 
        .ZN(n5440) );
  OAI221_X1 U6573 ( .B1(REIP_REG_21__SCAN_IN), .B2(n5441), .C1(n6537), .C2(
        n5762), .A(n5440), .ZN(n5442) );
  AOI21_X1 U6574 ( .B1(n5443), .B2(n5961), .A(n5442), .ZN(n5444) );
  OAI21_X1 U6575 ( .B1(n5445), .B2(n5946), .A(n5444), .ZN(U2806) );
  NAND2_X1 U6576 ( .A1(n6002), .A2(n5937), .ZN(n5453) );
  NOR2_X1 U6577 ( .A1(n5942), .A2(n5446), .ZN(n5764) );
  OAI21_X1 U6578 ( .B1(REIP_REG_17__SCAN_IN), .B2(n5447), .A(n5764), .ZN(n5452) );
  AOI22_X1 U6579 ( .A1(EBX_REG_17__SCAN_IN), .A2(n5967), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n5987), .ZN(n5451) );
  NAND2_X1 U6580 ( .A1(n5968), .A2(n5822), .ZN(n5448) );
  OAI211_X1 U6581 ( .C1(n5842), .C2(n5982), .A(n3095), .B(n5448), .ZN(n5449)
         );
  INV_X1 U6582 ( .A(n5449), .ZN(n5450) );
  NAND4_X1 U6583 ( .A1(n5453), .A2(n5452), .A3(n5451), .A4(n5450), .ZN(U2810)
         );
  INV_X1 U6584 ( .A(n5454), .ZN(n5456) );
  OAI22_X1 U6585 ( .A1(n5456), .A2(n5773), .B1(n5455), .B2(n5997), .ZN(U2828)
         );
  INV_X1 U6586 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5457) );
  OAI222_X1 U6587 ( .A1(n5480), .A2(n5458), .B1(n5773), .B2(n5590), .C1(n5457), 
        .C2(n5997), .ZN(U2830) );
  OAI22_X1 U6588 ( .A1(n5600), .A2(n5773), .B1(n5459), .B2(n5997), .ZN(n5460)
         );
  AOI21_X1 U6589 ( .B1(n5783), .B2(n4286), .A(n5460), .ZN(n5461) );
  INV_X1 U6590 ( .A(n5461), .ZN(U2831) );
  INV_X1 U6591 ( .A(n5532), .ZN(n5496) );
  OAI222_X1 U6592 ( .A1(n5773), .A2(n5462), .B1(n5997), .B2(n6625), .C1(n5496), 
        .C2(n5480), .ZN(U2833) );
  AOI21_X1 U6593 ( .B1(n5464), .B2(n5406), .A(n2973), .ZN(n5809) );
  INV_X1 U6594 ( .A(n5809), .ZN(n5470) );
  INV_X1 U6595 ( .A(n5408), .ZN(n5468) );
  INV_X1 U6596 ( .A(n5465), .ZN(n5467) );
  OAI21_X1 U6597 ( .B1(n5468), .B2(n5467), .A(n5466), .ZN(n5738) );
  INV_X1 U6598 ( .A(n5738), .ZN(n5828) );
  AOI22_X1 U6599 ( .A1(n5828), .A2(n5995), .B1(n5490), .B2(EBX_REG_25__SCAN_IN), .ZN(n5469) );
  OAI21_X1 U6600 ( .B1(n5470), .B2(n5480), .A(n5469), .ZN(U2834) );
  INV_X1 U6601 ( .A(n5471), .ZN(n5791) );
  OAI22_X1 U6602 ( .A1(n5625), .A2(n5773), .B1(n6750), .B2(n5997), .ZN(n5472)
         );
  AOI21_X1 U6603 ( .B1(n5791), .B2(n4286), .A(n5472), .ZN(n5473) );
  INV_X1 U6604 ( .A(n5473), .ZN(U2835) );
  NOR2_X1 U6605 ( .A1(n5419), .A2(n5474), .ZN(n5475) );
  OR2_X1 U6606 ( .A1(n5405), .A2(n5475), .ZN(n5749) );
  INV_X1 U6607 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5479) );
  NOR2_X1 U6608 ( .A1(n5477), .A2(n5476), .ZN(n5478) );
  OR2_X1 U6609 ( .A1(n5409), .A2(n5478), .ZN(n5748) );
  OAI222_X1 U6610 ( .A1(n5480), .A2(n5749), .B1(n5997), .B2(n5479), .C1(n5748), 
        .C2(n5773), .ZN(U2836) );
  OAI222_X1 U6611 ( .A1(n5480), .A2(n5555), .B1(n5997), .B2(n5428), .C1(n5637), 
        .C2(n5773), .ZN(U2837) );
  OAI22_X1 U6612 ( .A1(n5649), .A2(n5773), .B1(n5481), .B2(n5997), .ZN(n5482)
         );
  AOI21_X1 U6613 ( .B1(n5797), .B2(n4286), .A(n5482), .ZN(n5483) );
  INV_X1 U6614 ( .A(n5483), .ZN(U2838) );
  AND2_X1 U6615 ( .A1(n5486), .A2(n5485), .ZN(n5487) );
  NOR2_X1 U6616 ( .A1(n5484), .A2(n5487), .ZN(n5813) );
  INV_X1 U6617 ( .A(n5813), .ZN(n5493) );
  XNOR2_X1 U6618 ( .A(n5489), .B(n5488), .ZN(n5767) );
  INV_X1 U6619 ( .A(n5767), .ZN(n5491) );
  AOI22_X1 U6620 ( .A1(n5491), .A2(n5995), .B1(n5490), .B2(EBX_REG_19__SCAN_IN), .ZN(n5492) );
  OAI21_X1 U6621 ( .B1(n5493), .B2(n5480), .A(n5492), .ZN(U2840) );
  AOI22_X1 U6622 ( .A1(n6005), .A2(DATAI_26_), .B1(n6008), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U6623 ( .A1(n6009), .A2(DATAI_10_), .ZN(n5494) );
  OAI211_X1 U6624 ( .C1(n5496), .C2(n5499), .A(n5495), .B(n5494), .ZN(U2865)
         );
  AOI22_X1 U6625 ( .A1(n6005), .A2(DATAI_22_), .B1(n6008), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U6626 ( .A1(n6009), .A2(DATAI_6_), .ZN(n5497) );
  OAI211_X1 U6627 ( .C1(n5555), .C2(n5499), .A(n5498), .B(n5497), .ZN(U2869)
         );
  INV_X1 U6628 ( .A(n5506), .ZN(n5516) );
  XNOR2_X1 U6629 ( .A(n5501), .B(n5586), .ZN(n5594) );
  NAND2_X1 U6630 ( .A1(n2971), .A2(REIP_REG_29__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U6631 ( .A1(n6142), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5502)
         );
  OAI211_X1 U6632 ( .C1(n6139), .C2(n5503), .A(n5588), .B(n5502), .ZN(n5504)
         );
  AOI21_X1 U6633 ( .B1(n5780), .B2(n6133), .A(n5504), .ZN(n5505) );
  OAI21_X1 U6634 ( .B1(n5594), .B2(n6137), .A(n5505), .ZN(U2957) );
  INV_X1 U6635 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U6636 ( .A1(n5607), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5509) );
  INV_X1 U6637 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5596) );
  NAND3_X1 U6638 ( .A1(n5516), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5596), .ZN(n5508) );
  OAI211_X1 U6639 ( .C1(n5507), .C2(n5509), .A(n5508), .B(n4289), .ZN(n5510)
         );
  AOI21_X1 U6640 ( .B1(n5587), .B2(n5506), .A(n5510), .ZN(n5603) );
  NAND2_X1 U6641 ( .A1(n5821), .A2(n5511), .ZN(n5512) );
  NAND2_X1 U6642 ( .A1(n2971), .A2(REIP_REG_28__SCAN_IN), .ZN(n5598) );
  OAI211_X1 U6643 ( .C1(n5824), .C2(n5513), .A(n5512), .B(n5598), .ZN(n5514)
         );
  AOI21_X1 U6644 ( .B1(n5783), .B2(n6133), .A(n5514), .ZN(n5515) );
  OAI21_X1 U6645 ( .B1(n5603), .B2(n6137), .A(n5515), .ZN(U2958) );
  NOR2_X1 U6646 ( .A1(n5516), .A2(n5507), .ZN(n5517) );
  XNOR2_X1 U6647 ( .A(n5517), .B(n5607), .ZN(n5614) );
  AND2_X1 U6648 ( .A1(n5395), .A2(n5518), .ZN(n5519) );
  NAND2_X1 U6649 ( .A1(n2971), .A2(REIP_REG_27__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U6650 ( .A1(n6142), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5520)
         );
  OAI211_X1 U6651 ( .C1(n6139), .C2(n5725), .A(n5609), .B(n5520), .ZN(n5521)
         );
  AOI21_X1 U6652 ( .B1(n5786), .B2(n6133), .A(n5521), .ZN(n5522) );
  OAI21_X1 U6653 ( .B1(n5614), .B2(n6137), .A(n5522), .ZN(U2959) );
  INV_X1 U6654 ( .A(n5523), .ZN(n5527) );
  NOR2_X1 U6655 ( .A1(n5525), .A2(n5524), .ZN(n5526) );
  XNOR2_X1 U6656 ( .A(n5527), .B(n5526), .ZN(n5622) );
  NAND2_X1 U6657 ( .A1(n5821), .A2(n5528), .ZN(n5529) );
  NAND2_X1 U6658 ( .A1(n2971), .A2(REIP_REG_26__SCAN_IN), .ZN(n5616) );
  OAI211_X1 U6659 ( .C1(n5824), .C2(n5530), .A(n5529), .B(n5616), .ZN(n5531)
         );
  AOI21_X1 U6660 ( .B1(n5532), .B2(n6133), .A(n5531), .ZN(n5533) );
  OAI21_X1 U6661 ( .B1(n5622), .B2(n6137), .A(n5533), .ZN(U2960) );
  OAI21_X1 U6662 ( .B1(n5534), .B2(n5679), .A(n5539), .ZN(n5535) );
  XNOR2_X1 U6663 ( .A(n5539), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5568)
         );
  INV_X1 U6664 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5536) );
  OR2_X1 U6665 ( .A1(n5539), .A2(n5536), .ZN(n5537) );
  INV_X1 U6666 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5639) );
  XNOR2_X1 U6667 ( .A(n5539), .B(n5639), .ZN(n5562) );
  INV_X1 U6668 ( .A(n5560), .ZN(n5538) );
  OAI21_X1 U6669 ( .B1(n2986), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5538), 
        .ZN(n5553) );
  NAND3_X1 U6670 ( .A1(n5539), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5540) );
  NOR2_X1 U6671 ( .A1(n5539), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5551)
         );
  NAND2_X1 U6672 ( .A1(n2971), .A2(REIP_REG_24__SCAN_IN), .ZN(n5624) );
  NAND2_X1 U6673 ( .A1(n6142), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5541)
         );
  OAI211_X1 U6674 ( .C1(n6139), .C2(n5542), .A(n5624), .B(n5541), .ZN(n5543)
         );
  AOI21_X1 U6675 ( .B1(n5791), .B2(n6133), .A(n5543), .ZN(n5544) );
  OAI21_X1 U6676 ( .B1(n5629), .B2(n6137), .A(n5544), .ZN(U2962) );
  OAI21_X1 U6677 ( .B1(n5567), .B2(n5546), .A(n5545), .ZN(n5547) );
  XNOR2_X1 U6678 ( .A(n5547), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5636)
         );
  INV_X1 U6679 ( .A(n5749), .ZN(n5794) );
  NAND2_X1 U6680 ( .A1(n2971), .A2(REIP_REG_23__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U6681 ( .A1(n6142), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5548)
         );
  OAI211_X1 U6682 ( .C1(n6139), .C2(n5745), .A(n5630), .B(n5548), .ZN(n5549)
         );
  AOI21_X1 U6683 ( .B1(n5794), .B2(n6133), .A(n5549), .ZN(n5550) );
  OAI21_X1 U6684 ( .B1(n5636), .B2(n6137), .A(n5550), .ZN(U2963) );
  AOI21_X1 U6685 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5539), .A(n5551), 
        .ZN(n5552) );
  XNOR2_X1 U6686 ( .A(n5553), .B(n5552), .ZN(n5647) );
  NAND2_X1 U6687 ( .A1(n2971), .A2(REIP_REG_22__SCAN_IN), .ZN(n5638) );
  OAI21_X1 U6688 ( .B1(n5824), .B2(n5554), .A(n5638), .ZN(n5557) );
  NOR2_X1 U6689 ( .A1(n5555), .A2(n6145), .ZN(n5556) );
  AOI211_X1 U6690 ( .C1(n5821), .C2(n5558), .A(n5557), .B(n5556), .ZN(n5559)
         );
  OAI21_X1 U6691 ( .B1(n5647), .B2(n6137), .A(n5559), .ZN(U2964) );
  AOI21_X1 U6692 ( .B1(n5562), .B2(n5561), .A(n5560), .ZN(n5654) );
  NAND2_X1 U6693 ( .A1(n2971), .A2(REIP_REG_21__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U6694 ( .A1(n6142), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5563)
         );
  OAI211_X1 U6695 ( .C1(n6139), .C2(n5564), .A(n5648), .B(n5563), .ZN(n5565)
         );
  AOI21_X1 U6696 ( .B1(n5797), .B2(n6133), .A(n5565), .ZN(n5566) );
  OAI21_X1 U6697 ( .B1(n5654), .B2(n6137), .A(n5566), .ZN(U2965) );
  OAI21_X1 U6698 ( .B1(n3093), .B2(n5568), .A(n5567), .ZN(n5669) );
  XOR2_X1 U6699 ( .A(n5569), .B(n5484), .Z(n5800) );
  INV_X1 U6700 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5756) );
  NAND2_X1 U6701 ( .A1(n5821), .A2(n5758), .ZN(n5570) );
  NAND2_X1 U6702 ( .A1(n2971), .A2(REIP_REG_20__SCAN_IN), .ZN(n5665) );
  OAI211_X1 U6703 ( .C1(n5824), .C2(n5756), .A(n5570), .B(n5665), .ZN(n5571)
         );
  AOI21_X1 U6704 ( .B1(n5800), .B2(n6133), .A(n5571), .ZN(n5572) );
  OAI21_X1 U6705 ( .B1(n5669), .B2(n6137), .A(n5572), .ZN(U2966) );
  NOR2_X1 U6706 ( .A1(n2986), .A2(n5857), .ZN(n5819) );
  NAND2_X1 U6707 ( .A1(n5819), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5575) );
  NOR2_X1 U6708 ( .A1(n5539), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5818)
         );
  NAND3_X1 U6709 ( .A1(n5573), .A2(n5818), .A3(n5834), .ZN(n5574) );
  OAI21_X1 U6710 ( .B1(n5573), .B2(n5575), .A(n5574), .ZN(n5576) );
  XNOR2_X1 U6711 ( .A(n5576), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5836)
         );
  INV_X1 U6712 ( .A(n5891), .ZN(n5578) );
  AOI22_X1 U6713 ( .A1(n6142), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .B1(n2971), 
        .B2(REIP_REG_18__SCAN_IN), .ZN(n5577) );
  OAI21_X1 U6714 ( .B1(n5578), .B2(n6139), .A(n5577), .ZN(n5579) );
  AOI21_X1 U6715 ( .B1(n5999), .B2(n6133), .A(n5579), .ZN(n5580) );
  OAI21_X1 U6716 ( .B1(n5836), .B2(n6137), .A(n5580), .ZN(U2968) );
  NOR2_X1 U6717 ( .A1(n5819), .A2(n5818), .ZN(n5581) );
  XNOR2_X1 U6718 ( .A(n5573), .B(n5581), .ZN(n5852) );
  INV_X1 U6719 ( .A(n5900), .ZN(n5583) );
  AOI22_X1 U6720 ( .A1(n6142), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n2971), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5582) );
  OAI21_X1 U6721 ( .B1(n5583), .B2(n6139), .A(n5582), .ZN(n5584) );
  AOI21_X1 U6722 ( .B1(n6007), .B2(n6133), .A(n5584), .ZN(n5585) );
  OAI21_X1 U6723 ( .B1(n5852), .B2(n6137), .A(n5585), .ZN(U2970) );
  NAND3_X1 U6724 ( .A1(n5608), .A2(n5587), .A3(n5586), .ZN(n5589) );
  OAI211_X1 U6725 ( .C1(n5590), .C2(n6213), .A(n5589), .B(n5588), .ZN(n5591)
         );
  AOI21_X1 U6726 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5592), .A(n5591), 
        .ZN(n5593) );
  OAI21_X1 U6727 ( .B1(n5594), .B2(n6198), .A(n5593), .ZN(U2989) );
  INV_X1 U6728 ( .A(n5595), .ZN(n5612) );
  XNOR2_X1 U6729 ( .A(n5596), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5597)
         );
  NAND2_X1 U6730 ( .A1(n5608), .A2(n5597), .ZN(n5599) );
  OAI211_X1 U6731 ( .C1(n6213), .C2(n5600), .A(n5599), .B(n5598), .ZN(n5601)
         );
  AOI21_X1 U6732 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n5612), .A(n5601), 
        .ZN(n5602) );
  OAI21_X1 U6733 ( .B1(n5603), .B2(n6198), .A(n5602), .ZN(U2990) );
  NOR2_X1 U6734 ( .A1(n5605), .A2(n5604), .ZN(n5606) );
  NAND2_X1 U6735 ( .A1(n5608), .A2(n5607), .ZN(n5610) );
  OAI211_X1 U6736 ( .C1(n6213), .C2(n5774), .A(n5610), .B(n5609), .ZN(n5611)
         );
  AOI21_X1 U6737 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5612), .A(n5611), 
        .ZN(n5613) );
  OAI21_X1 U6738 ( .B1(n5614), .B2(n6198), .A(n5613), .ZN(U2991) );
  OAI21_X1 U6739 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5827), .ZN(n5618) );
  NAND2_X1 U6740 ( .A1(n5615), .A2(n4302), .ZN(n5617) );
  OAI211_X1 U6741 ( .C1(n5619), .C2(n5618), .A(n5617), .B(n5616), .ZN(n5620)
         );
  AOI21_X1 U6742 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n5826), .A(n5620), 
        .ZN(n5621) );
  OAI21_X1 U6743 ( .B1(n5622), .B2(n6198), .A(n5621), .ZN(U2992) );
  OAI21_X1 U6744 ( .B1(n5631), .B2(n5623), .A(n6633), .ZN(n5627) );
  OAI21_X1 U6745 ( .B1(n5625), .B2(n6213), .A(n5624), .ZN(n5626) );
  AOI21_X1 U6746 ( .B1(n5826), .B2(n5627), .A(n5626), .ZN(n5628) );
  OAI21_X1 U6747 ( .B1(n5629), .B2(n6198), .A(n5628), .ZN(U2994) );
  OAI21_X1 U6748 ( .B1(n5748), .B2(n6213), .A(n5630), .ZN(n5633) );
  NOR2_X1 U6749 ( .A1(n5631), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5632)
         );
  AOI211_X1 U6750 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5634), .A(n5633), .B(n5632), .ZN(n5635) );
  OAI21_X1 U6751 ( .B1(n5636), .B2(n6198), .A(n5635), .ZN(U2995) );
  INV_X1 U6752 ( .A(n5637), .ZN(n5642) );
  INV_X1 U6753 ( .A(n5638), .ZN(n5641) );
  NOR3_X1 U6754 ( .A1(n5644), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n5639), 
        .ZN(n5640) );
  AOI211_X1 U6755 ( .C1(n4302), .C2(n5642), .A(n5641), .B(n5640), .ZN(n5646)
         );
  INV_X1 U6756 ( .A(n5643), .ZN(n5652) );
  NOR2_X1 U6757 ( .A1(n5644), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5650)
         );
  OAI21_X1 U6758 ( .B1(n5652), .B2(n5650), .A(INSTADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n5645) );
  OAI211_X1 U6759 ( .C1(n5647), .C2(n6198), .A(n5646), .B(n5645), .ZN(U2996)
         );
  OAI21_X1 U6760 ( .B1(n5649), .B2(n6213), .A(n5648), .ZN(n5651) );
  AOI211_X1 U6761 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5652), .A(n5651), .B(n5650), .ZN(n5653) );
  OAI21_X1 U6762 ( .B1(n5654), .B2(n6198), .A(n5653), .ZN(U2997) );
  AOI221_X1 U6763 ( .B1(n5656), .B2(n5834), .C1(n5655), .C2(n5834), .A(n5845), 
        .ZN(n5840) );
  OAI21_X1 U6764 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5686), .A(n5840), 
        .ZN(n5670) );
  MUX2_X1 U6765 ( .A(n5659), .B(n5658), .S(n5657), .Z(n5661) );
  XNOR2_X1 U6766 ( .A(n5661), .B(n5660), .ZN(n5759) );
  NOR2_X1 U6767 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5662) );
  NOR2_X1 U6768 ( .A1(n5663), .A2(n5662), .ZN(n5664) );
  NAND2_X1 U6769 ( .A1(n5676), .A2(n5664), .ZN(n5666) );
  OAI211_X1 U6770 ( .C1(n6213), .C2(n5759), .A(n5666), .B(n5665), .ZN(n5667)
         );
  AOI21_X1 U6771 ( .B1(n5670), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5667), 
        .ZN(n5668) );
  OAI21_X1 U6772 ( .B1(n5669), .B2(n6198), .A(n5668), .ZN(U2998) );
  INV_X1 U6773 ( .A(n5670), .ZN(n5680) );
  OAI21_X1 U6774 ( .B1(n5671), .B2(n5679), .A(n5672), .ZN(n5673) );
  XNOR2_X1 U6775 ( .A(n5673), .B(n2986), .ZN(n5814) );
  NAND2_X1 U6776 ( .A1(n5814), .A2(n6218), .ZN(n5678) );
  INV_X1 U6777 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5674) );
  OAI22_X1 U6778 ( .A1(n5767), .A2(n6213), .B1(n3095), .B2(n5674), .ZN(n5675)
         );
  AOI21_X1 U6779 ( .B1(n5676), .B2(n5679), .A(n5675), .ZN(n5677) );
  OAI211_X1 U6780 ( .C1(n5680), .C2(n5679), .A(n5678), .B(n5677), .ZN(U2999)
         );
  INV_X1 U6781 ( .A(n5681), .ZN(n5682) );
  AOI22_X1 U6782 ( .A1(n5684), .A2(n5683), .B1(n6209), .B2(n5682), .ZN(n6222)
         );
  OAI21_X1 U6783 ( .B1(n5686), .B2(n5685), .A(n6222), .ZN(n6183) );
  OAI21_X1 U6784 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n5687), .A(n6183), 
        .ZN(n5697) );
  NAND3_X1 U6785 ( .A1(n5689), .A2(n6217), .A3(n5688), .ZN(n5696) );
  AOI22_X1 U6786 ( .A1(n4302), .A2(n5690), .B1(n2971), .B2(REIP_REG_5__SCAN_IN), .ZN(n5695) );
  OAI21_X1 U6787 ( .B1(n5693), .B2(n5692), .A(n5691), .ZN(n6114) );
  OR2_X1 U6788 ( .A1(n6114), .A2(n6198), .ZN(n5694) );
  NAND4_X1 U6789 ( .A1(n5697), .A2(n5696), .A3(n5695), .A4(n5694), .ZN(U3013)
         );
  INV_X1 U6790 ( .A(n5698), .ZN(n5706) );
  OAI22_X1 U6791 ( .A1(n6213), .A2(n5699), .B1(n6593), .B2(n3095), .ZN(n5700)
         );
  AOI21_X1 U6792 ( .B1(n6218), .B2(n5701), .A(n5700), .ZN(n5705) );
  OAI21_X1 U6793 ( .B1(n5703), .B2(n5702), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5704) );
  NAND3_X1 U6794 ( .A1(n5706), .A2(n5705), .A3(n5704), .ZN(U3018) );
  OAI211_X1 U6795 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n5707), .A(n5710), .B(
        n6312), .ZN(n5708) );
  OAI21_X1 U6796 ( .B1(n5711), .B2(n5715), .A(n5708), .ZN(n5709) );
  MUX2_X1 U6797 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5709), .S(n6223), 
        .Z(U3464) );
  XNOR2_X1 U6798 ( .A(n5710), .B(n4429), .ZN(n5712) );
  OAI22_X1 U6799 ( .A1(n5712), .A2(n6364), .B1(n4426), .B2(n5711), .ZN(n5713)
         );
  MUX2_X1 U6800 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5713), .S(n6223), 
        .Z(U3463) );
  NOR3_X1 U6801 ( .A1(n6431), .A2(n5714), .A3(n4538), .ZN(n5717) );
  NOR2_X1 U6802 ( .A1(n5715), .A2(n6430), .ZN(n5716) );
  AOI211_X1 U6803 ( .C1(n6434), .C2(n3754), .A(n5717), .B(n5716), .ZN(n6437)
         );
  INV_X1 U6804 ( .A(n5718), .ZN(n6580) );
  AOI22_X1 U6805 ( .A1(n5721), .A2(n6580), .B1(n5720), .B2(n5719), .ZN(n5722)
         );
  OAI21_X1 U6806 ( .B1(n6437), .B2(n6586), .A(n5722), .ZN(n5723) );
  MUX2_X1 U6807 ( .A(n5723), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(n6583), 
        .Z(U3460) );
  AND2_X1 U6808 ( .A1(n6032), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  NOR2_X1 U6809 ( .A1(n5724), .A2(REIP_REG_27__SCAN_IN), .ZN(n5730) );
  INV_X1 U6810 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5728) );
  INV_X1 U6811 ( .A(n5725), .ZN(n5726) );
  AOI22_X1 U6812 ( .A1(n5968), .A2(n5726), .B1(n5967), .B2(EBX_REG_27__SCAN_IN), .ZN(n5727) );
  OAI21_X1 U6813 ( .B1(n5963), .B2(n5728), .A(n5727), .ZN(n5729) );
  AOI211_X1 U6814 ( .C1(n5786), .C2(n5937), .A(n5730), .B(n5729), .ZN(n5733)
         );
  INV_X1 U6815 ( .A(n5774), .ZN(n5731) );
  NAND2_X1 U6816 ( .A1(n5731), .A2(n5961), .ZN(n5732) );
  OAI211_X1 U6817 ( .C1(n5734), .C2(n6547), .A(n5733), .B(n5732), .ZN(U2800)
         );
  INV_X1 U6818 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6545) );
  OAI22_X1 U6819 ( .A1(n5993), .A2(n5812), .B1(n5735), .B2(n5981), .ZN(n5736)
         );
  AOI21_X1 U6820 ( .B1(PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n5987), .A(n5736), 
        .ZN(n5737) );
  OAI21_X1 U6821 ( .B1(n5738), .B2(n5982), .A(n5737), .ZN(n5739) );
  AOI21_X1 U6822 ( .B1(n5809), .B2(n5937), .A(n5739), .ZN(n5740) );
  OAI221_X1 U6823 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5742), .C1(n6545), .C2(
        n5741), .A(n5740), .ZN(U2802) );
  AOI21_X1 U6824 ( .B1(n5744), .B2(n5743), .A(REIP_REG_23__SCAN_IN), .ZN(n5754) );
  INV_X1 U6825 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5746) );
  OAI22_X1 U6826 ( .A1(n5746), .A2(n5963), .B1(n5745), .B2(n5993), .ZN(n5747)
         );
  AOI21_X1 U6827 ( .B1(EBX_REG_23__SCAN_IN), .B2(n5967), .A(n5747), .ZN(n5752)
         );
  OAI22_X1 U6828 ( .A1(n5749), .A2(n5946), .B1(n5748), .B2(n5982), .ZN(n5750)
         );
  INV_X1 U6829 ( .A(n5750), .ZN(n5751) );
  OAI211_X1 U6830 ( .C1(n5754), .C2(n5753), .A(n5752), .B(n5751), .ZN(U2804)
         );
  NOR2_X1 U6831 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5755), .ZN(n5763) );
  INV_X1 U6832 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5779) );
  OAI22_X1 U6833 ( .A1(n5779), .A2(n5981), .B1(n5756), .B2(n5963), .ZN(n5757)
         );
  AOI21_X1 U6834 ( .B1(n5758), .B2(n5968), .A(n5757), .ZN(n5761) );
  INV_X1 U6835 ( .A(n5759), .ZN(n5777) );
  AOI22_X1 U6836 ( .A1(n5800), .A2(n5937), .B1(n5961), .B2(n5777), .ZN(n5760)
         );
  OAI211_X1 U6837 ( .C1(n5763), .C2(n5762), .A(n5761), .B(n5760), .ZN(U2807)
         );
  INV_X1 U6838 ( .A(n5764), .ZN(n5893) );
  OAI22_X1 U6839 ( .A1(n5817), .A2(n5993), .B1(n5674), .B2(n5893), .ZN(n5765)
         );
  AOI211_X1 U6840 ( .C1(n5987), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n2971), 
        .B(n5765), .ZN(n5771) );
  OAI21_X1 U6841 ( .B1(REIP_REG_19__SCAN_IN), .B2(REIP_REG_18__SCAN_IN), .A(
        n5766), .ZN(n5768) );
  OAI22_X1 U6842 ( .A1(n5898), .A2(n5768), .B1(n5982), .B2(n5767), .ZN(n5769)
         );
  AOI21_X1 U6843 ( .B1(n5813), .B2(n5937), .A(n5769), .ZN(n5770) );
  OAI211_X1 U6844 ( .C1(n5772), .C2(n5981), .A(n5771), .B(n5770), .ZN(U2808)
         );
  NOR2_X1 U6845 ( .A1(n5774), .A2(n5773), .ZN(n5775) );
  AOI21_X1 U6846 ( .B1(n5786), .B2(n4286), .A(n5775), .ZN(n5776) );
  OAI21_X1 U6847 ( .B1(n6690), .B2(n5997), .A(n5776), .ZN(U2832) );
  AOI22_X1 U6848 ( .A1(n5800), .A2(n4286), .B1(n5995), .B2(n5777), .ZN(n5778)
         );
  OAI21_X1 U6849 ( .B1(n5779), .B2(n5997), .A(n5778), .ZN(U2839) );
  AOI22_X1 U6850 ( .A1(n5780), .A2(n6006), .B1(n6005), .B2(DATAI_29_), .ZN(
        n5782) );
  AOI22_X1 U6851 ( .A1(n6009), .A2(DATAI_13_), .B1(n6008), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5781) );
  NAND2_X1 U6852 ( .A1(n5782), .A2(n5781), .ZN(U2862) );
  AOI22_X1 U6853 ( .A1(n5783), .A2(n6006), .B1(n6005), .B2(DATAI_28_), .ZN(
        n5785) );
  AOI22_X1 U6854 ( .A1(n6009), .A2(DATAI_12_), .B1(n6008), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5784) );
  NAND2_X1 U6855 ( .A1(n5785), .A2(n5784), .ZN(U2863) );
  AOI22_X1 U6856 ( .A1(n5786), .A2(n6006), .B1(n6005), .B2(DATAI_27_), .ZN(
        n5788) );
  AOI22_X1 U6857 ( .A1(n6009), .A2(DATAI_11_), .B1(n6008), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5787) );
  NAND2_X1 U6858 ( .A1(n5788), .A2(n5787), .ZN(U2864) );
  AOI22_X1 U6859 ( .A1(n5809), .A2(n6006), .B1(n6005), .B2(DATAI_25_), .ZN(
        n5790) );
  AOI22_X1 U6860 ( .A1(n6009), .A2(DATAI_9_), .B1(n6008), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U6861 ( .A1(n5790), .A2(n5789), .ZN(U2866) );
  AOI22_X1 U6862 ( .A1(n5791), .A2(n6006), .B1(n6005), .B2(DATAI_24_), .ZN(
        n5793) );
  AOI22_X1 U6863 ( .A1(n6009), .A2(DATAI_8_), .B1(n6008), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U6864 ( .A1(n5793), .A2(n5792), .ZN(U2867) );
  AOI22_X1 U6865 ( .A1(n5794), .A2(n6006), .B1(n6005), .B2(DATAI_23_), .ZN(
        n5796) );
  AOI22_X1 U6866 ( .A1(n6009), .A2(DATAI_7_), .B1(n6008), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U6867 ( .A1(n5796), .A2(n5795), .ZN(U2868) );
  AOI22_X1 U6868 ( .A1(n5797), .A2(n6006), .B1(n6005), .B2(DATAI_21_), .ZN(
        n5799) );
  AOI22_X1 U6869 ( .A1(n6009), .A2(DATAI_5_), .B1(n6008), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U6870 ( .A1(n5799), .A2(n5798), .ZN(U2870) );
  AOI22_X1 U6871 ( .A1(n5800), .A2(n6006), .B1(n6005), .B2(DATAI_20_), .ZN(
        n5802) );
  AOI22_X1 U6872 ( .A1(n6009), .A2(DATAI_4_), .B1(n6008), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U6873 ( .A1(n5802), .A2(n5801), .ZN(U2871) );
  AOI22_X1 U6874 ( .A1(n5813), .A2(n6006), .B1(n6005), .B2(DATAI_19_), .ZN(
        n5804) );
  AOI22_X1 U6875 ( .A1(n6009), .A2(DATAI_3_), .B1(n6008), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5803) );
  NAND2_X1 U6876 ( .A1(n5804), .A2(n5803), .ZN(U2872) );
  AOI22_X1 U6877 ( .A1(n2971), .A2(REIP_REG_25__SCAN_IN), .B1(n6142), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5811) );
  INV_X1 U6878 ( .A(n5805), .ZN(n5806) );
  OAI21_X1 U6879 ( .B1(n5808), .B2(n5807), .A(n5806), .ZN(n5829) );
  AOI22_X1 U6880 ( .A1(n5809), .A2(n6133), .B1(n4310), .B2(n5829), .ZN(n5810)
         );
  OAI211_X1 U6881 ( .C1(n6139), .C2(n5812), .A(n5811), .B(n5810), .ZN(U2961)
         );
  AOI22_X1 U6882 ( .A1(n2971), .A2(REIP_REG_19__SCAN_IN), .B1(n6142), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5816) );
  AOI22_X1 U6883 ( .A1(n5814), .A2(n4310), .B1(n6133), .B2(n5813), .ZN(n5815)
         );
  OAI211_X1 U6884 ( .C1(n6139), .C2(n5817), .A(n5816), .B(n5815), .ZN(U2967)
         );
  INV_X1 U6885 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5825) );
  MUX2_X1 U6886 ( .A(n5819), .B(n5818), .S(n5573), .Z(n5820) );
  XNOR2_X1 U6887 ( .A(n5820), .B(n5834), .ZN(n5841) );
  AOI222_X1 U6888 ( .A1(n5841), .A2(n4310), .B1(n6133), .B2(n6002), .C1(n5822), 
        .C2(n5821), .ZN(n5823) );
  NAND2_X1 U6889 ( .A1(n2971), .A2(REIP_REG_17__SCAN_IN), .ZN(n5846) );
  OAI211_X1 U6890 ( .C1(n5825), .C2(n5824), .A(n5823), .B(n5846), .ZN(U2969)
         );
  INV_X1 U6891 ( .A(n5826), .ZN(n5832) );
  AOI22_X1 U6892 ( .A1(REIP_REG_25__SCAN_IN), .A2(n2971), .B1(n5827), .B2(
        n6674), .ZN(n5831) );
  AOI22_X1 U6893 ( .A1(n5829), .A2(n6218), .B1(n4302), .B2(n5828), .ZN(n5830)
         );
  OAI211_X1 U6894 ( .C1(n5832), .C2(n6674), .A(n5831), .B(n5830), .ZN(U2993)
         );
  INV_X1 U6895 ( .A(n5833), .ZN(n5848) );
  NOR3_X1 U6896 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5834), .A3(n5848), 
        .ZN(n5835) );
  AOI21_X1 U6897 ( .B1(REIP_REG_18__SCAN_IN), .B2(n2971), .A(n5835), .ZN(n5839) );
  INV_X1 U6898 ( .A(n5836), .ZN(n5837) );
  AOI22_X1 U6899 ( .A1(n5837), .A2(n6218), .B1(n4302), .B2(n5895), .ZN(n5838)
         );
  OAI211_X1 U6900 ( .C1(n5840), .C2(n6737), .A(n5839), .B(n5838), .ZN(U3000)
         );
  INV_X1 U6901 ( .A(n5841), .ZN(n5843) );
  OAI22_X1 U6902 ( .A1(n5843), .A2(n6198), .B1(n6213), .B2(n5842), .ZN(n5844)
         );
  AOI21_X1 U6903 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5845), .A(n5844), 
        .ZN(n5847) );
  OAI211_X1 U6904 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5848), .A(n5847), .B(n5846), .ZN(U3001) );
  AOI22_X1 U6905 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .B1(n5857), .B2(n5849), .ZN(n5850)
         );
  AOI22_X1 U6906 ( .A1(n2971), .A2(REIP_REG_16__SCAN_IN), .B1(n5851), .B2(
        n5850), .ZN(n5856) );
  INV_X1 U6907 ( .A(n5852), .ZN(n5854) );
  INV_X1 U6908 ( .A(n5853), .ZN(n5903) );
  AOI22_X1 U6909 ( .A1(n5854), .A2(n6218), .B1(n4302), .B2(n5903), .ZN(n5855)
         );
  OAI211_X1 U6910 ( .C1(n5858), .C2(n5857), .A(n5856), .B(n5855), .ZN(U3002)
         );
  OR2_X1 U6911 ( .A1(n5859), .A2(n6151), .ZN(n5867) );
  INV_X1 U6912 ( .A(n5860), .ZN(n5862) );
  AOI21_X1 U6913 ( .B1(n5862), .B2(n4302), .A(n5861), .ZN(n5866) );
  AOI22_X1 U6914 ( .A1(n5864), .A2(n6218), .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n5863), .ZN(n5865) );
  OAI211_X1 U6915 ( .C1(INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n5867), .A(n5866), .B(n5865), .ZN(U3004) );
  INV_X1 U6916 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6501) );
  INV_X1 U6917 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6695) );
  AOI21_X1 U6918 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6501), .A(n6695), .ZN(n5872) );
  INV_X1 U6919 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5868) );
  NOR2_X1 U6920 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6708), .ZN(n6611) );
  AOI21_X1 U6921 ( .B1(n5872), .B2(n5868), .A(n6611), .ZN(U2789) );
  OAI21_X1 U6922 ( .B1(n5869), .B2(n6474), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5870) );
  OAI21_X1 U6923 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6475), .A(n5870), .ZN(
        U2790) );
  NOR2_X1 U6924 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5873) );
  OAI21_X1 U6925 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5873), .A(n6597), .ZN(n5871)
         );
  OAI21_X1 U6926 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6597), .A(n5871), .ZN(
        U2791) );
  NOR2_X1 U6927 ( .A1(n6611), .A2(n5872), .ZN(n6564) );
  OAI21_X1 U6928 ( .B1(BS16_N), .B2(n5873), .A(n6564), .ZN(n6562) );
  OAI21_X1 U6929 ( .B1(n6564), .B2(n6602), .A(n6562), .ZN(U2792) );
  OAI21_X1 U6930 ( .B1(n5875), .B2(n5874), .A(n6137), .ZN(U2793) );
  NOR4_X1 U6931 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n5879) );
  NOR4_X1 U6932 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n5878) );
  NOR4_X1 U6933 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5877) );
  NOR4_X1 U6934 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5876) );
  NAND4_X1 U6935 ( .A1(n5879), .A2(n5878), .A3(n5877), .A4(n5876), .ZN(n5885)
         );
  NOR4_X1 U6936 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(n5883) );
  AOI211_X1 U6937 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_18__SCAN_IN), .B(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n5882) );
  NOR4_X1 U6938 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(n5881)
         );
  NOR4_X1 U6939 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n5880) );
  NAND4_X1 U6940 ( .A1(n5883), .A2(n5882), .A3(n5881), .A4(n5880), .ZN(n5884)
         );
  NOR2_X1 U6941 ( .A1(n5885), .A2(n5884), .ZN(n6591) );
  INV_X1 U6942 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5887) );
  NOR3_X1 U6943 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), 
        .A3(DATAWIDTH_REG_1__SCAN_IN), .ZN(n5888) );
  OAI21_X1 U6944 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5888), .A(n6591), .ZN(n5886)
         );
  OAI21_X1 U6945 ( .B1(n6591), .B2(n5887), .A(n5886), .ZN(U2794) );
  INV_X1 U6946 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6563) );
  AOI21_X1 U6947 ( .B1(n6587), .B2(n6563), .A(n5888), .ZN(n5890) );
  INV_X1 U6948 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5889) );
  INV_X1 U6949 ( .A(n6591), .ZN(n6594) );
  AOI22_X1 U6950 ( .A1(n6591), .A2(n5890), .B1(n5889), .B2(n6594), .ZN(U2795)
         );
  INV_X1 U6951 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6533) );
  AOI22_X1 U6952 ( .A1(EBX_REG_18__SCAN_IN), .A2(n5967), .B1(n5891), .B2(n5968), .ZN(n5892) );
  OAI21_X1 U6953 ( .B1(n6533), .B2(n5893), .A(n5892), .ZN(n5894) );
  AOI211_X1 U6954 ( .C1(n5987), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n2971), 
        .B(n5894), .ZN(n5897) );
  AOI22_X1 U6955 ( .A1(n5999), .A2(n5937), .B1(n5961), .B2(n5895), .ZN(n5896)
         );
  OAI211_X1 U6956 ( .C1(REIP_REG_18__SCAN_IN), .C2(n5898), .A(n5897), .B(n5896), .ZN(U2809) );
  OAI21_X1 U6957 ( .B1(REIP_REG_16__SCAN_IN), .B2(REIP_REG_15__SCAN_IN), .A(
        n5899), .ZN(n5906) );
  INV_X1 U6958 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6529) );
  AOI22_X1 U6959 ( .A1(EBX_REG_16__SCAN_IN), .A2(n5967), .B1(n5900), .B2(n5968), .ZN(n5901) );
  OAI21_X1 U6960 ( .B1(n6529), .B2(n5910), .A(n5901), .ZN(n5902) );
  AOI211_X1 U6961 ( .C1(n5987), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n2971), 
        .B(n5902), .ZN(n5905) );
  AOI22_X1 U6962 ( .A1(n6007), .A2(n5937), .B1(n5961), .B2(n5903), .ZN(n5904)
         );
  OAI211_X1 U6963 ( .C1(n5918), .C2(n5906), .A(n5905), .B(n5904), .ZN(U2811)
         );
  OAI21_X1 U6964 ( .B1(n5963), .B2(n5907), .A(n3095), .ZN(n5912) );
  INV_X1 U6965 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6527) );
  INV_X1 U6966 ( .A(n5908), .ZN(n5909) );
  OAI22_X1 U6967 ( .A1(n5910), .A2(n6527), .B1(n5982), .B2(n5909), .ZN(n5911)
         );
  AOI211_X1 U6968 ( .C1(EBX_REG_15__SCAN_IN), .C2(n5967), .A(n5912), .B(n5911), 
        .ZN(n5917) );
  INV_X1 U6969 ( .A(n5913), .ZN(n5915) );
  AOI22_X1 U6970 ( .A1(n5915), .A2(n5937), .B1(n5968), .B2(n5914), .ZN(n5916)
         );
  OAI211_X1 U6971 ( .C1(REIP_REG_15__SCAN_IN), .C2(n5918), .A(n5917), .B(n5916), .ZN(U2812) );
  AOI22_X1 U6972 ( .A1(n5920), .A2(n5937), .B1(n5919), .B2(n5968), .ZN(n5928)
         );
  INV_X1 U6973 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6521) );
  AOI22_X1 U6974 ( .A1(n5921), .A2(n5961), .B1(n5967), .B2(EBX_REG_12__SCAN_IN), .ZN(n5922) );
  OAI211_X1 U6975 ( .C1(n5963), .C2(n5923), .A(n5922), .B(n3095), .ZN(n5924)
         );
  AOI221_X1 U6976 ( .B1(n5926), .B2(REIP_REG_12__SCAN_IN), .C1(n5925), .C2(
        n6521), .A(n5924), .ZN(n5927) );
  NAND2_X1 U6977 ( .A1(n5928), .A2(n5927), .ZN(U2815) );
  XNOR2_X1 U6978 ( .A(n5930), .B(n5929), .ZN(n5994) );
  AOI21_X1 U6979 ( .B1(n5967), .B2(EBX_REG_7__SCAN_IN), .A(n2971), .ZN(n5931)
         );
  OAI21_X1 U6980 ( .B1(n5994), .B2(n5982), .A(n5931), .ZN(n5932) );
  AOI21_X1 U6981 ( .B1(n5987), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n5932), 
        .ZN(n5933) );
  OAI21_X1 U6982 ( .B1(n5934), .B2(REIP_REG_7__SCAN_IN), .A(n5933), .ZN(n5935)
         );
  INV_X1 U6983 ( .A(n5935), .ZN(n5940) );
  INV_X1 U6984 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6511) );
  NAND2_X1 U6985 ( .A1(n5936), .A2(n6511), .ZN(n5950) );
  OAI21_X1 U6986 ( .B1(n5941), .B2(n5942), .A(n5950), .ZN(n5938) );
  AOI22_X1 U6987 ( .A1(n5938), .A2(REIP_REG_7__SCAN_IN), .B1(n5937), .B2(n6110), .ZN(n5939) );
  OAI211_X1 U6988 ( .C1(n6113), .C2(n5993), .A(n5940), .B(n5939), .ZN(U2820)
         );
  OR2_X1 U6989 ( .A1(n5942), .A2(n5941), .ZN(n5952) );
  AOI21_X1 U6990 ( .B1(n5967), .B2(EBX_REG_6__SCAN_IN), .A(n2971), .ZN(n5943)
         );
  OAI21_X1 U6991 ( .B1(n6177), .B2(n5982), .A(n5943), .ZN(n5944) );
  AOI21_X1 U6992 ( .B1(n5987), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n5944), 
        .ZN(n5945) );
  OAI21_X1 U6993 ( .B1(n5947), .B2(n5946), .A(n5945), .ZN(n5948) );
  AOI21_X1 U6994 ( .B1(n5949), .B2(n5968), .A(n5948), .ZN(n5951) );
  OAI211_X1 U6995 ( .C1(n5952), .C2(n6511), .A(n5951), .B(n5950), .ZN(U2821)
         );
  NAND2_X1 U6996 ( .A1(n5987), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5956)
         );
  AOI21_X1 U6997 ( .B1(n5953), .B2(n6509), .A(n5952), .ZN(n5954) );
  AOI211_X1 U6998 ( .C1(n5967), .C2(EBX_REG_5__SCAN_IN), .A(n2971), .B(n5954), 
        .ZN(n5955) );
  OAI211_X1 U6999 ( .C1(n5957), .C2(n5982), .A(n5956), .B(n5955), .ZN(n5958)
         );
  AOI21_X1 U7000 ( .B1(n6115), .B2(n5986), .A(n5958), .ZN(n5959) );
  OAI21_X1 U7001 ( .B1(n6119), .B2(n5993), .A(n5959), .ZN(U2822) );
  INV_X1 U7002 ( .A(n5960), .ZN(n6191) );
  AOI22_X1 U7003 ( .A1(n5962), .A2(n5984), .B1(n5961), .B2(n6191), .ZN(n5976)
         );
  INV_X1 U7004 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6507) );
  OAI22_X1 U7005 ( .A1(n5965), .A2(n6507), .B1(n5964), .B2(n5963), .ZN(n5966)
         );
  AOI211_X1 U7006 ( .C1(n5967), .C2(EBX_REG_4__SCAN_IN), .A(n2971), .B(n5966), 
        .ZN(n5975) );
  AOI22_X1 U7007 ( .A1(n5970), .A2(n5986), .B1(n5969), .B2(n5968), .ZN(n5974)
         );
  NAND3_X1 U7008 ( .A1(n5972), .A2(n5971), .A3(n6507), .ZN(n5973) );
  NAND4_X1 U7009 ( .A1(n5976), .A2(n5975), .A3(n5974), .A4(n5973), .ZN(U2823)
         );
  OAI21_X1 U7010 ( .B1(n5977), .B2(n6587), .A(n6503), .ZN(n5978) );
  NAND2_X1 U7011 ( .A1(n5979), .A2(n5978), .ZN(n5991) );
  INV_X1 U7012 ( .A(n4426), .ZN(n5985) );
  OAI22_X1 U7013 ( .A1(n6212), .A2(n5982), .B1(n5981), .B2(n5980), .ZN(n5983)
         );
  AOI21_X1 U7014 ( .B1(n5985), .B2(n5984), .A(n5983), .ZN(n5990) );
  NAND2_X1 U7015 ( .A1(n5986), .A2(n6132), .ZN(n5989) );
  NAND2_X1 U7016 ( .A1(n5987), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5988)
         );
  AND4_X1 U7017 ( .A1(n5991), .A2(n5990), .A3(n5989), .A4(n5988), .ZN(n5992)
         );
  OAI21_X1 U7018 ( .B1(n6136), .B2(n5993), .A(n5992), .ZN(U2825) );
  INV_X1 U7019 ( .A(n5994), .ZN(n6170) );
  AOI22_X1 U7020 ( .A1(n6110), .A2(n4286), .B1(n5995), .B2(n6170), .ZN(n5996)
         );
  OAI21_X1 U7021 ( .B1(n5998), .B2(n5997), .A(n5996), .ZN(U2852) );
  AOI22_X1 U7022 ( .A1(n5999), .A2(n6006), .B1(n6005), .B2(DATAI_18_), .ZN(
        n6001) );
  AOI22_X1 U7023 ( .A1(n6009), .A2(DATAI_2_), .B1(n6008), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7024 ( .A1(n6001), .A2(n6000), .ZN(U2873) );
  AOI22_X1 U7025 ( .A1(n6002), .A2(n6006), .B1(n6005), .B2(DATAI_17_), .ZN(
        n6004) );
  AOI22_X1 U7026 ( .A1(n6009), .A2(DATAI_1_), .B1(n6008), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7027 ( .A1(n6004), .A2(n6003), .ZN(U2874) );
  AOI22_X1 U7028 ( .A1(n6007), .A2(n6006), .B1(n6005), .B2(DATAI_16_), .ZN(
        n6011) );
  AOI22_X1 U7029 ( .A1(n6009), .A2(DATAI_0_), .B1(n6008), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7030 ( .A1(n6011), .A2(n6010), .ZN(U2875) );
  INV_X1 U7031 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n6680) );
  INV_X1 U7032 ( .A(n6012), .ZN(n6013) );
  AOI22_X1 U7033 ( .A1(n6032), .A2(DATAO_REG_20__SCAN_IN), .B1(n6013), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6014) );
  OAI21_X1 U7034 ( .B1(n6600), .B2(n6680), .A(n6014), .ZN(U2903) );
  INV_X1 U7035 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6105) );
  AOI22_X1 U7036 ( .A1(n6030), .A2(LWORD_REG_15__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6015) );
  OAI21_X1 U7037 ( .B1(n6105), .B2(n6038), .A(n6015), .ZN(U2908) );
  INV_X1 U7038 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6100) );
  AOI22_X1 U7039 ( .A1(n6030), .A2(LWORD_REG_14__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6016) );
  OAI21_X1 U7040 ( .B1(n6100), .B2(n6038), .A(n6016), .ZN(U2909) );
  AOI22_X1 U7041 ( .A1(n6030), .A2(LWORD_REG_13__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6017) );
  OAI21_X1 U7042 ( .B1(n6018), .B2(n6038), .A(n6017), .ZN(U2910) );
  AOI22_X1 U7043 ( .A1(n6030), .A2(LWORD_REG_12__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6019) );
  OAI21_X1 U7044 ( .B1(n5074), .B2(n6038), .A(n6019), .ZN(U2911) );
  INV_X1 U7045 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6091) );
  AOI22_X1 U7046 ( .A1(n6030), .A2(LWORD_REG_11__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6020) );
  OAI21_X1 U7047 ( .B1(n6091), .B2(n6038), .A(n6020), .ZN(U2912) );
  INV_X1 U7048 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6087) );
  AOI22_X1 U7049 ( .A1(n6030), .A2(LWORD_REG_10__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6021) );
  OAI21_X1 U7050 ( .B1(n6087), .B2(n6038), .A(n6021), .ZN(U2913) );
  AOI22_X1 U7051 ( .A1(n6030), .A2(LWORD_REG_9__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6022) );
  OAI21_X1 U7052 ( .B1(n6023), .B2(n6038), .A(n6022), .ZN(U2914) );
  INV_X1 U7053 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6083) );
  AOI22_X1 U7054 ( .A1(n6030), .A2(LWORD_REG_8__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6024) );
  OAI21_X1 U7055 ( .B1(n6083), .B2(n6038), .A(n6024), .ZN(U2915) );
  INV_X1 U7056 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6026) );
  AOI22_X1 U7057 ( .A1(n6030), .A2(LWORD_REG_7__SCAN_IN), .B1(
        DATAO_REG_7__SCAN_IN), .B2(n6032), .ZN(n6025) );
  OAI21_X1 U7058 ( .B1(n6026), .B2(n6038), .A(n6025), .ZN(U2916) );
  AOI22_X1 U7059 ( .A1(n6030), .A2(LWORD_REG_6__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6027) );
  OAI21_X1 U7060 ( .B1(n6028), .B2(n6038), .A(n6027), .ZN(U2917) );
  AOI22_X1 U7061 ( .A1(n6030), .A2(LWORD_REG_5__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6029) );
  OAI21_X1 U7062 ( .B1(n4987), .B2(n6038), .A(n6029), .ZN(U2918) );
  AOI22_X1 U7063 ( .A1(n6030), .A2(LWORD_REG_4__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6031) );
  OAI21_X1 U7064 ( .B1(n6616), .B2(n6038), .A(n6031), .ZN(U2919) );
  INV_X1 U7065 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n6620) );
  AOI22_X1 U7066 ( .A1(EAX_REG_3__SCAN_IN), .A2(n6040), .B1(n6032), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6033) );
  OAI21_X1 U7067 ( .B1(n6600), .B2(n6620), .A(n6033), .ZN(U2920) );
  AOI22_X1 U7068 ( .A1(n6036), .A2(LWORD_REG_2__SCAN_IN), .B1(n6032), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6034) );
  OAI21_X1 U7069 ( .B1(n6035), .B2(n6038), .A(n6034), .ZN(U2921) );
  AOI22_X1 U7070 ( .A1(n6036), .A2(LWORD_REG_1__SCAN_IN), .B1(
        DATAO_REG_1__SCAN_IN), .B2(n6032), .ZN(n6037) );
  OAI21_X1 U7071 ( .B1(n6039), .B2(n6038), .A(n6037), .ZN(U2922) );
  INV_X1 U7072 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n6671) );
  AOI22_X1 U7073 ( .A1(EAX_REG_0__SCAN_IN), .A2(n6040), .B1(
        DATAO_REG_0__SCAN_IN), .B2(n6032), .ZN(n6041) );
  OAI21_X1 U7074 ( .B1(n6600), .B2(n6671), .A(n6041), .ZN(U2923) );
  OAI21_X1 U7075 ( .B1(n2984), .B2(n6491), .A(n6042), .ZN(n6089) );
  AOI22_X1 U7076 ( .A1(n6101), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n6094), .ZN(n6044) );
  OAI21_X1 U7077 ( .B1(n6097), .B2(n6067), .A(n6044), .ZN(U2924) );
  AOI22_X1 U7078 ( .A1(n6089), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n6094), .ZN(n6045) );
  OAI21_X1 U7079 ( .B1(n6097), .B2(n6069), .A(n6045), .ZN(U2925) );
  AOI22_X1 U7080 ( .A1(n6089), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6094), .ZN(n6046) );
  OAI21_X1 U7081 ( .B1(n6097), .B2(n6071), .A(n6046), .ZN(U2926) );
  AOI22_X1 U7082 ( .A1(n6089), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6094), .ZN(n6047) );
  OAI21_X1 U7083 ( .B1(n6097), .B2(n6073), .A(n6047), .ZN(U2927) );
  AOI22_X1 U7084 ( .A1(n6089), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6094), .ZN(n6048) );
  OAI21_X1 U7085 ( .B1(n6097), .B2(n6075), .A(n6048), .ZN(U2928) );
  AOI22_X1 U7086 ( .A1(n6101), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6094), .ZN(n6049) );
  OAI21_X1 U7087 ( .B1(n6097), .B2(n4986), .A(n6049), .ZN(U2929) );
  AOI22_X1 U7088 ( .A1(n6089), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6094), .ZN(n6050) );
  OAI21_X1 U7089 ( .B1(n6097), .B2(n6078), .A(n6050), .ZN(U2930) );
  AOI22_X1 U7090 ( .A1(n6101), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6094), .ZN(n6051) );
  OAI21_X1 U7091 ( .B1(n6097), .B2(n6080), .A(n6051), .ZN(U2931) );
  INV_X1 U7092 ( .A(DATAI_8_), .ZN(n6052) );
  NOR2_X1 U7093 ( .A1(n6097), .A2(n6052), .ZN(n6081) );
  AOI21_X1 U7094 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6101), .A(n6081), .ZN(n6053) );
  OAI21_X1 U7095 ( .B1(n4117), .B2(n6104), .A(n6053), .ZN(U2932) );
  AOI22_X1 U7096 ( .A1(n6101), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n6094), .ZN(n6054) );
  OAI21_X1 U7097 ( .B1(n6097), .B2(n6740), .A(n6054), .ZN(U2933) );
  INV_X1 U7098 ( .A(DATAI_10_), .ZN(n6055) );
  NOR2_X1 U7099 ( .A1(n6097), .A2(n6055), .ZN(n6085) );
  AOI21_X1 U7100 ( .B1(UWORD_REG_10__SCAN_IN), .B2(n6101), .A(n6085), .ZN(
        n6056) );
  OAI21_X1 U7101 ( .B1(n6057), .B2(n6104), .A(n6056), .ZN(U2934) );
  INV_X1 U7102 ( .A(DATAI_11_), .ZN(n6058) );
  NOR2_X1 U7103 ( .A1(n6097), .A2(n6058), .ZN(n6088) );
  AOI21_X1 U7104 ( .B1(UWORD_REG_11__SCAN_IN), .B2(n6101), .A(n6088), .ZN(
        n6059) );
  OAI21_X1 U7105 ( .B1(n4178), .B2(n6104), .A(n6059), .ZN(U2935) );
  NOR2_X1 U7106 ( .A1(n6097), .A2(n6060), .ZN(n6092) );
  AOI21_X1 U7107 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6101), .A(n6092), .ZN(
        n6061) );
  OAI21_X1 U7108 ( .B1(n6062), .B2(n6104), .A(n6061), .ZN(U2936) );
  AOI22_X1 U7109 ( .A1(n6101), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n6094), .ZN(n6063) );
  OAI21_X1 U7110 ( .B1(n6097), .B2(n6096), .A(n6063), .ZN(U2937) );
  INV_X1 U7111 ( .A(DATAI_14_), .ZN(n6064) );
  NOR2_X1 U7112 ( .A1(n6097), .A2(n6064), .ZN(n6098) );
  AOI21_X1 U7113 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6101), .A(n6098), .ZN(
        n6065) );
  OAI21_X1 U7114 ( .B1(n4253), .B2(n6104), .A(n6065), .ZN(U2938) );
  AOI22_X1 U7115 ( .A1(n6101), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6094), .ZN(n6066) );
  OAI21_X1 U7116 ( .B1(n6097), .B2(n6067), .A(n6066), .ZN(U2939) );
  AOI22_X1 U7117 ( .A1(n6101), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6094), .ZN(n6068) );
  OAI21_X1 U7118 ( .B1(n6097), .B2(n6069), .A(n6068), .ZN(U2940) );
  AOI22_X1 U7119 ( .A1(n6101), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6094), .ZN(n6070) );
  OAI21_X1 U7120 ( .B1(n6097), .B2(n6071), .A(n6070), .ZN(U2941) );
  AOI22_X1 U7121 ( .A1(n6101), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6094), .ZN(n6072) );
  OAI21_X1 U7122 ( .B1(n6097), .B2(n6073), .A(n6072), .ZN(U2942) );
  AOI22_X1 U7123 ( .A1(n6101), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6094), .ZN(n6074) );
  OAI21_X1 U7124 ( .B1(n6097), .B2(n6075), .A(n6074), .ZN(U2943) );
  AOI22_X1 U7125 ( .A1(n6101), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6094), .ZN(n6076) );
  OAI21_X1 U7126 ( .B1(n6097), .B2(n4986), .A(n6076), .ZN(U2944) );
  AOI22_X1 U7127 ( .A1(n6101), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6094), .ZN(n6077) );
  OAI21_X1 U7128 ( .B1(n6097), .B2(n6078), .A(n6077), .ZN(U2945) );
  AOI22_X1 U7129 ( .A1(n6101), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6094), .ZN(n6079) );
  OAI21_X1 U7130 ( .B1(n6097), .B2(n6080), .A(n6079), .ZN(U2946) );
  AOI21_X1 U7131 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6101), .A(n6081), .ZN(n6082) );
  OAI21_X1 U7132 ( .B1(n6083), .B2(n6104), .A(n6082), .ZN(U2947) );
  AOI22_X1 U7133 ( .A1(n6101), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n6094), .ZN(n6084) );
  OAI21_X1 U7134 ( .B1(n6097), .B2(n6740), .A(n6084), .ZN(U2948) );
  AOI21_X1 U7135 ( .B1(LWORD_REG_10__SCAN_IN), .B2(n6101), .A(n6085), .ZN(
        n6086) );
  OAI21_X1 U7136 ( .B1(n6087), .B2(n6104), .A(n6086), .ZN(U2949) );
  AOI21_X1 U7137 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6089), .A(n6088), .ZN(
        n6090) );
  OAI21_X1 U7138 ( .B1(n6091), .B2(n6104), .A(n6090), .ZN(U2950) );
  AOI21_X1 U7139 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6101), .A(n6092), .ZN(
        n6093) );
  OAI21_X1 U7140 ( .B1(n5074), .B2(n6104), .A(n6093), .ZN(U2951) );
  AOI22_X1 U7141 ( .A1(n6101), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n6094), .ZN(n6095) );
  OAI21_X1 U7142 ( .B1(n6097), .B2(n6096), .A(n6095), .ZN(U2952) );
  AOI21_X1 U7143 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6101), .A(n6098), .ZN(
        n6099) );
  OAI21_X1 U7144 ( .B1(n6100), .B2(n6104), .A(n6099), .ZN(U2953) );
  AOI22_X1 U7145 ( .A1(n6102), .A2(DATAI_15_), .B1(n6101), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n6103) );
  OAI21_X1 U7146 ( .B1(n6105), .B2(n6104), .A(n6103), .ZN(U2954) );
  AOI22_X1 U7147 ( .A1(n2971), .A2(REIP_REG_7__SCAN_IN), .B1(n6142), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6112) );
  OAI21_X1 U7148 ( .B1(n6108), .B2(n6107), .A(n6106), .ZN(n6109) );
  INV_X1 U7149 ( .A(n6109), .ZN(n6171) );
  AOI22_X1 U7150 ( .A1(n6171), .A2(n4310), .B1(n6133), .B2(n6110), .ZN(n6111)
         );
  OAI211_X1 U7151 ( .C1(n6139), .C2(n6113), .A(n6112), .B(n6111), .ZN(U2979)
         );
  AOI22_X1 U7152 ( .A1(n2971), .A2(REIP_REG_5__SCAN_IN), .B1(n6142), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6118) );
  INV_X1 U7153 ( .A(n6114), .ZN(n6116) );
  AOI22_X1 U7154 ( .A1(n6116), .A2(n4310), .B1(n6133), .B2(n6115), .ZN(n6117)
         );
  OAI211_X1 U7155 ( .C1(n6139), .C2(n6119), .A(n6118), .B(n6117), .ZN(U2981)
         );
  AOI22_X1 U7156 ( .A1(n2971), .A2(REIP_REG_3__SCAN_IN), .B1(n6142), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6127) );
  OAI21_X1 U7157 ( .B1(n6122), .B2(n6121), .A(n6120), .ZN(n6199) );
  INV_X1 U7158 ( .A(n6199), .ZN(n6125) );
  INV_X1 U7159 ( .A(n6123), .ZN(n6124) );
  AOI22_X1 U7160 ( .A1(n4310), .A2(n6125), .B1(n6124), .B2(n6133), .ZN(n6126)
         );
  OAI211_X1 U7161 ( .C1(n6139), .C2(n6128), .A(n6127), .B(n6126), .ZN(U2983)
         );
  AOI22_X1 U7162 ( .A1(n2971), .A2(REIP_REG_2__SCAN_IN), .B1(n6142), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6135) );
  XOR2_X1 U7163 ( .A(n6129), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n6130) );
  XNOR2_X1 U7164 ( .A(n6131), .B(n6130), .ZN(n6219) );
  AOI22_X1 U7165 ( .A1(n6219), .A2(n4310), .B1(n6133), .B2(n6132), .ZN(n6134)
         );
  OAI211_X1 U7166 ( .C1(n6139), .C2(n6136), .A(n6135), .B(n6134), .ZN(U2984)
         );
  OAI22_X1 U7167 ( .A1(n6139), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6138), 
        .B2(n6137), .ZN(n6140) );
  AOI211_X1 U7168 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6142), .A(n6141), 
        .B(n6140), .ZN(n6143) );
  OAI21_X1 U7169 ( .B1(n6145), .B2(n6144), .A(n6143), .ZN(U2985) );
  INV_X1 U7170 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6519) );
  OAI222_X1 U7171 ( .A1(n6147), .A2(n6213), .B1(n3095), .B2(n6519), .C1(n6198), 
        .C2(n6146), .ZN(n6148) );
  INV_X1 U7172 ( .A(n6148), .ZN(n6149) );
  OAI221_X1 U7173 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6151), .C1(
        n3517), .C2(n6150), .A(n6149), .ZN(U3007) );
  AOI21_X1 U7174 ( .B1(n4302), .B2(n6153), .A(n6152), .ZN(n6157) );
  AOI22_X1 U7175 ( .A1(n6155), .A2(n6218), .B1(n6154), .B2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6156) );
  OAI211_X1 U7176 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6158), .A(n6157), 
        .B(n6156), .ZN(U3009) );
  INV_X1 U7177 ( .A(n6159), .ZN(n6162) );
  INV_X1 U7178 ( .A(n6160), .ZN(n6161) );
  AOI21_X1 U7179 ( .B1(n4302), .B2(n6162), .A(n6161), .ZN(n6168) );
  INV_X1 U7180 ( .A(n6163), .ZN(n6166) );
  AOI21_X1 U7181 ( .B1(n6175), .B2(n6169), .A(n6164), .ZN(n6165) );
  AOI22_X1 U7182 ( .A1(n6166), .A2(n6218), .B1(n6172), .B2(n6165), .ZN(n6167)
         );
  OAI211_X1 U7183 ( .C1(n6176), .C2(n6169), .A(n6168), .B(n6167), .ZN(U3010)
         );
  AOI22_X1 U7184 ( .A1(n4302), .A2(n6170), .B1(n2971), .B2(REIP_REG_7__SCAN_IN), .ZN(n6174) );
  AOI22_X1 U7185 ( .A1(n6172), .A2(n6175), .B1(n6171), .B2(n6218), .ZN(n6173)
         );
  OAI211_X1 U7186 ( .C1(n6176), .C2(n6175), .A(n6174), .B(n6173), .ZN(U3011)
         );
  INV_X1 U7187 ( .A(n6177), .ZN(n6180) );
  INV_X1 U7188 ( .A(n6178), .ZN(n6179) );
  AOI21_X1 U7189 ( .B1(n4302), .B2(n6180), .A(n6179), .ZN(n6185) );
  INV_X1 U7190 ( .A(n6181), .ZN(n6182) );
  AOI22_X1 U7191 ( .A1(n6183), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .B1(n6218), 
        .B2(n6182), .ZN(n6184) );
  OAI211_X1 U7192 ( .C1(INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n6186), .A(n6185), 
        .B(n6184), .ZN(U3012) );
  NAND2_X1 U7193 ( .A1(n6187), .A2(n6206), .ZN(n6204) );
  OAI21_X1 U7194 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6188), .ZN(n6196) );
  INV_X1 U7195 ( .A(n6189), .ZN(n6190) );
  AOI21_X1 U7196 ( .B1(n4302), .B2(n6191), .A(n6190), .ZN(n6195) );
  OAI21_X1 U7197 ( .B1(n6206), .B2(n6209), .A(n6222), .ZN(n6201) );
  INV_X1 U7198 ( .A(n6192), .ZN(n6193) );
  AOI22_X1 U7199 ( .A1(n6201), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .B1(n6218), 
        .B2(n6193), .ZN(n6194) );
  OAI211_X1 U7200 ( .C1(n6204), .C2(n6196), .A(n6195), .B(n6194), .ZN(U3014)
         );
  AOI22_X1 U7201 ( .A1(n4302), .A2(n6197), .B1(n2971), .B2(REIP_REG_3__SCAN_IN), .ZN(n6203) );
  NOR2_X1 U7202 ( .A1(n6199), .A2(n6198), .ZN(n6200) );
  AOI21_X1 U7203 ( .B1(n6201), .B2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6200), 
        .ZN(n6202) );
  OAI211_X1 U7204 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n6204), .A(n6203), 
        .B(n6202), .ZN(U3015) );
  INV_X1 U7205 ( .A(n6206), .ZN(n6207) );
  AOI21_X1 U7206 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n3351), .A(n6207), 
        .ZN(n6208) );
  OR2_X1 U7207 ( .A1(n6209), .A2(n6208), .ZN(n6211) );
  NAND2_X1 U7208 ( .A1(n2971), .A2(REIP_REG_2__SCAN_IN), .ZN(n6210) );
  OAI211_X1 U7209 ( .C1(n6213), .C2(n6212), .A(n6211), .B(n6210), .ZN(n6214)
         );
  INV_X1 U7210 ( .A(n6214), .ZN(n6221) );
  NOR2_X1 U7211 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n6215), .ZN(n6216)
         );
  AOI22_X1 U7212 ( .A1(n6219), .A2(n6218), .B1(n6217), .B2(n6216), .ZN(n6220)
         );
  OAI211_X1 U7213 ( .C1(n6222), .C2(n6758), .A(n6221), .B(n6220), .ZN(U3016)
         );
  NOR2_X1 U7214 ( .A1(n6459), .A2(n6223), .ZN(U3019) );
  OR2_X1 U7215 ( .A1(n6225), .A2(n6224), .ZN(n6227) );
  NOR2_X1 U7216 ( .A1(n6356), .A2(n6231), .ZN(n6253) );
  INV_X1 U7217 ( .A(n6253), .ZN(n6226) );
  AND2_X1 U7218 ( .A1(n6227), .A2(n6226), .ZN(n6232) );
  AND2_X1 U7219 ( .A1(n6230), .A2(n6232), .ZN(n6228) );
  INV_X1 U7220 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n6706) );
  NOR2_X2 U7221 ( .A1(n6260), .A2(n6229), .ZN(n6296) );
  AOI22_X1 U7222 ( .A1(n6418), .A2(n6253), .B1(n6360), .B2(n6296), .ZN(n6236)
         );
  INV_X1 U7223 ( .A(n6230), .ZN(n6233) );
  OAI22_X1 U7224 ( .A1(n6233), .A2(n6232), .B1(n6601), .B2(n6231), .ZN(n6255)
         );
  AOI22_X1 U7225 ( .A1(n6255), .A2(n6421), .B1(n6368), .B2(n6254), .ZN(n6235)
         );
  OAI211_X1 U7226 ( .C1(n6259), .C2(n6706), .A(n6236), .B(n6235), .ZN(U3060)
         );
  INV_X1 U7227 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6749) );
  AOI22_X1 U7228 ( .A1(n6373), .A2(n6253), .B1(n6372), .B2(n6296), .ZN(n6238)
         );
  AOI22_X1 U7229 ( .A1(n6255), .A2(n6335), .B1(n6374), .B2(n6254), .ZN(n6237)
         );
  OAI211_X1 U7230 ( .C1(n6259), .C2(n6749), .A(n6238), .B(n6237), .ZN(U3061)
         );
  INV_X1 U7231 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6241) );
  AOI22_X1 U7232 ( .A1(n6379), .A2(n6253), .B1(n6378), .B2(n6296), .ZN(n6240)
         );
  AOI22_X1 U7233 ( .A1(n6255), .A2(n6339), .B1(n6380), .B2(n6254), .ZN(n6239)
         );
  OAI211_X1 U7234 ( .C1(n6259), .C2(n6241), .A(n6240), .B(n6239), .ZN(U3062)
         );
  INV_X1 U7235 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n6244) );
  AOI22_X1 U7236 ( .A1(n6385), .A2(n6253), .B1(n6386), .B2(n6296), .ZN(n6243)
         );
  AOI22_X1 U7237 ( .A1(n6255), .A2(n6279), .B1(n6384), .B2(n6254), .ZN(n6242)
         );
  OAI211_X1 U7238 ( .C1(n6259), .C2(n6244), .A(n6243), .B(n6242), .ZN(U3063)
         );
  INV_X1 U7239 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n6247) );
  AOI22_X1 U7240 ( .A1(n6391), .A2(n6253), .B1(n6392), .B2(n6296), .ZN(n6246)
         );
  AOI22_X1 U7241 ( .A1(n6255), .A2(n6343), .B1(n6390), .B2(n6254), .ZN(n6245)
         );
  OAI211_X1 U7242 ( .C1(n6259), .C2(n6247), .A(n6246), .B(n6245), .ZN(U3064)
         );
  INV_X1 U7243 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n6733) );
  AOI22_X1 U7244 ( .A1(n6397), .A2(n6253), .B1(n6396), .B2(n6296), .ZN(n6249)
         );
  AOI22_X1 U7245 ( .A1(n6255), .A2(n6286), .B1(n6398), .B2(n6254), .ZN(n6248)
         );
  OAI211_X1 U7246 ( .C1(n6259), .C2(n6733), .A(n6249), .B(n6248), .ZN(U3065)
         );
  INV_X1 U7247 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6252) );
  AOI22_X1 U7248 ( .A1(n6403), .A2(n6253), .B1(n6404), .B2(n6296), .ZN(n6251)
         );
  AOI22_X1 U7249 ( .A1(n6255), .A2(n6290), .B1(n6402), .B2(n6254), .ZN(n6250)
         );
  OAI211_X1 U7250 ( .C1(n6259), .C2(n6252), .A(n6251), .B(n6250), .ZN(U3066)
         );
  INV_X1 U7251 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n6258) );
  AOI22_X1 U7252 ( .A1(n2999), .A2(n6253), .B1(n6783), .B2(n6296), .ZN(n6257)
         );
  AOI22_X1 U7253 ( .A1(n6255), .A2(n6350), .B1(n6412), .B2(n6254), .ZN(n6256)
         );
  OAI211_X1 U7254 ( .C1(n6259), .C2(n6258), .A(n6257), .B(n6256), .ZN(U3067)
         );
  AOI22_X1 U7255 ( .A1(n6264), .A2(n6304), .B1(n6263), .B2(n6262), .ZN(n6265)
         );
  AND2_X1 U7256 ( .A1(n6356), .A2(n6313), .ZN(n6294) );
  AOI22_X1 U7257 ( .A1(n6421), .A2(n6295), .B1(n6418), .B2(n6294), .ZN(n6272)
         );
  NOR2_X1 U7258 ( .A1(n6303), .A2(n6364), .ZN(n6269) );
  OAI21_X1 U7259 ( .B1(n6330), .B2(n6296), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6268) );
  AOI211_X1 U7260 ( .C1(n6269), .C2(n6268), .A(n6267), .B(n6266), .ZN(n6270)
         );
  OAI211_X1 U7261 ( .C1(n6294), .C2(n6718), .A(n6270), .B(n6446), .ZN(n6297)
         );
  AOI22_X1 U7262 ( .A1(n6297), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6368), 
        .B2(n6296), .ZN(n6271) );
  OAI211_X1 U7263 ( .C1(n6422), .C2(n6300), .A(n6272), .B(n6271), .ZN(U3068)
         );
  AOI22_X1 U7264 ( .A1(n6373), .A2(n6294), .B1(n6335), .B2(n6295), .ZN(n6274)
         );
  AOI22_X1 U7265 ( .A1(n6297), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6374), 
        .B2(n6296), .ZN(n6273) );
  OAI211_X1 U7266 ( .C1(n6275), .C2(n6300), .A(n6274), .B(n6273), .ZN(U3069)
         );
  AOI22_X1 U7267 ( .A1(n6379), .A2(n6294), .B1(n6339), .B2(n6295), .ZN(n6277)
         );
  AOI22_X1 U7268 ( .A1(n6297), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6380), 
        .B2(n6296), .ZN(n6276) );
  OAI211_X1 U7269 ( .C1(n6278), .C2(n6300), .A(n6277), .B(n6276), .ZN(U3070)
         );
  AOI22_X1 U7270 ( .A1(n6385), .A2(n6294), .B1(n6279), .B2(n6295), .ZN(n6281)
         );
  AOI22_X1 U7271 ( .A1(n6297), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6384), 
        .B2(n6296), .ZN(n6280) );
  OAI211_X1 U7272 ( .C1(n6282), .C2(n6300), .A(n6281), .B(n6280), .ZN(U3071)
         );
  AOI22_X1 U7273 ( .A1(n6391), .A2(n6294), .B1(n6343), .B2(n6295), .ZN(n6284)
         );
  AOI22_X1 U7274 ( .A1(n6297), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6390), 
        .B2(n6296), .ZN(n6283) );
  OAI211_X1 U7275 ( .C1(n6285), .C2(n6300), .A(n6284), .B(n6283), .ZN(U3072)
         );
  AOI22_X1 U7276 ( .A1(n6286), .A2(n6295), .B1(n6397), .B2(n6294), .ZN(n6288)
         );
  AOI22_X1 U7277 ( .A1(n6297), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6398), 
        .B2(n6296), .ZN(n6287) );
  OAI211_X1 U7278 ( .C1(n6289), .C2(n6300), .A(n6288), .B(n6287), .ZN(U3073)
         );
  AOI22_X1 U7279 ( .A1(n6403), .A2(n6294), .B1(n6290), .B2(n6295), .ZN(n6292)
         );
  AOI22_X1 U7280 ( .A1(n6297), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6402), 
        .B2(n6296), .ZN(n6291) );
  OAI211_X1 U7281 ( .C1(n6293), .C2(n6300), .A(n6292), .B(n6291), .ZN(U3074)
         );
  AOI22_X1 U7282 ( .A1(n6350), .A2(n6295), .B1(n2999), .B2(n6294), .ZN(n6299)
         );
  AOI22_X1 U7283 ( .A1(n6297), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6412), 
        .B2(n6296), .ZN(n6298) );
  OAI211_X1 U7284 ( .C1(n6301), .C2(n6300), .A(n6299), .B(n6298), .ZN(U3075)
         );
  AND2_X1 U7285 ( .A1(n6302), .A2(n6312), .ZN(n6309) );
  NAND3_X1 U7286 ( .A1(n6304), .A2(n6303), .A3(n3763), .ZN(n6305) );
  NAND2_X1 U7287 ( .A1(n6305), .A2(n6306), .ZN(n6307) );
  AOI22_X1 U7288 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6313), .B1(n6309), .B2(
        n6307), .ZN(n6334) );
  INV_X1 U7289 ( .A(n6306), .ZN(n6329) );
  AOI22_X1 U7290 ( .A1(n6418), .A2(n6329), .B1(n6360), .B2(n6328), .ZN(n6315)
         );
  INV_X1 U7291 ( .A(n6307), .ZN(n6308) );
  NAND2_X1 U7292 ( .A1(n6309), .A2(n6308), .ZN(n6311) );
  OAI211_X1 U7293 ( .C1(n6313), .C2(n6312), .A(n6311), .B(n6310), .ZN(n6331)
         );
  AOI22_X1 U7294 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6331), .B1(n6368), 
        .B2(n6330), .ZN(n6314) );
  OAI211_X1 U7295 ( .C1(n6334), .C2(n6371), .A(n6315), .B(n6314), .ZN(U3076)
         );
  AOI22_X1 U7296 ( .A1(n6373), .A2(n6329), .B1(n6372), .B2(n6328), .ZN(n6317)
         );
  AOI22_X1 U7297 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6331), .B1(n6374), 
        .B2(n6330), .ZN(n6316) );
  OAI211_X1 U7298 ( .C1(n6334), .C2(n6377), .A(n6317), .B(n6316), .ZN(U3077)
         );
  AOI22_X1 U7299 ( .A1(n6379), .A2(n6329), .B1(n6380), .B2(n6330), .ZN(n6319)
         );
  AOI22_X1 U7300 ( .A1(n6331), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n6378), 
        .B2(n6328), .ZN(n6318) );
  OAI211_X1 U7301 ( .C1(n6334), .C2(n6383), .A(n6319), .B(n6318), .ZN(U3078)
         );
  AOI22_X1 U7302 ( .A1(n6385), .A2(n6329), .B1(n6384), .B2(n6330), .ZN(n6321)
         );
  AOI22_X1 U7303 ( .A1(n6331), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n6386), 
        .B2(n6328), .ZN(n6320) );
  OAI211_X1 U7304 ( .C1(n6334), .C2(n6389), .A(n6321), .B(n6320), .ZN(U3079)
         );
  AOI22_X1 U7305 ( .A1(n6391), .A2(n6329), .B1(n6390), .B2(n6330), .ZN(n6323)
         );
  AOI22_X1 U7306 ( .A1(n6331), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n6392), 
        .B2(n6328), .ZN(n6322) );
  OAI211_X1 U7307 ( .C1(n6334), .C2(n6395), .A(n6323), .B(n6322), .ZN(U3080)
         );
  AOI22_X1 U7308 ( .A1(n6397), .A2(n6329), .B1(n6396), .B2(n6328), .ZN(n6325)
         );
  AOI22_X1 U7309 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6331), .B1(n6398), 
        .B2(n6330), .ZN(n6324) );
  OAI211_X1 U7310 ( .C1(n6334), .C2(n6401), .A(n6325), .B(n6324), .ZN(U3081)
         );
  AOI22_X1 U7311 ( .A1(n6403), .A2(n6329), .B1(n6402), .B2(n6330), .ZN(n6327)
         );
  AOI22_X1 U7312 ( .A1(n6331), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n6404), 
        .B2(n6328), .ZN(n6326) );
  OAI211_X1 U7313 ( .C1(n6334), .C2(n6407), .A(n6327), .B(n6326), .ZN(U3082)
         );
  AOI22_X1 U7314 ( .A1(n2999), .A2(n6329), .B1(n6783), .B2(n6328), .ZN(n6333)
         );
  AOI22_X1 U7315 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6331), .B1(n6412), 
        .B2(n6330), .ZN(n6332) );
  OAI211_X1 U7316 ( .C1(n6334), .C2(n6786), .A(n6333), .B(n6332), .ZN(U3083)
         );
  AOI22_X1 U7317 ( .A1(n6373), .A2(n6348), .B1(n6347), .B2(n6372), .ZN(n6337)
         );
  AOI22_X1 U7318 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6351), .B1(n6335), 
        .B2(n6349), .ZN(n6336) );
  OAI211_X1 U7319 ( .C1(n6338), .C2(n6354), .A(n6337), .B(n6336), .ZN(U3109)
         );
  AOI22_X1 U7320 ( .A1(n6379), .A2(n6348), .B1(n6347), .B2(n6378), .ZN(n6341)
         );
  AOI22_X1 U7321 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6351), .B1(n6339), 
        .B2(n6349), .ZN(n6340) );
  OAI211_X1 U7322 ( .C1(n6342), .C2(n6354), .A(n6341), .B(n6340), .ZN(U3110)
         );
  AOI22_X1 U7323 ( .A1(n6391), .A2(n6348), .B1(n6347), .B2(n6392), .ZN(n6345)
         );
  AOI22_X1 U7324 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6351), .B1(n6343), 
        .B2(n6349), .ZN(n6344) );
  OAI211_X1 U7325 ( .C1(n6346), .C2(n6354), .A(n6345), .B(n6344), .ZN(U3112)
         );
  AOI22_X1 U7326 ( .A1(n2999), .A2(n6348), .B1(n6347), .B2(n6783), .ZN(n6353)
         );
  AOI22_X1 U7327 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6351), .B1(n6350), 
        .B2(n6349), .ZN(n6352) );
  OAI211_X1 U7328 ( .C1(n6778), .C2(n6354), .A(n6353), .B(n6352), .ZN(U3115)
         );
  OR2_X1 U7329 ( .A1(n6355), .A2(n6364), .ZN(n6367) );
  NOR2_X1 U7330 ( .A1(n6356), .A2(n6363), .ZN(n6409) );
  AOI21_X1 U7331 ( .B1(n6358), .B2(n6357), .A(n6409), .ZN(n6361) );
  OAI22_X1 U7332 ( .A1(n6601), .A2(n6363), .B1(n6367), .B2(n6361), .ZN(n6359)
         );
  AOI22_X1 U7333 ( .A1(n6418), .A2(n6409), .B1(n6360), .B2(n6408), .ZN(n6370)
         );
  INV_X1 U7334 ( .A(n6361), .ZN(n6366) );
  AOI21_X1 U7335 ( .B1(n6364), .B2(n6363), .A(n6362), .ZN(n6365) );
  OAI21_X1 U7336 ( .B1(n6367), .B2(n6366), .A(n6365), .ZN(n6413) );
  AOI22_X1 U7337 ( .A1(n6413), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n6368), 
        .B2(n6411), .ZN(n6369) );
  OAI211_X1 U7338 ( .C1(n6416), .C2(n6371), .A(n6370), .B(n6369), .ZN(U3124)
         );
  AOI22_X1 U7339 ( .A1(n6373), .A2(n6409), .B1(n6372), .B2(n6408), .ZN(n6376)
         );
  AOI22_X1 U7340 ( .A1(n6413), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n6374), 
        .B2(n6411), .ZN(n6375) );
  OAI211_X1 U7341 ( .C1(n6416), .C2(n6377), .A(n6376), .B(n6375), .ZN(U3125)
         );
  AOI22_X1 U7342 ( .A1(n6379), .A2(n6409), .B1(n6378), .B2(n6408), .ZN(n6382)
         );
  AOI22_X1 U7343 ( .A1(n6413), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n6380), 
        .B2(n6411), .ZN(n6381) );
  OAI211_X1 U7344 ( .C1(n6416), .C2(n6383), .A(n6382), .B(n6381), .ZN(U3126)
         );
  AOI22_X1 U7345 ( .A1(n6385), .A2(n6409), .B1(n6384), .B2(n6411), .ZN(n6388)
         );
  AOI22_X1 U7346 ( .A1(n6413), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n6386), 
        .B2(n6408), .ZN(n6387) );
  OAI211_X1 U7347 ( .C1(n6416), .C2(n6389), .A(n6388), .B(n6387), .ZN(U3127)
         );
  AOI22_X1 U7348 ( .A1(n6391), .A2(n6409), .B1(n6390), .B2(n6411), .ZN(n6394)
         );
  AOI22_X1 U7349 ( .A1(n6413), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n6392), 
        .B2(n6408), .ZN(n6393) );
  OAI211_X1 U7350 ( .C1(n6416), .C2(n6395), .A(n6394), .B(n6393), .ZN(U3128)
         );
  AOI22_X1 U7351 ( .A1(n6397), .A2(n6409), .B1(n6396), .B2(n6408), .ZN(n6400)
         );
  AOI22_X1 U7352 ( .A1(n6413), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n6398), 
        .B2(n6411), .ZN(n6399) );
  OAI211_X1 U7353 ( .C1(n6416), .C2(n6401), .A(n6400), .B(n6399), .ZN(U3129)
         );
  AOI22_X1 U7354 ( .A1(n6403), .A2(n6409), .B1(n6402), .B2(n6411), .ZN(n6406)
         );
  AOI22_X1 U7355 ( .A1(n6413), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n6404), 
        .B2(n6408), .ZN(n6405) );
  OAI211_X1 U7356 ( .C1(n6416), .C2(n6407), .A(n6406), .B(n6405), .ZN(U3130)
         );
  AOI22_X1 U7357 ( .A1(n2999), .A2(n6409), .B1(n6783), .B2(n6408), .ZN(n6415)
         );
  AOI22_X1 U7358 ( .A1(n6413), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n6412), 
        .B2(n6411), .ZN(n6414) );
  OAI211_X1 U7359 ( .C1(n6416), .C2(n6786), .A(n6415), .B(n6414), .ZN(U3131)
         );
  INV_X1 U7360 ( .A(n6417), .ZN(n6429) );
  INV_X1 U7361 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n6626) );
  AOI22_X1 U7362 ( .A1(n6421), .A2(n6420), .B1(n6419), .B2(n6418), .ZN(n6428)
         );
  OAI22_X1 U7363 ( .A1(n6425), .A2(n6424), .B1(n6423), .B2(n6422), .ZN(n6426)
         );
  INV_X1 U7364 ( .A(n6426), .ZN(n6427) );
  OAI211_X1 U7365 ( .C1(n6429), .C2(n6626), .A(n6428), .B(n6427), .ZN(U3140)
         );
  INV_X1 U7366 ( .A(n6430), .ZN(n6433) );
  NOR2_X1 U7367 ( .A1(n6431), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6432)
         );
  AOI21_X1 U7368 ( .B1(n3763), .B2(n6433), .A(n6432), .ZN(n6576) );
  NAND2_X1 U7369 ( .A1(n6434), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6585) );
  AND2_X1 U7370 ( .A1(n6585), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6435)
         );
  AND2_X1 U7371 ( .A1(n6576), .A2(n6435), .ZN(n6440) );
  AOI211_X1 U7372 ( .C1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n6440), .A(n6437), .B(n6436), .ZN(n6438) );
  INV_X1 U7373 ( .A(n6438), .ZN(n6439) );
  OAI21_X1 U7374 ( .B1(n6440), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6439), 
        .ZN(n6443) );
  INV_X1 U7375 ( .A(n6443), .ZN(n6445) );
  AOI21_X1 U7376 ( .B1(n6443), .B2(n6442), .A(n6441), .ZN(n6444) );
  AOI21_X1 U7377 ( .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6445), .A(n6444), 
        .ZN(n6448) );
  INV_X1 U7378 ( .A(n6448), .ZN(n6451) );
  INV_X1 U7379 ( .A(n6447), .ZN(n6450) );
  OAI21_X1 U7380 ( .B1(n6448), .B2(n6447), .A(n6446), .ZN(n6449) );
  OAI21_X1 U7381 ( .B1(n6451), .B2(n6450), .A(n6449), .ZN(n6460) );
  OAI21_X1 U7382 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6452), 
        .ZN(n6453) );
  NAND4_X1 U7383 ( .A1(n6456), .A2(n6455), .A3(n6454), .A4(n6453), .ZN(n6457)
         );
  AOI211_X1 U7384 ( .C1(n6460), .C2(n6459), .A(n6458), .B(n6457), .ZN(n6461)
         );
  INV_X1 U7385 ( .A(n6461), .ZN(n6466) );
  OAI22_X1 U7386 ( .A1(n6466), .A2(n6474), .B1(n6491), .B2(n6600), .ZN(n6462)
         );
  OAI21_X1 U7387 ( .B1(n6464), .B2(n6463), .A(n6462), .ZN(n6568) );
  OAI21_X1 U7388 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6491), .A(n6568), .ZN(
        n6477) );
  AOI211_X1 U7389 ( .C1(n6467), .C2(n6466), .A(n6465), .B(n6477), .ZN(n6472)
         );
  INV_X1 U7390 ( .A(n6468), .ZN(n6469) );
  OAI211_X1 U7391 ( .C1(n6469), .C2(n6471), .A(n6603), .B(n6568), .ZN(n6470)
         );
  OAI221_X1 U7392 ( .B1(n6603), .B2(n6472), .C1(n6603), .C2(n6471), .A(n6470), 
        .ZN(U3148) );
  INV_X1 U7393 ( .A(n6473), .ZN(n6480) );
  NOR2_X1 U7394 ( .A1(n6603), .A2(n6634), .ZN(n6481) );
  OAI21_X1 U7395 ( .B1(READY_N), .B2(n6475), .A(n6474), .ZN(n6476) );
  AOI22_X1 U7396 ( .A1(n6481), .A2(n6477), .B1(n6568), .B2(n6476), .ZN(n6479)
         );
  OAI211_X1 U7397 ( .C1(n6480), .C2(n6568), .A(n6479), .B(n6478), .ZN(U3149)
         );
  INV_X1 U7398 ( .A(n6566), .ZN(n6484) );
  AOI21_X1 U7399 ( .B1(n6481), .B2(n6491), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n6483) );
  OAI21_X1 U7400 ( .B1(n6484), .B2(n6483), .A(n6482), .ZN(U3150) );
  AND2_X1 U7401 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6560), .ZN(U3151) );
  AND2_X1 U7402 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6560), .ZN(U3152) );
  AND2_X1 U7403 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6560), .ZN(U3153) );
  AND2_X1 U7404 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6560), .ZN(U3154) );
  AND2_X1 U7405 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6560), .ZN(U3155) );
  AND2_X1 U7406 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6560), .ZN(U3156) );
  AND2_X1 U7407 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6560), .ZN(U3157) );
  AND2_X1 U7408 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6560), .ZN(U3158) );
  AND2_X1 U7409 ( .A1(n6560), .A2(DATAWIDTH_REG_23__SCAN_IN), .ZN(U3159) );
  AND2_X1 U7410 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6560), .ZN(U3160) );
  AND2_X1 U7411 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6560), .ZN(U3161) );
  AND2_X1 U7412 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6560), .ZN(U3162) );
  AND2_X1 U7413 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6560), .ZN(U3163) );
  AND2_X1 U7414 ( .A1(n6560), .A2(DATAWIDTH_REG_18__SCAN_IN), .ZN(U3164) );
  INV_X1 U7415 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6701) );
  NOR2_X1 U7416 ( .A1(n6564), .A2(n6701), .ZN(U3165) );
  AND2_X1 U7417 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6560), .ZN(U3166) );
  AND2_X1 U7418 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6560), .ZN(U3167) );
  AND2_X1 U7419 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6560), .ZN(U3168) );
  AND2_X1 U7420 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6560), .ZN(U3169) );
  AND2_X1 U7421 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6560), .ZN(U3170) );
  AND2_X1 U7422 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6560), .ZN(U3171) );
  AND2_X1 U7423 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6560), .ZN(U3172) );
  AND2_X1 U7424 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6560), .ZN(U3173) );
  AND2_X1 U7425 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6560), .ZN(U3174) );
  AND2_X1 U7426 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6560), .ZN(U3175) );
  AND2_X1 U7427 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6560), .ZN(U3176) );
  AND2_X1 U7428 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6560), .ZN(U3177) );
  AND2_X1 U7429 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6560), .ZN(U3178) );
  AND2_X1 U7430 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6560), .ZN(U3179) );
  AND2_X1 U7431 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6560), .ZN(U3180) );
  INV_X1 U7432 ( .A(n6499), .ZN(n6486) );
  AOI22_X1 U7433 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6500) );
  OAI221_X1 U7434 ( .B1(n6501), .B2(NA_N), .C1(n6501), .C2(n6708), .A(n6695), 
        .ZN(n6496) );
  AND2_X1 U7435 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6487) );
  INV_X1 U7436 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6609) );
  OAI21_X1 U7437 ( .B1(n6487), .B2(n6609), .A(n6597), .ZN(n6485) );
  OAI211_X1 U7438 ( .C1(n6486), .C2(n6500), .A(n6496), .B(n6485), .ZN(U3181)
         );
  NOR2_X1 U7439 ( .A1(n6695), .A2(n6609), .ZN(n6488) );
  NAND2_X1 U7440 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6493) );
  OAI21_X1 U7441 ( .B1(n6488), .B2(n6487), .A(n6493), .ZN(n6489) );
  OAI211_X1 U7442 ( .C1(n6708), .C2(n6491), .A(n6490), .B(n6489), .ZN(U3182)
         );
  NOR4_X1 U7443 ( .A1(NA_N), .A2(n6695), .A3(n6491), .A4(n6609), .ZN(n6497) );
  NOR2_X1 U7444 ( .A1(NA_N), .A2(n6491), .ZN(n6492) );
  OAI211_X1 U7445 ( .C1(n6492), .C2(n6708), .A(HOLD), .B(n6609), .ZN(n6494) );
  NAND3_X1 U7446 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6494), .A3(n6493), .ZN(
        n6495) );
  AOI22_X1 U7447 ( .A1(STATE_REG_1__SCAN_IN), .A2(n6497), .B1(n6496), .B2(
        n6495), .ZN(n6498) );
  OAI21_X1 U7448 ( .B1(n6500), .B2(n6499), .A(n6498), .ZN(U3183) );
  NAND2_X1 U7449 ( .A1(n6611), .A2(n6501), .ZN(n6517) );
  NOR2_X1 U7450 ( .A1(n6501), .A2(n6597), .ZN(n6548) );
  INV_X1 U7451 ( .A(n6548), .ZN(n6553) );
  AOI22_X1 U7452 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6555), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6597), .ZN(n6502) );
  OAI21_X1 U7453 ( .B1(n6503), .B2(n6517), .A(n6502), .ZN(U3184) );
  AOI22_X1 U7454 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6555), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6597), .ZN(n6504) );
  OAI21_X1 U7455 ( .B1(n6505), .B2(n6517), .A(n6504), .ZN(U3185) );
  AOI22_X1 U7456 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6555), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6597), .ZN(n6506) );
  OAI21_X1 U7457 ( .B1(n6507), .B2(n6517), .A(n6506), .ZN(U3186) );
  AOI22_X1 U7458 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6555), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6597), .ZN(n6508) );
  OAI21_X1 U7459 ( .B1(n6509), .B2(n6517), .A(n6508), .ZN(U3187) );
  AOI22_X1 U7460 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6555), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6597), .ZN(n6510) );
  OAI21_X1 U7461 ( .B1(n6511), .B2(n6517), .A(n6510), .ZN(U3188) );
  AOI22_X1 U7462 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6555), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6597), .ZN(n6512) );
  OAI21_X1 U7463 ( .B1(n6513), .B2(n6517), .A(n6512), .ZN(U3189) );
  INV_X1 U7464 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6725) );
  AOI22_X1 U7465 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6555), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6597), .ZN(n6514) );
  OAI21_X1 U7466 ( .B1(n6725), .B2(n6517), .A(n6514), .ZN(U3190) );
  AOI22_X1 U7467 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6555), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6597), .ZN(n6515) );
  OAI21_X1 U7468 ( .B1(n6721), .B2(n6517), .A(n6515), .ZN(U3191) );
  INV_X1 U7469 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6756) );
  AOI22_X1 U7470 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6555), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6597), .ZN(n6516) );
  OAI21_X1 U7471 ( .B1(n6756), .B2(n6517), .A(n6516), .ZN(U3192) );
  INV_X1 U7472 ( .A(n6517), .ZN(n6551) );
  INV_X1 U7473 ( .A(n6551), .ZN(n6557) );
  AOI22_X1 U7474 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6555), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6597), .ZN(n6518) );
  OAI21_X1 U7475 ( .B1(n6519), .B2(n6557), .A(n6518), .ZN(U3193) );
  AOI22_X1 U7476 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6555), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6597), .ZN(n6520) );
  OAI21_X1 U7477 ( .B1(n6521), .B2(n6557), .A(n6520), .ZN(U3194) );
  AOI22_X1 U7478 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6555), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6597), .ZN(n6522) );
  OAI21_X1 U7479 ( .B1(n6523), .B2(n6557), .A(n6522), .ZN(U3195) );
  AOI22_X1 U7480 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6555), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6597), .ZN(n6524) );
  OAI21_X1 U7481 ( .B1(n6525), .B2(n6557), .A(n6524), .ZN(U3196) );
  AOI22_X1 U7482 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6548), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6597), .ZN(n6526) );
  OAI21_X1 U7483 ( .B1(n6527), .B2(n6557), .A(n6526), .ZN(U3197) );
  AOI22_X1 U7484 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6548), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6597), .ZN(n6528) );
  OAI21_X1 U7485 ( .B1(n6529), .B2(n6557), .A(n6528), .ZN(U3198) );
  AOI22_X1 U7486 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6548), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6597), .ZN(n6530) );
  OAI21_X1 U7487 ( .B1(n6531), .B2(n6557), .A(n6530), .ZN(U3199) );
  AOI22_X1 U7488 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6548), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6597), .ZN(n6532) );
  OAI21_X1 U7489 ( .B1(n6533), .B2(n6557), .A(n6532), .ZN(U3200) );
  AOI22_X1 U7490 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6548), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6597), .ZN(n6534) );
  OAI21_X1 U7491 ( .B1(n5674), .B2(n6557), .A(n6534), .ZN(U3201) );
  AOI22_X1 U7492 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6551), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6597), .ZN(n6535) );
  OAI21_X1 U7493 ( .B1(n5674), .B2(n6553), .A(n6535), .ZN(U3202) );
  AOI22_X1 U7494 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6548), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6597), .ZN(n6536) );
  OAI21_X1 U7495 ( .B1(n6537), .B2(n6557), .A(n6536), .ZN(U3203) );
  AOI22_X1 U7496 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6548), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6597), .ZN(n6538) );
  OAI21_X1 U7497 ( .B1(n6540), .B2(n6557), .A(n6538), .ZN(U3204) );
  AOI22_X1 U7498 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6551), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6597), .ZN(n6539) );
  OAI21_X1 U7499 ( .B1(n6540), .B2(n6553), .A(n6539), .ZN(U3205) );
  AOI22_X1 U7500 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6548), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6597), .ZN(n6541) );
  OAI21_X1 U7501 ( .B1(n6542), .B2(n6557), .A(n6541), .ZN(U3206) );
  AOI22_X1 U7502 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6548), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6597), .ZN(n6543) );
  OAI21_X1 U7503 ( .B1(n6545), .B2(n6557), .A(n6543), .ZN(U3207) );
  AOI22_X1 U7504 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6551), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6597), .ZN(n6544) );
  OAI21_X1 U7505 ( .B1(n6545), .B2(n6553), .A(n6544), .ZN(U3208) );
  AOI22_X1 U7506 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6555), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6597), .ZN(n6546) );
  OAI21_X1 U7507 ( .B1(n6547), .B2(n6557), .A(n6546), .ZN(U3209) );
  AOI222_X1 U7508 ( .A1(n6548), .A2(REIP_REG_27__SCAN_IN), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6597), .C1(REIP_REG_28__SCAN_IN), .C2(
        n6551), .ZN(n6549) );
  INV_X1 U7509 ( .A(n6549), .ZN(U3210) );
  AOI22_X1 U7510 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6555), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6597), .ZN(n6550) );
  OAI21_X1 U7511 ( .B1(n6554), .B2(n6557), .A(n6550), .ZN(U3211) );
  AOI22_X1 U7512 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6551), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6597), .ZN(n6552) );
  OAI21_X1 U7513 ( .B1(n6554), .B2(n6553), .A(n6552), .ZN(U3212) );
  AOI22_X1 U7514 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6555), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6597), .ZN(n6556) );
  OAI21_X1 U7515 ( .B1(n6558), .B2(n6557), .A(n6556), .ZN(U3213) );
  MUX2_X1 U7516 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6611), .Z(U3445) );
  MUX2_X1 U7517 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6611), .Z(U3446) );
  MUX2_X1 U7518 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6611), .Z(U3447) );
  MUX2_X1 U7519 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6611), .Z(U3448) );
  INV_X1 U7520 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6561) );
  INV_X1 U7521 ( .A(n6562), .ZN(n6559) );
  AOI21_X1 U7522 ( .B1(n6561), .B2(n6560), .A(n6559), .ZN(U3451) );
  OAI21_X1 U7523 ( .B1(n6564), .B2(n6563), .A(n6562), .ZN(U3452) );
  INV_X1 U7524 ( .A(n6565), .ZN(n6567) );
  OAI211_X1 U7525 ( .C1(n6718), .C2(n6568), .A(n6567), .B(n6566), .ZN(U3453)
         );
  AOI22_X1 U7526 ( .A1(n6572), .A2(n6571), .B1(n6570), .B2(n6569), .ZN(n6573)
         );
  INV_X1 U7527 ( .A(n6573), .ZN(n6574) );
  OAI22_X1 U7528 ( .A1(n6581), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(n6574), .B2(n6583), .ZN(n6575) );
  INV_X1 U7529 ( .A(n6575), .ZN(U3456) );
  INV_X1 U7530 ( .A(n6576), .ZN(n6577) );
  AOI21_X1 U7531 ( .B1(n6577), .B2(n6718), .A(STATE2_REG_1__SCAN_IN), .ZN(
        n6579) );
  OAI22_X1 U7532 ( .A1(n6580), .A2(n6579), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6578), .ZN(n6582) );
  AOI22_X1 U7533 ( .A1(n6583), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(n6582), .B2(n6581), .ZN(n6584) );
  OAI21_X1 U7534 ( .B1(n6586), .B2(n6585), .A(n6584), .ZN(U3461) );
  AOI21_X1 U7535 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6588) );
  AOI22_X1 U7536 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6588), .B2(n6587), .ZN(n6590) );
  INV_X1 U7537 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6589) );
  AOI22_X1 U7538 ( .A1(n6591), .A2(n6590), .B1(n6589), .B2(n6594), .ZN(U3468)
         );
  INV_X1 U7539 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6595) );
  NOR2_X1 U7540 ( .A1(n6594), .A2(REIP_REG_1__SCAN_IN), .ZN(n6592) );
  AOI22_X1 U7541 ( .A1(n6595), .A2(n6594), .B1(n6593), .B2(n6592), .ZN(U3469)
         );
  NAND2_X1 U7542 ( .A1(n6597), .A2(W_R_N_REG_SCAN_IN), .ZN(n6596) );
  OAI21_X1 U7543 ( .B1(n6597), .B2(READREQUEST_REG_SCAN_IN), .A(n6596), .ZN(
        U3470) );
  OAI211_X1 U7544 ( .C1(READY_N), .C2(n6600), .A(n6599), .B(n6598), .ZN(n6610)
         );
  AOI21_X1 U7545 ( .B1(n2984), .B2(n6602), .A(n6601), .ZN(n6604) );
  AOI21_X1 U7546 ( .B1(n6605), .B2(n6604), .A(n6603), .ZN(n6606) );
  OAI21_X1 U7547 ( .B1(n6607), .B2(n6606), .A(n6610), .ZN(n6608) );
  OAI21_X1 U7548 ( .B1(n6610), .B2(n6609), .A(n6608), .ZN(U3472) );
  MUX2_X1 U7549 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6611), .Z(U3473) );
  OAI22_X1 U7550 ( .A1(n6613), .A2(keyinput46), .B1(n5074), .B2(keyinput27), 
        .ZN(n6612) );
  AOI221_X1 U7551 ( .B1(n6613), .B2(keyinput46), .C1(keyinput27), .C2(n5074), 
        .A(n6612), .ZN(n6775) );
  OAI22_X1 U7552 ( .A1(n3290), .A2(keyinput35), .B1(n4953), .B2(keyinput9), 
        .ZN(n6614) );
  AOI221_X1 U7553 ( .B1(n3290), .B2(keyinput35), .C1(keyinput9), .C2(n4953), 
        .A(n6614), .ZN(n6774) );
  OAI22_X1 U7554 ( .A1(n6617), .A2(keyinput34), .B1(n6616), .B2(keyinput39), 
        .ZN(n6615) );
  AOI221_X1 U7555 ( .B1(n6617), .B2(keyinput34), .C1(keyinput39), .C2(n6616), 
        .A(n6615), .ZN(n6630) );
  INV_X1 U7556 ( .A(keyinput38), .ZN(n6619) );
  OAI22_X1 U7557 ( .A1(keyinput15), .A2(n6620), .B1(n6619), .B2(
        ADDRESS_REG_28__SCAN_IN), .ZN(n6618) );
  AOI221_X1 U7558 ( .B1(n6620), .B2(keyinput15), .C1(n6619), .C2(
        ADDRESS_REG_28__SCAN_IN), .A(n6618), .ZN(n6629) );
  INV_X1 U7559 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n6623) );
  INV_X1 U7560 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n6622) );
  OAI22_X1 U7561 ( .A1(n6623), .A2(keyinput7), .B1(n6622), .B2(keyinput32), 
        .ZN(n6621) );
  AOI221_X1 U7562 ( .B1(n6623), .B2(keyinput7), .C1(keyinput32), .C2(n6622), 
        .A(n6621), .ZN(n6628) );
  OAI22_X1 U7563 ( .A1(n6626), .A2(keyinput59), .B1(n6625), .B2(keyinput28), 
        .ZN(n6624) );
  AOI221_X1 U7564 ( .B1(n6626), .B2(keyinput59), .C1(keyinput28), .C2(n6625), 
        .A(n6624), .ZN(n6627) );
  NAND4_X1 U7565 ( .A1(n6630), .A2(n6629), .A3(n6628), .A4(n6627), .ZN(n6638)
         );
  INV_X1 U7566 ( .A(keyinput17), .ZN(n6632) );
  AOI22_X1 U7567 ( .A1(n6633), .A2(keyinput42), .B1(DATAWIDTH_REG_0__SCAN_IN), 
        .B2(n6632), .ZN(n6631) );
  OAI221_X1 U7568 ( .B1(n6633), .B2(keyinput42), .C1(n6632), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(n6631), .ZN(n6637) );
  XOR2_X1 U7569 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .B(keyinput14), .Z(n6636)
         );
  XNOR2_X1 U7570 ( .A(n6634), .B(keyinput31), .ZN(n6635) );
  NOR4_X1 U7571 ( .A1(n6638), .A2(n6637), .A3(n6636), .A4(n6635), .ZN(n6773)
         );
  NOR2_X1 U7572 ( .A1(keyinput52), .A2(keyinput63), .ZN(n6639) );
  NAND3_X1 U7573 ( .A1(keyinput20), .A2(keyinput56), .A3(n6639), .ZN(n6644) );
  NAND3_X1 U7574 ( .A1(keyinput60), .A2(keyinput57), .A3(keyinput41), .ZN(
        n6643) );
  NOR4_X1 U7575 ( .A1(keyinput29), .A2(keyinput4), .A3(keyinput10), .A4(
        keyinput21), .ZN(n6641) );
  INV_X1 U7576 ( .A(keyinput8), .ZN(n6640) );
  NAND4_X1 U7577 ( .A1(keyinput5), .A2(keyinput33), .A3(n6641), .A4(n6640), 
        .ZN(n6642) );
  NOR4_X1 U7578 ( .A1(keyinput30), .A2(n6644), .A3(n6643), .A4(n6642), .ZN(
        n6667) );
  NAND3_X1 U7579 ( .A1(keyinput23), .A2(keyinput47), .A3(keyinput50), .ZN(
        n6650) );
  INV_X1 U7580 ( .A(keyinput16), .ZN(n6645) );
  NAND4_X1 U7581 ( .A1(keyinput54), .A2(keyinput19), .A3(keyinput49), .A4(
        n6645), .ZN(n6649) );
  NOR3_X1 U7582 ( .A1(keyinput3), .A2(keyinput43), .A3(keyinput13), .ZN(n6647)
         );
  NOR3_X1 U7583 ( .A1(keyinput12), .A2(keyinput62), .A3(keyinput2), .ZN(n6646)
         );
  NAND4_X1 U7584 ( .A1(keyinput0), .A2(n6647), .A3(keyinput45), .A4(n6646), 
        .ZN(n6648) );
  NOR4_X1 U7585 ( .A1(keyinput24), .A2(n6650), .A3(n6649), .A4(n6648), .ZN(
        n6666) );
  NAND3_X1 U7586 ( .A1(keyinput27), .A2(keyinput17), .A3(keyinput14), .ZN(
        n6657) );
  NOR2_X1 U7587 ( .A1(keyinput34), .A2(keyinput38), .ZN(n6651) );
  NAND3_X1 U7588 ( .A1(keyinput15), .A2(keyinput31), .A3(n6651), .ZN(n6656) );
  NOR3_X1 U7589 ( .A1(keyinput35), .A2(keyinput9), .A3(keyinput46), .ZN(n6654)
         );
  INV_X1 U7590 ( .A(keyinput59), .ZN(n6652) );
  NOR3_X1 U7591 ( .A1(keyinput28), .A2(keyinput7), .A3(n6652), .ZN(n6653) );
  NAND4_X1 U7592 ( .A1(keyinput11), .A2(n6654), .A3(keyinput39), .A4(n6653), 
        .ZN(n6655) );
  NOR4_X1 U7593 ( .A1(keyinput42), .A2(n6657), .A3(n6656), .A4(n6655), .ZN(
        n6665) );
  NAND3_X1 U7594 ( .A1(keyinput32), .A2(keyinput22), .A3(keyinput1), .ZN(n6663) );
  INV_X1 U7595 ( .A(keyinput53), .ZN(n6658) );
  NAND4_X1 U7596 ( .A1(keyinput61), .A2(keyinput55), .A3(keyinput48), .A4(
        n6658), .ZN(n6662) );
  NOR3_X1 U7597 ( .A1(keyinput36), .A2(keyinput40), .A3(keyinput18), .ZN(n6660) );
  INV_X1 U7598 ( .A(keyinput51), .ZN(n6679) );
  NOR3_X1 U7599 ( .A1(keyinput37), .A2(keyinput44), .A3(n6679), .ZN(n6659) );
  NAND4_X1 U7600 ( .A1(keyinput25), .A2(n6660), .A3(keyinput26), .A4(n6659), 
        .ZN(n6661) );
  NOR4_X1 U7601 ( .A1(keyinput58), .A2(n6663), .A3(n6662), .A4(n6661), .ZN(
        n6664) );
  NAND4_X1 U7602 ( .A1(n6667), .A2(n6666), .A3(n6665), .A4(n6664), .ZN(n6668)
         );
  AOI21_X1 U7603 ( .B1(keyinput6), .B2(n6668), .A(n6701), .ZN(n6771) );
  INV_X1 U7604 ( .A(keyinput37), .ZN(n6670) );
  OAI22_X1 U7605 ( .A1(keyinput18), .A2(n6671), .B1(n6670), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6669) );
  AOI221_X1 U7606 ( .B1(n6671), .B2(keyinput18), .C1(n6670), .C2(
        DATAO_REG_1__SCAN_IN), .A(n6669), .ZN(n6684) );
  INV_X1 U7607 ( .A(keyinput40), .ZN(n6673) );
  OAI22_X1 U7608 ( .A1(n6674), .A2(keyinput36), .B1(n6673), .B2(
        BYTEENABLE_REG_1__SCAN_IN), .ZN(n6672) );
  AOI221_X1 U7609 ( .B1(n6674), .B2(keyinput36), .C1(BYTEENABLE_REG_1__SCAN_IN), .C2(n6673), .A(n6672), .ZN(n6683) );
  INV_X1 U7610 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n6677) );
  INV_X1 U7611 ( .A(keyinput33), .ZN(n6676) );
  OAI22_X1 U7612 ( .A1(n6677), .A2(keyinput26), .B1(n6676), .B2(BS16_N), .ZN(
        n6675) );
  AOI221_X1 U7613 ( .B1(n6677), .B2(keyinput26), .C1(BS16_N), .C2(n6676), .A(
        n6675), .ZN(n6682) );
  OAI22_X1 U7614 ( .A1(keyinput44), .A2(n6680), .B1(n6679), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6678) );
  AOI221_X1 U7615 ( .B1(n6680), .B2(keyinput44), .C1(n6679), .C2(
        DATAO_REG_7__SCAN_IN), .A(n6678), .ZN(n6681) );
  NAND4_X1 U7616 ( .A1(n6684), .A2(n6683), .A3(n6682), .A4(n6681), .ZN(n6770)
         );
  INV_X1 U7617 ( .A(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n6687) );
  INV_X1 U7618 ( .A(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n6686) );
  OAI22_X1 U7619 ( .A1(n6687), .A2(keyinput1), .B1(n6686), .B2(keyinput61), 
        .ZN(n6685) );
  AOI221_X1 U7620 ( .B1(n6687), .B2(keyinput1), .C1(keyinput61), .C2(n6686), 
        .A(n6685), .ZN(n6700) );
  INV_X1 U7621 ( .A(keyinput58), .ZN(n6689) );
  OAI22_X1 U7622 ( .A1(n6690), .A2(keyinput22), .B1(n6689), .B2(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n6688) );
  AOI221_X1 U7623 ( .B1(n6690), .B2(keyinput22), .C1(DATAWIDTH_REG_23__SCAN_IN), .C2(n6689), .A(n6688), .ZN(n6699) );
  INV_X1 U7624 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n6693) );
  INV_X1 U7625 ( .A(keyinput25), .ZN(n6692) );
  OAI22_X1 U7626 ( .A1(n6693), .A2(keyinput48), .B1(n6692), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n6691) );
  AOI221_X1 U7627 ( .B1(n6693), .B2(keyinput48), .C1(DATAO_REG_16__SCAN_IN), 
        .C2(n6692), .A(n6691), .ZN(n6698) );
  OAI22_X1 U7628 ( .A1(n6696), .A2(keyinput53), .B1(n6695), .B2(keyinput55), 
        .ZN(n6694) );
  AOI221_X1 U7629 ( .B1(n6696), .B2(keyinput53), .C1(keyinput55), .C2(n6695), 
        .A(n6694), .ZN(n6697) );
  NAND4_X1 U7630 ( .A1(n6700), .A2(n6699), .A3(n6698), .A4(n6697), .ZN(n6769)
         );
  INV_X1 U7631 ( .A(keyinput52), .ZN(n6705) );
  AOI22_X1 U7632 ( .A1(n6706), .A2(keyinput8), .B1(DATAO_REG_0__SCAN_IN), .B2(
        n6705), .ZN(n6704) );
  OAI221_X1 U7633 ( .B1(n6706), .B2(keyinput8), .C1(n6705), .C2(
        DATAO_REG_0__SCAN_IN), .A(n6704), .ZN(n6714) );
  AOI22_X1 U7634 ( .A1(n4817), .A2(keyinput20), .B1(keyinput56), .B2(n6708), 
        .ZN(n6707) );
  OAI221_X1 U7635 ( .B1(n4817), .B2(keyinput20), .C1(n6708), .C2(keyinput56), 
        .A(n6707), .ZN(n6713) );
  INV_X1 U7636 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6711) );
  AOI22_X1 U7637 ( .A1(n6711), .A2(keyinput63), .B1(keyinput60), .B2(n6710), 
        .ZN(n6709) );
  OAI221_X1 U7638 ( .B1(n6711), .B2(keyinput63), .C1(n6710), .C2(keyinput60), 
        .A(n6709), .ZN(n6712) );
  NOR4_X1 U7639 ( .A1(n6715), .A2(n6714), .A3(n6713), .A4(n6712), .ZN(n6767)
         );
  INV_X1 U7640 ( .A(keyinput21), .ZN(n6717) );
  AOI22_X1 U7641 ( .A1(n6718), .A2(keyinput23), .B1(ADDRESS_REG_7__SCAN_IN), 
        .B2(n6717), .ZN(n6716) );
  OAI221_X1 U7642 ( .B1(n6718), .B2(keyinput23), .C1(n6717), .C2(
        ADDRESS_REG_7__SCAN_IN), .A(n6716), .ZN(n6731) );
  INV_X1 U7643 ( .A(DATAI_30_), .ZN(n6720) );
  AOI22_X1 U7644 ( .A1(n6721), .A2(keyinput57), .B1(keyinput30), .B2(n6720), 
        .ZN(n6719) );
  OAI221_X1 U7645 ( .B1(n6721), .B2(keyinput57), .C1(n6720), .C2(keyinput30), 
        .A(n6719), .ZN(n6730) );
  INV_X1 U7646 ( .A(keyinput41), .ZN(n6724) );
  INV_X1 U7647 ( .A(keyinput29), .ZN(n6723) );
  AOI22_X1 U7648 ( .A1(n6724), .A2(MEMORYFETCH_REG_SCAN_IN), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6723), .ZN(n6722) );
  OAI221_X1 U7649 ( .B1(n6724), .B2(MEMORYFETCH_REG_SCAN_IN), .C1(n6723), .C2(
        ADDRESS_REG_26__SCAN_IN), .A(n6722), .ZN(n6729) );
  XOR2_X1 U7650 ( .A(n6725), .B(keyinput10), .Z(n6727) );
  XNOR2_X1 U7651 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .B(keyinput4), .ZN(n6726)
         );
  NAND2_X1 U7652 ( .A1(n6727), .A2(n6726), .ZN(n6728) );
  NOR4_X1 U7653 ( .A1(n6731), .A2(n6730), .A3(n6729), .A4(n6728), .ZN(n6766)
         );
  INV_X1 U7654 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n6734) );
  AOI22_X1 U7655 ( .A1(n6734), .A2(keyinput24), .B1(keyinput47), .B2(n6733), 
        .ZN(n6732) );
  OAI221_X1 U7656 ( .B1(n6734), .B2(keyinput24), .C1(n6733), .C2(keyinput47), 
        .A(n6732), .ZN(n6747) );
  INV_X1 U7657 ( .A(keyinput50), .ZN(n6736) );
  AOI22_X1 U7658 ( .A1(n6737), .A2(keyinput3), .B1(UWORD_REG_6__SCAN_IN), .B2(
        n6736), .ZN(n6735) );
  OAI221_X1 U7659 ( .B1(n6737), .B2(keyinput3), .C1(n6736), .C2(
        UWORD_REG_6__SCAN_IN), .A(n6735), .ZN(n6746) );
  AOI22_X1 U7660 ( .A1(n6740), .A2(keyinput43), .B1(n6739), .B2(keyinput13), 
        .ZN(n6738) );
  OAI221_X1 U7661 ( .B1(n6740), .B2(keyinput43), .C1(n6739), .C2(keyinput13), 
        .A(n6738), .ZN(n6745) );
  INV_X1 U7662 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n6743) );
  INV_X1 U7663 ( .A(keyinput54), .ZN(n6742) );
  AOI22_X1 U7664 ( .A1(n6743), .A2(keyinput0), .B1(DATAO_REG_25__SCAN_IN), 
        .B2(n6742), .ZN(n6741) );
  OAI221_X1 U7665 ( .B1(n6743), .B2(keyinput0), .C1(n6742), .C2(
        DATAO_REG_25__SCAN_IN), .A(n6741), .ZN(n6744) );
  NOR4_X1 U7666 ( .A1(n6747), .A2(n6746), .A3(n6745), .A4(n6744), .ZN(n6765)
         );
  AOI22_X1 U7667 ( .A1(n6750), .A2(keyinput16), .B1(n6749), .B2(keyinput19), 
        .ZN(n6748) );
  OAI221_X1 U7668 ( .B1(n6750), .B2(keyinput16), .C1(n6749), .C2(keyinput19), 
        .A(n6748), .ZN(n6763) );
  INV_X1 U7669 ( .A(DATAI_28_), .ZN(n6753) );
  INV_X1 U7670 ( .A(keyinput49), .ZN(n6752) );
  AOI22_X1 U7671 ( .A1(n6753), .A2(keyinput12), .B1(DATAWIDTH_REG_18__SCAN_IN), 
        .B2(n6752), .ZN(n6751) );
  OAI221_X1 U7672 ( .B1(n6753), .B2(keyinput12), .C1(n6752), .C2(
        DATAWIDTH_REG_18__SCAN_IN), .A(n6751), .ZN(n6762) );
  INV_X1 U7673 ( .A(keyinput45), .ZN(n6755) );
  AOI22_X1 U7674 ( .A1(n6756), .A2(keyinput62), .B1(ADDRESS_REG_13__SCAN_IN), 
        .B2(n6755), .ZN(n6754) );
  OAI221_X1 U7675 ( .B1(n6756), .B2(keyinput62), .C1(n6755), .C2(
        ADDRESS_REG_13__SCAN_IN), .A(n6754), .ZN(n6761) );
  INV_X1 U7676 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n6759) );
  AOI22_X1 U7677 ( .A1(n6759), .A2(keyinput2), .B1(keyinput11), .B2(n6758), 
        .ZN(n6757) );
  OAI221_X1 U7678 ( .B1(n6759), .B2(keyinput2), .C1(n6758), .C2(keyinput11), 
        .A(n6757), .ZN(n6760) );
  NOR4_X1 U7679 ( .A1(n6763), .A2(n6762), .A3(n6761), .A4(n6760), .ZN(n6764)
         );
  NAND4_X1 U7680 ( .A1(n6767), .A2(n6766), .A3(n6765), .A4(n6764), .ZN(n6768)
         );
  NOR4_X1 U7681 ( .A1(n6771), .A2(n6770), .A3(n6769), .A4(n6768), .ZN(n6772)
         );
  NAND4_X1 U7682 ( .A1(n6775), .A2(n6774), .A3(n6773), .A4(n6772), .ZN(n6789)
         );
  NAND2_X1 U7683 ( .A1(n6776), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6785)
         );
  OAI22_X1 U7684 ( .A1(n6780), .A2(n6779), .B1(n6778), .B2(n6777), .ZN(n6781)
         );
  AOI21_X1 U7685 ( .B1(n6783), .B2(n6782), .A(n6781), .ZN(n6784) );
  OAI211_X1 U7686 ( .C1(n6787), .C2(n6786), .A(n6785), .B(n6784), .ZN(n6788)
         );
  XNOR2_X1 U7687 ( .A(n6789), .B(n6788), .ZN(U3139) );
  INV_X1 U4207 ( .A(n3346), .ZN(n3309) );
  BUF_X1 U4221 ( .A(n3895), .Z(n4081) );
  CLKBUF_X1 U3436 ( .A(n3239), .Z(n2983) );
  CLKBUF_X1 U3437 ( .A(n3310), .Z(n4277) );
  CLKBUF_X2 U3443 ( .A(n3255), .Z(n3227) );
  CLKBUF_X1 U34690 ( .A(n6030), .Z(n6036) );
  AOI211_X2 U3816 ( .C1(n6364), .C2(n6231), .A(n6228), .B(n6362), .ZN(n6259)
         );
endmodule

