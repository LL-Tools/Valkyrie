

module b22_C_SARLock_k_64_1 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6437, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410;

  OAI21_X1 U7186 ( .B1(n13015), .B2(n7351), .A(n13014), .ZN(n13258) );
  INV_X2 U7187 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7188 ( .A(n8639), .ZN(n9032) );
  OR2_X1 U7189 ( .A1(n10506), .A2(n13550), .ZN(n14788) );
  NAND2_X1 U7190 ( .A1(n7332), .A2(n14328), .ZN(n14329) );
  NAND2_X2 U7192 ( .A1(n8615), .A2(n6437), .ZN(n8644) );
  NAND2_X1 U7193 ( .A1(n6648), .A2(n6647), .ZN(n10722) );
  CLKBUF_X2 U7195 ( .A(n9211), .Z(n9513) );
  INV_X1 U7197 ( .A(n9429), .ZN(n9799) );
  AND3_X1 U7198 ( .A1(n6728), .A2(n9200), .A3(n6727), .ZN(n9135) );
  AND2_X1 U7199 ( .A1(n11430), .A2(n7254), .ZN(n6630) );
  INV_X2 U7200 ( .A(n7904), .ZN(n8423) );
  INV_X1 U7201 ( .A(n11836), .ZN(n11831) );
  INV_X2 U7202 ( .A(n11837), .ZN(n11827) );
  INV_X1 U7203 ( .A(n13514), .ZN(n9399) );
  INV_X1 U7204 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9286) );
  NAND2_X1 U7205 ( .A1(n11860), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8609) );
  INV_X1 U7206 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n9027) );
  INV_X1 U7207 ( .A(n8399), .ZN(n8385) );
  XNOR2_X1 U7208 ( .A(n13255), .B(n13027), .ZN(n13013) );
  INV_X1 U7209 ( .A(n13503), .ZN(n9560) );
  XNOR2_X1 U7210 ( .A(n14329), .B(n7331), .ZN(n14368) );
  NAND2_X1 U7211 ( .A1(n8649), .A2(n8648), .ZN(n15143) );
  NOR2_X1 U7213 ( .A1(n7823), .A2(n7822), .ZN(n14845) );
  MUX2_X1 U7214 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14258), .S(n14822), .Z(
        n14154) );
  NAND2_X2 U7215 ( .A1(n9439), .A2(n9438), .ZN(n14049) );
  NAND4_X1 U7216 ( .A1(n8734), .A2(n8733), .A3(n8732), .A4(n8731), .ZN(n12283)
         );
  XNOR2_X1 U7217 ( .A(n7742), .B(n7741), .ZN(n7757) );
  OAI21_X2 U7218 ( .B1(n13660), .B2(n13659), .A(n13658), .ZN(n13662) );
  NOR2_X4 U7219 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n10404) );
  AOI21_X2 U7220 ( .B1(n14164), .B2(n14793), .A(n13983), .ZN(n7139) );
  XNOR2_X2 U7221 ( .A(n11558), .B(n7064), .ZN(n7059) );
  OAI211_X1 U7222 ( .C1(n13671), .C2(n13668), .A(n13670), .B(n13667), .ZN(
        n13679) );
  INV_X1 U7223 ( .A(n8614), .ZN(n6437) );
  INV_X2 U7225 ( .A(n6437), .ZN(n6439) );
  NAND2_X2 U7226 ( .A1(n8233), .A2(n8232), .ZN(n13275) );
  NAND2_X2 U7227 ( .A1(n9276), .A2(n9275), .ZN(n13618) );
  NAND2_X2 U7228 ( .A1(n8259), .A2(n8258), .ZN(n13269) );
  NOR2_X2 U7229 ( .A1(n14426), .A2(n14389), .ZN(n14391) );
  OAI21_X2 U7230 ( .B1(n6446), .B2(P3_REG2_REG_1__SCAN_IN), .A(n6920), .ZN(
        n10415) );
  BUF_X8 U7231 ( .A(n12437), .Z(n6446) );
  XNOR2_X2 U7232 ( .A(n14049), .B(n13777), .ZN(n14054) );
  NAND2_X2 U7233 ( .A1(n9291), .A2(n9290), .ZN(n14563) );
  NAND2_X2 U7234 ( .A1(n8351), .A2(n8350), .ZN(n13255) );
  NOR2_X4 U7235 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7788) );
  XNOR2_X2 U7236 ( .A(n14326), .B(n7333), .ZN(n14370) );
  NAND2_X2 U7237 ( .A1(n14325), .A2(n6915), .ZN(n14326) );
  CLKBUF_X1 U7238 ( .A(n8395), .Z(n6440) );
  AND2_X1 U7239 ( .A1(n7279), .A2(n7757), .ZN(n8395) );
  NOR2_X2 U7240 ( .A1(n11961), .A2(n11960), .ZN(n11959) );
  OAI21_X2 U7241 ( .B1(n10985), .B2(n10991), .A(n6902), .ZN(n11961) );
  XNOR2_X2 U7242 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n14373) );
  AOI21_X1 U7243 ( .B1(n7338), .B2(n11722), .A(n6459), .ZN(n7337) );
  XNOR2_X1 U7244 ( .A(n6618), .B(n11644), .ZN(n12032) );
  NAND2_X1 U7245 ( .A1(n11903), .A2(n11637), .ZN(n12014) );
  NOR2_X1 U7246 ( .A1(n11559), .A2(n7062), .ZN(n7058) );
  NAND2_X2 U7247 ( .A1(n9921), .A2(n9922), .ZN(n9955) );
  INV_X1 U7248 ( .A(n15144), .ZN(n10328) );
  XNOR2_X1 U7249 ( .A(n10330), .B(n11622), .ZN(n10986) );
  INV_X1 U7250 ( .A(n14757), .ZN(n10058) );
  INV_X1 U7251 ( .A(n13795), .ZN(n10588) );
  NAND2_X1 U7252 ( .A1(n9776), .A2(n9775), .ZN(n13228) );
  INV_X1 U7253 ( .A(n13798), .ZN(n7185) );
  INV_X1 U7254 ( .A(n8664), .ZN(n8793) );
  INV_X2 U7255 ( .A(n9010), .ZN(n6443) );
  INV_X2 U7257 ( .A(n9272), .ZN(n13511) );
  CLKBUF_X2 U7258 ( .A(n13506), .Z(n9562) );
  INV_X1 U7259 ( .A(n10010), .ZN(n10167) );
  NAND2_X1 U7260 ( .A1(n6833), .A2(n8585), .ZN(n12437) );
  OR2_X1 U7261 ( .A1(n7736), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n8479) );
  INV_X8 U7262 ( .A(n9155), .ZN(n7171) );
  AND3_X1 U7263 ( .A1(n6896), .A2(n6867), .A3(n13759), .ZN(n13769) );
  AND2_X1 U7264 ( .A1(n13002), .A2(n13001), .ZN(n13252) );
  AND2_X1 U7265 ( .A1(n7350), .A2(n7352), .ZN(n13015) );
  AOI21_X1 U7266 ( .B1(n7030), .B2(n13228), .A(n7028), .ZN(n13257) );
  AND2_X1 U7267 ( .A1(n11588), .A2(n7389), .ZN(n7388) );
  OAI21_X1 U7268 ( .B1(n13026), .B2(n7284), .A(n7281), .ZN(n12998) );
  NAND2_X1 U7269 ( .A1(n6757), .A2(n6758), .ZN(n13035) );
  OAI211_X1 U7270 ( .C1(n11650), .C2(n6627), .A(n11652), .B(n6625), .ZN(n11943) );
  NAND2_X1 U7271 ( .A1(n13080), .A2(n7335), .ZN(n6757) );
  NAND2_X1 U7272 ( .A1(n7342), .A2(n11720), .ZN(n7341) );
  AND2_X1 U7273 ( .A1(n7297), .A2(n7296), .ZN(n13039) );
  AOI21_X1 U7274 ( .B1(n7337), .B2(n7339), .A(n6531), .ZN(n7335) );
  OR2_X1 U7275 ( .A1(n13090), .A2(n13091), .ZN(n13093) );
  OAI22_X1 U7276 ( .A1(n13117), .A2(n11717), .B1(n13122), .B2(n13140), .ZN(
        n13113) );
  NAND2_X1 U7277 ( .A1(n12014), .A2(n12013), .ZN(n12012) );
  OAI21_X1 U7278 ( .B1(n11710), .B2(n6750), .A(n6748), .ZN(n13133) );
  XNOR2_X1 U7279 ( .A(n8231), .B(n8230), .ZN(n14315) );
  NAND2_X1 U7280 ( .A1(n7058), .A2(n7063), .ZN(n12836) );
  NAND2_X1 U7281 ( .A1(n9462), .A2(n9461), .ZN(n14268) );
  NAND2_X1 U7282 ( .A1(n11953), .A2(n11627), .ZN(n7253) );
  AOI21_X1 U7283 ( .B1(n13201), .B2(n11682), .A(n11681), .ZN(n13185) );
  NAND2_X1 U7284 ( .A1(n13220), .A2(n11679), .ZN(n13201) );
  NAND2_X1 U7285 ( .A1(n7149), .A2(n14241), .ZN(n14143) );
  NAND2_X1 U7286 ( .A1(n8189), .A2(n8188), .ZN(n13286) );
  AND2_X1 U7287 ( .A1(n9414), .A2(n9413), .ZN(n14098) );
  NAND2_X1 U7288 ( .A1(n9416), .A2(n9415), .ZN(n14285) );
  XNOR2_X1 U7289 ( .A(n8250), .B(SI_22_), .ZN(n9428) );
  NAND2_X1 U7290 ( .A1(n13221), .A2(n13222), .ZN(n13220) );
  INV_X1 U7291 ( .A(n11534), .ZN(n7149) );
  NAND2_X1 U7292 ( .A1(n8121), .A2(n8120), .ZN(n13302) );
  OAI21_X1 U7293 ( .B1(n11703), .B2(n11702), .A(n11705), .ZN(n13216) );
  NAND2_X1 U7294 ( .A1(n8164), .A2(n8163), .ZN(n13290) );
  OAI21_X1 U7295 ( .B1(n11356), .B2(n11355), .A(n11357), .ZN(n11703) );
  NAND2_X1 U7296 ( .A1(n8187), .A2(n8186), .ZN(n8208) );
  AND2_X1 U7297 ( .A1(n7169), .A2(n7168), .ZN(n11221) );
  NOR2_X1 U7298 ( .A1(n11068), .A2(n15217), .ZN(n11401) );
  OR2_X1 U7299 ( .A1(n11063), .A2(n13529), .ZN(n11062) );
  XNOR2_X1 U7300 ( .A(n8555), .B(n11373), .ZN(n8635) );
  OR2_X1 U7301 ( .A1(n7685), .A2(n9701), .ZN(n7687) );
  OAI21_X1 U7302 ( .B1(n10874), .B2(n10873), .A(n10875), .ZN(n10913) );
  NAND2_X1 U7303 ( .A1(n7952), .A2(n7951), .ZN(n11089) );
  NAND2_X1 U7304 ( .A1(n7676), .A2(n7071), .ZN(n7968) );
  NAND3_X1 U7305 ( .A1(n7071), .A2(n7676), .A3(n7613), .ZN(n7970) );
  NOR2_X1 U7306 ( .A1(n15401), .A2(n14393), .ZN(n14396) );
  NAND2_X1 U7307 ( .A1(n7675), .A2(SI_10_), .ZN(n7676) );
  OR2_X1 U7308 ( .A1(n7675), .A2(SI_10_), .ZN(n7071) );
  NAND2_X1 U7309 ( .A1(n7948), .A2(n7674), .ZN(n7675) );
  INV_X2 U7310 ( .A(n15159), .ZN(n14498) );
  AOI21_X1 U7311 ( .B1(n11137), .B2(n11138), .A(n6514), .ZN(n6619) );
  NAND2_X1 U7312 ( .A1(n7946), .A2(n7945), .ZN(n7948) );
  OAI21_X1 U7313 ( .B1(n8826), .B2(n10179), .A(n8544), .ZN(n8839) );
  NAND2_X1 U7314 ( .A1(n15398), .A2(n14384), .ZN(n14386) );
  AND2_X1 U7315 ( .A1(n7886), .A2(n7885), .ZN(n9665) );
  AND2_X1 U7316 ( .A1(n9205), .A2(n9204), .ZN(n10507) );
  OR2_X1 U7317 ( .A1(n12283), .A2(n11167), .ZN(n12159) );
  NAND2_X1 U7318 ( .A1(n6623), .A2(n6486), .ZN(n7211) );
  NAND2_X1 U7319 ( .A1(n8666), .A2(n6853), .ZN(n15131) );
  INV_X1 U7320 ( .A(n12143), .ZN(n15174) );
  NAND2_X1 U7321 ( .A1(n6615), .A2(n10058), .ZN(n10580) );
  NAND2_X1 U7322 ( .A1(n7856), .A2(n7855), .ZN(n7858) );
  AND3_X1 U7323 ( .A1(n8756), .A2(n8755), .A3(n8754), .ZN(n11027) );
  OAI211_X1 U7324 ( .C1(n8793), .C2(SI_4_), .A(n8689), .B(n8688), .ZN(n12143)
         );
  OAI211_X1 U7325 ( .C1(n8793), .C2(SI_3_), .A(n8677), .B(n8676), .ZN(n15116)
         );
  NAND4_X1 U7326 ( .A1(n8660), .A2(n8659), .A3(n8658), .A4(n8657), .ZN(n15144)
         );
  OAI211_X1 U7327 ( .C1(n8793), .C2(n9640), .A(n8655), .B(n8654), .ZN(n10268)
         );
  AND2_X1 U7328 ( .A1(n7321), .A2(n6557), .ZN(n14382) );
  NAND2_X1 U7329 ( .A1(n9081), .A2(n9096), .ZN(n9085) );
  NAND2_X1 U7330 ( .A1(n7641), .A2(n7172), .ZN(n10168) );
  NAND2_X2 U7331 ( .A1(n9751), .A2(n13230), .ZN(n9771) );
  NAND2_X1 U7332 ( .A1(n9525), .A2(n13549), .ZN(n14730) );
  OR2_X1 U7333 ( .A1(n15397), .A2(n15396), .ZN(n7321) );
  NOR2_X1 U7334 ( .A1(n7264), .A2(n12108), .ZN(n7263) );
  INV_X1 U7336 ( .A(n9010), .ZN(n12079) );
  NAND2_X1 U7337 ( .A1(n14751), .A2(n14725), .ZN(n14726) );
  NAND2_X1 U7338 ( .A1(n7805), .A2(n6906), .ZN(n7807) );
  NAND2_X2 U7339 ( .A1(n9971), .A2(n9970), .ZN(n11837) );
  NAND2_X1 U7340 ( .A1(n6805), .A2(n6803), .ZN(n7840) );
  AND2_X2 U7341 ( .A1(n9971), .A2(n13564), .ZN(n11826) );
  OR2_X2 U7342 ( .A1(n6914), .A2(n15030), .ZN(n13194) );
  AND2_X1 U7343 ( .A1(n7770), .A2(n6794), .ZN(n8419) );
  OR2_X1 U7344 ( .A1(n10674), .A2(n10474), .ZN(n10676) );
  NOR2_X1 U7345 ( .A1(n8644), .A2(n10220), .ZN(n8645) );
  NAND4_X1 U7346 ( .A1(n7796), .A2(n7795), .A3(n7794), .A4(n7793), .ZN(n12916)
         );
  NAND2_X1 U7347 ( .A1(n10395), .A2(n9155), .ZN(n9010) );
  INV_X1 U7348 ( .A(n13560), .ZN(n14725) );
  OAI22_X1 U7349 ( .A1(n7803), .A2(n7658), .B1(n7801), .B2(SI_2_), .ZN(n7825)
         );
  AND2_X2 U7350 ( .A1(n9398), .A2(n6472), .ZN(n14082) );
  CLKBUF_X2 U7351 ( .A(n11222), .Z(n6914) );
  XNOR2_X1 U7352 ( .A(n9075), .B(n9074), .ZN(n11002) );
  INV_X1 U7353 ( .A(n9149), .ZN(n14302) );
  OAI21_X1 U7354 ( .B1(n9073), .B2(P3_IR_REG_24__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9075) );
  NAND2_X1 U7355 ( .A1(n9073), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9072) );
  INV_X1 U7356 ( .A(n10441), .ZN(n12127) );
  XNOR2_X1 U7357 ( .A(n9143), .B(n14296), .ZN(n9148) );
  OR2_X1 U7358 ( .A1(n7073), .A2(n9027), .ZN(n6987) );
  NAND2_X1 U7359 ( .A1(n8479), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6761) );
  XNOR2_X1 U7360 ( .A(n8612), .B(n8611), .ZN(n8614) );
  XNOR2_X1 U7361 ( .A(n9026), .B(n9025), .ZN(n10441) );
  MUX2_X1 U7362 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8584), .S(
        P3_IR_REG_27__SCAN_IN), .Z(n6833) );
  XNOR2_X1 U7363 ( .A(n8914), .B(n8913), .ZN(n12428) );
  XNOR2_X1 U7364 ( .A(n9030), .B(n9029), .ZN(n10181) );
  AND2_X1 U7365 ( .A1(n6804), .A2(n7662), .ZN(n6803) );
  NAND2_X1 U7366 ( .A1(n7743), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7744) );
  OR2_X1 U7367 ( .A1(n9028), .A2(n9027), .ZN(n9030) );
  NAND2_X1 U7368 ( .A1(n9153), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7145) );
  OR2_X1 U7369 ( .A1(n9024), .A2(n9027), .ZN(n9026) );
  NAND2_X1 U7370 ( .A1(n8486), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7709) );
  NAND2_X1 U7371 ( .A1(n14299), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9143) );
  NAND2_X1 U7372 ( .A1(n7317), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7742) );
  NAND2_X1 U7373 ( .A1(n9140), .A2(n9578), .ZN(n9153) );
  AND2_X1 U7374 ( .A1(n8897), .A2(n8913), .ZN(n9028) );
  AND2_X1 U7375 ( .A1(n7572), .A2(n6565), .ZN(n7251) );
  AND3_X2 U7376 ( .A1(n6838), .A2(n6837), .A3(n6835), .ZN(n8897) );
  AND2_X1 U7377 ( .A1(n7522), .A2(n7740), .ZN(n7316) );
  AND2_X1 U7378 ( .A1(n7573), .A2(n8913), .ZN(n7572) );
  AND3_X1 U7379 ( .A1(n7728), .A2(n7729), .A3(n7503), .ZN(n7731) );
  AND2_X1 U7380 ( .A1(n7523), .A2(n7708), .ZN(n7522) );
  NOR2_X1 U7381 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n7523) );
  AND2_X1 U7382 ( .A1(n8580), .A2(n6836), .ZN(n6835) );
  INV_X1 U7383 ( .A(n8687), .ZN(n6838) );
  AND2_X2 U7384 ( .A1(n7581), .A2(n7582), .ZN(n9619) );
  AND2_X1 U7385 ( .A1(n8583), .A2(n7574), .ZN(n7573) );
  AND3_X1 U7386 ( .A1(n8491), .A2(n7503), .A3(n7697), .ZN(n7704) );
  AND3_X1 U7387 ( .A1(n7726), .A2(n7694), .A3(n7693), .ZN(n8491) );
  NAND2_X1 U7388 ( .A1(n10404), .A2(n8665), .ZN(n8687) );
  AND4_X1 U7389 ( .A1(n8579), .A2(n8578), .A3(n8842), .A4(n8577), .ZN(n8580)
         );
  AND2_X1 U7390 ( .A1(n9129), .A2(n9190), .ZN(n7144) );
  NAND4_X1 U7391 ( .A1(n7652), .A2(n13935), .A3(n7651), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7581) );
  NAND2_X1 U7392 ( .A1(n7580), .A2(n7583), .ZN(n7582) );
  AND2_X1 U7393 ( .A1(n7721), .A2(n7698), .ZN(n6708) );
  AND2_X1 U7394 ( .A1(n6760), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14374) );
  AND3_X1 U7395 ( .A1(n7696), .A2(n7695), .A3(n7712), .ZN(n7503) );
  AND3_X1 U7396 ( .A1(n7701), .A2(n7700), .A3(n7699), .ZN(n7729) );
  INV_X1 U7397 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7574) );
  NOR2_X1 U7398 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n8573) );
  NOR2_X1 U7399 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n8575) );
  NOR2_X1 U7400 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n7726) );
  NOR2_X1 U7401 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n8574) );
  NOR2_X1 U7402 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n7696) );
  NOR2_X1 U7403 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n7695) );
  AND2_X1 U7404 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7583) );
  NOR2_X1 U7405 ( .A1(P3_ADDR_REG_19__SCAN_IN), .A2(P2_RD_REG_SCAN_IN), .ZN(
        n7580) );
  INV_X1 U7406 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n13935) );
  INV_X1 U7407 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7652) );
  INV_X4 U7408 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7409 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n8578) );
  NOR2_X1 U7410 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .ZN(
        n8579) );
  INV_X1 U7411 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9025) );
  INV_X1 U7412 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9129) );
  INV_X1 U7413 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7842) );
  NOR2_X1 U7414 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n7701) );
  NOR2_X1 U7415 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n7700) );
  NOR2_X1 U7416 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n7699) );
  INV_X1 U7417 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n9071) );
  NAND2_X2 U7418 ( .A1(n7212), .A2(n7211), .ZN(n12122) );
  OAI21_X2 U7419 ( .B1(n9271), .B2(n7904), .A(n7975), .ZN(n15027) );
  AOI21_X2 U7420 ( .B1(n7253), .B2(n6621), .A(n6551), .ZN(n11903) );
  NAND2_X2 U7421 ( .A1(n7846), .A2(n7845), .ZN(n10240) );
  AOI22_X1 U7422 ( .A1(n8146), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8145), .B2(
        n14858), .ZN(n7845) );
  INV_X4 U7423 ( .A(n7219), .ZN(n8638) );
  OR2_X1 U7424 ( .A1(n6914), .A2(n15030), .ZN(n6444) );
  XNOR2_X2 U7425 ( .A(n7707), .B(n7740), .ZN(n8497) );
  NOR2_X2 U7426 ( .A1(n14066), .A2(n14049), .ZN(n7159) );
  XNOR2_X2 U7428 ( .A(n7709), .B(n7708), .ZN(n13356) );
  NAND3_X2 U7429 ( .A1(n8640), .A2(n7213), .A3(n7215), .ZN(n15124) );
  OR2_X1 U7430 ( .A1(n8644), .A2(n15155), .ZN(n8640) );
  AND2_X1 U7431 ( .A1(n7214), .A2(n7217), .ZN(n7213) );
  AND2_X4 U7432 ( .A1(n9771), .A2(n9752), .ZN(n11584) );
  OAI21_X2 U7433 ( .B1(n12023), .B2(n12019), .A(n12020), .ZN(n11888) );
  NAND2_X2 U7434 ( .A1(n11932), .A2(n7087), .ZN(n12023) );
  OR2_X1 U7435 ( .A1(n8615), .A2(n6439), .ZN(n8639) );
  NOR2_X4 U7436 ( .A1(n10931), .A2(n6711), .ZN(n11049) );
  NOR2_X2 U7437 ( .A1(n10932), .A2(n10933), .ZN(n10931) );
  XNOR2_X2 U7438 ( .A(n6987), .B(n6986), .ZN(n9031) );
  NAND2_X1 U7439 ( .A1(n14004), .A2(n7154), .ZN(n13942) );
  NOR2_X4 U7440 ( .A1(n14035), .A2(n14268), .ZN(n14004) );
  AOI21_X2 U7441 ( .B1(n12836), .B2(n11564), .A(n12835), .ZN(n12827) );
  NAND2_X1 U7442 ( .A1(n12514), .A2(n11946), .ZN(n6831) );
  NAND2_X1 U7443 ( .A1(n6834), .A2(n7230), .ZN(n12553) );
  AOI21_X1 U7444 ( .B1(n6447), .B2(n12580), .A(n6588), .ZN(n7230) );
  NAND2_X1 U7445 ( .A1(n12579), .A2(n6447), .ZN(n6834) );
  INV_X1 U7446 ( .A(n12244), .ZN(n12260) );
  INV_X1 U7447 ( .A(n7545), .ZN(n6837) );
  NAND2_X1 U7448 ( .A1(n12863), .A2(n11583), .ZN(n11585) );
  INV_X1 U7449 ( .A(n11688), .ZN(n7024) );
  INV_X1 U7450 ( .A(n9148), .ZN(n9150) );
  OAI21_X1 U7451 ( .B1(n8297), .B2(n7619), .A(n7614), .ZN(n8349) );
  NOR2_X1 U7452 ( .A1(n7623), .A2(n7620), .ZN(n7619) );
  AND2_X1 U7453 ( .A1(n7617), .A2(n7615), .ZN(n7614) );
  NAND2_X1 U7454 ( .A1(n7623), .A2(n7618), .ZN(n7617) );
  NAND3_X1 U7455 ( .A1(n9135), .A2(n7428), .A3(n7429), .ZN(n7427) );
  INV_X1 U7456 ( .A(n8113), .ZN(n8115) );
  XNOR2_X1 U7457 ( .A(n7688), .B(SI_15_), .ZN(n8069) );
  NOR2_X1 U7458 ( .A1(n6877), .A2(n11876), .ZN(n11130) );
  NAND2_X1 U7459 ( .A1(n6879), .A2(n6878), .ZN(n6877) );
  AND3_X1 U7460 ( .A1(n8634), .A2(n8633), .A3(n8632), .ZN(n12222) );
  NAND2_X1 U7462 ( .A1(n9038), .A2(n12260), .ZN(n12646) );
  NAND2_X1 U7463 ( .A1(n10210), .A2(n12260), .ZN(n12642) );
  NAND2_X1 U7464 ( .A1(n9120), .A2(n12089), .ZN(n15149) );
  CLKBUF_X1 U7465 ( .A(n8653), .Z(n6883) );
  NAND2_X1 U7466 ( .A1(n7572), .A2(n8897), .ZN(n9079) );
  NAND2_X1 U7467 ( .A1(n8415), .A2(n7649), .ZN(n8369) );
  AOI21_X1 U7468 ( .B1(n7348), .B2(n11723), .A(n6537), .ZN(n7347) );
  AND2_X1 U7469 ( .A1(n13266), .A2(n12895), .ZN(n7032) );
  OAI211_X1 U7470 ( .C1(n10010), .C2(n7773), .A(n8427), .B(n6445), .ZN(n7775)
         );
  INV_X1 U7471 ( .A(n7810), .ZN(n6767) );
  NOR2_X1 U7472 ( .A1(n7987), .A2(n6533), .ZN(n7532) );
  INV_X1 U7473 ( .A(n8085), .ZN(n7049) );
  AOI21_X1 U7474 ( .B1(n8180), .B2(n7520), .A(n8178), .ZN(n7517) );
  OR2_X1 U7475 ( .A1(n13237), .A2(n12986), .ZN(n6913) );
  NAND2_X1 U7476 ( .A1(n7596), .A2(n7594), .ZN(n8276) );
  AOI21_X1 U7477 ( .B1(n7598), .B2(n7600), .A(n7595), .ZN(n7594) );
  INV_X1 U7478 ( .A(n8257), .ZN(n7595) );
  NAND2_X1 U7479 ( .A1(n9119), .A2(n10194), .ZN(n7260) );
  XNOR2_X1 U7480 ( .A(n15174), .B(n11622), .ZN(n10989) );
  AND2_X1 U7481 ( .A1(n6661), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n6657) );
  OR2_X1 U7482 ( .A1(n12659), .A2(n12472), .ZN(n12255) );
  AOI21_X1 U7483 ( .B1(n6828), .B2(n6826), .A(n12499), .ZN(n6824) );
  INV_X1 U7484 ( .A(n6826), .ZN(n6825) );
  OR2_X1 U7485 ( .A1(n12680), .A2(n12533), .ZN(n12110) );
  OR2_X1 U7486 ( .A1(n12690), .A2(n12556), .ZN(n12229) );
  NAND2_X1 U7487 ( .A1(n12545), .A2(n7239), .ZN(n7235) );
  OR2_X1 U7488 ( .A1(n12040), .A2(n11976), .ZN(n12206) );
  OR2_X1 U7489 ( .A1(n12284), .A2(n11112), .ZN(n12154) );
  XNOR2_X1 U7490 ( .A(n10328), .B(n15131), .ZN(n7210) );
  NAND2_X1 U7491 ( .A1(n8556), .A2(n7116), .ZN(n6670) );
  NOR2_X1 U7492 ( .A1(n6682), .A2(n6680), .ZN(n6679) );
  AND2_X1 U7493 ( .A1(n7111), .A2(n6681), .ZN(n6680) );
  INV_X1 U7494 ( .A(n7110), .ZN(n6682) );
  INV_X1 U7495 ( .A(n8838), .ZN(n6681) );
  OR2_X1 U7496 ( .A1(n8720), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8752) );
  NAND2_X1 U7497 ( .A1(n11721), .A2(n7340), .ZN(n7339) );
  INV_X1 U7498 ( .A(n6475), .ZN(n7022) );
  NOR2_X1 U7499 ( .A1(n13290), .A2(n13298), .ZN(n6949) );
  OAI211_X1 U7500 ( .C1(n13389), .C2(n7468), .A(n7466), .B(n10527), .ZN(n7460)
         );
  NAND2_X1 U7501 ( .A1(n7470), .A2(n7467), .ZN(n7466) );
  NAND2_X1 U7502 ( .A1(n7463), .A2(n7462), .ZN(n7461) );
  INV_X1 U7503 ( .A(n10297), .ZN(n7462) );
  INV_X1 U7504 ( .A(n10296), .ZN(n7463) );
  INV_X1 U7505 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9130) );
  NOR2_X1 U7506 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n9132) );
  NOR2_X1 U7507 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n9131) );
  NOR2_X1 U7508 ( .A1(n14290), .A2(n13781), .ZN(n7448) );
  NOR2_X1 U7509 ( .A1(n9377), .A2(n6969), .ZN(n6968) );
  INV_X1 U7510 ( .A(n9366), .ZN(n6969) );
  OR2_X1 U7511 ( .A1(n14248), .A2(n11752), .ZN(n13653) );
  NAND2_X1 U7512 ( .A1(n8319), .A2(n8318), .ZN(n8373) );
  INV_X1 U7513 ( .A(n8320), .ZN(n8318) );
  INV_X1 U7514 ( .A(n9134), .ZN(n7429) );
  INV_X1 U7515 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9382) );
  XNOR2_X1 U7516 ( .A(n8185), .B(SI_20_), .ZN(n7575) );
  NAND2_X1 U7517 ( .A1(n8135), .A2(n6581), .ZN(n7586) );
  INV_X1 U7518 ( .A(n7427), .ZN(n7426) );
  NAND2_X1 U7519 ( .A1(n9382), .A2(n7381), .ZN(n7380) );
  AND2_X1 U7520 ( .A1(n7136), .A2(n7691), .ZN(n7134) );
  XNOR2_X1 U7521 ( .A(n7683), .B(SI_13_), .ZN(n8027) );
  NAND2_X1 U7522 ( .A1(n6807), .A2(n6806), .ZN(n7827) );
  OAI21_X1 U7523 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n14348), .A(n14347), .ZN(
        n14362) );
  NAND2_X1 U7524 ( .A1(n7084), .A2(n6512), .ZN(n11666) );
  AOI21_X1 U7525 ( .B1(n7272), .B2(n7274), .A(n6540), .ZN(n7270) );
  NAND2_X1 U7526 ( .A1(n12012), .A2(n6506), .ZN(n11922) );
  INV_X1 U7527 ( .A(n11640), .ZN(n7275) );
  INV_X1 U7528 ( .A(n12521), .ZN(n11946) );
  INV_X1 U7529 ( .A(n12002), .ZN(n6870) );
  INV_X1 U7530 ( .A(n12060), .ZN(n7265) );
  XNOR2_X1 U7531 ( .A(n7119), .B(n12428), .ZN(n12109) );
  NAND2_X1 U7532 ( .A1(n12265), .A2(n7120), .ZN(n7119) );
  NOR2_X1 U7533 ( .A1(n12262), .A2(n12107), .ZN(n7120) );
  OR2_X1 U7534 ( .A1(n15054), .A2(n8730), .ZN(n6665) );
  NAND2_X1 U7535 ( .A1(n7165), .A2(n7164), .ZN(n15093) );
  INV_X1 U7536 ( .A(n15096), .ZN(n7164) );
  OR2_X1 U7537 ( .A1(n14485), .A2(n12352), .ZN(n7162) );
  INV_X1 U7538 ( .A(n6931), .ZN(n12351) );
  AND2_X1 U7539 ( .A1(n8975), .A2(n8974), .ZN(n12484) );
  NAND2_X1 U7540 ( .A1(n12519), .A2(n6827), .ZN(n6823) );
  NAND2_X1 U7541 ( .A1(n6822), .A2(n6824), .ZN(n12492) );
  OR2_X1 U7542 ( .A1(n12519), .A2(n6825), .ZN(n6822) );
  NAND2_X1 U7543 ( .A1(n12535), .A2(n7005), .ZN(n7541) );
  NOR2_X1 U7544 ( .A1(n12090), .A2(n7006), .ZN(n7005) );
  INV_X1 U7545 ( .A(n12234), .ZN(n7006) );
  OR2_X1 U7546 ( .A1(n12690), .A2(n12276), .ZN(n7238) );
  INV_X1 U7547 ( .A(n12218), .ZN(n7556) );
  NAND2_X1 U7548 ( .A1(n12585), .A2(n12206), .ZN(n12571) );
  AOI21_X1 U7549 ( .B1(n7002), .B2(n7004), .A(n7001), .ZN(n7000) );
  INV_X1 U7550 ( .A(n7003), .ZN(n7002) );
  OAI21_X1 U7551 ( .B1(n11334), .B2(n6590), .A(n8812), .ZN(n11385) );
  INV_X1 U7552 ( .A(n11436), .ZN(n14529) );
  AND2_X1 U7553 ( .A1(n10186), .A2(n9713), .ZN(n10392) );
  AOI21_X1 U7554 ( .B1(n8622), .B2(n7116), .A(n7115), .ZN(n7114) );
  INV_X1 U7555 ( .A(n8562), .ZN(n7115) );
  OAI211_X1 U7556 ( .C1(n8557), .C2(n6668), .A(n6667), .B(n8940), .ZN(n8943)
         );
  INV_X1 U7557 ( .A(n7114), .ZN(n6668) );
  NAND2_X1 U7558 ( .A1(n6670), .A2(n7114), .ZN(n6667) );
  INV_X1 U7559 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n6836) );
  NAND2_X1 U7560 ( .A1(n8557), .A2(n8556), .ZN(n8623) );
  AND2_X1 U7561 ( .A1(n6562), .A2(n7066), .ZN(n7065) );
  NAND2_X1 U7562 ( .A1(n11551), .A2(n11550), .ZN(n6704) );
  NOR2_X1 U7563 ( .A1(n8476), .A2(n11725), .ZN(n8478) );
  AND2_X1 U7564 ( .A1(n7510), .A2(n6568), .ZN(n7040) );
  NOR2_X1 U7565 ( .A1(n8310), .A2(n8309), .ZN(n8370) );
  NOR2_X1 U7566 ( .A1(n8272), .A2(n8271), .ZN(n6786) );
  INV_X1 U7567 ( .A(n7762), .ZN(n8504) );
  INV_X1 U7568 ( .A(n8450), .ZN(n7508) );
  INV_X1 U7569 ( .A(n8444), .ZN(n7509) );
  OAI21_X1 U7570 ( .B1(n14845), .B2(n10013), .A(n6715), .ZN(n14841) );
  NAND2_X1 U7571 ( .A1(n14845), .A2(n10013), .ZN(n6715) );
  NAND2_X1 U7572 ( .A1(n13003), .A2(n13011), .ZN(n7288) );
  NOR2_X1 U7573 ( .A1(n7290), .A2(n6457), .ZN(n7286) );
  OR2_X1 U7574 ( .A1(n7287), .A2(n6457), .ZN(n7285) );
  AOI21_X1 U7575 ( .B1(n7289), .B2(n6454), .A(n7351), .ZN(n7287) );
  AOI21_X1 U7576 ( .B1(n7298), .B2(n7300), .A(n13040), .ZN(n7297) );
  NAND2_X1 U7577 ( .A1(n13073), .A2(n11695), .ZN(n7302) );
  INV_X1 U7578 ( .A(n13139), .ZN(n13225) );
  INV_X1 U7579 ( .A(n10160), .ZN(n6926) );
  OR2_X1 U7580 ( .A1(n9648), .A2(n7904), .ZN(n7805) );
  NAND2_X1 U7581 ( .A1(n7731), .A2(n7730), .ZN(n7736) );
  NOR2_X1 U7582 ( .A1(n7841), .A2(n7725), .ZN(n7730) );
  INV_X1 U7583 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7723) );
  INV_X1 U7584 ( .A(n6983), .ZN(n6982) );
  OAI21_X1 U7585 ( .B1(n6985), .B2(n13485), .A(n6984), .ZN(n6983) );
  NAND2_X1 U7586 ( .A1(n13376), .A2(n6456), .ZN(n6984) );
  INV_X1 U7587 ( .A(n7484), .ZN(n7483) );
  OAI21_X1 U7588 ( .B1(n13485), .B2(n6456), .A(n13376), .ZN(n7484) );
  NAND2_X1 U7589 ( .A1(n11476), .A2(n7489), .ZN(n7488) );
  AND4_X1 U7590 ( .A1(n9310), .A2(n9309), .A3(n9308), .A4(n9307), .ZN(n11486)
         );
  NAND2_X1 U7591 ( .A1(n7451), .A2(n7450), .ZN(n7449) );
  INV_X1 U7592 ( .A(n14106), .ZN(n7451) );
  INV_X1 U7593 ( .A(n9577), .ZN(n9140) );
  AND2_X1 U7594 ( .A1(n9578), .A2(n9154), .ZN(n7454) );
  XNOR2_X1 U7595 ( .A(n9589), .B(n9588), .ZN(n9800) );
  INV_X1 U7596 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9588) );
  NAND2_X1 U7597 ( .A1(n7626), .A2(n7687), .ZN(n8070) );
  INV_X1 U7598 ( .A(n7033), .ZN(n7900) );
  OAI21_X1 U7599 ( .B1(SI_7_), .B2(n7034), .A(n7668), .ZN(n7033) );
  AOI21_X1 U7600 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n14344), .A(n14343), .ZN(
        n14364) );
  AND2_X1 U7601 ( .A1(n7328), .A2(n7327), .ZN(n14405) );
  OAI21_X1 U7602 ( .B1(n7330), .B2(n7329), .A(P2_ADDR_REG_11__SCAN_IN), .ZN(
        n7328) );
  XNOR2_X1 U7603 ( .A(n11648), .B(n11646), .ZN(n11895) );
  NAND2_X1 U7604 ( .A1(n12475), .A2(n6882), .ZN(n12665) );
  OR2_X1 U7605 ( .A1(n12664), .A2(n15153), .ZN(n6882) );
  NAND2_X1 U7606 ( .A1(n8916), .A2(n8915), .ZN(n12756) );
  NAND2_X1 U7607 ( .A1(n8284), .A2(n8283), .ZN(n13259) );
  NAND2_X1 U7608 ( .A1(n8362), .A2(n8361), .ZN(n13027) );
  NAND2_X1 U7609 ( .A1(n8292), .A2(n8291), .ZN(n13012) );
  NAND2_X1 U7610 ( .A1(n8305), .A2(n8304), .ZN(n13060) );
  NAND2_X1 U7611 ( .A1(n9574), .A2(n7471), .ZN(n9971) );
  NOR2_X1 U7612 ( .A1(n14310), .A2(n6976), .ZN(n7471) );
  NAND2_X1 U7613 ( .A1(n6451), .A2(n9585), .ZN(n6976) );
  NAND2_X1 U7614 ( .A1(n9486), .A2(n9485), .ZN(n14165) );
  NOR2_X1 U7615 ( .A1(n14432), .A2(n14893), .ZN(n14431) );
  OR2_X1 U7616 ( .A1(n13587), .A2(n13586), .ZN(n13588) );
  NAND2_X1 U7617 ( .A1(n7371), .A2(n13592), .ZN(n7370) );
  OAI211_X1 U7618 ( .C1(n7814), .C2(n7813), .A(n6765), .B(n6762), .ZN(n7834)
         );
  INV_X1 U7619 ( .A(n13617), .ZN(n7374) );
  INV_X1 U7620 ( .A(n13627), .ZN(n7364) );
  OR2_X1 U7621 ( .A1(n7944), .A2(n7943), .ZN(n7964) );
  AOI21_X1 U7622 ( .B1(n7942), .B2(n7941), .A(n7940), .ZN(n7944) );
  INV_X1 U7623 ( .A(n6549), .ZN(n7538) );
  INV_X1 U7624 ( .A(n8025), .ZN(n7536) );
  INV_X1 U7625 ( .A(n7527), .ZN(n7526) );
  OR2_X1 U7626 ( .A1(n7532), .A2(n7530), .ZN(n7529) );
  OAI21_X1 U7627 ( .B1(n7531), .B2(n7530), .A(n7528), .ZN(n7527) );
  NOR2_X1 U7628 ( .A1(n7042), .A2(n8004), .ZN(n7041) );
  INV_X1 U7629 ( .A(n7531), .ZN(n7042) );
  NOR2_X1 U7630 ( .A1(n7048), .A2(n7047), .ZN(n7046) );
  NOR2_X1 U7631 ( .A1(n7533), .A2(n8067), .ZN(n7047) );
  NOR2_X1 U7632 ( .A1(n6478), .A2(n7049), .ZN(n7048) );
  INV_X1 U7633 ( .A(n8065), .ZN(n7533) );
  OAI21_X1 U7634 ( .B1(n6799), .B2(n7360), .A(n6924), .ZN(n6798) );
  AND2_X1 U7635 ( .A1(n7359), .A2(n13701), .ZN(n6924) );
  NAND2_X1 U7636 ( .A1(n7358), .A2(n13700), .ZN(n7357) );
  AND2_X1 U7637 ( .A1(n8159), .A2(n6462), .ZN(n7521) );
  NAND2_X1 U7638 ( .A1(n7035), .A2(n6785), .ZN(n6784) );
  NAND2_X1 U7639 ( .A1(n8132), .A2(n8131), .ZN(n6785) );
  INV_X1 U7640 ( .A(n7521), .ZN(n7518) );
  NOR2_X1 U7641 ( .A1(n12239), .A2(n12493), .ZN(n6702) );
  NOR2_X1 U7642 ( .A1(n8202), .A2(n8205), .ZN(n7512) );
  INV_X1 U7643 ( .A(n8202), .ZN(n7511) );
  NAND2_X1 U7644 ( .A1(n10250), .A2(n7762), .ZN(n8245) );
  AND2_X1 U7645 ( .A1(n13714), .A2(n6818), .ZN(n6817) );
  INV_X1 U7646 ( .A(n13713), .ZN(n6818) );
  INV_X1 U7647 ( .A(n8210), .ZN(n7600) );
  INV_X1 U7648 ( .A(n11652), .ZN(n7086) );
  INV_X1 U7649 ( .A(n6997), .ZN(n6996) );
  OAI21_X1 U7650 ( .B1(n12092), .B2(n6998), .A(n12156), .ZN(n6997) );
  INV_X1 U7651 ( .A(n12154), .ZN(n6998) );
  NAND2_X1 U7652 ( .A1(n10395), .A2(n6461), .ZN(n7076) );
  INV_X1 U7653 ( .A(n8553), .ZN(n6692) );
  OAI21_X1 U7654 ( .B1(n8552), .B2(n6692), .A(n8910), .ZN(n6691) );
  NAND2_X1 U7655 ( .A1(n13551), .A2(n13548), .ZN(n13725) );
  INV_X1 U7656 ( .A(n13722), .ZN(n7368) );
  NOR2_X1 U7657 ( .A1(n14171), .A2(n14165), .ZN(n7157) );
  NOR2_X1 U7658 ( .A1(n7409), .A2(n7406), .ZN(n7405) );
  INV_X1 U7659 ( .A(n9540), .ZN(n7408) );
  INV_X1 U7660 ( .A(n8349), .ZN(n6876) );
  NAND2_X1 U7661 ( .A1(n6814), .A2(n6815), .ZN(n8185) );
  AOI21_X1 U7662 ( .B1(n6450), .B2(n7588), .A(n6816), .ZN(n6815) );
  NAND2_X1 U7663 ( .A1(n8113), .A2(n6450), .ZN(n6814) );
  INV_X1 U7664 ( .A(n8160), .ZN(n6816) );
  INV_X1 U7665 ( .A(n8114), .ZN(n8116) );
  OR2_X1 U7666 ( .A1(n9257), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n9288) );
  NAND2_X1 U7667 ( .A1(n7072), .A2(SI_5_), .ZN(n7665) );
  AND2_X1 U7668 ( .A1(n12049), .A2(n7273), .ZN(n7272) );
  OR2_X1 U7669 ( .A1(n11944), .A2(n7274), .ZN(n7273) );
  NAND2_X1 U7670 ( .A1(n11951), .A2(n12066), .ZN(n7252) );
  XNOR2_X1 U7671 ( .A(n11622), .B(n11963), .ZN(n10992) );
  OR2_X1 U7672 ( .A1(n12724), .A2(n12450), .ZN(n12263) );
  NAND2_X1 U7673 ( .A1(n7090), .A2(n7089), .ZN(n6888) );
  NAND2_X1 U7674 ( .A1(n11081), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7089) );
  NOR2_X1 U7675 ( .A1(n11411), .A2(n15071), .ZN(n11412) );
  AND2_X1 U7676 ( .A1(n15093), .A2(n12321), .ZN(n12328) );
  INV_X1 U7677 ( .A(n12368), .ZN(n7109) );
  NAND2_X1 U7678 ( .A1(n12350), .A2(n12357), .ZN(n6931) );
  OR2_X1 U7679 ( .A1(n8931), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8946) );
  AND2_X1 U7680 ( .A1(n6497), .A2(n8740), .ZN(n7228) );
  INV_X1 U7681 ( .A(n8527), .ZN(n6686) );
  INV_X1 U7682 ( .A(n6664), .ZN(n8718) );
  OR2_X1 U7683 ( .A1(n8687), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n6664) );
  INV_X1 U7684 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7651) );
  NAND2_X1 U7685 ( .A1(n13237), .A2(n8427), .ZN(n6912) );
  AOI21_X1 U7686 ( .B1(n7335), .B2(n7336), .A(n6518), .ZN(n6758) );
  INV_X1 U7687 ( .A(n7337), .ZN(n7336) );
  OR2_X1 U7688 ( .A1(n13280), .A2(n12861), .ZN(n11693) );
  NOR2_X1 U7689 ( .A1(n13123), .A2(n7023), .ZN(n7015) );
  NOR2_X1 U7690 ( .A1(n13174), .A2(n13302), .ZN(n11731) );
  INV_X1 U7691 ( .A(n11362), .ZN(n7312) );
  NOR2_X1 U7692 ( .A1(n10903), .A2(n15027), .ZN(n7168) );
  AOI21_X1 U7693 ( .B1(n10877), .B2(n7295), .A(n7294), .ZN(n7293) );
  INV_X1 U7694 ( .A(n10878), .ZN(n7295) );
  NAND3_X1 U7695 ( .A1(n13064), .A2(n13003), .A3(n6455), .ZN(n13005) );
  NAND2_X1 U7696 ( .A1(n13190), .A2(n13172), .ZN(n13174) );
  NOR2_X1 U7697 ( .A1(n13206), .A2(n13189), .ZN(n13190) );
  AND2_X1 U7698 ( .A1(n11222), .A2(n7762), .ZN(n7770) );
  INV_X1 U7699 ( .A(n10745), .ZN(n7492) );
  XNOR2_X1 U7700 ( .A(n6731), .B(n11838), .ZN(n10295) );
  NAND2_X1 U7701 ( .A1(n10289), .A2(n6732), .ZN(n6731) );
  NAND2_X1 U7702 ( .A1(n13797), .A2(n11827), .ZN(n6732) );
  INV_X1 U7703 ( .A(n11806), .ZN(n7476) );
  NAND2_X1 U7704 ( .A1(n7591), .A2(n7589), .ZN(n7593) );
  NOR2_X1 U7705 ( .A1(n13734), .A2(n7590), .ZN(n7589) );
  INV_X1 U7706 ( .A(n13502), .ZN(n7590) );
  INV_X1 U7707 ( .A(n13548), .ZN(n9566) );
  OR2_X1 U7708 ( .A1(n13505), .A2(n9810), .ZN(n7402) );
  NAND2_X1 U7709 ( .A1(n6958), .A2(n9473), .ZN(n6957) );
  INV_X1 U7710 ( .A(n6960), .ZN(n6958) );
  INV_X1 U7711 ( .A(n9473), .ZN(n6959) );
  INV_X1 U7712 ( .A(n7189), .ZN(n7188) );
  OAI21_X1 U7713 ( .B1(n13998), .B2(n7190), .A(n13980), .ZN(n7189) );
  INV_X1 U7714 ( .A(n13981), .ZN(n7190) );
  NOR2_X1 U7715 ( .A1(n14014), .A2(n6961), .ZN(n6960) );
  INV_X1 U7716 ( .A(n9460), .ZN(n6961) );
  NAND2_X1 U7717 ( .A1(n7129), .A2(n14054), .ZN(n7132) );
  NAND2_X1 U7718 ( .A1(n7199), .A2(n14054), .ZN(n7133) );
  NAND2_X1 U7719 ( .A1(n7203), .A2(n13539), .ZN(n7202) );
  NAND2_X1 U7720 ( .A1(n7204), .A2(n7206), .ZN(n7203) );
  XNOR2_X1 U7721 ( .A(n14281), .B(n7138), .ZN(n13539) );
  INV_X1 U7722 ( .A(n9535), .ZN(n7437) );
  NOR2_X1 U7723 ( .A1(n9220), .A2(n7194), .ZN(n7193) );
  INV_X1 U7724 ( .A(n9206), .ZN(n7194) );
  NAND2_X1 U7725 ( .A1(n6482), .A2(n9531), .ZN(n7433) );
  AND2_X1 U7726 ( .A1(n13519), .A2(n9530), .ZN(n7434) );
  INV_X1 U7727 ( .A(n13564), .ZN(n9970) );
  OR2_X1 U7728 ( .A1(n14729), .A2(n14725), .ZN(n13565) );
  AOI21_X1 U7729 ( .B1(n13644), .B2(n6955), .A(n6954), .ZN(n6953) );
  INV_X1 U7730 ( .A(n9327), .ZN(n6955) );
  INV_X1 U7731 ( .A(n13647), .ZN(n6954) );
  INV_X1 U7732 ( .A(n13644), .ZN(n6956) );
  INV_X1 U7733 ( .A(n7605), .ZN(n7604) );
  OAI21_X1 U7734 ( .B1(n8275), .B2(n8274), .A(n8277), .ZN(n8297) );
  XNOR2_X1 U7735 ( .A(n8276), .B(SI_24_), .ZN(n8275) );
  INV_X1 U7736 ( .A(n7127), .ZN(n7126) );
  OAI21_X1 U7737 ( .B1(n7612), .B2(n6452), .A(n8006), .ZN(n7127) );
  INV_X1 U7738 ( .A(SI_12_), .ZN(n7679) );
  OAI21_X1 U7739 ( .B1(n7610), .B2(SI_10_), .A(n7125), .ZN(n7124) );
  NAND2_X1 U7740 ( .A1(n7611), .A2(SI_10_), .ZN(n7125) );
  NAND2_X1 U7741 ( .A1(n6809), .A2(n6476), .ZN(n6813) );
  INV_X1 U7742 ( .A(n7675), .ZN(n6809) );
  INV_X1 U7743 ( .A(n7610), .ZN(n7128) );
  INV_X1 U7744 ( .A(n7988), .ZN(n7612) );
  NAND2_X1 U7745 ( .A1(n7858), .A2(n7665), .ZN(n7884) );
  NAND2_X1 U7746 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n6916), .ZN(n6915) );
  INV_X1 U7747 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6916) );
  NAND2_X1 U7748 ( .A1(n14330), .A2(n14331), .ZN(n14332) );
  XNOR2_X1 U7749 ( .A(n14332), .B(n7320), .ZN(n14381) );
  INV_X1 U7750 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7320) );
  AOI21_X2 U7751 ( .B1(n12032), .B2(n11928), .A(n6483), .ZN(n11648) );
  XNOR2_X1 U7752 ( .A(n15131), .B(n11622), .ZN(n10322) );
  INV_X1 U7753 ( .A(n7252), .ZN(n6622) );
  OR2_X1 U7754 ( .A1(n11951), .A2(n12066), .ZN(n11627) );
  OAI21_X1 U7755 ( .B1(n11989), .B2(n7079), .A(n10990), .ZN(n6902) );
  INV_X1 U7756 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11077) );
  NAND2_X1 U7757 ( .A1(n8598), .A2(n8597), .ZN(n8919) );
  INV_X1 U7758 ( .A(n8917), .ZN(n8598) );
  NAND2_X1 U7759 ( .A1(n7255), .A2(n12280), .ZN(n7254) );
  INV_X1 U7760 ( .A(n11431), .ZN(n7255) );
  NAND2_X1 U7761 ( .A1(n10272), .A2(n10271), .ZN(n10273) );
  XNOR2_X1 U7762 ( .A(n10322), .B(n10328), .ZN(n10274) );
  OR2_X1 U7763 ( .A1(n8901), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8917) );
  OR2_X1 U7764 ( .A1(n10992), .A2(n11993), .ZN(n6879) );
  NOR2_X1 U7765 ( .A1(n6990), .A2(n6989), .ZN(n6988) );
  AND2_X1 U7766 ( .A1(n12262), .A2(n12724), .ZN(n6989) );
  AOI21_X1 U7767 ( .B1(n12078), .B2(n12258), .A(n6991), .ZN(n6990) );
  NAND2_X1 U7768 ( .A1(n12265), .A2(n6992), .ZN(n6991) );
  NAND2_X1 U7769 ( .A1(n6640), .A2(n10653), .ZN(n10629) );
  NAND2_X1 U7770 ( .A1(n6642), .A2(n6641), .ZN(n6640) );
  OR2_X1 U7771 ( .A1(n10620), .A2(n6641), .ZN(n7096) );
  INV_X1 U7772 ( .A(n10619), .ZN(n7099) );
  NAND2_X1 U7773 ( .A1(n10620), .A2(n10619), .ZN(n7097) );
  NAND2_X1 U7774 ( .A1(n6665), .A2(n6480), .ZN(n7092) );
  NAND2_X1 U7775 ( .A1(n7092), .A2(n7091), .ZN(n7090) );
  INV_X1 U7776 ( .A(n10958), .ZN(n7091) );
  XNOR2_X1 U7777 ( .A(n7177), .B(n11423), .ZN(n11424) );
  NAND2_X1 U7778 ( .A1(n6654), .A2(n6652), .ZN(n7177) );
  AOI21_X1 U7779 ( .B1(n11421), .B2(n6655), .A(n6653), .ZN(n6652) );
  NAND2_X1 U7780 ( .A1(n11420), .A2(n6655), .ZN(n6654) );
  INV_X1 U7781 ( .A(n11422), .ZN(n6653) );
  NOR2_X1 U7782 ( .A1(n11424), .A2(n11336), .ZN(n12299) );
  OR2_X1 U7783 ( .A1(n15091), .A2(n15090), .ZN(n15088) );
  NOR2_X1 U7784 ( .A1(n11412), .A2(n11413), .ZN(n12308) );
  OR2_X1 U7785 ( .A1(n12318), .A2(n12319), .ZN(n7165) );
  INV_X1 U7786 ( .A(n6930), .ZN(n12317) );
  AND2_X1 U7787 ( .A1(n15088), .A2(n12303), .ZN(n12332) );
  OR2_X1 U7788 ( .A1(n14480), .A2(n12372), .ZN(n7107) );
  NAND2_X1 U7789 ( .A1(n7107), .A2(n7106), .ZN(n12387) );
  INV_X1 U7790 ( .A(n12375), .ZN(n7106) );
  NAND2_X1 U7791 ( .A1(n6659), .A2(n12406), .ZN(n6658) );
  INV_X1 U7792 ( .A(n12387), .ZN(n6659) );
  NAND2_X1 U7793 ( .A1(n12387), .A2(n6660), .ZN(n6656) );
  AND2_X1 U7794 ( .A1(n12417), .A2(n12386), .ZN(n6660) );
  INV_X1 U7795 ( .A(n12355), .ZN(n7161) );
  NAND2_X1 U7796 ( .A1(n7105), .A2(n7104), .ZN(n7103) );
  INV_X1 U7797 ( .A(n12420), .ZN(n7104) );
  OR2_X1 U7798 ( .A1(n8996), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9013) );
  NAND2_X1 U7799 ( .A1(n7247), .A2(n7246), .ZN(n12469) );
  AND2_X1 U7800 ( .A1(n7247), .A2(n7250), .ZN(n12470) );
  AND2_X1 U7801 ( .A1(n8988), .A2(n8987), .ZN(n12497) );
  NAND2_X1 U7802 ( .A1(n6552), .A2(n6831), .ZN(n6826) );
  OR2_X1 U7803 ( .A1(n8946), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8956) );
  AOI21_X1 U7804 ( .B1(n12518), .B2(n7544), .A(n7543), .ZN(n7542) );
  INV_X1 U7805 ( .A(n12110), .ZN(n7543) );
  INV_X1 U7806 ( .A(n12233), .ZN(n7544) );
  NAND2_X1 U7807 ( .A1(n12111), .A2(n12113), .ZN(n12510) );
  OR2_X1 U7808 ( .A1(n12037), .A2(n11928), .ZN(n12233) );
  NAND2_X1 U7809 ( .A1(n12037), .A2(n12543), .ZN(n7237) );
  OAI21_X1 U7810 ( .B1(n9050), .B2(n7009), .A(n7007), .ZN(n9052) );
  AOI21_X1 U7811 ( .B1(n7010), .B2(n7013), .A(n7008), .ZN(n7007) );
  OR2_X1 U7812 ( .A1(n8919), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8631) );
  AOI21_X1 U7813 ( .B1(n7555), .B2(n9051), .A(n7553), .ZN(n7552) );
  INV_X1 U7814 ( .A(n12224), .ZN(n7553) );
  OR2_X1 U7815 ( .A1(n12555), .A2(n7235), .ZN(n12541) );
  AND3_X1 U7816 ( .A1(n8629), .A2(n8628), .A3(n8627), .ZN(n12556) );
  AND4_X1 U7817 ( .A1(n8891), .A2(n8890), .A3(n8889), .A4(n8888), .ZN(n12583)
         );
  NAND2_X1 U7818 ( .A1(n8908), .A2(n8907), .ZN(n12577) );
  INV_X1 U7819 ( .A(n12579), .ZN(n8908) );
  NAND2_X1 U7820 ( .A1(n9050), .A2(n7012), .ZN(n12585) );
  INV_X1 U7821 ( .A(n12594), .ZN(n12599) );
  NAND2_X1 U7822 ( .A1(n6819), .A2(n7222), .ZN(n12609) );
  AOI21_X1 U7823 ( .B1(n12624), .B2(n7223), .A(n6586), .ZN(n7222) );
  NAND2_X1 U7824 ( .A1(n12641), .A2(n7220), .ZN(n6819) );
  INV_X1 U7825 ( .A(n8854), .ZN(n7223) );
  NAND2_X1 U7826 ( .A1(n12639), .A2(n8854), .ZN(n12625) );
  NAND2_X1 U7827 ( .A1(n7559), .A2(n7560), .ZN(n12631) );
  AOI21_X1 U7828 ( .B1(n7562), .B2(n9048), .A(n7561), .ZN(n7560) );
  NAND2_X1 U7829 ( .A1(n12631), .A2(n12630), .ZN(n12629) );
  AND4_X1 U7830 ( .A1(n8867), .A2(n8866), .A3(n8865), .A4(n8864), .ZN(n12647)
         );
  NAND2_X1 U7831 ( .A1(n12641), .A2(n12640), .ZN(n12639) );
  NAND2_X1 U7832 ( .A1(n11229), .A2(n6510), .ZN(n11331) );
  OR2_X1 U7833 ( .A1(n8775), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8796) );
  NAND2_X1 U7834 ( .A1(n11152), .A2(n12170), .ZN(n9046) );
  NAND2_X1 U7835 ( .A1(n9046), .A2(n7567), .ZN(n11229) );
  NOR2_X1 U7836 ( .A1(n12096), .A2(n7568), .ZN(n7567) );
  INV_X1 U7837 ( .A(n12169), .ZN(n7568) );
  OR2_X1 U7838 ( .A1(n8742), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8758) );
  AND3_X1 U7839 ( .A1(n8724), .A2(n8723), .A3(n8722), .ZN(n11112) );
  NAND2_X1 U7840 ( .A1(n8667), .A2(n7210), .ZN(n7208) );
  OR2_X1 U7841 ( .A1(n9010), .A2(n6852), .ZN(n8677) );
  INV_X1 U7842 ( .A(n9624), .ZN(n6852) );
  INV_X1 U7843 ( .A(n12642), .ZN(n15142) );
  OR2_X1 U7844 ( .A1(n14437), .A2(n10441), .ZN(n12244) );
  NAND2_X1 U7845 ( .A1(n8995), .A2(n8994), .ZN(n12659) );
  NAND2_X1 U7846 ( .A1(n8967), .A2(n8966), .ZN(n12240) );
  NOR2_X1 U7847 ( .A1(n9114), .A2(n9104), .ZN(n10208) );
  NOR2_X1 U7848 ( .A1(n9115), .A2(n9104), .ZN(n10212) );
  NAND2_X1 U7849 ( .A1(n14437), .A2(n10441), .ZN(n15138) );
  INV_X1 U7850 ( .A(n15138), .ZN(n15173) );
  INV_X1 U7851 ( .A(n12646), .ZN(n15145) );
  OAI21_X1 U7852 ( .B1(n9005), .B2(n9004), .A(n9006), .ZN(n9008) );
  OAI21_X1 U7853 ( .B1(n8977), .B2(n8570), .A(n8571), .ZN(n8991) );
  INV_X1 U7854 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n6628) );
  AND2_X1 U7855 ( .A1(n8564), .A2(n8563), .ZN(n8940) );
  INV_X1 U7856 ( .A(n6670), .ZN(n6669) );
  AND2_X1 U7857 ( .A1(n7278), .A2(n9025), .ZN(n7277) );
  INV_X1 U7858 ( .A(n8559), .ZN(n7117) );
  NAND2_X1 U7859 ( .A1(n8623), .A2(n8558), .ZN(n7118) );
  AND2_X1 U7860 ( .A1(n8913), .A2(n9029), .ZN(n7278) );
  INV_X1 U7861 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n9029) );
  AOI21_X1 U7862 ( .B1(n8548), .B2(n7112), .A(n6589), .ZN(n7111) );
  INV_X1 U7863 ( .A(n8546), .ZN(n7112) );
  OAI21_X1 U7864 ( .B1(n8785), .B2(n6582), .A(n6697), .ZN(n8814) );
  INV_X1 U7865 ( .A(n6698), .ZN(n6697) );
  OAI21_X1 U7866 ( .B1(n6582), .B2(n8536), .A(n8537), .ZN(n6698) );
  NAND2_X1 U7867 ( .A1(n8698), .A2(n8526), .ZN(n6688) );
  INV_X1 U7868 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n8702) );
  NAND2_X1 U7869 ( .A1(n6664), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8700) );
  NAND2_X1 U7870 ( .A1(n8663), .A2(n8662), .ZN(n8661) );
  INV_X1 U7871 ( .A(n11600), .ZN(n7398) );
  NOR2_X1 U7872 ( .A1(n12777), .A2(n7401), .ZN(n7400) );
  INV_X1 U7873 ( .A(n11604), .ZN(n7401) );
  XNOR2_X1 U7874 ( .A(n11584), .B(n10168), .ZN(n9757) );
  INV_X1 U7875 ( .A(n11585), .ZN(n11587) );
  NAND2_X1 U7876 ( .A1(n7385), .A2(n7387), .ZN(n7384) );
  XNOR2_X1 U7877 ( .A(n11582), .B(n11581), .ZN(n12862) );
  NAND2_X1 U7878 ( .A1(n12813), .A2(n11600), .ZN(n12885) );
  NAND2_X1 U7879 ( .A1(n14868), .A2(n14867), .ZN(n14866) );
  NOR2_X1 U7880 ( .A1(n14916), .A2(n14917), .ZN(n14915) );
  OR2_X1 U7881 ( .A1(n14953), .A2(n14952), .ZN(n6720) );
  NOR2_X1 U7882 ( .A1(n12992), .A2(n12991), .ZN(n12990) );
  AOI21_X1 U7883 ( .B1(n7285), .B2(n7283), .A(n7282), .ZN(n7281) );
  INV_X1 U7884 ( .A(n7286), .ZN(n7283) );
  NAND2_X1 U7885 ( .A1(n6759), .A2(n7344), .ZN(n12996) );
  AOI21_X1 U7886 ( .B1(n7347), .B2(n7345), .A(n12999), .ZN(n7344) );
  NAND2_X1 U7887 ( .A1(n6757), .A2(n6755), .ZN(n6759) );
  INV_X1 U7888 ( .A(n7348), .ZN(n7345) );
  INV_X1 U7889 ( .A(n13035), .ZN(n6904) );
  INV_X1 U7890 ( .A(n11723), .ZN(n6903) );
  OR2_X1 U7891 ( .A1(n13259), .A2(n13012), .ZN(n7352) );
  NOR2_X1 U7892 ( .A1(n13013), .A2(n7349), .ZN(n7348) );
  INV_X1 U7893 ( .A(n7352), .ZN(n7349) );
  OAI21_X1 U7894 ( .B1(n13026), .B2(n6454), .A(n7289), .ZN(n7031) );
  NAND2_X1 U7895 ( .A1(n13064), .A2(n13050), .ZN(n13046) );
  NOR2_X1 U7896 ( .A1(n13076), .A2(n13269), .ZN(n13064) );
  NOR2_X1 U7897 ( .A1(n11694), .A2(n7340), .ZN(n7301) );
  AND2_X1 U7898 ( .A1(n7302), .A2(n7305), .ZN(n13057) );
  NAND2_X1 U7899 ( .A1(n7176), .A2(n7175), .ZN(n13098) );
  NOR2_X1 U7900 ( .A1(n13123), .A2(n7019), .ZN(n7018) );
  NAND2_X1 U7901 ( .A1(n13153), .A2(n7023), .ZN(n7020) );
  INV_X1 U7902 ( .A(n13153), .ZN(n7026) );
  AOI21_X1 U7903 ( .B1(n6751), .B2(n13184), .A(n6749), .ZN(n6748) );
  INV_X1 U7904 ( .A(n6751), .ZN(n6750) );
  INV_X1 U7905 ( .A(n7353), .ZN(n6749) );
  NAND2_X1 U7906 ( .A1(n7753), .A2(n7752), .ZN(n8124) );
  AND2_X1 U7907 ( .A1(n13154), .A2(n11713), .ZN(n7355) );
  NAND2_X1 U7908 ( .A1(n13168), .A2(n13167), .ZN(n7356) );
  NAND2_X1 U7909 ( .A1(n13180), .A2(n11711), .ZN(n13168) );
  AND2_X1 U7910 ( .A1(n11678), .A2(n11675), .ZN(n11363) );
  NAND2_X1 U7911 ( .A1(n11211), .A2(n11210), .ZN(n11356) );
  NAND2_X1 U7912 ( .A1(n11192), .A2(n11191), .ZN(n11215) );
  AOI21_X1 U7913 ( .B1(n10912), .B2(n6754), .A(n6493), .ZN(n6753) );
  INV_X1 U7914 ( .A(n10867), .ZN(n6754) );
  NOR2_X1 U7915 ( .A1(n10342), .A2(n15001), .ZN(n10556) );
  AOI21_X1 U7916 ( .B1(n6550), .B2(n6939), .A(n6745), .ZN(n6744) );
  NOR2_X1 U7917 ( .A1(n10236), .A2(n12913), .ZN(n6745) );
  OR2_X1 U7918 ( .A1(n15030), .A2(n13230), .ZN(n9779) );
  NAND2_X1 U7919 ( .A1(n13355), .A2(n8423), .ZN(n8351) );
  NAND2_X1 U7920 ( .A1(n8030), .A2(n8029), .ZN(n11704) );
  NAND2_X1 U7921 ( .A1(n9629), .A2(n8423), .ZN(n6741) );
  AND2_X1 U7922 ( .A1(n7762), .A2(n11445), .ZN(n9772) );
  NAND2_X1 U7923 ( .A1(n6905), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7707) );
  NAND2_X1 U7924 ( .A1(n7706), .A2(n7522), .ZN(n6905) );
  NAND2_X1 U7925 ( .A1(n6708), .A2(n7788), .ZN(n7841) );
  OR2_X1 U7926 ( .A1(n9672), .A2(n9272), .ZN(n9235) );
  OR2_X1 U7927 ( .A1(n13376), .A2(n6456), .ZN(n6985) );
  NAND2_X1 U7928 ( .A1(n11742), .A2(n6515), .ZN(n15381) );
  AOI21_X1 U7929 ( .B1(n7483), .B2(n6456), .A(n6526), .ZN(n7482) );
  INV_X1 U7930 ( .A(n7460), .ZN(n7456) );
  NAND2_X1 U7931 ( .A1(n7464), .A2(n7461), .ZN(n10526) );
  INV_X1 U7932 ( .A(n14559), .ZN(n6733) );
  NAND2_X1 U7933 ( .A1(n7488), .A2(n6513), .ZN(n7486) );
  OAI21_X1 U7934 ( .B1(n13456), .B2(n7499), .A(n6729), .ZN(n13464) );
  AOI21_X1 U7935 ( .B1(n7498), .B2(n6730), .A(n6584), .ZN(n6729) );
  INV_X1 U7936 ( .A(n13455), .ZN(n6730) );
  NAND2_X1 U7937 ( .A1(n13464), .A2(n13465), .ZN(n13463) );
  OR2_X1 U7938 ( .A1(n11465), .A2(n11464), .ZN(n6972) );
  NAND2_X1 U7939 ( .A1(n13474), .A2(n13475), .ZN(n13473) );
  AND2_X1 U7940 ( .A1(n10546), .A2(n7461), .ZN(n7459) );
  NAND2_X1 U7941 ( .A1(n11826), .A2(n10641), .ZN(n11836) );
  AND4_X1 U7942 ( .A1(n9483), .A2(n9482), .A3(n9481), .A4(n9480), .ZN(n13419)
         );
  AND4_X1 U7943 ( .A1(n9365), .A2(n9364), .A3(n9363), .A4(n9362), .ZN(n13656)
         );
  AND4_X1 U7944 ( .A1(n9326), .A2(n9325), .A3(n9324), .A4(n9323), .ZN(n13636)
         );
  INV_X1 U7945 ( .A(n13506), .ZN(n9419) );
  AND4_X1 U7946 ( .A1(n9242), .A2(n9241), .A3(n9240), .A4(n9239), .ZN(n10791)
         );
  AND4_X1 U7947 ( .A1(n9230), .A2(n9229), .A3(n9228), .A4(n9227), .ZN(n13593)
         );
  NOR2_X1 U7948 ( .A1(n13942), .A2(n14155), .ZN(n13944) );
  OAI21_X1 U7949 ( .B1(n13997), .B2(n7190), .A(n7188), .ZN(n7142) );
  NAND2_X1 U7950 ( .A1(n14017), .A2(n9473), .ZN(n13997) );
  NAND2_X1 U7951 ( .A1(n14027), .A2(n6960), .ZN(n14017) );
  AND2_X1 U7952 ( .A1(n14014), .A2(n9549), .ZN(n7410) );
  NAND3_X1 U7953 ( .A1(n7133), .A2(n7132), .A3(n7130), .ZN(n14027) );
  NOR2_X1 U7954 ( .A1(n14024), .A2(n7131), .ZN(n7130) );
  INV_X1 U7955 ( .A(n9446), .ZN(n7131) );
  NAND2_X1 U7956 ( .A1(n7159), .A2(n7158), .ZN(n14035) );
  INV_X1 U7957 ( .A(n14272), .ZN(n7158) );
  INV_X1 U7958 ( .A(n13539), .ZN(n14061) );
  NOR2_X1 U7959 ( .A1(n14094), .A2(n14285), .ZN(n14077) );
  AOI21_X1 U7960 ( .B1(n7447), .B2(n14105), .A(n6477), .ZN(n7444) );
  INV_X1 U7961 ( .A(n7448), .ZN(n7446) );
  OR2_X1 U7962 ( .A1(n14110), .A2(n14215), .ZN(n14094) );
  AND2_X1 U7963 ( .A1(n14109), .A2(n13680), .ZN(n14091) );
  NAND2_X1 U7964 ( .A1(n14091), .A2(n14098), .ZN(n14090) );
  AOI21_X1 U7965 ( .B1(n7419), .B2(n7421), .A(n7417), .ZN(n7416) );
  AND2_X1 U7966 ( .A1(n14142), .A2(n14132), .ZN(n14127) );
  NAND2_X1 U7967 ( .A1(n14127), .A2(n14113), .ZN(n14110) );
  OR2_X1 U7968 ( .A1(n14107), .A2(n7450), .ZN(n14109) );
  NAND2_X1 U7969 ( .A1(n6967), .A2(n6964), .ZN(n14123) );
  NOR2_X1 U7970 ( .A1(n6965), .A2(n6509), .ZN(n6964) );
  NAND2_X1 U7971 ( .A1(n11533), .A2(n13535), .ZN(n11532) );
  OR2_X1 U7972 ( .A1(n11531), .A2(n13535), .ZN(n11529) );
  INV_X1 U7973 ( .A(n14248), .ZN(n11753) );
  NAND2_X1 U7974 ( .A1(n11517), .A2(n11753), .ZN(n11534) );
  OR2_X1 U7975 ( .A1(n11499), .A2(n13644), .ZN(n11501) );
  AND2_X1 U7976 ( .A1(n13647), .A2(n13645), .ZN(n13644) );
  NAND2_X1 U7977 ( .A1(n11317), .A2(n9311), .ZN(n14449) );
  NAND2_X1 U7978 ( .A1(n11062), .A2(n9284), .ZN(n11342) );
  NAND2_X1 U7979 ( .A1(n11341), .A2(n13530), .ZN(n11340) );
  NAND2_X1 U7980 ( .A1(n9261), .A2(n9260), .ZN(n14693) );
  NAND2_X1 U7981 ( .A1(n10789), .A2(n6970), .ZN(n14684) );
  AND2_X1 U7982 ( .A1(n13527), .A2(n9256), .ZN(n6970) );
  INV_X1 U7983 ( .A(n13603), .ZN(n10765) );
  AND2_X1 U7984 ( .A1(n9201), .A2(n6573), .ZN(n7375) );
  INV_X1 U7985 ( .A(n7380), .ZN(n7379) );
  NAND2_X1 U7986 ( .A1(n7196), .A2(n7195), .ZN(n10492) );
  INV_X1 U7987 ( .A(n10489), .ZN(n7196) );
  NAND2_X1 U7988 ( .A1(n10221), .A2(n7434), .ZN(n10504) );
  XNOR2_X1 U7989 ( .A(n13797), .B(n13578), .ZN(n10222) );
  AND2_X1 U7990 ( .A1(n13573), .A2(n13572), .ZN(n13569) );
  NAND2_X1 U7991 ( .A1(n9386), .A2(n9385), .ZN(n14230) );
  INV_X1 U7992 ( .A(n13594), .ZN(n14779) );
  INV_X1 U7993 ( .A(n14796), .ZN(n14758) );
  AND2_X1 U7994 ( .A1(n9583), .A2(n9582), .ZN(n9702) );
  XNOR2_X1 U7995 ( .A(n8422), .B(n8421), .ZN(n13512) );
  XNOR2_X1 U7996 ( .A(n6971), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9149) );
  OR2_X1 U7997 ( .A1(n9144), .A2(n9156), .ZN(n6971) );
  OAI21_X1 U7998 ( .B1(n9153), .B2(P1_IR_REG_27__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6613) );
  AND3_X1 U7999 ( .A1(n7428), .A2(n9135), .A3(n9575), .ZN(n7425) );
  INV_X1 U8000 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9578) );
  INV_X1 U8001 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9575) );
  NAND2_X1 U8002 ( .A1(n9201), .A2(n6481), .ZN(n7424) );
  AND2_X1 U8003 ( .A1(n9382), .A2(n7378), .ZN(n7501) );
  INV_X1 U8004 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7502) );
  NAND2_X1 U8005 ( .A1(n7585), .A2(n6450), .ZN(n8161) );
  NAND2_X1 U8006 ( .A1(n7585), .A2(n7586), .ZN(n8141) );
  AND2_X1 U8007 ( .A1(n9201), .A2(n7381), .ZN(n7376) );
  NAND2_X1 U8008 ( .A1(n7135), .A2(n7627), .ZN(n8087) );
  NAND2_X1 U8009 ( .A1(n7884), .A2(n7883), .ZN(n7886) );
  AND2_X1 U8010 ( .A1(n7900), .A2(n7056), .ZN(n7055) );
  NAND2_X1 U8011 ( .A1(n7666), .A2(n7667), .ZN(n7056) );
  INV_X1 U8012 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9190) );
  XNOR2_X1 U8013 ( .A(n14368), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n14369) );
  XNOR2_X1 U8014 ( .A(n14381), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n14383) );
  INV_X1 U8015 ( .A(n14595), .ZN(n7329) );
  OAI21_X1 U8016 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n14346), .A(n14345), .ZN(
        n14402) );
  NAND2_X1 U8017 ( .A1(n6768), .A2(n6774), .ZN(n6772) );
  INV_X1 U8018 ( .A(n14608), .ZN(n6773) );
  INV_X1 U8019 ( .A(n14612), .ZN(n6771) );
  NAND2_X1 U8020 ( .A1(n9099), .A2(n9098), .ZN(n10186) );
  NAND2_X1 U8021 ( .A1(n8625), .A2(n8624), .ZN(n12690) );
  AND4_X1 U8022 ( .A1(n8906), .A2(n8905), .A3(n8904), .A4(n8903), .ZN(n11976)
         );
  NAND2_X1 U8023 ( .A1(n10985), .A2(n7080), .ZN(n11990) );
  NAND2_X1 U8024 ( .A1(n6620), .A2(n6619), .ZN(n12001) );
  INV_X1 U8025 ( .A(n12277), .ZN(n12584) );
  INV_X1 U8026 ( .A(n12073), .ZN(n12041) );
  INV_X1 U8027 ( .A(n12533), .ZN(n12508) );
  INV_X1 U8028 ( .A(n12222), .ZN(n12568) );
  INV_X1 U8029 ( .A(n11976), .ZN(n12596) );
  NAND2_X1 U8030 ( .A1(n10704), .A2(n10703), .ZN(n10702) );
  NOR2_X1 U8031 ( .A1(n14481), .A2(n14482), .ZN(n14480) );
  NOR2_X1 U8032 ( .A1(n12385), .A2(n12709), .ZN(n12402) );
  INV_X1 U8033 ( .A(n7105), .ZN(n12421) );
  INV_X1 U8034 ( .A(n7103), .ZN(n12430) );
  AOI21_X1 U8035 ( .B1(n12423), .B2(n15100), .A(n12422), .ZN(n7179) );
  NAND2_X1 U8036 ( .A1(n7103), .A2(n12429), .ZN(n7102) );
  NOR2_X1 U8037 ( .A1(n12427), .A2(n12426), .ZN(n6935) );
  NOR2_X1 U8038 ( .A1(n6608), .A2(n6856), .ZN(n6855) );
  NAND2_X1 U8039 ( .A1(n6858), .A2(n15100), .ZN(n6857) );
  INV_X1 U8040 ( .A(n12444), .ZN(n6856) );
  NAND2_X1 U8041 ( .A1(n9012), .A2(n9011), .ZN(n11866) );
  AOI21_X1 U8042 ( .B1(n9041), .B2(n15149), .A(n9040), .ZN(n11867) );
  OAI21_X1 U8043 ( .B1(n6849), .B2(n12582), .A(n6847), .ZN(n12668) );
  INV_X1 U8044 ( .A(n6848), .ZN(n6847) );
  OAI22_X1 U8045 ( .A1(n12483), .A2(n12646), .B1(n12642), .B2(n12484), .ZN(
        n6848) );
  NAND2_X1 U8046 ( .A1(n8945), .A2(n8944), .ZN(n12680) );
  AND2_X1 U8047 ( .A1(n8811), .A2(n8810), .ZN(n11436) );
  NOR2_X1 U8048 ( .A1(n11237), .A2(n15138), .ZN(n14499) );
  NOR2_X1 U8049 ( .A1(n12665), .A2(n6495), .ZN(n12729) );
  OR2_X1 U8050 ( .A1(n11150), .A2(n9010), .ZN(n8979) );
  NAND2_X1 U8051 ( .A1(n9083), .A2(n9082), .ZN(n10261) );
  NAND2_X1 U8052 ( .A1(n8912), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8914) );
  NAND2_X1 U8053 ( .A1(n12885), .A2(n7400), .ZN(n12779) );
  OR2_X1 U8054 ( .A1(n10833), .A2(n10832), .ZN(n6711) );
  INV_X1 U8055 ( .A(n12821), .ZN(n7062) );
  OR2_X1 U8056 ( .A1(n12827), .A2(n7068), .ZN(n12872) );
  INV_X1 U8057 ( .A(n12860), .ZN(n12893) );
  OR2_X1 U8058 ( .A1(n8501), .A2(n8500), .ZN(n8502) );
  INV_X1 U8059 ( .A(n7040), .ZN(n7039) );
  AOI21_X1 U8060 ( .B1(n7040), .B2(n8369), .A(n7505), .ZN(n7038) );
  OAI21_X1 U8061 ( .B1(n8371), .B2(n8369), .A(n7040), .ZN(n7506) );
  INV_X1 U8062 ( .A(n6786), .ZN(n8371) );
  NOR2_X1 U8063 ( .A1(n7505), .A2(n8508), .ZN(n7504) );
  NAND2_X1 U8064 ( .A1(n7816), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7778) );
  NAND2_X1 U8065 ( .A1(n6440), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7779) );
  NAND2_X1 U8066 ( .A1(n14839), .A2(n9888), .ZN(n14853) );
  NAND2_X1 U8067 ( .A1(n6717), .A2(n6716), .ZN(n14882) );
  INV_X1 U8068 ( .A(n14879), .ZN(n6716) );
  INV_X1 U8069 ( .A(n14880), .ZN(n6717) );
  NAND2_X1 U8070 ( .A1(n8394), .A2(n8393), .ZN(n13244) );
  XNOR2_X1 U8071 ( .A(n13026), .B(n6910), .ZN(n13028) );
  INV_X1 U8072 ( .A(n13034), .ZN(n6910) );
  NAND2_X1 U8073 ( .A1(n7341), .A2(n7338), .ZN(n13055) );
  NAND2_X1 U8074 ( .A1(n7341), .A2(n11721), .ZN(n13053) );
  NAND2_X1 U8075 ( .A1(n7720), .A2(n7719), .ZN(n13307) );
  NAND2_X1 U8076 ( .A1(n8075), .A2(n8074), .ZN(n13318) );
  NOR2_X1 U8077 ( .A1(n10040), .A2(n6938), .ZN(n10370) );
  NAND2_X1 U8078 ( .A1(n13219), .A2(n10085), .ZN(n13236) );
  AND2_X1 U8079 ( .A1(n10378), .A2(n11580), .ZN(n13131) );
  AND2_X1 U8080 ( .A1(n7740), .A2(n7315), .ZN(n7314) );
  INV_X1 U8081 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7315) );
  MUX2_X1 U8082 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7733), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n7734) );
  NOR2_X1 U8083 ( .A1(n6980), .A2(n15379), .ZN(n6978) );
  AND2_X1 U8084 ( .A1(n6982), .A2(n6571), .ZN(n6980) );
  NAND2_X1 U8085 ( .A1(n6982), .A2(n6985), .ZN(n6981) );
  AOI21_X1 U8086 ( .B1(n6460), .B2(n7493), .A(n6548), .ZN(n7490) );
  INV_X1 U8087 ( .A(n13578), .ZN(n13394) );
  INV_X1 U8088 ( .A(n13485), .ZN(n6887) );
  NAND2_X1 U8089 ( .A1(n6722), .A2(n6721), .ZN(n13484) );
  NAND2_X1 U8090 ( .A1(n13381), .A2(n6724), .ZN(n6722) );
  AOI21_X1 U8091 ( .B1(n6724), .B2(n6726), .A(n6523), .ZN(n6721) );
  AOI21_X1 U8092 ( .B1(n7472), .B2(n7475), .A(n6725), .ZN(n6724) );
  AND2_X1 U8093 ( .A1(n10737), .A2(n14758), .ZN(n14562) );
  AND2_X1 U8094 ( .A1(n10288), .A2(n14316), .ZN(n15385) );
  AOI21_X1 U8095 ( .B1(n13764), .B2(n13763), .A(n6897), .ZN(n6896) );
  INV_X1 U8096 ( .A(n13760), .ZN(n6897) );
  OR3_X1 U8097 ( .A1(n9459), .A2(n9458), .A3(n9457), .ZN(n13776) );
  NAND2_X1 U8098 ( .A1(n6899), .A2(n13966), .ZN(n14162) );
  NAND2_X1 U8099 ( .A1(n6900), .A2(n13975), .ZN(n6899) );
  NAND2_X1 U8100 ( .A1(n7415), .A2(n9553), .ZN(n6900) );
  NAND2_X1 U8101 ( .A1(n9570), .A2(n6963), .ZN(n9612) );
  AND2_X1 U8102 ( .A1(n9569), .A2(n7644), .ZN(n6963) );
  XNOR2_X1 U8103 ( .A(n14369), .B(n14865), .ZN(n15397) );
  NAND2_X1 U8104 ( .A1(n15404), .A2(n6917), .ZN(n15396) );
  OAI21_X1 U8105 ( .B1(n15406), .B2(n15405), .A(n6918), .ZN(n6917) );
  OR2_X1 U8106 ( .A1(n14440), .A2(n6789), .ZN(n6787) );
  AND2_X1 U8107 ( .A1(n14440), .A2(n6789), .ZN(n6788) );
  NAND2_X1 U8108 ( .A1(n14613), .A2(n14612), .ZN(n14611) );
  OAI21_X1 U8109 ( .B1(n14473), .B2(n14474), .A(n14989), .ZN(n7324) );
  OR2_X1 U8110 ( .A1(n7371), .A2(n13592), .ZN(n7372) );
  AOI21_X1 U8111 ( .B1(n12916), .B2(n8363), .A(n7806), .ZN(n7814) );
  NAND2_X1 U8112 ( .A1(n13604), .A2(n13606), .ZN(n6894) );
  NOR2_X1 U8113 ( .A1(n6782), .A2(n7050), .ZN(n6781) );
  INV_X1 U8114 ( .A(n7854), .ZN(n6782) );
  OR2_X1 U8115 ( .A1(n7373), .A2(n13617), .ZN(n6865) );
  INV_X1 U8116 ( .A(n13616), .ZN(n7373) );
  NAND2_X1 U8117 ( .A1(n7877), .A2(n7878), .ZN(n7876) );
  NAND2_X1 U8118 ( .A1(n13629), .A2(n13627), .ZN(n7363) );
  NAND2_X1 U8119 ( .A1(n6775), .A2(n7043), .ZN(n7942) );
  NAND2_X1 U8120 ( .A1(n7922), .A2(n6502), .ZN(n7043) );
  NAND2_X1 U8121 ( .A1(n7525), .A2(n6467), .ZN(n7524) );
  OR2_X1 U8122 ( .A1(n13633), .A2(n13632), .ZN(n13634) );
  NAND2_X1 U8123 ( .A1(n13650), .A2(n13649), .ZN(n6923) );
  INV_X1 U8124 ( .A(n8003), .ZN(n7528) );
  INV_X1 U8125 ( .A(n8004), .ZN(n7530) );
  NAND2_X1 U8126 ( .A1(n6533), .A2(n7987), .ZN(n7531) );
  NAND2_X1 U8127 ( .A1(n6549), .A2(n8025), .ZN(n7537) );
  NAND2_X1 U8128 ( .A1(n7538), .A2(n7536), .ZN(n7535) );
  NOR2_X1 U8129 ( .A1(n8068), .A2(n8065), .ZN(n7534) );
  NAND2_X1 U8130 ( .A1(n13698), .A2(n13697), .ZN(n7359) );
  NAND2_X1 U8131 ( .A1(n6921), .A2(n13693), .ZN(n13694) );
  OR2_X1 U8132 ( .A1(n13692), .A2(n13691), .ZN(n13695) );
  INV_X1 U8133 ( .A(n7359), .ZN(n7358) );
  INV_X1 U8134 ( .A(n8112), .ZN(n7036) );
  NAND2_X1 U8135 ( .A1(n7361), .A2(n6521), .ZN(n13707) );
  INV_X1 U8136 ( .A(n13702), .ZN(n7362) );
  OAI21_X1 U8137 ( .B1(n8158), .B2(n7521), .A(n7519), .ZN(n8181) );
  INV_X1 U8138 ( .A(n7517), .ZN(n7516) );
  INV_X1 U8139 ( .A(n15148), .ZN(n10197) );
  NOR2_X1 U8140 ( .A1(n6795), .A2(n11445), .ZN(n6794) );
  AND2_X1 U8141 ( .A1(n8281), .A2(SI_26_), .ZN(n7622) );
  INV_X1 U8142 ( .A(n7599), .ZN(n7598) );
  OAI21_X1 U8143 ( .B1(n8207), .B2(n7600), .A(n8249), .ZN(n7599) );
  INV_X1 U8144 ( .A(SI_13_), .ZN(n7682) );
  NAND2_X1 U8145 ( .A1(n6812), .A2(n8027), .ZN(n6811) );
  INV_X1 U8146 ( .A(n7681), .ZN(n6812) );
  NAND2_X1 U8147 ( .A1(n6700), .A2(n12247), .ZN(n6699) );
  MUX2_X1 U8148 ( .A(n12246), .B(n12245), .S(n12244), .Z(n12247) );
  NOR2_X1 U8149 ( .A1(n12477), .A2(n7249), .ZN(n7248) );
  NAND2_X1 U8150 ( .A1(n6443), .A2(n6624), .ZN(n6623) );
  INV_X1 U8151 ( .A(n6610), .ZN(n6624) );
  OR2_X1 U8152 ( .A1(n9085), .A2(P3_D_REG_0__SCAN_IN), .ZN(n7258) );
  AOI21_X1 U8153 ( .B1(n7111), .B2(n8855), .A(n8868), .ZN(n7110) );
  INV_X1 U8154 ( .A(n10896), .ZN(n7294) );
  XNOR2_X1 U8155 ( .A(n14082), .B(n13553), .ZN(n13551) );
  AOI21_X1 U8156 ( .B1(n8296), .B2(n7622), .A(n7621), .ZN(n7620) );
  INV_X1 U8157 ( .A(n8311), .ZN(n7621) );
  AOI21_X1 U8158 ( .B1(n8296), .B2(n8281), .A(SI_26_), .ZN(n7623) );
  INV_X1 U8159 ( .A(n8281), .ZN(n7618) );
  NAND2_X1 U8160 ( .A1(n7620), .A2(n7616), .ZN(n7615) );
  INV_X1 U8161 ( .A(n7622), .ZN(n7616) );
  NAND2_X1 U8162 ( .A1(n7137), .A2(n8086), .ZN(n7136) );
  INV_X1 U8163 ( .A(n7627), .ZN(n7137) );
  NAND2_X1 U8164 ( .A1(n7611), .A2(n7613), .ZN(n7610) );
  INV_X1 U8165 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14327) );
  INV_X1 U8166 ( .A(n11655), .ZN(n7274) );
  OR2_X1 U8167 ( .A1(n11982), .A2(n7086), .ZN(n7085) );
  NAND2_X1 U8168 ( .A1(n6487), .A2(n7086), .ZN(n7083) );
  INV_X1 U8169 ( .A(n15143), .ZN(n9042) );
  INV_X1 U8170 ( .A(n7080), .ZN(n7079) );
  NAND2_X1 U8171 ( .A1(n11132), .A2(n11129), .ZN(n6878) );
  NAND2_X1 U8172 ( .A1(n14518), .A2(n12450), .ZN(n6992) );
  AND2_X1 U8173 ( .A1(n12263), .A2(n12085), .ZN(n12265) );
  NAND2_X1 U8174 ( .A1(n6446), .A2(n10412), .ZN(n6920) );
  NOR2_X1 U8175 ( .A1(n10619), .A2(n6641), .ZN(n7095) );
  NAND2_X1 U8176 ( .A1(n10626), .A2(n10625), .ZN(n10628) );
  INV_X1 U8177 ( .A(n15069), .ZN(n6634) );
  INV_X1 U8178 ( .A(n15063), .ZN(n6655) );
  OR2_X1 U8179 ( .A1(n11866), .A2(n12458), .ZN(n12258) );
  NOR2_X1 U8180 ( .A1(n7248), .A2(n7245), .ZN(n7244) );
  INV_X1 U8181 ( .A(n8989), .ZN(n7245) );
  OR2_X1 U8182 ( .A1(n7246), .A2(n7248), .ZN(n7243) );
  NAND2_X1 U8183 ( .A1(n9056), .A2(n12274), .ZN(n7250) );
  AND2_X1 U8184 ( .A1(n12471), .A2(n7250), .ZN(n7246) );
  OR2_X1 U8185 ( .A1(n9056), .A2(n12497), .ZN(n12245) );
  NOR2_X1 U8186 ( .A1(n8939), .A2(n7234), .ZN(n7233) );
  INV_X1 U8187 ( .A(n7238), .ZN(n7234) );
  NAND2_X1 U8188 ( .A1(n7235), .A2(n7233), .ZN(n7231) );
  INV_X1 U8189 ( .A(n7549), .ZN(n7008) );
  AOI21_X1 U8190 ( .B1(n7552), .B2(n7554), .A(n7550), .ZN(n7549) );
  INV_X1 U8191 ( .A(n12230), .ZN(n7550) );
  NOR2_X1 U8192 ( .A1(n7551), .A2(n7011), .ZN(n7010) );
  INV_X1 U8193 ( .A(n12206), .ZN(n7011) );
  INV_X1 U8194 ( .A(n12200), .ZN(n7004) );
  OAI21_X1 U8195 ( .B1(n12630), .B2(n7004), .A(n12614), .ZN(n7003) );
  OR2_X1 U8196 ( .A1(n8847), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8862) );
  NOR2_X1 U8197 ( .A1(n12630), .A2(n7221), .ZN(n7220) );
  INV_X1 U8198 ( .A(n12192), .ZN(n7561) );
  INV_X1 U8199 ( .A(n12188), .ZN(n7563) );
  OR2_X1 U8200 ( .A1(n12282), .A2(n11027), .ZN(n12165) );
  INV_X1 U8201 ( .A(n11021), .ZN(n12162) );
  AOI21_X1 U8202 ( .B1(n6996), .B2(n6998), .A(n6995), .ZN(n6994) );
  INV_X1 U8203 ( .A(n12159), .ZN(n6995) );
  NAND2_X1 U8204 ( .A1(n15121), .A2(n12130), .ZN(n15107) );
  NAND2_X1 U8205 ( .A1(n15122), .A2(n7210), .ZN(n15121) );
  NAND2_X1 U8206 ( .A1(n8943), .A2(n8564), .ZN(n8565) );
  NAND2_X1 U8207 ( .A1(n6693), .A2(n8554), .ZN(n8555) );
  OAI21_X1 U8208 ( .B1(n8894), .B2(n6692), .A(n6690), .ZN(n6693) );
  INV_X1 U8209 ( .A(n6691), .ZN(n6690) );
  INV_X1 U8210 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n8577) );
  NAND2_X1 U8211 ( .A1(n8814), .A2(n8538), .ZN(n8541) );
  INV_X1 U8212 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n8542) );
  INV_X1 U8213 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8539) );
  INV_X1 U8214 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7546) );
  NAND2_X1 U8215 ( .A1(n7393), .A2(n7068), .ZN(n7066) );
  XNOR2_X1 U8216 ( .A(n13290), .B(n11592), .ZN(n11575) );
  NAND2_X1 U8217 ( .A1(n6777), .A2(n7513), .ZN(n8270) );
  NAND2_X1 U8218 ( .A1(n8246), .A2(n6505), .ZN(n7513) );
  AOI21_X1 U8219 ( .B1(n8445), .B2(n8444), .A(n6504), .ZN(n7510) );
  NOR2_X1 U8220 ( .A1(n6756), .A2(n7346), .ZN(n6755) );
  INV_X1 U8221 ( .A(n7347), .ZN(n7346) );
  INV_X1 U8222 ( .A(n6758), .ZN(n6756) );
  NOR2_X1 U8223 ( .A1(n13266), .A2(n13259), .ZN(n6946) );
  AOI21_X1 U8224 ( .B1(n7355), .B2(n11712), .A(n6527), .ZN(n7353) );
  NOR2_X1 U8225 ( .A1(n7354), .A2(n6752), .ZN(n6751) );
  INV_X1 U8226 ( .A(n11711), .ZN(n6752) );
  INV_X1 U8227 ( .A(n7355), .ZN(n7354) );
  OR2_X1 U8228 ( .A1(n8077), .A2(n8076), .ZN(n8096) );
  AND2_X1 U8229 ( .A1(n13064), .A2(n6455), .ZN(n13018) );
  INV_X1 U8230 ( .A(n13318), .ZN(n6943) );
  NOR2_X1 U8231 ( .A1(n11361), .A2(n11704), .ZN(n6940) );
  INV_X1 U8232 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n7705) );
  INV_X1 U8233 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8480) );
  INV_X1 U8234 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7712) );
  INV_X1 U8235 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7711) );
  OR2_X1 U8236 ( .A1(n7949), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n7971) );
  OR2_X1 U8237 ( .A1(n7927), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n7949) );
  INV_X1 U8238 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7698) );
  OR2_X1 U8239 ( .A1(n11747), .A2(n11746), .ZN(n11748) );
  NAND2_X1 U8240 ( .A1(n13723), .A2(n7368), .ZN(n7367) );
  AND2_X1 U8241 ( .A1(n13736), .A2(n7366), .ZN(n7365) );
  OR2_X1 U8242 ( .A1(n13723), .A2(n7368), .ZN(n7366) );
  INV_X1 U8243 ( .A(n13665), .ZN(n7417) );
  NOR2_X1 U8244 ( .A1(n13663), .A2(n7423), .ZN(n7422) );
  INV_X1 U8245 ( .A(n9545), .ZN(n7423) );
  NOR2_X1 U8246 ( .A1(n7420), .A2(n6966), .ZN(n6965) );
  INV_X1 U8247 ( .A(n6968), .ZN(n6966) );
  NAND2_X1 U8248 ( .A1(n7185), .A2(n14757), .ZN(n13573) );
  NAND2_X1 U8249 ( .A1(n9977), .A2(n9173), .ZN(n13562) );
  NAND2_X1 U8250 ( .A1(n9566), .A2(n9590), .ZN(n13564) );
  NAND2_X1 U8251 ( .A1(n14004), .A2(n7157), .ZN(n13984) );
  NAND2_X1 U8252 ( .A1(n14004), .A2(n14005), .ZN(n14006) );
  NAND2_X1 U8253 ( .A1(n7404), .A2(n7407), .ZN(n14457) );
  AOI21_X1 U8254 ( .B1(n7408), .B2(n13532), .A(n6530), .ZN(n7407) );
  AOI21_X1 U8255 ( .B1(n8389), .B2(n7607), .A(n7606), .ZN(n7605) );
  INV_X1 U8256 ( .A(n8377), .ZN(n7606) );
  INV_X1 U8257 ( .A(n8372), .ZN(n7607) );
  NAND2_X1 U8258 ( .A1(n6876), .A2(n6602), .ZN(n8314) );
  INV_X1 U8259 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6728) );
  INV_X1 U8260 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6727) );
  OR2_X1 U8261 ( .A1(n8185), .A2(n10182), .ZN(n8186) );
  NAND2_X1 U8262 ( .A1(n8115), .A2(n7587), .ZN(n7585) );
  INV_X1 U8263 ( .A(n8142), .ZN(n8143) );
  NAND2_X1 U8264 ( .A1(n7629), .A2(n7628), .ZN(n7627) );
  INV_X1 U8265 ( .A(SI_15_), .ZN(n7628) );
  INV_X1 U8266 ( .A(n7688), .ZN(n7629) );
  INV_X1 U8267 ( .A(n8069), .ZN(n7624) );
  OR2_X1 U8268 ( .A1(n9288), .A2(n9287), .ZN(n9302) );
  INV_X1 U8269 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9285) );
  INV_X1 U8270 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9244) );
  NAND2_X1 U8271 ( .A1(n7034), .A2(SI_7_), .ZN(n7668) );
  NOR2_X1 U8272 ( .A1(n7576), .A2(n7122), .ZN(n7121) );
  NAND2_X1 U8273 ( .A1(n7840), .A2(n7663), .ZN(n7856) );
  OAI21_X1 U8274 ( .B1(SI_5_), .B2(n7072), .A(n7665), .ZN(n7664) );
  NAND2_X1 U8275 ( .A1(n7577), .A2(n7584), .ZN(n6796) );
  OAI21_X1 U8276 ( .B1(n7581), .B2(n7653), .A(n7579), .ZN(n7578) );
  NAND2_X1 U8277 ( .A1(n6796), .A2(SI_1_), .ZN(n7657) );
  INV_X1 U8278 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7331) );
  OAI21_X1 U8279 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n14342), .A(n14341), .ZN(
        n14366) );
  AOI21_X1 U8280 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n14660), .A(n14349), .ZN(
        n14360) );
  NOR2_X1 U8281 ( .A1(n14363), .A2(n14362), .ZN(n14349) );
  XNOR2_X1 U8282 ( .A(n11165), .B(n11622), .ZN(n11876) );
  NAND2_X1 U8283 ( .A1(n10268), .A2(n9042), .ZN(n12126) );
  INV_X1 U8284 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10618) );
  NAND2_X1 U8285 ( .A1(n7253), .A2(n7252), .ZN(n11973) );
  NAND2_X1 U8286 ( .A1(n10990), .A2(n6850), .ZN(n11989) );
  NAND2_X1 U8287 ( .A1(n6851), .A2(n15108), .ZN(n6850) );
  NAND2_X1 U8288 ( .A1(n11922), .A2(n11642), .ZN(n6618) );
  AND2_X1 U8289 ( .A1(n11434), .A2(n11435), .ZN(n11935) );
  NAND2_X1 U8290 ( .A1(n11888), .A2(n14507), .ZN(n7266) );
  NAND2_X1 U8291 ( .A1(n7268), .A2(n6494), .ZN(n7269) );
  NAND2_X1 U8292 ( .A1(n12019), .A2(n6485), .ZN(n7267) );
  NAND2_X1 U8293 ( .A1(n11871), .A2(n7216), .ZN(n7214) );
  NAND2_X1 U8294 ( .A1(n6646), .A2(n6645), .ZN(n10674) );
  OR2_X1 U8295 ( .A1(n10445), .A2(n10477), .ZN(n6645) );
  OAI21_X1 U8296 ( .B1(n10717), .B2(n10716), .A(n7640), .ZN(n10715) );
  OR2_X1 U8297 ( .A1(n10670), .A2(n10475), .ZN(n10672) );
  INV_X1 U8298 ( .A(n7095), .ZN(n7100) );
  NAND2_X1 U8299 ( .A1(n7182), .A2(n10658), .ZN(n6651) );
  NAND3_X1 U8300 ( .A1(n7093), .A2(n7094), .A3(n7096), .ZN(n10661) );
  NOR2_X1 U8301 ( .A1(n7095), .A2(n10614), .ZN(n7094) );
  NAND2_X1 U8302 ( .A1(n6639), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n10655) );
  NAND2_X1 U8303 ( .A1(n6638), .A2(n10652), .ZN(n10937) );
  NAND2_X1 U8304 ( .A1(n10655), .A2(n10653), .ZN(n6638) );
  XNOR2_X1 U8305 ( .A(n10938), .B(n15053), .ZN(n15057) );
  AND2_X1 U8306 ( .A1(n6651), .A2(n7181), .ZN(n10957) );
  NAND2_X1 U8307 ( .A1(n10956), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7181) );
  AND2_X1 U8308 ( .A1(n10937), .A2(n7167), .ZN(n10938) );
  NAND2_X1 U8309 ( .A1(n10956), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7167) );
  NOR2_X1 U8310 ( .A1(n11067), .A2(n6864), .ZN(n11400) );
  NOR2_X1 U8311 ( .A1(n11072), .A2(n10942), .ZN(n6864) );
  XNOR2_X1 U8312 ( .A(n6888), .B(n11069), .ZN(n11082) );
  OR2_X1 U8313 ( .A1(n8752), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8769) );
  NOR2_X1 U8314 ( .A1(n11401), .A2(n11402), .ZN(n15070) );
  NOR2_X1 U8315 ( .A1(n8760), .A2(n11082), .ZN(n11420) );
  INV_X1 U8316 ( .A(n6888), .ZN(n11418) );
  NAND2_X1 U8317 ( .A1(n6633), .A2(n6631), .ZN(n6930) );
  AOI21_X1 U8318 ( .B1(n11402), .B2(n6634), .A(n6632), .ZN(n6631) );
  NAND2_X1 U8319 ( .A1(n11401), .A2(n6634), .ZN(n6633) );
  INV_X1 U8320 ( .A(n11403), .ZN(n6632) );
  INV_X1 U8321 ( .A(n12338), .ZN(n7160) );
  INV_X1 U8322 ( .A(n12322), .ZN(n6644) );
  OR2_X1 U8323 ( .A1(n12334), .A2(n7108), .ZN(n6663) );
  INV_X1 U8324 ( .A(n12369), .ZN(n7108) );
  INV_X1 U8325 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n15254) );
  XNOR2_X1 U8326 ( .A(n6931), .B(n14484), .ZN(n14486) );
  OR2_X1 U8327 ( .A1(n12360), .A2(n12361), .ZN(n14489) );
  OR2_X1 U8328 ( .A1(n12417), .A2(n12386), .ZN(n6661) );
  INV_X1 U8329 ( .A(n6662), .ZN(n12418) );
  NAND2_X1 U8330 ( .A1(n6662), .A2(n6489), .ZN(n7105) );
  AND2_X1 U8331 ( .A1(n12387), .A2(n12386), .ZN(n12416) );
  INV_X1 U8332 ( .A(n12440), .ZN(n6859) );
  OAI21_X1 U8333 ( .B1(n12492), .B2(n7242), .A(n7240), .ZN(n12455) );
  INV_X1 U8334 ( .A(n7244), .ZN(n7242) );
  AND2_X1 U8335 ( .A1(n7243), .A2(n7241), .ZN(n7240) );
  NAND2_X1 U8336 ( .A1(n7244), .A2(n6534), .ZN(n7241) );
  OR2_X1 U8337 ( .A1(n8980), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8982) );
  NAND2_X1 U8338 ( .A1(n6821), .A2(n6820), .ZN(n12482) );
  AOI21_X1 U8339 ( .B1(n6824), .B2(n6825), .A(n6534), .ZN(n6820) );
  NAND2_X1 U8340 ( .A1(n12498), .A2(n9055), .ZN(n12485) );
  NOR2_X1 U8341 ( .A1(n7540), .A2(n12510), .ZN(n7539) );
  INV_X1 U8342 ( .A(n7542), .ZN(n7540) );
  NAND2_X1 U8343 ( .A1(n8602), .A2(n8601), .ZN(n8968) );
  INV_X1 U8344 ( .A(n8956), .ZN(n8602) );
  NAND2_X1 U8345 ( .A1(n8600), .A2(n8599), .ZN(n8931) );
  INV_X1 U8346 ( .A(n8631), .ZN(n8600) );
  NAND2_X1 U8347 ( .A1(n12593), .A2(n8892), .ZN(n12579) );
  NAND2_X1 U8348 ( .A1(n8596), .A2(n8595), .ZN(n8901) );
  INV_X1 U8349 ( .A(n8886), .ZN(n8596) );
  NAND2_X1 U8350 ( .A1(n12595), .A2(n12594), .ZN(n12593) );
  NAND2_X1 U8351 ( .A1(n8594), .A2(n15254), .ZN(n8873) );
  INV_X1 U8352 ( .A(n8862), .ZN(n8594) );
  OR2_X1 U8353 ( .A1(n8873), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8886) );
  NAND2_X1 U8354 ( .A1(n12609), .A2(n12608), .ZN(n12607) );
  NAND2_X1 U8355 ( .A1(n14504), .A2(n8837), .ZN(n12641) );
  NAND2_X1 U8356 ( .A1(n8593), .A2(n12024), .ZN(n8847) );
  INV_X1 U8357 ( .A(n8831), .ZN(n8593) );
  OAI21_X1 U8358 ( .B1(n11385), .B2(n12099), .A(n8825), .ZN(n14506) );
  NAND2_X1 U8359 ( .A1(n8592), .A2(n8591), .ZN(n8831) );
  INV_X1 U8360 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n8591) );
  INV_X1 U8361 ( .A(n8819), .ZN(n8592) );
  NAND2_X1 U8362 ( .A1(n11331), .A2(n12173), .ZN(n11387) );
  AND2_X1 U8363 ( .A1(n12180), .A2(n12184), .ZN(n12099) );
  OR2_X1 U8364 ( .A1(n8796), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8819) );
  NAND2_X1 U8365 ( .A1(n8795), .A2(n8794), .ZN(n11334) );
  NOR2_X1 U8366 ( .A1(n7227), .A2(n7225), .ZN(n7224) );
  AND2_X1 U8367 ( .A1(n7226), .A2(n6453), .ZN(n11230) );
  NAND2_X1 U8368 ( .A1(n8590), .A2(n11077), .ZN(n8775) );
  AND2_X1 U8369 ( .A1(n8741), .A2(n8740), .ZN(n11022) );
  NAND2_X1 U8370 ( .A1(n11116), .A2(n8726), .ZN(n11168) );
  NAND2_X1 U8371 ( .A1(n8589), .A2(n11878), .ZN(n8742) );
  INV_X1 U8372 ( .A(n8728), .ZN(n8589) );
  NAND2_X1 U8373 ( .A1(n11111), .A2(n12154), .ZN(n11166) );
  NAND2_X1 U8374 ( .A1(n10809), .A2(n7229), .ZN(n11116) );
  AND2_X1 U8375 ( .A1(n8725), .A2(n8706), .ZN(n7229) );
  NAND2_X1 U8376 ( .A1(n10809), .A2(n8706), .ZN(n11114) );
  OR2_X1 U8377 ( .A1(n8708), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8728) );
  NAND2_X1 U8378 ( .A1(n11109), .A2(n12092), .ZN(n11111) );
  INV_X1 U8379 ( .A(n10693), .ZN(n12141) );
  OR2_X1 U8380 ( .A1(n9010), .A2(n6901), .ZN(n8689) );
  INV_X1 U8381 ( .A(n9622), .ZN(n6901) );
  NAND2_X1 U8382 ( .A1(n12138), .A2(n12137), .ZN(n15110) );
  NAND2_X1 U8383 ( .A1(n15111), .A2(n15110), .ZN(n15109) );
  INV_X1 U8384 ( .A(n7210), .ZN(n15126) );
  NAND2_X1 U8385 ( .A1(n15127), .A2(n15126), .ZN(n15125) );
  INV_X1 U8386 ( .A(n12126), .ZN(n15141) );
  AND2_X1 U8387 ( .A1(n9065), .A2(n9116), .ZN(n15153) );
  INV_X1 U8388 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8611) );
  OAI21_X1 U8389 ( .B1(n8991), .B2(n8990), .A(n8992), .ZN(n9005) );
  OAI21_X1 U8390 ( .B1(n8965), .B2(n8568), .A(n8569), .ZN(n8977) );
  XNOR2_X1 U8391 ( .A(n8565), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n8953) );
  XNOR2_X1 U8392 ( .A(n9101), .B(n9069), .ZN(n10394) );
  NAND2_X1 U8393 ( .A1(n9100), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9101) );
  NAND2_X1 U8394 ( .A1(n6684), .A2(n8549), .ZN(n8881) );
  OAI21_X1 U8395 ( .B1(n8839), .B2(n6683), .A(n6679), .ZN(n6684) );
  INV_X1 U8396 ( .A(n7111), .ZN(n6683) );
  OR2_X1 U8397 ( .A1(n8858), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n8882) );
  XNOR2_X1 U8398 ( .A(n8543), .B(n8542), .ZN(n8826) );
  NOR2_X1 U8399 ( .A1(n8687), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n7547) );
  AND2_X1 U8400 ( .A1(n8534), .A2(n8533), .ZN(n8765) );
  AND2_X1 U8401 ( .A1(n8532), .A2(n8531), .ZN(n8748) );
  OAI21_X1 U8402 ( .B1(n6688), .B2(n6687), .A(n6685), .ZN(n8736) );
  INV_X1 U8403 ( .A(n8528), .ZN(n6687) );
  AOI21_X1 U8404 ( .B1(n6686), .B2(n8528), .A(n6545), .ZN(n6685) );
  AND2_X1 U8405 ( .A1(n8721), .A2(n8752), .ZN(n10657) );
  OAI21_X1 U8406 ( .B1(n8661), .B2(n8672), .A(n6694), .ZN(n8686) );
  AOI21_X1 U8407 ( .B1(n8519), .B2(n6696), .A(n6695), .ZN(n6694) );
  INV_X1 U8408 ( .A(n8520), .ZN(n6695) );
  INV_X1 U8409 ( .A(n8517), .ZN(n6696) );
  INV_X1 U8410 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8665) );
  NOR2_X1 U8411 ( .A1(n8665), .A2(n9027), .ZN(n6649) );
  XNOR2_X1 U8412 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8641) );
  AND2_X1 U8413 ( .A1(n8513), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8650) );
  OR2_X1 U8414 ( .A1(n7977), .A2(n7976), .ZN(n7995) );
  AND2_X1 U8415 ( .A1(n11569), .A2(n12793), .ZN(n7395) );
  NAND2_X1 U8416 ( .A1(n9755), .A2(n6444), .ZN(n9756) );
  INV_X1 U8417 ( .A(n8167), .ZN(n8165) );
  NAND2_X1 U8418 ( .A1(n7750), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8015) );
  INV_X1 U8419 ( .A(n7995), .ZN(n7750) );
  OR2_X1 U8420 ( .A1(n8015), .A2(n8014), .ZN(n8032) );
  NAND2_X1 U8421 ( .A1(n8213), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8235) );
  INV_X1 U8422 ( .A(n8215), .ZN(n8213) );
  NAND2_X1 U8423 ( .A1(n12873), .A2(n7070), .ZN(n7068) );
  AND2_X1 U8424 ( .A1(n8504), .A2(n9774), .ZN(n9744) );
  INV_X1 U8425 ( .A(n11445), .ZN(n9774) );
  INV_X1 U8426 ( .A(n7816), .ZN(n8399) );
  NAND2_X1 U8427 ( .A1(n14840), .A2(n14841), .ZN(n14839) );
  NAND2_X1 U8428 ( .A1(n14866), .A2(n9895), .ZN(n14880) );
  NOR2_X1 U8429 ( .A1(n14915), .A2(n6601), .ZN(n14927) );
  AND2_X1 U8430 ( .A1(n14927), .A2(n14926), .ZN(n14928) );
  NOR2_X1 U8431 ( .A1(n12976), .A2(n6719), .ZN(n14978) );
  AND2_X1 U8432 ( .A1(n12975), .A2(n14980), .ZN(n6719) );
  NAND2_X1 U8433 ( .A1(n8425), .A2(n8424), .ZN(n12992) );
  OR2_X1 U8434 ( .A1(n8355), .A2(n8326), .ZN(n11728) );
  AND2_X1 U8435 ( .A1(n8353), .A2(n8287), .ZN(n13031) );
  NAND2_X1 U8436 ( .A1(n13064), .A2(n6946), .ZN(n13029) );
  OR2_X1 U8437 ( .A1(n8260), .A2(n15315), .ZN(n8300) );
  AOI21_X1 U8438 ( .B1(n7301), .B2(n7299), .A(n7304), .ZN(n7298) );
  AND2_X1 U8439 ( .A1(n13269), .A2(n13044), .ZN(n7304) );
  INV_X1 U8440 ( .A(n11695), .ZN(n7299) );
  INV_X1 U8441 ( .A(n7301), .ZN(n7300) );
  INV_X1 U8442 ( .A(n13080), .ZN(n7342) );
  NAND2_X1 U8443 ( .A1(n7174), .A2(n7173), .ZN(n13076) );
  INV_X1 U8444 ( .A(n13098), .ZN(n7174) );
  AND2_X1 U8445 ( .A1(n11693), .A2(n8453), .ZN(n13091) );
  NOR2_X1 U8446 ( .A1(n13286), .A2(n6948), .ZN(n6947) );
  INV_X1 U8447 ( .A(n6949), .ZN(n6948) );
  AOI21_X1 U8448 ( .B1(n7015), .B2(n7021), .A(n7016), .ZN(n7014) );
  INV_X1 U8449 ( .A(n7018), .ZN(n7017) );
  INV_X1 U8450 ( .A(n11690), .ZN(n7016) );
  NAND2_X1 U8451 ( .A1(n11731), .A2(n6949), .ZN(n13118) );
  INV_X1 U8452 ( .A(n11731), .ZN(n13157) );
  NAND2_X1 U8453 ( .A1(n11731), .A2(n7027), .ZN(n13142) );
  INV_X1 U8454 ( .A(n8124), .ZN(n8122) );
  NAND2_X1 U8455 ( .A1(n11710), .A2(n11709), .ZN(n13180) );
  NAND2_X1 U8456 ( .A1(n7311), .A2(n7310), .ZN(n13221) );
  NAND2_X1 U8457 ( .A1(n6553), .A2(n11678), .ZN(n7310) );
  AND2_X1 U8458 ( .A1(n8456), .A2(n11679), .ZN(n13222) );
  NAND2_X1 U8459 ( .A1(n7751), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8055) );
  INV_X1 U8460 ( .A(n8032), .ZN(n7751) );
  OR2_X1 U8461 ( .A1(n8055), .A2(n8054), .ZN(n8077) );
  INV_X1 U8462 ( .A(n13222), .ZN(n13215) );
  NAND2_X1 U8463 ( .A1(n11221), .A2(n14543), .ZN(n11365) );
  NAND2_X1 U8464 ( .A1(n11197), .A2(n11196), .ZN(n11209) );
  INV_X1 U8465 ( .A(n11191), .ZN(n11198) );
  XNOR2_X1 U8466 ( .A(n11376), .B(n12907), .ZN(n11191) );
  INV_X1 U8467 ( .A(n7168), .ZN(n11202) );
  NAND2_X1 U8468 ( .A1(n10870), .A2(n10879), .ZN(n10894) );
  INV_X1 U8469 ( .A(n7292), .ZN(n10897) );
  AOI21_X1 U8470 ( .B1(n10915), .B2(n10878), .A(n10879), .ZN(n7292) );
  NAND2_X1 U8471 ( .A1(n15010), .A2(n10556), .ZN(n10922) );
  NAND2_X1 U8472 ( .A1(n10562), .A2(n10561), .ZN(n10874) );
  NAND2_X1 U8473 ( .A1(n10132), .A2(n6501), .ZN(n10342) );
  NAND2_X1 U8474 ( .A1(n10132), .A2(n10380), .ZN(n10344) );
  NAND2_X1 U8475 ( .A1(n6936), .A2(n10372), .ZN(n10039) );
  AND2_X1 U8476 ( .A1(n12991), .A2(n11732), .ZN(n13245) );
  INV_X1 U8477 ( .A(n15030), .ZN(n13291) );
  NAND2_X1 U8478 ( .A1(n7770), .A2(n11372), .ZN(n15023) );
  NAND2_X1 U8479 ( .A1(n7706), .A2(n7523), .ZN(n8486) );
  AND2_X1 U8480 ( .A1(n8495), .A2(n8488), .ZN(n9727) );
  OR2_X1 U8481 ( .A1(n8071), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n8088) );
  NAND2_X1 U8482 ( .A1(n6710), .A2(n6709), .ZN(n7905) );
  INV_X1 U8483 ( .A(n7859), .ZN(n6710) );
  OR2_X1 U8484 ( .A1(n9236), .A2(n10749), .ZN(n9249) );
  XNOR2_X1 U8485 ( .A(n10743), .B(n11838), .ZN(n10845) );
  INV_X1 U8486 ( .A(n10974), .ZN(n7494) );
  INV_X1 U8487 ( .A(n7496), .ZN(n7493) );
  NAND2_X1 U8488 ( .A1(n9387), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9402) );
  OR2_X1 U8489 ( .A1(n9402), .A2(n13405), .ZN(n9409) );
  NAND2_X1 U8490 ( .A1(n10845), .A2(n6885), .ZN(n7650) );
  INV_X1 U8491 ( .A(n10846), .ZN(n6885) );
  INV_X1 U8492 ( .A(n9976), .ZN(n9986) );
  MUX2_X1 U8493 ( .A(n6473), .B(n9995), .S(n9996), .Z(n9976) );
  AND2_X1 U8494 ( .A1(n9983), .A2(n9982), .ZN(n9984) );
  OR2_X1 U8495 ( .A1(n11789), .A2(n11788), .ZN(n7636) );
  NOR2_X1 U8496 ( .A1(n9357), .A2(n9356), .ZN(n9370) );
  INV_X1 U8497 ( .A(n7470), .ZN(n7469) );
  NOR2_X1 U8498 ( .A1(n9262), .A2(n15259), .ZN(n9277) );
  INV_X1 U8499 ( .A(n10545), .ZN(n7457) );
  AOI21_X1 U8500 ( .B1(n7474), .B2(n7476), .A(n6529), .ZN(n7472) );
  INV_X1 U8501 ( .A(n13418), .ZN(n6725) );
  INV_X1 U8502 ( .A(n7472), .ZN(n6726) );
  OR2_X1 U8503 ( .A1(n9346), .A2(n9345), .ZN(n9357) );
  NAND2_X1 U8504 ( .A1(n6738), .A2(n6737), .ZN(n6736) );
  INV_X1 U8505 ( .A(n11750), .ZN(n6737) );
  INV_X1 U8506 ( .A(n11751), .ZN(n6738) );
  NAND2_X1 U8507 ( .A1(n11751), .A2(n11750), .ZN(n11755) );
  AOI211_X1 U8508 ( .C1(n13756), .C2(n13755), .A(n13754), .B(n13753), .ZN(
        n13760) );
  AND2_X1 U8509 ( .A1(n14320), .A2(n9566), .ZN(n13555) );
  AND4_X1 U8510 ( .A1(n9471), .A2(n9470), .A3(n9469), .A4(n9468), .ZN(n13486)
         );
  AND4_X1 U8511 ( .A1(n9351), .A2(n9350), .A3(n9349), .A4(n9348), .ZN(n11752)
         );
  AND4_X1 U8512 ( .A1(n9300), .A2(n9299), .A3(n9298), .A4(n9297), .ZN(n11471)
         );
  OR2_X1 U8513 ( .A1(n13506), .A2(n9145), .ZN(n9147) );
  OR2_X1 U8514 ( .A1(n9341), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n9232) );
  INV_X1 U8515 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n15259) );
  INV_X1 U8516 ( .A(n7428), .ZN(n9133) );
  NOR2_X1 U8517 ( .A1(n13735), .A2(n7156), .ZN(n7154) );
  NAND2_X1 U8518 ( .A1(n7187), .A2(n7186), .ZN(n13976) );
  AOI21_X1 U8519 ( .B1(n7188), .B2(n7190), .A(n6498), .ZN(n7186) );
  OAI21_X1 U8520 ( .B1(n14027), .B2(n6959), .A(n6541), .ZN(n7187) );
  INV_X1 U8521 ( .A(n7202), .ZN(n7200) );
  NAND2_X1 U8522 ( .A1(n6919), .A2(n13541), .ZN(n14057) );
  INV_X1 U8523 ( .A(n14055), .ZN(n6919) );
  OAI211_X1 U8524 ( .C1(n7442), .C2(n14106), .A(n7440), .B(n7441), .ZN(n14062)
         );
  OR2_X1 U8525 ( .A1(n14285), .A2(n13779), .ZN(n7440) );
  NAND2_X1 U8526 ( .A1(n7444), .A2(n7443), .ZN(n7442) );
  AOI21_X1 U8527 ( .B1(n7422), .B2(n7420), .A(n6491), .ZN(n7419) );
  INV_X1 U8528 ( .A(n7422), .ZN(n7421) );
  AND2_X1 U8529 ( .A1(n9394), .A2(n9393), .ZN(n14122) );
  OR2_X1 U8530 ( .A1(n14788), .A2(n14082), .ZN(n10641) );
  NAND2_X1 U8531 ( .A1(n6617), .A2(n6616), .ZN(n14459) );
  OR2_X1 U8532 ( .A1(n9987), .A2(n9801), .ZN(n13487) );
  AND4_X1 U8533 ( .A1(n9283), .A2(n9282), .A3(n9281), .A4(n9280), .ZN(n11344)
         );
  NAND2_X1 U8534 ( .A1(n7436), .A2(n7435), .ZN(n14680) );
  NAND2_X1 U8535 ( .A1(n6544), .A2(n9537), .ZN(n7435) );
  AOI21_X1 U8536 ( .B1(n13519), .B2(n7193), .A(n6458), .ZN(n7192) );
  NAND2_X1 U8537 ( .A1(n10489), .A2(n7193), .ZN(n7191) );
  NAND2_X1 U8538 ( .A1(n10588), .A2(n7431), .ZN(n7430) );
  OR2_X1 U8539 ( .A1(n7433), .A2(n7434), .ZN(n7432) );
  INV_X1 U8540 ( .A(n13590), .ZN(n7431) );
  NAND2_X1 U8541 ( .A1(n10225), .A2(n13576), .ZN(n10224) );
  OR2_X1 U8542 ( .A1(n14788), .A2(n13929), .ZN(n10494) );
  NAND2_X1 U8543 ( .A1(n14090), .A2(n9414), .ZN(n14079) );
  NAND2_X1 U8544 ( .A1(n9408), .A2(n9407), .ZN(n14215) );
  NAND2_X1 U8545 ( .A1(n11529), .A2(n9366), .ZN(n14137) );
  AOI21_X1 U8546 ( .B1(n6953), .B2(n6956), .A(n6952), .ZN(n6951) );
  OAI21_X1 U8547 ( .B1(n14447), .B2(n6956), .A(n6953), .ZN(n11518) );
  AND2_X1 U8548 ( .A1(n9333), .A2(n9332), .ZN(n15383) );
  OR3_X1 U8549 ( .A1(n14320), .A2(n13550), .A3(n13929), .ZN(n14789) );
  NAND2_X1 U8550 ( .A1(n10492), .A2(n9206), .ZN(n10595) );
  INV_X1 U8551 ( .A(n14807), .ZN(n14762) );
  OR2_X1 U8552 ( .A1(n10506), .A2(n9608), .ZN(n14796) );
  NAND2_X1 U8553 ( .A1(n10573), .A2(n14789), .ZN(n14807) );
  AOI21_X1 U8554 ( .B1(n7603), .B2(n7608), .A(n6603), .ZN(n7602) );
  NAND2_X1 U8555 ( .A1(n8392), .A2(n8391), .ZN(n13349) );
  NAND2_X1 U8556 ( .A1(n8390), .A2(n8389), .ZN(n8392) );
  OR2_X1 U8557 ( .A1(n8390), .A2(n8389), .ZN(n8391) );
  XNOR2_X1 U8558 ( .A(n8349), .B(n8348), .ZN(n13355) );
  OAI21_X1 U8559 ( .B1(n8297), .B2(n8296), .A(n8281), .ZN(n8312) );
  AND2_X1 U8560 ( .A1(n9574), .A2(n6451), .ZN(n9586) );
  XNOR2_X1 U8561 ( .A(n9521), .B(n9520), .ZN(n13553) );
  NAND2_X1 U8562 ( .A1(n9571), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9521) );
  XNOR2_X1 U8563 ( .A(n9524), .B(P1_IR_REG_20__SCAN_IN), .ZN(n13550) );
  NAND2_X1 U8564 ( .A1(n6472), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9524) );
  XNOR2_X1 U8565 ( .A(n7575), .B(n8183), .ZN(n11371) );
  NOR2_X1 U8566 ( .A1(n9379), .A2(n7380), .ZN(n7377) );
  XNOR2_X1 U8567 ( .A(n8118), .B(n8117), .ZN(n11033) );
  NAND2_X1 U8568 ( .A1(n8115), .A2(n7648), .ZN(n8137) );
  NAND2_X1 U8569 ( .A1(n6810), .A2(n7681), .ZN(n8026) );
  OAI21_X1 U8570 ( .B1(n7968), .B2(n7967), .A(n6535), .ZN(n7609) );
  AND2_X1 U8571 ( .A1(n9259), .A2(n9273), .ZN(n9857) );
  AND2_X1 U8572 ( .A1(n9158), .A2(n9129), .ZN(n9189) );
  CLKBUF_X1 U8573 ( .A(n9158), .Z(n9159) );
  NAND2_X1 U8574 ( .A1(n6889), .A2(n6928), .ZN(n14372) );
  NAND2_X1 U8575 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n6929), .ZN(n6928) );
  INV_X1 U8576 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6929) );
  INV_X1 U8577 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7333) );
  NAND2_X1 U8578 ( .A1(n14334), .A2(n14333), .ZN(n14387) );
  NAND2_X1 U8579 ( .A1(n14429), .A2(n14398), .ZN(n14400) );
  AND2_X1 U8580 ( .A1(n14598), .A2(n14406), .ZN(n14407) );
  AND2_X1 U8581 ( .A1(n6783), .A2(n14600), .ZN(n14412) );
  AND2_X1 U8582 ( .A1(n11142), .A2(n11143), .ZN(n7256) );
  INV_X1 U8583 ( .A(n15116), .ZN(n10330) );
  NOR2_X1 U8584 ( .A1(n6536), .A2(n6622), .ZN(n6621) );
  AND2_X1 U8585 ( .A1(n11663), .A2(n12483), .ZN(n11664) );
  NAND2_X1 U8586 ( .A1(n11622), .A2(n12122), .ZN(n10196) );
  NAND2_X1 U8587 ( .A1(n15148), .A2(n11643), .ZN(n7074) );
  NAND2_X1 U8588 ( .A1(n12012), .A2(n11640), .ZN(n11924) );
  INV_X1 U8589 ( .A(n11982), .ZN(n6627) );
  NAND2_X1 U8590 ( .A1(n6626), .A2(n11982), .ZN(n6625) );
  INV_X1 U8591 ( .A(n11649), .ZN(n6626) );
  NAND2_X1 U8592 ( .A1(n11650), .A2(n11649), .ZN(n11981) );
  NOR2_X1 U8593 ( .A1(n11934), .A2(n6629), .ZN(n11434) );
  NOR2_X1 U8594 ( .A1(n6630), .A2(n6484), .ZN(n6629) );
  NOR2_X1 U8595 ( .A1(n6854), .A2(n6511), .ZN(n6853) );
  NOR2_X1 U8596 ( .A1(n9010), .A2(n9659), .ZN(n6854) );
  INV_X1 U8597 ( .A(n6879), .ZN(n11128) );
  INV_X1 U8598 ( .A(n12049), .ZN(n6932) );
  NAND2_X1 U8599 ( .A1(n10205), .A2(n10392), .ZN(n12073) );
  NAND2_X1 U8600 ( .A1(n7266), .A2(n7269), .ZN(n12059) );
  OAI211_X1 U8601 ( .C1(n6678), .C2(n12089), .A(n6674), .B(n6464), .ZN(n6673)
         );
  XNOR2_X1 U8602 ( .A(n6988), .B(n12442), .ZN(n6678) );
  INV_X1 U8603 ( .A(n12273), .ZN(n6672) );
  AOI21_X1 U8604 ( .B1(n12463), .B2(n9014), .A(n9000), .ZN(n12472) );
  INV_X1 U8605 ( .A(n12275), .ZN(n12285) );
  OR2_X1 U8606 ( .A1(n10406), .A2(n10412), .ZN(n10443) );
  OAI21_X1 U8607 ( .B1(n10722), .B2(n10469), .A(n7101), .ZN(n10704) );
  AOI21_X1 U8608 ( .B1(n10715), .B2(n10685), .A(n10684), .ZN(n10687) );
  INV_X1 U8609 ( .A(n6665), .ZN(n15055) );
  NOR2_X1 U8610 ( .A1(n10941), .A2(n10940), .ZN(n11067) );
  INV_X1 U8611 ( .A(n7092), .ZN(n10959) );
  INV_X1 U8612 ( .A(n7090), .ZN(n11080) );
  NOR2_X1 U8613 ( .A1(n11420), .A2(n11421), .ZN(n15064) );
  XNOR2_X1 U8614 ( .A(n6930), .B(n11423), .ZN(n11404) );
  NOR2_X1 U8615 ( .A1(n12299), .A2(n12300), .ZN(n15091) );
  INV_X1 U8616 ( .A(n7177), .ZN(n12298) );
  NOR2_X1 U8617 ( .A1(n12308), .A2(n6925), .ZN(n15101) );
  AND2_X1 U8618 ( .A1(n12309), .A2(n7166), .ZN(n6925) );
  INV_X1 U8619 ( .A(n7165), .ZN(n15095) );
  XNOR2_X1 U8620 ( .A(n12371), .B(n12370), .ZN(n14481) );
  INV_X1 U8621 ( .A(n7107), .ZN(n12376) );
  OAI211_X1 U8622 ( .C1(n12384), .C2(n12417), .A(n6636), .B(n6635), .ZN(n12385) );
  NAND2_X1 U8623 ( .A1(n6637), .A2(n12406), .ZN(n6636) );
  NAND2_X1 U8624 ( .A1(n12384), .A2(n6609), .ZN(n6635) );
  OAI21_X1 U8625 ( .B1(n12394), .B2(n12395), .A(n12393), .ZN(n12397) );
  NOR2_X1 U8626 ( .A1(n12397), .A2(n12396), .ZN(n12408) );
  INV_X1 U8627 ( .A(n12438), .ZN(n6934) );
  NAND2_X1 U8628 ( .A1(n6823), .A2(n6826), .ZN(n12494) );
  NAND2_X1 U8629 ( .A1(n7541), .A2(n7542), .ZN(n12511) );
  AND2_X1 U8630 ( .A1(n6829), .A2(n6832), .ZN(n12506) );
  NAND2_X1 U8631 ( .A1(n12519), .A2(n12090), .ZN(n6829) );
  NAND2_X1 U8632 ( .A1(n9053), .A2(n12233), .ZN(n12517) );
  NAND2_X1 U8633 ( .A1(n12535), .A2(n12234), .ZN(n9053) );
  NAND2_X1 U8634 ( .A1(n12541), .A2(n7238), .ZN(n12531) );
  NAND2_X1 U8635 ( .A1(n7548), .A2(n7552), .ZN(n12546) );
  NAND2_X1 U8636 ( .A1(n12571), .A2(n7555), .ZN(n7548) );
  NOR2_X1 U8637 ( .A1(n12555), .A2(n7236), .ZN(n12542) );
  OR3_X1 U8638 ( .A1(n12555), .A2(n12582), .A3(n12554), .ZN(n12559) );
  NAND2_X1 U8639 ( .A1(n7557), .A2(n12218), .ZN(n12561) );
  NAND2_X1 U8640 ( .A1(n7558), .A2(n12219), .ZN(n7557) );
  INV_X1 U8641 ( .A(n12571), .ZN(n7558) );
  NAND2_X1 U8642 ( .A1(n12577), .A2(n6447), .ZN(n12567) );
  NAND2_X1 U8643 ( .A1(n9050), .A2(n12209), .ZN(n12587) );
  NAND2_X1 U8644 ( .A1(n12629), .A2(n12200), .ZN(n12615) );
  NAND2_X1 U8645 ( .A1(n12625), .A2(n12624), .ZN(n12623) );
  NAND2_X1 U8646 ( .A1(n7564), .A2(n12188), .ZN(n12638) );
  NAND2_X1 U8647 ( .A1(n7565), .A2(n12189), .ZN(n7564) );
  INV_X1 U8648 ( .A(n14503), .ZN(n7565) );
  AND2_X1 U8649 ( .A1(n8817), .A2(n8816), .ZN(n11619) );
  INV_X1 U8650 ( .A(n14499), .ZN(n12650) );
  NAND2_X1 U8651 ( .A1(n11229), .A2(n12181), .ZN(n11333) );
  INV_X1 U8652 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15117) );
  INV_X1 U8653 ( .A(n15136), .ZN(n15154) );
  AND2_X1 U8654 ( .A1(n10266), .A2(n15140), .ZN(n15136) );
  NOR2_X1 U8655 ( .A1(n12450), .A2(n12449), .ZN(n14517) );
  NAND2_X1 U8656 ( .A1(n9067), .A2(n9066), .ZN(n9068) );
  AND2_X1 U8657 ( .A1(n12661), .A2(n12660), .ZN(n7631) );
  INV_X1 U8658 ( .A(n12240), .ZN(n12739) );
  INV_X1 U8659 ( .A(n12223), .ZN(n12753) );
  AND2_X1 U8660 ( .A1(n10394), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9713) );
  OAI22_X1 U8661 ( .A1(n11869), .A2(n11868), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n13513), .ZN(n11854) );
  INV_X1 U8662 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n6986) );
  INV_X1 U8663 ( .A(n8585), .ZN(n7073) );
  NAND2_X1 U8664 ( .A1(n9028), .A2(n8583), .ZN(n9077) );
  INV_X1 U8665 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9074) );
  NAND2_X1 U8666 ( .A1(n6666), .A2(n7114), .ZN(n8941) );
  NAND2_X1 U8667 ( .A1(n9100), .A2(n9023), .ZN(n14437) );
  NAND2_X1 U8668 ( .A1(n8897), .A2(n7277), .ZN(n9022) );
  NAND2_X1 U8669 ( .A1(n7118), .A2(n7116), .ZN(n8928) );
  NAND2_X1 U8670 ( .A1(n7118), .A2(n8559), .ZN(n8926) );
  AND2_X1 U8671 ( .A1(n8897), .A2(n7278), .ZN(n9024) );
  NAND2_X1 U8672 ( .A1(n6689), .A2(n8553), .ZN(n8911) );
  NAND2_X1 U8673 ( .A1(n8894), .A2(n8552), .ZN(n6689) );
  OAI21_X1 U8674 ( .B1(n8547), .B2(n8855), .A(n7111), .ZN(n8869) );
  NAND2_X1 U8675 ( .A1(n8547), .A2(n8546), .ZN(n8856) );
  INV_X1 U8676 ( .A(SI_11_), .ZN(n9656) );
  NAND2_X1 U8677 ( .A1(n8785), .A2(n8536), .ZN(n8804) );
  NAND2_X1 U8678 ( .A1(n6688), .A2(n8527), .ZN(n8716) );
  INV_X1 U8679 ( .A(n10657), .ZN(n10956) );
  NAND2_X1 U8680 ( .A1(n8700), .A2(n8699), .ZN(n8701) );
  NAND2_X1 U8681 ( .A1(n8661), .A2(n8517), .ZN(n8673) );
  OAI21_X1 U8682 ( .B1(n10404), .B2(n9027), .A(n8665), .ZN(n6647) );
  NAND2_X1 U8683 ( .A1(n6650), .A2(n6649), .ZN(n6648) );
  INV_X1 U8684 ( .A(n10404), .ZN(n6650) );
  NAND2_X1 U8685 ( .A1(n6707), .A2(n10315), .ZN(n10515) );
  NAND2_X1 U8686 ( .A1(n10062), .A2(n6874), .ZN(n6707) );
  NOR2_X1 U8687 ( .A1(n7384), .A2(n11183), .ZN(n7383) );
  NAND2_X1 U8688 ( .A1(n10827), .A2(n10826), .ZN(n10932) );
  INV_X1 U8689 ( .A(n7400), .ZN(n7399) );
  AOI21_X1 U8690 ( .B1(n7398), .B2(n7400), .A(n7397), .ZN(n7396) );
  INV_X1 U8691 ( .A(n11607), .ZN(n7397) );
  NAND2_X1 U8692 ( .A1(n7930), .A2(n7929), .ZN(n15018) );
  NAND2_X1 U8693 ( .A1(n7170), .A2(n9687), .ZN(n7172) );
  OAI22_X1 U8694 ( .A1(n9654), .A2(n9155), .B1(n9653), .B2(n7171), .ZN(n7170)
         );
  AND2_X1 U8695 ( .A1(n7391), .A2(n6466), .ZN(n12803) );
  INV_X1 U8696 ( .A(n11559), .ZN(n7061) );
  INV_X1 U8697 ( .A(n12840), .ZN(n7389) );
  NAND2_X1 U8698 ( .A1(n11589), .A2(n11588), .ZN(n7390) );
  INV_X1 U8699 ( .A(n7384), .ZN(n7382) );
  NAND2_X1 U8700 ( .A1(n6703), .A2(n6449), .ZN(n12863) );
  INV_X1 U8701 ( .A(n12862), .ZN(n6703) );
  XNOR2_X1 U8702 ( .A(n15027), .B(n11592), .ZN(n10829) );
  INV_X1 U8703 ( .A(n9916), .ZN(n9915) );
  NOR2_X1 U8704 ( .A1(n12827), .A2(n7069), .ZN(n12874) );
  NAND2_X1 U8705 ( .A1(n10062), .A2(n10061), .ZN(n10308) );
  NAND2_X1 U8706 ( .A1(n14882), .A2(n9897), .ZN(n9899) );
  NOR2_X1 U8707 ( .A1(n14928), .A2(n6712), .ZN(n14941) );
  NOR2_X1 U8708 ( .A1(n6714), .A2(n6713), .ZN(n6712) );
  AND2_X1 U8709 ( .A1(n6720), .A2(n6490), .ZN(n14962) );
  AND2_X1 U8710 ( .A1(n14978), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n14981) );
  XNOR2_X1 U8711 ( .A(n6718), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n12979) );
  NOR2_X1 U8712 ( .A1(n14981), .A2(n12976), .ZN(n6718) );
  NAND2_X1 U8713 ( .A1(n8384), .A2(n8383), .ZN(n13237) );
  INV_X1 U8714 ( .A(n11699), .ZN(n11700) );
  AOI22_X1 U8715 ( .A1(n13011), .A2(n13225), .B1(n12985), .B2(n12904), .ZN(
        n11699) );
  NAND2_X1 U8716 ( .A1(n7280), .A2(n7285), .ZN(n13000) );
  NAND2_X1 U8717 ( .A1(n13026), .A2(n7286), .ZN(n7280) );
  NAND2_X1 U8718 ( .A1(n7343), .A2(n7347), .ZN(n12997) );
  NAND2_X1 U8719 ( .A1(n13035), .A2(n7348), .ZN(n7343) );
  NAND2_X1 U8720 ( .A1(n7350), .A2(n7348), .ZN(n13014) );
  NAND2_X1 U8721 ( .A1(n6904), .A2(n6903), .ZN(n7350) );
  INV_X1 U8722 ( .A(n7029), .ZN(n7028) );
  XNOR2_X1 U8723 ( .A(n7031), .B(n13013), .ZN(n7030) );
  AOI22_X1 U8724 ( .A1(n13011), .A2(n13223), .B1(n13225), .B2(n13012), .ZN(
        n7029) );
  NAND2_X1 U8725 ( .A1(n7334), .A2(n7337), .ZN(n13038) );
  NAND2_X1 U8726 ( .A1(n13080), .A2(n7338), .ZN(n7334) );
  AND2_X1 U8727 ( .A1(n7302), .A2(n7301), .ZN(n13058) );
  NAND2_X1 U8728 ( .A1(n7020), .A2(n7018), .ZN(n13124) );
  NAND2_X1 U8729 ( .A1(n7025), .A2(n11688), .ZN(n13134) );
  NAND2_X1 U8730 ( .A1(n7026), .A2(n6475), .ZN(n7025) );
  NAND2_X1 U8731 ( .A1(n7356), .A2(n11713), .ZN(n13151) );
  NAND2_X1 U8732 ( .A1(n8093), .A2(n8092), .ZN(n13189) );
  NAND2_X1 U8733 ( .A1(n8053), .A2(n8052), .ZN(n13323) );
  NAND2_X1 U8734 ( .A1(n7313), .A2(n11362), .ZN(n11677) );
  NAND2_X1 U8735 ( .A1(n11359), .A2(n11358), .ZN(n7313) );
  NAND2_X1 U8736 ( .A1(n10911), .A2(n10912), .ZN(n10910) );
  NAND2_X1 U8737 ( .A1(n10868), .A2(n10867), .ZN(n10911) );
  NAND2_X1 U8738 ( .A1(n6743), .A2(n6744), .ZN(n10553) );
  NAND2_X1 U8739 ( .A1(n7309), .A2(n10007), .ZN(n10127) );
  INV_X1 U8740 ( .A(n7807), .ZN(n10372) );
  INV_X1 U8741 ( .A(n10168), .ZN(n10362) );
  NAND2_X1 U8742 ( .A1(n14998), .A2(n9734), .ZN(n13217) );
  AND2_X1 U8743 ( .A1(n13219), .A2(n10090), .ZN(n13234) );
  OR2_X1 U8744 ( .A1(n13263), .A2(n13327), .ZN(n6909) );
  AOI21_X1 U8745 ( .B1(n10370), .B2(n13291), .A(n6937), .ZN(n10041) );
  INV_X1 U8746 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n7741) );
  INV_X1 U8747 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n7739) );
  INV_X1 U8748 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11373) );
  INV_X1 U8749 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10820) );
  AND2_X1 U8750 ( .A1(n7718), .A2(n8493), .ZN(n12974) );
  INV_X1 U8751 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10804) );
  INV_X1 U8752 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10510) );
  INV_X1 U8753 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10060) );
  INV_X1 U8754 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9930) );
  INV_X1 U8755 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9769) );
  INV_X1 U8756 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9684) );
  INV_X1 U8757 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9679) );
  INV_X1 U8758 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9671) );
  INV_X1 U8759 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9667) );
  INV_X1 U8760 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9652) );
  INV_X1 U8761 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9647) );
  INV_X1 U8762 ( .A(n7841), .ZN(n7822) );
  INV_X1 U8763 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9649) );
  NAND2_X1 U8764 ( .A1(n10740), .A2(n6528), .ZN(n10746) );
  NAND2_X1 U8765 ( .A1(n10746), .A2(n10745), .ZN(n10847) );
  NAND2_X1 U8766 ( .A1(n11742), .A2(n11741), .ZN(n15378) );
  NAND2_X1 U8767 ( .A1(n13463), .A2(n11799), .ZN(n13381) );
  NAND2_X1 U8768 ( .A1(n13473), .A2(n11776), .ZN(n13400) );
  NOR2_X1 U8769 ( .A1(n7485), .A2(n7483), .ZN(n7480) );
  NAND2_X1 U8770 ( .A1(n7482), .A2(n11842), .ZN(n7481) );
  NAND2_X1 U8771 ( .A1(n13454), .A2(n7636), .ZN(n13409) );
  NAND2_X1 U8772 ( .A1(n6974), .A2(n7488), .ZN(n14549) );
  NOR2_X1 U8773 ( .A1(n14558), .A2(n11476), .ZN(n14551) );
  NAND2_X1 U8774 ( .A1(n6723), .A2(n7472), .ZN(n13417) );
  NAND2_X1 U8775 ( .A1(n13381), .A2(n7474), .ZN(n6723) );
  NOR2_X1 U8776 ( .A1(n7456), .A2(n10526), .ZN(n10547) );
  NAND2_X1 U8777 ( .A1(n9369), .A2(n9368), .ZN(n14235) );
  NAND2_X1 U8778 ( .A1(n7473), .A2(n11806), .ZN(n13446) );
  NAND2_X1 U8779 ( .A1(n13381), .A2(n13382), .ZN(n7473) );
  NAND2_X1 U8780 ( .A1(n13401), .A2(n7646), .ZN(n13456) );
  OR2_X1 U8781 ( .A1(n11784), .A2(n11783), .ZN(n7646) );
  NAND2_X1 U8782 ( .A1(n13456), .A2(n13455), .ZN(n13454) );
  NAND2_X1 U8783 ( .A1(n6974), .A2(n6898), .ZN(n11742) );
  NOR2_X1 U8784 ( .A1(n7486), .A2(n6975), .ZN(n6898) );
  INV_X1 U8785 ( .A(n11484), .ZN(n6975) );
  NOR2_X1 U8786 ( .A1(n7487), .A2(n7486), .ZN(n11485) );
  NAND2_X1 U8787 ( .A1(n6734), .A2(n6520), .ZN(n14559) );
  NAND2_X1 U8788 ( .A1(n11463), .A2(n6972), .ZN(n6734) );
  NOR2_X1 U8789 ( .A1(n14559), .A2(n14560), .ZN(n14558) );
  INV_X1 U8790 ( .A(n15388), .ZN(n14566) );
  NAND2_X1 U8791 ( .A1(n7458), .A2(n6735), .ZN(n10740) );
  AND2_X1 U8792 ( .A1(n10549), .A2(n7457), .ZN(n6735) );
  NAND2_X1 U8793 ( .A1(n11755), .A2(n6736), .ZN(n13494) );
  NAND2_X1 U8794 ( .A1(n6869), .A2(n6868), .ZN(n6867) );
  INV_X1 U8795 ( .A(n13762), .ZN(n6868) );
  INV_X1 U8796 ( .A(n13761), .ZN(n6869) );
  OR2_X1 U8797 ( .A1(n9376), .A2(n9375), .ZN(n13783) );
  NAND2_X1 U8798 ( .A1(n13503), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9188) );
  OR2_X1 U8799 ( .A1(n13505), .A2(n9809), .ZN(n9176) );
  CLKBUF_X1 U8800 ( .A(n9981), .Z(n14728) );
  OR2_X1 U8801 ( .A1(n13506), .A2(n9165), .ZN(n9168) );
  AOI21_X1 U8802 ( .B1(n6448), .B2(n13980), .A(n6517), .ZN(n7414) );
  NAND2_X1 U8803 ( .A1(n7141), .A2(n14730), .ZN(n7140) );
  NAND2_X1 U8804 ( .A1(n13982), .A2(n7142), .ZN(n7141) );
  NAND2_X1 U8805 ( .A1(n14027), .A2(n9460), .ZN(n14015) );
  AND2_X1 U8806 ( .A1(n14034), .A2(n9549), .ZN(n14013) );
  NAND2_X1 U8807 ( .A1(n7201), .A2(n7204), .ZN(n14060) );
  NAND2_X1 U8808 ( .A1(n14090), .A2(n7205), .ZN(n7201) );
  NAND2_X1 U8809 ( .A1(n7439), .A2(n7444), .ZN(n14074) );
  NAND2_X1 U8810 ( .A1(n14106), .A2(n7447), .ZN(n7439) );
  NAND2_X1 U8811 ( .A1(n7449), .A2(n7447), .ZN(n14101) );
  NAND2_X1 U8812 ( .A1(n7449), .A2(n7446), .ZN(n14099) );
  AND2_X1 U8813 ( .A1(n14093), .A2(n14092), .ZN(n14216) );
  INV_X1 U8814 ( .A(n14230), .ZN(n14132) );
  NAND2_X1 U8815 ( .A1(n11532), .A2(n9545), .ZN(n14135) );
  NAND2_X1 U8816 ( .A1(n9344), .A2(n9343), .ZN(n14248) );
  NAND2_X1 U8817 ( .A1(n11501), .A2(n9542), .ZN(n11516) );
  NAND2_X1 U8818 ( .A1(n11495), .A2(n13644), .ZN(n11494) );
  NAND2_X1 U8819 ( .A1(n14447), .A2(n9327), .ZN(n11495) );
  NAND2_X1 U8820 ( .A1(n11325), .A2(n13532), .ZN(n11324) );
  NAND2_X1 U8821 ( .A1(n11340), .A2(n9540), .ZN(n11325) );
  NAND2_X1 U8822 ( .A1(n10789), .A2(n9256), .ZN(n14682) );
  NAND2_X1 U8823 ( .A1(n7438), .A2(n9535), .ZN(n10788) );
  NAND2_X1 U8824 ( .A1(n10757), .A2(n9534), .ZN(n7438) );
  NAND2_X1 U8825 ( .A1(n10504), .A2(n9531), .ZN(n10589) );
  INV_X1 U8826 ( .A(n14739), .ZN(n14694) );
  OR2_X1 U8827 ( .A1(n14746), .A2(n14453), .ZN(n14739) );
  NOR2_X1 U8828 ( .A1(n14710), .A2(n14704), .ZN(n14118) );
  NAND2_X1 U8829 ( .A1(n13516), .A2(n13515), .ZN(n14155) );
  NAND2_X1 U8830 ( .A1(n14808), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7152) );
  NAND2_X1 U8831 ( .A1(n6488), .A2(n14153), .ZN(n14258) );
  NAND2_X1 U8832 ( .A1(n9448), .A2(n9447), .ZN(n14272) );
  NAND2_X1 U8833 ( .A1(n14321), .A2(n9429), .ZN(n14281) );
  NAND2_X1 U8834 ( .A1(n9401), .A2(n9400), .ZN(n14290) );
  NAND2_X1 U8835 ( .A1(n13511), .A2(n9629), .ZN(n6614) );
  INV_X1 U8836 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14296) );
  NOR2_X1 U8837 ( .A1(n7453), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n7452) );
  NAND2_X1 U8838 ( .A1(n7454), .A2(n9142), .ZN(n7453) );
  INV_X1 U8839 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9142) );
  XNOR2_X1 U8841 ( .A(n9579), .B(n9578), .ZN(n14309) );
  XNOR2_X1 U8842 ( .A(n9576), .B(n9575), .ZN(n14310) );
  XNOR2_X1 U8843 ( .A(n6802), .B(n8560), .ZN(n14321) );
  NOR2_X1 U8844 ( .A1(n9428), .A2(n7171), .ZN(n6802) );
  INV_X1 U8845 ( .A(n13553), .ZN(n14320) );
  XNOR2_X1 U8846 ( .A(n9523), .B(n9522), .ZN(n13548) );
  AND2_X1 U8847 ( .A1(n7502), .A2(n7501), .ZN(n7500) );
  INV_X1 U8848 ( .A(n13550), .ZN(n9590) );
  INV_X1 U8849 ( .A(n14082), .ZN(n13929) );
  INV_X1 U8850 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11034) );
  INV_X1 U8851 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10819) );
  INV_X1 U8852 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10803) );
  INV_X1 U8853 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10756) );
  INV_X1 U8854 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9770) );
  INV_X1 U8855 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9682) );
  INV_X1 U8856 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9677) );
  INV_X1 U8857 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9673) );
  NAND2_X1 U8858 ( .A1(n7903), .A2(n7902), .ZN(n9672) );
  INV_X1 U8859 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9669) );
  INV_X1 U8860 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7653) );
  INV_X1 U8861 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14375) );
  NOR2_X1 U8862 ( .A1(n15408), .A2(n14379), .ZN(n14423) );
  XNOR2_X1 U8863 ( .A(n14382), .B(n7319), .ZN(n15399) );
  NAND2_X1 U8864 ( .A1(n15399), .A2(n12931), .ZN(n15398) );
  XNOR2_X1 U8865 ( .A(n14386), .B(n14385), .ZN(n14428) );
  NOR2_X1 U8866 ( .A1(n14428), .A2(n14427), .ZN(n14426) );
  INV_X1 U8867 ( .A(n14397), .ZN(n7325) );
  XNOR2_X1 U8868 ( .A(n14400), .B(n14399), .ZN(n14432) );
  XNOR2_X1 U8869 ( .A(n14405), .B(n7326), .ZN(n14599) );
  INV_X1 U8870 ( .A(n14404), .ZN(n7326) );
  NAND2_X1 U8871 ( .A1(n14599), .A2(n14923), .ZN(n14598) );
  NAND2_X1 U8872 ( .A1(n14407), .A2(n14408), .ZN(n14602) );
  NAND2_X1 U8873 ( .A1(n14602), .A2(n14935), .ZN(n14600) );
  NOR2_X1 U8874 ( .A1(n14412), .A2(n14411), .ZN(n14604) );
  NAND2_X1 U8875 ( .A1(n14412), .A2(n14411), .ZN(n14606) );
  OAI21_X1 U8876 ( .B1(n6769), .B2(n6770), .A(n14974), .ZN(n7318) );
  NAND2_X1 U8877 ( .A1(n6772), .A2(n6771), .ZN(n6770) );
  INV_X1 U8878 ( .A(n14607), .ZN(n6769) );
  INV_X1 U8879 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n14476) );
  NAND2_X1 U8880 ( .A1(n7088), .A2(n11620), .ZN(n7087) );
  INV_X1 U8881 ( .A(n11621), .ZN(n7088) );
  OAI21_X1 U8882 ( .B1(n12424), .B2(n15097), .A(n7178), .ZN(P3_U3200) );
  AND2_X1 U8883 ( .A1(n7180), .A2(n7179), .ZN(n7178) );
  OAI21_X1 U8884 ( .B1(n12430), .B2(n6463), .A(n15089), .ZN(n7180) );
  XNOR2_X1 U8885 ( .A(n7102), .B(n12436), .ZN(n12446) );
  INV_X1 U8886 ( .A(n7570), .ZN(n7569) );
  OAI21_X1 U8887 ( .B1(n11864), .B2(n12653), .A(n7571), .ZN(n7570) );
  AOI21_X1 U8888 ( .B1(n11866), .B2(n14499), .A(n11865), .ZN(n7571) );
  NAND2_X1 U8889 ( .A1(n6846), .A2(n6844), .ZN(P3_U3486) );
  INV_X1 U8890 ( .A(n6845), .ZN(n6844) );
  OR2_X1 U8891 ( .A1(n12729), .A2(n15219), .ZN(n6846) );
  OAI22_X1 U8892 ( .A1(n12731), .A2(n12722), .B1(n15222), .B2(n12667), .ZN(
        n6845) );
  NAND2_X1 U8893 ( .A1(n9056), .A2(n6842), .ZN(n6841) );
  OAI21_X1 U8894 ( .B1(n12729), .B2(n15205), .A(n6839), .ZN(P3_U3454) );
  INV_X1 U8895 ( .A(n6840), .ZN(n6839) );
  OAI22_X1 U8896 ( .A1(n12731), .A2(n12776), .B1(n15206), .B2(n12730), .ZN(
        n6840) );
  NAND2_X1 U8897 ( .A1(n9056), .A2(n12723), .ZN(n6843) );
  INV_X1 U8898 ( .A(n6872), .ZN(n6871) );
  OAI21_X1 U8899 ( .B1(n6945), .B2(n12883), .A(n12783), .ZN(n6872) );
  NAND2_X1 U8900 ( .A1(n7391), .A2(n7392), .ZN(n12858) );
  INV_X1 U8901 ( .A(n7060), .ZN(n11560) );
  NAND2_X1 U8902 ( .A1(n7506), .A2(n7504), .ZN(n8510) );
  AOI21_X1 U8903 ( .B1(n8509), .B2(n8503), .A(n8502), .ZN(n8511) );
  AND2_X1 U8904 ( .A1(n6908), .A2(n6907), .ZN(n13037) );
  AOI21_X1 U8905 ( .B1(n13260), .B2(n13131), .A(n13036), .ZN(n6907) );
  OR2_X1 U8906 ( .A1(n13263), .A2(n13236), .ZN(n6908) );
  INV_X1 U8907 ( .A(n9709), .ZN(n9618) );
  NAND2_X1 U8908 ( .A1(n6981), .A2(n14564), .ZN(n6979) );
  OAI21_X1 U8909 ( .B1(n6886), .B2(n15379), .A(n13491), .ZN(P1_U3240) );
  XNOR2_X1 U8910 ( .A(n13484), .B(n6887), .ZN(n6886) );
  OAI21_X1 U8911 ( .B1(n9612), .B2(n9605), .A(n9606), .ZN(n6962) );
  OR2_X1 U8912 ( .A1(n14822), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6860) );
  NAND2_X1 U8913 ( .A1(n7153), .A2(n7150), .ZN(P1_U3526) );
  INV_X1 U8914 ( .A(n7151), .ZN(n7150) );
  NAND2_X1 U8915 ( .A1(n14258), .A2(n14810), .ZN(n7153) );
  OAI21_X1 U8916 ( .B1(n14260), .B2(n14282), .A(n7152), .ZN(n7151) );
  OR2_X1 U8917 ( .A1(n14810), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6862) );
  INV_X1 U8918 ( .A(n7321), .ZN(n15395) );
  NOR2_X1 U8919 ( .A1(n14439), .A2(n14440), .ZN(n14438) );
  INV_X1 U8920 ( .A(n7330), .ZN(n14596) );
  INV_X1 U8921 ( .A(n7327), .ZN(n14594) );
  XNOR2_X1 U8922 ( .A(n14479), .B(n14478), .ZN(n7322) );
  AND2_X1 U8923 ( .A1(n6465), .A2(n8909), .ZN(n6447) );
  AND2_X1 U8924 ( .A1(n13967), .A2(n9553), .ZN(n6448) );
  NAND2_X1 U8925 ( .A1(n6941), .A2(n11730), .ZN(n13229) );
  AND2_X1 U8926 ( .A1(n13105), .A2(n13194), .ZN(n6449) );
  INV_X1 U8927 ( .A(n13618), .ZN(n7148) );
  AND2_X1 U8928 ( .A1(n7586), .A2(n8143), .ZN(n6450) );
  OR2_X1 U8929 ( .A1(n7424), .A2(n7427), .ZN(n6451) );
  NOR2_X1 U8930 ( .A1(n11689), .A2(n7024), .ZN(n7023) );
  INV_X1 U8931 ( .A(n13535), .ZN(n7420) );
  INV_X1 U8932 ( .A(n13532), .ZN(n7409) );
  AND2_X1 U8933 ( .A1(n7678), .A2(n9656), .ZN(n6452) );
  NAND2_X1 U8934 ( .A1(n8637), .A2(n8636), .ZN(n12223) );
  INV_X1 U8935 ( .A(n14105), .ZN(n7450) );
  MUX2_X1 U8936 ( .A(n9694), .B(n13374), .S(n9687), .Z(n10010) );
  OR2_X1 U8937 ( .A1(n8773), .A2(n11154), .ZN(n6453) );
  NOR2_X1 U8938 ( .A1(n13259), .A2(n13043), .ZN(n6454) );
  INV_X1 U8939 ( .A(n10350), .ZN(n6939) );
  INV_X1 U8940 ( .A(n12640), .ZN(n7221) );
  NAND2_X2 U8941 ( .A1(n9031), .A2(n12437), .ZN(n10395) );
  AND2_X1 U8942 ( .A1(n6946), .A2(n6945), .ZN(n6455) );
  AND2_X1 U8943 ( .A1(n11825), .A2(n11824), .ZN(n6456) );
  AND2_X1 U8944 ( .A1(n13255), .A2(n12891), .ZN(n6457) );
  AND2_X1 U8945 ( .A1(n13590), .A2(n10588), .ZN(n6458) );
  AND2_X1 U8946 ( .A1(n13269), .A2(n13074), .ZN(n6459) );
  AND2_X1 U8947 ( .A1(n7491), .A2(n7494), .ZN(n6460) );
  INV_X1 U8948 ( .A(n12999), .ZN(n7282) );
  AND2_X1 U8949 ( .A1(n7171), .A2(SI_1_), .ZN(n6461) );
  INV_X1 U8950 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9156) );
  NAND2_X1 U8951 ( .A1(n8324), .A2(n8323), .ZN(n13250) );
  XNOR2_X1 U8952 ( .A(n14165), .B(n13773), .ZN(n13980) );
  INV_X1 U8953 ( .A(n11712), .ZN(n13167) );
  AND2_X1 U8954 ( .A1(n8157), .A2(n8156), .ZN(n6462) );
  INV_X1 U8955 ( .A(n12477), .ZN(n12731) );
  NAND2_X1 U8956 ( .A1(n8587), .A2(n8586), .ZN(n12477) );
  INV_X1 U8957 ( .A(n12096), .ZN(n7225) );
  NAND2_X1 U8958 ( .A1(n9511), .A2(n9510), .ZN(n13735) );
  AND2_X1 U8959 ( .A1(n12421), .A2(n12420), .ZN(n6463) );
  OR2_X1 U8960 ( .A1(n12109), .A2(n12108), .ZN(n6464) );
  INV_X1 U8961 ( .A(n7667), .ZN(n7576) );
  NAND2_X1 U8962 ( .A1(n7143), .A2(SI_6_), .ZN(n7667) );
  NAND2_X1 U8963 ( .A1(n12218), .A2(n12219), .ZN(n6465) );
  NAND2_X1 U8964 ( .A1(n8930), .A2(n8929), .ZN(n12037) );
  AND2_X1 U8965 ( .A1(n7392), .A2(n6559), .ZN(n6466) );
  AND2_X1 U8966 ( .A1(n7898), .A2(n7897), .ZN(n6467) );
  XNOR2_X1 U8967 ( .A(n9755), .B(n10168), .ZN(n10160) );
  AND2_X1 U8968 ( .A1(n7522), .A2(n7314), .ZN(n6468) );
  OR2_X1 U8969 ( .A1(n14078), .A2(n9427), .ZN(n7204) );
  INV_X1 U8970 ( .A(n13778), .ZN(n7138) );
  INV_X1 U8971 ( .A(n13298), .ZN(n7027) );
  AND4_X1 U8972 ( .A1(n8574), .A2(n8575), .A3(n8573), .A4(n8702), .ZN(n6469)
         );
  INV_X1 U8973 ( .A(n12580), .ZN(n8907) );
  AND2_X1 U8974 ( .A1(n12206), .A2(n12211), .ZN(n12580) );
  NAND2_X1 U8975 ( .A1(n8221), .A2(n8220), .ZN(n13105) );
  INV_X1 U8976 ( .A(n9056), .ZN(n12735) );
  NAND2_X1 U8977 ( .A1(n8979), .A2(n8978), .ZN(n9056) );
  NAND2_X1 U8978 ( .A1(n9316), .A2(n9315), .ZN(n13638) );
  INV_X1 U8979 ( .A(n13638), .ZN(n6616) );
  INV_X1 U8980 ( .A(n14553), .ZN(n7146) );
  NAND2_X1 U8981 ( .A1(n7148), .A2(n7147), .ZN(n6470) );
  INV_X1 U8982 ( .A(n6944), .ZN(n6941) );
  OR2_X1 U8983 ( .A1(n12339), .A2(n6607), .ZN(n6471) );
  AND2_X1 U8984 ( .A1(n12553), .A2(n12552), .ZN(n12555) );
  NAND2_X1 U8985 ( .A1(n7686), .A2(n7630), .ZN(n7626) );
  NAND2_X1 U8986 ( .A1(n7426), .A2(n7375), .ZN(n6472) );
  INV_X1 U8987 ( .A(n7815), .ZN(n8429) );
  INV_X1 U8988 ( .A(n12182), .ZN(n7566) );
  AND2_X1 U8989 ( .A1(n9556), .A2(n13564), .ZN(n6473) );
  INV_X1 U8990 ( .A(n13530), .ZN(n7406) );
  NAND2_X1 U8991 ( .A1(n9687), .A2(n7171), .ZN(n7904) );
  NAND2_X1 U8992 ( .A1(n12872), .A2(n7393), .ZN(n7391) );
  INV_X1 U8993 ( .A(n13056), .ZN(n7340) );
  NAND2_X1 U8994 ( .A1(n8955), .A2(n8954), .ZN(n12676) );
  NAND2_X1 U8995 ( .A1(n12082), .A2(n12081), .ZN(n12724) );
  NAND4_X1 U8996 ( .A1(n7768), .A2(n7767), .A3(n7766), .A4(n7765), .ZN(n8459)
         );
  XNOR2_X1 U8997 ( .A(n12916), .B(n7807), .ZN(n10036) );
  OR2_X1 U8998 ( .A1(n12340), .A2(n6471), .ZN(n6474) );
  OR2_X1 U8999 ( .A1(n13302), .A2(n13138), .ZN(n6475) );
  AND2_X1 U9000 ( .A1(n7128), .A2(SI_10_), .ZN(n6476) );
  NAND2_X1 U9001 ( .A1(n8839), .A2(n8838), .ZN(n8547) );
  AND2_X1 U9002 ( .A1(n14215), .A2(n13780), .ZN(n6477) );
  AND2_X1 U9003 ( .A1(n8084), .A2(n8083), .ZN(n6478) );
  NAND2_X1 U9004 ( .A1(n14004), .A2(n7155), .ZN(n6479) );
  AOI21_X1 U9005 ( .B1(n7510), .B2(n7509), .A(n7508), .ZN(n7507) );
  OR2_X1 U9006 ( .A1(n15053), .A2(n10957), .ZN(n6480) );
  AND4_X1 U9007 ( .A1(n9139), .A2(n9138), .A3(n9137), .A4(n9136), .ZN(n6481)
         );
  NAND2_X1 U9008 ( .A1(n13590), .A2(n13795), .ZN(n6482) );
  AND2_X1 U9009 ( .A1(n6618), .A2(n11645), .ZN(n6483) );
  XOR2_X1 U9010 ( .A(n11622), .B(n14529), .Z(n6484) );
  AND2_X1 U9011 ( .A1(n12020), .A2(n12025), .ZN(n6485) );
  INV_X1 U9012 ( .A(n10395), .ZN(n8653) );
  AND2_X1 U9013 ( .A1(n8643), .A2(n7076), .ZN(n6486) );
  AND2_X1 U9014 ( .A1(n7272), .A2(n7085), .ZN(n6487) );
  OR3_X1 U9015 ( .A1(n13943), .A2(n13944), .A3(n14788), .ZN(n6488) );
  NAND4_X1 U9016 ( .A1(n9179), .A2(n9178), .A3(n9177), .A4(n9176), .ZN(n13798)
         );
  NAND2_X1 U9017 ( .A1(n9355), .A2(n9354), .ZN(n13657) );
  OR2_X1 U9018 ( .A1(n12417), .A2(n12416), .ZN(n6489) );
  INV_X1 U9019 ( .A(n13519), .ZN(n7195) );
  NAND2_X1 U9020 ( .A1(n9493), .A2(n9492), .ZN(n13968) );
  INV_X1 U9021 ( .A(n13968), .ZN(n14263) );
  NAND4_X1 U9022 ( .A1(n9147), .A2(n9146), .A3(n7402), .A4(n9152), .ZN(n9981)
         );
  INV_X1 U9023 ( .A(n9981), .ZN(n9173) );
  INV_X1 U9024 ( .A(n15124), .ZN(n7212) );
  OR2_X1 U9025 ( .A1(n11287), .A2(n11306), .ZN(n6490) );
  NAND2_X1 U9026 ( .A1(n7970), .A2(n7969), .ZN(n9271) );
  AND2_X1 U9027 ( .A1(n14235), .A2(n13783), .ZN(n6491) );
  AND3_X1 U9028 ( .A1(n13644), .A2(n13643), .A3(n13642), .ZN(n6492) );
  AND2_X1 U9029 ( .A1(n15018), .A2(n12910), .ZN(n6493) );
  AND2_X1 U9030 ( .A1(n11886), .A2(n7267), .ZN(n6494) );
  NAND2_X1 U9031 ( .A1(n8299), .A2(n8298), .ZN(n13266) );
  AND2_X1 U9032 ( .A1(n12666), .A2(n15203), .ZN(n6495) );
  OR2_X1 U9033 ( .A1(n14473), .A2(n14474), .ZN(n6496) );
  INV_X1 U9034 ( .A(n7021), .ZN(n7019) );
  AOI21_X1 U9035 ( .B1(n7022), .B2(n7023), .A(n6547), .ZN(n7021) );
  NOR2_X1 U9036 ( .A1(n12162), .A2(n8773), .ZN(n6497) );
  AND2_X1 U9037 ( .A1(n14165), .A2(n13488), .ZN(n6498) );
  NAND2_X1 U9038 ( .A1(n8148), .A2(n8147), .ZN(n13298) );
  NAND4_X1 U9039 ( .A1(n8684), .A2(n8683), .A3(n8682), .A4(n8681), .ZN(n15108)
         );
  NAND2_X1 U9040 ( .A1(n9475), .A2(n9474), .ZN(n14171) );
  NAND4_X1 U9041 ( .A1(n8671), .A2(n8670), .A3(n8669), .A4(n8668), .ZN(n15123)
         );
  INV_X1 U9042 ( .A(n11842), .ZN(n7485) );
  AND2_X1 U9043 ( .A1(n12676), .A2(n12521), .ZN(n6499) );
  AND2_X1 U9044 ( .A1(n6619), .A2(n6870), .ZN(n6500) );
  NAND2_X1 U9045 ( .A1(n7597), .A2(n8210), .ZN(n8250) );
  AND2_X1 U9046 ( .A1(n10380), .A2(n6939), .ZN(n6501) );
  AND2_X1 U9047 ( .A1(n7919), .A2(n7918), .ZN(n6502) );
  INV_X1 U9048 ( .A(n7475), .ZN(n7474) );
  OAI21_X1 U9049 ( .B1(n13382), .B2(n7476), .A(n13447), .ZN(n7475) );
  NOR2_X1 U9050 ( .A1(n10860), .A2(n10411), .ZN(n6503) );
  AND2_X1 U9051 ( .A1(n8447), .A2(n8446), .ZN(n6504) );
  AND2_X1 U9052 ( .A1(n8243), .A2(n8242), .ZN(n6505) );
  NOR2_X1 U9053 ( .A1(n11925), .A2(n7275), .ZN(n6506) );
  NOR2_X1 U9054 ( .A1(n11250), .A2(n11242), .ZN(n6507) );
  NOR2_X1 U9055 ( .A1(n14550), .A2(n14560), .ZN(n6508) );
  INV_X1 U9056 ( .A(n7159), .ZN(n14048) );
  INV_X1 U9057 ( .A(n7520), .ZN(n7519) );
  NOR2_X1 U9058 ( .A1(n8159), .A2(n6462), .ZN(n7520) );
  NOR2_X1 U9059 ( .A1(n14235), .A2(n9378), .ZN(n6509) );
  AND2_X1 U9060 ( .A1(n7566), .A2(n12181), .ZN(n6510) );
  NAND2_X1 U9061 ( .A1(n7788), .A2(n7698), .ZN(n7799) );
  AND2_X1 U9062 ( .A1(n8653), .A2(n10722), .ZN(n6511) );
  INV_X1 U9063 ( .A(n7013), .ZN(n7012) );
  NAND2_X1 U9064 ( .A1(n12580), .A2(n12209), .ZN(n7013) );
  AND2_X1 U9065 ( .A1(n7083), .A2(n7270), .ZN(n6512) );
  NAND2_X1 U9066 ( .A1(n11480), .A2(n11479), .ZN(n6513) );
  AND2_X1 U9067 ( .A1(n11136), .A2(n12282), .ZN(n6514) );
  AND2_X1 U9068 ( .A1(n11745), .A2(n11741), .ZN(n6515) );
  OR2_X1 U9069 ( .A1(n8043), .A2(n8042), .ZN(n6516) );
  AND2_X1 U9070 ( .A1(n13968), .A2(n9506), .ZN(n6517) );
  AND2_X1 U9071 ( .A1(n13266), .A2(n13060), .ZN(n6518) );
  AND2_X1 U9072 ( .A1(n7277), .A2(n7276), .ZN(n6519) );
  INV_X1 U9073 ( .A(n7070), .ZN(n7069) );
  OR2_X1 U9074 ( .A1(n11467), .A2(n11466), .ZN(n6520) );
  OR2_X1 U9075 ( .A1(n7362), .A2(n13703), .ZN(n6521) );
  INV_X1 U9076 ( .A(n7339), .ZN(n7338) );
  AND2_X1 U9077 ( .A1(n8110), .A2(n8109), .ZN(n6522) );
  AND2_X1 U9078 ( .A1(n11818), .A2(n11817), .ZN(n6523) );
  AND2_X1 U9079 ( .A1(n13454), .A2(n7498), .ZN(n6524) );
  INV_X1 U9080 ( .A(n7290), .ZN(n7289) );
  NOR2_X1 U9081 ( .A1(n13033), .A2(n13012), .ZN(n7290) );
  AND2_X1 U9082 ( .A1(n10129), .A2(n10128), .ZN(n6525) );
  AND2_X1 U9083 ( .A1(n11834), .A2(n11833), .ZN(n6526) );
  INV_X1 U9084 ( .A(n7967), .ZN(n7613) );
  NOR2_X1 U9085 ( .A1(n13302), .A2(n13165), .ZN(n6527) );
  OR2_X1 U9086 ( .A1(n10741), .A2(n10742), .ZN(n6528) );
  NOR2_X1 U9087 ( .A1(n11812), .A2(n11811), .ZN(n6529) );
  NOR2_X1 U9088 ( .A1(n14553), .A2(n13788), .ZN(n6530) );
  NOR2_X1 U9089 ( .A1(n13266), .A2(n13060), .ZN(n6531) );
  INV_X1 U9090 ( .A(n7206), .ZN(n7205) );
  NAND2_X1 U9091 ( .A1(n9414), .A2(n7207), .ZN(n7206) );
  AND2_X1 U9092 ( .A1(n7827), .A2(n7660), .ZN(n6532) );
  AND2_X1 U9093 ( .A1(n7984), .A2(n7983), .ZN(n6533) );
  NOR2_X1 U9094 ( .A1(n12739), .A2(n12484), .ZN(n6534) );
  AND2_X1 U9095 ( .A1(n7676), .A2(n7612), .ZN(n6535) );
  INV_X1 U9096 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6709) );
  OR2_X1 U9097 ( .A1(n11972), .A2(n11630), .ZN(n6536) );
  AND2_X1 U9098 ( .A1(n13255), .A2(n13027), .ZN(n6537) );
  AND2_X1 U9099 ( .A1(n7020), .A2(n7021), .ZN(n6538) );
  NAND2_X1 U9100 ( .A1(n9383), .A2(n7500), .ZN(n6539) );
  AND2_X1 U9101 ( .A1(n11657), .A2(n12497), .ZN(n6540) );
  AND2_X1 U9102 ( .A1(n7188), .A2(n6957), .ZN(n6541) );
  INV_X1 U9103 ( .A(n7156), .ZN(n7155) );
  NAND2_X1 U9104 ( .A1(n7157), .A2(n14263), .ZN(n7156) );
  AND2_X1 U9105 ( .A1(n13653), .A2(n13652), .ZN(n13534) );
  INV_X1 U9106 ( .A(n13534), .ZN(n6952) );
  OR2_X1 U9107 ( .A1(n12238), .A2(n12237), .ZN(n6542) );
  INV_X1 U9108 ( .A(n6452), .ZN(n7611) );
  INV_X1 U9109 ( .A(n7499), .ZN(n7498) );
  NAND2_X1 U9110 ( .A1(n11791), .A2(n7636), .ZN(n7499) );
  NAND2_X1 U9111 ( .A1(n11597), .A2(n12809), .ZN(n12813) );
  AND3_X1 U9112 ( .A1(n8702), .A2(n7546), .A3(n8576), .ZN(n6543) );
  OR2_X1 U9113 ( .A1(n7437), .A2(n9536), .ZN(n6544) );
  AND2_X1 U9114 ( .A1(n9667), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6545) );
  OR2_X1 U9115 ( .A1(n14281), .A2(n13778), .ZN(n6546) );
  INV_X1 U9116 ( .A(n6828), .ZN(n6827) );
  NAND2_X1 U9117 ( .A1(n6831), .A2(n12090), .ZN(n6828) );
  AND2_X1 U9118 ( .A1(n7027), .A2(n13126), .ZN(n6547) );
  AND2_X1 U9119 ( .A1(n11008), .A2(n10973), .ZN(n6548) );
  INV_X1 U9120 ( .A(n7199), .ZN(n7198) );
  OAI21_X1 U9121 ( .B1(n7202), .B2(n7204), .A(n6546), .ZN(n7199) );
  AND2_X1 U9122 ( .A1(n8022), .A2(n8021), .ZN(n6549) );
  NAND2_X1 U9123 ( .A1(n10236), .A2(n12913), .ZN(n6550) );
  INV_X1 U9124 ( .A(n7758), .ZN(n7279) );
  NAND2_X1 U9125 ( .A1(n11635), .A2(n11634), .ZN(n6551) );
  INV_X1 U9126 ( .A(n7468), .ZN(n7467) );
  NAND2_X1 U9127 ( .A1(n10296), .A2(n10297), .ZN(n7468) );
  OR2_X1 U9128 ( .A1(n6499), .A2(n6830), .ZN(n6552) );
  OR2_X1 U9129 ( .A1(n11676), .A2(n7312), .ZN(n6553) );
  INV_X1 U9130 ( .A(n13591), .ZN(n7371) );
  AND2_X1 U9131 ( .A1(n7624), .A2(n8086), .ZN(n6554) );
  OR2_X1 U9132 ( .A1(n9687), .A2(n12924), .ZN(n6555) );
  AND2_X1 U9133 ( .A1(n9537), .A2(n9534), .ZN(n6556) );
  OR2_X1 U9134 ( .A1(n14369), .A2(n14865), .ZN(n6557) );
  AND2_X1 U9135 ( .A1(n12384), .A2(n12383), .ZN(n6558) );
  OR2_X1 U9136 ( .A1(n11575), .A2(n11574), .ZN(n6559) );
  AND3_X1 U9137 ( .A1(n7502), .A2(n7501), .A3(n9522), .ZN(n6560) );
  OR2_X1 U9138 ( .A1(n8246), .A2(n6505), .ZN(n6561) );
  AND2_X1 U9139 ( .A1(n6466), .A2(n12802), .ZN(n6562) );
  INV_X1 U9140 ( .A(n7211), .ZN(n15139) );
  AND2_X1 U9141 ( .A1(n11678), .A2(n11358), .ZN(n6563) );
  AND2_X1 U9142 ( .A1(n7126), .A2(n8027), .ZN(n6564) );
  NOR2_X1 U9143 ( .A1(P3_IR_REG_27__SCAN_IN), .A2(P3_IR_REG_28__SCAN_IN), .ZN(
        n6565) );
  INV_X1 U9144 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7276) );
  AND2_X1 U9145 ( .A1(n7485), .A2(n7483), .ZN(n6566) );
  NOR2_X1 U9146 ( .A1(n9049), .A2(n7563), .ZN(n7562) );
  AND2_X1 U9147 ( .A1(n6952), .A2(n9542), .ZN(n6567) );
  OR2_X1 U9148 ( .A1(n8369), .A2(n8370), .ZN(n6568) );
  OR2_X1 U9149 ( .A1(n13606), .A2(n13604), .ZN(n6569) );
  OR2_X1 U9150 ( .A1(n7374), .A2(n13616), .ZN(n6570) );
  NAND2_X1 U9151 ( .A1(n13376), .A2(n13485), .ZN(n6571) );
  OR2_X1 U9152 ( .A1(n7922), .A2(n6502), .ZN(n6572) );
  AND2_X1 U9153 ( .A1(n7379), .A2(n7378), .ZN(n6573) );
  OR2_X1 U9154 ( .A1(n13702), .A2(n13704), .ZN(n6574) );
  AND2_X1 U9155 ( .A1(n6811), .A2(n7684), .ZN(n6575) );
  OR2_X1 U9156 ( .A1(n7525), .A2(n6467), .ZN(n6576) );
  AND2_X1 U9157 ( .A1(n7231), .A2(n7237), .ZN(n6577) );
  AND2_X1 U9158 ( .A1(n6478), .A2(n7049), .ZN(n6578) );
  INV_X1 U9159 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7381) );
  INV_X1 U9160 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7378) );
  INV_X1 U9161 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8513) );
  NAND2_X1 U9162 ( .A1(n13628), .A2(n7364), .ZN(n6579) );
  AND2_X1 U9163 ( .A1(n9141), .A2(n7454), .ZN(n6580) );
  INV_X1 U9165 ( .A(n13255), .ZN(n6945) );
  AND2_X1 U9166 ( .A1(n8621), .A2(n8620), .ZN(n12483) );
  INV_X1 U9167 ( .A(n12483), .ZN(n7249) );
  XNOR2_X1 U9168 ( .A(n8642), .B(P3_IR_REG_1__SCAN_IN), .ZN(n10414) );
  AND2_X1 U9169 ( .A1(n7547), .A2(n6469), .ZN(n8788) );
  INV_X1 U9170 ( .A(n13013), .ZN(n7351) );
  OR2_X1 U9171 ( .A1(n8136), .A2(SI_18_), .ZN(n6581) );
  XNOR2_X1 U9172 ( .A(n14285), .B(n13779), .ZN(n14078) );
  INV_X1 U9173 ( .A(n14078), .ZN(n7443) );
  NAND2_X1 U9174 ( .A1(n8897), .A2(n6519), .ZN(n9100) );
  AND2_X1 U9175 ( .A1(n9930), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n6582) );
  INV_X1 U9176 ( .A(n13275), .ZN(n7173) );
  INV_X1 U9177 ( .A(n12201), .ZN(n7001) );
  AND4_X1 U9178 ( .A1(n8878), .A2(n8877), .A3(n8876), .A4(n8875), .ZN(n12066)
         );
  OR2_X1 U9179 ( .A1(n9134), .A2(n9133), .ZN(n6583) );
  AND2_X1 U9180 ( .A1(n10167), .A2(n8459), .ZN(n10158) );
  INV_X1 U9181 ( .A(n10158), .ZN(n6927) );
  INV_X1 U9182 ( .A(n7447), .ZN(n7445) );
  NOR2_X1 U9183 ( .A1(n14098), .A2(n7448), .ZN(n7447) );
  NAND2_X1 U9184 ( .A1(n8212), .A2(n8211), .ZN(n13280) );
  INV_X1 U9185 ( .A(n13280), .ZN(n7175) );
  AND2_X1 U9186 ( .A1(n11792), .A2(n11793), .ZN(n6584) );
  INV_X1 U9187 ( .A(n12543), .ZN(n11928) );
  NAND2_X1 U9188 ( .A1(n8938), .A2(n8937), .ZN(n12543) );
  AND2_X1 U9189 ( .A1(n9046), .A2(n12169), .ZN(n6585) );
  INV_X1 U9190 ( .A(n7555), .ZN(n7554) );
  NOR2_X1 U9191 ( .A1(n12552), .A2(n7556), .ZN(n7555) );
  INV_X1 U9192 ( .A(n7588), .ZN(n7587) );
  NAND2_X1 U9193 ( .A1(n7648), .A2(n6581), .ZN(n7588) );
  INV_X1 U9194 ( .A(n6706), .ZN(n11243) );
  NAND2_X1 U9195 ( .A1(n7386), .A2(n7383), .ZN(n6706) );
  AND2_X1 U9196 ( .A1(n12067), .A2(n12610), .ZN(n6586) );
  INV_X1 U9197 ( .A(n7176), .ZN(n13108) );
  AND2_X1 U9198 ( .A1(n11731), .A2(n6947), .ZN(n7176) );
  AND2_X1 U9199 ( .A1(n7356), .A2(n7355), .ZN(n6587) );
  NOR2_X1 U9200 ( .A1(n12756), .A2(n12584), .ZN(n6588) );
  INV_X1 U9201 ( .A(n7239), .ZN(n7236) );
  NAND2_X1 U9202 ( .A1(n12223), .A2(n12568), .ZN(n7239) );
  NOR2_X1 U9203 ( .A1(n14407), .A2(n14408), .ZN(n14601) );
  INV_X1 U9204 ( .A(n14601), .ZN(n6783) );
  AND2_X1 U9205 ( .A1(n10756), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n6589) );
  AND2_X1 U9206 ( .A1(n12279), .A2(n11436), .ZN(n6590) );
  INV_X1 U9207 ( .A(n6974), .ZN(n7487) );
  NAND2_X1 U9208 ( .A1(n6733), .A2(n6508), .ZN(n6974) );
  NOR2_X1 U9209 ( .A1(n12333), .A2(n12334), .ZN(n6591) );
  AND2_X1 U9210 ( .A1(n8180), .A2(n7518), .ZN(n6592) );
  NOR2_X1 U9211 ( .A1(n11680), .A2(n11580), .ZN(n6593) );
  NOR2_X1 U9212 ( .A1(n12329), .A2(n12330), .ZN(n6594) );
  AND2_X1 U9213 ( .A1(n7060), .A2(n7061), .ZN(n6595) );
  AND2_X1 U9214 ( .A1(n11781), .A2(n11776), .ZN(n6596) );
  AND2_X1 U9215 ( .A1(n12577), .A2(n8909), .ZN(n6597) );
  INV_X1 U9216 ( .A(n6832), .ZN(n6830) );
  NAND2_X1 U9217 ( .A1(n12680), .A2(n12508), .ZN(n6832) );
  INV_X1 U9218 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9645) );
  NAND2_X1 U9219 ( .A1(n7734), .A2(n7736), .ZN(n11372) );
  INV_X1 U9220 ( .A(n11372), .ZN(n6795) );
  INV_X1 U9221 ( .A(n12722), .ZN(n6842) );
  INV_X1 U9222 ( .A(n10558), .ZN(n6742) );
  NAND2_X1 U9223 ( .A1(n7706), .A2(n7705), .ZN(n8484) );
  AND3_X1 U9224 ( .A1(n7148), .A2(n7147), .A3(n14575), .ZN(n6598) );
  NAND2_X1 U9225 ( .A1(n7258), .A2(n9908), .ZN(n10195) );
  INV_X1 U9226 ( .A(n11423), .ZN(n7166) );
  INV_X1 U9227 ( .A(n11376), .ZN(n7169) );
  INV_X1 U9228 ( .A(n13194), .ZN(n11580) );
  NOR2_X1 U9229 ( .A1(n8925), .A2(n7117), .ZN(n7116) );
  NOR2_X1 U9230 ( .A1(n15064), .A2(n15063), .ZN(n6599) );
  NOR2_X1 U9231 ( .A1(n15070), .A2(n15069), .ZN(n6600) );
  AND2_X1 U9232 ( .A1(n14909), .A2(n11285), .ZN(n6601) );
  OR2_X1 U9233 ( .A1(n8346), .A2(SI_27_), .ZN(n6602) );
  NAND2_X1 U9234 ( .A1(n6706), .A2(n6507), .ZN(n6705) );
  NAND2_X1 U9235 ( .A1(n6598), .A2(n7146), .ZN(n14458) );
  INV_X1 U9236 ( .A(n14458), .ZN(n6617) );
  AND2_X1 U9237 ( .A1(n8378), .A2(SI_30_), .ZN(n6603) );
  NAND2_X1 U9238 ( .A1(n10847), .A2(n7496), .ZN(n7495) );
  INV_X1 U9239 ( .A(n7147), .ZN(n14687) );
  NOR2_X2 U9240 ( .A1(n14686), .A2(n14693), .ZN(n7147) );
  AND2_X1 U9241 ( .A1(n10221), .A2(n9530), .ZN(n6604) );
  AND2_X1 U9242 ( .A1(n7458), .A2(n7457), .ZN(n6605) );
  NOR2_X1 U9243 ( .A1(n8420), .A2(n7604), .ZN(n7603) );
  INV_X1 U9244 ( .A(n6453), .ZN(n7227) );
  OR2_X1 U9245 ( .A1(n7109), .A2(n7108), .ZN(n6606) );
  INV_X1 U9246 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6713) );
  INV_X2 U9247 ( .A(n15205), .ZN(n15206) );
  NAND2_X1 U9248 ( .A1(n9743), .A2(n9733), .ZN(n12902) );
  AND2_X1 U9249 ( .A1(n10407), .A2(n10398), .ZN(n15089) );
  AND2_X1 U9250 ( .A1(n12337), .A2(n12336), .ZN(n6607) );
  OR2_X1 U9251 ( .A1(n15205), .A2(n15138), .ZN(n12776) );
  INV_X1 U9252 ( .A(n14730), .ZN(n14704) );
  AND2_X1 U9253 ( .A1(n15084), .A2(n12442), .ZN(n6608) );
  INV_X1 U9254 ( .A(n12370), .ZN(n14484) );
  INV_X1 U9255 ( .A(n10166), .ZN(n6936) );
  AND2_X1 U9256 ( .A1(n12383), .A2(n12417), .ZN(n6609) );
  OR3_X1 U9257 ( .A1(n9989), .A2(n13766), .A3(n9988), .ZN(n15379) );
  INV_X1 U9258 ( .A(n13757), .ZN(n7592) );
  INV_X1 U9259 ( .A(SI_26_), .ZN(n15289) );
  INV_X1 U9260 ( .A(n8389), .ZN(n7608) );
  INV_X1 U9261 ( .A(n11300), .ZN(n6714) );
  INV_X1 U9262 ( .A(n12428), .ZN(n12442) );
  INV_X1 U9263 ( .A(n15140), .ZN(n6677) );
  XOR2_X1 U9264 ( .A(n8650), .B(n8641), .Z(n6610) );
  INV_X1 U9265 ( .A(SI_1_), .ZN(n7077) );
  INV_X1 U9266 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n6774) );
  INV_X1 U9267 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n7218) );
  INV_X1 U9268 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n6789) );
  INV_X1 U9269 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6918) );
  NOR2_X1 U9270 ( .A1(n7171), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11855) );
  NAND2_X1 U9271 ( .A1(n10628), .A2(n10627), .ZN(n10653) );
  NOR2_X1 U9272 ( .A1(n7099), .A2(n10627), .ZN(n7098) );
  NAND2_X1 U9273 ( .A1(n7097), .A2(n10627), .ZN(n10659) );
  XNOR2_X1 U9274 ( .A(n12328), .B(n12336), .ZN(n12322) );
  XNOR2_X1 U9275 ( .A(n12332), .B(n12336), .ZN(n12304) );
  AND2_X2 U9276 ( .A1(n6612), .A2(n6611), .ZN(n7428) );
  NOR2_X2 U9277 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n6611) );
  NOR2_X2 U9278 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n6612) );
  XNOR2_X1 U9279 ( .A(n6613), .B(n9141), .ZN(n9567) );
  NOR2_X2 U9280 ( .A1(n10580), .A2(n13394), .ZN(n10488) );
  AND3_X2 U9281 ( .A1(n6614), .A2(n9193), .A3(n9192), .ZN(n13578) );
  INV_X1 U9282 ( .A(n14726), .ZN(n6615) );
  AND3_X2 U9283 ( .A1(n9163), .A2(n9164), .A3(n9162), .ZN(n14751) );
  NOR2_X2 U9284 ( .A1(n14459), .A2(n11506), .ZN(n11517) );
  NAND2_X1 U9285 ( .A1(n10273), .A2(n10274), .ZN(n10325) );
  NAND3_X1 U9286 ( .A1(n10200), .A2(n7075), .A3(n15147), .ZN(n10272) );
  NAND2_X1 U9287 ( .A1(n7074), .A2(n10196), .ZN(n10200) );
  NAND2_X2 U9288 ( .A1(n6620), .A2(n6500), .ZN(n11999) );
  OR2_X2 U9289 ( .A1(n11139), .A2(n11959), .ZN(n6620) );
  NAND3_X1 U9290 ( .A1(n6623), .A2(n6486), .A3(n15124), .ZN(n12118) );
  NAND2_X2 U9291 ( .A1(n12122), .A2(n12118), .ZN(n15148) );
  NAND2_X1 U9292 ( .A1(n11943), .A2(n11944), .ZN(n7271) );
  NAND3_X1 U9293 ( .A1(n8897), .A2(n7572), .A3(n6628), .ZN(n8585) );
  AND2_X2 U9294 ( .A1(n6630), .A2(n6484), .ZN(n11934) );
  INV_X1 U9295 ( .A(n12383), .ZN(n6637) );
  NOR2_X1 U9296 ( .A1(n12402), .A2(n12403), .ZN(n12405) );
  INV_X1 U9297 ( .A(n10629), .ZN(n6639) );
  INV_X1 U9298 ( .A(n10627), .ZN(n6641) );
  INV_X1 U9299 ( .A(n10628), .ZN(n6642) );
  INV_X1 U9300 ( .A(n7162), .ZN(n12356) );
  NOR2_X1 U9301 ( .A1(n14486), .A2(n14487), .ZN(n14485) );
  NOR2_X1 U9302 ( .A1(n12322), .A2(n12305), .ZN(n12329) );
  OAI211_X1 U9303 ( .C1(n12330), .C2(n6644), .A(n6643), .B(n7160), .ZN(n12350)
         );
  OR2_X1 U9304 ( .A1(n12330), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n6643) );
  INV_X1 U9305 ( .A(n6646), .ZN(n10448) );
  NAND2_X1 U9306 ( .A1(n10445), .A2(n10477), .ZN(n6646) );
  NAND2_X1 U9307 ( .A1(n10676), .A2(n6646), .ZN(n10446) );
  NAND2_X1 U9308 ( .A1(n6651), .A2(n10662), .ZN(n10663) );
  NAND3_X1 U9309 ( .A1(n6658), .A2(n6661), .A3(n6656), .ZN(n12388) );
  NAND3_X1 U9310 ( .A1(n6658), .A2(n6657), .A3(n6656), .ZN(n6662) );
  OAI21_X1 U9311 ( .B1(n12333), .B2(n6663), .A(n6606), .ZN(n12371) );
  NAND2_X1 U9312 ( .A1(n8557), .A2(n6669), .ZN(n6666) );
  NAND2_X1 U9313 ( .A1(n6671), .A2(n12272), .ZN(P3_U3296) );
  NAND2_X1 U9314 ( .A1(n6673), .A2(n6672), .ZN(n6671) );
  INV_X1 U9315 ( .A(n6675), .ZN(n6674) );
  OAI21_X1 U9316 ( .B1(n12266), .B2(n6677), .A(n6676), .ZN(n6675) );
  NAND2_X1 U9317 ( .A1(n12266), .A2(n12267), .ZN(n6676) );
  NAND2_X1 U9318 ( .A1(n12248), .A2(n6699), .ZN(n12250) );
  NAND3_X1 U9319 ( .A1(n12243), .A2(n12242), .A3(n6701), .ZN(n6700) );
  NAND2_X1 U9320 ( .A1(n6542), .A2(n6702), .ZN(n6701) );
  AND2_X2 U9321 ( .A1(n6705), .A2(n6704), .ZN(n11558) );
  NAND2_X1 U9322 ( .A1(n10026), .A2(n10027), .ZN(n10062) );
  NAND2_X1 U9323 ( .A1(n10025), .A2(n10024), .ZN(n10026) );
  NAND3_X1 U9324 ( .A1(n6708), .A2(n7788), .A3(n7842), .ZN(n7859) );
  OR2_X1 U9325 ( .A1(n9757), .A2(n9756), .ZN(n9758) );
  NAND3_X1 U9326 ( .A1(n10780), .A2(n10781), .A3(n10778), .ZN(n10827) );
  INV_X1 U9327 ( .A(n6720), .ZN(n14951) );
  NOR2_X1 U9328 ( .A1(n14962), .A2(n14961), .ZN(n14959) );
  XNOR2_X1 U9329 ( .A(n11287), .B(n11306), .ZN(n14953) );
  NAND2_X1 U9330 ( .A1(n6460), .A2(n10746), .ZN(n6973) );
  NAND3_X1 U9331 ( .A1(n11755), .A2(n11754), .A3(n6736), .ZN(n13492) );
  AND2_X2 U9332 ( .A1(n9149), .A2(n9148), .ZN(n13503) );
  INV_X2 U9333 ( .A(n8162), .ZN(n8146) );
  NAND2_X2 U9334 ( .A1(n6741), .A2(n6739), .ZN(n10128) );
  AOI21_X1 U9335 ( .B1(n8145), .B2(n14845), .A(n6740), .ZN(n6739) );
  NOR2_X1 U9336 ( .A1(n8162), .A2(n9645), .ZN(n6740) );
  NAND2_X2 U9337 ( .A1(n9687), .A2(n9155), .ZN(n8162) );
  NAND3_X1 U9338 ( .A1(n6743), .A2(n6744), .A3(n6742), .ZN(n6747) );
  OR2_X1 U9339 ( .A1(n10237), .A2(n6746), .ZN(n6743) );
  NAND2_X1 U9340 ( .A1(n10237), .A2(n10236), .ZN(n10334) );
  NOR2_X1 U9341 ( .A1(n6939), .A2(n10244), .ZN(n6746) );
  NAND2_X1 U9342 ( .A1(n6747), .A2(n10554), .ZN(n10555) );
  NAND2_X1 U9343 ( .A1(n13133), .A2(n11714), .ZN(n11716) );
  OAI21_X1 U9344 ( .B1(n10868), .B2(n10869), .A(n6753), .ZN(n10870) );
  NAND2_X1 U9345 ( .A1(n12996), .A2(n11724), .ZN(n11726) );
  NAND2_X1 U9346 ( .A1(n14373), .A2(n14374), .ZN(n6889) );
  INV_X1 U9347 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6760) );
  XNOR2_X2 U9348 ( .A(n6761), .B(n7739), .ZN(n7762) );
  NAND2_X1 U9349 ( .A1(n7514), .A2(n7834), .ZN(n7052) );
  NAND2_X1 U9350 ( .A1(n6764), .A2(n6763), .ZN(n6762) );
  INV_X1 U9351 ( .A(n7811), .ZN(n6763) );
  INV_X1 U9352 ( .A(n7812), .ZN(n6764) );
  NAND2_X1 U9353 ( .A1(n6767), .A2(n6766), .ZN(n6765) );
  NAND2_X1 U9354 ( .A1(n7812), .A2(n7811), .ZN(n6766) );
  NAND2_X1 U9355 ( .A1(n14607), .A2(n6772), .ZN(n14613) );
  NAND3_X1 U9356 ( .A1(n14603), .A2(n6773), .A3(n14605), .ZN(n6768) );
  NAND2_X1 U9357 ( .A1(n14603), .A2(n14605), .ZN(n14609) );
  NAND3_X1 U9358 ( .A1(n6776), .A2(n7524), .A3(n6572), .ZN(n6775) );
  NAND3_X1 U9359 ( .A1(n7882), .A2(n6576), .A3(n7881), .ZN(n6776) );
  NAND3_X1 U9360 ( .A1(n6779), .A2(n6561), .A3(n6778), .ZN(n6777) );
  OR2_X1 U9361 ( .A1(n8226), .A2(n8225), .ZN(n6778) );
  NAND2_X1 U9362 ( .A1(n6780), .A2(n7054), .ZN(n6779) );
  NAND2_X1 U9363 ( .A1(n8226), .A2(n8225), .ZN(n6780) );
  OAI22_X1 U9364 ( .A1(n7051), .A2(n6781), .B1(n7854), .B2(n7853), .ZN(n7877)
         );
  OAI22_X1 U9365 ( .A1(n6784), .A2(n6522), .B1(n8132), .B2(n8131), .ZN(n8158)
         );
  OAI21_X2 U9366 ( .B1(n6786), .B2(n7039), .A(n7038), .ZN(n8509) );
  OAI21_X2 U9367 ( .B1(n14439), .B2(n6788), .A(n6787), .ZN(n7330) );
  NAND2_X1 U9368 ( .A1(n7330), .A2(n7329), .ZN(n7327) );
  NAND2_X1 U9369 ( .A1(n6790), .A2(n7537), .ZN(n8043) );
  NAND3_X1 U9370 ( .A1(n6792), .A2(n6791), .A3(n7535), .ZN(n6790) );
  OAI21_X1 U9371 ( .B1(n6793), .B2(n7529), .A(n7526), .ZN(n6791) );
  OAI21_X1 U9372 ( .B1(n6793), .B2(n7532), .A(n7041), .ZN(n6792) );
  OR2_X1 U9373 ( .A1(n7966), .A2(n7965), .ZN(n6793) );
  NAND3_X1 U9374 ( .A1(n7580), .A2(n7583), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n7579) );
  OAI21_X1 U9375 ( .B1(SI_1_), .B2(n6796), .A(n7657), .ZN(n7784) );
  NOR2_X1 U9376 ( .A1(n7360), .A2(n13701), .ZN(n6797) );
  NAND3_X1 U9377 ( .A1(n6797), .A2(n13694), .A3(n13695), .ZN(n6801) );
  NAND3_X1 U9378 ( .A1(n6800), .A2(n6574), .A3(n6798), .ZN(n7361) );
  NAND2_X1 U9379 ( .A1(n13695), .A2(n13694), .ZN(n6799) );
  NAND3_X1 U9380 ( .A1(n6801), .A2(n7357), .A3(n13699), .ZN(n6800) );
  NAND2_X1 U9381 ( .A1(n7824), .A2(n7660), .ZN(n6804) );
  NAND2_X1 U9382 ( .A1(n7825), .A2(n7660), .ZN(n6805) );
  INV_X1 U9383 ( .A(n7824), .ZN(n6806) );
  INV_X1 U9384 ( .A(n7825), .ZN(n6807) );
  NAND2_X1 U9385 ( .A1(n6808), .A2(n6575), .ZN(n7685) );
  NAND3_X1 U9386 ( .A1(n6813), .A2(n6564), .A3(n7123), .ZN(n6808) );
  NAND3_X1 U9387 ( .A1(n6813), .A2(n7123), .A3(n7126), .ZN(n6810) );
  INV_X1 U9388 ( .A(n13718), .ZN(n13721) );
  OAI22_X2 U9389 ( .A1(n13715), .A2(n6817), .B1(n6818), .B2(n13714), .ZN(
        n13718) );
  NAND2_X1 U9390 ( .A1(n12519), .A2(n6824), .ZN(n6821) );
  AND2_X4 U9391 ( .A1(n10395), .A2(n7171), .ZN(n8664) );
  NAND3_X1 U9392 ( .A1(n6837), .A2(n6838), .A3(n8580), .ZN(n8895) );
  NOR2_X1 U9393 ( .A1(n7545), .A2(n8687), .ZN(n8807) );
  NAND2_X1 U9394 ( .A1(n12671), .A2(n6841), .ZN(P3_U3485) );
  NAND2_X1 U9395 ( .A1(n12734), .A2(n6843), .ZN(P3_U3453) );
  NAND2_X1 U9396 ( .A1(n7209), .A2(n7208), .ZN(n15111) );
  NAND2_X1 U9397 ( .A1(n7232), .A2(n6577), .ZN(n12519) );
  XNOR2_X1 U9398 ( .A(n12482), .B(n12486), .ZN(n6849) );
  NAND2_X1 U9399 ( .A1(n10810), .A2(n12146), .ZN(n10809) );
  NAND4_X1 U9400 ( .A1(n6543), .A2(n8574), .A3(n8575), .A4(n8573), .ZN(n7545)
         );
  NAND3_X1 U9401 ( .A1(n9042), .A2(n12118), .A3(n10268), .ZN(n10198) );
  INV_X1 U9402 ( .A(n10989), .ZN(n6851) );
  XNOR2_X1 U9403 ( .A(n12441), .B(n6859), .ZN(n6858) );
  NAND2_X1 U9404 ( .A1(n6857), .A2(n6855), .ZN(n12445) );
  NOR2_X1 U9405 ( .A1(n12313), .A2(n12312), .ZN(n12340) );
  NOR2_X1 U9406 ( .A1(n12359), .A2(n14484), .ZN(n12361) );
  NOR2_X1 U9407 ( .A1(n15072), .A2(n15073), .ZN(n15071) );
  NOR2_X1 U9408 ( .A1(n10483), .A2(n10482), .ZN(n10610) );
  XNOR2_X1 U9409 ( .A(n12431), .B(n12432), .ZN(n12413) );
  AOI21_X1 U9410 ( .B1(n10777), .B2(n10775), .A(n10774), .ZN(n10780) );
  INV_X4 U9411 ( .A(n11584), .ZN(n11592) );
  OAI21_X2 U9412 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(n14415), .A(n14466), .ZN(
        n14473) );
  NOR2_X1 U9413 ( .A1(n14468), .A2(n14467), .ZN(n14415) );
  NAND2_X1 U9414 ( .A1(n7318), .A2(n14611), .ZN(n14468) );
  NAND2_X1 U9415 ( .A1(n6861), .A2(n6860), .ZN(n14163) );
  OR2_X1 U9416 ( .A1(n14261), .A2(n9605), .ZN(n6861) );
  NAND2_X1 U9417 ( .A1(n6863), .A2(n6862), .ZN(n14262) );
  OR2_X1 U9418 ( .A1(n14261), .A2(n14808), .ZN(n6863) );
  NOR2_X1 U9419 ( .A1(n15057), .A2(n8727), .ZN(n15056) );
  NAND2_X1 U9420 ( .A1(n7162), .A2(n7161), .ZN(n12384) );
  OAI21_X1 U9421 ( .B1(n10722), .B2(n10468), .A(n7163), .ZN(n10707) );
  INV_X1 U9422 ( .A(n7285), .ZN(n7284) );
  OAI21_X1 U9423 ( .B1(n11912), .B2(n11134), .A(n11876), .ZN(n11137) );
  NAND2_X1 U9424 ( .A1(n14473), .A2(n14474), .ZN(n14475) );
  NAND2_X1 U9425 ( .A1(n7271), .A2(n11655), .ZN(n6933) );
  INV_X1 U9426 ( .A(n10126), .ZN(n10003) );
  XNOR2_X1 U9427 ( .A(n11726), .B(n11725), .ZN(n13248) );
  INV_X1 U9428 ( .A(n7706), .ZN(n8488) );
  AND2_X4 U9429 ( .A1(n7704), .A2(n8007), .ZN(n7706) );
  OAI21_X1 U9430 ( .B1(n13200), .B2(n13202), .A(n11708), .ZN(n13182) );
  NAND2_X1 U9431 ( .A1(n13707), .A2(n13708), .ZN(n13706) );
  NAND2_X1 U9432 ( .A1(n6866), .A2(n6865), .ZN(n13621) );
  NAND3_X1 U9433 ( .A1(n13615), .A2(n13614), .A3(n6570), .ZN(n6866) );
  NAND2_X1 U9434 ( .A1(n13687), .A2(n13688), .ZN(n13689) );
  NAND2_X1 U9435 ( .A1(n13683), .A2(n13682), .ZN(n13687) );
  MUX2_X1 U9436 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14322), .S(n9429), .Z(n13560)
         );
  NAND2_X1 U9437 ( .A1(n6895), .A2(n6894), .ZN(n13610) );
  NAND2_X2 U9438 ( .A1(n13356), .A2(n8497), .ZN(n9687) );
  OR2_X1 U9439 ( .A1(n7884), .A2(n7883), .ZN(n7885) );
  NAND2_X1 U9440 ( .A1(n12801), .A2(n11579), .ZN(n11582) );
  NAND2_X1 U9441 ( .A1(n6873), .A2(n6871), .ZN(P2_U3186) );
  AND2_X1 U9442 ( .A1(n10310), .A2(n10061), .ZN(n6874) );
  NAND3_X1 U9443 ( .A1(n6880), .A2(n12871), .A3(n12779), .ZN(n6873) );
  NAND2_X1 U9444 ( .A1(n11587), .A2(n11586), .ZN(n11588) );
  NAND2_X1 U9445 ( .A1(n11999), .A2(n7256), .ZN(n11430) );
  NAND2_X1 U9446 ( .A1(n6875), .A2(n7134), .ZN(n8113) );
  NAND3_X1 U9447 ( .A1(n7687), .A2(n7626), .A3(n6554), .ZN(n6875) );
  NAND2_X1 U9448 ( .A1(n8541), .A2(n8540), .ZN(n8543) );
  INV_X1 U9449 ( .A(n7552), .ZN(n7551) );
  NAND2_X1 U9450 ( .A1(n8567), .A2(n8566), .ZN(n8965) );
  INV_X1 U9451 ( .A(n7010), .ZN(n7009) );
  INV_X1 U9452 ( .A(n7507), .ZN(n7505) );
  NAND2_X2 U9453 ( .A1(n13093), .A2(n11719), .ZN(n13080) );
  NAND2_X1 U9454 ( .A1(n7113), .A2(n8551), .ZN(n8894) );
  NAND2_X1 U9455 ( .A1(n6926), .A2(n6927), .ZN(n10156) );
  NAND2_X1 U9456 ( .A1(n8524), .A2(n8523), .ZN(n8698) );
  NAND2_X1 U9457 ( .A1(n8783), .A2(n8782), .ZN(n8785) );
  NAND2_X1 U9458 ( .A1(n12778), .A2(n12777), .ZN(n6880) );
  NAND2_X1 U9459 ( .A1(n7065), .A2(n7067), .ZN(n12801) );
  XNOR2_X1 U9460 ( .A(n14373), .B(n6881), .ZN(n14377) );
  INV_X1 U9461 ( .A(n14374), .ZN(n6881) );
  NAND2_X1 U9462 ( .A1(n15406), .A2(n15405), .ZN(n15404) );
  OAI21_X1 U9463 ( .B1(n14380), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n14422), .ZN(
        n15406) );
  NAND2_X1 U9464 ( .A1(n15222), .A2(n15173), .ZN(n12722) );
  INV_X1 U9465 ( .A(n14383), .ZN(n7319) );
  NAND2_X1 U9466 ( .A1(n14370), .A2(n14327), .ZN(n7332) );
  NAND2_X1 U9467 ( .A1(n7082), .A2(n10325), .ZN(n10985) );
  NAND2_X1 U9468 ( .A1(n10198), .A2(n11622), .ZN(n7075) );
  NAND2_X1 U9469 ( .A1(n12998), .A2(n7288), .ZN(n11696) );
  NAND2_X1 U9470 ( .A1(n6884), .A2(n7365), .ZN(n13749) );
  NAND3_X1 U9471 ( .A1(n6893), .A2(n7367), .A3(n6892), .ZN(n6884) );
  NOR2_X1 U9472 ( .A1(n13697), .A2(n13698), .ZN(n7360) );
  NAND2_X1 U9473 ( .A1(n13712), .A2(n13711), .ZN(n13715) );
  NAND2_X1 U9474 ( .A1(n7490), .A2(n6973), .ZN(n11463) );
  NAND2_X1 U9475 ( .A1(n7886), .A2(n7667), .ZN(n7901) );
  NAND2_X1 U9476 ( .A1(n7496), .A2(n7492), .ZN(n7491) );
  NOR2_X1 U9477 ( .A1(n12304), .A2(n12306), .ZN(n12333) );
  NAND2_X1 U9478 ( .A1(n11049), .A2(n11047), .ZN(n7386) );
  NAND2_X2 U9479 ( .A1(n7889), .A2(n7888), .ZN(n15001) );
  NAND2_X1 U9480 ( .A1(n7045), .A2(n7044), .ZN(n8104) );
  OAI211_X1 U9481 ( .C1(n7836), .C2(n7837), .A(n7053), .B(n7052), .ZN(n7051)
         );
  NAND2_X1 U9482 ( .A1(n8044), .A2(n6516), .ZN(n8066) );
  OAI22_X1 U9483 ( .A1(n8203), .A2(n7512), .B1(n7511), .B2(n8204), .ZN(n8226)
         );
  NAND2_X1 U9484 ( .A1(n14430), .A2(n14878), .ZN(n14429) );
  NOR2_X2 U9485 ( .A1(n14431), .A2(n14401), .ZN(n14439) );
  NAND2_X1 U9486 ( .A1(n10706), .A2(n10707), .ZN(n10705) );
  XNOR2_X1 U9487 ( .A(n11400), .B(n11419), .ZN(n11068) );
  XNOR2_X1 U9488 ( .A(n14396), .B(n7325), .ZN(n14430) );
  NAND2_X1 U9489 ( .A1(n6496), .A2(n14475), .ZN(n6890) );
  NAND2_X1 U9490 ( .A1(n7324), .A2(n14475), .ZN(n7323) );
  NOR2_X1 U9491 ( .A1(n14423), .A2(n14424), .ZN(n14380) );
  XNOR2_X1 U9492 ( .A(n6890), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  NAND2_X1 U9493 ( .A1(n14372), .A2(n14371), .ZN(n14325) );
  NAND2_X1 U9494 ( .A1(n12261), .A2(n12257), .ZN(n12259) );
  NAND2_X1 U9495 ( .A1(n12251), .A2(n12461), .ZN(n12261) );
  NAND2_X1 U9496 ( .A1(n6891), .A2(n7363), .ZN(n13633) );
  NAND3_X1 U9497 ( .A1(n13626), .A2(n6579), .A3(n13625), .ZN(n6891) );
  NAND2_X1 U9498 ( .A1(n13721), .A2(n13720), .ZN(n6892) );
  NAND2_X1 U9499 ( .A1(n13717), .A2(n13716), .ZN(n6893) );
  NAND3_X1 U9500 ( .A1(n13602), .A2(n13601), .A3(n6569), .ZN(n6895) );
  INV_X1 U9501 ( .A(n7377), .ZN(n9397) );
  INV_X4 U9502 ( .A(n13734), .ZN(n13732) );
  NAND2_X1 U9503 ( .A1(n15381), .A2(n11748), .ZN(n11751) );
  NAND2_X1 U9504 ( .A1(n7609), .A2(n7611), .ZN(n8005) );
  INV_X1 U9505 ( .A(n14550), .ZN(n7489) );
  NAND4_X1 U9506 ( .A1(n7425), .A2(n7429), .A3(n6481), .A4(n9201), .ZN(n9577)
         );
  NAND2_X1 U9507 ( .A1(n9552), .A2(n9551), .ZN(n13979) );
  NAND2_X1 U9508 ( .A1(n14077), .A2(n14281), .ZN(n14066) );
  OR2_X2 U9509 ( .A1(n10590), .A2(n13590), .ZN(n14713) );
  AND2_X2 U9510 ( .A1(n14714), .A2(n10765), .ZN(n10795) );
  INV_X1 U9511 ( .A(n8610), .ZN(n8608) );
  XNOR2_X1 U9512 ( .A(n6933), .B(n6932), .ZN(n12056) );
  OAI21_X1 U9513 ( .B1(n13113), .B2(n13104), .A(n11718), .ZN(n13090) );
  AND2_X1 U9514 ( .A1(n7804), .A2(n6555), .ZN(n6906) );
  NAND2_X1 U9515 ( .A1(n11716), .A2(n11715), .ZN(n13117) );
  NAND3_X1 U9516 ( .A1(n6909), .A2(n13262), .A3(n13261), .ZN(n13333) );
  NAND2_X1 U9517 ( .A1(n7782), .A2(n7656), .ZN(n7786) );
  NOR2_X1 U9518 ( .A1(n7655), .A2(n9640), .ZN(n7782) );
  NAND3_X1 U9519 ( .A1(n6913), .A2(n6912), .A3(n8449), .ZN(n8443) );
  NAND2_X1 U9520 ( .A1(n8008), .A2(n7711), .ZN(n7716) );
  INV_X1 U9521 ( .A(n7716), .ZN(n7717) );
  NAND2_X1 U9522 ( .A1(n15101), .A2(n15102), .ZN(n15099) );
  OAI21_X1 U9523 ( .B1(n10648), .B2(n10647), .A(n10646), .ZN(n10650) );
  XNOR2_X1 U9524 ( .A(n7323), .B(n7322), .ZN(SUB_1596_U4) );
  XNOR2_X1 U9525 ( .A(n14377), .B(n14378), .ZN(n15409) );
  NAND2_X1 U9526 ( .A1(n10894), .A2(n10893), .ZN(n11195) );
  NAND2_X1 U9527 ( .A1(n11707), .A2(n11706), .ZN(n13200) );
  NAND2_X1 U9528 ( .A1(n14606), .A2(n14947), .ZN(n14603) );
  NAND2_X1 U9529 ( .A1(n10555), .A2(n10563), .ZN(n10868) );
  XNOR2_X2 U9530 ( .A(n12915), .B(n10128), .ZN(n10126) );
  NAND2_X1 U9531 ( .A1(n12057), .A2(n11626), .ZN(n11953) );
  INV_X1 U9532 ( .A(n9908), .ZN(n7264) );
  NAND3_X1 U9533 ( .A1(n7266), .A2(n7265), .A3(n7269), .ZN(n12057) );
  INV_X1 U9534 ( .A(n11151), .ZN(n9096) );
  NAND2_X1 U9535 ( .A1(n9080), .A2(n9079), .ZN(n11151) );
  NAND2_X1 U9536 ( .A1(n6962), .A2(n9610), .ZN(P1_U3557) );
  NAND2_X1 U9537 ( .A1(n14034), .A2(n7410), .ZN(n14012) );
  NAND2_X1 U9538 ( .A1(n7415), .A2(n6448), .ZN(n13966) );
  NAND2_X1 U9539 ( .A1(n7903), .A2(n7668), .ZN(n7924) );
  NAND2_X1 U9540 ( .A1(n15050), .A2(n15051), .ZN(n15049) );
  NAND2_X1 U9541 ( .A1(n9008), .A2(n9007), .ZN(n11852) );
  NAND2_X1 U9542 ( .A1(n8953), .A2(n11547), .ZN(n8567) );
  OAI21_X1 U9543 ( .B1(n8736), .B2(n8735), .A(n8530), .ZN(n8749) );
  AOI21_X1 U9544 ( .B1(n11407), .B2(n11406), .A(n11405), .ZN(n15072) );
  AOI21_X1 U9545 ( .B1(n10612), .B2(n10611), .A(n10610), .ZN(n10648) );
  NAND2_X1 U9546 ( .A1(n8749), .A2(n8748), .ZN(n8751) );
  NAND2_X1 U9547 ( .A1(n12885), .A2(n11604), .ZN(n12778) );
  NAND2_X1 U9548 ( .A1(n13692), .A2(n13691), .ZN(n6921) );
  NAND2_X1 U9549 ( .A1(n13651), .A2(n6922), .ZN(n13655) );
  NOR2_X1 U9550 ( .A1(n6492), .A2(n6923), .ZN(n6922) );
  INV_X1 U9551 ( .A(n15383), .ZN(n11506) );
  NAND2_X1 U9552 ( .A1(n9619), .A2(n8513), .ZN(n7654) );
  NAND2_X1 U9553 ( .A1(n7057), .A2(n7055), .ZN(n7903) );
  NAND2_X1 U9554 ( .A1(n7625), .A2(n7687), .ZN(n8048) );
  NAND2_X1 U9555 ( .A1(n7411), .A2(n14024), .ZN(n14034) );
  NAND2_X1 U9556 ( .A1(n7412), .A2(n9554), .ZN(n7415) );
  NAND2_X1 U9557 ( .A1(n7858), .A2(n7121), .ZN(n7057) );
  INV_X1 U9558 ( .A(n13182), .ZN(n11710) );
  XNOR2_X1 U9559 ( .A(n14391), .B(n14392), .ZN(n15402) );
  XNOR2_X1 U9560 ( .A(n6935), .B(n6934), .ZN(n12448) );
  NOR2_X1 U9561 ( .A1(n10939), .A2(n15056), .ZN(n10941) );
  NAND2_X4 U9562 ( .A1(n7259), .A2(n7257), .ZN(n11622) );
  NAND2_X1 U9563 ( .A1(n7575), .A2(n8184), .ZN(n8187) );
  OAI21_X1 U9564 ( .B1(n9619), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n7654), .ZN(
        n7655) );
  NOR2_X1 U9565 ( .A1(n11404), .A2(n8798), .ZN(n12318) );
  NAND2_X1 U9566 ( .A1(n7807), .A2(n8363), .ZN(n7808) );
  NAND2_X1 U9567 ( .A1(n10162), .A2(n7807), .ZN(n10007) );
  XNOR2_X1 U9568 ( .A(n7807), .B(n11584), .ZN(n9916) );
  AND2_X1 U9569 ( .A1(n7807), .A2(n15019), .ZN(n6937) );
  AND2_X1 U9570 ( .A1(n10166), .A2(n7807), .ZN(n6938) );
  NAND2_X1 U9571 ( .A1(n11221), .A2(n6940), .ZN(n6944) );
  INV_X1 U9572 ( .A(n13229), .ZN(n6942) );
  NAND2_X1 U9573 ( .A1(n6942), .A2(n6943), .ZN(n13206) );
  NAND2_X1 U9574 ( .A1(n14447), .A2(n6953), .ZN(n6950) );
  NAND2_X1 U9575 ( .A1(n6950), .A2(n6951), .ZN(n14249) );
  NAND2_X1 U9576 ( .A1(n11531), .A2(n6968), .ZN(n6967) );
  NAND2_X1 U9577 ( .A1(n14684), .A2(n9270), .ZN(n11063) );
  NAND2_X1 U9578 ( .A1(n13484), .A2(n6978), .ZN(n6977) );
  OAI211_X1 U9579 ( .C1(n13484), .C2(n6979), .A(n13380), .B(n6977), .ZN(
        P1_U3214) );
  NAND2_X1 U9580 ( .A1(n11109), .A2(n6996), .ZN(n6993) );
  NAND2_X1 U9581 ( .A1(n6993), .A2(n6994), .ZN(n11019) );
  NAND2_X1 U9582 ( .A1(n12631), .A2(n7002), .ZN(n6999) );
  NAND2_X1 U9583 ( .A1(n6999), .A2(n7000), .ZN(n12600) );
  NAND2_X1 U9584 ( .A1(n7541), .A2(n7539), .ZN(n9054) );
  OAI21_X1 U9585 ( .B1(n13153), .B2(n7017), .A(n7014), .ZN(n13103) );
  NOR2_X2 U9586 ( .A1(n13039), .A2(n7032), .ZN(n13026) );
  NAND2_X2 U9587 ( .A1(n7993), .A2(n7992), .ZN(n11376) );
  NAND2_X1 U9588 ( .A1(n7970), .A2(n7676), .ZN(n7989) );
  MUX2_X1 U9589 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n9155), .Z(n7034) );
  NAND2_X1 U9590 ( .A1(n7037), .A2(n7036), .ZN(n7035) );
  INV_X1 U9591 ( .A(n8111), .ZN(n7037) );
  NOR2_X1 U9592 ( .A1(n7942), .A2(n7941), .ZN(n7943) );
  AOI21_X1 U9593 ( .B1(n7046), .B2(n7534), .A(n6578), .ZN(n7044) );
  NAND2_X1 U9594 ( .A1(n8066), .A2(n7046), .ZN(n7045) );
  INV_X1 U9595 ( .A(n7853), .ZN(n7050) );
  NAND2_X1 U9596 ( .A1(n7834), .A2(n7833), .ZN(n7053) );
  NOR2_X1 U9597 ( .A1(n8270), .A2(n8269), .ZN(n8271) );
  INV_X1 U9598 ( .A(n8224), .ZN(n7054) );
  AND3_X2 U9599 ( .A1(n7703), .A2(n7702), .A3(n7729), .ZN(n8007) );
  XNOR2_X2 U9600 ( .A(n11585), .B(n11586), .ZN(n12785) );
  NAND2_X1 U9601 ( .A1(n7059), .A2(n6593), .ZN(n7063) );
  CLKBUF_X1 U9602 ( .A(n7063), .Z(n7060) );
  INV_X1 U9603 ( .A(n11557), .ZN(n7064) );
  NAND2_X1 U9604 ( .A1(n12827), .A2(n7393), .ZN(n7067) );
  NAND2_X1 U9605 ( .A1(n11566), .A2(n11565), .ZN(n7070) );
  MUX2_X1 U9606 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n9155), .Z(n7072) );
  NAND2_X1 U9607 ( .A1(n15143), .A2(n10268), .ZN(n15147) );
  AND2_X1 U9608 ( .A1(n7078), .A2(n10985), .ZN(n11988) );
  NOR2_X1 U9609 ( .A1(n11989), .A2(n7079), .ZN(n7078) );
  NAND2_X1 U9610 ( .A1(n7081), .A2(n15123), .ZN(n7080) );
  INV_X1 U9611 ( .A(n10986), .ZN(n7081) );
  AND2_X1 U9612 ( .A1(n10326), .A2(n10324), .ZN(n7082) );
  NAND2_X1 U9613 ( .A1(n11981), .A2(n6487), .ZN(n7084) );
  NAND2_X1 U9614 ( .A1(n10620), .A2(n7098), .ZN(n7093) );
  NAND3_X1 U9615 ( .A1(n7096), .A2(n7100), .A3(n7093), .ZN(n10621) );
  NAND2_X1 U9616 ( .A1(n10722), .A2(n10469), .ZN(n7101) );
  NAND2_X1 U9617 ( .A1(n8686), .A2(n8522), .ZN(n8524) );
  NAND2_X1 U9618 ( .A1(n8881), .A2(n8550), .ZN(n7113) );
  INV_X1 U9619 ( .A(n7665), .ZN(n7122) );
  NAND2_X1 U9620 ( .A1(n7675), .A2(n7124), .ZN(n7123) );
  INV_X1 U9621 ( .A(n7197), .ZN(n7129) );
  NAND3_X1 U9622 ( .A1(n7133), .A2(n7132), .A3(n9446), .ZN(n14025) );
  NAND2_X1 U9623 ( .A1(n14045), .A2(n14054), .ZN(n14044) );
  NAND2_X1 U9624 ( .A1(n7197), .A2(n7198), .ZN(n14045) );
  NAND3_X1 U9625 ( .A1(n7626), .A2(n7687), .A3(n7624), .ZN(n7135) );
  AND2_X2 U9626 ( .A1(n7140), .A2(n7139), .ZN(n14168) );
  OAI21_X1 U9627 ( .B1(SI_6_), .B2(n7143), .A(n7667), .ZN(n7666) );
  MUX2_X1 U9628 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n9155), .Z(n7143) );
  AND2_X2 U9629 ( .A1(n7144), .A2(n9158), .ZN(n9201) );
  NAND2_X4 U9630 ( .A1(n9429), .A2(n7171), .ZN(n13514) );
  NAND2_X2 U9631 ( .A1(n9567), .A2(n14617), .ZN(n9429) );
  XNOR2_X2 U9632 ( .A(n7145), .B(n9154), .ZN(n14617) );
  NOR2_X2 U9633 ( .A1(n14143), .A2(n14235), .ZN(n14142) );
  NAND2_X1 U9634 ( .A1(n10722), .A2(n10468), .ZN(n7163) );
  NAND2_X1 U9635 ( .A1(n10705), .A2(n10444), .ZN(n10445) );
  NOR2_X2 U9636 ( .A1(n10039), .A2(n10128), .ZN(n10132) );
  NAND2_X1 U9637 ( .A1(n10702), .A2(n10453), .ZN(n10454) );
  NAND2_X1 U9638 ( .A1(n10661), .A2(n10659), .ZN(n7182) );
  NAND2_X1 U9639 ( .A1(n9395), .A2(n9394), .ZN(n14107) );
  OAI211_X2 U9640 ( .C1(n9429), .C2(n13819), .A(n7184), .B(n7183), .ZN(n14757)
         );
  OR2_X1 U9641 ( .A1(n9272), .A2(n9648), .ZN(n7183) );
  OR2_X1 U9642 ( .A1(n13514), .A2(n9628), .ZN(n7184) );
  NAND2_X1 U9643 ( .A1(n13997), .A2(n13998), .ZN(n13996) );
  AOI21_X1 U9644 ( .B1(n14702), .B2(n13522), .A(n9231), .ZN(n10759) );
  NAND2_X1 U9645 ( .A1(n7191), .A2(n7192), .ZN(n14702) );
  NAND2_X1 U9646 ( .A1(n14090), .A2(n7200), .ZN(n7197) );
  INV_X1 U9647 ( .A(n9427), .ZN(n7207) );
  NAND3_X1 U9648 ( .A1(n15146), .A2(n8656), .A3(n8667), .ZN(n7209) );
  NAND2_X1 U9649 ( .A1(n15146), .A2(n8656), .ZN(n15127) );
  NAND3_X1 U9650 ( .A1(n11871), .A2(n6439), .A3(P3_REG0_REG_1__SCAN_IN), .ZN(
        n7215) );
  NAND2_X2 U9651 ( .A1(n11871), .A2(n6439), .ZN(n7219) );
  NOR2_X1 U9652 ( .A1(n6439), .A2(n10412), .ZN(n7216) );
  NAND2_X2 U9653 ( .A1(n6439), .A2(n8615), .ZN(n10860) );
  NAND3_X1 U9654 ( .A1(n6439), .A2(n8615), .A3(P3_REG2_REG_1__SCAN_IN), .ZN(
        n7217) );
  NAND2_X1 U9655 ( .A1(n7226), .A2(n7224), .ZN(n8795) );
  NAND2_X1 U9656 ( .A1(n8741), .A2(n7228), .ZN(n7226) );
  INV_X1 U9657 ( .A(n11022), .ZN(n11020) );
  NAND2_X1 U9658 ( .A1(n12555), .A2(n7233), .ZN(n7232) );
  NAND2_X1 U9659 ( .A1(n12482), .A2(n8989), .ZN(n7247) );
  NAND2_X1 U9660 ( .A1(n7251), .A2(n8897), .ZN(n8610) );
  NAND2_X1 U9661 ( .A1(n9085), .A2(n7263), .ZN(n7257) );
  AOI21_X2 U9662 ( .B1(n9908), .B2(n7261), .A(n7260), .ZN(n7259) );
  NOR2_X1 U9663 ( .A1(n12108), .A2(n7262), .ZN(n7261) );
  INV_X1 U9664 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n7262) );
  NAND2_X1 U9665 ( .A1(n12023), .A2(n6485), .ZN(n7268) );
  OR2_X2 U9666 ( .A1(n7757), .A2(n7279), .ZN(n8169) );
  NOR2_X2 U9667 ( .A1(n7757), .A2(n7758), .ZN(n7816) );
  NAND2_X1 U9668 ( .A1(n7291), .A2(n10895), .ZN(n11190) );
  OAI21_X1 U9669 ( .B1(n10915), .B2(n10879), .A(n7293), .ZN(n7291) );
  NAND2_X1 U9670 ( .A1(n13073), .A2(n7298), .ZN(n7296) );
  OAI21_X1 U9671 ( .B1(n13073), .B2(n7300), .A(n7298), .ZN(n7303) );
  INV_X1 U9672 ( .A(n7303), .ZN(n13041) );
  INV_X1 U9673 ( .A(n11694), .ZN(n7305) );
  NAND2_X1 U9674 ( .A1(n7307), .A2(n7306), .ZN(n10239) );
  AOI21_X1 U9675 ( .B1(n7308), .B2(n10126), .A(n6525), .ZN(n7306) );
  NAND3_X1 U9676 ( .A1(n10037), .A2(n10036), .A3(n10126), .ZN(n7307) );
  NAND2_X1 U9677 ( .A1(n10037), .A2(n10036), .ZN(n7309) );
  INV_X1 U9678 ( .A(n10007), .ZN(n7308) );
  NAND2_X1 U9679 ( .A1(n11359), .A2(n6563), .ZN(n7311) );
  NAND2_X1 U9680 ( .A1(n7706), .A2(n6468), .ZN(n7317) );
  NAND2_X1 U9681 ( .A1(n7706), .A2(n7316), .ZN(n7743) );
  NAND2_X2 U9682 ( .A1(n11687), .A2(n11686), .ZN(n13153) );
  INV_X1 U9683 ( .A(n10913), .ZN(n10876) );
  NAND2_X1 U9684 ( .A1(n13610), .A2(n13611), .ZN(n13609) );
  NAND2_X1 U9685 ( .A1(n7369), .A2(n7372), .ZN(n13597) );
  NAND3_X1 U9686 ( .A1(n13588), .A2(n13589), .A3(n7370), .ZN(n7369) );
  NAND2_X1 U9687 ( .A1(n13621), .A2(n13622), .ZN(n13620) );
  NAND2_X1 U9688 ( .A1(n7426), .A2(n9201), .ZN(n9379) );
  AND2_X1 U9689 ( .A1(n7426), .A2(n7376), .ZN(n9383) );
  OAI21_X1 U9690 ( .B1(n11049), .B2(n11042), .A(n11047), .ZN(n11179) );
  NAND2_X1 U9691 ( .A1(n7386), .A2(n7382), .ZN(n11182) );
  NAND2_X1 U9692 ( .A1(n11042), .A2(n11047), .ZN(n7385) );
  OR2_X1 U9693 ( .A1(n11180), .A2(n11181), .ZN(n7387) );
  NAND2_X1 U9694 ( .A1(n11589), .A2(n7388), .ZN(n12808) );
  AOI21_X1 U9695 ( .B1(n7390), .B2(n12840), .A(n12902), .ZN(n12841) );
  NAND2_X1 U9696 ( .A1(n12872), .A2(n7395), .ZN(n12855) );
  OR2_X1 U9697 ( .A1(n12854), .A2(n11572), .ZN(n7392) );
  NOR2_X1 U9698 ( .A1(n12854), .A2(n7394), .ZN(n7393) );
  INV_X1 U9699 ( .A(n7395), .ZN(n7394) );
  OAI21_X1 U9700 ( .B1(n12813), .B2(n7399), .A(n7396), .ZN(n11611) );
  NAND2_X1 U9701 ( .A1(n7403), .A2(n9615), .ZN(P1_U3525) );
  OAI21_X1 U9702 ( .B1(n9612), .B2(n14808), .A(n9613), .ZN(n7403) );
  NAND2_X1 U9703 ( .A1(n11341), .A2(n7405), .ZN(n7404) );
  INV_X1 U9704 ( .A(n14031), .ZN(n7411) );
  INV_X1 U9705 ( .A(n13979), .ZN(n7412) );
  NAND2_X1 U9706 ( .A1(n13979), .A2(n6448), .ZN(n7413) );
  NAND2_X1 U9707 ( .A1(n7413), .A2(n7414), .ZN(n9555) );
  OAI21_X1 U9708 ( .B1(n11533), .B2(n7421), .A(n7419), .ZN(n14121) );
  NAND2_X1 U9709 ( .A1(n7418), .A2(n7416), .ZN(n9546) );
  NAND2_X1 U9710 ( .A1(n11533), .A2(n7419), .ZN(n7418) );
  OAI211_X1 U9711 ( .C1(n10221), .C2(n7433), .A(n7432), .B(n7430), .ZN(n14700)
         );
  NAND2_X1 U9712 ( .A1(n11501), .A2(n6567), .ZN(n9544) );
  NAND2_X1 U9713 ( .A1(n10757), .A2(n6556), .ZN(n7436) );
  NAND3_X1 U9714 ( .A1(n7444), .A2(n7445), .A3(n7443), .ZN(n7441) );
  AND2_X1 U9715 ( .A1(n9140), .A2(n6580), .ZN(n9144) );
  NAND2_X1 U9716 ( .A1(n9140), .A2(n7452), .ZN(n14299) );
  NAND2_X1 U9717 ( .A1(n7455), .A2(n10050), .ZN(n10051) );
  NAND2_X1 U9718 ( .A1(n9986), .A2(n9985), .ZN(n7455) );
  OAI21_X1 U9719 ( .B1(n9985), .B2(n9986), .A(n7455), .ZN(n9990) );
  NAND3_X1 U9720 ( .A1(n7460), .A2(n7464), .A3(n7459), .ZN(n7458) );
  NAND2_X1 U9721 ( .A1(n13389), .A2(n7469), .ZN(n13390) );
  NAND2_X1 U9722 ( .A1(n7465), .A2(n13389), .ZN(n7464) );
  NOR2_X1 U9723 ( .A1(n7470), .A2(n10297), .ZN(n7465) );
  NAND2_X1 U9724 ( .A1(n13390), .A2(n7467), .ZN(n10528) );
  NAND2_X1 U9725 ( .A1(n13391), .A2(n13388), .ZN(n7470) );
  OAI211_X1 U9726 ( .C1(n13484), .C2(n7481), .A(n7478), .B(n7477), .ZN(n11849)
         );
  NAND2_X1 U9727 ( .A1(n13484), .A2(n6566), .ZN(n7477) );
  OAI22_X1 U9728 ( .A1(n7480), .A2(n7479), .B1(n7485), .B2(n7482), .ZN(n7478)
         );
  INV_X1 U9729 ( .A(n7482), .ZN(n7479) );
  NAND2_X1 U9730 ( .A1(n10847), .A2(n7650), .ZN(n10848) );
  INV_X1 U9731 ( .A(n7495), .ZN(n11005) );
  NOR2_X1 U9732 ( .A1(n10849), .A2(n7497), .ZN(n7496) );
  INV_X1 U9733 ( .A(n7650), .ZN(n7497) );
  NAND2_X1 U9734 ( .A1(n13473), .A2(n6596), .ZN(n13401) );
  NAND2_X1 U9735 ( .A1(n9383), .A2(n6560), .ZN(n9571) );
  NAND2_X1 U9736 ( .A1(n7717), .A2(n7503), .ZN(n8493) );
  AND2_X1 U9737 ( .A1(n7830), .A2(n7832), .ZN(n7514) );
  INV_X1 U9738 ( .A(n8158), .ZN(n7515) );
  AOI21_X1 U9739 ( .B1(n7515), .B2(n6592), .A(n7516), .ZN(n8179) );
  INV_X1 U9740 ( .A(n7899), .ZN(n7525) );
  NAND2_X1 U9741 ( .A1(n6469), .A2(n6838), .ZN(n8786) );
  NAND2_X1 U9742 ( .A1(n14503), .A2(n7562), .ZN(n7559) );
  OAI21_X1 U9743 ( .B1(n11867), .B2(n14498), .A(n7569), .ZN(P3_U3204) );
  XNOR2_X1 U9744 ( .A(n12078), .B(n9059), .ZN(n11864) );
  INV_X1 U9745 ( .A(n7578), .ZN(n7577) );
  NAND3_X1 U9746 ( .A1(n7582), .A2(n7581), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n7584) );
  NAND2_X1 U9747 ( .A1(n13501), .A2(n13511), .ZN(n7591) );
  NAND2_X1 U9748 ( .A1(n7591), .A2(n13502), .ZN(n13936) );
  XNOR2_X1 U9749 ( .A(n7593), .B(n7592), .ZN(n13752) );
  INV_X1 U9750 ( .A(n7593), .ZN(n13751) );
  NAND2_X1 U9751 ( .A1(n8208), .A2(n7598), .ZN(n7596) );
  NAND2_X1 U9752 ( .A1(n8208), .A2(n8207), .ZN(n7597) );
  NAND2_X1 U9753 ( .A1(n8373), .A2(n7603), .ZN(n7601) );
  NAND2_X1 U9754 ( .A1(n7601), .A2(n7602), .ZN(n8381) );
  OAI21_X1 U9755 ( .B1(n8373), .B2(n7608), .A(n7605), .ZN(n8422) );
  NAND2_X1 U9756 ( .A1(n8373), .A2(n8372), .ZN(n8390) );
  INV_X1 U9757 ( .A(n7626), .ZN(n7625) );
  NAND2_X1 U9758 ( .A1(n7687), .A2(n7686), .ZN(n8046) );
  INV_X1 U9759 ( .A(n8045), .ZN(n7630) );
  NAND2_X1 U9760 ( .A1(n13976), .A2(n9507), .ZN(n9509) );
  NAND2_X1 U9761 ( .A1(n12662), .A2(n7631), .ZN(n12728) );
  INV_X1 U9762 ( .A(n12657), .ZN(n12662) );
  NAND2_X1 U9763 ( .A1(n14249), .A2(n13653), .ZN(n11531) );
  NAND2_X1 U9764 ( .A1(n9528), .A2(n9527), .ZN(n10575) );
  OR2_X1 U9765 ( .A1(n12658), .A2(n14530), .ZN(n12661) );
  NAND2_X1 U9766 ( .A1(n12457), .A2(n15149), .ZN(n12460) );
  NAND2_X1 U9767 ( .A1(n9124), .A2(n15206), .ZN(n9111) );
  NAND2_X1 U9768 ( .A1(n8610), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8612) );
  NAND4_X4 U9769 ( .A1(n9170), .A2(n9169), .A3(n9168), .A4(n9167), .ZN(n14729)
         );
  XNOR2_X1 U9770 ( .A(n9980), .B(n11838), .ZN(n9983) );
  NAND2_X1 U9771 ( .A1(n13963), .A2(n14730), .ZN(n9570) );
  NAND2_X1 U9772 ( .A1(n9971), .A2(n9709), .ZN(n13766) );
  OAI21_X1 U9773 ( .B1(n8509), .B2(n6795), .A(n7645), .ZN(n8512) );
  INV_X1 U9774 ( .A(n11864), .ZN(n9067) );
  INV_X1 U9775 ( .A(n8321), .ZN(n8319) );
  INV_X1 U9776 ( .A(n13936), .ZN(n14257) );
  NOR2_X1 U9777 ( .A1(n12456), .A2(n12455), .ZN(n7632) );
  AND2_X2 U9778 ( .A1(n10265), .A2(n9123), .ZN(n15222) );
  INV_X1 U9779 ( .A(n10181), .ZN(n10193) );
  AND2_X1 U9780 ( .A1(n15153), .A2(n12663), .ZN(n14530) );
  INV_X1 U9781 ( .A(n14530), .ZN(n9066) );
  XOR2_X1 U9782 ( .A(n15139), .B(n11622), .Z(n7633) );
  AND2_X1 U9783 ( .A1(n13798), .A2(n14757), .ZN(n7634) );
  OR2_X1 U9784 ( .A1(n13798), .A2(n14757), .ZN(n7635) );
  INV_X1 U9785 ( .A(n15026), .ZN(n15037) );
  AND2_X2 U9786 ( .A1(n10016), .A2(n10015), .ZN(n15026) );
  NAND2_X1 U9787 ( .A1(n10016), .A2(n9782), .ZN(n15045) );
  AND2_X1 U9788 ( .A1(n12459), .A2(n7639), .ZN(n7637) );
  AND2_X1 U9789 ( .A1(n15219), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n7638) );
  NAND2_X2 U9790 ( .A1(n10083), .A2(n13217), .ZN(n13219) );
  OR2_X1 U9791 ( .A1(n12458), .A2(n12646), .ZN(n7639) );
  AND2_X1 U9792 ( .A1(n10685), .A2(n10473), .ZN(n7640) );
  INV_X1 U9793 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7708) );
  OR2_X1 U9794 ( .A1(n9687), .A2(n9885), .ZN(n7641) );
  INV_X1 U9795 ( .A(n10869), .ZN(n10912) );
  XOR2_X1 U9796 ( .A(n12992), .B(n8451), .Z(n7642) );
  INV_X1 U9797 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n11850) );
  INV_X1 U9798 ( .A(n8725), .ZN(n12092) );
  AND2_X1 U9799 ( .A1(n10010), .A2(n7773), .ZN(n7643) );
  INV_X1 U9800 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7710) );
  NAND2_X1 U9801 ( .A1(n10502), .A2(n14708), .ZN(n14691) );
  INV_X1 U9802 ( .A(n11622), .ZN(n11643) );
  AND3_X1 U9803 ( .A1(n13961), .A2(n13949), .A3(n13956), .ZN(n7644) );
  INV_X1 U9804 ( .A(n13735), .ZN(n13957) );
  AND4_X1 U9805 ( .A1(n8483), .A2(n6914), .A3(n8505), .A4(n11445), .ZN(n7645)
         );
  OR2_X1 U9806 ( .A1(n8181), .A2(n8180), .ZN(n7647) );
  OR2_X1 U9807 ( .A1(n8116), .A2(SI_17_), .ZN(n7648) );
  AND2_X1 U9808 ( .A1(n8368), .A2(n8367), .ZN(n7649) );
  INV_X1 U9809 ( .A(n13980), .ZN(n9554) );
  INV_X1 U9810 ( .A(n14282), .ZN(n9614) );
  NAND2_X1 U9811 ( .A1(n7792), .A2(n7791), .ZN(n7811) );
  OAI21_X1 U9812 ( .B1(n10431), .B2(n8419), .A(n7831), .ZN(n7835) );
  MUX2_X1 U9813 ( .A(n13580), .B(n13579), .S(n13732), .Z(n13581) );
  OAI21_X1 U9814 ( .B1(n13642), .B2(n13643), .A(n13644), .ZN(n13639) );
  INV_X1 U9815 ( .A(n13639), .ZN(n13640) );
  OAI21_X1 U9816 ( .B1(n13687), .B2(n13688), .A(n13686), .ZN(n13690) );
  INV_X1 U9817 ( .A(n8204), .ZN(n8205) );
  NAND2_X1 U9818 ( .A1(n12127), .A2(n10181), .ZN(n10194) );
  AND4_X1 U9819 ( .A1(n8582), .A2(n8581), .A3(n9025), .A4(n7276), .ZN(n8583)
         );
  AND2_X1 U9820 ( .A1(n8417), .A2(n8416), .ZN(n8418) );
  INV_X1 U9821 ( .A(n11737), .ZN(n11740) );
  INV_X1 U9822 ( .A(n13377), .ZN(n9506) );
  INV_X1 U9823 ( .A(n8206), .ZN(n8207) );
  INV_X1 U9824 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n12024) );
  INV_X1 U9825 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8576) );
  XNOR2_X1 U9826 ( .A(n13237), .B(n12986), .ZN(n8477) );
  NAND2_X1 U9827 ( .A1(n8477), .A2(n8418), .ZN(n8445) );
  INV_X1 U9828 ( .A(n8096), .ZN(n7753) );
  INV_X1 U9829 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8014) );
  INV_X1 U9830 ( .A(n13184), .ZN(n11709) );
  NAND2_X1 U9831 ( .A1(n11215), .A2(n11214), .ZN(n11359) );
  INV_X1 U9832 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7721) );
  NAND2_X1 U9833 ( .A1(n14263), .A2(n9506), .ZN(n9507) );
  INV_X1 U9834 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8545) );
  AND2_X1 U9835 ( .A1(n7801), .A2(SI_2_), .ZN(n7658) );
  INV_X1 U9836 ( .A(n8968), .ZN(n8604) );
  NAND2_X1 U9837 ( .A1(n7633), .A2(n7212), .ZN(n10271) );
  NAND2_X1 U9838 ( .A1(n12659), .A2(n9001), .ZN(n9002) );
  OR2_X1 U9839 ( .A1(n8565), .A2(n13368), .ZN(n8566) );
  INV_X1 U9840 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7740) );
  OR2_X1 U9841 ( .A1(n8300), .A2(n8285), .ZN(n8353) );
  NAND2_X1 U9842 ( .A1(n8165), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8191) );
  AND2_X1 U9843 ( .A1(n11302), .A2(n14944), .ZN(n11304) );
  NAND2_X1 U9844 ( .A1(n8122), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8150) );
  INV_X1 U9845 ( .A(n9779), .ZN(n9734) );
  INV_X1 U9846 ( .A(n15377), .ZN(n11745) );
  OR2_X1 U9847 ( .A1(n11798), .A2(n11797), .ZN(n11799) );
  OR2_X1 U9848 ( .A1(n11775), .A2(n11774), .ZN(n11776) );
  OR2_X1 U9849 ( .A1(n11760), .A2(n11759), .ZN(n11761) );
  INV_X1 U9850 ( .A(n11826), .ZN(n11835) );
  INV_X1 U9851 ( .A(n9431), .ZN(n9432) );
  OR2_X1 U9852 ( .A1(n9249), .A2(n10850), .ZN(n9262) );
  INV_X1 U9853 ( .A(n9440), .ZN(n9449) );
  AND2_X1 U9854 ( .A1(n9370), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9387) );
  NOR2_X1 U9855 ( .A1(n9320), .A2(n9319), .ZN(n9335) );
  INV_X1 U9856 ( .A(n13782), .ZN(n13672) );
  AND2_X1 U9857 ( .A1(n8377), .A2(n8376), .ZN(n8389) );
  OR2_X1 U9858 ( .A1(n14336), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n14335) );
  NOR2_X1 U9859 ( .A1(n14367), .A2(n14366), .ZN(n14343) );
  INV_X1 U9860 ( .A(n12456), .ZN(n12461) );
  NAND2_X1 U9861 ( .A1(n8604), .A2(n8603), .ZN(n8980) );
  INV_X1 U9862 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10463) );
  INV_X1 U9863 ( .A(n9038), .ZN(n10210) );
  OR2_X1 U9864 ( .A1(n10211), .A2(n10210), .ZN(n12065) );
  INV_X1 U9865 ( .A(n9013), .ZN(n11863) );
  INV_X1 U9866 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n11878) );
  AND2_X1 U9867 ( .A1(n10419), .A2(n10417), .ZN(n10407) );
  OR2_X1 U9868 ( .A1(n14437), .A2(n12428), .ZN(n9120) );
  AND2_X1 U9869 ( .A1(n10181), .A2(n12442), .ZN(n15140) );
  OR2_X1 U9870 ( .A1(n10261), .A2(n10195), .ZN(n9115) );
  AND2_X1 U9871 ( .A1(n10863), .A2(n10862), .ZN(n12450) );
  NAND2_X1 U9872 ( .A1(n9070), .A2(n9069), .ZN(n9073) );
  INV_X1 U9873 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8842) );
  AND2_X1 U9874 ( .A1(n8536), .A2(n8535), .ZN(n8782) );
  OR2_X1 U9875 ( .A1(n8235), .A2(n8234), .ZN(n8260) );
  OR2_X1 U9876 ( .A1(n8191), .A2(n8190), .ZN(n8215) );
  NAND2_X1 U9877 ( .A1(n10520), .A2(n10519), .ZN(n10777) );
  INV_X1 U9878 ( .A(n13105), .ZN(n12861) );
  AND2_X1 U9879 ( .A1(n9918), .A2(n9954), .ZN(n9922) );
  OR2_X1 U9880 ( .A1(n11613), .A2(n13139), .ZN(n12896) );
  AND2_X1 U9881 ( .A1(n11728), .A2(n8327), .ZN(n13006) );
  OR2_X1 U9882 ( .A1(n8150), .A2(n8149), .ZN(n8167) );
  INV_X1 U9883 ( .A(n8356), .ZN(n8328) );
  OR2_X1 U9884 ( .A1(n9882), .A2(n9883), .ZN(n11294) );
  OR2_X1 U9885 ( .A1(n14900), .A2(n14899), .ZN(n14902) );
  OR2_X1 U9886 ( .A1(n11304), .A2(n11303), .ZN(n14937) );
  OR2_X1 U9887 ( .A1(n14967), .A2(n14966), .ZN(n14963) );
  AND2_X1 U9888 ( .A1(n9697), .A2(n13351), .ZN(n9691) );
  NAND2_X1 U9889 ( .A1(n8498), .A2(n9744), .ZN(n13139) );
  INV_X1 U9890 ( .A(n13399), .ZN(n11781) );
  INV_X1 U9891 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10850) );
  INV_X1 U9892 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9212) );
  INV_X1 U9893 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9292) );
  AND2_X1 U9894 ( .A1(n13555), .A2(n9801), .ZN(n13478) );
  NOR2_X1 U9895 ( .A1(n9409), .A2(n13459), .ZN(n9417) );
  INV_X1 U9896 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10749) );
  OR2_X1 U9897 ( .A1(n14627), .A2(n9807), .ZN(n14672) );
  NAND2_X1 U9898 ( .A1(n9584), .A2(n9707), .ZN(n10500) );
  NAND2_X1 U9899 ( .A1(n10496), .A2(n10495), .ZN(n14708) );
  INV_X1 U9900 ( .A(n14822), .ZN(n9605) );
  OR2_X1 U9901 ( .A1(n10505), .A2(n14082), .ZN(n10573) );
  AOI21_X1 U9902 ( .B1(n9529), .B2(n7635), .A(n7634), .ZN(n10223) );
  XNOR2_X1 U9903 ( .A(n8381), .B(n8380), .ZN(n13501) );
  INV_X1 U9904 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9520) );
  AOI22_X1 U9905 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14336), .B1(n14387), .B2(
        n14335), .ZN(n14338) );
  OAI22_X1 U9906 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14351), .B1(n14360), 
        .B2(n14350), .ZN(n14410) );
  AND2_X1 U9907 ( .A1(n9097), .A2(n9096), .ZN(n9099) );
  INV_X1 U9908 ( .A(n11619), .ZN(n14524) );
  INV_X1 U9909 ( .A(n12065), .ZN(n12050) );
  AND2_X1 U9910 ( .A1(n10209), .A2(n10210), .ZN(n12062) );
  INV_X1 U9911 ( .A(n12068), .ZN(n12036) );
  NAND2_X1 U9912 ( .A1(n10192), .A2(n10191), .ZN(n12071) );
  INV_X1 U9913 ( .A(n8644), .ZN(n9014) );
  AND2_X1 U9914 ( .A1(n8952), .A2(n8951), .ZN(n12533) );
  AND4_X1 U9915 ( .A1(n8836), .A2(n8835), .A3(n8834), .A4(n8833), .ZN(n12643)
         );
  MUX2_X1 U9916 ( .A(n10407), .B(P3_U3897), .S(n12268), .Z(n15084) );
  INV_X1 U9917 ( .A(n15074), .ZN(n15100) );
  INV_X1 U9918 ( .A(n12090), .ZN(n12518) );
  INV_X1 U9919 ( .A(n12653), .ZN(n12635) );
  NAND2_X1 U9920 ( .A1(n10265), .A2(n10264), .ZN(n10267) );
  AND3_X1 U9921 ( .A1(n9115), .A2(n9114), .A3(n9113), .ZN(n10265) );
  INV_X1 U9922 ( .A(n12663), .ZN(n15203) );
  INV_X1 U9923 ( .A(n9085), .ZN(n9784) );
  INV_X1 U9924 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8913) );
  AND2_X1 U9925 ( .A1(n8859), .A2(n8882), .ZN(n12370) );
  INV_X1 U9926 ( .A(n12890), .ZN(n12848) );
  NAND2_X1 U9927 ( .A1(n9735), .A2(n13217), .ZN(n12900) );
  OR2_X1 U9928 ( .A1(n13095), .A2(n8356), .ZN(n8221) );
  INV_X1 U9929 ( .A(n6441), .ZN(n8432) );
  NAND2_X1 U9930 ( .A1(n6442), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7795) );
  INV_X1 U9931 ( .A(n14960), .ZN(n14977) );
  INV_X1 U9932 ( .A(n14985), .ZN(n14965) );
  OR2_X1 U9933 ( .A1(n14925), .A2(n14924), .ZN(n14931) );
  INV_X1 U9934 ( .A(n14979), .ZN(n14971) );
  AND2_X1 U9935 ( .A1(n10894), .A2(n10871), .ZN(n11088) );
  INV_X1 U9936 ( .A(n13141), .ZN(n13223) );
  NOR2_X1 U9937 ( .A1(n14994), .A2(n10081), .ZN(n9782) );
  AND2_X1 U9938 ( .A1(n9771), .A2(n15023), .ZN(n13327) );
  AND2_X1 U9939 ( .A1(n10014), .A2(n14994), .ZN(n10015) );
  AND2_X1 U9940 ( .A1(n9724), .A2(n9723), .ZN(n14990) );
  OR2_X1 U9941 ( .A1(n9293), .A2(n9292), .ZN(n9320) );
  INV_X1 U9942 ( .A(n15379), .ZN(n14564) );
  OR2_X1 U9943 ( .A1(n9991), .A2(n9969), .ZN(n9989) );
  AND4_X1 U9944 ( .A1(n9505), .A2(n9504), .A3(n9503), .A4(n9502), .ZN(n13377)
         );
  INV_X1 U9945 ( .A(n13799), .ZN(n14666) );
  OR2_X1 U9946 ( .A1(n13663), .A2(n6491), .ZN(n14136) );
  INV_X1 U9947 ( .A(n9534), .ZN(n13523) );
  INV_X1 U9948 ( .A(n14696), .ZN(n14742) );
  INV_X1 U9949 ( .A(n14205), .ZN(n9609) );
  INV_X1 U9950 ( .A(n10582), .ZN(n13950) );
  INV_X1 U9951 ( .A(n10573), .ZN(n14793) );
  NAND2_X1 U9952 ( .A1(n9604), .A2(n9704), .ZN(n10582) );
  INV_X1 U9953 ( .A(n13766), .ZN(n10496) );
  INV_X1 U9954 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9154) );
  INV_X1 U9955 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9522) );
  XNOR2_X1 U9956 ( .A(n9331), .B(P1_IR_REG_14__SCAN_IN), .ZN(n13894) );
  INV_X1 U9957 ( .A(n9713), .ZN(n9909) );
  NAND2_X1 U9958 ( .A1(n10213), .A2(n10266), .ZN(n12068) );
  AND2_X1 U9959 ( .A1(n10863), .A2(n9018), .ZN(n12458) );
  NAND2_X1 U9960 ( .A1(n8963), .A2(n8962), .ZN(n12521) );
  INV_X1 U9961 ( .A(n12066), .ZN(n12626) );
  INV_X1 U9962 ( .A(n15084), .ZN(n15068) );
  INV_X1 U9963 ( .A(n15089), .ZN(n15081) );
  OR2_X1 U9964 ( .A1(n10409), .A2(n10408), .ZN(n15097) );
  NAND2_X2 U9965 ( .A1(n10267), .A2(n15154), .ZN(n15159) );
  INV_X1 U9966 ( .A(n15222), .ZN(n15219) );
  NOR2_X1 U9967 ( .A1(n9109), .A2(n9108), .ZN(n9110) );
  INV_X1 U9968 ( .A(n12037), .ZN(n12748) );
  AND2_X1 U9969 ( .A1(n9106), .A2(n9105), .ZN(n15205) );
  NOR2_X1 U9970 ( .A1(n9784), .A2(n9909), .ZN(n10094) );
  INV_X1 U9971 ( .A(SI_14_), .ZN(n9701) );
  INV_X1 U9972 ( .A(n11072), .ZN(n11081) );
  NOR2_X1 U9973 ( .A1(n9697), .A2(P2_U3088), .ZN(n14823) );
  INV_X1 U9974 ( .A(n12888), .ZN(n12877) );
  INV_X1 U9975 ( .A(n12900), .ZN(n12883) );
  NAND2_X1 U9976 ( .A1(n8334), .A2(n8333), .ZN(n13011) );
  OAI21_X1 U9977 ( .B1(n13065), .B2(n8356), .A(n8265), .ZN(n13074) );
  INV_X1 U9978 ( .A(n14823), .ZN(n14988) );
  INV_X1 U9979 ( .A(n13234), .ZN(n13147) );
  AND2_X1 U9980 ( .A1(n13089), .A2(n13088), .ZN(n13283) );
  INV_X2 U9981 ( .A(n15045), .ZN(n15047) );
  NOR2_X1 U9982 ( .A1(n14995), .A2(n14990), .ZN(n14991) );
  INV_X1 U9983 ( .A(n14998), .ZN(n14995) );
  INV_X1 U9984 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13358) );
  INV_X1 U9985 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10179) );
  OR2_X1 U9986 ( .A1(n9991), .A2(n10501), .ZN(n15388) );
  INV_X1 U9987 ( .A(n14562), .ZN(n15382) );
  INV_X1 U9988 ( .A(n13939), .ZN(n13770) );
  OR2_X1 U9989 ( .A1(n9392), .A2(n9391), .ZN(n13782) );
  INV_X1 U9990 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14644) );
  OR2_X1 U9991 ( .A1(n14627), .A2(n13810), .ZN(n13799) );
  INV_X1 U9992 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14660) );
  INV_X1 U9993 ( .A(n14624), .ZN(n14677) );
  AND2_X1 U9994 ( .A1(n11498), .A2(n15387), .ZN(n14586) );
  OR2_X1 U9995 ( .A1(n14746), .A2(n10505), .ZN(n14461) );
  INV_X1 U9996 ( .A(n14691), .ZN(n14746) );
  AND2_X2 U9997 ( .A1(n9611), .A2(n13950), .ZN(n14822) );
  AND3_X1 U9998 ( .A1(n14586), .A2(n14585), .A3(n14584), .ZN(n14592) );
  INV_X1 U9999 ( .A(n14810), .ZN(n14808) );
  AND2_X2 U10000 ( .A1(n9611), .A2(n10582), .ZN(n14810) );
  AND2_X1 U10001 ( .A1(n9800), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9709) );
  INV_X1 U10002 ( .A(n9586), .ZN(n11546) );
  INV_X1 U10003 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11125) );
  INV_X1 U10004 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n15329) );
  NOR2_X2 U10005 ( .A1(n10186), .A2(n9909), .ZN(P3_U3897) );
  AND2_X1 U10006 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9689), .ZN(P2_U3947) );
  NOR2_X1 U10007 ( .A1(n9971), .A2(n9618), .ZN(P1_U4016) );
  INV_X1 U10008 ( .A(n7784), .ZN(n7656) );
  INV_X1 U10009 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9171) );
  INV_X1 U10010 ( .A(SI_0_), .ZN(n9640) );
  NAND2_X1 U10011 ( .A1(n7786), .A2(n7657), .ZN(n7803) );
  MUX2_X1 U10012 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n9619), .Z(n7801) );
  MUX2_X1 U10013 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n9619), .Z(n7659) );
  NAND2_X1 U10014 ( .A1(n7659), .A2(SI_3_), .ZN(n7660) );
  OAI21_X1 U10015 ( .B1(n7659), .B2(SI_3_), .A(n7660), .ZN(n7824) );
  MUX2_X1 U10016 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n9619), .Z(n7661) );
  NAND2_X1 U10017 ( .A1(n7661), .A2(SI_4_), .ZN(n7663) );
  OAI21_X1 U10018 ( .B1(n7661), .B2(SI_4_), .A(n7663), .ZN(n7838) );
  INV_X1 U10019 ( .A(n7838), .ZN(n7662) );
  INV_X2 U10020 ( .A(n9619), .ZN(n9155) );
  INV_X1 U10021 ( .A(n7664), .ZN(n7855) );
  INV_X1 U10022 ( .A(n7666), .ZN(n7883) );
  MUX2_X1 U10023 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n7171), .Z(n7669) );
  NAND2_X1 U10024 ( .A1(n7669), .A2(SI_8_), .ZN(n7671) );
  OAI21_X1 U10025 ( .B1(n7669), .B2(SI_8_), .A(n7671), .ZN(n7670) );
  INV_X1 U10026 ( .A(n7670), .ZN(n7923) );
  NAND2_X1 U10027 ( .A1(n7924), .A2(n7923), .ZN(n7926) );
  NAND2_X1 U10028 ( .A1(n7926), .A2(n7671), .ZN(n7946) );
  MUX2_X1 U10029 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n7171), .Z(n7672) );
  NAND2_X1 U10030 ( .A1(n7672), .A2(SI_9_), .ZN(n7674) );
  OAI21_X1 U10031 ( .B1(n7672), .B2(SI_9_), .A(n7674), .ZN(n7673) );
  INV_X1 U10032 ( .A(n7673), .ZN(n7945) );
  MUX2_X1 U10033 ( .A(n9770), .B(n9769), .S(n7171), .Z(n7967) );
  MUX2_X1 U10034 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n7171), .Z(n7677) );
  XNOR2_X1 U10035 ( .A(n7677), .B(SI_11_), .ZN(n7988) );
  INV_X1 U10036 ( .A(n7677), .ZN(n7678) );
  MUX2_X1 U10037 ( .A(n8539), .B(n10060), .S(n7171), .Z(n7680) );
  XNOR2_X1 U10038 ( .A(n7680), .B(SI_12_), .ZN(n8006) );
  NAND2_X1 U10039 ( .A1(n7680), .A2(n7679), .ZN(n7681) );
  MUX2_X1 U10040 ( .A(n8542), .B(n10179), .S(n7171), .Z(n7683) );
  NAND2_X1 U10041 ( .A1(n7683), .A2(n7682), .ZN(n7684) );
  NAND2_X1 U10042 ( .A1(n7685), .A2(n9701), .ZN(n7686) );
  MUX2_X1 U10043 ( .A(n8545), .B(n10510), .S(n7171), .Z(n8045) );
  MUX2_X1 U10044 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n7171), .Z(n7688) );
  MUX2_X1 U10045 ( .A(n10803), .B(n10804), .S(n9619), .Z(n7690) );
  XNOR2_X1 U10046 ( .A(n7690), .B(SI_16_), .ZN(n8086) );
  INV_X1 U10047 ( .A(SI_16_), .ZN(n7689) );
  NAND2_X1 U10048 ( .A1(n7690), .A2(n7689), .ZN(n7691) );
  MUX2_X1 U10049 ( .A(n10819), .B(n10820), .S(n7171), .Z(n8114) );
  XNOR2_X1 U10050 ( .A(n8114), .B(SI_17_), .ZN(n7692) );
  XNOR2_X1 U10051 ( .A(n8113), .B(n7692), .ZN(n10818) );
  NOR2_X1 U10052 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n7694) );
  NOR2_X1 U10053 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n7693) );
  NOR2_X1 U10054 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n7697) );
  INV_X1 U10055 ( .A(n7799), .ZN(n7703) );
  NAND2_X1 U10056 ( .A1(n6709), .A2(n7842), .ZN(n7722) );
  NOR2_X1 U10057 ( .A1(n7722), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n7702) );
  NAND2_X1 U10058 ( .A1(n10818), .A2(n8423), .ZN(n7720) );
  NOR2_X1 U10059 ( .A1(n7716), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U10060 ( .A1(n8049), .A2(n7712), .ZN(n8071) );
  INV_X1 U10061 ( .A(n8088), .ZN(n7714) );
  INV_X1 U10062 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7713) );
  NAND2_X1 U10063 ( .A1(n7714), .A2(n7713), .ZN(n8090) );
  NAND2_X1 U10064 ( .A1(n8090), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7715) );
  MUX2_X1 U10065 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7715), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n7718) );
  INV_X2 U10066 ( .A(n9687), .ZN(n8145) );
  AOI22_X1 U10067 ( .A1(n8146), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n12974), 
        .B2(n8145), .ZN(n7719) );
  INV_X1 U10068 ( .A(n7722), .ZN(n7724) );
  NAND2_X1 U10069 ( .A1(n7724), .A2(n7723), .ZN(n7725) );
  INV_X1 U10070 ( .A(n7726), .ZN(n7727) );
  NOR2_X1 U10071 ( .A1(n7727), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n7728) );
  INV_X1 U10072 ( .A(n7731), .ZN(n7732) );
  OAI21_X1 U10073 ( .B1(n7905), .B2(n7732), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n7733) );
  NAND2_X1 U10074 ( .A1(n7736), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7735) );
  MUX2_X1 U10075 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7735), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n7737) );
  NAND2_X2 U10076 ( .A1(n7737), .A2(n8479), .ZN(n11445) );
  AND2_X2 U10077 ( .A1(n11372), .A2(n9774), .ZN(n9750) );
  OAI21_X2 U10078 ( .B1(n8493), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7738) );
  XNOR2_X2 U10079 ( .A(n7738), .B(P2_IR_REG_19__SCAN_IN), .ZN(n11222) );
  AND2_X1 U10080 ( .A1(n9750), .A2(n11222), .ZN(n10250) );
  INV_X4 U10081 ( .A(n8245), .ZN(n8363) );
  NAND2_X1 U10082 ( .A1(n13307), .A2(n8363), .ZN(n7764) );
  INV_X1 U10083 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n7761) );
  NAND2_X1 U10084 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7865) );
  INV_X1 U10085 ( .A(n7865), .ZN(n7745) );
  NAND2_X1 U10086 ( .A1(n7745), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7891) );
  INV_X1 U10087 ( .A(n7891), .ZN(n7746) );
  NAND2_X1 U10088 ( .A1(n7746), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7912) );
  INV_X1 U10089 ( .A(n7912), .ZN(n7747) );
  NAND2_X1 U10090 ( .A1(n7747), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7932) );
  INV_X1 U10091 ( .A(n7932), .ZN(n7748) );
  NAND2_X1 U10092 ( .A1(n7748), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7954) );
  INV_X1 U10093 ( .A(n7954), .ZN(n7749) );
  NAND2_X1 U10094 ( .A1(n7749), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7977) );
  INV_X1 U10095 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7976) );
  INV_X1 U10096 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8054) );
  INV_X1 U10097 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8076) );
  AND2_X1 U10098 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n7752) );
  INV_X1 U10099 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7755) );
  INV_X1 U10100 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7754) );
  OAI21_X1 U10101 ( .B1(n8096), .B2(n7755), .A(n7754), .ZN(n7756) );
  NAND2_X1 U10102 ( .A1(n8124), .A2(n7756), .ZN(n13169) );
  OR2_X1 U10103 ( .A1(n13169), .A2(n8169), .ZN(n7760) );
  AND2_X2 U10104 ( .A1(n7757), .A2(n7758), .ZN(n7815) );
  AOI22_X1 U10105 ( .A1(n8385), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n7815), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n7759) );
  OAI211_X1 U10106 ( .C1(n8432), .C2(n7761), .A(n7760), .B(n7759), .ZN(n13186)
         );
  INV_X2 U10107 ( .A(n8419), .ZN(n8403) );
  NAND2_X1 U10108 ( .A1(n13186), .A2(n8403), .ZN(n7763) );
  NAND2_X1 U10109 ( .A1(n7764), .A2(n7763), .ZN(n8112) );
  NAND2_X1 U10110 ( .A1(n6442), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7768) );
  NAND2_X1 U10111 ( .A1(n7816), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7767) );
  NAND2_X1 U10112 ( .A1(n7815), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7766) );
  INV_X1 U10113 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10086) );
  OR2_X1 U10114 ( .A1(n8169), .A2(n10086), .ZN(n7765) );
  INV_X1 U10115 ( .A(n6445), .ZN(n7772) );
  INV_X1 U10116 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9694) );
  NAND2_X1 U10117 ( .A1(n7171), .A2(SI_0_), .ZN(n7769) );
  XNOR2_X1 U10118 ( .A(n7769), .B(n8513), .ZN(n13374) );
  INV_X1 U10119 ( .A(n7770), .ZN(n7771) );
  NAND2_X1 U10120 ( .A1(n7771), .A2(n9750), .ZN(n7773) );
  NAND2_X1 U10121 ( .A1(n7772), .A2(n7643), .ZN(n7776) );
  NAND2_X1 U10122 ( .A1(n10167), .A2(n8363), .ZN(n7774) );
  NAND3_X1 U10123 ( .A1(n7776), .A2(n7775), .A3(n7774), .ZN(n7812) );
  INV_X1 U10124 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7777) );
  OR2_X1 U10125 ( .A1(n8169), .A2(n7777), .ZN(n7781) );
  NAND2_X1 U10126 ( .A1(n7815), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7780) );
  NAND4_X2 U10127 ( .A1(n7781), .A2(n7780), .A3(n7779), .A4(n7778), .ZN(n9755)
         );
  NAND2_X1 U10128 ( .A1(n9755), .A2(n8427), .ZN(n7792) );
  INV_X1 U10129 ( .A(n7782), .ZN(n7783) );
  NAND2_X1 U10130 ( .A1(n7784), .A2(n7783), .ZN(n7785) );
  NAND2_X1 U10131 ( .A1(n7786), .A2(n7785), .ZN(n9654) );
  INV_X1 U10132 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9653) );
  NAND2_X1 U10133 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n7787) );
  MUX2_X1 U10134 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7787), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n7790) );
  INV_X1 U10135 ( .A(n7788), .ZN(n7789) );
  NAND2_X1 U10136 ( .A1(n7790), .A2(n7789), .ZN(n9885) );
  NAND2_X1 U10137 ( .A1(n10168), .A2(n8363), .ZN(n7791) );
  INV_X1 U10138 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10367) );
  OR2_X1 U10139 ( .A1(n8169), .A2(n10367), .ZN(n7796) );
  NAND2_X1 U10140 ( .A1(n7816), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7794) );
  NAND2_X1 U10141 ( .A1(n7815), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7793) );
  NOR2_X1 U10142 ( .A1(n7788), .A2(n7710), .ZN(n7797) );
  MUX2_X1 U10143 ( .A(n7710), .B(n7797), .S(P2_IR_REG_2__SCAN_IN), .Z(n7798)
         );
  INV_X1 U10144 ( .A(n7798), .ZN(n7800) );
  NAND2_X1 U10145 ( .A1(n7800), .A2(n7799), .ZN(n12924) );
  INV_X1 U10146 ( .A(SI_2_), .ZN(n9660) );
  XNOR2_X1 U10147 ( .A(n7801), .B(n9660), .ZN(n7802) );
  XNOR2_X1 U10148 ( .A(n7803), .B(n7802), .ZN(n9648) );
  OR2_X1 U10149 ( .A1(n8162), .A2(n9649), .ZN(n7804) );
  INV_X1 U10150 ( .A(n8419), .ZN(n8427) );
  AND2_X1 U10151 ( .A1(n7807), .A2(n8403), .ZN(n7806) );
  NAND2_X1 U10152 ( .A1(n12916), .A2(n8427), .ZN(n7809) );
  NAND2_X1 U10153 ( .A1(n7809), .A2(n7808), .ZN(n7813) );
  AOI22_X1 U10154 ( .A1(n9755), .A2(n8363), .B1(n10168), .B2(n8427), .ZN(n7810) );
  NAND2_X1 U10155 ( .A1(n7814), .A2(n7813), .ZN(n7832) );
  OR2_X1 U10156 ( .A1(n8169), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7820) );
  NAND2_X1 U10157 ( .A1(n7815), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7819) );
  NAND2_X1 U10158 ( .A1(n6441), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7818) );
  NAND2_X1 U10159 ( .A1(n7816), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7817) );
  NAND4_X1 U10160 ( .A1(n7820), .A2(n7819), .A3(n7818), .A4(n7817), .ZN(n12915) );
  NAND2_X1 U10161 ( .A1(n12915), .A2(n8403), .ZN(n7829) );
  NOR2_X1 U10162 ( .A1(n7703), .A2(n7710), .ZN(n7821) );
  MUX2_X1 U10163 ( .A(n7710), .B(n7821), .S(P2_IR_REG_3__SCAN_IN), .Z(n7823)
         );
  NAND2_X1 U10164 ( .A1(n7825), .A2(n7824), .ZN(n7826) );
  AND2_X1 U10165 ( .A1(n7827), .A2(n7826), .ZN(n9629) );
  NAND2_X1 U10166 ( .A1(n10128), .A2(n8363), .ZN(n7828) );
  NAND2_X1 U10167 ( .A1(n7829), .A2(n7828), .ZN(n7836) );
  INV_X1 U10168 ( .A(n7836), .ZN(n7830) );
  INV_X1 U10169 ( .A(n10128), .ZN(n10431) );
  NAND2_X1 U10170 ( .A1(n12915), .A2(n8363), .ZN(n7831) );
  AND2_X1 U10171 ( .A1(n7832), .A2(n7835), .ZN(n7833) );
  INV_X1 U10172 ( .A(n7835), .ZN(n7837) );
  NAND2_X1 U10173 ( .A1(n6532), .A2(n7838), .ZN(n7839) );
  AND2_X1 U10174 ( .A1(n7840), .A2(n7839), .ZN(n9636) );
  NAND2_X1 U10175 ( .A1(n9636), .A2(n8423), .ZN(n7846) );
  NAND2_X1 U10176 ( .A1(n7841), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7843) );
  MUX2_X1 U10177 ( .A(n7843), .B(P2_IR_REG_31__SCAN_IN), .S(n7842), .Z(n7844)
         );
  NAND2_X1 U10178 ( .A1(n7844), .A2(n7859), .ZN(n9889) );
  INV_X1 U10179 ( .A(n9889), .ZN(n14858) );
  NAND2_X1 U10180 ( .A1(n10240), .A2(n8403), .ZN(n7852) );
  NAND2_X1 U10181 ( .A1(n7816), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7850) );
  OAI21_X1 U10182 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n7865), .ZN(n10379) );
  OR2_X1 U10183 ( .A1(n8169), .A2(n10379), .ZN(n7849) );
  INV_X2 U10184 ( .A(n8429), .ZN(n8396) );
  NAND2_X1 U10185 ( .A1(n8396), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7848) );
  NAND2_X1 U10186 ( .A1(n6442), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7847) );
  NAND4_X1 U10187 ( .A1(n7850), .A2(n7849), .A3(n7848), .A4(n7847), .ZN(n12914) );
  NAND2_X1 U10188 ( .A1(n12914), .A2(n8363), .ZN(n7851) );
  NAND2_X1 U10189 ( .A1(n7852), .A2(n7851), .ZN(n7854) );
  AOI22_X1 U10190 ( .A1(n10240), .A2(n8363), .B1(n12914), .B2(n8427), .ZN(
        n7853) );
  OR2_X1 U10191 ( .A1(n7856), .A2(n7855), .ZN(n7857) );
  AND2_X1 U10192 ( .A1(n7858), .A2(n7857), .ZN(n9641) );
  NAND2_X1 U10193 ( .A1(n9641), .A2(n8423), .ZN(n7863) );
  NAND2_X1 U10194 ( .A1(n7859), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7860) );
  MUX2_X1 U10195 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7860), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n7861) );
  AND2_X1 U10196 ( .A1(n7861), .A2(n7905), .ZN(n12933) );
  AOI22_X1 U10197 ( .A1(n8146), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8145), .B2(
        n12933), .ZN(n7862) );
  NAND2_X1 U10198 ( .A1(n7863), .A2(n7862), .ZN(n10350) );
  NAND2_X1 U10199 ( .A1(n10350), .A2(n8363), .ZN(n7872) );
  NAND2_X1 U10200 ( .A1(n7816), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7870) );
  INV_X1 U10201 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7864) );
  NAND2_X1 U10202 ( .A1(n7865), .A2(n7864), .ZN(n7866) );
  NAND2_X1 U10203 ( .A1(n7891), .A2(n7866), .ZN(n10345) );
  OR2_X1 U10204 ( .A1(n8169), .A2(n10345), .ZN(n7869) );
  NAND2_X1 U10205 ( .A1(n8396), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7868) );
  NAND2_X1 U10206 ( .A1(n6442), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7867) );
  NAND4_X1 U10207 ( .A1(n7870), .A2(n7869), .A3(n7868), .A4(n7867), .ZN(n12913) );
  NAND2_X1 U10208 ( .A1(n12913), .A2(n8403), .ZN(n7871) );
  NAND2_X1 U10209 ( .A1(n7872), .A2(n7871), .ZN(n7878) );
  NAND2_X1 U10210 ( .A1(n10350), .A2(n8403), .ZN(n7874) );
  NAND2_X1 U10211 ( .A1(n12913), .A2(n8363), .ZN(n7873) );
  NAND2_X1 U10212 ( .A1(n7874), .A2(n7873), .ZN(n7875) );
  NAND2_X1 U10213 ( .A1(n7876), .A2(n7875), .ZN(n7882) );
  INV_X1 U10214 ( .A(n7877), .ZN(n7880) );
  INV_X1 U10215 ( .A(n7878), .ZN(n7879) );
  NAND2_X1 U10216 ( .A1(n7880), .A2(n7879), .ZN(n7881) );
  NAND2_X1 U10217 ( .A1(n9665), .A2(n8423), .ZN(n7889) );
  NAND2_X1 U10218 ( .A1(n7905), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7887) );
  XNOR2_X1 U10219 ( .A(n7887), .B(P2_IR_REG_6__SCAN_IN), .ZN(n12945) );
  AOI22_X1 U10220 ( .A1(n8146), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8145), .B2(
        n12945), .ZN(n7888) );
  NAND2_X1 U10221 ( .A1(n15001), .A2(n8403), .ZN(n7898) );
  NAND2_X1 U10222 ( .A1(n8396), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7896) );
  INV_X1 U10223 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7890) );
  NAND2_X1 U10224 ( .A1(n7891), .A2(n7890), .ZN(n7892) );
  NAND2_X1 U10225 ( .A1(n7912), .A2(n7892), .ZN(n10252) );
  OR2_X1 U10226 ( .A1(n8356), .A2(n10252), .ZN(n7895) );
  NAND2_X1 U10227 ( .A1(n7816), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7894) );
  NAND2_X1 U10228 ( .A1(n6441), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7893) );
  NAND4_X1 U10229 ( .A1(n7896), .A2(n7895), .A3(n7894), .A4(n7893), .ZN(n12912) );
  NAND2_X1 U10230 ( .A1(n12912), .A2(n8363), .ZN(n7897) );
  AOI22_X1 U10231 ( .A1(n15001), .A2(n8363), .B1(n12912), .B2(n8427), .ZN(
        n7899) );
  OR2_X1 U10232 ( .A1(n7901), .A2(n7900), .ZN(n7902) );
  OR2_X1 U10233 ( .A1(n9672), .A2(n7904), .ZN(n7910) );
  INV_X1 U10234 ( .A(n7905), .ZN(n7907) );
  INV_X1 U10235 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7906) );
  NAND2_X1 U10236 ( .A1(n7907), .A2(n7906), .ZN(n7927) );
  NAND2_X1 U10237 ( .A1(n7927), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7908) );
  XNOR2_X1 U10238 ( .A(n7908), .B(P2_IR_REG_7__SCAN_IN), .ZN(n12957) );
  AOI22_X1 U10239 ( .A1(n8146), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8145), .B2(
        n12957), .ZN(n7909) );
  NAND2_X1 U10240 ( .A1(n7910), .A2(n7909), .ZN(n10872) );
  NAND2_X1 U10241 ( .A1(n10872), .A2(n8363), .ZN(n7919) );
  NAND2_X1 U10242 ( .A1(n7816), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7917) );
  INV_X1 U10243 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7911) );
  NAND2_X1 U10244 ( .A1(n7912), .A2(n7911), .ZN(n7913) );
  NAND2_X1 U10245 ( .A1(n7932), .A2(n7913), .ZN(n10316) );
  OR2_X1 U10246 ( .A1(n8356), .A2(n10316), .ZN(n7916) );
  NAND2_X1 U10247 ( .A1(n8396), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7915) );
  NAND2_X1 U10248 ( .A1(n6442), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7914) );
  NAND4_X1 U10249 ( .A1(n7917), .A2(n7916), .A3(n7915), .A4(n7914), .ZN(n12911) );
  NAND2_X1 U10250 ( .A1(n12911), .A2(n8403), .ZN(n7918) );
  NAND2_X1 U10251 ( .A1(n10872), .A2(n8403), .ZN(n7921) );
  NAND2_X1 U10252 ( .A1(n12911), .A2(n8363), .ZN(n7920) );
  NAND2_X1 U10253 ( .A1(n7921), .A2(n7920), .ZN(n7922) );
  OR2_X1 U10254 ( .A1(n7924), .A2(n7923), .ZN(n7925) );
  NAND2_X1 U10255 ( .A1(n7926), .A2(n7925), .ZN(n9678) );
  OR2_X1 U10256 ( .A1(n9678), .A2(n7904), .ZN(n7930) );
  NAND2_X1 U10257 ( .A1(n7949), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7928) );
  XNOR2_X1 U10258 ( .A(n7928), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9894) );
  AOI22_X1 U10259 ( .A1(n8146), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8145), .B2(
        n9894), .ZN(n7929) );
  NAND2_X1 U10260 ( .A1(n15018), .A2(n8403), .ZN(n7939) );
  NAND2_X1 U10261 ( .A1(n8385), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7937) );
  INV_X1 U10262 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7931) );
  NAND2_X1 U10263 ( .A1(n7932), .A2(n7931), .ZN(n7933) );
  NAND2_X1 U10264 ( .A1(n7954), .A2(n7933), .ZN(n10923) );
  OR2_X1 U10265 ( .A1(n8356), .A2(n10923), .ZN(n7936) );
  NAND2_X1 U10266 ( .A1(n8396), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7935) );
  NAND2_X1 U10267 ( .A1(n6441), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7934) );
  NAND4_X1 U10268 ( .A1(n7937), .A2(n7936), .A3(n7935), .A4(n7934), .ZN(n12910) );
  NAND2_X1 U10269 ( .A1(n12910), .A2(n8363), .ZN(n7938) );
  NAND2_X1 U10270 ( .A1(n7939), .A2(n7938), .ZN(n7941) );
  AOI22_X1 U10271 ( .A1(n15018), .A2(n8363), .B1(n12910), .B2(n8427), .ZN(
        n7940) );
  OR2_X1 U10272 ( .A1(n7946), .A2(n7945), .ZN(n7947) );
  NAND2_X1 U10273 ( .A1(n7948), .A2(n7947), .ZN(n9683) );
  OR2_X1 U10274 ( .A1(n9683), .A2(n7904), .ZN(n7952) );
  NAND2_X1 U10275 ( .A1(n7971), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7950) );
  XNOR2_X1 U10276 ( .A(n7950), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9896) );
  AOI22_X1 U10277 ( .A1(n8146), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8145), .B2(
        n9896), .ZN(n7951) );
  NAND2_X1 U10278 ( .A1(n11089), .A2(n8363), .ZN(n7961) );
  NAND2_X1 U10279 ( .A1(n8396), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7959) );
  INV_X1 U10280 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7953) );
  NAND2_X1 U10281 ( .A1(n7954), .A2(n7953), .ZN(n7955) );
  NAND2_X1 U10282 ( .A1(n7977), .A2(n7955), .ZN(n10886) );
  OR2_X1 U10283 ( .A1(n8356), .A2(n10886), .ZN(n7958) );
  NAND2_X1 U10284 ( .A1(n8385), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7957) );
  NAND2_X1 U10285 ( .A1(n6441), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7956) );
  NAND4_X1 U10286 ( .A1(n7959), .A2(n7958), .A3(n7957), .A4(n7956), .ZN(n12909) );
  NAND2_X1 U10287 ( .A1(n12909), .A2(n8403), .ZN(n7960) );
  NAND2_X1 U10288 ( .A1(n7961), .A2(n7960), .ZN(n7963) );
  AOI22_X1 U10289 ( .A1(n11089), .A2(n8403), .B1(n8363), .B2(n12909), .ZN(
        n7962) );
  AOI21_X1 U10290 ( .B1(n7964), .B2(n7963), .A(n7962), .ZN(n7966) );
  NOR2_X1 U10291 ( .A1(n7964), .A2(n7963), .ZN(n7965) );
  NAND2_X1 U10292 ( .A1(n7968), .A2(n7967), .ZN(n7969) );
  INV_X1 U10293 ( .A(n7971), .ZN(n7973) );
  INV_X1 U10294 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7972) );
  NAND2_X1 U10295 ( .A1(n7973), .A2(n7972), .ZN(n7990) );
  NAND2_X1 U10296 ( .A1(n7990), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7974) );
  XNOR2_X1 U10297 ( .A(n7974), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11292) );
  AOI22_X1 U10298 ( .A1(n8146), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n11292), 
        .B2(n8145), .ZN(n7975) );
  NAND2_X1 U10299 ( .A1(n15027), .A2(n8403), .ZN(n7984) );
  NAND2_X1 U10300 ( .A1(n8385), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7982) );
  NAND2_X1 U10301 ( .A1(n7977), .A2(n7976), .ZN(n7978) );
  NAND2_X1 U10302 ( .A1(n7995), .A2(n7978), .ZN(n10930) );
  OR2_X1 U10303 ( .A1(n8356), .A2(n10930), .ZN(n7981) );
  NAND2_X1 U10304 ( .A1(n8396), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7980) );
  NAND2_X1 U10305 ( .A1(n6442), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7979) );
  NAND4_X1 U10306 ( .A1(n7982), .A2(n7981), .A3(n7980), .A4(n7979), .ZN(n12908) );
  NAND2_X1 U10307 ( .A1(n12908), .A2(n8363), .ZN(n7983) );
  NAND2_X1 U10308 ( .A1(n15027), .A2(n8363), .ZN(n7986) );
  NAND2_X1 U10309 ( .A1(n12908), .A2(n8403), .ZN(n7985) );
  NAND2_X1 U10310 ( .A1(n7986), .A2(n7985), .ZN(n7987) );
  XNOR2_X1 U10311 ( .A(n7989), .B(n7988), .ZN(n9929) );
  NAND2_X1 U10312 ( .A1(n9929), .A2(n8423), .ZN(n7993) );
  OAI21_X1 U10313 ( .B1(n7990), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7991) );
  XNOR2_X1 U10314 ( .A(n7991), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11295) );
  AOI22_X1 U10315 ( .A1(n11295), .A2(n8145), .B1(n8146), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n7992) );
  NAND2_X1 U10316 ( .A1(n11376), .A2(n8363), .ZN(n8002) );
  NAND2_X1 U10317 ( .A1(n8385), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8000) );
  INV_X1 U10318 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7994) );
  NAND2_X1 U10319 ( .A1(n7995), .A2(n7994), .ZN(n7996) );
  NAND2_X1 U10320 ( .A1(n8015), .A2(n7996), .ZN(n11203) );
  OR2_X1 U10321 ( .A1(n8356), .A2(n11203), .ZN(n7999) );
  NAND2_X1 U10322 ( .A1(n8396), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7998) );
  NAND2_X1 U10323 ( .A1(n6441), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7997) );
  NAND4_X1 U10324 ( .A1(n8000), .A2(n7999), .A3(n7998), .A4(n7997), .ZN(n12907) );
  NAND2_X1 U10325 ( .A1(n12907), .A2(n8403), .ZN(n8001) );
  NAND2_X1 U10326 ( .A1(n8002), .A2(n8001), .ZN(n8004) );
  AOI22_X1 U10327 ( .A1(n11376), .A2(n8403), .B1(n8363), .B2(n12907), .ZN(
        n8003) );
  XNOR2_X1 U10328 ( .A(n8005), .B(n8006), .ZN(n9999) );
  NAND2_X1 U10329 ( .A1(n9999), .A2(n8423), .ZN(n8013) );
  CLKBUF_X1 U10330 ( .A(n8007), .Z(n8008) );
  INV_X1 U10331 ( .A(n8008), .ZN(n8009) );
  NAND2_X1 U10332 ( .A1(n8009), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8010) );
  MUX2_X1 U10333 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8010), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8011) );
  AND2_X1 U10334 ( .A1(n8011), .A2(n7716), .ZN(n11297) );
  AOI22_X1 U10335 ( .A1(n8146), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8145), 
        .B2(n11297), .ZN(n8012) );
  NAND2_X2 U10336 ( .A1(n8013), .A2(n8012), .ZN(n11361) );
  NAND2_X1 U10337 ( .A1(n11361), .A2(n8403), .ZN(n8022) );
  NAND2_X1 U10338 ( .A1(n8015), .A2(n8014), .ZN(n8016) );
  NAND2_X1 U10339 ( .A1(n8032), .A2(n8016), .ZN(n11224) );
  OR2_X1 U10340 ( .A1(n8356), .A2(n11224), .ZN(n8020) );
  NAND2_X1 U10341 ( .A1(n8396), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8019) );
  NAND2_X1 U10342 ( .A1(n6442), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8018) );
  NAND2_X1 U10343 ( .A1(n8385), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8017) );
  NAND4_X1 U10344 ( .A1(n8020), .A2(n8019), .A3(n8018), .A4(n8017), .ZN(n12906) );
  NAND2_X1 U10345 ( .A1(n12906), .A2(n8363), .ZN(n8021) );
  NAND2_X1 U10346 ( .A1(n11361), .A2(n8363), .ZN(n8024) );
  NAND2_X1 U10347 ( .A1(n12906), .A2(n8403), .ZN(n8023) );
  NAND2_X1 U10348 ( .A1(n8024), .A2(n8023), .ZN(n8025) );
  XNOR2_X1 U10349 ( .A(n8026), .B(n8027), .ZN(n10076) );
  NAND2_X1 U10350 ( .A1(n10076), .A2(n8423), .ZN(n8030) );
  NAND2_X1 U10351 ( .A1(n7716), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8028) );
  XNOR2_X1 U10352 ( .A(n8028), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11300) );
  AOI22_X1 U10353 ( .A1(n8146), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8145), 
        .B2(n11300), .ZN(n8029) );
  NAND2_X1 U10354 ( .A1(n11704), .A2(n8363), .ZN(n8039) );
  NAND2_X1 U10355 ( .A1(n7815), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8037) );
  INV_X1 U10356 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8031) );
  NAND2_X1 U10357 ( .A1(n8032), .A2(n8031), .ZN(n8033) );
  NAND2_X1 U10358 ( .A1(n8055), .A2(n8033), .ZN(n11184) );
  OR2_X1 U10359 ( .A1(n8169), .A2(n11184), .ZN(n8036) );
  NAND2_X1 U10360 ( .A1(n8385), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8035) );
  NAND2_X1 U10361 ( .A1(n6442), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8034) );
  NAND4_X1 U10362 ( .A1(n8037), .A2(n8036), .A3(n8035), .A4(n8034), .ZN(n13226) );
  NAND2_X1 U10363 ( .A1(n13226), .A2(n8403), .ZN(n8038) );
  NAND2_X1 U10364 ( .A1(n8039), .A2(n8038), .ZN(n8042) );
  AOI22_X1 U10365 ( .A1(n11704), .A2(n8403), .B1(n8363), .B2(n13226), .ZN(
        n8040) );
  AOI21_X1 U10366 ( .B1(n8043), .B2(n8042), .A(n8040), .ZN(n8041) );
  INV_X1 U10367 ( .A(n8041), .ZN(n8044) );
  NAND2_X1 U10368 ( .A1(n8046), .A2(n8045), .ZN(n8047) );
  AND2_X1 U10369 ( .A1(n8048), .A2(n8047), .ZN(n10389) );
  NAND2_X1 U10370 ( .A1(n10389), .A2(n8423), .ZN(n8053) );
  INV_X1 U10371 ( .A(n8049), .ZN(n8050) );
  NAND2_X1 U10372 ( .A1(n8050), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8051) );
  XNOR2_X1 U10373 ( .A(n8051), .B(P2_IR_REG_14__SCAN_IN), .ZN(n14944) );
  AOI22_X1 U10374 ( .A1(n8146), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8145), 
        .B2(n14944), .ZN(n8052) );
  NAND2_X1 U10375 ( .A1(n13323), .A2(n8403), .ZN(n8062) );
  NAND2_X1 U10376 ( .A1(n7815), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8060) );
  NAND2_X1 U10377 ( .A1(n8055), .A2(n8054), .ZN(n8056) );
  NAND2_X1 U10378 ( .A1(n8077), .A2(n8056), .ZN(n13218) );
  OR2_X1 U10379 ( .A1(n8356), .A2(n13218), .ZN(n8059) );
  NAND2_X1 U10380 ( .A1(n6442), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8058) );
  NAND2_X1 U10381 ( .A1(n8385), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8057) );
  NAND4_X1 U10382 ( .A1(n8060), .A2(n8059), .A3(n8058), .A4(n8057), .ZN(n13203) );
  NAND2_X1 U10383 ( .A1(n13203), .A2(n8363), .ZN(n8061) );
  NAND2_X1 U10384 ( .A1(n8062), .A2(n8061), .ZN(n8067) );
  NAND2_X1 U10385 ( .A1(n13323), .A2(n8363), .ZN(n8064) );
  NAND2_X1 U10386 ( .A1(n13203), .A2(n8403), .ZN(n8063) );
  NAND2_X1 U10387 ( .A1(n8064), .A2(n8063), .ZN(n8065) );
  INV_X1 U10388 ( .A(n8067), .ZN(n8068) );
  XNOR2_X1 U10389 ( .A(n8070), .B(n8069), .ZN(n10753) );
  NAND2_X1 U10390 ( .A1(n10753), .A2(n8423), .ZN(n8075) );
  NAND2_X1 U10391 ( .A1(n8071), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8073) );
  INV_X1 U10392 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8072) );
  XNOR2_X1 U10393 ( .A(n8073), .B(n8072), .ZN(n11306) );
  INV_X1 U10394 ( .A(n11306), .ZN(n14956) );
  AOI22_X1 U10395 ( .A1(n8146), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8145), 
        .B2(n14956), .ZN(n8074) );
  NAND2_X1 U10396 ( .A1(n13318), .A2(n8363), .ZN(n8084) );
  NAND2_X1 U10397 ( .A1(n8077), .A2(n8076), .ZN(n8078) );
  AND2_X1 U10398 ( .A1(n8096), .A2(n8078), .ZN(n13208) );
  NAND2_X1 U10399 ( .A1(n13208), .A2(n8328), .ZN(n8082) );
  INV_X1 U10400 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14952) );
  OR2_X1 U10401 ( .A1(n8429), .A2(n14952), .ZN(n8081) );
  NAND2_X1 U10402 ( .A1(n8385), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8080) );
  NAND2_X1 U10403 ( .A1(n6442), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n8079) );
  NAND4_X1 U10404 ( .A1(n8082), .A2(n8081), .A3(n8080), .A4(n8079), .ZN(n13224) );
  NAND2_X1 U10405 ( .A1(n13224), .A2(n8403), .ZN(n8083) );
  AOI22_X1 U10406 ( .A1(n13318), .A2(n8403), .B1(n8363), .B2(n13224), .ZN(
        n8085) );
  XNOR2_X1 U10407 ( .A(n8087), .B(n8086), .ZN(n10802) );
  NAND2_X1 U10408 ( .A1(n10802), .A2(n8423), .ZN(n8093) );
  NAND2_X1 U10409 ( .A1(n8088), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8089) );
  MUX2_X1 U10410 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8089), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n8091) );
  NAND2_X1 U10411 ( .A1(n8091), .A2(n8090), .ZN(n11309) );
  INV_X1 U10412 ( .A(n11309), .ZN(n14970) );
  AOI22_X1 U10413 ( .A1(n8146), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8145), 
        .B2(n14970), .ZN(n8092) );
  NAND2_X1 U10414 ( .A1(n13189), .A2(n8403), .ZN(n8101) );
  INV_X1 U10415 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8099) );
  NAND2_X1 U10416 ( .A1(n7815), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8095) );
  NAND2_X1 U10417 ( .A1(n8385), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8094) );
  AND2_X1 U10418 ( .A1(n8095), .A2(n8094), .ZN(n8098) );
  XNOR2_X1 U10419 ( .A(n8096), .B(P2_REG3_REG_16__SCAN_IN), .ZN(n13192) );
  NAND2_X1 U10420 ( .A1(n13192), .A2(n8328), .ZN(n8097) );
  OAI211_X1 U10421 ( .C1(n8432), .C2(n8099), .A(n8098), .B(n8097), .ZN(n13204)
         );
  NAND2_X1 U10422 ( .A1(n13204), .A2(n8363), .ZN(n8100) );
  NAND2_X1 U10423 ( .A1(n8101), .A2(n8100), .ZN(n8103) );
  AOI22_X1 U10424 ( .A1(n13189), .A2(n8363), .B1(n13204), .B2(n8427), .ZN(
        n8102) );
  AOI21_X1 U10425 ( .B1(n8104), .B2(n8103), .A(n8102), .ZN(n8106) );
  NOR2_X1 U10426 ( .A1(n8104), .A2(n8103), .ZN(n8105) );
  OR2_X1 U10427 ( .A1(n8106), .A2(n8105), .ZN(n8111) );
  NAND2_X1 U10428 ( .A1(n8111), .A2(n8112), .ZN(n8110) );
  NAND2_X1 U10429 ( .A1(n13307), .A2(n8403), .ZN(n8108) );
  NAND2_X1 U10430 ( .A1(n13186), .A2(n8363), .ZN(n8107) );
  NAND2_X1 U10431 ( .A1(n8108), .A2(n8107), .ZN(n8109) );
  NAND2_X1 U10432 ( .A1(n8116), .A2(SI_17_), .ZN(n8133) );
  NAND2_X1 U10433 ( .A1(n8137), .A2(n8133), .ZN(n8118) );
  MUX2_X1 U10434 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9619), .Z(n8136) );
  XNOR2_X1 U10435 ( .A(n8136), .B(SI_18_), .ZN(n8117) );
  NAND2_X1 U10436 ( .A1(n11033), .A2(n8423), .ZN(n8121) );
  NAND2_X1 U10437 ( .A1(n8493), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8119) );
  XNOR2_X1 U10438 ( .A(n8119), .B(P2_IR_REG_18__SCAN_IN), .ZN(n12969) );
  AOI22_X1 U10439 ( .A1(n8146), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8145), 
        .B2(n12969), .ZN(n8120) );
  NAND2_X1 U10440 ( .A1(n13302), .A2(n8403), .ZN(n8130) );
  INV_X1 U10441 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8128) );
  INV_X1 U10442 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8123) );
  NAND2_X1 U10443 ( .A1(n8124), .A2(n8123), .ZN(n8125) );
  NAND2_X1 U10444 ( .A1(n8150), .A2(n8125), .ZN(n13160) );
  OR2_X1 U10445 ( .A1(n13160), .A2(n8356), .ZN(n8127) );
  AOI22_X1 U10446 ( .A1(n8385), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n7815), .B2(
        P2_REG1_REG_18__SCAN_IN), .ZN(n8126) );
  OAI211_X1 U10447 ( .C1(n8432), .C2(n8128), .A(n8127), .B(n8126), .ZN(n13165)
         );
  NAND2_X1 U10448 ( .A1(n13165), .A2(n8363), .ZN(n8129) );
  NAND2_X1 U10449 ( .A1(n8130), .A2(n8129), .ZN(n8132) );
  AOI22_X1 U10450 ( .A1(n13302), .A2(n8363), .B1(n13165), .B2(n8427), .ZN(
        n8131) );
  INV_X1 U10451 ( .A(n8136), .ZN(n8134) );
  INV_X1 U10452 ( .A(SI_18_), .ZN(n9941) );
  OAI21_X1 U10453 ( .B1(n8134), .B2(n9941), .A(n8133), .ZN(n8135) );
  INV_X1 U10454 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11127) );
  MUX2_X1 U10455 ( .A(n11125), .B(n11127), .S(n9619), .Z(n8138) );
  INV_X1 U10456 ( .A(SI_19_), .ZN(n9942) );
  NAND2_X1 U10457 ( .A1(n8138), .A2(n9942), .ZN(n8160) );
  INV_X1 U10458 ( .A(n8138), .ZN(n8139) );
  NAND2_X1 U10459 ( .A1(n8139), .A2(SI_19_), .ZN(n8140) );
  NAND2_X1 U10460 ( .A1(n8160), .A2(n8140), .ZN(n8142) );
  NAND2_X1 U10461 ( .A1(n8141), .A2(n8142), .ZN(n8144) );
  NAND2_X1 U10462 ( .A1(n8144), .A2(n8161), .ZN(n11124) );
  NAND2_X1 U10463 ( .A1(n11124), .A2(n8423), .ZN(n8148) );
  AOI22_X1 U10464 ( .A1(n8146), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8145), 
        .B2(n6914), .ZN(n8147) );
  NAND2_X1 U10465 ( .A1(n13298), .A2(n8363), .ZN(n8155) );
  INV_X1 U10466 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8149) );
  NAND2_X1 U10467 ( .A1(n8150), .A2(n8149), .ZN(n8151) );
  NAND2_X1 U10468 ( .A1(n8167), .A2(n8151), .ZN(n13144) );
  AOI22_X1 U10469 ( .A1(n6441), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n8396), .B2(
        P2_REG1_REG_19__SCAN_IN), .ZN(n8153) );
  NAND2_X1 U10470 ( .A1(n8385), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8152) );
  OAI211_X1 U10471 ( .C1(n13144), .C2(n8356), .A(n8153), .B(n8152), .ZN(n13126) );
  NAND2_X1 U10472 ( .A1(n13126), .A2(n8403), .ZN(n8154) );
  NAND2_X1 U10473 ( .A1(n8155), .A2(n8154), .ZN(n8159) );
  NAND2_X1 U10474 ( .A1(n13298), .A2(n8403), .ZN(n8157) );
  NAND2_X1 U10475 ( .A1(n13126), .A2(n8363), .ZN(n8156) );
  INV_X1 U10476 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11375) );
  MUX2_X1 U10477 ( .A(n11375), .B(n11373), .S(n7171), .Z(n8183) );
  NAND2_X1 U10478 ( .A1(n11371), .A2(n8423), .ZN(n8164) );
  OR2_X1 U10479 ( .A1(n8162), .A2(n11373), .ZN(n8163) );
  NAND2_X1 U10480 ( .A1(n13290), .A2(n8403), .ZN(n8177) );
  INV_X1 U10481 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8166) );
  NAND2_X1 U10482 ( .A1(n8167), .A2(n8166), .ZN(n8168) );
  NAND2_X1 U10483 ( .A1(n8191), .A2(n8168), .ZN(n12846) );
  OR2_X1 U10484 ( .A1(n12846), .A2(n8169), .ZN(n8175) );
  INV_X1 U10485 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8172) );
  NAND2_X1 U10486 ( .A1(n8385), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8171) );
  NAND2_X1 U10487 ( .A1(n7815), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8170) );
  OAI211_X1 U10488 ( .C1(n8172), .C2(n8432), .A(n8171), .B(n8170), .ZN(n8173)
         );
  INV_X1 U10489 ( .A(n8173), .ZN(n8174) );
  NAND2_X1 U10490 ( .A1(n8175), .A2(n8174), .ZN(n13106) );
  NAND2_X1 U10491 ( .A1(n13106), .A2(n8363), .ZN(n8176) );
  NAND2_X1 U10492 ( .A1(n8177), .A2(n8176), .ZN(n8180) );
  AOI22_X1 U10493 ( .A1(n13290), .A2(n8363), .B1(n13106), .B2(n8403), .ZN(
        n8178) );
  INV_X1 U10494 ( .A(n8179), .ZN(n8182) );
  NAND2_X1 U10495 ( .A1(n8182), .A2(n7647), .ZN(n8203) );
  INV_X1 U10496 ( .A(n8183), .ZN(n8184) );
  INV_X1 U10497 ( .A(SI_20_), .ZN(n10182) );
  MUX2_X1 U10498 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n7171), .Z(n8209) );
  XNOR2_X1 U10499 ( .A(n8209), .B(SI_21_), .ZN(n8206) );
  XNOR2_X1 U10500 ( .A(n8208), .B(n8206), .ZN(n11444) );
  NAND2_X1 U10501 ( .A1(n11444), .A2(n8423), .ZN(n8189) );
  INV_X1 U10502 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11446) );
  OR2_X1 U10503 ( .A1(n8162), .A2(n11446), .ZN(n8188) );
  NAND2_X1 U10504 ( .A1(n13286), .A2(n8363), .ZN(n8200) );
  INV_X1 U10505 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8190) );
  NAND2_X1 U10506 ( .A1(n8191), .A2(n8190), .ZN(n8192) );
  AND2_X1 U10507 ( .A1(n8215), .A2(n8192), .ZN(n13109) );
  NAND2_X1 U10508 ( .A1(n13109), .A2(n8328), .ZN(n8198) );
  INV_X1 U10509 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8195) );
  NAND2_X1 U10510 ( .A1(n8396), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8194) );
  NAND2_X1 U10511 ( .A1(n8385), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8193) );
  OAI211_X1 U10512 ( .C1(n8195), .C2(n8432), .A(n8194), .B(n8193), .ZN(n8196)
         );
  INV_X1 U10513 ( .A(n8196), .ZN(n8197) );
  NAND2_X1 U10514 ( .A1(n8198), .A2(n8197), .ZN(n13127) );
  NAND2_X1 U10515 ( .A1(n13127), .A2(n8403), .ZN(n8199) );
  NAND2_X1 U10516 ( .A1(n8200), .A2(n8199), .ZN(n8204) );
  INV_X1 U10517 ( .A(n13127), .ZN(n12865) );
  NAND2_X1 U10518 ( .A1(n13286), .A2(n8403), .ZN(n8201) );
  OAI21_X1 U10519 ( .B1(n12865), .B2(n8245), .A(n8201), .ZN(n8202) );
  NAND2_X1 U10520 ( .A1(n8209), .A2(SI_21_), .ZN(n8210) );
  MUX2_X1 U10521 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n7171), .Z(n8251) );
  XNOR2_X1 U10522 ( .A(n9428), .B(n8251), .ZN(n11617) );
  NAND2_X1 U10523 ( .A1(n11617), .A2(n8423), .ZN(n8212) );
  INV_X1 U10524 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n15239) );
  OR2_X1 U10525 ( .A1(n8162), .A2(n15239), .ZN(n8211) );
  NAND2_X1 U10526 ( .A1(n13280), .A2(n8403), .ZN(n8223) );
  INV_X1 U10527 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8214) );
  NAND2_X1 U10528 ( .A1(n8215), .A2(n8214), .ZN(n8216) );
  NAND2_X1 U10529 ( .A1(n8235), .A2(n8216), .ZN(n13095) );
  INV_X1 U10530 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n15302) );
  NAND2_X1 U10531 ( .A1(n7815), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8218) );
  NAND2_X1 U10532 ( .A1(n8385), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8217) );
  OAI211_X1 U10533 ( .C1(n15302), .C2(n8432), .A(n8218), .B(n8217), .ZN(n8219)
         );
  INV_X1 U10534 ( .A(n8219), .ZN(n8220) );
  NAND2_X1 U10535 ( .A1(n13105), .A2(n8363), .ZN(n8222) );
  NAND2_X1 U10536 ( .A1(n8223), .A2(n8222), .ZN(n8225) );
  AOI22_X1 U10537 ( .A1(n13280), .A2(n8363), .B1(n13105), .B2(n8403), .ZN(
        n8224) );
  INV_X1 U10538 ( .A(n9428), .ZN(n8227) );
  NAND2_X1 U10539 ( .A1(n8227), .A2(n8251), .ZN(n8229) );
  NAND2_X1 U10540 ( .A1(n8250), .A2(SI_22_), .ZN(n8228) );
  NAND2_X1 U10541 ( .A1(n8229), .A2(n8228), .ZN(n8231) );
  MUX2_X1 U10542 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n7171), .Z(n8254) );
  XNOR2_X1 U10543 ( .A(n8254), .B(SI_23_), .ZN(n8230) );
  NAND2_X1 U10544 ( .A1(n14315), .A2(n8423), .ZN(n8233) );
  INV_X1 U10545 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n13373) );
  OR2_X1 U10546 ( .A1(n8162), .A2(n13373), .ZN(n8232) );
  NAND2_X1 U10547 ( .A1(n13275), .A2(n8363), .ZN(n8243) );
  INV_X1 U10548 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8234) );
  NAND2_X1 U10549 ( .A1(n8235), .A2(n8234), .ZN(n8236) );
  AND2_X1 U10550 ( .A1(n8260), .A2(n8236), .ZN(n13078) );
  NAND2_X1 U10551 ( .A1(n13078), .A2(n8328), .ZN(n8241) );
  INV_X1 U10552 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n15260) );
  NAND2_X1 U10553 ( .A1(n8396), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8238) );
  NAND2_X1 U10554 ( .A1(n8385), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8237) );
  OAI211_X1 U10555 ( .C1(n8432), .C2(n15260), .A(n8238), .B(n8237), .ZN(n8239)
         );
  INV_X1 U10556 ( .A(n8239), .ZN(n8240) );
  NAND2_X1 U10557 ( .A1(n8241), .A2(n8240), .ZN(n13087) );
  NAND2_X1 U10558 ( .A1(n13087), .A2(n8427), .ZN(n8242) );
  INV_X1 U10559 ( .A(n13087), .ZN(n12866) );
  NAND2_X1 U10560 ( .A1(n13275), .A2(n8403), .ZN(n8244) );
  OAI21_X1 U10561 ( .B1(n12866), .B2(n8245), .A(n8244), .ZN(n8246) );
  INV_X1 U10562 ( .A(n8254), .ZN(n8247) );
  INV_X1 U10563 ( .A(SI_23_), .ZN(n10773) );
  NAND2_X1 U10564 ( .A1(n8247), .A2(n10773), .ZN(n8255) );
  OAI21_X1 U10565 ( .B1(SI_22_), .B2(n8251), .A(n8255), .ZN(n8248) );
  INV_X1 U10566 ( .A(n8248), .ZN(n8249) );
  INV_X1 U10567 ( .A(n8251), .ZN(n8253) );
  INV_X1 U10568 ( .A(SI_22_), .ZN(n8252) );
  NOR2_X1 U10569 ( .A1(n8253), .A2(n8252), .ZN(n8256) );
  AOI22_X1 U10570 ( .A1(n8256), .A2(n8255), .B1(n8254), .B2(SI_23_), .ZN(n8257) );
  MUX2_X1 U10571 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9619), .Z(n8273) );
  XNOR2_X1 U10572 ( .A(n8275), .B(n8273), .ZN(n11545) );
  NAND2_X1 U10573 ( .A1(n11545), .A2(n8423), .ZN(n8259) );
  INV_X1 U10574 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13368) );
  OR2_X1 U10575 ( .A1(n8162), .A2(n13368), .ZN(n8258) );
  NAND2_X1 U10576 ( .A1(n13269), .A2(n8403), .ZN(n8267) );
  INV_X1 U10577 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n15315) );
  NAND2_X1 U10578 ( .A1(n8260), .A2(n15315), .ZN(n8261) );
  NAND2_X1 U10579 ( .A1(n8300), .A2(n8261), .ZN(n13065) );
  INV_X1 U10580 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n15245) );
  NAND2_X1 U10581 ( .A1(n7815), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U10582 ( .A1(n8385), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8262) );
  OAI211_X1 U10583 ( .C1(n8432), .C2(n15245), .A(n8263), .B(n8262), .ZN(n8264)
         );
  INV_X1 U10584 ( .A(n8264), .ZN(n8265) );
  NAND2_X1 U10585 ( .A1(n13074), .A2(n8363), .ZN(n8266) );
  NAND2_X1 U10586 ( .A1(n8267), .A2(n8266), .ZN(n8269) );
  AOI22_X1 U10587 ( .A1(n13269), .A2(n8363), .B1(n13074), .B2(n8403), .ZN(
        n8268) );
  AOI21_X1 U10588 ( .B1(n8270), .B2(n8269), .A(n8268), .ZN(n8272) );
  INV_X1 U10589 ( .A(n8273), .ZN(n8274) );
  NAND2_X1 U10590 ( .A1(n8276), .A2(SI_24_), .ZN(n8277) );
  INV_X1 U10591 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14313) );
  INV_X1 U10592 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13364) );
  MUX2_X1 U10593 ( .A(n14313), .B(n13364), .S(n7171), .Z(n8278) );
  INV_X1 U10594 ( .A(SI_25_), .ZN(n11003) );
  NAND2_X1 U10595 ( .A1(n8278), .A2(n11003), .ZN(n8281) );
  INV_X1 U10596 ( .A(n8278), .ZN(n8279) );
  NAND2_X1 U10597 ( .A1(n8279), .A2(SI_25_), .ZN(n8280) );
  NAND2_X1 U10598 ( .A1(n8281), .A2(n8280), .ZN(n8296) );
  INV_X1 U10599 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14307) );
  INV_X1 U10600 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13360) );
  MUX2_X1 U10601 ( .A(n14307), .B(n13360), .S(n7171), .Z(n8311) );
  XNOR2_X1 U10602 ( .A(n8311), .B(SI_26_), .ZN(n8282) );
  XNOR2_X1 U10603 ( .A(n8312), .B(n8282), .ZN(n13359) );
  NAND2_X1 U10604 ( .A1(n13359), .A2(n8423), .ZN(n8284) );
  OR2_X1 U10605 ( .A1(n8162), .A2(n13360), .ZN(n8283) );
  NAND2_X1 U10606 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n8285) );
  INV_X1 U10607 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n12816) );
  INV_X1 U10608 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8286) );
  OAI21_X1 U10609 ( .B1(n8300), .B2(n12816), .A(n8286), .ZN(n8287) );
  NAND2_X1 U10610 ( .A1(n13031), .A2(n8328), .ZN(n8292) );
  INV_X1 U10611 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n15257) );
  NAND2_X1 U10612 ( .A1(n8385), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8289) );
  NAND2_X1 U10613 ( .A1(n7815), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8288) );
  OAI211_X1 U10614 ( .C1(n15257), .C2(n8432), .A(n8289), .B(n8288), .ZN(n8290)
         );
  INV_X1 U10615 ( .A(n8290), .ZN(n8291) );
  AND2_X1 U10616 ( .A1(n13012), .A2(n8427), .ZN(n8293) );
  AOI21_X1 U10617 ( .B1(n13259), .B2(n8363), .A(n8293), .ZN(n8341) );
  NAND2_X1 U10618 ( .A1(n13259), .A2(n8403), .ZN(n8295) );
  NAND2_X1 U10619 ( .A1(n13012), .A2(n8363), .ZN(n8294) );
  NAND2_X1 U10620 ( .A1(n8295), .A2(n8294), .ZN(n8340) );
  NAND2_X1 U10621 ( .A1(n8341), .A2(n8340), .ZN(n8345) );
  INV_X1 U10622 ( .A(n8345), .ZN(n8310) );
  XNOR2_X1 U10623 ( .A(n8297), .B(n8296), .ZN(n13362) );
  NAND2_X1 U10624 ( .A1(n13362), .A2(n8423), .ZN(n8299) );
  OR2_X1 U10625 ( .A1(n8162), .A2(n13364), .ZN(n8298) );
  NAND2_X1 U10626 ( .A1(n13266), .A2(n8363), .ZN(n8307) );
  XNOR2_X1 U10627 ( .A(n8300), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n13047) );
  NAND2_X1 U10628 ( .A1(n13047), .A2(n8328), .ZN(n8305) );
  INV_X1 U10629 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n15332) );
  NAND2_X1 U10630 ( .A1(n8385), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8302) );
  NAND2_X1 U10631 ( .A1(n8396), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8301) );
  OAI211_X1 U10632 ( .C1(n15332), .C2(n8432), .A(n8302), .B(n8301), .ZN(n8303)
         );
  INV_X1 U10633 ( .A(n8303), .ZN(n8304) );
  NAND2_X1 U10634 ( .A1(n13060), .A2(n8403), .ZN(n8306) );
  NAND2_X1 U10635 ( .A1(n8307), .A2(n8306), .ZN(n8338) );
  AND2_X1 U10636 ( .A1(n13060), .A2(n8363), .ZN(n8308) );
  AOI21_X1 U10637 ( .B1(n13266), .B2(n8427), .A(n8308), .ZN(n8339) );
  NOR2_X1 U10638 ( .A1(n8338), .A2(n8339), .ZN(n8309) );
  MUX2_X1 U10639 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n7171), .Z(n8346) );
  NAND2_X1 U10640 ( .A1(n8346), .A2(SI_27_), .ZN(n8313) );
  NAND2_X1 U10641 ( .A1(n8314), .A2(n8313), .ZN(n8321) );
  INV_X1 U10642 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11549) );
  INV_X1 U10643 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9003) );
  MUX2_X1 U10644 ( .A(n11549), .B(n9003), .S(n9619), .Z(n8315) );
  INV_X1 U10645 ( .A(SI_28_), .ZN(n11512) );
  NAND2_X1 U10646 ( .A1(n8315), .A2(n11512), .ZN(n8372) );
  INV_X1 U10647 ( .A(n8315), .ZN(n8316) );
  NAND2_X1 U10648 ( .A1(n8316), .A2(SI_28_), .ZN(n8317) );
  NAND2_X1 U10649 ( .A1(n8372), .A2(n8317), .ZN(n8320) );
  NAND2_X1 U10650 ( .A1(n8321), .A2(n8320), .ZN(n8322) );
  NAND2_X1 U10651 ( .A1(n8373), .A2(n8322), .ZN(n11548) );
  NAND2_X1 U10652 ( .A1(n11548), .A2(n8423), .ZN(n8324) );
  OR2_X1 U10653 ( .A1(n8162), .A2(n9003), .ZN(n8323) );
  INV_X1 U10654 ( .A(n8353), .ZN(n8325) );
  NAND2_X1 U10655 ( .A1(n8325), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8355) );
  INV_X1 U10656 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8326) );
  NAND2_X1 U10657 ( .A1(n8355), .A2(n8326), .ZN(n8327) );
  NAND2_X1 U10658 ( .A1(n13006), .A2(n8328), .ZN(n8334) );
  INV_X1 U10659 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8331) );
  NAND2_X1 U10660 ( .A1(n7815), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8330) );
  NAND2_X1 U10661 ( .A1(n8385), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8329) );
  OAI211_X1 U10662 ( .C1(n8331), .C2(n8432), .A(n8330), .B(n8329), .ZN(n8332)
         );
  INV_X1 U10663 ( .A(n8332), .ZN(n8333) );
  AND2_X1 U10664 ( .A1(n13011), .A2(n8363), .ZN(n8335) );
  AOI21_X1 U10665 ( .B1(n13250), .B2(n8403), .A(n8335), .ZN(n8411) );
  NAND2_X1 U10666 ( .A1(n13250), .A2(n8363), .ZN(n8337) );
  NAND2_X1 U10667 ( .A1(n13011), .A2(n8403), .ZN(n8336) );
  NAND2_X1 U10668 ( .A1(n8337), .A2(n8336), .ZN(n8410) );
  NAND2_X1 U10669 ( .A1(n8411), .A2(n8410), .ZN(n8415) );
  AND2_X1 U10670 ( .A1(n8339), .A2(n8338), .ZN(n8344) );
  INV_X1 U10671 ( .A(n8340), .ZN(n8343) );
  INV_X1 U10672 ( .A(n8341), .ZN(n8342) );
  AOI22_X1 U10673 ( .A1(n8345), .A2(n8344), .B1(n8343), .B2(n8342), .ZN(n8368)
         );
  INV_X1 U10674 ( .A(n8346), .ZN(n8347) );
  XNOR2_X1 U10675 ( .A(n8347), .B(SI_27_), .ZN(n8348) );
  OR2_X1 U10676 ( .A1(n8162), .A2(n13358), .ZN(n8350) );
  INV_X1 U10677 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8352) );
  NAND2_X1 U10678 ( .A1(n8353), .A2(n8352), .ZN(n8354) );
  NAND2_X1 U10679 ( .A1(n8355), .A2(n8354), .ZN(n12780) );
  OR2_X1 U10680 ( .A1(n12780), .A2(n8356), .ZN(n8362) );
  INV_X1 U10681 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8359) );
  NAND2_X1 U10682 ( .A1(n8385), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8358) );
  NAND2_X1 U10683 ( .A1(n8396), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8357) );
  OAI211_X1 U10684 ( .C1(n8359), .C2(n8432), .A(n8358), .B(n8357), .ZN(n8360)
         );
  INV_X1 U10685 ( .A(n8360), .ZN(n8361) );
  AND2_X1 U10686 ( .A1(n13027), .A2(n8363), .ZN(n8364) );
  AOI21_X1 U10687 ( .B1(n13255), .B2(n8403), .A(n8364), .ZN(n8407) );
  NAND2_X1 U10688 ( .A1(n13255), .A2(n8363), .ZN(n8366) );
  NAND2_X1 U10689 ( .A1(n13027), .A2(n8403), .ZN(n8365) );
  NAND2_X1 U10690 ( .A1(n8366), .A2(n8365), .ZN(n8406) );
  NAND2_X1 U10691 ( .A1(n8407), .A2(n8406), .ZN(n8367) );
  INV_X1 U10692 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14304) );
  INV_X1 U10693 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13350) );
  MUX2_X1 U10694 ( .A(n14304), .B(n13350), .S(n9619), .Z(n8374) );
  INV_X1 U10695 ( .A(SI_29_), .ZN(n11515) );
  NAND2_X1 U10696 ( .A1(n8374), .A2(n11515), .ZN(n8377) );
  INV_X1 U10697 ( .A(n8374), .ZN(n8375) );
  NAND2_X1 U10698 ( .A1(n8375), .A2(SI_29_), .ZN(n8376) );
  MUX2_X1 U10699 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7171), .Z(n8378) );
  XNOR2_X1 U10700 ( .A(n8378), .B(SI_30_), .ZN(n8420) );
  MUX2_X1 U10701 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7171), .Z(n8379) );
  XNOR2_X1 U10702 ( .A(n8379), .B(SI_31_), .ZN(n8380) );
  NAND2_X1 U10703 ( .A1(n13501), .A2(n8423), .ZN(n8384) );
  INV_X1 U10704 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8382) );
  OR2_X1 U10705 ( .A1(n8162), .A2(n8382), .ZN(n8383) );
  INV_X1 U10706 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8388) );
  NAND2_X1 U10707 ( .A1(n8385), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8387) );
  NAND2_X1 U10708 ( .A1(n7815), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8386) );
  OAI211_X1 U10709 ( .C1(n8432), .C2(n8388), .A(n8387), .B(n8386), .ZN(n12986)
         );
  NAND2_X1 U10710 ( .A1(n13349), .A2(n8423), .ZN(n8394) );
  OR2_X1 U10711 ( .A1(n8162), .A2(n13350), .ZN(n8393) );
  INV_X1 U10712 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n11727) );
  NAND2_X1 U10713 ( .A1(n6441), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8398) );
  NAND2_X1 U10714 ( .A1(n8396), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8397) );
  OAI211_X1 U10715 ( .C1(n8399), .C2(n11727), .A(n8398), .B(n8397), .ZN(n8400)
         );
  INV_X1 U10716 ( .A(n8400), .ZN(n8401) );
  OAI21_X1 U10717 ( .B1(n11728), .B2(n8356), .A(n8401), .ZN(n12905) );
  AND2_X1 U10718 ( .A1(n12905), .A2(n8427), .ZN(n8402) );
  AOI21_X1 U10719 ( .B1(n13244), .B2(n8363), .A(n8402), .ZN(n8441) );
  NAND2_X1 U10720 ( .A1(n13244), .A2(n8403), .ZN(n8405) );
  NAND2_X1 U10721 ( .A1(n12905), .A2(n8363), .ZN(n8404) );
  NAND2_X1 U10722 ( .A1(n8405), .A2(n8404), .ZN(n8440) );
  NAND2_X1 U10723 ( .A1(n8441), .A2(n8440), .ZN(n8417) );
  INV_X1 U10724 ( .A(n8406), .ZN(n8409) );
  INV_X1 U10725 ( .A(n8407), .ZN(n8408) );
  AND2_X1 U10726 ( .A1(n8409), .A2(n8408), .ZN(n8414) );
  INV_X1 U10727 ( .A(n8410), .ZN(n8413) );
  INV_X1 U10728 ( .A(n8411), .ZN(n8412) );
  AOI22_X1 U10729 ( .A1(n8415), .A2(n8414), .B1(n8413), .B2(n8412), .ZN(n8416)
         );
  NAND2_X1 U10730 ( .A1(n12986), .A2(n8363), .ZN(n8449) );
  INV_X1 U10731 ( .A(n8420), .ZN(n8421) );
  NAND2_X1 U10732 ( .A1(n13512), .A2(n8423), .ZN(n8425) );
  INV_X1 U10733 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n11861) );
  OR2_X1 U10734 ( .A1(n8162), .A2(n11861), .ZN(n8424) );
  NAND2_X1 U10735 ( .A1(n6914), .A2(n8504), .ZN(n9776) );
  INV_X2 U10736 ( .A(n11222), .ZN(n13230) );
  NAND2_X1 U10737 ( .A1(n13230), .A2(n11372), .ZN(n9741) );
  OAI211_X1 U10738 ( .C1(n9776), .C2(n6795), .A(n9774), .B(n9741), .ZN(n8426)
         );
  AOI21_X1 U10739 ( .B1(n12986), .B2(n8427), .A(n8426), .ZN(n8436) );
  INV_X1 U10740 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8428) );
  OR2_X1 U10741 ( .A1(n8429), .A2(n8428), .ZN(n8435) );
  INV_X1 U10742 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8430) );
  OR2_X1 U10743 ( .A1(n8399), .A2(n8430), .ZN(n8434) );
  INV_X1 U10744 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8431) );
  OR2_X1 U10745 ( .A1(n8432), .A2(n8431), .ZN(n8433) );
  AND3_X1 U10746 ( .A1(n8435), .A2(n8434), .A3(n8433), .ZN(n8451) );
  NOR2_X1 U10747 ( .A1(n8436), .A2(n8451), .ZN(n8437) );
  AOI21_X1 U10748 ( .B1(n12992), .B2(n8363), .A(n8437), .ZN(n8447) );
  NAND2_X1 U10749 ( .A1(n12992), .A2(n8403), .ZN(n8439) );
  INV_X1 U10750 ( .A(n8451), .ZN(n12904) );
  NAND2_X1 U10751 ( .A1(n12904), .A2(n8363), .ZN(n8438) );
  NAND2_X1 U10752 ( .A1(n8439), .A2(n8438), .ZN(n8446) );
  OAI22_X1 U10753 ( .A1(n8447), .A2(n8446), .B1(n8441), .B2(n8440), .ZN(n8442)
         );
  NAND2_X1 U10754 ( .A1(n8443), .A2(n8442), .ZN(n8444) );
  OR2_X1 U10755 ( .A1(n12986), .A2(n8363), .ZN(n8448) );
  MUX2_X1 U10756 ( .A(n8449), .B(n8448), .S(n13237), .Z(n8450) );
  NAND2_X1 U10757 ( .A1(n13250), .A2(n13011), .ZN(n11724) );
  OR2_X1 U10758 ( .A1(n13250), .A2(n13011), .ZN(n8452) );
  NAND2_X1 U10759 ( .A1(n11724), .A2(n8452), .ZN(n12999) );
  INV_X1 U10760 ( .A(n13060), .ZN(n12895) );
  XNOR2_X1 U10761 ( .A(n13266), .B(n12895), .ZN(n13040) );
  XNOR2_X1 U10762 ( .A(n13269), .B(n13074), .ZN(n13056) );
  NAND2_X1 U10763 ( .A1(n13280), .A2(n12861), .ZN(n8453) );
  XNOR2_X1 U10764 ( .A(n13286), .B(n12865), .ZN(n13112) );
  INV_X1 U10765 ( .A(n13106), .ZN(n13140) );
  NAND2_X1 U10766 ( .A1(n13290), .A2(n13140), .ZN(n11690) );
  OR2_X1 U10767 ( .A1(n13290), .A2(n13140), .ZN(n8454) );
  NAND2_X1 U10768 ( .A1(n11690), .A2(n8454), .ZN(n13123) );
  INV_X1 U10769 ( .A(n13165), .ZN(n13138) );
  XNOR2_X1 U10770 ( .A(n13302), .B(n13138), .ZN(n13154) );
  OR2_X1 U10771 ( .A1(n13298), .A2(n13126), .ZN(n11715) );
  NAND2_X1 U10772 ( .A1(n13298), .A2(n13126), .ZN(n11714) );
  NAND2_X1 U10773 ( .A1(n11715), .A2(n11714), .ZN(n13135) );
  INV_X1 U10774 ( .A(n13224), .ZN(n11680) );
  XNOR2_X1 U10775 ( .A(n13318), .B(n11680), .ZN(n13199) );
  INV_X1 U10776 ( .A(n13323), .ZN(n11730) );
  NAND2_X1 U10777 ( .A1(n11730), .A2(n13203), .ZN(n8456) );
  INV_X1 U10778 ( .A(n13203), .ZN(n8455) );
  NAND2_X1 U10779 ( .A1(n13323), .A2(n8455), .ZN(n11679) );
  INV_X1 U10780 ( .A(n13226), .ZN(n8457) );
  OR2_X1 U10781 ( .A1(n11704), .A2(n8457), .ZN(n11678) );
  NAND2_X1 U10782 ( .A1(n11704), .A2(n8457), .ZN(n11675) );
  INV_X1 U10783 ( .A(n12907), .ZN(n11213) );
  NAND2_X1 U10784 ( .A1(n15027), .A2(n12908), .ZN(n11196) );
  OR2_X1 U10785 ( .A1(n15027), .A2(n12908), .ZN(n8458) );
  NAND2_X1 U10786 ( .A1(n11196), .A2(n8458), .ZN(n10895) );
  INV_X1 U10787 ( .A(n12911), .ZN(n10917) );
  XNOR2_X1 U10788 ( .A(n10872), .B(n10917), .ZN(n10563) );
  XNOR2_X1 U10789 ( .A(n15001), .B(n12912), .ZN(n10558) );
  NAND2_X1 U10790 ( .A1(n10126), .A2(n10036), .ZN(n8461) );
  OAI21_X1 U10791 ( .B1(n6445), .B2(n10167), .A(n6927), .ZN(n10093) );
  NAND3_X1 U10792 ( .A1(n10160), .A2(n10093), .A3(n6795), .ZN(n8460) );
  NOR2_X1 U10793 ( .A1(n8461), .A2(n8460), .ZN(n8462) );
  XNOR2_X1 U10794 ( .A(n10350), .B(n12913), .ZN(n10333) );
  XNOR2_X1 U10795 ( .A(n10240), .B(n12914), .ZN(n10238) );
  NAND4_X1 U10796 ( .A1(n10558), .A2(n8462), .A3(n10333), .A4(n10238), .ZN(
        n8463) );
  NOR2_X1 U10797 ( .A1(n10563), .A2(n8463), .ZN(n8465) );
  XNOR2_X1 U10798 ( .A(n15018), .B(n12910), .ZN(n10869) );
  NAND2_X1 U10799 ( .A1(n11089), .A2(n12909), .ZN(n10893) );
  OR2_X1 U10800 ( .A1(n11089), .A2(n12909), .ZN(n8464) );
  NAND2_X1 U10801 ( .A1(n10893), .A2(n8464), .ZN(n10877) );
  NAND4_X1 U10802 ( .A1(n10895), .A2(n8465), .A3(n10869), .A4(n10877), .ZN(
        n8466) );
  NOR2_X1 U10803 ( .A1(n11198), .A2(n8466), .ZN(n8467) );
  XNOR2_X1 U10804 ( .A(n11361), .B(n12906), .ZN(n11216) );
  NAND4_X1 U10805 ( .A1(n13222), .A2(n11363), .A3(n8467), .A4(n11216), .ZN(
        n8468) );
  NOR2_X1 U10806 ( .A1(n13199), .A2(n8468), .ZN(n8469) );
  XNOR2_X1 U10807 ( .A(n13307), .B(n13186), .ZN(n11712) );
  XNOR2_X1 U10808 ( .A(n13189), .B(n13204), .ZN(n13184) );
  NAND4_X1 U10809 ( .A1(n13135), .A2(n8469), .A3(n11712), .A4(n13184), .ZN(
        n8470) );
  OR3_X1 U10810 ( .A1(n13123), .A2(n13154), .A3(n8470), .ZN(n8471) );
  NOR2_X1 U10811 ( .A1(n13112), .A2(n8471), .ZN(n8472) );
  OR2_X1 U10812 ( .A1(n13275), .A2(n13087), .ZN(n11721) );
  NAND2_X1 U10813 ( .A1(n13275), .A2(n13087), .ZN(n11720) );
  NAND2_X1 U10814 ( .A1(n11721), .A2(n11720), .ZN(n13081) );
  NAND4_X1 U10815 ( .A1(n13056), .A2(n13091), .A3(n8472), .A4(n13081), .ZN(
        n8473) );
  NOR2_X1 U10816 ( .A1(n13040), .A2(n8473), .ZN(n8474) );
  XNOR2_X1 U10817 ( .A(n13259), .B(n13012), .ZN(n13034) );
  NAND4_X1 U10818 ( .A1(n12999), .A2(n8474), .A3(n13013), .A4(n13034), .ZN(
        n8476) );
  INV_X1 U10819 ( .A(n12905), .ZN(n8475) );
  XNOR2_X1 U10820 ( .A(n13244), .B(n8475), .ZN(n11725) );
  NAND3_X1 U10821 ( .A1(n7642), .A2(n8478), .A3(n8477), .ZN(n8483) );
  OAI21_X1 U10822 ( .B1(n8479), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8481) );
  XNOR2_X1 U10823 ( .A(n8481), .B(n8480), .ZN(n9685) );
  INV_X1 U10824 ( .A(n9685), .ZN(n9616) );
  NAND2_X1 U10825 ( .A1(n9616), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13370) );
  INV_X1 U10826 ( .A(n13370), .ZN(n8505) );
  MUX2_X1 U10827 ( .A(n11445), .B(n7762), .S(n11372), .Z(n8482) );
  NOR3_X1 U10828 ( .A1(n8482), .A2(n13370), .A3(n13230), .ZN(n8503) );
  NOR4_X1 U10829 ( .A1(n8483), .A2(n9774), .A3(n6914), .A4(n13370), .ZN(n8501)
         );
  INV_X1 U10830 ( .A(P2_B_REG_SCAN_IN), .ZN(n11697) );
  NAND2_X1 U10831 ( .A1(n8484), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8485) );
  MUX2_X1 U10832 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8485), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8487) );
  NAND2_X1 U10833 ( .A1(n8487), .A2(n8486), .ZN(n13361) );
  NAND2_X1 U10834 ( .A1(n8488), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8489) );
  MUX2_X1 U10835 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8489), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8490) );
  NAND2_X1 U10836 ( .A1(n8490), .A2(n8484), .ZN(n13363) );
  NOR2_X1 U10837 ( .A1(n13361), .A2(n13363), .ZN(n8496) );
  INV_X1 U10838 ( .A(n8491), .ZN(n8492) );
  OAI21_X1 U10839 ( .B1(n8493), .B2(n8492), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8494) );
  MUX2_X1 U10840 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8494), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8495) );
  NAND2_X1 U10841 ( .A1(n8496), .A2(n9727), .ZN(n9617) );
  AND2_X1 U10842 ( .A1(n9617), .A2(n9685), .ZN(n9738) );
  AND2_X1 U10843 ( .A1(n9738), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14998) );
  INV_X1 U10844 ( .A(n8497), .ZN(n8498) );
  NOR4_X1 U10845 ( .A1(n14995), .A2(n13356), .A3(n9741), .A4(n13139), .ZN(
        n8499) );
  AOI211_X1 U10846 ( .C1(n8505), .C2(n7762), .A(n11697), .B(n8499), .ZN(n8500)
         );
  INV_X1 U10847 ( .A(n9750), .ZN(n9752) );
  NOR2_X1 U10848 ( .A1(n9752), .A2(n8504), .ZN(n8507) );
  OAI21_X1 U10849 ( .B1(n6914), .B2(n11445), .A(n9741), .ZN(n8506) );
  OAI21_X1 U10850 ( .B1(n8507), .B2(n8506), .A(n8505), .ZN(n8508) );
  NAND3_X1 U10851 ( .A1(n8512), .A2(n8511), .A3(n8510), .ZN(P2_U3328) );
  NAND2_X1 U10852 ( .A1(n8641), .A2(n8650), .ZN(n8515) );
  NAND2_X1 U10853 ( .A1(n9653), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8514) );
  NAND2_X1 U10854 ( .A1(n8515), .A2(n8514), .ZN(n8663) );
  NAND2_X1 U10855 ( .A1(n9649), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8517) );
  INV_X1 U10856 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9628) );
  NAND2_X1 U10857 ( .A1(n9628), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8516) );
  AND2_X1 U10858 ( .A1(n8517), .A2(n8516), .ZN(n8662) );
  NAND2_X1 U10859 ( .A1(n9645), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8520) );
  INV_X1 U10860 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9630) );
  NAND2_X1 U10861 ( .A1(n9630), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U10862 ( .A1(n8520), .A2(n8518), .ZN(n8672) );
  INV_X1 U10863 ( .A(n8672), .ZN(n8519) );
  NAND2_X1 U10864 ( .A1(n9647), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8523) );
  INV_X1 U10865 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9637) );
  NAND2_X1 U10866 ( .A1(n9637), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8521) );
  NAND2_X1 U10867 ( .A1(n8523), .A2(n8521), .ZN(n8685) );
  INV_X1 U10868 ( .A(n8685), .ZN(n8522) );
  NAND2_X1 U10869 ( .A1(n9652), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8527) );
  INV_X1 U10870 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9642) );
  NAND2_X1 U10871 ( .A1(n9642), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8525) );
  NAND2_X1 U10872 ( .A1(n8527), .A2(n8525), .ZN(n8697) );
  INV_X1 U10873 ( .A(n8697), .ZN(n8526) );
  NAND2_X1 U10874 ( .A1(n9669), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8528) );
  NAND2_X1 U10875 ( .A1(n9673), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8530) );
  NAND2_X1 U10876 ( .A1(n9671), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8529) );
  NAND2_X1 U10877 ( .A1(n8530), .A2(n8529), .ZN(n8735) );
  NAND2_X1 U10878 ( .A1(n9677), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8532) );
  NAND2_X1 U10879 ( .A1(n9679), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8531) );
  NAND2_X1 U10880 ( .A1(n8751), .A2(n8532), .ZN(n8766) );
  NAND2_X1 U10881 ( .A1(n9682), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8534) );
  NAND2_X1 U10882 ( .A1(n9684), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U10883 ( .A1(n8766), .A2(n8765), .ZN(n8768) );
  NAND2_X1 U10884 ( .A1(n8768), .A2(n8534), .ZN(n8783) );
  NAND2_X1 U10885 ( .A1(n9770), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8536) );
  NAND2_X1 U10886 ( .A1(n9769), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8535) );
  NAND2_X1 U10887 ( .A1(n15329), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8537) );
  XNOR2_X1 U10888 ( .A(n8539), .B(P1_DATAO_REG_12__SCAN_IN), .ZN(n8813) );
  INV_X1 U10889 ( .A(n8813), .ZN(n8538) );
  NAND2_X1 U10890 ( .A1(n8539), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8540) );
  NAND2_X1 U10891 ( .A1(n8543), .A2(n8542), .ZN(n8544) );
  XNOR2_X1 U10892 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8838) );
  NAND2_X1 U10893 ( .A1(n8545), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8546) );
  XNOR2_X1 U10894 ( .A(n10756), .B(P1_DATAO_REG_15__SCAN_IN), .ZN(n8855) );
  INV_X1 U10895 ( .A(n8855), .ZN(n8548) );
  XNOR2_X1 U10896 ( .A(n10803), .B(P1_DATAO_REG_16__SCAN_IN), .ZN(n8868) );
  NAND2_X1 U10897 ( .A1(n10803), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8549) );
  XNOR2_X1 U10898 ( .A(n10819), .B(P1_DATAO_REG_17__SCAN_IN), .ZN(n8880) );
  INV_X1 U10899 ( .A(n8880), .ZN(n8550) );
  NAND2_X1 U10900 ( .A1(n10819), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8551) );
  XNOR2_X1 U10901 ( .A(n11034), .B(P1_DATAO_REG_18__SCAN_IN), .ZN(n8893) );
  INV_X1 U10902 ( .A(n8893), .ZN(n8552) );
  NAND2_X1 U10903 ( .A1(n11034), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8553) );
  XNOR2_X1 U10904 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .ZN(n8910) );
  NAND2_X1 U10905 ( .A1(n11125), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8554) );
  NAND2_X1 U10906 ( .A1(n8635), .A2(n11375), .ZN(n8557) );
  NAND2_X1 U10907 ( .A1(n8555), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8556) );
  INV_X1 U10908 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11448) );
  XNOR2_X1 U10909 ( .A(n11448), .B(P1_DATAO_REG_21__SCAN_IN), .ZN(n8622) );
  INV_X1 U10910 ( .A(n8622), .ZN(n8558) );
  NAND2_X1 U10911 ( .A1(n11448), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8559) );
  NAND2_X1 U10912 ( .A1(n15239), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8562) );
  INV_X1 U10913 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8560) );
  NAND2_X1 U10914 ( .A1(n8560), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U10915 ( .A1(n8562), .A2(n8561), .ZN(n8925) );
  NAND2_X1 U10916 ( .A1(n13373), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8564) );
  INV_X1 U10917 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n14319) );
  NAND2_X1 U10918 ( .A1(n14319), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8563) );
  INV_X1 U10919 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11547) );
  AND2_X1 U10920 ( .A1(n14313), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8568) );
  NAND2_X1 U10921 ( .A1(n13364), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8569) );
  NOR2_X1 U10922 ( .A1(n14307), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8570) );
  NAND2_X1 U10923 ( .A1(n14307), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8571) );
  INV_X1 U10924 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14306) );
  AOI22_X1 U10925 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n13358), .B2(n14306), .ZN(n8572) );
  XNOR2_X1 U10926 ( .A(n8991), .B(n8572), .ZN(n11253) );
  NOR2_X1 U10927 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), 
        .ZN(n8582) );
  NOR2_X1 U10928 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), 
        .ZN(n8581) );
  NAND2_X1 U10929 ( .A1(n9079), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8584) );
  NAND2_X1 U10930 ( .A1(n11253), .A2(n12079), .ZN(n8587) );
  NAND2_X1 U10931 ( .A1(n8664), .A2(SI_27_), .ZN(n8586) );
  NAND2_X1 U10932 ( .A1(n15117), .A2(n10463), .ZN(n8691) );
  INV_X1 U10933 ( .A(n8691), .ZN(n8588) );
  NAND2_X1 U10934 ( .A1(n8588), .A2(n10618), .ZN(n8708) );
  INV_X1 U10935 ( .A(n8758), .ZN(n8590) );
  INV_X1 U10936 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8595) );
  INV_X1 U10937 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8597) );
  INV_X1 U10938 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8599) );
  INV_X1 U10939 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8601) );
  INV_X1 U10940 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8603) );
  INV_X1 U10941 ( .A(n8982), .ZN(n8606) );
  INV_X1 U10942 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8605) );
  NAND2_X1 U10943 ( .A1(n8606), .A2(n8605), .ZN(n8996) );
  NAND2_X1 U10944 ( .A1(n8982), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8607) );
  NAND2_X1 U10945 ( .A1(n8996), .A2(n8607), .ZN(n12476) );
  NAND2_X1 U10946 ( .A1(n8608), .A2(n8611), .ZN(n11860) );
  XNOR2_X2 U10947 ( .A(n8609), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8615) );
  NAND2_X1 U10948 ( .A1(n12476), .A2(n9014), .ZN(n8621) );
  INV_X1 U10949 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n8618) );
  NAND2_X1 U10950 ( .A1(n9032), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8617) );
  NAND2_X1 U10951 ( .A1(n8638), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8616) );
  OAI211_X1 U10952 ( .C1(n8618), .C2(n10860), .A(n8617), .B(n8616), .ZN(n8619)
         );
  INV_X1 U10953 ( .A(n8619), .ZN(n8620) );
  XNOR2_X1 U10954 ( .A(n8623), .B(n8622), .ZN(n10438) );
  NAND2_X1 U10955 ( .A1(n10438), .A2(n6443), .ZN(n8625) );
  NAND2_X1 U10956 ( .A1(n8664), .A2(SI_21_), .ZN(n8624) );
  NAND2_X1 U10957 ( .A1(n8631), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U10958 ( .A1(n8931), .A2(n8626), .ZN(n12547) );
  NAND2_X1 U10959 ( .A1(n12547), .A2(n9014), .ZN(n8629) );
  AOI22_X1 U10960 ( .A1(n9032), .A2(P3_REG1_REG_21__SCAN_IN), .B1(n8638), .B2(
        P3_REG0_REG_21__SCAN_IN), .ZN(n8628) );
  INV_X1 U10961 ( .A(n10860), .ZN(n9033) );
  NAND2_X1 U10962 ( .A1(n9033), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8627) );
  INV_X1 U10963 ( .A(n12556), .ZN(n12276) );
  NAND2_X1 U10964 ( .A1(n8919), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8630) );
  NAND2_X1 U10965 ( .A1(n8631), .A2(n8630), .ZN(n12562) );
  NAND2_X1 U10966 ( .A1(n12562), .A2(n9014), .ZN(n8634) );
  AOI22_X1 U10967 ( .A1(n9032), .A2(P3_REG1_REG_20__SCAN_IN), .B1(n8638), .B2(
        P3_REG0_REG_20__SCAN_IN), .ZN(n8633) );
  NAND2_X1 U10968 ( .A1(n9033), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8632) );
  XNOR2_X1 U10969 ( .A(n8635), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n10180) );
  NAND2_X1 U10970 ( .A1(n10180), .A2(n6443), .ZN(n8637) );
  NAND2_X1 U10971 ( .A1(n8664), .A2(SI_20_), .ZN(n8636) );
  INV_X1 U10972 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10413) );
  INV_X1 U10973 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15155) );
  INV_X1 U10974 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10412) );
  NAND2_X1 U10975 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8642) );
  NAND2_X1 U10976 ( .A1(n8653), .A2(n10414), .ZN(n8643) );
  INV_X1 U10977 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10220) );
  INV_X1 U10978 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10411) );
  NOR2_X1 U10979 ( .A1(n8645), .A2(n6503), .ZN(n8649) );
  INV_X1 U10980 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n12287) );
  OR2_X1 U10981 ( .A1(n8639), .A2(n12287), .ZN(n8647) );
  NAND2_X1 U10982 ( .A1(n8638), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8646) );
  AND2_X1 U10983 ( .A1(n8647), .A2(n8646), .ZN(n8648) );
  INV_X1 U10984 ( .A(n8650), .ZN(n8652) );
  NAND2_X1 U10985 ( .A1(n9171), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U10986 ( .A1(n8652), .A2(n8651), .ZN(n9638) );
  NAND2_X1 U10987 ( .A1(n6443), .A2(n9638), .ZN(n8655) );
  NAND2_X1 U10988 ( .A1(n8653), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n8654) );
  NAND2_X1 U10989 ( .A1(n15148), .A2(n15147), .ZN(n15146) );
  OR2_X1 U10990 ( .A1(n15124), .A2(n7211), .ZN(n8656) );
  NAND2_X1 U10991 ( .A1(n8638), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8660) );
  INV_X1 U10992 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10710) );
  OR2_X1 U10993 ( .A1(n8644), .A2(n10710), .ZN(n8659) );
  INV_X1 U10994 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10469) );
  OR2_X1 U10995 ( .A1(n10860), .A2(n10469), .ZN(n8658) );
  INV_X1 U10996 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10468) );
  OR2_X1 U10997 ( .A1(n8639), .A2(n10468), .ZN(n8657) );
  OAI21_X1 U10998 ( .B1(n8663), .B2(n8662), .A(n8661), .ZN(n9659) );
  NAND2_X1 U10999 ( .A1(n8664), .A2(n9660), .ZN(n8666) );
  NAND2_X1 U11000 ( .A1(n10328), .A2(n15131), .ZN(n8667) );
  NAND2_X1 U11001 ( .A1(n8638), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8671) );
  OR2_X1 U11002 ( .A1(n8644), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8670) );
  INV_X1 U11003 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10475) );
  OR2_X1 U11004 ( .A1(n10860), .A2(n10475), .ZN(n8669) );
  INV_X1 U11005 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10474) );
  OR2_X1 U11006 ( .A1(n8639), .A2(n10474), .ZN(n8668) );
  XNOR2_X1 U11007 ( .A(n8673), .B(n8672), .ZN(n9624) );
  NAND2_X1 U11008 ( .A1(n8687), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8675) );
  INV_X1 U11009 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8674) );
  XNOR2_X1 U11010 ( .A(n8675), .B(n8674), .ZN(n10477) );
  NAND2_X1 U11011 ( .A1(n8653), .A2(n10477), .ZN(n8676) );
  OR2_X1 U11012 ( .A1(n15123), .A2(n15116), .ZN(n12138) );
  NAND2_X1 U11013 ( .A1(n15123), .A2(n15116), .ZN(n12137) );
  INV_X1 U11014 ( .A(n15110), .ZN(n12093) );
  NAND2_X1 U11015 ( .A1(n15123), .A2(n10330), .ZN(n8678) );
  NAND2_X1 U11016 ( .A1(n15109), .A2(n8678), .ZN(n10694) );
  NAND2_X1 U11017 ( .A1(n9032), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8684) );
  INV_X1 U11018 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8679) );
  OR2_X1 U11019 ( .A1(n7219), .A2(n8679), .ZN(n8683) );
  NAND2_X1 U11020 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8680) );
  AND2_X1 U11021 ( .A1(n8691), .A2(n8680), .ZN(n10698) );
  OR2_X1 U11022 ( .A1(n8644), .A2(n10698), .ZN(n8682) );
  OR2_X1 U11023 ( .A1(n10860), .A2(n10455), .ZN(n8681) );
  XNOR2_X1 U11024 ( .A(n8686), .B(n8685), .ZN(n9622) );
  INV_X1 U11025 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8699) );
  XNOR2_X1 U11026 ( .A(n8700), .B(n8699), .ZN(n10624) );
  NAND2_X1 U11027 ( .A1(n8653), .A2(n10624), .ZN(n8688) );
  XNOR2_X1 U11028 ( .A(n12143), .B(n15108), .ZN(n10693) );
  AND2_X1 U11029 ( .A1(n15108), .A2(n15174), .ZN(n8690) );
  AOI21_X1 U11030 ( .B1(n10694), .B2(n10693), .A(n8690), .ZN(n10810) );
  NAND2_X1 U11031 ( .A1(n8638), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8696) );
  INV_X1 U11032 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10613) );
  OR2_X1 U11033 ( .A1(n8639), .A2(n10613), .ZN(n8695) );
  NAND2_X1 U11034 ( .A1(n8691), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8692) );
  AND2_X1 U11035 ( .A1(n8708), .A2(n8692), .ZN(n10815) );
  OR2_X1 U11036 ( .A1(n8644), .A2(n10815), .ZN(n8694) );
  INV_X1 U11037 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10614) );
  OR2_X1 U11038 ( .A1(n10860), .A2(n10614), .ZN(n8693) );
  NAND4_X1 U11039 ( .A1(n8696), .A2(n8695), .A3(n8694), .A4(n8693), .ZN(n11993) );
  XNOR2_X1 U11040 ( .A(n8698), .B(n8697), .ZN(n9626) );
  NAND2_X1 U11041 ( .A1(n6443), .A2(n9626), .ZN(n8705) );
  NAND2_X1 U11042 ( .A1(n8701), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8703) );
  XNOR2_X1 U11043 ( .A(n8702), .B(n8703), .ZN(n10627) );
  NAND2_X1 U11044 ( .A1(n8653), .A2(n10627), .ZN(n8704) );
  OAI211_X1 U11045 ( .C1(n8793), .C2(SI_5_), .A(n8705), .B(n8704), .ZN(n11963)
         );
  OR2_X1 U11046 ( .A1(n11993), .A2(n11963), .ZN(n12149) );
  NAND2_X1 U11047 ( .A1(n11993), .A2(n11963), .ZN(n12150) );
  NAND2_X1 U11048 ( .A1(n12149), .A2(n12150), .ZN(n12146) );
  INV_X1 U11049 ( .A(n11993), .ZN(n10995) );
  NAND2_X1 U11050 ( .A1(n10995), .A2(n11963), .ZN(n8706) );
  NAND2_X1 U11051 ( .A1(n9032), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8714) );
  INV_X1 U11052 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8707) );
  OR2_X1 U11053 ( .A1(n7219), .A2(n8707), .ZN(n8713) );
  NAND2_X1 U11054 ( .A1(n8708), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8709) );
  AND2_X1 U11055 ( .A1(n8728), .A2(n8709), .ZN(n11113) );
  OR2_X1 U11056 ( .A1(n8644), .A2(n11113), .ZN(n8712) );
  INV_X1 U11057 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n8710) );
  OR2_X1 U11058 ( .A1(n10860), .A2(n8710), .ZN(n8711) );
  NAND4_X1 U11059 ( .A1(n8714), .A2(n8713), .A3(n8712), .A4(n8711), .ZN(n12284) );
  NAND2_X1 U11060 ( .A1(n8664), .A2(SI_6_), .ZN(n8724) );
  XNOR2_X1 U11061 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n8715) );
  XNOR2_X1 U11062 ( .A(n8716), .B(n8715), .ZN(n9662) );
  NAND2_X1 U11063 ( .A1(n12079), .A2(n9662), .ZN(n8723) );
  NOR2_X1 U11064 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n8717) );
  NAND2_X1 U11065 ( .A1(n8718), .A2(n8717), .ZN(n8720) );
  NAND2_X1 U11066 ( .A1(n8720), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8719) );
  MUX2_X1 U11067 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8719), .S(
        P3_IR_REG_6__SCAN_IN), .Z(n8721) );
  NAND2_X1 U11068 ( .A1(n8653), .A2(n10657), .ZN(n8722) );
  NAND2_X1 U11069 ( .A1(n12284), .A2(n11112), .ZN(n12153) );
  NAND2_X1 U11070 ( .A1(n12154), .A2(n12153), .ZN(n8725) );
  INV_X1 U11071 ( .A(n11112), .ZN(n10998) );
  NAND2_X1 U11072 ( .A1(n12284), .A2(n10998), .ZN(n8726) );
  NAND2_X1 U11073 ( .A1(n8638), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8734) );
  INV_X1 U11074 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n8727) );
  OR2_X1 U11075 ( .A1(n8639), .A2(n8727), .ZN(n8733) );
  NAND2_X1 U11076 ( .A1(n8728), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8729) );
  AND2_X1 U11077 ( .A1(n8742), .A2(n8729), .ZN(n11880) );
  OR2_X1 U11078 ( .A1(n8644), .A2(n11880), .ZN(n8732) );
  INV_X1 U11079 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n8730) );
  OR2_X1 U11080 ( .A1(n10860), .A2(n8730), .ZN(n8731) );
  XNOR2_X1 U11081 ( .A(n8736), .B(n8735), .ZN(n9620) );
  NAND2_X1 U11082 ( .A1(n12079), .A2(n9620), .ZN(n8739) );
  NAND2_X1 U11083 ( .A1(n8752), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8737) );
  XNOR2_X1 U11084 ( .A(n8737), .B(P3_IR_REG_7__SCAN_IN), .ZN(n15053) );
  INV_X1 U11085 ( .A(n15053), .ZN(n10944) );
  NAND2_X1 U11086 ( .A1(n8653), .A2(n10944), .ZN(n8738) );
  OAI211_X1 U11087 ( .C1(n8793), .C2(SI_7_), .A(n8739), .B(n8738), .ZN(n11167)
         );
  NAND2_X1 U11088 ( .A1(n12283), .A2(n11167), .ZN(n12160) );
  NAND2_X2 U11089 ( .A1(n12159), .A2(n12160), .ZN(n11165) );
  NAND2_X1 U11090 ( .A1(n11168), .A2(n11165), .ZN(n8741) );
  INV_X1 U11091 ( .A(n11167), .ZN(n11879) );
  NAND2_X1 U11092 ( .A1(n12283), .A2(n11879), .ZN(n8740) );
  NAND2_X1 U11093 ( .A1(n8638), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8747) );
  INV_X1 U11094 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n10942) );
  OR2_X1 U11095 ( .A1(n8639), .A2(n10942), .ZN(n8746) );
  NAND2_X1 U11096 ( .A1(n8742), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8743) );
  AND2_X1 U11097 ( .A1(n8758), .A2(n8743), .ZN(n11028) );
  OR2_X1 U11098 ( .A1(n8644), .A2(n11028), .ZN(n8745) );
  INV_X1 U11099 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10943) );
  OR2_X1 U11100 ( .A1(n10860), .A2(n10943), .ZN(n8744) );
  NAND4_X1 U11101 ( .A1(n8747), .A2(n8746), .A3(n8745), .A4(n8744), .ZN(n12282) );
  NAND2_X1 U11102 ( .A1(n8664), .A2(SI_8_), .ZN(n8756) );
  OR2_X1 U11103 ( .A1(n8749), .A2(n8748), .ZN(n8750) );
  AND2_X1 U11104 ( .A1(n8751), .A2(n8750), .ZN(n9631) );
  NAND2_X1 U11105 ( .A1(n12079), .A2(n9631), .ZN(n8755) );
  NAND2_X1 U11106 ( .A1(n8769), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8753) );
  XNOR2_X1 U11107 ( .A(n8753), .B(P3_IR_REG_8__SCAN_IN), .ZN(n11072) );
  NAND2_X1 U11108 ( .A1(n8653), .A2(n11072), .ZN(n8754) );
  NAND2_X1 U11109 ( .A1(n12282), .A2(n11027), .ZN(n12164) );
  NAND2_X1 U11110 ( .A1(n12165), .A2(n12164), .ZN(n11021) );
  NAND2_X1 U11111 ( .A1(n9032), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8764) );
  INV_X1 U11112 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n8757) );
  OR2_X1 U11113 ( .A1(n7219), .A2(n8757), .ZN(n8763) );
  NAND2_X1 U11114 ( .A1(n8758), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8759) );
  AND2_X1 U11115 ( .A1(n8775), .A2(n8759), .ZN(n12006) );
  OR2_X1 U11116 ( .A1(n8644), .A2(n12006), .ZN(n8762) );
  INV_X1 U11117 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n8760) );
  OR2_X1 U11118 ( .A1(n10860), .A2(n8760), .ZN(n8761) );
  NAND4_X1 U11119 ( .A1(n8764), .A2(n8763), .A3(n8762), .A4(n8761), .ZN(n12281) );
  OR2_X1 U11120 ( .A1(n8766), .A2(n8765), .ZN(n8767) );
  NAND2_X1 U11121 ( .A1(n8768), .A2(n8767), .ZN(n9634) );
  NAND2_X1 U11122 ( .A1(n12079), .A2(n9634), .ZN(n8772) );
  OAI21_X1 U11123 ( .B1(n8769), .B2(P3_IR_REG_8__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8770) );
  XNOR2_X1 U11124 ( .A(n8770), .B(P3_IR_REG_9__SCAN_IN), .ZN(n11419) );
  INV_X1 U11125 ( .A(n11419), .ZN(n11069) );
  NAND2_X1 U11126 ( .A1(n6883), .A2(n11069), .ZN(n8771) );
  OAI211_X1 U11127 ( .C1(n8793), .C2(SI_9_), .A(n8772), .B(n8771), .ZN(n11160)
         );
  INV_X1 U11128 ( .A(n11160), .ZN(n12005) );
  AND2_X1 U11129 ( .A1(n12281), .A2(n12005), .ZN(n8773) );
  OR2_X1 U11130 ( .A1(n12281), .A2(n11160), .ZN(n12169) );
  NAND2_X1 U11131 ( .A1(n12281), .A2(n11160), .ZN(n12170) );
  NAND2_X1 U11132 ( .A1(n12169), .A2(n12170), .ZN(n12091) );
  INV_X1 U11133 ( .A(n11027), .ZN(n11916) );
  OR2_X1 U11134 ( .A1(n12282), .A2(n11916), .ZN(n11153) );
  AND2_X1 U11135 ( .A1(n12091), .A2(n11153), .ZN(n11154) );
  NAND2_X1 U11136 ( .A1(n9032), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8781) );
  INV_X1 U11137 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n8774) );
  OR2_X1 U11138 ( .A1(n7219), .A2(n8774), .ZN(n8780) );
  NAND2_X1 U11139 ( .A1(n8775), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8776) );
  AND2_X1 U11140 ( .A1(n8796), .A2(n8776), .ZN(n11235) );
  OR2_X1 U11141 ( .A1(n8644), .A2(n11235), .ZN(n8779) );
  INV_X1 U11142 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n8777) );
  OR2_X1 U11143 ( .A1(n10860), .A2(n8777), .ZN(n8778) );
  NAND4_X1 U11144 ( .A1(n8781), .A2(n8780), .A3(n8779), .A4(n8778), .ZN(n12280) );
  OR2_X1 U11145 ( .A1(n8783), .A2(n8782), .ZN(n8784) );
  NAND2_X1 U11146 ( .A1(n8785), .A2(n8784), .ZN(n9657) );
  NAND2_X1 U11147 ( .A1(n12079), .A2(n9657), .ZN(n8792) );
  NAND2_X1 U11148 ( .A1(n8786), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8787) );
  MUX2_X1 U11149 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8787), .S(
        P3_IR_REG_10__SCAN_IN), .Z(n8790) );
  INV_X1 U11150 ( .A(n8788), .ZN(n8789) );
  NAND2_X1 U11151 ( .A1(n8790), .A2(n8789), .ZN(n15067) );
  NAND2_X1 U11152 ( .A1(n6883), .A2(n15067), .ZN(n8791) );
  OAI211_X1 U11153 ( .C1(n8793), .C2(SI_10_), .A(n8792), .B(n8791), .ZN(n11234) );
  OR2_X1 U11154 ( .A1(n12280), .A2(n11234), .ZN(n12174) );
  NAND2_X1 U11155 ( .A1(n12280), .A2(n11234), .ZN(n12181) );
  NAND2_X1 U11156 ( .A1(n12174), .A2(n12181), .ZN(n12096) );
  INV_X1 U11157 ( .A(n11234), .ZN(n11147) );
  NAND2_X1 U11158 ( .A1(n12280), .A2(n11147), .ZN(n8794) );
  NAND2_X1 U11159 ( .A1(n8638), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8802) );
  INV_X1 U11160 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11336) );
  OR2_X1 U11161 ( .A1(n10860), .A2(n11336), .ZN(n8801) );
  NAND2_X1 U11162 ( .A1(n8796), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8797) );
  AND2_X1 U11163 ( .A1(n8819), .A2(n8797), .ZN(n11440) );
  OR2_X1 U11164 ( .A1(n8644), .A2(n11440), .ZN(n8800) );
  INV_X1 U11165 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n8798) );
  OR2_X1 U11166 ( .A1(n8639), .A2(n8798), .ZN(n8799) );
  NAND4_X1 U11167 ( .A1(n8802), .A2(n8801), .A3(n8800), .A4(n8799), .ZN(n12279) );
  XNOR2_X1 U11168 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8803) );
  XNOR2_X1 U11169 ( .A(n8804), .B(n8803), .ZN(n9655) );
  NAND2_X1 U11170 ( .A1(n9655), .A2(n12079), .ZN(n8811) );
  NOR2_X1 U11171 ( .A1(n8788), .A2(n9027), .ZN(n8805) );
  MUX2_X1 U11172 ( .A(n9027), .B(n8805), .S(P3_IR_REG_11__SCAN_IN), .Z(n8806)
         );
  INV_X1 U11173 ( .A(n8806), .ZN(n8809) );
  INV_X1 U11174 ( .A(n8807), .ZN(n8808) );
  NAND2_X1 U11175 ( .A1(n8809), .A2(n8808), .ZN(n11423) );
  AOI22_X1 U11176 ( .A1(n8664), .A2(n9656), .B1(n6883), .B2(n11423), .ZN(n8810) );
  INV_X1 U11177 ( .A(n12279), .ZN(n11435) );
  NAND2_X1 U11178 ( .A1(n11435), .A2(n14529), .ZN(n8812) );
  XNOR2_X1 U11179 ( .A(n8814), .B(n8813), .ZN(n9675) );
  NAND2_X1 U11180 ( .A1(n9675), .A2(n12079), .ZN(n8817) );
  OR2_X1 U11181 ( .A1(n8807), .A2(n9027), .ZN(n8815) );
  XNOR2_X1 U11182 ( .A(n8815), .B(P3_IR_REG_12__SCAN_IN), .ZN(n15083) );
  AOI22_X1 U11183 ( .A1(n8664), .A2(SI_12_), .B1(n6883), .B2(n15083), .ZN(
        n8816) );
  NAND2_X1 U11184 ( .A1(n9032), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8824) );
  INV_X1 U11185 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n8818) );
  OR2_X1 U11186 ( .A1(n7219), .A2(n8818), .ZN(n8823) );
  NAND2_X1 U11187 ( .A1(n8819), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8820) );
  AND2_X1 U11188 ( .A1(n8831), .A2(n8820), .ZN(n11942) );
  OR2_X1 U11189 ( .A1(n8644), .A2(n11942), .ZN(n8822) );
  INV_X1 U11190 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12301) );
  OR2_X1 U11191 ( .A1(n10860), .A2(n12301), .ZN(n8821) );
  NAND4_X1 U11192 ( .A1(n8824), .A2(n8823), .A3(n8822), .A4(n8821), .ZN(n14508) );
  NAND2_X1 U11193 ( .A1(n11619), .A2(n14508), .ZN(n12180) );
  INV_X1 U11194 ( .A(n14508), .ZN(n11620) );
  NAND2_X1 U11195 ( .A1(n11620), .A2(n14524), .ZN(n12184) );
  NAND2_X1 U11196 ( .A1(n14524), .A2(n14508), .ZN(n8825) );
  XNOR2_X1 U11197 ( .A(n8826), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n9680) );
  NAND2_X1 U11198 ( .A1(n9680), .A2(n12079), .ZN(n8830) );
  INV_X1 U11199 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8827) );
  NAND2_X1 U11200 ( .A1(n8807), .A2(n8827), .ZN(n8840) );
  NAND2_X1 U11201 ( .A1(n8840), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8828) );
  XNOR2_X1 U11202 ( .A(n8828), .B(P3_IR_REG_13__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U11203 ( .A1(n8664), .A2(SI_13_), .B1(n6883), .B2(n12336), .ZN(
        n8829) );
  NAND2_X1 U11204 ( .A1(n8830), .A2(n8829), .ZN(n14512) );
  NAND2_X1 U11205 ( .A1(n8638), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8836) );
  INV_X1 U11206 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12305) );
  OR2_X1 U11207 ( .A1(n8639), .A2(n12305), .ZN(n8835) );
  NAND2_X1 U11208 ( .A1(n8831), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8832) );
  AND2_X1 U11209 ( .A1(n8847), .A2(n8832), .ZN(n14513) );
  OR2_X1 U11210 ( .A1(n8644), .A2(n14513), .ZN(n8834) );
  INV_X1 U11211 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12306) );
  OR2_X1 U11212 ( .A1(n10860), .A2(n12306), .ZN(n8833) );
  OR2_X1 U11213 ( .A1(n14512), .A2(n12643), .ZN(n12188) );
  NAND2_X1 U11214 ( .A1(n14512), .A2(n12643), .ZN(n12189) );
  NAND2_X1 U11215 ( .A1(n12188), .A2(n12189), .ZN(n14505) );
  NAND2_X1 U11216 ( .A1(n14506), .A2(n14505), .ZN(n14504) );
  INV_X1 U11217 ( .A(n12643), .ZN(n12278) );
  NAND2_X1 U11218 ( .A1(n14512), .A2(n12278), .ZN(n8837) );
  XNOR2_X1 U11219 ( .A(n8839), .B(n8838), .ZN(n9700) );
  NAND2_X1 U11220 ( .A1(n9700), .A2(n12079), .ZN(n8846) );
  NOR2_X1 U11221 ( .A1(n8840), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n8843) );
  OR2_X1 U11222 ( .A1(n8843), .A2(n9027), .ZN(n8841) );
  MUX2_X1 U11223 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8841), .S(
        P3_IR_REG_14__SCAN_IN), .Z(n8844) );
  NAND2_X1 U11224 ( .A1(n8843), .A2(n8842), .ZN(n8858) );
  NAND2_X1 U11225 ( .A1(n8844), .A2(n8858), .ZN(n12344) );
  AOI22_X1 U11226 ( .A1(n8664), .A2(n9701), .B1(n6883), .B2(n12344), .ZN(n8845) );
  NAND2_X1 U11227 ( .A1(n8846), .A2(n8845), .ZN(n12775) );
  NAND2_X1 U11228 ( .A1(n9032), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8853) );
  INV_X1 U11229 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12773) );
  OR2_X1 U11230 ( .A1(n7219), .A2(n12773), .ZN(n8852) );
  NAND2_X1 U11231 ( .A1(n8847), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8848) );
  AND2_X1 U11232 ( .A1(n8862), .A2(n8848), .ZN(n11889) );
  OR2_X1 U11233 ( .A1(n8644), .A2(n11889), .ZN(n8851) );
  INV_X1 U11234 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n8849) );
  OR2_X1 U11235 ( .A1(n10860), .A2(n8849), .ZN(n8850) );
  NAND4_X1 U11236 ( .A1(n8853), .A2(n8852), .A3(n8851), .A4(n8850), .ZN(n14507) );
  OR2_X1 U11237 ( .A1(n12775), .A2(n14507), .ZN(n12192) );
  NAND2_X1 U11238 ( .A1(n12775), .A2(n14507), .ZN(n12193) );
  NAND2_X1 U11239 ( .A1(n12192), .A2(n12193), .ZN(n12640) );
  INV_X1 U11240 ( .A(n14507), .ZN(n12025) );
  OR2_X1 U11241 ( .A1(n12775), .A2(n12025), .ZN(n8854) );
  XNOR2_X1 U11242 ( .A(n8856), .B(n8855), .ZN(n9748) );
  NAND2_X1 U11243 ( .A1(n9748), .A2(n6443), .ZN(n8861) );
  NAND2_X1 U11244 ( .A1(n8858), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8857) );
  MUX2_X1 U11245 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8857), .S(
        P3_IR_REG_15__SCAN_IN), .Z(n8859) );
  AOI22_X1 U11246 ( .A1(n8664), .A2(SI_15_), .B1(n6883), .B2(n12370), .ZN(
        n8860) );
  NAND2_X1 U11247 ( .A1(n8861), .A2(n8860), .ZN(n12067) );
  NAND2_X1 U11248 ( .A1(n8638), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8867) );
  INV_X1 U11249 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14482) );
  OR2_X1 U11250 ( .A1(n10860), .A2(n14482), .ZN(n8866) );
  NAND2_X1 U11251 ( .A1(n8862), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8863) );
  AND2_X1 U11252 ( .A1(n8873), .A2(n8863), .ZN(n12061) );
  OR2_X1 U11253 ( .A1(n8644), .A2(n12061), .ZN(n8865) );
  INV_X1 U11254 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14487) );
  OR2_X1 U11255 ( .A1(n8639), .A2(n14487), .ZN(n8864) );
  OR2_X1 U11256 ( .A1(n12067), .A2(n12647), .ZN(n12196) );
  NAND2_X1 U11257 ( .A1(n12067), .A2(n12647), .ZN(n12200) );
  NAND2_X1 U11258 ( .A1(n12196), .A2(n12200), .ZN(n12624) );
  INV_X1 U11259 ( .A(n12647), .ZN(n12610) );
  XNOR2_X1 U11260 ( .A(n8869), .B(n8868), .ZN(n9788) );
  NAND2_X1 U11261 ( .A1(n9788), .A2(n12079), .ZN(n8872) );
  NAND2_X1 U11262 ( .A1(n8882), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8870) );
  XNOR2_X1 U11263 ( .A(n8870), .B(P3_IR_REG_16__SCAN_IN), .ZN(n12373) );
  AOI22_X1 U11264 ( .A1(n8664), .A2(SI_16_), .B1(n6883), .B2(n12373), .ZN(
        n8871) );
  NAND2_X1 U11265 ( .A1(n8872), .A2(n8871), .ZN(n12616) );
  NAND2_X1 U11266 ( .A1(n8638), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8878) );
  INV_X1 U11267 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12713) );
  OR2_X1 U11268 ( .A1(n8639), .A2(n12713), .ZN(n8877) );
  NAND2_X1 U11269 ( .A1(n8873), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8874) );
  AND2_X1 U11270 ( .A1(n8886), .A2(n8874), .ZN(n12617) );
  OR2_X1 U11271 ( .A1(n8644), .A2(n12617), .ZN(n8876) );
  INV_X1 U11272 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12618) );
  OR2_X1 U11273 ( .A1(n10860), .A2(n12618), .ZN(n8875) );
  OR2_X1 U11274 ( .A1(n12616), .A2(n12066), .ZN(n12202) );
  NAND2_X1 U11275 ( .A1(n12616), .A2(n12066), .ZN(n12201) );
  NAND2_X1 U11276 ( .A1(n12202), .A2(n12201), .ZN(n12608) );
  NAND2_X1 U11277 ( .A1(n12616), .A2(n12626), .ZN(n8879) );
  NAND2_X1 U11278 ( .A1(n12607), .A2(n8879), .ZN(n12595) );
  XNOR2_X1 U11279 ( .A(n8881), .B(n8880), .ZN(n9911) );
  NAND2_X1 U11280 ( .A1(n9911), .A2(n6443), .ZN(n8885) );
  OAI21_X1 U11281 ( .B1(n8882), .B2(P3_IR_REG_16__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8883) );
  XNOR2_X1 U11282 ( .A(n8883), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12417) );
  AOI22_X1 U11283 ( .A1(n8664), .A2(SI_17_), .B1(n6883), .B2(n12417), .ZN(
        n8884) );
  NAND2_X1 U11284 ( .A1(n8885), .A2(n8884), .ZN(n11971) );
  NAND2_X1 U11285 ( .A1(n8638), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8891) );
  INV_X1 U11286 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12602) );
  OR2_X1 U11287 ( .A1(n10860), .A2(n12602), .ZN(n8890) );
  NAND2_X1 U11288 ( .A1(n8886), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8887) );
  AND2_X1 U11289 ( .A1(n8901), .A2(n8887), .ZN(n12601) );
  OR2_X1 U11290 ( .A1(n8644), .A2(n12601), .ZN(n8889) );
  INV_X1 U11291 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12709) );
  OR2_X1 U11292 ( .A1(n8639), .A2(n12709), .ZN(n8888) );
  OR2_X1 U11293 ( .A1(n11971), .A2(n12583), .ZN(n12207) );
  NAND2_X1 U11294 ( .A1(n11971), .A2(n12583), .ZN(n12209) );
  NAND2_X1 U11295 ( .A1(n12207), .A2(n12209), .ZN(n12594) );
  INV_X1 U11296 ( .A(n12583), .ZN(n12611) );
  NAND2_X1 U11297 ( .A1(n11971), .A2(n12611), .ZN(n8892) );
  XNOR2_X1 U11298 ( .A(n8894), .B(n8893), .ZN(n9939) );
  NAND2_X1 U11299 ( .A1(n9939), .A2(n6443), .ZN(n8900) );
  NAND2_X1 U11300 ( .A1(n8895), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8896) );
  MUX2_X1 U11301 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8896), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n8898) );
  INV_X1 U11302 ( .A(n8897), .ZN(n8912) );
  AND2_X1 U11303 ( .A1(n8898), .A2(n8912), .ZN(n12432) );
  AOI22_X1 U11304 ( .A1(n8664), .A2(SI_18_), .B1(n6883), .B2(n12432), .ZN(
        n8899) );
  NAND2_X1 U11305 ( .A1(n8900), .A2(n8899), .ZN(n12040) );
  NAND2_X1 U11306 ( .A1(n8901), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8902) );
  NAND2_X1 U11307 ( .A1(n8917), .A2(n8902), .ZN(n12588) );
  NAND2_X1 U11308 ( .A1(n9014), .A2(n12588), .ZN(n8906) );
  INV_X1 U11309 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12705) );
  OR2_X1 U11310 ( .A1(n8639), .A2(n12705), .ZN(n8905) );
  INV_X1 U11311 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n15282) );
  OR2_X1 U11312 ( .A1(n7219), .A2(n15282), .ZN(n8904) );
  INV_X1 U11313 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12411) );
  OR2_X1 U11314 ( .A1(n10860), .A2(n12411), .ZN(n8903) );
  NAND2_X1 U11315 ( .A1(n12040), .A2(n11976), .ZN(n12211) );
  OR2_X1 U11316 ( .A1(n12040), .A2(n12596), .ZN(n8909) );
  XNOR2_X1 U11317 ( .A(n8911), .B(n8910), .ZN(n9943) );
  NAND2_X1 U11318 ( .A1(n9943), .A2(n6443), .ZN(n8916) );
  AOI22_X1 U11319 ( .A1(n8664), .A2(n9942), .B1(n6883), .B2(n12428), .ZN(n8915) );
  NAND2_X1 U11320 ( .A1(n8917), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8918) );
  NAND2_X1 U11321 ( .A1(n8919), .A2(n8918), .ZN(n12572) );
  NAND2_X1 U11322 ( .A1(n12572), .A2(n9014), .ZN(n8924) );
  NAND2_X1 U11323 ( .A1(n9032), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8923) );
  INV_X1 U11324 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n15280) );
  OR2_X1 U11325 ( .A1(n7219), .A2(n15280), .ZN(n8922) );
  INV_X1 U11326 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n8920) );
  OR2_X1 U11327 ( .A1(n10860), .A2(n8920), .ZN(n8921) );
  NAND4_X1 U11328 ( .A1(n8924), .A2(n8923), .A3(n8922), .A4(n8921), .ZN(n12277) );
  OR2_X1 U11329 ( .A1(n12756), .A2(n12277), .ZN(n12218) );
  NAND2_X1 U11330 ( .A1(n12756), .A2(n12277), .ZN(n12219) );
  XNOR2_X1 U11331 ( .A(n12223), .B(n12222), .ZN(n12552) );
  NAND2_X1 U11332 ( .A1(n12690), .A2(n12556), .ZN(n12230) );
  NAND2_X1 U11333 ( .A1(n12229), .A2(n12230), .ZN(n12545) );
  NAND2_X1 U11334 ( .A1(n8926), .A2(n8925), .ZN(n8927) );
  NAND2_X1 U11335 ( .A1(n8928), .A2(n8927), .ZN(n14435) );
  NAND2_X1 U11336 ( .A1(n14435), .A2(n6443), .ZN(n8930) );
  NAND2_X1 U11337 ( .A1(n8664), .A2(SI_22_), .ZN(n8929) );
  NAND2_X1 U11338 ( .A1(n8931), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8932) );
  NAND2_X1 U11339 ( .A1(n8946), .A2(n8932), .ZN(n12536) );
  NAND2_X1 U11340 ( .A1(n12536), .A2(n9014), .ZN(n8938) );
  INV_X1 U11341 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n8935) );
  NAND2_X1 U11342 ( .A1(n9032), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8934) );
  NAND2_X1 U11343 ( .A1(n8638), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8933) );
  OAI211_X1 U11344 ( .C1(n8935), .C2(n10860), .A(n8934), .B(n8933), .ZN(n8936)
         );
  INV_X1 U11345 ( .A(n8936), .ZN(n8937) );
  NOR2_X1 U11346 ( .A1(n12037), .A2(n12543), .ZN(n8939) );
  OR2_X1 U11347 ( .A1(n8941), .A2(n8940), .ZN(n8942) );
  NAND2_X1 U11348 ( .A1(n8943), .A2(n8942), .ZN(n10771) );
  NAND2_X1 U11349 ( .A1(n10771), .A2(n6443), .ZN(n8945) );
  NAND2_X1 U11350 ( .A1(n8664), .A2(SI_23_), .ZN(n8944) );
  NAND2_X1 U11351 ( .A1(n8946), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8947) );
  NAND2_X1 U11352 ( .A1(n8956), .A2(n8947), .ZN(n12524) );
  NAND2_X1 U11353 ( .A1(n12524), .A2(n9014), .ZN(n8952) );
  INV_X1 U11354 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12526) );
  NAND2_X1 U11355 ( .A1(n9032), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8949) );
  NAND2_X1 U11356 ( .A1(n8638), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8948) );
  OAI211_X1 U11357 ( .C1(n12526), .C2(n10860), .A(n8949), .B(n8948), .ZN(n8950) );
  INV_X1 U11358 ( .A(n8950), .ZN(n8951) );
  NAND2_X1 U11359 ( .A1(n12680), .A2(n12533), .ZN(n12114) );
  NAND2_X1 U11360 ( .A1(n12110), .A2(n12114), .ZN(n12090) );
  XNOR2_X1 U11361 ( .A(n8953), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n11036) );
  NAND2_X1 U11362 ( .A1(n11036), .A2(n6443), .ZN(n8955) );
  NAND2_X1 U11363 ( .A1(n8664), .A2(SI_24_), .ZN(n8954) );
  NAND2_X1 U11364 ( .A1(n8956), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8957) );
  NAND2_X1 U11365 ( .A1(n8968), .A2(n8957), .ZN(n12512) );
  NAND2_X1 U11366 ( .A1(n12512), .A2(n9014), .ZN(n8963) );
  INV_X1 U11367 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n8960) );
  NAND2_X1 U11368 ( .A1(n9032), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8959) );
  NAND2_X1 U11369 ( .A1(n8638), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8958) );
  OAI211_X1 U11370 ( .C1(n8960), .C2(n10860), .A(n8959), .B(n8958), .ZN(n8961)
         );
  INV_X1 U11371 ( .A(n8961), .ZN(n8962) );
  INV_X1 U11372 ( .A(n12676), .ZN(n12514) );
  XNOR2_X1 U11373 ( .A(n13364), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8964) );
  XNOR2_X1 U11374 ( .A(n8965), .B(n8964), .ZN(n11001) );
  NAND2_X1 U11375 ( .A1(n11001), .A2(n6443), .ZN(n8967) );
  NAND2_X1 U11376 ( .A1(n8664), .A2(SI_25_), .ZN(n8966) );
  NAND2_X1 U11377 ( .A1(n8968), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8969) );
  NAND2_X1 U11378 ( .A1(n8980), .A2(n8969), .ZN(n12501) );
  NAND2_X1 U11379 ( .A1(n12501), .A2(n9014), .ZN(n8975) );
  INV_X1 U11380 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n8972) );
  NAND2_X1 U11381 ( .A1(n9032), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8971) );
  NAND2_X1 U11382 ( .A1(n8638), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8970) );
  OAI211_X1 U11383 ( .C1(n8972), .C2(n10860), .A(n8971), .B(n8970), .ZN(n8973)
         );
  INV_X1 U11384 ( .A(n8973), .ZN(n8974) );
  XNOR2_X1 U11385 ( .A(n12240), .B(n12484), .ZN(n12493) );
  AOI22_X1 U11386 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(
        P1_DATAO_REG_26__SCAN_IN), .B1(n13360), .B2(n14307), .ZN(n8976) );
  XNOR2_X1 U11387 ( .A(n8977), .B(n8976), .ZN(n11150) );
  NAND2_X1 U11388 ( .A1(n8664), .A2(SI_26_), .ZN(n8978) );
  NAND2_X1 U11389 ( .A1(n8980), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8981) );
  NAND2_X1 U11390 ( .A1(n8982), .A2(n8981), .ZN(n12487) );
  NAND2_X1 U11391 ( .A1(n12487), .A2(n9014), .ZN(n8988) );
  INV_X1 U11392 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n8985) );
  NAND2_X1 U11393 ( .A1(n8638), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8984) );
  NAND2_X1 U11394 ( .A1(n9032), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8983) );
  OAI211_X1 U11395 ( .C1(n8985), .C2(n10860), .A(n8984), .B(n8983), .ZN(n8986)
         );
  INV_X1 U11396 ( .A(n8986), .ZN(n8987) );
  NAND2_X1 U11397 ( .A1(n12735), .A2(n12497), .ZN(n8989) );
  INV_X1 U11398 ( .A(n12497), .ZN(n12274) );
  XNOR2_X1 U11399 ( .A(n12477), .B(n12483), .ZN(n12471) );
  NOR2_X1 U11400 ( .A1(n13358), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8990) );
  NAND2_X1 U11401 ( .A1(n13358), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8992) );
  XNOR2_X1 U11402 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .ZN(n8993) );
  XNOR2_X1 U11403 ( .A(n9005), .B(n8993), .ZN(n11511) );
  NAND2_X1 U11404 ( .A1(n11511), .A2(n6443), .ZN(n8995) );
  NAND2_X1 U11405 ( .A1(n8664), .A2(SI_28_), .ZN(n8994) );
  NAND2_X1 U11406 ( .A1(n8996), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8997) );
  NAND2_X1 U11407 ( .A1(n9013), .A2(n8997), .ZN(n12463) );
  INV_X1 U11408 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n15319) );
  NAND2_X1 U11409 ( .A1(n9032), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8999) );
  NAND2_X1 U11410 ( .A1(n9033), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8998) );
  OAI211_X1 U11411 ( .C1(n7219), .C2(n15319), .A(n8999), .B(n8998), .ZN(n9000)
         );
  NAND2_X1 U11412 ( .A1(n12659), .A2(n12472), .ZN(n12254) );
  NAND2_X1 U11413 ( .A1(n12255), .A2(n12254), .ZN(n12456) );
  NAND2_X1 U11414 ( .A1(n12455), .A2(n12456), .ZN(n12457) );
  INV_X1 U11415 ( .A(n12659), .ZN(n11670) );
  INV_X1 U11416 ( .A(n12472), .ZN(n9001) );
  NAND2_X1 U11417 ( .A1(n12457), .A2(n9002), .ZN(n9020) );
  AND2_X1 U11418 ( .A1(n9003), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9004) );
  NAND2_X1 U11419 ( .A1(n11549), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9006) );
  XNOR2_X1 U11420 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n9007) );
  OR2_X1 U11421 ( .A1(n9008), .A2(n9007), .ZN(n9009) );
  NAND2_X1 U11422 ( .A1(n11852), .A2(n9009), .ZN(n11514) );
  OR2_X1 U11423 ( .A1(n11514), .A2(n9010), .ZN(n9012) );
  NAND2_X1 U11424 ( .A1(n8664), .A2(SI_29_), .ZN(n9011) );
  NAND2_X1 U11425 ( .A1(n11863), .A2(n9014), .ZN(n10863) );
  INV_X1 U11426 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n15246) );
  NAND2_X1 U11427 ( .A1(n8638), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9016) );
  NAND2_X1 U11428 ( .A1(n9032), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9015) );
  OAI211_X1 U11429 ( .C1(n15246), .C2(n10860), .A(n9016), .B(n9015), .ZN(n9017) );
  INV_X1 U11430 ( .A(n9017), .ZN(n9018) );
  NAND2_X1 U11431 ( .A1(n11866), .A2(n12458), .ZN(n12083) );
  NAND2_X1 U11432 ( .A1(n12258), .A2(n12083), .ZN(n9059) );
  INV_X1 U11433 ( .A(n9059), .ZN(n9019) );
  XNOR2_X1 U11434 ( .A(n9020), .B(n9019), .ZN(n9041) );
  NAND2_X1 U11435 ( .A1(n9022), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9021) );
  MUX2_X1 U11436 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9021), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n9023) );
  NAND2_X1 U11437 ( .A1(n12127), .A2(n10193), .ZN(n12089) );
  INV_X1 U11438 ( .A(n9031), .ZN(n12268) );
  INV_X1 U11439 ( .A(n6446), .ZN(n10408) );
  NAND2_X1 U11440 ( .A1(n12268), .A2(n10408), .ZN(n10397) );
  NAND2_X1 U11441 ( .A1(n10397), .A2(n10395), .ZN(n9038) );
  INV_X1 U11442 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14534) );
  NAND2_X1 U11443 ( .A1(n9032), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9035) );
  NAND2_X1 U11444 ( .A1(n9033), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9034) );
  OAI211_X1 U11445 ( .C1(n7219), .C2(n14534), .A(n9035), .B(n9034), .ZN(n9036)
         );
  INV_X1 U11446 ( .A(n9036), .ZN(n9037) );
  AND2_X1 U11447 ( .A1(n10863), .A2(n9037), .ZN(n12086) );
  AND2_X1 U11448 ( .A1(n12268), .A2(P3_B_REG_SCAN_IN), .ZN(n9039) );
  OR2_X1 U11449 ( .A1(n12646), .A2(n9039), .ZN(n12449) );
  OAI22_X1 U11450 ( .A1(n12472), .A2(n12642), .B1(n12086), .B2(n12449), .ZN(
        n9040) );
  INV_X1 U11451 ( .A(n10268), .ZN(n10284) );
  NAND2_X1 U11452 ( .A1(n10198), .A2(n12122), .ZN(n15122) );
  OR2_X1 U11453 ( .A1(n15144), .A2(n15131), .ZN(n12130) );
  NAND2_X1 U11454 ( .A1(n15107), .A2(n12093), .ZN(n9043) );
  NAND2_X1 U11455 ( .A1(n9043), .A2(n12138), .ZN(n10690) );
  NAND2_X1 U11456 ( .A1(n10690), .A2(n12141), .ZN(n10692) );
  OR2_X1 U11457 ( .A1(n15108), .A2(n12143), .ZN(n12145) );
  NAND2_X1 U11458 ( .A1(n10692), .A2(n12145), .ZN(n10808) );
  INV_X1 U11459 ( .A(n12146), .ZN(n12095) );
  NAND2_X1 U11460 ( .A1(n10808), .A2(n12095), .ZN(n9044) );
  NAND2_X1 U11461 ( .A1(n9044), .A2(n12149), .ZN(n11109) );
  INV_X1 U11462 ( .A(n11165), .ZN(n12156) );
  NAND2_X1 U11463 ( .A1(n11019), .A2(n12162), .ZN(n9045) );
  NAND2_X1 U11464 ( .A1(n9045), .A2(n12165), .ZN(n11152) );
  XNOR2_X1 U11465 ( .A(n12279), .B(n14529), .ZN(n12182) );
  OR2_X1 U11466 ( .A1(n12279), .A2(n14529), .ZN(n12173) );
  NAND2_X1 U11467 ( .A1(n11387), .A2(n12099), .ZN(n9047) );
  NAND2_X1 U11468 ( .A1(n9047), .A2(n12184), .ZN(n14503) );
  INV_X1 U11469 ( .A(n12189), .ZN(n9048) );
  INV_X1 U11470 ( .A(n12193), .ZN(n9049) );
  INV_X1 U11471 ( .A(n12624), .ZN(n12630) );
  INV_X1 U11472 ( .A(n12608), .ZN(n12614) );
  NAND2_X1 U11473 ( .A1(n12600), .A2(n12599), .ZN(n9050) );
  INV_X1 U11474 ( .A(n12219), .ZN(n9051) );
  OR2_X1 U11475 ( .A1(n12223), .A2(n12222), .ZN(n12224) );
  NAND2_X1 U11476 ( .A1(n9052), .A2(n12229), .ZN(n12535) );
  NAND2_X1 U11477 ( .A1(n12037), .A2(n11928), .ZN(n12234) );
  OR2_X1 U11478 ( .A1(n12676), .A2(n11946), .ZN(n12111) );
  NAND2_X1 U11479 ( .A1(n12676), .A2(n11946), .ZN(n12113) );
  NAND2_X1 U11480 ( .A1(n9054), .A2(n12113), .ZN(n12500) );
  INV_X1 U11481 ( .A(n12493), .ZN(n12499) );
  NAND2_X1 U11482 ( .A1(n12500), .A2(n12499), .ZN(n12498) );
  NAND2_X1 U11483 ( .A1(n12240), .A2(n12484), .ZN(n9055) );
  NAND2_X1 U11484 ( .A1(n12485), .A2(n12245), .ZN(n9057) );
  NAND2_X1 U11485 ( .A1(n9056), .A2(n12497), .ZN(n12246) );
  NAND2_X1 U11486 ( .A1(n9057), .A2(n12246), .ZN(n12468) );
  INV_X1 U11487 ( .A(n12471), .ZN(n12248) );
  AND2_X1 U11488 ( .A1(n12477), .A2(n12483), .ZN(n12252) );
  AOI21_X1 U11489 ( .B1(n12468), .B2(n12248), .A(n12252), .ZN(n12462) );
  INV_X1 U11490 ( .A(n12255), .ZN(n9058) );
  AOI21_X1 U11491 ( .B1(n12462), .B2(n12254), .A(n9058), .ZN(n12078) );
  NAND2_X1 U11492 ( .A1(n10441), .A2(n10181), .ZN(n9117) );
  INV_X1 U11493 ( .A(n9117), .ZN(n9060) );
  XNOR2_X1 U11494 ( .A(n9060), .B(n14437), .ZN(n9062) );
  NAND2_X1 U11495 ( .A1(n10441), .A2(n12428), .ZN(n9061) );
  NAND2_X1 U11496 ( .A1(n9062), .A2(n9061), .ZN(n10201) );
  NAND2_X1 U11497 ( .A1(n10181), .A2(n12428), .ZN(n9119) );
  INV_X1 U11498 ( .A(n9119), .ZN(n12267) );
  AND2_X1 U11499 ( .A1(n15138), .A2(n12267), .ZN(n9063) );
  NAND2_X1 U11500 ( .A1(n10201), .A2(n9063), .ZN(n9065) );
  NAND2_X1 U11501 ( .A1(n10193), .A2(n12428), .ZN(n9064) );
  OR2_X1 U11502 ( .A1(n14437), .A2(n9064), .ZN(n9116) );
  NAND2_X1 U11503 ( .A1(n14437), .A2(n15140), .ZN(n12663) );
  NAND2_X1 U11504 ( .A1(n11867), .A2(n9068), .ZN(n9124) );
  INV_X1 U11505 ( .A(n9100), .ZN(n9070) );
  INV_X1 U11506 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9069) );
  XNOR2_X2 U11507 ( .A(n9072), .B(n9071), .ZN(n9084) );
  XNOR2_X1 U11508 ( .A(n9084), .B(P3_B_REG_SCAN_IN), .ZN(n9076) );
  NAND2_X1 U11509 ( .A1(n9076), .A2(n11002), .ZN(n9081) );
  NAND2_X1 U11510 ( .A1(n9077), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9078) );
  MUX2_X1 U11511 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9078), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n9080) );
  INV_X1 U11512 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n15298) );
  NAND2_X1 U11513 ( .A1(n9784), .A2(n15298), .ZN(n9083) );
  NAND2_X1 U11514 ( .A1(n11002), .A2(n11151), .ZN(n9082) );
  NAND2_X1 U11515 ( .A1(n9084), .A2(n11151), .ZN(n9908) );
  NOR2_X1 U11516 ( .A1(P3_D_REG_5__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .ZN(
        n9089) );
  NOR4_X1 U11517 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_22__SCAN_IN), .ZN(n9088) );
  NOR4_X1 U11518 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n9087) );
  NOR4_X1 U11519 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n9086) );
  NAND4_X1 U11520 ( .A1(n9089), .A2(n9088), .A3(n9087), .A4(n9086), .ZN(n9095)
         );
  NOR4_X1 U11521 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n9093) );
  NOR4_X1 U11522 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_31__SCAN_IN), .A3(
        P3_D_REG_14__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n9092) );
  NOR4_X1 U11523 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9091) );
  NOR4_X1 U11524 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n9090) );
  NAND4_X1 U11525 ( .A1(n9093), .A2(n9092), .A3(n9091), .A4(n9090), .ZN(n9094)
         );
  OAI21_X1 U11526 ( .B1(n9095), .B2(n9094), .A(n9784), .ZN(n9112) );
  INV_X1 U11527 ( .A(n9112), .ZN(n9104) );
  INV_X1 U11528 ( .A(n9084), .ZN(n9097) );
  INV_X1 U11529 ( .A(n11002), .ZN(n9098) );
  NOR2_X1 U11530 ( .A1(n12244), .A2(n9119), .ZN(n10258) );
  NAND2_X1 U11531 ( .A1(n10392), .A2(n10258), .ZN(n10207) );
  NAND2_X1 U11532 ( .A1(n10441), .A2(n10193), .ZN(n12108) );
  NOR2_X1 U11533 ( .A1(n9120), .A2(n12108), .ZN(n10202) );
  NAND2_X1 U11534 ( .A1(n10392), .A2(n10202), .ZN(n9102) );
  NAND2_X1 U11535 ( .A1(n10207), .A2(n9102), .ZN(n9103) );
  NAND2_X1 U11536 ( .A1(n10212), .A2(n9103), .ZN(n9106) );
  NAND2_X1 U11537 ( .A1(n10261), .A2(n10195), .ZN(n9114) );
  NAND3_X1 U11538 ( .A1(n10208), .A2(n10392), .A3(n10201), .ZN(n9105) );
  INV_X1 U11539 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9107) );
  NOR2_X1 U11540 ( .A1(n15206), .A2(n9107), .ZN(n9109) );
  INV_X1 U11541 ( .A(n11866), .ZN(n9125) );
  NOR2_X1 U11542 ( .A1(n9125), .A2(n12776), .ZN(n9108) );
  NAND2_X1 U11543 ( .A1(n9111), .A2(n9110), .ZN(P3_U3456) );
  AND2_X1 U11544 ( .A1(n9112), .A2(n10392), .ZN(n9113) );
  NAND2_X1 U11545 ( .A1(n12260), .A2(n9119), .ZN(n10185) );
  NAND2_X1 U11546 ( .A1(n12244), .A2(n9116), .ZN(n10260) );
  AND2_X1 U11547 ( .A1(n10185), .A2(n10260), .ZN(n10262) );
  NAND2_X1 U11548 ( .A1(n14437), .A2(n9117), .ZN(n9118) );
  NAND3_X1 U11549 ( .A1(n9120), .A2(n9119), .A3(n9118), .ZN(n9121) );
  AND2_X1 U11550 ( .A1(n9121), .A2(n12244), .ZN(n9122) );
  MUX2_X1 U11551 ( .A(n10262), .B(n9122), .S(n10261), .Z(n9123) );
  NAND2_X1 U11552 ( .A1(n9124), .A2(n15222), .ZN(n9128) );
  NOR2_X1 U11553 ( .A1(n9125), .A2(n12722), .ZN(n9126) );
  NOR2_X1 U11554 ( .A1(n7638), .A2(n9126), .ZN(n9127) );
  NAND2_X1 U11555 ( .A1(n9128), .A2(n9127), .ZN(P3_U3488) );
  NOR2_X2 U11556 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9158) );
  NAND4_X1 U11557 ( .A1(n9132), .A2(n9131), .A3(n9130), .A4(n9286), .ZN(n9134)
         );
  NOR2_X1 U11558 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n9139) );
  NOR2_X1 U11559 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n9138) );
  NOR2_X1 U11560 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), 
        .ZN(n9137) );
  NOR2_X1 U11561 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n9136) );
  INV_X1 U11562 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9141) );
  NAND2_X2 U11563 ( .A1(n9148), .A2(n14302), .ZN(n13506) );
  INV_X1 U11564 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9145) );
  NAND2_X1 U11565 ( .A1(n13503), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9146) );
  NAND2_X4 U11566 ( .A1(n9150), .A2(n14302), .ZN(n13505) );
  INV_X1 U11567 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9810) );
  NAND2_X1 U11568 ( .A1(n9150), .A2(n9149), .ZN(n9211) );
  INV_X1 U11569 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9151) );
  OR2_X1 U11570 ( .A1(n9211), .A2(n9151), .ZN(n9152) );
  OR2_X1 U11571 ( .A1(n13514), .A2(n7653), .ZN(n9164) );
  NAND2_X2 U11572 ( .A1(n9429), .A2(n9155), .ZN(n9272) );
  OR2_X1 U11573 ( .A1(n9272), .A2(n9654), .ZN(n9163) );
  NAND2_X1 U11574 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9157) );
  MUX2_X1 U11575 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9157), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9161) );
  INV_X1 U11576 ( .A(n9159), .ZN(n9160) );
  NAND2_X1 U11577 ( .A1(n9161), .A2(n9160), .ZN(n9812) );
  OR2_X1 U11578 ( .A1(n9429), .A2(n9812), .ZN(n9162) );
  NAND2_X1 U11579 ( .A1(n9981), .A2(n14751), .ZN(n9526) );
  INV_X1 U11580 ( .A(n9526), .ZN(n13566) );
  NAND2_X1 U11581 ( .A1(n13503), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9170) );
  INV_X1 U11582 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10639) );
  OR2_X1 U11583 ( .A1(n9211), .A2(n10639), .ZN(n9169) );
  INV_X1 U11584 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9165) );
  INV_X1 U11585 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9166) );
  OR2_X1 U11586 ( .A1(n13505), .A2(n9166), .ZN(n9167) );
  NOR2_X1 U11587 ( .A1(n7171), .A2(n9640), .ZN(n9172) );
  XNOR2_X1 U11588 ( .A(n9172), .B(n9171), .ZN(n14322) );
  OAI21_X1 U11589 ( .B1(n13566), .B2(n13565), .A(n13562), .ZN(n10577) );
  NAND2_X1 U11590 ( .A1(n13503), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9179) );
  INV_X1 U11591 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9174) );
  OR2_X1 U11592 ( .A1(n9211), .A2(n9174), .ZN(n9178) );
  INV_X1 U11593 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9175) );
  OR2_X1 U11594 ( .A1(n13506), .A2(n9175), .ZN(n9177) );
  INV_X1 U11595 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9809) );
  NOR2_X1 U11596 ( .A1(n9159), .A2(n9156), .ZN(n9180) );
  MUX2_X1 U11597 ( .A(n9156), .B(n9180), .S(P1_IR_REG_2__SCAN_IN), .Z(n9181)
         );
  INV_X1 U11598 ( .A(n9181), .ZN(n9183) );
  INV_X1 U11599 ( .A(n9189), .ZN(n9182) );
  NAND2_X1 U11600 ( .A1(n9183), .A2(n9182), .ZN(n13819) );
  NAND2_X1 U11601 ( .A1(n13798), .A2(n10058), .ZN(n13572) );
  NAND2_X1 U11602 ( .A1(n10577), .A2(n13569), .ZN(n10576) );
  NAND2_X1 U11603 ( .A1(n10576), .A2(n13573), .ZN(n10225) );
  INV_X1 U11604 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9813) );
  OR2_X1 U11605 ( .A1(n13505), .A2(n9813), .ZN(n9187) );
  INV_X1 U11606 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9184) );
  OR2_X1 U11607 ( .A1(n13506), .A2(n9184), .ZN(n9186) );
  OR2_X1 U11608 ( .A1(n9211), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9185) );
  NAND4_X1 U11609 ( .A1(n9188), .A2(n9187), .A3(n9186), .A4(n9185), .ZN(n13797) );
  OR2_X1 U11610 ( .A1(n13514), .A2(n9630), .ZN(n9193) );
  OR2_X1 U11611 ( .A1(n9189), .A2(n9156), .ZN(n9191) );
  XNOR2_X1 U11612 ( .A(n9191), .B(n9190), .ZN(n13834) );
  OR2_X1 U11613 ( .A1(n9429), .A2(n13834), .ZN(n9192) );
  INV_X1 U11614 ( .A(n10222), .ZN(n13576) );
  OR2_X1 U11615 ( .A1(n13797), .A2(n13578), .ZN(n13579) );
  NAND2_X1 U11616 ( .A1(n10224), .A2(n13579), .ZN(n10489) );
  NAND2_X1 U11617 ( .A1(n13503), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9198) );
  INV_X1 U11618 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9194) );
  OR2_X1 U11619 ( .A1(n13506), .A2(n9194), .ZN(n9197) );
  NAND2_X1 U11620 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9213) );
  OAI21_X1 U11621 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n9213), .ZN(n10497) );
  OR2_X1 U11622 ( .A1(n9211), .A2(n10497), .ZN(n9196) );
  INV_X1 U11623 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9808) );
  OR2_X1 U11624 ( .A1(n13505), .A2(n9808), .ZN(n9195) );
  NAND4_X1 U11625 ( .A1(n9198), .A2(n9197), .A3(n9196), .A4(n9195), .ZN(n13796) );
  NAND2_X1 U11626 ( .A1(n9636), .A2(n13511), .ZN(n9205) );
  NOR2_X1 U11627 ( .A1(n9201), .A2(n9156), .ZN(n9199) );
  MUX2_X1 U11628 ( .A(n9156), .B(n9199), .S(P1_IR_REG_4__SCAN_IN), .Z(n9203)
         );
  INV_X1 U11629 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9200) );
  NAND2_X1 U11630 ( .A1(n9201), .A2(n9200), .ZN(n9341) );
  INV_X1 U11631 ( .A(n9341), .ZN(n9202) );
  NOR2_X1 U11632 ( .A1(n9203), .A2(n9202), .ZN(n14633) );
  AOI22_X1 U11633 ( .A1(n9399), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9799), .B2(
        n14633), .ZN(n9204) );
  XNOR2_X1 U11634 ( .A(n13796), .B(n10507), .ZN(n13519) );
  NAND2_X1 U11635 ( .A1(n13796), .A2(n10507), .ZN(n9206) );
  NAND2_X1 U11636 ( .A1(n9641), .A2(n13511), .ZN(n9210) );
  NAND2_X1 U11637 ( .A1(n9341), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9207) );
  MUX2_X1 U11638 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9207), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n9208) );
  AND2_X1 U11639 ( .A1(n9208), .A2(n9232), .ZN(n9819) );
  AOI22_X1 U11640 ( .A1(n9399), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9799), .B2(
        n9819), .ZN(n9209) );
  NAND2_X1 U11641 ( .A1(n9210), .A2(n9209), .ZN(n13590) );
  NAND2_X1 U11642 ( .A1(n9512), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9219) );
  INV_X1 U11643 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9828) );
  OR2_X1 U11644 ( .A1(n9560), .A2(n9828), .ZN(n9218) );
  AND2_X1 U11645 ( .A1(n9213), .A2(n9212), .ZN(n9214) );
  NOR2_X1 U11646 ( .A1(n9213), .A2(n9212), .ZN(n9224) );
  OR2_X1 U11647 ( .A1(n9214), .A2(n9224), .ZN(n10592) );
  OR2_X1 U11648 ( .A1(n9513), .A2(n10592), .ZN(n9217) );
  INV_X1 U11649 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9215) );
  OR2_X1 U11650 ( .A1(n9562), .A2(n9215), .ZN(n9216) );
  NAND4_X1 U11651 ( .A1(n9219), .A2(n9218), .A3(n9217), .A4(n9216), .ZN(n13795) );
  NOR2_X1 U11652 ( .A1(n13590), .A2(n10588), .ZN(n9220) );
  NAND2_X1 U11653 ( .A1(n9665), .A2(n13511), .ZN(n9223) );
  NAND2_X1 U11654 ( .A1(n9232), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9221) );
  XNOR2_X1 U11655 ( .A(n9221), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9837) );
  AOI22_X1 U11656 ( .A1(n9399), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9799), .B2(
        n9837), .ZN(n9222) );
  NAND2_X1 U11657 ( .A1(n9223), .A2(n9222), .ZN(n13594) );
  NAND2_X1 U11658 ( .A1(n13503), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9230) );
  INV_X1 U11659 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9836) );
  OR2_X1 U11660 ( .A1(n13505), .A2(n9836), .ZN(n9229) );
  NAND2_X1 U11661 ( .A1(n9224), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9236) );
  OR2_X1 U11662 ( .A1(n9224), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9225) );
  NAND2_X1 U11663 ( .A1(n9236), .A2(n9225), .ZN(n14707) );
  OR2_X1 U11664 ( .A1(n9513), .A2(n14707), .ZN(n9228) );
  INV_X1 U11665 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9226) );
  OR2_X1 U11666 ( .A1(n13506), .A2(n9226), .ZN(n9227) );
  XNOR2_X1 U11667 ( .A(n13594), .B(n13593), .ZN(n14701) );
  INV_X1 U11668 ( .A(n14701), .ZN(n13522) );
  AND2_X1 U11669 ( .A1(n13594), .A2(n13593), .ZN(n9231) );
  NOR2_X1 U11670 ( .A1(n9232), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n9245) );
  OR2_X1 U11671 ( .A1(n9245), .A2(n9156), .ZN(n9233) );
  XNOR2_X1 U11672 ( .A(n9233), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9838) );
  AOI22_X1 U11673 ( .A1(n9399), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9799), .B2(
        n9838), .ZN(n9234) );
  NAND2_X1 U11674 ( .A1(n9235), .A2(n9234), .ZN(n13603) );
  NAND2_X1 U11675 ( .A1(n9512), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9242) );
  INV_X1 U11676 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9829) );
  OR2_X1 U11677 ( .A1(n9560), .A2(n9829), .ZN(n9241) );
  NAND2_X1 U11678 ( .A1(n9236), .A2(n10749), .ZN(n9237) );
  NAND2_X1 U11679 ( .A1(n9249), .A2(n9237), .ZN(n10764) );
  OR2_X1 U11680 ( .A1(n9513), .A2(n10764), .ZN(n9240) );
  INV_X1 U11681 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9238) );
  OR2_X1 U11682 ( .A1(n9562), .A2(n9238), .ZN(n9239) );
  XNOR2_X1 U11683 ( .A(n13603), .B(n10791), .ZN(n9534) );
  NAND2_X1 U11684 ( .A1(n10759), .A2(n13523), .ZN(n10758) );
  INV_X1 U11685 ( .A(n10791), .ZN(n13793) );
  NAND2_X1 U11686 ( .A1(n10765), .A2(n13793), .ZN(n9243) );
  NAND2_X1 U11687 ( .A1(n10758), .A2(n9243), .ZN(n10790) );
  OR2_X1 U11688 ( .A1(n9678), .A2(n9272), .ZN(n9248) );
  NAND2_X1 U11689 ( .A1(n9245), .A2(n9244), .ZN(n9257) );
  NAND2_X1 U11690 ( .A1(n9257), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9246) );
  XNOR2_X1 U11691 ( .A(n9246), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9856) );
  AOI22_X1 U11692 ( .A1(n9399), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9799), .B2(
        n9856), .ZN(n9247) );
  NAND2_X1 U11693 ( .A1(n9248), .A2(n9247), .ZN(n13607) );
  NAND2_X1 U11694 ( .A1(n9512), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9255) );
  INV_X1 U11695 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9850) );
  OR2_X1 U11696 ( .A1(n9560), .A2(n9850), .ZN(n9254) );
  NAND2_X1 U11697 ( .A1(n9249), .A2(n10850), .ZN(n9250) );
  NAND2_X1 U11698 ( .A1(n9262), .A2(n9250), .ZN(n10796) );
  OR2_X1 U11699 ( .A1(n9513), .A2(n10796), .ZN(n9253) );
  INV_X1 U11700 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9251) );
  OR2_X1 U11701 ( .A1(n13506), .A2(n9251), .ZN(n9252) );
  NAND4_X1 U11702 ( .A1(n9255), .A2(n9254), .A3(n9253), .A4(n9252), .ZN(n13792) );
  XNOR2_X1 U11703 ( .A(n13607), .B(n13792), .ZN(n13525) );
  NAND2_X1 U11704 ( .A1(n10790), .A2(n13525), .ZN(n10789) );
  INV_X1 U11705 ( .A(n13607), .ZN(n14797) );
  NAND2_X1 U11706 ( .A1(n14797), .A2(n13792), .ZN(n9256) );
  OR2_X1 U11707 ( .A1(n9683), .A2(n9272), .ZN(n9261) );
  NAND2_X1 U11708 ( .A1(n9288), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9258) );
  OR2_X1 U11709 ( .A1(n9258), .A2(n9286), .ZN(n9259) );
  NAND2_X1 U11710 ( .A1(n9258), .A2(n9286), .ZN(n9273) );
  AOI22_X1 U11711 ( .A1(n9399), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9799), .B2(
        n9857), .ZN(n9260) );
  NAND2_X1 U11712 ( .A1(n9419), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9268) );
  INV_X1 U11713 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n14690) );
  OR2_X1 U11714 ( .A1(n13505), .A2(n14690), .ZN(n9267) );
  INV_X1 U11715 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10139) );
  OR2_X1 U11716 ( .A1(n9560), .A2(n10139), .ZN(n9266) );
  INV_X1 U11717 ( .A(n9277), .ZN(n9264) );
  NAND2_X1 U11718 ( .A1(n9262), .A2(n15259), .ZN(n9263) );
  NAND2_X1 U11719 ( .A1(n9264), .A2(n9263), .ZN(n14689) );
  OR2_X1 U11720 ( .A1(n9513), .A2(n14689), .ZN(n9265) );
  NAND4_X1 U11721 ( .A1(n9268), .A2(n9267), .A3(n9266), .A4(n9265), .ZN(n13791) );
  XNOR2_X1 U11722 ( .A(n14693), .B(n13791), .ZN(n13527) );
  INV_X1 U11723 ( .A(n13527), .ZN(n14681) );
  INV_X1 U11724 ( .A(n13791), .ZN(n9269) );
  NAND2_X1 U11725 ( .A1(n14693), .A2(n9269), .ZN(n9270) );
  OR2_X1 U11726 ( .A1(n9271), .A2(n9272), .ZN(n9276) );
  NAND2_X1 U11727 ( .A1(n9273), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9274) );
  XNOR2_X1 U11728 ( .A(n9274), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10148) );
  AOI22_X1 U11729 ( .A1(n9399), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n9799), 
        .B2(n10148), .ZN(n9275) );
  NAND2_X1 U11730 ( .A1(n13503), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9283) );
  INV_X1 U11731 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10147) );
  OR2_X1 U11732 ( .A1(n13505), .A2(n10147), .ZN(n9282) );
  NAND2_X1 U11733 ( .A1(n9277), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9293) );
  OR2_X1 U11734 ( .A1(n9277), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9278) );
  NAND2_X1 U11735 ( .A1(n9293), .A2(n9278), .ZN(n11056) );
  OR2_X1 U11736 ( .A1(n9513), .A2(n11056), .ZN(n9281) );
  INV_X1 U11737 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9279) );
  OR2_X1 U11738 ( .A1(n9562), .A2(n9279), .ZN(n9280) );
  XNOR2_X1 U11739 ( .A(n13618), .B(n11344), .ZN(n13529) );
  OR2_X1 U11740 ( .A1(n13618), .A2(n11344), .ZN(n9284) );
  NAND2_X1 U11741 ( .A1(n9929), .A2(n13511), .ZN(n9291) );
  NAND2_X1 U11742 ( .A1(n9286), .A2(n9285), .ZN(n9287) );
  NAND2_X1 U11743 ( .A1(n9302), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9289) );
  XNOR2_X1 U11744 ( .A(n9289), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10728) );
  AOI22_X1 U11745 ( .A1(n9399), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9799), 
        .B2(n10728), .ZN(n9290) );
  NAND2_X1 U11746 ( .A1(n9419), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9300) );
  NAND2_X1 U11747 ( .A1(n9293), .A2(n9292), .ZN(n9294) );
  NAND2_X1 U11748 ( .A1(n9320), .A2(n9294), .ZN(n14571) );
  OR2_X1 U11749 ( .A1(n9513), .A2(n14571), .ZN(n9299) );
  INV_X1 U11750 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9295) );
  OR2_X1 U11751 ( .A1(n9560), .A2(n9295), .ZN(n9298) );
  INV_X1 U11752 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9296) );
  OR2_X1 U11753 ( .A1(n13505), .A2(n9296), .ZN(n9297) );
  XNOR2_X1 U11754 ( .A(n14563), .B(n11471), .ZN(n13530) );
  NAND2_X1 U11755 ( .A1(n11342), .A2(n7406), .ZN(n11347) );
  OR2_X1 U11756 ( .A1(n14563), .A2(n11471), .ZN(n9301) );
  NAND2_X1 U11757 ( .A1(n11347), .A2(n9301), .ZN(n11318) );
  NAND2_X1 U11758 ( .A1(n9999), .A2(n13511), .ZN(n9304) );
  OAI21_X1 U11759 ( .B1(n9302), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9313) );
  XNOR2_X1 U11760 ( .A(n9313), .B(P1_IR_REG_12__SCAN_IN), .ZN(n14655) );
  AOI22_X1 U11761 ( .A1(n9399), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n14655), 
        .B2(n9799), .ZN(n9303) );
  NAND2_X2 U11762 ( .A1(n9304), .A2(n9303), .ZN(n14553) );
  NAND2_X1 U11763 ( .A1(n13503), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9310) );
  INV_X1 U11764 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11326) );
  OR2_X1 U11765 ( .A1(n13505), .A2(n11326), .ZN(n9309) );
  INV_X1 U11766 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9305) );
  OR2_X1 U11767 ( .A1(n9562), .A2(n9305), .ZN(n9308) );
  INV_X1 U11768 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9306) );
  XNOR2_X1 U11769 ( .A(n9320), .B(n9306), .ZN(n14557) );
  OR2_X1 U11770 ( .A1(n9513), .A2(n14557), .ZN(n9307) );
  XNOR2_X1 U11771 ( .A(n14553), .B(n11486), .ZN(n13532) );
  NAND2_X1 U11772 ( .A1(n11318), .A2(n7409), .ZN(n11317) );
  OR2_X1 U11773 ( .A1(n14553), .A2(n11486), .ZN(n9311) );
  NAND2_X1 U11774 ( .A1(n10076), .A2(n13511), .ZN(n9316) );
  INV_X1 U11775 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9312) );
  NAND2_X1 U11776 ( .A1(n9313), .A2(n9312), .ZN(n9314) );
  NAND2_X1 U11777 ( .A1(n9314), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9329) );
  XNOR2_X1 U11778 ( .A(n9329), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11266) );
  AOI22_X1 U11779 ( .A1(n11266), .A2(n9799), .B1(n9399), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n9315) );
  NAND2_X1 U11780 ( .A1(n13503), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9326) );
  INV_X1 U11781 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9317) );
  OR2_X1 U11782 ( .A1(n13505), .A2(n9317), .ZN(n9325) );
  INV_X1 U11783 ( .A(n9320), .ZN(n9318) );
  AOI21_X1 U11784 ( .B1(n9318), .B2(P1_REG3_REG_12__SCAN_IN), .A(
        P1_REG3_REG_13__SCAN_IN), .ZN(n9321) );
  NAND2_X1 U11785 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n9319) );
  OR2_X1 U11786 ( .A1(n9321), .A2(n9335), .ZN(n14452) );
  OR2_X1 U11787 ( .A1(n9513), .A2(n14452), .ZN(n9324) );
  INV_X1 U11788 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9322) );
  OR2_X1 U11789 ( .A1(n9562), .A2(n9322), .ZN(n9323) );
  XNOR2_X1 U11790 ( .A(n13638), .B(n13636), .ZN(n14456) );
  INV_X1 U11791 ( .A(n14456), .ZN(n14448) );
  NAND2_X1 U11792 ( .A1(n14449), .A2(n14448), .ZN(n14447) );
  OR2_X1 U11793 ( .A1(n13638), .A2(n13636), .ZN(n9327) );
  NAND2_X1 U11794 ( .A1(n10389), .A2(n13511), .ZN(n9333) );
  INV_X1 U11795 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9328) );
  NAND2_X1 U11796 ( .A1(n9329), .A2(n9328), .ZN(n9330) );
  NAND2_X1 U11797 ( .A1(n9330), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9331) );
  AOI22_X1 U11798 ( .A1(n13894), .A2(n9799), .B1(n9399), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9332) );
  NAND2_X1 U11799 ( .A1(n9419), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9340) );
  INV_X1 U11800 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11257) );
  OR2_X1 U11801 ( .A1(n9560), .A2(n11257), .ZN(n9339) );
  INV_X1 U11802 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9334) );
  OR2_X1 U11803 ( .A1(n13505), .A2(n9334), .ZN(n9338) );
  NAND2_X1 U11804 ( .A1(n9335), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9346) );
  OR2_X1 U11805 ( .A1(n9335), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9336) );
  NAND2_X1 U11806 ( .A1(n9346), .A2(n9336), .ZN(n15384) );
  OR2_X1 U11807 ( .A1(n9513), .A2(n15384), .ZN(n9337) );
  NAND4_X1 U11808 ( .A1(n9340), .A2(n9339), .A3(n9338), .A4(n9337), .ZN(n13786) );
  NAND2_X1 U11809 ( .A1(n15383), .A2(n13786), .ZN(n13647) );
  INV_X1 U11810 ( .A(n13786), .ZN(n11744) );
  NAND2_X1 U11811 ( .A1(n11506), .A2(n11744), .ZN(n13645) );
  NAND2_X1 U11812 ( .A1(n10753), .A2(n13511), .ZN(n9344) );
  OR2_X1 U11813 ( .A1(n9341), .A2(n6583), .ZN(n9352) );
  NAND2_X1 U11814 ( .A1(n9352), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9342) );
  XNOR2_X1 U11815 ( .A(n9342), .B(P1_IR_REG_15__SCAN_IN), .ZN(n14668) );
  AOI22_X1 U11816 ( .A1(n9399), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9799), 
        .B2(n14668), .ZN(n9343) );
  NAND2_X1 U11817 ( .A1(n9419), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n9351) );
  INV_X1 U11818 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11519) );
  OR2_X1 U11819 ( .A1(n13505), .A2(n11519), .ZN(n9350) );
  INV_X1 U11820 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14664) );
  OR2_X1 U11821 ( .A1(n9560), .A2(n14664), .ZN(n9349) );
  INV_X1 U11822 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9345) );
  NAND2_X1 U11823 ( .A1(n9346), .A2(n9345), .ZN(n9347) );
  NAND2_X1 U11824 ( .A1(n9357), .A2(n9347), .ZN(n13497) );
  OR2_X1 U11825 ( .A1(n9513), .A2(n13497), .ZN(n9348) );
  NAND2_X1 U11826 ( .A1(n14248), .A2(n11752), .ZN(n13652) );
  NAND2_X1 U11827 ( .A1(n10802), .A2(n13511), .ZN(n9355) );
  OAI21_X1 U11828 ( .B1(n9352), .B2(P1_IR_REG_15__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9353) );
  XNOR2_X1 U11829 ( .A(n9353), .B(P1_IR_REG_16__SCAN_IN), .ZN(n11456) );
  AOI22_X1 U11830 ( .A1(n9399), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9799), 
        .B2(n11456), .ZN(n9354) );
  INV_X1 U11831 ( .A(n9513), .ZN(n9359) );
  INV_X1 U11832 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9356) );
  AND2_X1 U11833 ( .A1(n9357), .A2(n9356), .ZN(n9358) );
  NOR2_X1 U11834 ( .A1(n9370), .A2(n9358), .ZN(n13432) );
  NAND2_X1 U11835 ( .A1(n9359), .A2(n13432), .ZN(n9365) );
  INV_X1 U11836 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11536) );
  OR2_X1 U11837 ( .A1(n13505), .A2(n11536), .ZN(n9364) );
  INV_X1 U11838 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9360) );
  OR2_X1 U11839 ( .A1(n9560), .A2(n9360), .ZN(n9363) );
  INV_X1 U11840 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9361) );
  OR2_X1 U11841 ( .A1(n9562), .A2(n9361), .ZN(n9362) );
  XNOR2_X1 U11842 ( .A(n13657), .B(n13656), .ZN(n13535) );
  NAND2_X1 U11843 ( .A1(n13657), .A2(n13656), .ZN(n9366) );
  NAND2_X1 U11844 ( .A1(n10818), .A2(n13511), .ZN(n9369) );
  NAND2_X1 U11845 ( .A1(n9379), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9367) );
  XNOR2_X1 U11846 ( .A(n9367), .B(P1_IR_REG_17__SCAN_IN), .ZN(n13906) );
  AOI22_X1 U11847 ( .A1(n9399), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9799), 
        .B2(n13906), .ZN(n9368) );
  NOR2_X1 U11848 ( .A1(n9370), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9371) );
  OR2_X1 U11849 ( .A1(n9387), .A2(n9371), .ZN(n14140) );
  NAND2_X1 U11850 ( .A1(n9419), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9372) );
  OAI21_X1 U11851 ( .B1(n14140), .B2(n9513), .A(n9372), .ZN(n9376) );
  INV_X1 U11852 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9374) );
  INV_X1 U11853 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14144) );
  OR2_X1 U11854 ( .A1(n13505), .A2(n14144), .ZN(n9373) );
  OAI21_X1 U11855 ( .B1(n9560), .B2(n9374), .A(n9373), .ZN(n9375) );
  INV_X1 U11856 ( .A(n13783), .ZN(n9378) );
  AND2_X1 U11857 ( .A1(n14235), .A2(n9378), .ZN(n9377) );
  NAND2_X1 U11858 ( .A1(n11033), .A2(n13511), .ZN(n9386) );
  INV_X1 U11859 ( .A(n9383), .ZN(n9380) );
  NAND2_X1 U11860 ( .A1(n9380), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9381) );
  MUX2_X1 U11861 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9381), .S(
        P1_IR_REG_18__SCAN_IN), .Z(n9384) );
  NAND2_X1 U11862 ( .A1(n9384), .A2(n9397), .ZN(n13914) );
  INV_X1 U11863 ( .A(n13914), .ZN(n13920) );
  AOI22_X1 U11864 ( .A1(n9399), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9799), 
        .B2(n13920), .ZN(n9385) );
  OR2_X1 U11865 ( .A1(n9387), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9388) );
  NAND2_X1 U11866 ( .A1(n9402), .A2(n9388), .ZN(n13477) );
  NAND2_X1 U11867 ( .A1(n9419), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n9389) );
  OAI21_X1 U11868 ( .B1(n13477), .B2(n9513), .A(n9389), .ZN(n9392) );
  INV_X1 U11869 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n13908) );
  INV_X1 U11870 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9390) );
  OAI22_X1 U11871 ( .A1(n9560), .A2(n13908), .B1(n13505), .B2(n9390), .ZN(
        n9391) );
  OR2_X1 U11872 ( .A1(n14230), .A2(n13672), .ZN(n9394) );
  NAND2_X1 U11873 ( .A1(n14230), .A2(n13672), .ZN(n9393) );
  NAND2_X1 U11874 ( .A1(n14123), .A2(n14122), .ZN(n9395) );
  NAND2_X1 U11875 ( .A1(n11124), .A2(n13511), .ZN(n9401) );
  NAND2_X1 U11876 ( .A1(n9397), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9396) );
  MUX2_X1 U11877 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9396), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n9398) );
  AOI22_X1 U11878 ( .A1(n9399), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14082), 
        .B2(n9799), .ZN(n9400) );
  INV_X1 U11879 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9406) );
  INV_X1 U11880 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n13405) );
  NAND2_X1 U11881 ( .A1(n9402), .A2(n13405), .ZN(n9403) );
  NAND2_X1 U11882 ( .A1(n9409), .A2(n9403), .ZN(n14112) );
  OR2_X1 U11883 ( .A1(n14112), .A2(n9513), .ZN(n9405) );
  AOI22_X1 U11884 ( .A1(n13503), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n9512), 
        .B2(P1_REG2_REG_19__SCAN_IN), .ZN(n9404) );
  OAI211_X1 U11885 ( .C1(n9562), .C2(n9406), .A(n9405), .B(n9404), .ZN(n13781)
         );
  XNOR2_X1 U11886 ( .A(n14290), .B(n13781), .ZN(n14105) );
  INV_X1 U11887 ( .A(n13781), .ZN(n13669) );
  NAND2_X1 U11888 ( .A1(n14290), .A2(n13669), .ZN(n13680) );
  NAND2_X1 U11889 ( .A1(n11371), .A2(n13511), .ZN(n9408) );
  OR2_X1 U11890 ( .A1(n13514), .A2(n11375), .ZN(n9407) );
  INV_X1 U11891 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13459) );
  AND2_X1 U11892 ( .A1(n9409), .A2(n13459), .ZN(n9410) );
  OR2_X1 U11893 ( .A1(n9417), .A2(n9410), .ZN(n13457) );
  AOI22_X1 U11894 ( .A1(n13503), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n9512), 
        .B2(P1_REG2_REG_20__SCAN_IN), .ZN(n9412) );
  NAND2_X1 U11895 ( .A1(n9419), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9411) );
  OAI211_X1 U11896 ( .C1(n13457), .C2(n9513), .A(n9412), .B(n9411), .ZN(n13780) );
  INV_X1 U11897 ( .A(n13780), .ZN(n13685) );
  OR2_X1 U11898 ( .A1(n14215), .A2(n13685), .ZN(n9414) );
  NAND2_X1 U11899 ( .A1(n14215), .A2(n13685), .ZN(n9413) );
  NAND2_X1 U11900 ( .A1(n11444), .A2(n13511), .ZN(n9416) );
  OR2_X1 U11901 ( .A1(n13514), .A2(n11448), .ZN(n9415) );
  OR2_X1 U11902 ( .A1(n9417), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9418) );
  NAND2_X1 U11903 ( .A1(n9417), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9431) );
  NAND2_X1 U11904 ( .A1(n9418), .A2(n9431), .ZN(n14084) );
  OR2_X1 U11905 ( .A1(n14084), .A2(n9513), .ZN(n9425) );
  INV_X1 U11906 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9422) );
  NAND2_X1 U11907 ( .A1(n9512), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9421) );
  NAND2_X1 U11908 ( .A1(n9419), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9420) );
  OAI211_X1 U11909 ( .C1(n9560), .C2(n9422), .A(n9421), .B(n9420), .ZN(n9423)
         );
  INV_X1 U11910 ( .A(n9423), .ZN(n9424) );
  NAND2_X1 U11911 ( .A1(n9425), .A2(n9424), .ZN(n13779) );
  INV_X1 U11912 ( .A(n13779), .ZN(n9426) );
  NOR2_X1 U11913 ( .A1(n14285), .A2(n9426), .ZN(n9427) );
  NAND2_X1 U11914 ( .A1(n13503), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n9437) );
  INV_X1 U11915 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9430) );
  OR2_X1 U11916 ( .A1(n13505), .A2(n9430), .ZN(n9436) );
  NAND2_X1 U11917 ( .A1(n9432), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9440) );
  OAI21_X1 U11918 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n9432), .A(n9440), .ZN(
        n14067) );
  OR2_X1 U11919 ( .A1(n9513), .A2(n14067), .ZN(n9435) );
  INV_X1 U11920 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9433) );
  OR2_X1 U11921 ( .A1(n13506), .A2(n9433), .ZN(n9434) );
  NAND4_X1 U11922 ( .A1(n9437), .A2(n9436), .A3(n9435), .A4(n9434), .ZN(n13778) );
  NAND2_X1 U11923 ( .A1(n14315), .A2(n13511), .ZN(n9439) );
  OR2_X1 U11924 ( .A1(n13514), .A2(n14319), .ZN(n9438) );
  NAND2_X1 U11925 ( .A1(n13503), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9444) );
  INV_X1 U11926 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n14275) );
  OR2_X1 U11927 ( .A1(n9562), .A2(n14275), .ZN(n9443) );
  XNOR2_X1 U11928 ( .A(P1_REG3_REG_23__SCAN_IN), .B(n9449), .ZN(n14050) );
  OR2_X1 U11929 ( .A1(n9513), .A2(n14050), .ZN(n9442) );
  INV_X1 U11930 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14051) );
  OR2_X1 U11931 ( .A1(n13505), .A2(n14051), .ZN(n9441) );
  NAND4_X1 U11932 ( .A1(n9444), .A2(n9443), .A3(n9442), .A4(n9441), .ZN(n13777) );
  INV_X1 U11933 ( .A(n13777), .ZN(n9445) );
  NAND2_X1 U11934 ( .A1(n14049), .A2(n9445), .ZN(n9446) );
  NAND2_X1 U11935 ( .A1(n11545), .A2(n13511), .ZN(n9448) );
  OR2_X1 U11936 ( .A1(n13514), .A2(n11547), .ZN(n9447) );
  NAND2_X1 U11937 ( .A1(n9512), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9454) );
  NAND3_X1 U11938 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(P1_REG3_REG_24__SCAN_IN), 
        .A3(n9449), .ZN(n9465) );
  INV_X1 U11939 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9451) );
  NAND2_X1 U11940 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n9449), .ZN(n9450) );
  NAND2_X1 U11941 ( .A1(n9451), .A2(n9450), .ZN(n9452) );
  NAND2_X1 U11942 ( .A1(n9465), .A2(n9452), .ZN(n14037) );
  OR2_X1 U11943 ( .A1(n9513), .A2(n14037), .ZN(n9453) );
  NAND2_X1 U11944 ( .A1(n9454), .A2(n9453), .ZN(n9459) );
  INV_X1 U11945 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9455) );
  NOR2_X1 U11946 ( .A1(n9560), .A2(n9455), .ZN(n9458) );
  INV_X1 U11947 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9456) );
  NOR2_X1 U11948 ( .A1(n9562), .A2(n9456), .ZN(n9457) );
  XNOR2_X1 U11949 ( .A(n14272), .B(n13776), .ZN(n14032) );
  INV_X1 U11950 ( .A(n14032), .ZN(n14024) );
  INV_X1 U11951 ( .A(n13776), .ZN(n13383) );
  OR2_X1 U11952 ( .A1(n13383), .A2(n14272), .ZN(n9460) );
  NAND2_X1 U11953 ( .A1(n13362), .A2(n13511), .ZN(n9462) );
  OR2_X1 U11954 ( .A1(n13514), .A2(n14313), .ZN(n9461) );
  NAND2_X1 U11955 ( .A1(n9512), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9471) );
  INV_X1 U11956 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9463) );
  OR2_X1 U11957 ( .A1(n9560), .A2(n9463), .ZN(n9470) );
  INV_X1 U11958 ( .A(n9465), .ZN(n9464) );
  NAND2_X1 U11959 ( .A1(n9464), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9478) );
  INV_X1 U11960 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n15244) );
  NAND2_X1 U11961 ( .A1(n9465), .A2(n15244), .ZN(n9466) );
  NAND2_X1 U11962 ( .A1(n9478), .A2(n9466), .ZN(n14018) );
  OR2_X1 U11963 ( .A1(n9513), .A2(n14018), .ZN(n9469) );
  INV_X1 U11964 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9467) );
  OR2_X1 U11965 ( .A1(n9562), .A2(n9467), .ZN(n9468) );
  NAND2_X1 U11966 ( .A1(n14268), .A2(n13486), .ZN(n9473) );
  OR2_X1 U11967 ( .A1(n14268), .A2(n13486), .ZN(n9472) );
  NAND2_X1 U11968 ( .A1(n9473), .A2(n9472), .ZN(n14014) );
  NAND2_X1 U11969 ( .A1(n13359), .A2(n13511), .ZN(n9475) );
  OR2_X1 U11970 ( .A1(n13514), .A2(n14307), .ZN(n9474) );
  NAND2_X1 U11971 ( .A1(n9512), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9483) );
  INV_X1 U11972 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9476) );
  OR2_X1 U11973 ( .A1(n9560), .A2(n9476), .ZN(n9482) );
  INV_X1 U11974 ( .A(n9478), .ZN(n9477) );
  NAND2_X1 U11975 ( .A1(n9477), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9497) );
  INV_X1 U11976 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n15228) );
  NAND2_X1 U11977 ( .A1(n9478), .A2(n15228), .ZN(n9479) );
  NAND2_X1 U11978 ( .A1(n9497), .A2(n9479), .ZN(n14002) );
  OR2_X1 U11979 ( .A1(n9513), .A2(n14002), .ZN(n9481) );
  INV_X1 U11980 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n15297) );
  OR2_X1 U11981 ( .A1(n13506), .A2(n15297), .ZN(n9480) );
  NAND2_X1 U11982 ( .A1(n14171), .A2(n13419), .ZN(n13981) );
  OR2_X1 U11983 ( .A1(n14171), .A2(n13419), .ZN(n9484) );
  NAND2_X1 U11984 ( .A1(n13981), .A2(n9484), .ZN(n13994) );
  INV_X1 U11985 ( .A(n13994), .ZN(n13998) );
  NAND2_X1 U11986 ( .A1(n13355), .A2(n13511), .ZN(n9486) );
  OR2_X1 U11987 ( .A1(n13514), .A2(n14306), .ZN(n9485) );
  NAND2_X1 U11988 ( .A1(n9512), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9491) );
  INV_X1 U11989 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n15318) );
  OR2_X1 U11990 ( .A1(n9560), .A2(n15318), .ZN(n9490) );
  INV_X1 U11991 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9496) );
  XNOR2_X1 U11992 ( .A(n9497), .B(n9496), .ZN(n13987) );
  OR2_X1 U11993 ( .A1(n9513), .A2(n13987), .ZN(n9489) );
  INV_X1 U11994 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9487) );
  OR2_X1 U11995 ( .A1(n13506), .A2(n9487), .ZN(n9488) );
  NAND4_X1 U11996 ( .A1(n9491), .A2(n9490), .A3(n9489), .A4(n9488), .ZN(n13773) );
  INV_X1 U11997 ( .A(n13773), .ZN(n13488) );
  NAND2_X1 U11998 ( .A1(n11548), .A2(n13511), .ZN(n9493) );
  OR2_X1 U11999 ( .A1(n13514), .A2(n11549), .ZN(n9492) );
  NAND2_X1 U12000 ( .A1(n13503), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9505) );
  INV_X1 U12001 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9494) );
  OR2_X1 U12002 ( .A1(n13505), .A2(n9494), .ZN(n9504) );
  INV_X1 U12003 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9495) );
  OAI21_X1 U12004 ( .B1(n9497), .B2(n9496), .A(n9495), .ZN(n9500) );
  INV_X1 U12005 ( .A(n9497), .ZN(n9499) );
  AND2_X1 U12006 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n9498) );
  NAND2_X1 U12007 ( .A1(n9499), .A2(n9498), .ZN(n13951) );
  NAND2_X1 U12008 ( .A1(n9500), .A2(n13951), .ZN(n13970) );
  OR2_X1 U12009 ( .A1(n9513), .A2(n13970), .ZN(n9503) );
  INV_X1 U12010 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9501) );
  OR2_X1 U12011 ( .A1(n9562), .A2(n9501), .ZN(n9502) );
  NAND2_X1 U12012 ( .A1(n13968), .A2(n13377), .ZN(n9508) );
  NAND2_X1 U12013 ( .A1(n9509), .A2(n9508), .ZN(n9519) );
  NAND2_X1 U12014 ( .A1(n13349), .A2(n13511), .ZN(n9511) );
  OR2_X1 U12015 ( .A1(n13514), .A2(n14304), .ZN(n9510) );
  NAND2_X1 U12016 ( .A1(n13503), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9518) );
  NAND2_X1 U12017 ( .A1(n9512), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9517) );
  OR2_X1 U12018 ( .A1(n9513), .A2(n13951), .ZN(n9516) );
  INV_X1 U12019 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9514) );
  OR2_X1 U12020 ( .A1(n9562), .A2(n9514), .ZN(n9515) );
  NAND4_X1 U12021 ( .A1(n9518), .A2(n9517), .A3(n9516), .A4(n9515), .ZN(n13772) );
  XNOR2_X1 U12022 ( .A(n13735), .B(n13772), .ZN(n13510) );
  XNOR2_X1 U12023 ( .A(n9519), .B(n13510), .ZN(n13963) );
  NAND2_X1 U12024 ( .A1(n14320), .A2(n14082), .ZN(n9525) );
  NAND2_X1 U12025 ( .A1(n6539), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9523) );
  NAND2_X1 U12026 ( .A1(n9566), .A2(n13550), .ZN(n13549) );
  NAND2_X1 U12027 ( .A1(n13562), .A2(n9526), .ZN(n14724) );
  NAND2_X1 U12028 ( .A1(n14729), .A2(n13560), .ZN(n14721) );
  NAND2_X1 U12029 ( .A1(n14724), .A2(n14721), .ZN(n9528) );
  INV_X1 U12030 ( .A(n14751), .ZN(n9977) );
  OR2_X1 U12031 ( .A1(n14728), .A2(n9977), .ZN(n9527) );
  INV_X1 U12032 ( .A(n10575), .ZN(n9529) );
  NAND2_X1 U12033 ( .A1(n10223), .A2(n10222), .ZN(n10221) );
  OR2_X1 U12034 ( .A1(n13797), .A2(n13394), .ZN(n9530) );
  INV_X1 U12035 ( .A(n10507), .ZN(n13583) );
  NAND2_X1 U12036 ( .A1(n13796), .A2(n13583), .ZN(n9531) );
  NAND2_X1 U12037 ( .A1(n14700), .A2(n14701), .ZN(n9533) );
  NAND2_X1 U12038 ( .A1(n14779), .A2(n13593), .ZN(n9532) );
  NAND2_X1 U12039 ( .A1(n9533), .A2(n9532), .ZN(n10757) );
  NAND2_X1 U12040 ( .A1(n10765), .A2(n10791), .ZN(n9535) );
  NOR2_X1 U12041 ( .A1(n13607), .A2(n13792), .ZN(n9536) );
  NAND2_X1 U12042 ( .A1(n13607), .A2(n13792), .ZN(n9537) );
  NAND2_X1 U12043 ( .A1(n14680), .A2(n14681), .ZN(n14679) );
  OR2_X1 U12044 ( .A1(n14693), .A2(n13791), .ZN(n9538) );
  NAND2_X1 U12045 ( .A1(n14679), .A2(n9538), .ZN(n11054) );
  NAND2_X1 U12046 ( .A1(n11054), .A2(n13529), .ZN(n11053) );
  INV_X1 U12047 ( .A(n11344), .ZN(n13790) );
  OR2_X1 U12048 ( .A1(n13618), .A2(n13790), .ZN(n9539) );
  NAND2_X1 U12049 ( .A1(n11053), .A2(n9539), .ZN(n11341) );
  INV_X1 U12050 ( .A(n11471), .ZN(n13789) );
  OR2_X1 U12051 ( .A1(n14563), .A2(n13789), .ZN(n9540) );
  INV_X1 U12052 ( .A(n11486), .ZN(n13788) );
  NAND2_X1 U12053 ( .A1(n14457), .A2(n14456), .ZN(n14455) );
  INV_X1 U12054 ( .A(n13636), .ZN(n13787) );
  OR2_X1 U12055 ( .A1(n13638), .A2(n13787), .ZN(n9541) );
  NAND2_X1 U12056 ( .A1(n14455), .A2(n9541), .ZN(n11499) );
  NAND2_X1 U12057 ( .A1(n11506), .A2(n13786), .ZN(n9542) );
  INV_X1 U12058 ( .A(n11752), .ZN(n13785) );
  OR2_X1 U12059 ( .A1(n14248), .A2(n13785), .ZN(n9543) );
  NAND2_X1 U12060 ( .A1(n9544), .A2(n9543), .ZN(n11533) );
  INV_X1 U12061 ( .A(n13656), .ZN(n13784) );
  OR2_X1 U12062 ( .A1(n13657), .A2(n13784), .ZN(n9545) );
  NOR2_X1 U12063 ( .A1(n14235), .A2(n13783), .ZN(n13663) );
  OR2_X1 U12064 ( .A1(n14230), .A2(n13782), .ZN(n13665) );
  NAND2_X1 U12065 ( .A1(n14230), .A2(n13782), .ZN(n13664) );
  NAND2_X1 U12066 ( .A1(n9546), .A2(n13664), .ZN(n14106) );
  NAND2_X1 U12067 ( .A1(n14062), .A2(n14061), .ZN(n14064) );
  NAND2_X1 U12068 ( .A1(n14281), .A2(n7138), .ZN(n9547) );
  NAND2_X1 U12069 ( .A1(n14064), .A2(n9547), .ZN(n14055) );
  NAND2_X1 U12070 ( .A1(n14049), .A2(n13777), .ZN(n9548) );
  NAND2_X1 U12071 ( .A1(n14057), .A2(n9548), .ZN(n14031) );
  OR2_X1 U12072 ( .A1(n13776), .A2(n14272), .ZN(n9549) );
  INV_X1 U12073 ( .A(n13486), .ZN(n13775) );
  NAND2_X1 U12074 ( .A1(n14268), .A2(n13775), .ZN(n9550) );
  NAND2_X1 U12075 ( .A1(n14012), .A2(n9550), .ZN(n13995) );
  NAND2_X1 U12076 ( .A1(n13995), .A2(n13994), .ZN(n9552) );
  INV_X1 U12077 ( .A(n13419), .ZN(n13774) );
  NAND2_X1 U12078 ( .A1(n14171), .A2(n13774), .ZN(n9551) );
  OR2_X1 U12079 ( .A1(n14165), .A2(n13773), .ZN(n9553) );
  XNOR2_X1 U12080 ( .A(n13968), .B(n13377), .ZN(n13967) );
  XNOR2_X1 U12081 ( .A(n9555), .B(n13510), .ZN(n13948) );
  NAND2_X1 U12082 ( .A1(n14320), .A2(n13929), .ZN(n9556) );
  NAND2_X1 U12083 ( .A1(n14320), .A2(n9970), .ZN(n9557) );
  NAND2_X1 U12084 ( .A1(n11838), .A2(n9557), .ZN(n10505) );
  NAND2_X1 U12085 ( .A1(n13948), .A2(n14807), .ZN(n9569) );
  INV_X1 U12086 ( .A(n14563), .ZN(n14575) );
  NAND2_X1 U12087 ( .A1(n10488), .A2(n10507), .ZN(n10590) );
  NOR2_X2 U12088 ( .A1(n14713), .A2(n13594), .ZN(n14714) );
  NAND2_X1 U12089 ( .A1(n10795), .A2(n14797), .ZN(n14686) );
  INV_X1 U12090 ( .A(n14290), .ZN(n14113) );
  INV_X1 U12091 ( .A(n14171), .ZN(n14005) );
  NAND2_X1 U12092 ( .A1(n13553), .A2(n13548), .ZN(n10506) );
  AOI21_X1 U12093 ( .B1(n13735), .B2(n6479), .A(n14788), .ZN(n9558) );
  NAND2_X1 U12094 ( .A1(n9558), .A2(n13942), .ZN(n13961) );
  INV_X1 U12095 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9559) );
  NOR2_X1 U12096 ( .A1(n9560), .A2(n9559), .ZN(n9565) );
  INV_X1 U12097 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9561) );
  NOR2_X1 U12098 ( .A1(n13505), .A2(n9561), .ZN(n9564) );
  INV_X1 U12099 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14259) );
  NOR2_X1 U12100 ( .A1(n9562), .A2(n14259), .ZN(n9563) );
  OR3_X1 U12101 ( .A1(n9565), .A2(n9564), .A3(n9563), .ZN(n13771) );
  INV_X1 U12102 ( .A(n13555), .ZN(n9987) );
  INV_X1 U12103 ( .A(n13815), .ZN(n9801) );
  INV_X1 U12104 ( .A(n14617), .ZN(n13810) );
  AND2_X1 U12105 ( .A1(n13810), .A2(P1_B_REG_SCAN_IN), .ZN(n9568) );
  NOR2_X1 U12106 ( .A1(n13487), .A2(n9568), .ZN(n13937) );
  NAND2_X1 U12107 ( .A1(n13771), .A2(n13937), .ZN(n13949) );
  NAND2_X1 U12108 ( .A1(n9506), .A2(n13478), .ZN(n13956) );
  INV_X1 U12109 ( .A(n9571), .ZN(n9572) );
  NAND2_X1 U12110 ( .A1(n9572), .A2(n9520), .ZN(n9587) );
  OAI21_X1 U12111 ( .B1(n9587), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9573) );
  MUX2_X1 U12112 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9573), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n9574) );
  NAND2_X1 U12113 ( .A1(n6451), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9576) );
  AND2_X1 U12114 ( .A1(n14310), .A2(P1_B_REG_SCAN_IN), .ZN(n9580) );
  NAND2_X1 U12115 ( .A1(n9577), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9579) );
  AOI21_X1 U12116 ( .B1(n11546), .B2(n9580), .A(n14309), .ZN(n9583) );
  INV_X1 U12117 ( .A(P1_B_REG_SCAN_IN), .ZN(n9581) );
  NAND2_X1 U12118 ( .A1(n9586), .A2(n9581), .ZN(n9582) );
  INV_X1 U12119 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9710) );
  NAND2_X1 U12120 ( .A1(n9702), .A2(n9710), .ZN(n9584) );
  NAND2_X1 U12121 ( .A1(n14309), .A2(n14310), .ZN(n9707) );
  NAND2_X1 U12122 ( .A1(n10500), .A2(n10494), .ZN(n9603) );
  INV_X1 U12123 ( .A(n14309), .ZN(n9585) );
  NAND2_X1 U12124 ( .A1(n9587), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9589) );
  NAND2_X1 U12125 ( .A1(n9590), .A2(n13929), .ZN(n9607) );
  AND2_X1 U12126 ( .A1(n13555), .A2(n9607), .ZN(n13765) );
  NOR2_X1 U12127 ( .A1(n13766), .A2(n13765), .ZN(n9602) );
  NOR4_X1 U12128 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9594) );
  NOR4_X1 U12129 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n9593) );
  NOR4_X1 U12130 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9592) );
  NOR4_X1 U12131 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9591) );
  AND4_X1 U12132 ( .A1(n9594), .A2(n9593), .A3(n9592), .A4(n9591), .ZN(n9600)
         );
  NOR2_X1 U12133 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .ZN(
        n9598) );
  NOR4_X1 U12134 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n9597) );
  NOR4_X1 U12135 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n9596) );
  NOR4_X1 U12136 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n9595) );
  AND4_X1 U12137 ( .A1(n9598), .A2(n9597), .A3(n9596), .A4(n9595), .ZN(n9599)
         );
  NAND2_X1 U12138 ( .A1(n9600), .A2(n9599), .ZN(n9601) );
  NAND2_X1 U12139 ( .A1(n9702), .A2(n9601), .ZN(n9968) );
  NAND2_X1 U12140 ( .A1(n9602), .A2(n9968), .ZN(n10501) );
  NOR2_X1 U12141 ( .A1(n9603), .A2(n10501), .ZN(n9611) );
  INV_X1 U12142 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9706) );
  NAND2_X1 U12143 ( .A1(n9702), .A2(n9706), .ZN(n9604) );
  NAND2_X1 U12144 ( .A1(n11546), .A2(n14309), .ZN(n9704) );
  OR2_X1 U12145 ( .A1(n14822), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9606) );
  INV_X1 U12146 ( .A(n9607), .ZN(n9608) );
  NAND2_X1 U12147 ( .A1(n14822), .A2(n14758), .ZN(n14205) );
  NAND2_X1 U12148 ( .A1(n13735), .A2(n9609), .ZN(n9610) );
  OR2_X1 U12149 ( .A1(n14810), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9613) );
  NAND2_X1 U12150 ( .A1(n14810), .A2(n14758), .ZN(n14282) );
  NAND2_X1 U12151 ( .A1(n13735), .A2(n9614), .ZN(n9615) );
  NOR2_X1 U12152 ( .A1(n9617), .A2(n9616), .ZN(n9689) );
  INV_X2 U12153 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U12154 ( .A(n11855), .ZN(n14434) );
  NAND2_X1 U12155 ( .A1(n9619), .A2(P3_U3151), .ZN(n14433) );
  INV_X1 U12156 ( .A(n10414), .ZN(n10426) );
  OAI222_X1 U12157 ( .A1(n14434), .A2(n6610), .B1(n14433), .B2(n7077), .C1(
        P3_U3151), .C2(n10426), .ZN(P3_U3294) );
  INV_X1 U12158 ( .A(SI_7_), .ZN(n9621) );
  OAI222_X1 U12159 ( .A1(P3_U3151), .A2(n10944), .B1(n14433), .B2(n9621), .C1(
        n14434), .C2(n9620), .ZN(P3_U3288) );
  INV_X1 U12160 ( .A(SI_4_), .ZN(n9623) );
  OAI222_X1 U12161 ( .A1(P3_U3151), .A2(n10624), .B1(n14433), .B2(n9623), .C1(
        n14434), .C2(n9622), .ZN(P3_U3291) );
  INV_X1 U12162 ( .A(SI_3_), .ZN(n9625) );
  OAI222_X1 U12163 ( .A1(P3_U3151), .A2(n10477), .B1(n14433), .B2(n9625), .C1(
        n14434), .C2(n9624), .ZN(P3_U3292) );
  INV_X1 U12164 ( .A(SI_5_), .ZN(n9627) );
  OAI222_X1 U12165 ( .A1(P3_U3151), .A2(n10627), .B1(n14433), .B2(n9627), .C1(
        n14434), .C2(n9626), .ZN(P3_U3290) );
  AND2_X1 U12166 ( .A1(n7171), .A2(P1_U3086), .ZN(n10390) );
  INV_X2 U12167 ( .A(n10390), .ZN(n14318) );
  NOR2_X1 U12168 ( .A1(n7171), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14314) );
  INV_X2 U12169 ( .A(n14314), .ZN(n14312) );
  OAI222_X1 U12170 ( .A1(n14318), .A2(n9628), .B1(n14312), .B2(n9648), .C1(
        P1_U3086), .C2(n13819), .ZN(P1_U3353) );
  OAI222_X1 U12171 ( .A1(n14312), .A2(n9654), .B1(n14318), .B2(n7653), .C1(
        P1_U3086), .C2(n9812), .ZN(P1_U3354) );
  INV_X1 U12172 ( .A(n9629), .ZN(n9644) );
  OAI222_X1 U12173 ( .A1(P1_U3086), .A2(n13834), .B1(n14312), .B2(n9644), .C1(
        n9630), .C2(n14318), .ZN(P1_U3352) );
  INV_X1 U12174 ( .A(n9631), .ZN(n9633) );
  INV_X1 U12175 ( .A(SI_8_), .ZN(n9632) );
  OAI222_X1 U12176 ( .A1(n14434), .A2(n9633), .B1(n14433), .B2(n9632), .C1(
        P3_U3151), .C2(n11081), .ZN(P3_U3287) );
  INV_X1 U12177 ( .A(SI_9_), .ZN(n9635) );
  OAI222_X1 U12178 ( .A1(P3_U3151), .A2(n11069), .B1(n14433), .B2(n9635), .C1(
        n14434), .C2(n9634), .ZN(P3_U3286) );
  INV_X1 U12179 ( .A(n14633), .ZN(n9796) );
  INV_X1 U12180 ( .A(n9636), .ZN(n9646) );
  OAI222_X1 U12181 ( .A1(P1_U3086), .A2(n9796), .B1(n14312), .B2(n9646), .C1(
        n9637), .C2(n14318), .ZN(P1_U3351) );
  INV_X1 U12182 ( .A(n14433), .ZN(n11856) );
  INV_X1 U12183 ( .A(n11856), .ZN(n11873) );
  AOI22_X1 U12184 ( .A1(n11855), .A2(n9638), .B1(P3_IR_REG_0__SCAN_IN), .B2(
        P3_STATE_REG_SCAN_IN), .ZN(n9639) );
  OAI21_X1 U12185 ( .B1(n9640), .B2(n11873), .A(n9639), .ZN(P3_U3295) );
  INV_X1 U12186 ( .A(n9641), .ZN(n9651) );
  INV_X1 U12187 ( .A(n9819), .ZN(n9835) );
  OAI222_X1 U12188 ( .A1(n14318), .A2(n9642), .B1(n14312), .B2(n9651), .C1(
        n9835), .C2(P1_U3086), .ZN(P1_U3350) );
  NOR2_X1 U12189 ( .A1(n7171), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13352) );
  INV_X2 U12190 ( .A(n13352), .ZN(n13372) );
  NAND2_X1 U12191 ( .A1(n7171), .A2(P2_U3088), .ZN(n13367) );
  INV_X1 U12192 ( .A(n13367), .ZN(n13369) );
  INV_X1 U12193 ( .A(n13369), .ZN(n13357) );
  INV_X1 U12194 ( .A(n14845), .ZN(n9643) );
  OAI222_X1 U12195 ( .A1(n13372), .A2(n9645), .B1(n13357), .B2(n9644), .C1(
        n9643), .C2(P2_U3088), .ZN(P2_U3324) );
  OAI222_X1 U12196 ( .A1(n13372), .A2(n9647), .B1(n13357), .B2(n9646), .C1(
        n9889), .C2(P2_U3088), .ZN(P2_U3323) );
  OAI222_X1 U12197 ( .A1(n13372), .A2(n9649), .B1(n13357), .B2(n9648), .C1(
        P2_U3088), .C2(n12924), .ZN(P2_U3325) );
  INV_X1 U12198 ( .A(n12933), .ZN(n9650) );
  OAI222_X1 U12199 ( .A1(n13372), .A2(n9652), .B1(n13357), .B2(n9651), .C1(
        n9650), .C2(P2_U3088), .ZN(P2_U3322) );
  OAI222_X1 U12200 ( .A1(P2_U3088), .A2(n9885), .B1(n13367), .B2(n9654), .C1(
        n9653), .C2(n13372), .ZN(P2_U3326) );
  OAI222_X1 U12201 ( .A1(P3_U3151), .A2(n11423), .B1(n11873), .B2(n9656), .C1(
        n14434), .C2(n9655), .ZN(P3_U3284) );
  INV_X1 U12202 ( .A(SI_10_), .ZN(n9658) );
  OAI222_X1 U12203 ( .A1(P3_U3151), .A2(n15067), .B1(n11873), .B2(n9658), .C1(
        n14434), .C2(n9657), .ZN(P3_U3285) );
  INV_X1 U12204 ( .A(n9659), .ZN(n9661) );
  OAI222_X1 U12205 ( .A1(P3_U3151), .A2(n10722), .B1(n14434), .B2(n9661), .C1(
        n9660), .C2(n11873), .ZN(P3_U3293) );
  INV_X1 U12206 ( .A(n9662), .ZN(n9664) );
  INV_X1 U12207 ( .A(SI_6_), .ZN(n9663) );
  OAI222_X1 U12208 ( .A1(P3_U3151), .A2(n10956), .B1(n14434), .B2(n9664), .C1(
        n9663), .C2(n11873), .ZN(P3_U3289) );
  INV_X1 U12209 ( .A(n9665), .ZN(n9668) );
  INV_X1 U12210 ( .A(n12945), .ZN(n9666) );
  OAI222_X1 U12211 ( .A1(n13372), .A2(n9667), .B1(n13357), .B2(n9668), .C1(
        n9666), .C2(P2_U3088), .ZN(P2_U3321) );
  INV_X1 U12212 ( .A(n9837), .ZN(n13843) );
  OAI222_X1 U12213 ( .A1(n14318), .A2(n9669), .B1(n14312), .B2(n9668), .C1(
        n13843), .C2(P1_U3086), .ZN(P1_U3349) );
  INV_X1 U12214 ( .A(n12957), .ZN(n9670) );
  OAI222_X1 U12215 ( .A1(n13372), .A2(n9671), .B1(n13357), .B2(n9672), .C1(
        n9670), .C2(P2_U3088), .ZN(P2_U3320) );
  INV_X1 U12216 ( .A(n9838), .ZN(n13856) );
  OAI222_X1 U12217 ( .A1(n14318), .A2(n9673), .B1(n14312), .B2(n9672), .C1(
        n13856), .C2(P1_U3086), .ZN(P1_U3348) );
  NAND2_X1 U12218 ( .A1(n6445), .A2(P2_U3947), .ZN(n9674) );
  OAI21_X1 U12219 ( .B1(n9171), .B2(P2_U3947), .A(n9674), .ZN(P2_U3531) );
  AOI222_X1 U12220 ( .A1(n9675), .A2(n11855), .B1(n15083), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_12_), .C2(n11856), .ZN(n9676) );
  INV_X1 U12221 ( .A(n9676), .ZN(P3_U3283) );
  INV_X1 U12222 ( .A(n9856), .ZN(n9851) );
  OAI222_X1 U12223 ( .A1(n14318), .A2(n9677), .B1(n14312), .B2(n9678), .C1(
        n9851), .C2(P1_U3086), .ZN(P1_U3347) );
  INV_X1 U12224 ( .A(n9894), .ZN(n14874) );
  OAI222_X1 U12225 ( .A1(n13372), .A2(n9679), .B1(n13357), .B2(n9678), .C1(
        n14874), .C2(P2_U3088), .ZN(P2_U3319) );
  AOI222_X1 U12226 ( .A1(n9680), .A2(n11855), .B1(n12336), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_13_), .C2(n11856), .ZN(n9681) );
  INV_X1 U12227 ( .A(n9681), .ZN(P3_U3282) );
  INV_X1 U12228 ( .A(n9857), .ZN(n10146) );
  OAI222_X1 U12229 ( .A1(n14318), .A2(n9682), .B1(n14312), .B2(n9683), .C1(
        n10146), .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U12230 ( .A(n9896), .ZN(n14887) );
  OAI222_X1 U12231 ( .A1(n13372), .A2(n9684), .B1(n13357), .B2(n9683), .C1(
        n14887), .C2(P2_U3088), .ZN(P2_U3318) );
  NAND2_X1 U12232 ( .A1(n9744), .A2(n9685), .ZN(n9686) );
  AND2_X1 U12233 ( .A1(n9687), .A2(n9686), .ZN(n9688) );
  OR2_X1 U12234 ( .A1(n9689), .A2(n9688), .ZN(n9697) );
  NOR2_X1 U12235 ( .A1(n8497), .A2(P2_U3088), .ZN(n13351) );
  NAND2_X1 U12236 ( .A1(n9691), .A2(n13356), .ZN(n14960) );
  INV_X1 U12237 ( .A(n13356), .ZN(n9690) );
  AND2_X1 U12238 ( .A1(n9691), .A2(n9690), .ZN(n14985) );
  INV_X1 U12239 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10087) );
  NAND2_X1 U12240 ( .A1(n14985), .A2(n10087), .ZN(n9692) );
  AND2_X1 U12241 ( .A1(n8497), .A2(n9697), .ZN(n14908) );
  NAND2_X1 U12242 ( .A1(n14908), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14979) );
  OAI211_X1 U12243 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n14960), .A(n9692), .B(
        n14979), .ZN(n9693) );
  INV_X1 U12244 ( .A(n9693), .ZN(n9696) );
  AOI22_X1 U12245 ( .A1(n14977), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n14985), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n9695) );
  MUX2_X1 U12246 ( .A(n9696), .B(n9695), .S(n9694), .Z(n9699) );
  AOI22_X1 U12247 ( .A1(n14823), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n9698) );
  NAND2_X1 U12248 ( .A1(n9699), .A2(n9698), .ZN(P2_U3214) );
  OAI222_X1 U12249 ( .A1(P3_U3151), .A2(n12344), .B1(n11873), .B2(n9701), .C1(
        n14434), .C2(n9700), .ZN(P3_U3281) );
  INV_X1 U12250 ( .A(n9702), .ZN(n9703) );
  NAND2_X1 U12251 ( .A1(n9703), .A2(n10496), .ZN(n14748) );
  INV_X1 U12252 ( .A(n9704), .ZN(n9705) );
  AOI22_X1 U12253 ( .A1(n14748), .A2(n9706), .B1(n9705), .B2(n9709), .ZN(
        P1_U3445) );
  INV_X1 U12254 ( .A(n9707), .ZN(n9708) );
  AOI22_X1 U12255 ( .A1(n14748), .A2(n9710), .B1(n9709), .B2(n9708), .ZN(
        P1_U3446) );
  INV_X1 U12256 ( .A(n10261), .ZN(n9711) );
  NAND2_X1 U12257 ( .A1(n9711), .A2(n9713), .ZN(n9712) );
  OAI21_X1 U12258 ( .B1(n9713), .B2(n15298), .A(n9712), .ZN(P3_U3377) );
  NOR4_X1 U12259 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9717) );
  NOR4_X1 U12260 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n9716) );
  NOR4_X1 U12261 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9715) );
  NOR4_X1 U12262 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9714) );
  NAND4_X1 U12263 ( .A1(n9717), .A2(n9716), .A3(n9715), .A4(n9714), .ZN(n9726)
         );
  NOR2_X1 U12264 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .ZN(
        n9721) );
  NOR4_X1 U12265 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n9720) );
  NOR4_X1 U12266 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9719) );
  NOR4_X1 U12267 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n9718) );
  NAND4_X1 U12268 ( .A1(n9721), .A2(n9720), .A3(n9719), .A4(n9718), .ZN(n9725)
         );
  XNOR2_X1 U12269 ( .A(n9727), .B(n11697), .ZN(n9722) );
  NAND2_X1 U12270 ( .A1(n9722), .A2(n13363), .ZN(n9724) );
  INV_X1 U12271 ( .A(n13361), .ZN(n9723) );
  OAI21_X1 U12272 ( .B1(n9726), .B2(n9725), .A(n14990), .ZN(n10078) );
  INV_X1 U12273 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14993) );
  NAND2_X1 U12274 ( .A1(n14990), .A2(n14993), .ZN(n9729) );
  INV_X1 U12275 ( .A(n9727), .ZN(n13365) );
  NAND2_X1 U12276 ( .A1(n13365), .A2(n13361), .ZN(n9728) );
  NAND2_X1 U12277 ( .A1(n9729), .A2(n9728), .ZN(n14994) );
  NOR2_X1 U12278 ( .A1(n14994), .A2(n14995), .ZN(n9732) );
  INV_X1 U12279 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14996) );
  NAND2_X1 U12280 ( .A1(n14990), .A2(n14996), .ZN(n9731) );
  NAND2_X1 U12281 ( .A1(n13361), .A2(n13363), .ZN(n9730) );
  NAND2_X1 U12282 ( .A1(n9731), .A2(n9730), .ZN(n14997) );
  INV_X1 U12283 ( .A(n14997), .ZN(n10079) );
  AND3_X1 U12284 ( .A1(n10078), .A2(n9732), .A3(n10079), .ZN(n9743) );
  AND2_X2 U12285 ( .A1(n9741), .A2(n9772), .ZN(n15019) );
  NOR2_X1 U12286 ( .A1(n15019), .A2(n9744), .ZN(n9733) );
  INV_X1 U12287 ( .A(n12902), .ZN(n12871) );
  NAND2_X2 U12288 ( .A1(n9772), .A2(n11372), .ZN(n15030) );
  NAND2_X1 U12289 ( .A1(n10158), .A2(n13194), .ZN(n9754) );
  AND3_X1 U12290 ( .A1(n6795), .A2(n11445), .A3(n7762), .ZN(n10090) );
  NAND2_X1 U12291 ( .A1(n9743), .A2(n10090), .ZN(n9735) );
  AOI21_X1 U12292 ( .B1(n12871), .B2(n9754), .A(n12900), .ZN(n9747) );
  NOR2_X1 U12293 ( .A1(n14994), .A2(n14997), .ZN(n9736) );
  NAND2_X1 U12294 ( .A1(n10078), .A2(n9736), .ZN(n9737) );
  NAND2_X1 U12295 ( .A1(n9737), .A2(n9779), .ZN(n9740) );
  NAND2_X1 U12296 ( .A1(n9741), .A2(n9744), .ZN(n9781) );
  AND2_X1 U12297 ( .A1(n9738), .A2(n9781), .ZN(n9739) );
  NAND2_X1 U12298 ( .A1(n9740), .A2(n9739), .ZN(n9934) );
  NOR2_X1 U12299 ( .A1(n9934), .A2(P2_U3088), .ZN(n9924) );
  INV_X1 U12300 ( .A(n9924), .ZN(n9764) );
  INV_X1 U12301 ( .A(n9741), .ZN(n9742) );
  NAND2_X1 U12302 ( .A1(n9743), .A2(n9742), .ZN(n11613) );
  NAND2_X1 U12303 ( .A1(n8497), .A2(n9744), .ZN(n13141) );
  OR2_X1 U12304 ( .A1(n11613), .A2(n13141), .ZN(n12890) );
  AOI22_X1 U12305 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n9764), .B1(n12848), .B2(
        n9755), .ZN(n9746) );
  OR2_X1 U12306 ( .A1(n12902), .A2(n11580), .ZN(n12860) );
  NAND3_X1 U12307 ( .A1(n12893), .A2(n6445), .A3(n6927), .ZN(n9745) );
  OAI211_X1 U12308 ( .C1(n9747), .C2(n10010), .A(n9746), .B(n9745), .ZN(
        P2_U3204) );
  AOI222_X1 U12309 ( .A1(n9748), .A2(n11855), .B1(n12370), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_15_), .C2(n11856), .ZN(n9749) );
  INV_X1 U12310 ( .A(n9749), .ZN(P3_U3280) );
  XNOR2_X1 U12311 ( .A(n9750), .B(n7762), .ZN(n9751) );
  NAND2_X1 U12312 ( .A1(n11584), .A2(n10010), .ZN(n9753) );
  NAND2_X1 U12313 ( .A1(n9754), .A2(n9753), .ZN(n9763) );
  NAND2_X1 U12314 ( .A1(n9756), .A2(n9757), .ZN(n9919) );
  NAND2_X1 U12315 ( .A1(n9919), .A2(n9758), .ZN(n9762) );
  INV_X1 U12316 ( .A(n9762), .ZN(n9760) );
  INV_X1 U12317 ( .A(n9763), .ZN(n9759) );
  NAND2_X1 U12318 ( .A1(n9760), .A2(n9759), .ZN(n9920) );
  INV_X1 U12319 ( .A(n9920), .ZN(n9761) );
  AOI21_X1 U12320 ( .B1(n9763), .B2(n9762), .A(n9761), .ZN(n9767) );
  AOI22_X1 U12321 ( .A1(n9764), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n10168), .B2(
        n12900), .ZN(n9766) );
  INV_X1 U12322 ( .A(n12896), .ZN(n12847) );
  AOI22_X1 U12323 ( .A1(n12848), .A2(n12916), .B1(n12847), .B2(n6445), .ZN(
        n9765) );
  OAI211_X1 U12324 ( .C1(n9767), .C2(n12902), .A(n9766), .B(n9765), .ZN(
        P2_U3194) );
  INV_X1 U12325 ( .A(n11292), .ZN(n9768) );
  OAI222_X1 U12326 ( .A1(n13372), .A2(n9769), .B1(n13357), .B2(n9271), .C1(
        n9768), .C2(P2_U3088), .ZN(P2_U3317) );
  INV_X1 U12327 ( .A(n10148), .ZN(n13875) );
  OAI222_X1 U12328 ( .A1(P1_U3086), .A2(n13875), .B1(n14312), .B2(n9271), .C1(
        n9770), .C2(n14318), .ZN(P1_U3345) );
  INV_X1 U12329 ( .A(n15023), .ZN(n15033) );
  INV_X1 U12330 ( .A(n10093), .ZN(n9778) );
  INV_X1 U12331 ( .A(n9772), .ZN(n9773) );
  OAI22_X1 U12332 ( .A1(n10093), .A2(n9771), .B1(n9773), .B2(n10010), .ZN(
        n9777) );
  NAND2_X1 U12333 ( .A1(n6795), .A2(n9774), .ZN(n9775) );
  INV_X1 U12334 ( .A(n13228), .ZN(n13137) );
  INV_X1 U12335 ( .A(n9755), .ZN(n9923) );
  OAI22_X1 U12336 ( .A1(n10093), .A2(n13137), .B1(n9923), .B2(n13141), .ZN(
        n10089) );
  AOI211_X1 U12337 ( .C1(n15033), .C2(n9778), .A(n9777), .B(n10089), .ZN(
        n15000) );
  AND2_X1 U12338 ( .A1(n14997), .A2(n9779), .ZN(n9780) );
  AND2_X1 U12339 ( .A1(n10078), .A2(n9780), .ZN(n10016) );
  NAND2_X1 U12340 ( .A1(n14998), .A2(n9781), .ZN(n10081) );
  NAND2_X1 U12341 ( .A1(n15045), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9783) );
  OAI21_X1 U12342 ( .B1(n15000), .B2(n15045), .A(n9783), .ZN(P2_U3499) );
  INV_X1 U12343 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9785) );
  NOR2_X1 U12344 ( .A1(n10094), .A2(n9785), .ZN(P3_U3258) );
  INV_X1 U12345 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n15225) );
  NOR2_X1 U12346 ( .A1(n10094), .A2(n15225), .ZN(P3_U3260) );
  INV_X1 U12347 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9786) );
  NOR2_X1 U12348 ( .A1(n10094), .A2(n9786), .ZN(P3_U3259) );
  INV_X1 U12349 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9787) );
  NOR2_X1 U12350 ( .A1(n10094), .A2(n9787), .ZN(P3_U3247) );
  AOI222_X1 U12351 ( .A1(n9788), .A2(n11855), .B1(n12373), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_16_), .C2(n11856), .ZN(n9789) );
  INV_X1 U12352 ( .A(n9789), .ZN(P3_U3279) );
  MUX2_X1 U12353 ( .A(n9828), .B(P1_REG1_REG_5__SCAN_IN), .S(n9819), .Z(n9798)
         );
  INV_X1 U12354 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9795) );
  INV_X1 U12355 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n14813) );
  MUX2_X1 U12356 ( .A(n14813), .B(P1_REG1_REG_2__SCAN_IN), .S(n13819), .Z(
        n13823) );
  INV_X1 U12357 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n14811) );
  MUX2_X1 U12358 ( .A(n14811), .B(P1_REG1_REG_1__SCAN_IN), .S(n9812), .Z(
        n13802) );
  AND2_X1 U12359 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n13801) );
  NAND2_X1 U12360 ( .A1(n13802), .A2(n13801), .ZN(n13800) );
  INV_X1 U12361 ( .A(n9812), .ZN(n13805) );
  NAND2_X1 U12362 ( .A1(n13805), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9790) );
  NAND2_X1 U12363 ( .A1(n13800), .A2(n9790), .ZN(n13822) );
  NAND2_X1 U12364 ( .A1(n13823), .A2(n13822), .ZN(n13821) );
  OR2_X1 U12365 ( .A1(n13819), .A2(n14813), .ZN(n9791) );
  NAND2_X1 U12366 ( .A1(n13821), .A2(n9791), .ZN(n13832) );
  INV_X1 U12367 ( .A(n13834), .ZN(n9816) );
  NAND2_X1 U12368 ( .A1(n9816), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9794) );
  INV_X1 U12369 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9792) );
  NAND2_X1 U12370 ( .A1(n13834), .A2(n9792), .ZN(n9793) );
  AND2_X1 U12371 ( .A1(n9794), .A2(n9793), .ZN(n13833) );
  NAND2_X1 U12372 ( .A1(n13832), .A2(n13833), .ZN(n13831) );
  NAND2_X1 U12373 ( .A1(n13831), .A2(n9794), .ZN(n14635) );
  XNOR2_X1 U12374 ( .A(n14633), .B(n9795), .ZN(n14636) );
  NAND2_X1 U12375 ( .A1(n14635), .A2(n14636), .ZN(n14634) );
  OAI21_X1 U12376 ( .B1(n9796), .B2(n9795), .A(n14634), .ZN(n9797) );
  NOR2_X1 U12377 ( .A1(n9797), .A2(n9798), .ZN(n9827) );
  AOI21_X1 U12378 ( .B1(n9798), .B2(n9797), .A(n9827), .ZN(n9826) );
  OR2_X1 U12379 ( .A1(n9800), .A2(P1_U3086), .ZN(n14316) );
  NAND2_X1 U12380 ( .A1(n13766), .A2(n14316), .ZN(n9804) );
  AOI21_X1 U12381 ( .B1(n13555), .B2(n9800), .A(n9799), .ZN(n9802) );
  NAND2_X1 U12382 ( .A1(n9804), .A2(n9802), .ZN(n14627) );
  OR2_X1 U12383 ( .A1(n14627), .A2(n9801), .ZN(n13924) );
  INV_X1 U12384 ( .A(n13924), .ZN(n14669) );
  INV_X1 U12385 ( .A(n9802), .ZN(n9803) );
  AND2_X1 U12386 ( .A1(n9804), .A2(n9803), .ZN(n14624) );
  INV_X1 U12387 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9805) );
  NAND2_X1 U12388 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10541) );
  OAI21_X1 U12389 ( .B1(n14677), .B2(n9805), .A(n10541), .ZN(n9806) );
  AOI21_X1 U12390 ( .B1(n9819), .B2(n14669), .A(n9806), .ZN(n9825) );
  OR2_X1 U12391 ( .A1(n13815), .A2(n14617), .ZN(n9807) );
  INV_X1 U12392 ( .A(n14672), .ZN(n14656) );
  MUX2_X1 U12393 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9808), .S(n14633), .Z(n9818) );
  MUX2_X1 U12394 ( .A(n9809), .B(P1_REG2_REG_2__SCAN_IN), .S(n13819), .Z(
        n13825) );
  MUX2_X1 U12395 ( .A(n9810), .B(P1_REG2_REG_1__SCAN_IN), .S(n9812), .Z(n13804) );
  AND2_X1 U12396 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9811) );
  NAND2_X1 U12397 ( .A1(n13804), .A2(n9811), .ZN(n13803) );
  OAI21_X1 U12398 ( .B1(n9810), .B2(n9812), .A(n13803), .ZN(n13824) );
  NAND2_X1 U12399 ( .A1(n13825), .A2(n13824), .ZN(n13837) );
  OR2_X1 U12400 ( .A1(n13819), .A2(n9809), .ZN(n13836) );
  NAND2_X1 U12401 ( .A1(n13837), .A2(n13836), .ZN(n9815) );
  MUX2_X1 U12402 ( .A(n9813), .B(P1_REG2_REG_3__SCAN_IN), .S(n13834), .Z(n9814) );
  NAND2_X1 U12403 ( .A1(n9815), .A2(n9814), .ZN(n14629) );
  NAND2_X1 U12404 ( .A1(n9816), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14628) );
  NAND2_X1 U12405 ( .A1(n14629), .A2(n14628), .ZN(n9817) );
  NAND2_X1 U12406 ( .A1(n9818), .A2(n9817), .ZN(n14632) );
  NAND2_X1 U12407 ( .A1(n14633), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9821) );
  INV_X1 U12408 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9834) );
  MUX2_X1 U12409 ( .A(n9834), .B(P1_REG2_REG_5__SCAN_IN), .S(n9819), .Z(n9820)
         );
  AOI21_X1 U12410 ( .B1(n14632), .B2(n9821), .A(n9820), .ZN(n13851) );
  INV_X1 U12411 ( .A(n13851), .ZN(n9823) );
  NAND3_X1 U12412 ( .A1(n14632), .A2(n9821), .A3(n9820), .ZN(n9822) );
  NAND3_X1 U12413 ( .A1(n14656), .A2(n9823), .A3(n9822), .ZN(n9824) );
  OAI211_X1 U12414 ( .C1(n9826), .C2(n13799), .A(n9825), .B(n9824), .ZN(
        P1_U3248) );
  MUX2_X1 U12415 ( .A(n9850), .B(P1_REG1_REG_8__SCAN_IN), .S(n9856), .Z(n9831)
         );
  AOI21_X1 U12416 ( .B1(n9835), .B2(n9828), .A(n9827), .ZN(n13847) );
  INV_X1 U12417 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14817) );
  MUX2_X1 U12418 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n14817), .S(n9837), .Z(
        n13848) );
  NAND2_X1 U12419 ( .A1(n13847), .A2(n13848), .ZN(n13846) );
  OAI21_X1 U12420 ( .B1(n14817), .B2(n13843), .A(n13846), .ZN(n13860) );
  MUX2_X1 U12421 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9829), .S(n9838), .Z(n13861) );
  NAND2_X1 U12422 ( .A1(n13860), .A2(n13861), .ZN(n13859) );
  OAI21_X1 U12423 ( .B1(n9829), .B2(n13856), .A(n13859), .ZN(n9830) );
  NOR2_X1 U12424 ( .A1(n9830), .A2(n9831), .ZN(n9849) );
  AOI21_X1 U12425 ( .B1(n9831), .B2(n9830), .A(n9849), .ZN(n9848) );
  NOR2_X1 U12426 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10850), .ZN(n9833) );
  NOR2_X1 U12427 ( .A1(n13924), .A2(n9851), .ZN(n9832) );
  AOI211_X1 U12428 ( .C1(n14624), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n9833), .B(
        n9832), .ZN(n9847) );
  NOR2_X1 U12429 ( .A1(n9835), .A2(n9834), .ZN(n13849) );
  MUX2_X1 U12430 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9836), .S(n9837), .Z(n13850) );
  OAI21_X1 U12431 ( .B1(n13851), .B2(n13849), .A(n13850), .ZN(n13865) );
  NAND2_X1 U12432 ( .A1(n9837), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n13864) );
  INV_X1 U12433 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9839) );
  MUX2_X1 U12434 ( .A(n9839), .B(P1_REG2_REG_7__SCAN_IN), .S(n9838), .Z(n13863) );
  AOI21_X1 U12435 ( .B1(n13865), .B2(n13864), .A(n13863), .ZN(n13862) );
  NOR2_X1 U12436 ( .A1(n13856), .A2(n9839), .ZN(n9844) );
  INV_X1 U12437 ( .A(n9844), .ZN(n9842) );
  INV_X1 U12438 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9840) );
  MUX2_X1 U12439 ( .A(n9840), .B(P1_REG2_REG_8__SCAN_IN), .S(n9856), .Z(n9841)
         );
  NAND2_X1 U12440 ( .A1(n9842), .A2(n9841), .ZN(n9845) );
  MUX2_X1 U12441 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n9840), .S(n9856), .Z(n9843)
         );
  OAI21_X1 U12442 ( .B1(n13862), .B2(n9844), .A(n9843), .ZN(n9860) );
  OAI211_X1 U12443 ( .C1(n13862), .C2(n9845), .A(n14656), .B(n9860), .ZN(n9846) );
  OAI211_X1 U12444 ( .C1(n9848), .C2(n13799), .A(n9847), .B(n9846), .ZN(
        P1_U3251) );
  MUX2_X1 U12445 ( .A(n10139), .B(P1_REG1_REG_9__SCAN_IN), .S(n9857), .Z(n9853) );
  AOI21_X1 U12446 ( .B1(n9851), .B2(n9850), .A(n9849), .ZN(n9852) );
  NOR2_X1 U12447 ( .A1(n9852), .A2(n9853), .ZN(n10138) );
  AOI21_X1 U12448 ( .B1(n9853), .B2(n9852), .A(n10138), .ZN(n9865) );
  NOR2_X1 U12449 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n15259), .ZN(n9855) );
  NOR2_X1 U12450 ( .A1(n13924), .A2(n10146), .ZN(n9854) );
  AOI211_X1 U12451 ( .C1(n14624), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n9855), .B(
        n9854), .ZN(n9864) );
  NAND2_X1 U12452 ( .A1(n9856), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9859) );
  MUX2_X1 U12453 ( .A(n14690), .B(P1_REG2_REG_9__SCAN_IN), .S(n9857), .Z(n9858) );
  AOI21_X1 U12454 ( .B1(n9860), .B2(n9859), .A(n9858), .ZN(n13880) );
  INV_X1 U12455 ( .A(n13880), .ZN(n9862) );
  NAND3_X1 U12456 ( .A1(n9860), .A2(n9859), .A3(n9858), .ZN(n9861) );
  NAND3_X1 U12457 ( .A1(n9862), .A2(n14656), .A3(n9861), .ZN(n9863) );
  OAI211_X1 U12458 ( .C1(n9865), .C2(n13799), .A(n9864), .B(n9863), .ZN(
        P1_U3252) );
  INV_X1 U12459 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9866) );
  MUX2_X1 U12460 ( .A(n9866), .B(P2_REG2_REG_10__SCAN_IN), .S(n11292), .Z(
        n9883) );
  INV_X1 U12461 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10368) );
  MUX2_X1 U12462 ( .A(n10368), .B(P2_REG2_REG_2__SCAN_IN), .S(n12924), .Z(
        n12920) );
  INV_X1 U12463 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10358) );
  MUX2_X1 U12464 ( .A(n10358), .B(P2_REG2_REG_1__SCAN_IN), .S(n9885), .Z(
        n14828) );
  NAND2_X1 U12465 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n14829) );
  INV_X1 U12466 ( .A(n14829), .ZN(n9867) );
  NAND2_X1 U12467 ( .A1(n14828), .A2(n9867), .ZN(n14832) );
  INV_X1 U12468 ( .A(n9885), .ZN(n14827) );
  NAND2_X1 U12469 ( .A1(n14827), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9868) );
  NAND2_X1 U12470 ( .A1(n14832), .A2(n9868), .ZN(n12919) );
  NAND2_X1 U12471 ( .A1(n12920), .A2(n12919), .ZN(n12918) );
  OR2_X1 U12472 ( .A1(n12924), .A2(n10368), .ZN(n9869) );
  NAND2_X1 U12473 ( .A1(n12918), .A2(n9869), .ZN(n14843) );
  INV_X1 U12474 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10430) );
  MUX2_X1 U12475 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10430), .S(n14845), .Z(
        n14844) );
  NAND2_X1 U12476 ( .A1(n14843), .A2(n14844), .ZN(n14842) );
  NAND2_X1 U12477 ( .A1(n14845), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9870) );
  NAND2_X1 U12478 ( .A1(n14842), .A2(n9870), .ZN(n14856) );
  INV_X1 U12479 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9871) );
  MUX2_X1 U12480 ( .A(n9871), .B(P2_REG2_REG_4__SCAN_IN), .S(n9889), .Z(n14857) );
  NAND2_X1 U12481 ( .A1(n14856), .A2(n14857), .ZN(n14855) );
  NAND2_X1 U12482 ( .A1(n14858), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9872) );
  NAND2_X1 U12483 ( .A1(n14855), .A2(n9872), .ZN(n12938) );
  INV_X1 U12484 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9873) );
  MUX2_X1 U12485 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n9873), .S(n12933), .Z(
        n12939) );
  NAND2_X1 U12486 ( .A1(n12938), .A2(n12939), .ZN(n12937) );
  NAND2_X1 U12487 ( .A1(n12933), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9874) );
  NAND2_X1 U12488 ( .A1(n12937), .A2(n9874), .ZN(n12947) );
  INV_X1 U12489 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10253) );
  XNOR2_X1 U12490 ( .A(n12945), .B(n10253), .ZN(n12948) );
  NAND2_X1 U12491 ( .A1(n12947), .A2(n12948), .ZN(n12946) );
  NAND2_X1 U12492 ( .A1(n12945), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9875) );
  NAND2_X1 U12493 ( .A1(n12946), .A2(n9875), .ZN(n12960) );
  INV_X1 U12494 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9876) );
  MUX2_X1 U12495 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9876), .S(n12957), .Z(
        n12959) );
  NAND2_X1 U12496 ( .A1(n12960), .A2(n12959), .ZN(n12958) );
  NAND2_X1 U12497 ( .A1(n12957), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9877) );
  NAND2_X1 U12498 ( .A1(n12958), .A2(n9877), .ZN(n14871) );
  INV_X1 U12499 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9878) );
  MUX2_X1 U12500 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n9878), .S(n9894), .Z(n14870) );
  NAND2_X1 U12501 ( .A1(n14871), .A2(n14870), .ZN(n14869) );
  NAND2_X1 U12502 ( .A1(n9894), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9879) );
  NAND2_X1 U12503 ( .A1(n14869), .A2(n9879), .ZN(n14884) );
  XNOR2_X1 U12504 ( .A(n9896), .B(P2_REG2_REG_9__SCAN_IN), .ZN(n14883) );
  OR2_X1 U12505 ( .A1(n14884), .A2(n14883), .ZN(n14886) );
  INV_X1 U12506 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10887) );
  NAND2_X1 U12507 ( .A1(n14887), .A2(n10887), .ZN(n9880) );
  NAND2_X1 U12508 ( .A1(n14886), .A2(n9880), .ZN(n9882) );
  INV_X1 U12509 ( .A(n11294), .ZN(n9881) );
  AOI211_X1 U12510 ( .C1(n9883), .C2(n9882), .A(n14965), .B(n9881), .ZN(n9904)
         );
  INV_X1 U12511 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9884) );
  MUX2_X1 U12512 ( .A(n9884), .B(P2_REG1_REG_10__SCAN_IN), .S(n11292), .Z(
        n9900) );
  INV_X1 U12513 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10044) );
  MUX2_X1 U12514 ( .A(n10044), .B(P2_REG1_REG_2__SCAN_IN), .S(n12924), .Z(
        n12923) );
  INV_X1 U12515 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10174) );
  MUX2_X1 U12516 ( .A(n10174), .B(P2_REG1_REG_1__SCAN_IN), .S(n9885), .Z(
        n14826) );
  AND2_X1 U12517 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14825) );
  NAND2_X1 U12518 ( .A1(n14826), .A2(n14825), .ZN(n14824) );
  NAND2_X1 U12519 ( .A1(n14827), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9886) );
  NAND2_X1 U12520 ( .A1(n14824), .A2(n9886), .ZN(n12922) );
  NAND2_X1 U12521 ( .A1(n12923), .A2(n12922), .ZN(n12921) );
  OR2_X1 U12522 ( .A1(n12924), .A2(n10044), .ZN(n9887) );
  NAND2_X1 U12523 ( .A1(n12921), .A2(n9887), .ZN(n14840) );
  INV_X1 U12524 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10013) );
  NAND2_X1 U12525 ( .A1(n14845), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9888) );
  INV_X1 U12526 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10137) );
  MUX2_X1 U12527 ( .A(n10137), .B(P2_REG1_REG_4__SCAN_IN), .S(n9889), .Z(
        n14854) );
  NAND2_X1 U12528 ( .A1(n14853), .A2(n14854), .ZN(n14852) );
  NAND2_X1 U12529 ( .A1(n14858), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9890) );
  NAND2_X1 U12530 ( .A1(n14852), .A2(n9890), .ZN(n12935) );
  INV_X1 U12531 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10356) );
  MUX2_X1 U12532 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10356), .S(n12933), .Z(
        n12936) );
  NAND2_X1 U12533 ( .A1(n12935), .A2(n12936), .ZN(n12934) );
  NAND2_X1 U12534 ( .A1(n12933), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9891) );
  NAND2_X1 U12535 ( .A1(n12934), .A2(n9891), .ZN(n12950) );
  INV_X1 U12536 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n15039) );
  MUX2_X1 U12537 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n15039), .S(n12945), .Z(
        n12951) );
  NAND2_X1 U12538 ( .A1(n12950), .A2(n12951), .ZN(n12949) );
  NAND2_X1 U12539 ( .A1(n12945), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9892) );
  NAND2_X1 U12540 ( .A1(n12949), .A2(n9892), .ZN(n12962) );
  INV_X1 U12541 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n15041) );
  MUX2_X1 U12542 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n15041), .S(n12957), .Z(
        n12963) );
  NAND2_X1 U12543 ( .A1(n12962), .A2(n12963), .ZN(n12961) );
  NAND2_X1 U12544 ( .A1(n12957), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9893) );
  NAND2_X1 U12545 ( .A1(n12961), .A2(n9893), .ZN(n14868) );
  INV_X1 U12546 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n15043) );
  MUX2_X1 U12547 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n15043), .S(n9894), .Z(
        n14867) );
  NAND2_X1 U12548 ( .A1(n9894), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9895) );
  INV_X1 U12549 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n11095) );
  MUX2_X1 U12550 ( .A(n11095), .B(P2_REG1_REG_9__SCAN_IN), .S(n9896), .Z(
        n14879) );
  NAND2_X1 U12551 ( .A1(n14887), .A2(n11095), .ZN(n9897) );
  OR2_X1 U12552 ( .A1(n9899), .A2(n9900), .ZN(n11283) );
  INV_X1 U12553 ( .A(n11283), .ZN(n9898) );
  AOI211_X1 U12554 ( .C1(n9900), .C2(n9899), .A(n14960), .B(n9898), .ZN(n9903)
         );
  NAND2_X1 U12555 ( .A1(n14971), .A2(n11292), .ZN(n9901) );
  NAND2_X1 U12556 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n10928)
         );
  OAI211_X1 U12557 ( .C1(n14988), .C2(n6789), .A(n9901), .B(n10928), .ZN(n9902) );
  OR3_X1 U12558 ( .A1(n9904), .A2(n9903), .A3(n9902), .ZN(P2_U3224) );
  CLKBUF_X2 U12559 ( .A(P1_U4016), .Z(n13814) );
  NOR2_X1 U12560 ( .A1(n14624), .A2(n13814), .ZN(P1_U3085) );
  XNOR2_X1 U12561 ( .A(n14729), .B(n13560), .ZN(n13517) );
  INV_X1 U12562 ( .A(n13517), .ZN(n9905) );
  OAI21_X1 U12563 ( .B1(n14730), .B2(n14807), .A(n9905), .ZN(n9906) );
  INV_X1 U12564 ( .A(n13487), .ZN(n13479) );
  NAND2_X1 U12565 ( .A1(n14728), .A2(n13479), .ZN(n10640) );
  OAI211_X1 U12566 ( .C1(n10506), .C2(n14725), .A(n9906), .B(n10640), .ZN(
        n9932) );
  NAND2_X1 U12567 ( .A1(n14810), .A2(n9932), .ZN(n9907) );
  OAI21_X1 U12568 ( .B1(n14810), .B2(n9165), .A(n9907), .ZN(P1_U3459) );
  OAI22_X1 U12569 ( .A1(n10094), .A2(P3_D_REG_0__SCAN_IN), .B1(n9909), .B2(
        n9908), .ZN(n9910) );
  INV_X1 U12570 ( .A(n9910), .ZN(P3_U3376) );
  INV_X1 U12571 ( .A(n12417), .ZN(n12406) );
  INV_X1 U12572 ( .A(SI_17_), .ZN(n9913) );
  INV_X1 U12573 ( .A(n9911), .ZN(n9912) );
  OAI222_X1 U12574 ( .A1(P3_U3151), .A2(n12406), .B1(n14433), .B2(n9913), .C1(
        n14434), .C2(n9912), .ZN(P3_U3278) );
  AND2_X1 U12575 ( .A1(n12916), .A2(n13194), .ZN(n9914) );
  NAND2_X1 U12576 ( .A1(n9914), .A2(n9915), .ZN(n9918) );
  INV_X1 U12577 ( .A(n9914), .ZN(n9917) );
  NAND2_X1 U12578 ( .A1(n9917), .A2(n9916), .ZN(n9954) );
  NAND2_X1 U12579 ( .A1(n9920), .A2(n9919), .ZN(n9921) );
  OAI21_X1 U12580 ( .B1(n9922), .B2(n9921), .A(n9955), .ZN(n9927) );
  INV_X1 U12581 ( .A(n12915), .ZN(n10129) );
  OAI22_X1 U12582 ( .A1(n10129), .A2(n12890), .B1(n12896), .B2(n9923), .ZN(
        n9926) );
  OAI22_X1 U12583 ( .A1(n12883), .A2(n10372), .B1(n9924), .B2(n10367), .ZN(
        n9925) );
  AOI211_X1 U12584 ( .C1(n12871), .C2(n9927), .A(n9926), .B(n9925), .ZN(n9928)
         );
  INV_X1 U12585 ( .A(n9928), .ZN(P2_U3209) );
  INV_X1 U12586 ( .A(n9929), .ZN(n9931) );
  INV_X1 U12587 ( .A(n11295), .ZN(n14898) );
  OAI222_X1 U12588 ( .A1(n13372), .A2(n9930), .B1(n13357), .B2(n9931), .C1(
        P2_U3088), .C2(n14898), .ZN(P2_U3316) );
  INV_X1 U12589 ( .A(n10728), .ZN(n10143) );
  OAI222_X1 U12590 ( .A1(n14318), .A2(n15329), .B1(n14312), .B2(n9931), .C1(
        P1_U3086), .C2(n10143), .ZN(P1_U3344) );
  INV_X1 U12591 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n14616) );
  NAND2_X1 U12592 ( .A1(n14822), .A2(n9932), .ZN(n9933) );
  OAI21_X1 U12593 ( .B1(n14822), .B2(n14616), .A(n9933), .ZN(P1_U3528) );
  AND2_X1 U12594 ( .A1(n9955), .A2(n9954), .ZN(n9947) );
  XNOR2_X1 U12595 ( .A(n10128), .B(n11592), .ZN(n9945) );
  NAND2_X1 U12596 ( .A1(n12915), .A2(n13194), .ZN(n9944) );
  XNOR2_X1 U12597 ( .A(n9945), .B(n9944), .ZN(n9953) );
  XNOR2_X1 U12598 ( .A(n9953), .B(n9947), .ZN(n9938) );
  AND2_X1 U12599 ( .A1(n9934), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12888) );
  INV_X1 U12600 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10429) );
  INV_X1 U12601 ( .A(n11613), .ZN(n12880) );
  INV_X1 U12602 ( .A(n12916), .ZN(n10162) );
  INV_X1 U12603 ( .A(n12914), .ZN(n10241) );
  OAI22_X1 U12604 ( .A1(n10162), .A2(n13139), .B1(n10241), .B2(n13141), .ZN(
        n10008) );
  AOI22_X1 U12605 ( .A1(n12880), .A2(n10008), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9935) );
  OAI21_X1 U12606 ( .B1(n10431), .B2(n12883), .A(n9935), .ZN(n9936) );
  AOI21_X1 U12607 ( .B1(n12888), .B2(n10429), .A(n9936), .ZN(n9937) );
  OAI21_X1 U12608 ( .B1(n9938), .B2(n12902), .A(n9937), .ZN(P2_U3190) );
  INV_X1 U12609 ( .A(n12432), .ZN(n12419) );
  INV_X1 U12610 ( .A(n9939), .ZN(n9940) );
  OAI222_X1 U12611 ( .A1(P3_U3151), .A2(n12419), .B1(n14433), .B2(n9941), .C1(
        n14434), .C2(n9940), .ZN(P3_U3277) );
  OAI222_X1 U12612 ( .A1(n14434), .A2(n9943), .B1(n14433), .B2(n9942), .C1(
        P3_U3151), .C2(n12428), .ZN(P3_U3276) );
  INV_X1 U12613 ( .A(n9944), .ZN(n9946) );
  AND2_X1 U12614 ( .A1(n9946), .A2(n9945), .ZN(n9956) );
  AOI21_X1 U12615 ( .B1(n9947), .B2(n9953), .A(n9956), .ZN(n9961) );
  XNOR2_X1 U12616 ( .A(n10240), .B(n11584), .ZN(n9948) );
  NAND2_X1 U12617 ( .A1(n12914), .A2(n13194), .ZN(n9949) );
  NAND2_X1 U12618 ( .A1(n9948), .A2(n9949), .ZN(n10024) );
  INV_X1 U12619 ( .A(n9948), .ZN(n9951) );
  INV_X1 U12620 ( .A(n9949), .ZN(n9950) );
  NAND2_X1 U12621 ( .A1(n9951), .A2(n9950), .ZN(n9952) );
  NAND2_X1 U12622 ( .A1(n10024), .A2(n9952), .ZN(n9957) );
  INV_X1 U12623 ( .A(n9957), .ZN(n9960) );
  NAND3_X1 U12624 ( .A1(n9955), .A2(n9954), .A3(n9953), .ZN(n9959) );
  NOR2_X1 U12625 ( .A1(n9957), .A2(n9956), .ZN(n9958) );
  NAND2_X1 U12626 ( .A1(n9959), .A2(n9958), .ZN(n10025) );
  OAI21_X1 U12627 ( .B1(n9961), .B2(n9960), .A(n10025), .ZN(n9962) );
  NAND2_X1 U12628 ( .A1(n9962), .A2(n12871), .ZN(n9966) );
  INV_X1 U12629 ( .A(n12913), .ZN(n10244) );
  OAI22_X1 U12630 ( .A1(n10129), .A2(n13139), .B1(n10244), .B2(n13141), .ZN(
        n10130) );
  INV_X1 U12631 ( .A(n10130), .ZN(n9963) );
  NAND2_X1 U12632 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n14863) );
  OAI21_X1 U12633 ( .B1(n11613), .B2(n9963), .A(n14863), .ZN(n9964) );
  AOI21_X1 U12634 ( .B1(n10240), .B2(n12900), .A(n9964), .ZN(n9965) );
  OAI211_X1 U12635 ( .C1(n12877), .C2(n10379), .A(n9966), .B(n9965), .ZN(
        P2_U3202) );
  INV_X1 U12636 ( .A(n10500), .ZN(n9967) );
  NAND2_X1 U12637 ( .A1(n13950), .A2(n9967), .ZN(n9991) );
  INV_X1 U12638 ( .A(n9968), .ZN(n9969) );
  NAND2_X1 U12639 ( .A1(n9989), .A2(n10494), .ZN(n10286) );
  AND2_X1 U12640 ( .A1(n10286), .A2(n10496), .ZN(n10737) );
  INV_X1 U12641 ( .A(n14729), .ZN(n14723) );
  INV_X1 U12642 ( .A(n9971), .ZN(n9973) );
  AOI22_X1 U12643 ( .A1(n11827), .A2(n13560), .B1(n9973), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n9972) );
  OAI21_X1 U12644 ( .B1(n11836), .B2(n14723), .A(n9972), .ZN(n9995) );
  NAND2_X1 U12645 ( .A1(n11827), .A2(n14729), .ZN(n9975) );
  NAND2_X1 U12646 ( .A1(n9973), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9974) );
  OAI211_X1 U12647 ( .C1(n11835), .C2(n14725), .A(n9975), .B(n9974), .ZN(n9996) );
  NAND2_X1 U12648 ( .A1(n11827), .A2(n9981), .ZN(n9979) );
  NAND2_X1 U12649 ( .A1(n11826), .A2(n9977), .ZN(n9978) );
  NAND2_X1 U12650 ( .A1(n9979), .A2(n9978), .ZN(n9980) );
  OAI22_X1 U12651 ( .A1(n11836), .A2(n9173), .B1(n14751), .B2(n11837), .ZN(
        n9982) );
  NOR2_X1 U12652 ( .A1(n9983), .A2(n9982), .ZN(n10049) );
  NOR2_X1 U12653 ( .A1(n9984), .A2(n10049), .ZN(n9985) );
  NAND2_X1 U12654 ( .A1(n9987), .A2(n14796), .ZN(n9988) );
  NAND2_X1 U12655 ( .A1(n9990), .A2(n14564), .ZN(n9994) );
  INV_X1 U12656 ( .A(n13765), .ZN(n10285) );
  NAND2_X1 U12657 ( .A1(n10737), .A2(n10285), .ZN(n10055) );
  INV_X1 U12658 ( .A(n13478), .ZN(n14734) );
  NAND2_X1 U12659 ( .A1(n13798), .A2(n13479), .ZN(n14722) );
  OAI21_X1 U12660 ( .B1(n14723), .B2(n14734), .A(n14722), .ZN(n9992) );
  AOI22_X1 U12661 ( .A1(n10055), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n14566), 
        .B2(n9992), .ZN(n9993) );
  OAI211_X1 U12662 ( .C1(n14751), .C2(n15382), .A(n9994), .B(n9993), .ZN(
        P1_U3222) );
  AOI22_X1 U12663 ( .A1(n14562), .A2(n13560), .B1(n10055), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n9998) );
  XOR2_X1 U12664 ( .A(n9996), .B(n9995), .Z(n13812) );
  NAND2_X1 U12665 ( .A1(n14564), .A2(n13812), .ZN(n9997) );
  OAI211_X1 U12666 ( .C1(n15388), .C2(n10640), .A(n9998), .B(n9997), .ZN(
        P1_U3232) );
  INV_X1 U12667 ( .A(n9999), .ZN(n10059) );
  AOI22_X1 U12668 ( .A1(n14655), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10390), .ZN(n10000) );
  OAI21_X1 U12669 ( .B1(n10059), .B2(n14312), .A(n10000), .ZN(P1_U3343) );
  OR2_X1 U12670 ( .A1(n9755), .A2(n10168), .ZN(n10001) );
  NAND2_X1 U12671 ( .A1(n10156), .A2(n10001), .ZN(n10035) );
  INV_X1 U12672 ( .A(n10036), .ZN(n10034) );
  NAND2_X1 U12673 ( .A1(n10035), .A2(n10034), .ZN(n10033) );
  NAND2_X1 U12674 ( .A1(n10162), .A2(n10372), .ZN(n10002) );
  NAND2_X1 U12675 ( .A1(n10033), .A2(n10002), .ZN(n10004) );
  NAND2_X1 U12676 ( .A1(n10004), .A2(n10003), .ZN(n10122) );
  OAI21_X1 U12677 ( .B1(n10004), .B2(n10003), .A(n10122), .ZN(n10005) );
  INV_X1 U12678 ( .A(n10005), .ZN(n10432) );
  NOR2_X1 U12679 ( .A1(n6445), .A2(n10010), .ZN(n10161) );
  NAND2_X1 U12680 ( .A1(n10160), .A2(n10161), .ZN(n10159) );
  OR2_X1 U12681 ( .A1(n9755), .A2(n10362), .ZN(n10006) );
  NAND2_X1 U12682 ( .A1(n10159), .A2(n10006), .ZN(n10037) );
  XNOR2_X1 U12683 ( .A(n10127), .B(n10126), .ZN(n10009) );
  AOI21_X1 U12684 ( .B1(n10009), .B2(n13228), .A(n10008), .ZN(n10427) );
  NAND2_X1 U12685 ( .A1(n10362), .A2(n10010), .ZN(n10166) );
  AOI211_X1 U12686 ( .C1(n10128), .C2(n10039), .A(n15030), .B(n10132), .ZN(
        n10435) );
  AOI21_X1 U12687 ( .B1(n15019), .B2(n10128), .A(n10435), .ZN(n10011) );
  OAI211_X1 U12688 ( .C1(n10432), .C2(n13327), .A(n10427), .B(n10011), .ZN(
        n10017) );
  NAND2_X1 U12689 ( .A1(n10017), .A2(n15047), .ZN(n10012) );
  OAI21_X1 U12690 ( .B1(n15047), .B2(n10013), .A(n10012), .ZN(P2_U3502) );
  INV_X1 U12691 ( .A(n10081), .ZN(n10014) );
  INV_X1 U12692 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15283) );
  NAND2_X1 U12693 ( .A1(n10017), .A2(n15026), .ZN(n10018) );
  OAI21_X1 U12694 ( .B1(n15026), .B2(n15283), .A(n10018), .ZN(P2_U3439) );
  XNOR2_X1 U12695 ( .A(n10350), .B(n6911), .ZN(n10019) );
  NAND2_X1 U12696 ( .A1(n12913), .A2(n13194), .ZN(n10020) );
  NAND2_X1 U12697 ( .A1(n10019), .A2(n10020), .ZN(n10061) );
  INV_X1 U12698 ( .A(n10019), .ZN(n10022) );
  INV_X1 U12699 ( .A(n10020), .ZN(n10021) );
  NAND2_X1 U12700 ( .A1(n10022), .A2(n10021), .ZN(n10023) );
  AND2_X1 U12701 ( .A1(n10061), .A2(n10023), .ZN(n10027) );
  OAI21_X1 U12702 ( .B1(n10027), .B2(n10026), .A(n10062), .ZN(n10031) );
  INV_X1 U12703 ( .A(n12912), .ZN(n10560) );
  OAI22_X1 U12704 ( .A1(n12877), .A2(n10345), .B1(n12890), .B2(n10560), .ZN(
        n10030) );
  NAND2_X1 U12705 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n12930) );
  NAND2_X1 U12706 ( .A1(n12900), .A2(n10350), .ZN(n10028) );
  OAI211_X1 U12707 ( .C1(n12896), .C2(n10241), .A(n12930), .B(n10028), .ZN(
        n10029) );
  AOI211_X1 U12708 ( .C1(n10031), .C2(n12871), .A(n10030), .B(n10029), .ZN(
        n10032) );
  INV_X1 U12709 ( .A(n10032), .ZN(P2_U3199) );
  OAI21_X1 U12710 ( .B1(n10035), .B2(n10034), .A(n10033), .ZN(n10374) );
  INV_X1 U12711 ( .A(n10374), .ZN(n10042) );
  XNOR2_X1 U12712 ( .A(n10036), .B(n10037), .ZN(n10038) );
  AOI222_X1 U12713 ( .A1(n13228), .A2(n10038), .B1(n9755), .B2(n13225), .C1(
        n12915), .C2(n13223), .ZN(n10376) );
  INV_X1 U12714 ( .A(n10039), .ZN(n10040) );
  OAI211_X1 U12715 ( .C1(n13327), .C2(n10042), .A(n10376), .B(n10041), .ZN(
        n10045) );
  NAND2_X1 U12716 ( .A1(n10045), .A2(n15047), .ZN(n10043) );
  OAI21_X1 U12717 ( .B1(n15047), .B2(n10044), .A(n10043), .ZN(P2_U3501) );
  INV_X1 U12718 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10047) );
  NAND2_X1 U12719 ( .A1(n10045), .A2(n15026), .ZN(n10046) );
  OAI21_X1 U12720 ( .B1(n15026), .B2(n10047), .A(n10046), .ZN(P2_U3436) );
  AOI22_X1 U12721 ( .A1(n11827), .A2(n13798), .B1(n11826), .B2(n14757), .ZN(
        n10048) );
  XNOR2_X1 U12722 ( .A(n10048), .B(n11838), .ZN(n10292) );
  OAI22_X1 U12723 ( .A1(n11836), .A2(n7185), .B1(n10058), .B2(n11837), .ZN(
        n10290) );
  XNOR2_X1 U12724 ( .A(n10292), .B(n10290), .ZN(n10052) );
  INV_X1 U12725 ( .A(n10049), .ZN(n10050) );
  NAND2_X1 U12726 ( .A1(n10051), .A2(n10052), .ZN(n13389) );
  OAI21_X1 U12727 ( .B1(n10052), .B2(n10051), .A(n13389), .ZN(n10053) );
  NAND2_X1 U12728 ( .A1(n10053), .A2(n14564), .ZN(n10057) );
  INV_X1 U12729 ( .A(n13797), .ZN(n10054) );
  OAI22_X1 U12730 ( .A1(n9173), .A2(n14734), .B1(n10054), .B2(n13487), .ZN(
        n10578) );
  AOI22_X1 U12731 ( .A1(n10055), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n14566), 
        .B2(n10578), .ZN(n10056) );
  OAI211_X1 U12732 ( .C1(n10058), .C2(n15382), .A(n10057), .B(n10056), .ZN(
        P1_U3237) );
  INV_X1 U12733 ( .A(n11297), .ZN(n14909) );
  OAI222_X1 U12734 ( .A1(n13372), .A2(n10060), .B1(n13357), .B2(n10059), .C1(
        n14909), .C2(P2_U3088), .ZN(P2_U3315) );
  XNOR2_X1 U12735 ( .A(n15001), .B(n6911), .ZN(n10311) );
  NAND2_X1 U12736 ( .A1(n12912), .A2(n13194), .ZN(n10312) );
  XNOR2_X1 U12737 ( .A(n10311), .B(n10312), .ZN(n10309) );
  XNOR2_X1 U12738 ( .A(n10309), .B(n10308), .ZN(n10069) );
  NAND2_X1 U12739 ( .A1(n12911), .A2(n13223), .ZN(n10064) );
  NAND2_X1 U12740 ( .A1(n12913), .A2(n13225), .ZN(n10063) );
  AND2_X1 U12741 ( .A1(n10064), .A2(n10063), .ZN(n10247) );
  INV_X1 U12742 ( .A(n10247), .ZN(n10065) );
  AOI22_X1 U12743 ( .A1(n12880), .A2(n10065), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10066) );
  OAI21_X1 U12744 ( .B1(n10252), .B2(n12877), .A(n10066), .ZN(n10067) );
  AOI21_X1 U12745 ( .B1(n15001), .B2(n12900), .A(n10067), .ZN(n10068) );
  OAI21_X1 U12746 ( .B1(n10069), .B2(n12902), .A(n10068), .ZN(P2_U3211) );
  INV_X1 U12747 ( .A(P3_U3897), .ZN(n12275) );
  INV_X1 U12748 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n10071) );
  NAND2_X1 U12749 ( .A1(n15143), .A2(n12285), .ZN(n10070) );
  OAI21_X1 U12750 ( .B1(n12285), .B2(n10071), .A(n10070), .ZN(P3_U3491) );
  INV_X1 U12751 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n10073) );
  NAND2_X1 U12752 ( .A1(n11993), .A2(n12285), .ZN(n10072) );
  OAI21_X1 U12753 ( .B1(n12285), .B2(n10073), .A(n10072), .ZN(P3_U3496) );
  INV_X1 U12754 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n10075) );
  NAND2_X1 U12755 ( .A1(n15123), .A2(n12285), .ZN(n10074) );
  OAI21_X1 U12756 ( .B1(n12285), .B2(n10075), .A(n10074), .ZN(P3_U3494) );
  INV_X1 U12757 ( .A(n10076), .ZN(n10178) );
  AOI22_X1 U12758 ( .A1(n11266), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10390), .ZN(n10077) );
  OAI21_X1 U12759 ( .B1(n10178), .B2(n14312), .A(n10077), .ZN(P1_U3342) );
  NAND2_X1 U12760 ( .A1(n10079), .A2(n10078), .ZN(n10080) );
  NOR2_X1 U12761 ( .A1(n10081), .A2(n10080), .ZN(n10082) );
  AND2_X1 U12762 ( .A1(n10082), .A2(n14994), .ZN(n10378) );
  INV_X1 U12763 ( .A(n10378), .ZN(n10083) );
  INV_X1 U12764 ( .A(n10250), .ZN(n10084) );
  NAND2_X1 U12765 ( .A1(n9771), .A2(n10084), .ZN(n10085) );
  OAI22_X1 U12766 ( .A1(n13219), .A2(n10087), .B1(n10086), .B2(n13217), .ZN(
        n10088) );
  AOI21_X1 U12767 ( .B1(n10089), .B2(n13219), .A(n10088), .ZN(n10092) );
  OAI21_X1 U12768 ( .B1(n13234), .B2(n13131), .A(n10167), .ZN(n10091) );
  OAI211_X1 U12769 ( .C1(n13236), .C2(n10093), .A(n10092), .B(n10091), .ZN(
        P2_U3265) );
  CLKBUF_X2 U12770 ( .A(n10094), .Z(n10120) );
  INV_X1 U12771 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10095) );
  NOR2_X1 U12772 ( .A1(n10120), .A2(n10095), .ZN(P3_U3245) );
  INV_X1 U12773 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10096) );
  NOR2_X1 U12774 ( .A1(n10120), .A2(n10096), .ZN(P3_U3242) );
  INV_X1 U12775 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10097) );
  NOR2_X1 U12776 ( .A1(n10120), .A2(n10097), .ZN(P3_U3235) );
  INV_X1 U12777 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10098) );
  NOR2_X1 U12778 ( .A1(n10120), .A2(n10098), .ZN(P3_U3244) );
  INV_X1 U12779 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10099) );
  NOR2_X1 U12780 ( .A1(n10120), .A2(n10099), .ZN(P3_U3246) );
  INV_X1 U12781 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10100) );
  NOR2_X1 U12782 ( .A1(n10120), .A2(n10100), .ZN(P3_U3252) );
  INV_X1 U12783 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10101) );
  NOR2_X1 U12784 ( .A1(n10120), .A2(n10101), .ZN(P3_U3238) );
  INV_X1 U12785 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10102) );
  NOR2_X1 U12786 ( .A1(n10120), .A2(n10102), .ZN(P3_U3250) );
  INV_X1 U12787 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10103) );
  NOR2_X1 U12788 ( .A1(n10120), .A2(n10103), .ZN(P3_U3234) );
  INV_X1 U12789 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10104) );
  NOR2_X1 U12790 ( .A1(n10120), .A2(n10104), .ZN(P3_U3237) );
  INV_X1 U12791 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10105) );
  NOR2_X1 U12792 ( .A1(n10120), .A2(n10105), .ZN(P3_U3257) );
  INV_X1 U12793 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10106) );
  NOR2_X1 U12794 ( .A1(n10120), .A2(n10106), .ZN(P3_U3255) );
  INV_X1 U12795 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10107) );
  NOR2_X1 U12796 ( .A1(n10120), .A2(n10107), .ZN(P3_U3241) );
  INV_X1 U12797 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10108) );
  NOR2_X1 U12798 ( .A1(n10120), .A2(n10108), .ZN(P3_U3240) );
  INV_X1 U12799 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10109) );
  NOR2_X1 U12800 ( .A1(n10120), .A2(n10109), .ZN(P3_U3239) );
  INV_X1 U12801 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10110) );
  NOR2_X1 U12802 ( .A1(n10120), .A2(n10110), .ZN(P3_U3253) );
  INV_X1 U12803 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10111) );
  NOR2_X1 U12804 ( .A1(n10120), .A2(n10111), .ZN(P3_U3251) );
  INV_X1 U12805 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10112) );
  NOR2_X1 U12806 ( .A1(n10120), .A2(n10112), .ZN(P3_U3236) );
  INV_X1 U12807 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10113) );
  NOR2_X1 U12808 ( .A1(n10120), .A2(n10113), .ZN(P3_U3254) );
  INV_X1 U12809 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10114) );
  NOR2_X1 U12810 ( .A1(n10120), .A2(n10114), .ZN(P3_U3263) );
  INV_X1 U12811 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10115) );
  NOR2_X1 U12812 ( .A1(n10120), .A2(n10115), .ZN(P3_U3262) );
  INV_X1 U12813 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10116) );
  NOR2_X1 U12814 ( .A1(n10120), .A2(n10116), .ZN(P3_U3256) );
  INV_X1 U12815 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10117) );
  NOR2_X1 U12816 ( .A1(n10120), .A2(n10117), .ZN(P3_U3261) );
  INV_X1 U12817 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10118) );
  NOR2_X1 U12818 ( .A1(n10120), .A2(n10118), .ZN(P3_U3243) );
  INV_X1 U12819 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10119) );
  NOR2_X1 U12820 ( .A1(n10120), .A2(n10119), .ZN(P3_U3248) );
  INV_X1 U12821 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n15224) );
  NOR2_X1 U12822 ( .A1(n10120), .A2(n15224), .ZN(P3_U3249) );
  NAND2_X1 U12823 ( .A1(n10129), .A2(n10431), .ZN(n10121) );
  NAND2_X1 U12824 ( .A1(n10122), .A2(n10121), .ZN(n10124) );
  INV_X1 U12825 ( .A(n10238), .ZN(n10123) );
  NAND2_X1 U12826 ( .A1(n10124), .A2(n10123), .ZN(n10237) );
  OAI21_X1 U12827 ( .B1(n10124), .B2(n10123), .A(n10237), .ZN(n10125) );
  INV_X1 U12828 ( .A(n10125), .ZN(n10385) );
  XNOR2_X1 U12829 ( .A(n10239), .B(n10238), .ZN(n10131) );
  AOI21_X1 U12830 ( .B1(n10131), .B2(n13228), .A(n10130), .ZN(n10377) );
  INV_X1 U12831 ( .A(n10132), .ZN(n10134) );
  INV_X1 U12832 ( .A(n10240), .ZN(n10380) );
  INV_X1 U12833 ( .A(n10344), .ZN(n10133) );
  AOI211_X1 U12834 ( .C1(n10240), .C2(n10134), .A(n15030), .B(n10133), .ZN(
        n10382) );
  AOI21_X1 U12835 ( .B1(n15019), .B2(n10240), .A(n10382), .ZN(n10135) );
  OAI211_X1 U12836 ( .C1(n10385), .C2(n13327), .A(n10377), .B(n10135), .ZN(
        n10175) );
  NAND2_X1 U12837 ( .A1(n10175), .A2(n15047), .ZN(n10136) );
  OAI21_X1 U12838 ( .B1(n15047), .B2(n10137), .A(n10136), .ZN(P2_U3503) );
  MUX2_X1 U12839 ( .A(n9295), .B(P1_REG1_REG_11__SCAN_IN), .S(n10728), .Z(
        n10142) );
  INV_X1 U12840 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10140) );
  AOI21_X1 U12841 ( .B1(n10146), .B2(n10139), .A(n10138), .ZN(n13873) );
  MUX2_X1 U12842 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n10140), .S(n10148), .Z(
        n13872) );
  NAND2_X1 U12843 ( .A1(n13873), .A2(n13872), .ZN(n13871) );
  OAI21_X1 U12844 ( .B1(n10140), .B2(n13875), .A(n13871), .ZN(n10141) );
  NOR2_X1 U12845 ( .A1(n10141), .A2(n10142), .ZN(n14653) );
  AOI21_X1 U12846 ( .B1(n10142), .B2(n10141), .A(n14653), .ZN(n10155) );
  NAND2_X1 U12847 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14568)
         );
  INV_X1 U12848 ( .A(n14568), .ZN(n10145) );
  NOR2_X1 U12849 ( .A1(n13924), .A2(n10143), .ZN(n10144) );
  AOI211_X1 U12850 ( .C1(n14624), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10145), 
        .B(n10144), .ZN(n10154) );
  NOR2_X1 U12851 ( .A1(n10146), .A2(n14690), .ZN(n13879) );
  MUX2_X1 U12852 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10147), .S(n10148), .Z(
        n13878) );
  OAI21_X1 U12853 ( .B1(n13880), .B2(n13879), .A(n13878), .ZN(n13882) );
  NAND2_X1 U12854 ( .A1(n10148), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10150) );
  MUX2_X1 U12855 ( .A(n9296), .B(P1_REG2_REG_11__SCAN_IN), .S(n10728), .Z(
        n10149) );
  AOI21_X1 U12856 ( .B1(n13882), .B2(n10150), .A(n10149), .ZN(n10723) );
  INV_X1 U12857 ( .A(n10723), .ZN(n10152) );
  NAND3_X1 U12858 ( .A1(n13882), .A2(n10150), .A3(n10149), .ZN(n10151) );
  NAND3_X1 U12859 ( .A1(n10152), .A2(n14656), .A3(n10151), .ZN(n10153) );
  OAI211_X1 U12860 ( .C1(n10155), .C2(n13799), .A(n10154), .B(n10153), .ZN(
        P1_U3254) );
  INV_X1 U12861 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10171) );
  INV_X1 U12862 ( .A(n10156), .ZN(n10157) );
  AOI21_X1 U12863 ( .B1(n10158), .B2(n10160), .A(n10157), .ZN(n10357) );
  OAI21_X1 U12864 ( .B1(n10161), .B2(n10160), .A(n10159), .ZN(n10165) );
  OAI22_X1 U12865 ( .A1(n10162), .A2(n13141), .B1(n7772), .B2(n13139), .ZN(
        n10164) );
  NOR2_X1 U12866 ( .A1(n10357), .A2(n9771), .ZN(n10163) );
  AOI211_X1 U12867 ( .C1(n13228), .C2(n10165), .A(n10164), .B(n10163), .ZN(
        n10366) );
  AOI21_X1 U12868 ( .B1(n10167), .B2(n10168), .A(n6936), .ZN(n10360) );
  AOI22_X1 U12869 ( .A1(n10360), .A2(n13291), .B1(n15019), .B2(n10168), .ZN(
        n10169) );
  OAI211_X1 U12870 ( .C1(n10357), .C2(n15023), .A(n10366), .B(n10169), .ZN(
        n10172) );
  NAND2_X1 U12871 ( .A1(n10172), .A2(n15026), .ZN(n10170) );
  OAI21_X1 U12872 ( .B1(n15026), .B2(n10171), .A(n10170), .ZN(P2_U3433) );
  NAND2_X1 U12873 ( .A1(n10172), .A2(n15047), .ZN(n10173) );
  OAI21_X1 U12874 ( .B1(n15047), .B2(n10174), .A(n10173), .ZN(P2_U3500) );
  INV_X1 U12875 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10177) );
  NAND2_X1 U12876 ( .A1(n10175), .A2(n15026), .ZN(n10176) );
  OAI21_X1 U12877 ( .B1(n15026), .B2(n10177), .A(n10176), .ZN(P2_U3442) );
  OAI222_X1 U12878 ( .A1(n13372), .A2(n10179), .B1(n13367), .B2(n10178), .C1(
        n6714), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U12879 ( .A(n10180), .ZN(n10183) );
  OAI222_X1 U12880 ( .A1(n14434), .A2(n10183), .B1(n14433), .B2(n10182), .C1(
        P3_U3151), .C2(n10181), .ZN(P3_U3275) );
  INV_X1 U12881 ( .A(n10201), .ZN(n10189) );
  INV_X1 U12882 ( .A(n10202), .ZN(n10184) );
  OR2_X1 U12883 ( .A1(n10208), .A2(n10184), .ZN(n10188) );
  AND3_X1 U12884 ( .A1(n10186), .A2(n10394), .A3(n10185), .ZN(n10187) );
  OAI211_X1 U12885 ( .C1(n10212), .C2(n10189), .A(n10188), .B(n10187), .ZN(
        n10190) );
  NAND2_X1 U12886 ( .A1(n10190), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10192) );
  OR2_X1 U12887 ( .A1(n10208), .A2(n10207), .ZN(n10191) );
  NOR2_X1 U12888 ( .A1(n12071), .A2(P3_U3151), .ZN(n10279) );
  NAND3_X1 U12889 ( .A1(n11622), .A2(n12126), .A3(n15148), .ZN(n10199) );
  OAI211_X1 U12890 ( .C1(n10200), .C2(n15147), .A(n10272), .B(n10199), .ZN(
        n10206) );
  NAND3_X1 U12891 ( .A1(n10212), .A2(n10201), .A3(n15138), .ZN(n10204) );
  NAND2_X1 U12892 ( .A1(n10208), .A2(n10202), .ZN(n10203) );
  NAND2_X1 U12893 ( .A1(n10204), .A2(n10203), .ZN(n10205) );
  NAND2_X1 U12894 ( .A1(n10206), .A2(n12041), .ZN(n10216) );
  INV_X1 U12895 ( .A(n10207), .ZN(n12269) );
  AND2_X1 U12896 ( .A1(n10208), .A2(n12269), .ZN(n10209) );
  INV_X1 U12897 ( .A(n10209), .ZN(n10211) );
  OR2_X1 U12898 ( .A1(n10212), .A2(n15140), .ZN(n10213) );
  AND2_X1 U12899 ( .A1(n10392), .A2(n15173), .ZN(n10266) );
  OAI22_X1 U12900 ( .A1(n12065), .A2(n10328), .B1(n12068), .B2(n15139), .ZN(
        n10214) );
  AOI21_X1 U12901 ( .B1(n12062), .B2(n15143), .A(n10214), .ZN(n10215) );
  OAI211_X1 U12902 ( .C1(n10279), .C2(n15155), .A(n10216), .B(n10215), .ZN(
        P3_U3162) );
  AOI22_X1 U12903 ( .A1(n12050), .A2(n15124), .B1(n12036), .B2(n10268), .ZN(
        n10219) );
  AND2_X1 U12904 ( .A1(n15143), .A2(n10284), .ZN(n12119) );
  NOR2_X1 U12905 ( .A1(n15141), .A2(n12119), .ZN(n12094) );
  INV_X1 U12906 ( .A(n12094), .ZN(n10217) );
  NAND2_X1 U12907 ( .A1(n12041), .A2(n10217), .ZN(n10218) );
  OAI211_X1 U12908 ( .C1(n10279), .C2(n10220), .A(n10219), .B(n10218), .ZN(
        P3_U3172) );
  INV_X1 U12909 ( .A(n14789), .ZN(n14784) );
  OAI21_X1 U12910 ( .B1(n10223), .B2(n10222), .A(n10221), .ZN(n10607) );
  AOI211_X1 U12911 ( .C1(n13394), .C2(n10580), .A(n14788), .B(n10488), .ZN(
        n10602) );
  NAND2_X1 U12912 ( .A1(n10607), .A2(n14793), .ZN(n10230) );
  OAI21_X1 U12913 ( .B1(n10225), .B2(n13576), .A(n10224), .ZN(n10228) );
  NAND2_X1 U12914 ( .A1(n13798), .A2(n13478), .ZN(n10227) );
  NAND2_X1 U12915 ( .A1(n13796), .A2(n13479), .ZN(n10226) );
  NAND2_X1 U12916 ( .A1(n10227), .A2(n10226), .ZN(n13393) );
  AOI21_X1 U12917 ( .B1(n10228), .B2(n14730), .A(n13393), .ZN(n10229) );
  NAND2_X1 U12918 ( .A1(n10230), .A2(n10229), .ZN(n10604) );
  AOI211_X1 U12919 ( .C1(n14784), .C2(n10607), .A(n10602), .B(n10604), .ZN(
        n10235) );
  OAI22_X1 U12920 ( .A1(n14282), .A2(n13578), .B1(n14810), .B2(n9184), .ZN(
        n10231) );
  INV_X1 U12921 ( .A(n10231), .ZN(n10232) );
  OAI21_X1 U12922 ( .B1(n10235), .B2(n14808), .A(n10232), .ZN(P1_U3468) );
  OAI22_X1 U12923 ( .A1(n14205), .A2(n13578), .B1(n14822), .B2(n9792), .ZN(
        n10233) );
  INV_X1 U12924 ( .A(n10233), .ZN(n10234) );
  OAI21_X1 U12925 ( .B1(n10235), .B2(n9605), .A(n10234), .ZN(P1_U3531) );
  NAND2_X1 U12926 ( .A1(n10380), .A2(n10241), .ZN(n10236) );
  XNOR2_X1 U12927 ( .A(n10553), .B(n6742), .ZN(n15005) );
  INV_X1 U12928 ( .A(n9771), .ZN(n11212) );
  NAND2_X1 U12929 ( .A1(n10239), .A2(n10238), .ZN(n10243) );
  NAND2_X1 U12930 ( .A1(n10241), .A2(n10240), .ZN(n10242) );
  NAND2_X1 U12931 ( .A1(n10243), .A2(n10242), .ZN(n10336) );
  NAND2_X1 U12932 ( .A1(n10336), .A2(n10333), .ZN(n10246) );
  NAND2_X1 U12933 ( .A1(n10350), .A2(n10244), .ZN(n10245) );
  NAND2_X1 U12934 ( .A1(n10246), .A2(n10245), .ZN(n10559) );
  XNOR2_X1 U12935 ( .A(n10559), .B(n6742), .ZN(n10248) );
  OAI21_X1 U12936 ( .B1(n10248), .B2(n13137), .A(n10247), .ZN(n10249) );
  AOI21_X1 U12937 ( .B1(n15005), .B2(n11212), .A(n10249), .ZN(n15007) );
  INV_X2 U12938 ( .A(n13219), .ZN(n13212) );
  NAND2_X1 U12939 ( .A1(n13219), .A2(n10250), .ZN(n13072) );
  INV_X1 U12940 ( .A(n13072), .ZN(n10908) );
  AND2_X1 U12941 ( .A1(n10342), .A2(n15001), .ZN(n10251) );
  OR2_X1 U12942 ( .A1(n10251), .A2(n10556), .ZN(n15003) );
  INV_X1 U12943 ( .A(n13131), .ZN(n12989) );
  OAI22_X1 U12944 ( .A1(n13219), .A2(n10253), .B1(n10252), .B2(n13217), .ZN(
        n10254) );
  AOI21_X1 U12945 ( .B1(n15001), .B2(n13234), .A(n10254), .ZN(n10255) );
  OAI21_X1 U12946 ( .B1(n15003), .B2(n12989), .A(n10255), .ZN(n10256) );
  AOI21_X1 U12947 ( .B1(n15005), .B2(n10908), .A(n10256), .ZN(n10257) );
  OAI21_X1 U12948 ( .B1(n15007), .B2(n13212), .A(n10257), .ZN(P2_U3259) );
  NOR3_X1 U12949 ( .A1(n12094), .A2(n15173), .A3(n10258), .ZN(n10259) );
  AOI21_X1 U12950 ( .B1(n15145), .B2(n15124), .A(n10259), .ZN(n10282) );
  INV_X1 U12951 ( .A(n10260), .ZN(n10263) );
  MUX2_X1 U12952 ( .A(n10263), .B(n10262), .S(n10261), .Z(n10264) );
  MUX2_X1 U12953 ( .A(n10411), .B(n10282), .S(n15159), .Z(n10270) );
  OR2_X1 U12954 ( .A1(n10267), .A2(n15140), .ZN(n11237) );
  AOI22_X1 U12955 ( .A1(n14499), .A2(n10268), .B1(n15136), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n10269) );
  NAND2_X1 U12956 ( .A1(n10270), .A2(n10269), .ZN(P3_U3233) );
  OAI21_X1 U12957 ( .B1(n10274), .B2(n10273), .A(n10325), .ZN(n10275) );
  NAND2_X1 U12958 ( .A1(n10275), .A2(n12041), .ZN(n10278) );
  INV_X1 U12959 ( .A(n15123), .ZN(n10987) );
  OAI22_X1 U12960 ( .A1(n12065), .A2(n10987), .B1(n12068), .B2(n15131), .ZN(
        n10276) );
  AOI21_X1 U12961 ( .B1(n12062), .B2(n15124), .A(n10276), .ZN(n10277) );
  OAI211_X1 U12962 ( .C1(n10279), .C2(n10710), .A(n10278), .B(n10277), .ZN(
        P3_U3177) );
  INV_X1 U12963 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10280) );
  MUX2_X1 U12964 ( .A(n10280), .B(n10282), .S(n15206), .Z(n10281) );
  OAI21_X1 U12965 ( .B1(n10284), .B2(n12776), .A(n10281), .ZN(P3_U3390) );
  MUX2_X1 U12966 ( .A(n12287), .B(n10282), .S(n15222), .Z(n10283) );
  OAI21_X1 U12967 ( .B1(n10284), .B2(n12722), .A(n10283), .ZN(P3_U3459) );
  NAND3_X1 U12968 ( .A1(n10286), .A2(n10285), .A3(n9971), .ZN(n10287) );
  NAND2_X1 U12969 ( .A1(n10287), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10288) );
  AOI22_X1 U12970 ( .A1(n11831), .A2(n13797), .B1(n11827), .B2(n13394), .ZN(
        n10293) );
  NAND2_X1 U12971 ( .A1(n11826), .A2(n13394), .ZN(n10289) );
  XNOR2_X1 U12972 ( .A(n10293), .B(n10295), .ZN(n13391) );
  INV_X1 U12973 ( .A(n10290), .ZN(n10291) );
  NAND2_X1 U12974 ( .A1(n10292), .A2(n10291), .ZN(n13388) );
  INV_X1 U12975 ( .A(n10293), .ZN(n10294) );
  NAND2_X1 U12976 ( .A1(n10295), .A2(n10294), .ZN(n10296) );
  AOI22_X1 U12977 ( .A1(n11831), .A2(n13796), .B1(n13583), .B2(n11827), .ZN(
        n10297) );
  INV_X1 U12978 ( .A(n10526), .ZN(n10298) );
  NAND2_X1 U12979 ( .A1(n10298), .A2(n10528), .ZN(n10300) );
  AOI22_X1 U12980 ( .A1(n13583), .A2(n11826), .B1(n11827), .B2(n13796), .ZN(
        n10299) );
  XOR2_X1 U12981 ( .A(n11838), .B(n10299), .Z(n10527) );
  XNOR2_X1 U12982 ( .A(n10300), .B(n10527), .ZN(n10301) );
  NAND2_X1 U12983 ( .A1(n10301), .A2(n14564), .ZN(n10307) );
  NOR2_X1 U12984 ( .A1(n10507), .A2(n14796), .ZN(n14765) );
  NAND2_X1 U12985 ( .A1(n13797), .A2(n13478), .ZN(n10303) );
  NAND2_X1 U12986 ( .A1(n13795), .A2(n13479), .ZN(n10302) );
  AND2_X1 U12987 ( .A1(n10303), .A2(n10302), .ZN(n10490) );
  INV_X1 U12988 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n10304) );
  OAI22_X1 U12989 ( .A1(n15388), .A2(n10490), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10304), .ZN(n10305) );
  AOI21_X1 U12990 ( .B1(n10737), .B2(n14765), .A(n10305), .ZN(n10306) );
  OAI211_X1 U12991 ( .C1(n15385), .C2(n10497), .A(n10307), .B(n10306), .ZN(
        P1_U3230) );
  INV_X1 U12992 ( .A(n10309), .ZN(n10310) );
  INV_X1 U12993 ( .A(n10311), .ZN(n10314) );
  INV_X1 U12994 ( .A(n10312), .ZN(n10313) );
  NAND2_X1 U12995 ( .A1(n10314), .A2(n10313), .ZN(n10315) );
  XNOR2_X1 U12996 ( .A(n10872), .B(n11592), .ZN(n10518) );
  NAND2_X1 U12997 ( .A1(n12911), .A2(n13194), .ZN(n10516) );
  XNOR2_X1 U12998 ( .A(n10518), .B(n10516), .ZN(n10514) );
  XOR2_X1 U12999 ( .A(n10515), .B(n10514), .Z(n10320) );
  INV_X1 U13000 ( .A(n10872), .ZN(n15010) );
  AOI22_X1 U13001 ( .A1(n12848), .A2(n12910), .B1(n12847), .B2(n12912), .ZN(
        n10318) );
  INV_X1 U13002 ( .A(n10316), .ZN(n10570) );
  AOI22_X1 U13003 ( .A1(n12888), .A2(n10570), .B1(P2_REG3_REG_7__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10317) );
  OAI211_X1 U13004 ( .C1(n15010), .C2(n12883), .A(n10318), .B(n10317), .ZN(
        n10319) );
  AOI21_X1 U13005 ( .B1(n10320), .B2(n12871), .A(n10319), .ZN(n10321) );
  INV_X1 U13006 ( .A(n10321), .ZN(P2_U3185) );
  INV_X1 U13007 ( .A(n12071), .ZN(n12028) );
  INV_X1 U13008 ( .A(n10322), .ZN(n10323) );
  NAND2_X1 U13009 ( .A1(n10323), .A2(n10328), .ZN(n10324) );
  AND2_X1 U13010 ( .A1(n10325), .A2(n10324), .ZN(n10327) );
  XNOR2_X1 U13011 ( .A(n10986), .B(n15123), .ZN(n10326) );
  OAI211_X1 U13012 ( .C1(n10327), .C2(n10326), .A(n12041), .B(n10985), .ZN(
        n10332) );
  NOR2_X1 U13013 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15117), .ZN(n10678) );
  INV_X1 U13014 ( .A(n12062), .ZN(n12052) );
  INV_X1 U13015 ( .A(n15108), .ZN(n10988) );
  OAI22_X1 U13016 ( .A1(n12052), .A2(n10328), .B1(n10988), .B2(n12065), .ZN(
        n10329) );
  AOI211_X1 U13017 ( .C1(n12036), .C2(n10330), .A(n10678), .B(n10329), .ZN(
        n10331) );
  OAI211_X1 U13018 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12028), .A(n10332), .B(
        n10331), .ZN(P3_U3158) );
  INV_X1 U13019 ( .A(n10333), .ZN(n10335) );
  XNOR2_X1 U13020 ( .A(n10334), .B(n10335), .ZN(n10337) );
  INV_X1 U13021 ( .A(n10337), .ZN(n10354) );
  XNOR2_X1 U13022 ( .A(n10336), .B(n10335), .ZN(n10340) );
  NAND2_X1 U13023 ( .A1(n10337), .A2(n11212), .ZN(n10339) );
  AOI22_X1 U13024 ( .A1(n13225), .A2(n12914), .B1(n12912), .B2(n13223), .ZN(
        n10338) );
  OAI211_X1 U13025 ( .C1(n13137), .C2(n10340), .A(n10339), .B(n10338), .ZN(
        n10349) );
  MUX2_X1 U13026 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10349), .S(n13219), .Z(
        n10341) );
  INV_X1 U13027 ( .A(n10341), .ZN(n10348) );
  INV_X1 U13028 ( .A(n10342), .ZN(n10343) );
  AOI21_X1 U13029 ( .B1(n10350), .B2(n10344), .A(n10343), .ZN(n10351) );
  OAI22_X1 U13030 ( .A1(n13147), .A2(n6939), .B1(n13217), .B2(n10345), .ZN(
        n10346) );
  AOI21_X1 U13031 ( .B1(n10351), .B2(n13131), .A(n10346), .ZN(n10347) );
  OAI211_X1 U13032 ( .C1(n10354), .C2(n13072), .A(n10348), .B(n10347), .ZN(
        P2_U3260) );
  INV_X1 U13033 ( .A(n10349), .ZN(n10353) );
  AOI22_X1 U13034 ( .A1(n10351), .A2(n13291), .B1(n15019), .B2(n10350), .ZN(
        n10352) );
  OAI211_X1 U13035 ( .C1(n15023), .C2(n10354), .A(n10353), .B(n10352), .ZN(
        n10386) );
  NAND2_X1 U13036 ( .A1(n10386), .A2(n15047), .ZN(n10355) );
  OAI21_X1 U13037 ( .B1(n15047), .B2(n10356), .A(n10355), .ZN(P2_U3504) );
  INV_X1 U13038 ( .A(n10357), .ZN(n10364) );
  OAI22_X1 U13039 ( .A1(n13219), .A2(n10358), .B1(n7777), .B2(n13217), .ZN(
        n10359) );
  AOI21_X1 U13040 ( .B1(n10360), .B2(n13131), .A(n10359), .ZN(n10361) );
  OAI21_X1 U13041 ( .B1(n10362), .B2(n13147), .A(n10361), .ZN(n10363) );
  AOI21_X1 U13042 ( .B1(n10364), .B2(n10908), .A(n10363), .ZN(n10365) );
  OAI21_X1 U13043 ( .B1(n10366), .B2(n13212), .A(n10365), .ZN(P2_U3264) );
  INV_X1 U13044 ( .A(n13236), .ZN(n13023) );
  OAI22_X1 U13045 ( .A1(n13219), .A2(n10368), .B1(n10367), .B2(n13217), .ZN(
        n10369) );
  AOI21_X1 U13046 ( .B1(n10370), .B2(n13131), .A(n10369), .ZN(n10371) );
  OAI21_X1 U13047 ( .B1(n10372), .B2(n13147), .A(n10371), .ZN(n10373) );
  AOI21_X1 U13048 ( .B1(n13023), .B2(n10374), .A(n10373), .ZN(n10375) );
  OAI21_X1 U13049 ( .B1(n10376), .B2(n13212), .A(n10375), .ZN(P2_U3263) );
  MUX2_X1 U13050 ( .A(n9871), .B(n10377), .S(n13219), .Z(n10384) );
  AND2_X1 U13051 ( .A1(n10378), .A2(n13230), .ZN(n13175) );
  OAI22_X1 U13052 ( .A1(n13147), .A2(n10380), .B1(n13217), .B2(n10379), .ZN(
        n10381) );
  AOI21_X1 U13053 ( .B1(n10382), .B2(n13175), .A(n10381), .ZN(n10383) );
  OAI211_X1 U13054 ( .C1(n13236), .C2(n10385), .A(n10384), .B(n10383), .ZN(
        P2_U3261) );
  INV_X1 U13055 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10388) );
  NAND2_X1 U13056 ( .A1(n10386), .A2(n15026), .ZN(n10387) );
  OAI21_X1 U13057 ( .B1(n15026), .B2(n10388), .A(n10387), .ZN(P2_U3445) );
  INV_X1 U13058 ( .A(n10389), .ZN(n10511) );
  AOI22_X1 U13059 ( .A1(n13894), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10390), .ZN(n10391) );
  OAI21_X1 U13060 ( .B1(n10511), .B2(n14312), .A(n10391), .ZN(P1_U3341) );
  INV_X1 U13061 ( .A(n10392), .ZN(n10393) );
  OR2_X1 U13062 ( .A1(n10394), .A2(P3_U3151), .ZN(n12273) );
  NAND2_X1 U13063 ( .A1(n10393), .A2(n12273), .ZN(n10419) );
  NAND2_X1 U13064 ( .A1(n12260), .A2(n10394), .ZN(n10396) );
  AND2_X1 U13065 ( .A1(n10396), .A2(n10395), .ZN(n10417) );
  INV_X1 U13066 ( .A(n10397), .ZN(n10398) );
  INV_X1 U13067 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n12289) );
  NAND2_X1 U13068 ( .A1(n12289), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10399) );
  NAND2_X1 U13069 ( .A1(n10414), .A2(n10399), .ZN(n10400) );
  NAND2_X1 U13070 ( .A1(n10404), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10451) );
  NAND2_X1 U13071 ( .A1(n10400), .A2(n10451), .ZN(n10401) );
  INV_X1 U13072 ( .A(n10401), .ZN(n10402) );
  OR2_X1 U13073 ( .A1(n10401), .A2(n10413), .ZN(n10452) );
  OAI21_X1 U13074 ( .B1(n10402), .B2(P3_REG2_REG_1__SCAN_IN), .A(n10452), .ZN(
        n10424) );
  NAND2_X1 U13075 ( .A1(n12289), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10403) );
  NAND2_X1 U13076 ( .A1(n10414), .A2(n10403), .ZN(n10405) );
  NAND2_X1 U13077 ( .A1(n10404), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n10442) );
  NAND2_X1 U13078 ( .A1(n10405), .A2(n10442), .ZN(n10406) );
  NAND2_X1 U13079 ( .A1(n10406), .A2(n10412), .ZN(n10410) );
  INV_X1 U13080 ( .A(n10407), .ZN(n10409) );
  AOI21_X1 U13081 ( .B1(n10443), .B2(n10410), .A(n15097), .ZN(n10423) );
  MUX2_X1 U13082 ( .A(n10411), .B(n12287), .S(n6446), .Z(n12286) );
  NAND2_X1 U13083 ( .A1(n12286), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n12292) );
  NAND2_X1 U13084 ( .A1(n10415), .A2(n10414), .ZN(n10467) );
  OAI21_X1 U13085 ( .B1(n10415), .B2(n10414), .A(n10467), .ZN(n10416) );
  NOR2_X1 U13086 ( .A1(n10416), .A2(n12292), .ZN(n10717) );
  AOI21_X1 U13087 ( .B1(n12292), .B2(n10416), .A(n10717), .ZN(n10421) );
  NAND2_X1 U13088 ( .A1(n12285), .A2(n9031), .ZN(n15074) );
  INV_X1 U13089 ( .A(n10417), .ZN(n10418) );
  AND2_X1 U13090 ( .A1(n10419), .A2(n10418), .ZN(n15087) );
  AOI22_X1 U13091 ( .A1(n15087), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10420) );
  OAI21_X1 U13092 ( .B1(n10421), .B2(n15074), .A(n10420), .ZN(n10422) );
  AOI211_X1 U13093 ( .C1(n15089), .C2(n10424), .A(n10423), .B(n10422), .ZN(
        n10425) );
  OAI21_X1 U13094 ( .B1(n10426), .B2(n15068), .A(n10425), .ZN(P3_U3183) );
  INV_X1 U13095 ( .A(n13217), .ZN(n13209) );
  INV_X1 U13096 ( .A(n10427), .ZN(n10428) );
  AOI21_X1 U13097 ( .B1(n13209), .B2(n10429), .A(n10428), .ZN(n10437) );
  OAI22_X1 U13098 ( .A1(n13147), .A2(n10431), .B1(n10430), .B2(n13219), .ZN(
        n10434) );
  NOR2_X1 U13099 ( .A1(n10432), .A2(n13236), .ZN(n10433) );
  AOI211_X1 U13100 ( .C1(n10435), .C2(n13175), .A(n10434), .B(n10433), .ZN(
        n10436) );
  OAI21_X1 U13101 ( .B1(n13212), .B2(n10437), .A(n10436), .ZN(P2_U3262) );
  INV_X1 U13102 ( .A(SI_21_), .ZN(n10440) );
  INV_X1 U13103 ( .A(n10438), .ZN(n10439) );
  OAI222_X1 U13104 ( .A1(P3_U3151), .A2(n10441), .B1(n14433), .B2(n10440), 
        .C1(n14434), .C2(n10439), .ZN(P3_U3274) );
  INV_X1 U13105 ( .A(n10624), .ZN(n10612) );
  NAND2_X1 U13106 ( .A1(n10443), .A2(n10442), .ZN(n10706) );
  NAND2_X1 U13107 ( .A1(n10722), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10444) );
  INV_X1 U13108 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15210) );
  MUX2_X1 U13109 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n15210), .S(n10624), .Z(
        n10447) );
  NAND2_X1 U13110 ( .A1(n10446), .A2(n10447), .ZN(n10626) );
  NOR2_X1 U13111 ( .A1(n10448), .A2(n10447), .ZN(n10449) );
  NAND2_X1 U13112 ( .A1(n10676), .A2(n10449), .ZN(n10450) );
  AND2_X1 U13113 ( .A1(n10626), .A2(n10450), .ZN(n10466) );
  NAND2_X1 U13114 ( .A1(n10452), .A2(n10451), .ZN(n10703) );
  NAND2_X1 U13115 ( .A1(n10722), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10453) );
  NAND2_X1 U13116 ( .A1(n10454), .A2(n10477), .ZN(n10457) );
  OAI21_X1 U13117 ( .B1(n10454), .B2(n10477), .A(n10457), .ZN(n10670) );
  NAND2_X1 U13118 ( .A1(n10672), .A2(n10457), .ZN(n10456) );
  INV_X1 U13119 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10455) );
  MUX2_X1 U13120 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n10455), .S(n10624), .Z(
        n10458) );
  NAND2_X1 U13121 ( .A1(n10456), .A2(n10458), .ZN(n10620) );
  INV_X1 U13122 ( .A(n10457), .ZN(n10459) );
  NOR2_X1 U13123 ( .A1(n10459), .A2(n10458), .ZN(n10460) );
  NAND2_X1 U13124 ( .A1(n10672), .A2(n10460), .ZN(n10461) );
  NAND2_X1 U13125 ( .A1(n10620), .A2(n10461), .ZN(n10462) );
  NAND2_X1 U13126 ( .A1(n15089), .A2(n10462), .ZN(n10465) );
  NOR2_X1 U13127 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10463), .ZN(n11992) );
  AOI21_X1 U13128 ( .B1(n15087), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n11992), .ZN(
        n10464) );
  OAI211_X1 U13129 ( .C1(n10466), .C2(n15097), .A(n10465), .B(n10464), .ZN(
        n10486) );
  INV_X1 U13130 ( .A(n10467), .ZN(n10716) );
  MUX2_X1 U13131 ( .A(n10469), .B(n10468), .S(n6446), .Z(n10471) );
  INV_X1 U13132 ( .A(n10722), .ZN(n10470) );
  NAND2_X1 U13133 ( .A1(n10471), .A2(n10470), .ZN(n10685) );
  INV_X1 U13134 ( .A(n10471), .ZN(n10472) );
  NAND2_X1 U13135 ( .A1(n10472), .A2(n10722), .ZN(n10473) );
  MUX2_X1 U13136 ( .A(n10475), .B(n10474), .S(n6446), .Z(n10476) );
  INV_X1 U13137 ( .A(n10477), .ZN(n10683) );
  NAND2_X1 U13138 ( .A1(n10476), .A2(n10683), .ZN(n10480) );
  INV_X1 U13139 ( .A(n10476), .ZN(n10478) );
  NAND2_X1 U13140 ( .A1(n10478), .A2(n10477), .ZN(n10479) );
  NAND2_X1 U13141 ( .A1(n10480), .A2(n10479), .ZN(n10684) );
  INV_X1 U13142 ( .A(n10480), .ZN(n10481) );
  NOR2_X1 U13143 ( .A1(n10687), .A2(n10481), .ZN(n10483) );
  MUX2_X1 U13144 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n6446), .Z(n10609) );
  XNOR2_X1 U13145 ( .A(n10609), .B(n10624), .ZN(n10482) );
  AOI21_X1 U13146 ( .B1(n10483), .B2(n10482), .A(n10610), .ZN(n10484) );
  NOR2_X1 U13147 ( .A1(n10484), .A2(n15074), .ZN(n10485) );
  AOI211_X1 U13148 ( .C1(n15084), .C2(n10612), .A(n10486), .B(n10485), .ZN(
        n10487) );
  INV_X1 U13149 ( .A(n10487), .ZN(P3_U3186) );
  INV_X1 U13150 ( .A(n14788), .ZN(n14715) );
  OAI211_X1 U13151 ( .C1(n10488), .C2(n10507), .A(n10590), .B(n14715), .ZN(
        n14766) );
  AOI21_X1 U13152 ( .B1(n10489), .B2(n13519), .A(n14704), .ZN(n10493) );
  INV_X1 U13153 ( .A(n10490), .ZN(n10491) );
  AOI21_X1 U13154 ( .B1(n10493), .B2(n10492), .A(n10491), .ZN(n14768) );
  INV_X1 U13155 ( .A(n10494), .ZN(n10495) );
  INV_X1 U13156 ( .A(n14708), .ZN(n14737) );
  INV_X1 U13157 ( .A(n10497), .ZN(n10498) );
  NAND2_X1 U13158 ( .A1(n14737), .A2(n10498), .ZN(n10499) );
  OAI211_X1 U13159 ( .C1(n14082), .C2(n14766), .A(n14768), .B(n10499), .ZN(
        n10503) );
  NOR2_X1 U13160 ( .A1(n10501), .A2(n10500), .ZN(n13954) );
  NAND2_X1 U13161 ( .A1(n13954), .A2(n10582), .ZN(n10502) );
  MUX2_X1 U13162 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10503), .S(n14691), .Z(
        n10509) );
  OAI21_X1 U13163 ( .B1(n6604), .B2(n13519), .A(n10504), .ZN(n14764) );
  OR2_X1 U13164 ( .A1(n10506), .A2(n9590), .ZN(n14453) );
  OAI22_X1 U13165 ( .A1(n14764), .A2(n14461), .B1(n10507), .B2(n14739), .ZN(
        n10508) );
  OR2_X1 U13166 ( .A1(n10509), .A2(n10508), .ZN(P1_U3289) );
  INV_X1 U13167 ( .A(n14944), .ZN(n10512) );
  OAI222_X1 U13168 ( .A1(P2_U3088), .A2(n10512), .B1(n13367), .B2(n10511), 
        .C1(n10510), .C2(n13372), .ZN(P2_U3313) );
  AND2_X1 U13169 ( .A1(n12910), .A2(n13194), .ZN(n10776) );
  XNOR2_X1 U13170 ( .A(n15018), .B(n11592), .ZN(n10775) );
  AND2_X1 U13171 ( .A1(n10775), .A2(n10776), .ZN(n10774) );
  INV_X1 U13172 ( .A(n10774), .ZN(n10513) );
  OAI21_X1 U13173 ( .B1(n10776), .B2(n10775), .A(n10513), .ZN(n10521) );
  NAND2_X1 U13174 ( .A1(n10515), .A2(n10514), .ZN(n10520) );
  INV_X1 U13175 ( .A(n10516), .ZN(n10517) );
  NAND2_X1 U13176 ( .A1(n10518), .A2(n10517), .ZN(n10519) );
  XOR2_X1 U13177 ( .A(n10521), .B(n10777), .Z(n10525) );
  AOI22_X1 U13178 ( .A1(n12847), .A2(n12911), .B1(n12848), .B2(n12909), .ZN(
        n10522) );
  NAND2_X1 U13179 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n14876) );
  OAI211_X1 U13180 ( .C1(n10923), .C2(n12877), .A(n10522), .B(n14876), .ZN(
        n10523) );
  AOI21_X1 U13181 ( .B1(n15018), .B2(n12900), .A(n10523), .ZN(n10524) );
  OAI21_X1 U13182 ( .B1(n10525), .B2(n12902), .A(n10524), .ZN(P2_U3193) );
  NAND2_X1 U13183 ( .A1(n13590), .A2(n11826), .ZN(n10530) );
  NAND2_X1 U13184 ( .A1(n11827), .A2(n13795), .ZN(n10529) );
  NAND2_X1 U13185 ( .A1(n10530), .A2(n10529), .ZN(n10531) );
  XNOR2_X1 U13186 ( .A(n10531), .B(n6473), .ZN(n10535) );
  INV_X1 U13187 ( .A(n10535), .ZN(n10533) );
  AOI22_X1 U13188 ( .A1(n11831), .A2(n13795), .B1(n13590), .B2(n11827), .ZN(
        n10534) );
  INV_X1 U13189 ( .A(n10534), .ZN(n10532) );
  NAND2_X1 U13190 ( .A1(n10533), .A2(n10532), .ZN(n10546) );
  INV_X1 U13191 ( .A(n10546), .ZN(n10536) );
  AND2_X1 U13192 ( .A1(n10535), .A2(n10534), .ZN(n10545) );
  NOR2_X1 U13193 ( .A1(n10536), .A2(n10545), .ZN(n10537) );
  XNOR2_X1 U13194 ( .A(n10547), .B(n10537), .ZN(n10538) );
  NAND2_X1 U13195 ( .A1(n10538), .A2(n14564), .ZN(n10544) );
  AND2_X1 U13196 ( .A1(n13590), .A2(n14758), .ZN(n14771) );
  OR2_X1 U13197 ( .A1(n13593), .A2(n13487), .ZN(n10540) );
  NAND2_X1 U13198 ( .A1(n13796), .A2(n13478), .ZN(n10539) );
  AND2_X1 U13199 ( .A1(n10540), .A2(n10539), .ZN(n14774) );
  OAI21_X1 U13200 ( .B1(n15388), .B2(n14774), .A(n10541), .ZN(n10542) );
  AOI21_X1 U13201 ( .B1(n10737), .B2(n14771), .A(n10542), .ZN(n10543) );
  OAI211_X1 U13202 ( .C1(n15385), .C2(n10592), .A(n10544), .B(n10543), .ZN(
        P1_U3227) );
  OAI22_X1 U13203 ( .A1(n14779), .A2(n11837), .B1(n13593), .B2(n11836), .ZN(
        n10738) );
  OAI22_X1 U13204 ( .A1(n14779), .A2(n11835), .B1(n13593), .B2(n11837), .ZN(
        n10548) );
  XNOR2_X1 U13205 ( .A(n10548), .B(n11838), .ZN(n10739) );
  XOR2_X1 U13206 ( .A(n10738), .B(n10739), .Z(n10549) );
  OAI211_X1 U13207 ( .C1(n6605), .C2(n10549), .A(n10740), .B(n14564), .ZN(
        n10552) );
  AOI22_X1 U13208 ( .A1(n13793), .A2(n13479), .B1(n13478), .B2(n13795), .ZN(
        n14703) );
  INV_X1 U13209 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n13842) );
  OAI22_X1 U13210 ( .A1(n15388), .A2(n14703), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13842), .ZN(n10550) );
  AOI21_X1 U13211 ( .B1(n14562), .B2(n13594), .A(n10550), .ZN(n10551) );
  OAI211_X1 U13212 ( .C1(n15385), .C2(n14707), .A(n10552), .B(n10551), .ZN(
        P1_U3239) );
  NAND2_X1 U13213 ( .A1(n15001), .A2(n12912), .ZN(n10554) );
  OAI21_X1 U13214 ( .B1(n10555), .B2(n10563), .A(n10868), .ZN(n15009) );
  OR2_X1 U13215 ( .A1(n15010), .A2(n10556), .ZN(n10557) );
  NAND2_X1 U13216 ( .A1(n10922), .A2(n10557), .ZN(n15011) );
  INV_X1 U13217 ( .A(n15011), .ZN(n10568) );
  NAND2_X1 U13218 ( .A1(n10559), .A2(n10558), .ZN(n10562) );
  NAND2_X1 U13219 ( .A1(n15001), .A2(n10560), .ZN(n10561) );
  INV_X1 U13220 ( .A(n10563), .ZN(n10564) );
  XNOR2_X1 U13221 ( .A(n10874), .B(n10564), .ZN(n10565) );
  NAND2_X1 U13222 ( .A1(n10565), .A2(n13228), .ZN(n10567) );
  AOI22_X1 U13223 ( .A1(n13223), .A2(n12910), .B1(n12912), .B2(n13225), .ZN(
        n10566) );
  NAND2_X1 U13224 ( .A1(n10567), .A2(n10566), .ZN(n15012) );
  AOI21_X1 U13225 ( .B1(n11580), .B2(n10568), .A(n15012), .ZN(n10569) );
  MUX2_X1 U13226 ( .A(n9876), .B(n10569), .S(n13219), .Z(n10572) );
  AOI22_X1 U13227 ( .A1(n10872), .A2(n13234), .B1(n13209), .B2(n10570), .ZN(
        n10571) );
  OAI211_X1 U13228 ( .C1(n13236), .C2(n15009), .A(n10572), .B(n10571), .ZN(
        P2_U3258) );
  INV_X2 U13229 ( .A(n14691), .ZN(n14710) );
  OR2_X1 U13230 ( .A1(n13564), .A2(n13929), .ZN(n13556) );
  NOR2_X1 U13231 ( .A1(n14710), .A2(n13556), .ZN(n14743) );
  NOR2_X1 U13232 ( .A1(n14710), .A2(n10573), .ZN(n10574) );
  OR2_X1 U13233 ( .A1(n14743), .A2(n10574), .ZN(n14042) );
  INV_X1 U13234 ( .A(n14042), .ZN(n10770) );
  XNOR2_X1 U13235 ( .A(n10575), .B(n13569), .ZN(n14761) );
  OAI21_X1 U13236 ( .B1(n13569), .B2(n10577), .A(n10576), .ZN(n10579) );
  AOI21_X1 U13237 ( .B1(n10579), .B2(n14730), .A(n10578), .ZN(n14759) );
  NOR2_X1 U13238 ( .A1(n14759), .A2(n14710), .ZN(n10586) );
  INV_X1 U13239 ( .A(n10580), .ZN(n10581) );
  AOI211_X1 U13240 ( .C1(n14757), .C2(n14726), .A(n14788), .B(n10581), .ZN(
        n14756) );
  AND2_X1 U13241 ( .A1(n10582), .A2(n13929), .ZN(n10583) );
  NAND2_X1 U13242 ( .A1(n13954), .A2(n10583), .ZN(n14696) );
  AOI22_X1 U13243 ( .A1(n14756), .A2(n14742), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n14737), .ZN(n10584) );
  OAI21_X1 U13244 ( .B1(n14691), .B2(n9809), .A(n10584), .ZN(n10585) );
  AOI211_X1 U13245 ( .C1(n14694), .C2(n14757), .A(n10586), .B(n10585), .ZN(
        n10587) );
  OAI21_X1 U13246 ( .B1(n10770), .B2(n14761), .A(n10587), .ZN(P1_U3291) );
  XNOR2_X1 U13247 ( .A(n13590), .B(n10588), .ZN(n13520) );
  XOR2_X1 U13248 ( .A(n13520), .B(n10589), .Z(n14777) );
  INV_X1 U13249 ( .A(n14777), .ZN(n10600) );
  AOI21_X1 U13250 ( .B1(n10590), .B2(n13590), .A(n14788), .ZN(n10591) );
  NAND2_X1 U13251 ( .A1(n10591), .A2(n14713), .ZN(n14772) );
  NAND2_X1 U13252 ( .A1(n14710), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10594) );
  OR2_X1 U13253 ( .A1(n14708), .A2(n10592), .ZN(n10593) );
  OAI211_X1 U13254 ( .C1(n14772), .C2(n14696), .A(n10594), .B(n10593), .ZN(
        n10598) );
  XNOR2_X1 U13255 ( .A(n10595), .B(n13520), .ZN(n10596) );
  NAND2_X1 U13256 ( .A1(n10596), .A2(n14730), .ZN(n14775) );
  AOI21_X1 U13257 ( .B1(n14775), .B2(n14774), .A(n14710), .ZN(n10597) );
  AOI211_X1 U13258 ( .C1(n14694), .C2(n13590), .A(n10598), .B(n10597), .ZN(
        n10599) );
  OAI21_X1 U13259 ( .B1(n10770), .B2(n10600), .A(n10599), .ZN(P1_U3288) );
  INV_X1 U13260 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10601) );
  AOI22_X1 U13261 ( .A1(n10602), .A2(n14742), .B1(n14737), .B2(n10601), .ZN(
        n10603) );
  OAI21_X1 U13262 ( .B1(n13578), .B2(n14739), .A(n10603), .ZN(n10606) );
  MUX2_X1 U13263 ( .A(n10604), .B(P1_REG2_REG_3__SCAN_IN), .S(n14746), .Z(
        n10605) );
  AOI211_X1 U13264 ( .C1(n14743), .C2(n10607), .A(n10606), .B(n10605), .ZN(
        n10608) );
  INV_X1 U13265 ( .A(n10608), .ZN(P1_U3290) );
  INV_X1 U13266 ( .A(n10609), .ZN(n10611) );
  MUX2_X1 U13267 ( .A(n10614), .B(n10613), .S(n6446), .Z(n10615) );
  NOR2_X1 U13268 ( .A1(n10615), .A2(n6641), .ZN(n10647) );
  INV_X1 U13269 ( .A(n10647), .ZN(n10616) );
  NAND2_X1 U13270 ( .A1(n10615), .A2(n6641), .ZN(n10646) );
  NAND2_X1 U13271 ( .A1(n10616), .A2(n10646), .ZN(n10617) );
  XNOR2_X1 U13272 ( .A(n10648), .B(n10617), .ZN(n10637) );
  NAND2_X1 U13273 ( .A1(n15084), .A2(n6641), .ZN(n10635) );
  NOR2_X1 U13274 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10618), .ZN(n11964) );
  AOI21_X1 U13275 ( .B1(n15087), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n11964), .ZN(
        n10634) );
  NAND2_X1 U13276 ( .A1(n10624), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n10619) );
  NAND2_X1 U13277 ( .A1(n10621), .A2(n10614), .ZN(n10622) );
  NAND2_X1 U13278 ( .A1(n10661), .A2(n10622), .ZN(n10623) );
  NAND2_X1 U13279 ( .A1(n15089), .A2(n10623), .ZN(n10633) );
  INV_X1 U13280 ( .A(n15097), .ZN(n10709) );
  NAND2_X1 U13281 ( .A1(n10624), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10625) );
  NAND2_X1 U13282 ( .A1(n10629), .A2(n10613), .ZN(n10630) );
  NAND2_X1 U13283 ( .A1(n10655), .A2(n10630), .ZN(n10631) );
  NAND2_X1 U13284 ( .A1(n10709), .A2(n10631), .ZN(n10632) );
  NAND4_X1 U13285 ( .A1(n10635), .A2(n10634), .A3(n10633), .A4(n10632), .ZN(
        n10636) );
  AOI21_X1 U13286 ( .B1(n10637), .B2(n15100), .A(n10636), .ZN(n10638) );
  INV_X1 U13287 ( .A(n10638), .ZN(P3_U3187) );
  INV_X1 U13288 ( .A(n14461), .ZN(n14578) );
  NOR2_X1 U13289 ( .A1(n14118), .A2(n14578), .ZN(n10645) );
  OAI22_X1 U13290 ( .A1(n14746), .A2(n10640), .B1(n10639), .B2(n14708), .ZN(
        n10643) );
  OR2_X1 U13291 ( .A1(n14746), .A2(n10641), .ZN(n14460) );
  AOI21_X1 U13292 ( .B1(n14739), .B2(n14460), .A(n14725), .ZN(n10642) );
  AOI211_X1 U13293 ( .C1(n14710), .C2(P1_REG2_REG_0__SCAN_IN), .A(n10643), .B(
        n10642), .ZN(n10644) );
  OAI21_X1 U13294 ( .B1(n13517), .B2(n10645), .A(n10644), .ZN(P1_U3293) );
  MUX2_X1 U13295 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n6446), .Z(n10946) );
  XNOR2_X1 U13296 ( .A(n10946), .B(n10657), .ZN(n10649) );
  NAND2_X1 U13297 ( .A1(n10649), .A2(n10650), .ZN(n10947) );
  OAI21_X1 U13298 ( .B1(n10650), .B2(n10649), .A(n10947), .ZN(n10651) );
  NAND2_X1 U13299 ( .A1(n10651), .A2(n15100), .ZN(n10669) );
  INV_X1 U13300 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15213) );
  MUX2_X1 U13301 ( .A(n15213), .B(P3_REG1_REG_6__SCAN_IN), .S(n10657), .Z(
        n10652) );
  INV_X1 U13302 ( .A(n10652), .ZN(n10654) );
  NAND3_X1 U13303 ( .A1(n10655), .A2(n10654), .A3(n10653), .ZN(n10656) );
  AND2_X1 U13304 ( .A1(n10937), .A2(n10656), .ZN(n10666) );
  MUX2_X1 U13305 ( .A(n8710), .B(P3_REG2_REG_6__SCAN_IN), .S(n10657), .Z(
        n10658) );
  INV_X1 U13306 ( .A(n10658), .ZN(n10660) );
  NAND3_X1 U13307 ( .A1(n10661), .A2(n10660), .A3(n10659), .ZN(n10662) );
  NAND2_X1 U13308 ( .A1(n15089), .A2(n10663), .ZN(n10665) );
  AND2_X1 U13309 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n10997) );
  AOI21_X1 U13310 ( .B1(n15087), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n10997), .ZN(
        n10664) );
  OAI211_X1 U13311 ( .C1(n10666), .C2(n15097), .A(n10665), .B(n10664), .ZN(
        n10667) );
  INV_X1 U13312 ( .A(n10667), .ZN(n10668) );
  OAI211_X1 U13313 ( .C1(n15068), .C2(n10956), .A(n10669), .B(n10668), .ZN(
        P3_U3188) );
  NAND2_X1 U13314 ( .A1(n10670), .A2(n10475), .ZN(n10671) );
  NAND2_X1 U13315 ( .A1(n10672), .A2(n10671), .ZN(n10673) );
  NAND2_X1 U13316 ( .A1(n15089), .A2(n10673), .ZN(n10681) );
  NAND2_X1 U13317 ( .A1(n10674), .A2(n10474), .ZN(n10675) );
  NAND2_X1 U13318 ( .A1(n10676), .A2(n10675), .ZN(n10677) );
  NAND2_X1 U13319 ( .A1(n10709), .A2(n10677), .ZN(n10680) );
  AOI21_X1 U13320 ( .B1(n15087), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10678), .ZN(
        n10679) );
  NAND3_X1 U13321 ( .A1(n10681), .A2(n10680), .A3(n10679), .ZN(n10682) );
  AOI21_X1 U13322 ( .B1(n10683), .B2(n15084), .A(n10682), .ZN(n10689) );
  AND3_X1 U13323 ( .A1(n10715), .A2(n10685), .A3(n10684), .ZN(n10686) );
  OAI21_X1 U13324 ( .B1(n10687), .B2(n10686), .A(n15100), .ZN(n10688) );
  NAND2_X1 U13325 ( .A1(n10689), .A2(n10688), .ZN(P3_U3185) );
  OR2_X1 U13326 ( .A1(n10690), .A2(n12141), .ZN(n10691) );
  NAND2_X1 U13327 ( .A1(n10692), .A2(n10691), .ZN(n15175) );
  INV_X1 U13328 ( .A(n15175), .ZN(n10701) );
  NAND2_X1 U13329 ( .A1(n12127), .A2(n15140), .ZN(n15133) );
  INV_X1 U13330 ( .A(n15133), .ZN(n15115) );
  NAND2_X1 U13331 ( .A1(n15159), .A2(n15115), .ZN(n15156) );
  INV_X1 U13332 ( .A(n15153), .ZN(n11117) );
  OAI22_X1 U13333 ( .A1(n10995), .A2(n12646), .B1(n10987), .B2(n12642), .ZN(
        n10697) );
  XNOR2_X1 U13334 ( .A(n10694), .B(n10693), .ZN(n10695) );
  INV_X1 U13335 ( .A(n15149), .ZN(n12582) );
  NOR2_X1 U13336 ( .A1(n10695), .A2(n12582), .ZN(n10696) );
  AOI211_X1 U13337 ( .C1(n11117), .C2(n15175), .A(n10697), .B(n10696), .ZN(
        n15177) );
  MUX2_X1 U13338 ( .A(n10455), .B(n15177), .S(n15159), .Z(n10700) );
  INV_X1 U13339 ( .A(n10698), .ZN(n11994) );
  AOI22_X1 U13340 ( .A1(n14499), .A2(n15174), .B1(n15136), .B2(n11994), .ZN(
        n10699) );
  OAI211_X1 U13341 ( .C1(n10701), .C2(n15156), .A(n10700), .B(n10699), .ZN(
        P3_U3229) );
  OAI21_X1 U13342 ( .B1(n10704), .B2(n10703), .A(n10702), .ZN(n10714) );
  OAI21_X1 U13343 ( .B1(n10707), .B2(n10706), .A(n10705), .ZN(n10708) );
  AND2_X1 U13344 ( .A1(n10709), .A2(n10708), .ZN(n10713) );
  INV_X1 U13345 ( .A(n15087), .ZN(n15065) );
  INV_X1 U13346 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10711) );
  OAI22_X1 U13347 ( .A1(n15065), .A2(n10711), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10710), .ZN(n10712) );
  AOI211_X1 U13348 ( .C1(n15089), .C2(n10714), .A(n10713), .B(n10712), .ZN(
        n10721) );
  INV_X1 U13349 ( .A(n10715), .ZN(n10719) );
  NOR3_X1 U13350 ( .A1(n10717), .A2(n10716), .A3(n7640), .ZN(n10718) );
  OAI21_X1 U13351 ( .B1(n10719), .B2(n10718), .A(n15100), .ZN(n10720) );
  OAI211_X1 U13352 ( .C1(n15068), .C2(n10722), .A(n10721), .B(n10720), .ZN(
        P3_U3184) );
  MUX2_X1 U13353 ( .A(n9317), .B(P1_REG2_REG_13__SCAN_IN), .S(n11266), .Z(
        n11267) );
  AOI21_X1 U13354 ( .B1(n10728), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10723), 
        .ZN(n14646) );
  MUX2_X1 U13355 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n11326), .S(n14655), .Z(
        n14647) );
  NAND2_X1 U13356 ( .A1(n14646), .A2(n14647), .ZN(n14645) );
  OAI21_X1 U13357 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n14655), .A(n14645), 
        .ZN(n11268) );
  XOR2_X1 U13358 ( .A(n11267), .B(n11268), .Z(n10735) );
  INV_X1 U13359 ( .A(n11266), .ZN(n10726) );
  NAND2_X1 U13360 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n11489)
         );
  INV_X1 U13361 ( .A(n11489), .ZN(n10724) );
  AOI21_X1 U13362 ( .B1(n14624), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10724), 
        .ZN(n10725) );
  OAI21_X1 U13363 ( .B1(n13924), .B2(n10726), .A(n10725), .ZN(n10734) );
  INV_X1 U13364 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10727) );
  MUX2_X1 U13365 ( .A(n10727), .B(P1_REG1_REG_13__SCAN_IN), .S(n11266), .Z(
        n10732) );
  NOR2_X1 U13366 ( .A1(n10728), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n14648) );
  INV_X1 U13367 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10729) );
  MUX2_X1 U13368 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10729), .S(n14655), .Z(
        n10730) );
  OAI21_X1 U13369 ( .B1(n14653), .B2(n14648), .A(n10730), .ZN(n14651) );
  OAI21_X1 U13370 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n14655), .A(n14651), 
        .ZN(n10731) );
  NOR2_X1 U13371 ( .A1(n10731), .A2(n10732), .ZN(n11258) );
  AOI211_X1 U13372 ( .C1(n10732), .C2(n10731), .A(n13799), .B(n11258), .ZN(
        n10733) );
  AOI211_X1 U13373 ( .C1(n14656), .C2(n10735), .A(n10734), .B(n10733), .ZN(
        n10736) );
  INV_X1 U13374 ( .A(n10736), .ZN(P1_U3256) );
  INV_X1 U13375 ( .A(n10737), .ZN(n11018) );
  NAND2_X1 U13376 ( .A1(n13603), .A2(n14758), .ZN(n14785) );
  INV_X1 U13377 ( .A(n10738), .ZN(n10742) );
  INV_X1 U13378 ( .A(n10739), .ZN(n10741) );
  OAI22_X1 U13379 ( .A1(n10765), .A2(n11835), .B1(n10791), .B2(n11837), .ZN(
        n10743) );
  NOR2_X1 U13380 ( .A1(n11836), .A2(n10791), .ZN(n10744) );
  AOI21_X1 U13381 ( .B1(n13603), .B2(n11827), .A(n10744), .ZN(n10846) );
  XNOR2_X1 U13382 ( .A(n10845), .B(n10846), .ZN(n10745) );
  OAI211_X1 U13383 ( .C1(n10746), .C2(n10745), .A(n10847), .B(n14564), .ZN(
        n10752) );
  OR2_X1 U13384 ( .A1(n13593), .A2(n14734), .ZN(n10748) );
  NAND2_X1 U13385 ( .A1(n13792), .A2(n13479), .ZN(n10747) );
  NAND2_X1 U13386 ( .A1(n10748), .A2(n10747), .ZN(n10760) );
  NOR2_X1 U13387 ( .A1(n10749), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13858) );
  NOR2_X1 U13388 ( .A1(n15385), .A2(n10764), .ZN(n10750) );
  AOI211_X1 U13389 ( .C1(n14566), .C2(n10760), .A(n13858), .B(n10750), .ZN(
        n10751) );
  OAI211_X1 U13390 ( .C1(n11018), .C2(n14785), .A(n10752), .B(n10751), .ZN(
        P1_U3213) );
  INV_X1 U13391 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10754) );
  INV_X1 U13392 ( .A(n10753), .ZN(n10755) );
  OAI222_X1 U13393 ( .A1(n13372), .A2(n10754), .B1(n13367), .B2(n10755), .C1(
        P2_U3088), .C2(n11306), .ZN(P2_U3312) );
  INV_X1 U13394 ( .A(n14668), .ZN(n11273) );
  OAI222_X1 U13395 ( .A1(n14318), .A2(n10756), .B1(n14312), .B2(n10755), .C1(
        P1_U3086), .C2(n11273), .ZN(P1_U3340) );
  XNOR2_X1 U13396 ( .A(n10757), .B(n13523), .ZN(n14790) );
  OAI211_X1 U13397 ( .C1(n10759), .C2(n13523), .A(n10758), .B(n14730), .ZN(
        n10762) );
  INV_X1 U13398 ( .A(n10760), .ZN(n10761) );
  AND2_X1 U13399 ( .A1(n10762), .A2(n10761), .ZN(n14786) );
  MUX2_X1 U13400 ( .A(n9839), .B(n14786), .S(n14691), .Z(n10769) );
  INV_X1 U13401 ( .A(n10795), .ZN(n10763) );
  OAI21_X1 U13402 ( .B1(n10765), .B2(n14714), .A(n10763), .ZN(n14787) );
  INV_X1 U13403 ( .A(n14787), .ZN(n10767) );
  INV_X1 U13404 ( .A(n14460), .ZN(n13986) );
  OAI22_X1 U13405 ( .A1(n14739), .A2(n10765), .B1(n14708), .B2(n10764), .ZN(
        n10766) );
  AOI21_X1 U13406 ( .B1(n10767), .B2(n13986), .A(n10766), .ZN(n10768) );
  OAI211_X1 U13407 ( .C1(n10770), .C2(n14790), .A(n10769), .B(n10768), .ZN(
        P1_U3286) );
  NAND2_X1 U13408 ( .A1(n10771), .A2(n11855), .ZN(n10772) );
  OAI211_X1 U13409 ( .C1(n10773), .C2(n11873), .A(n10772), .B(n12273), .ZN(
        P3_U3272) );
  NAND2_X1 U13410 ( .A1(n10777), .A2(n10776), .ZN(n10778) );
  XNOR2_X1 U13411 ( .A(n11089), .B(n11592), .ZN(n10823) );
  NAND2_X1 U13412 ( .A1(n12909), .A2(n13194), .ZN(n10824) );
  XNOR2_X1 U13413 ( .A(n10823), .B(n10824), .ZN(n10781) );
  AOI22_X1 U13414 ( .A1(n12847), .A2(n12910), .B1(n12848), .B2(n12908), .ZN(
        n10779) );
  NAND2_X1 U13415 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n14891) );
  OAI211_X1 U13416 ( .C1(n10886), .C2(n12877), .A(n10779), .B(n14891), .ZN(
        n10785) );
  OR2_X1 U13417 ( .A1(n10780), .A2(n12902), .ZN(n10783) );
  NAND3_X1 U13418 ( .A1(n10777), .A2(n12893), .A3(n12910), .ZN(n10782) );
  AOI21_X1 U13419 ( .B1(n10783), .B2(n10782), .A(n10781), .ZN(n10784) );
  AOI211_X1 U13420 ( .C1(n11089), .C2(n12900), .A(n10785), .B(n10784), .ZN(
        n10786) );
  OAI21_X1 U13421 ( .B1(n10827), .B2(n12902), .A(n10786), .ZN(P2_U3203) );
  NAND2_X1 U13422 ( .A1(n12275), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n10787) );
  OAI21_X1 U13423 ( .B1(n12472), .B2(n12275), .A(n10787), .ZN(P3_U3519) );
  XOR2_X1 U13424 ( .A(n10788), .B(n13525), .Z(n14800) );
  INV_X1 U13425 ( .A(n14800), .ZN(n10801) );
  OAI211_X1 U13426 ( .C1(n10790), .C2(n13525), .A(n10789), .B(n14730), .ZN(
        n10794) );
  OR2_X1 U13427 ( .A1(n10791), .A2(n14734), .ZN(n10793) );
  NAND2_X1 U13428 ( .A1(n13791), .A2(n13479), .ZN(n10792) );
  AND2_X1 U13429 ( .A1(n10793), .A2(n10792), .ZN(n10851) );
  NAND2_X1 U13430 ( .A1(n10794), .A2(n10851), .ZN(n14798) );
  OAI211_X1 U13431 ( .C1(n10795), .C2(n14797), .A(n14715), .B(n14686), .ZN(
        n14795) );
  INV_X1 U13432 ( .A(n10796), .ZN(n10853) );
  AOI22_X1 U13433 ( .A1(n14710), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n10853), 
        .B2(n14737), .ZN(n10798) );
  NAND2_X1 U13434 ( .A1(n14694), .A2(n13607), .ZN(n10797) );
  OAI211_X1 U13435 ( .C1(n14795), .C2(n14696), .A(n10798), .B(n10797), .ZN(
        n10799) );
  AOI21_X1 U13436 ( .B1(n14798), .B2(n14691), .A(n10799), .ZN(n10800) );
  OAI21_X1 U13437 ( .B1(n10801), .B2(n14461), .A(n10800), .ZN(P1_U3285) );
  INV_X1 U13438 ( .A(n10802), .ZN(n10805) );
  INV_X1 U13439 ( .A(n11456), .ZN(n11276) );
  OAI222_X1 U13440 ( .A1(n14318), .A2(n10803), .B1(n14312), .B2(n10805), .C1(
        n11276), .C2(P1_U3086), .ZN(P1_U3339) );
  OAI222_X1 U13441 ( .A1(P2_U3088), .A2(n11309), .B1(n13367), .B2(n10805), 
        .C1(n10804), .C2(n13372), .ZN(P2_U3311) );
  NAND2_X1 U13442 ( .A1(n12275), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10806) );
  OAI21_X1 U13443 ( .B1(n12086), .B2(n12275), .A(n10806), .ZN(P3_U3521) );
  NAND2_X1 U13444 ( .A1(n12275), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n10807) );
  OAI21_X1 U13445 ( .B1(n12458), .B2(n12275), .A(n10807), .ZN(P3_U3520) );
  XNOR2_X1 U13446 ( .A(n10808), .B(n12146), .ZN(n15178) );
  OAI21_X1 U13447 ( .B1(n10810), .B2(n12146), .A(n10809), .ZN(n10811) );
  NAND2_X1 U13448 ( .A1(n10811), .A2(n15149), .ZN(n10813) );
  AOI22_X1 U13449 ( .A1(n15145), .A2(n12284), .B1(n15108), .B2(n15142), .ZN(
        n10812) );
  OAI211_X1 U13450 ( .C1(n15178), .C2(n15153), .A(n10813), .B(n10812), .ZN(
        n15179) );
  MUX2_X1 U13451 ( .A(P3_REG2_REG_5__SCAN_IN), .B(n15179), .S(n15159), .Z(
        n10814) );
  INV_X1 U13452 ( .A(n10814), .ZN(n10817) );
  INV_X1 U13453 ( .A(n11237), .ZN(n15118) );
  NOR2_X1 U13454 ( .A1(n11963), .A2(n15138), .ZN(n15180) );
  INV_X1 U13455 ( .A(n10815), .ZN(n11966) );
  AOI22_X1 U13456 ( .A1(n15118), .A2(n15180), .B1(n15136), .B2(n11966), .ZN(
        n10816) );
  OAI211_X1 U13457 ( .C1(n15178), .C2(n15156), .A(n10817), .B(n10816), .ZN(
        P3_U3228) );
  INV_X1 U13458 ( .A(n10818), .ZN(n10821) );
  INV_X1 U13459 ( .A(n13906), .ZN(n13903) );
  OAI222_X1 U13460 ( .A1(n14318), .A2(n10819), .B1(n14312), .B2(n10821), .C1(
        n13903), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U13461 ( .A(n12974), .ZN(n10822) );
  OAI222_X1 U13462 ( .A1(P2_U3088), .A2(n10822), .B1(n13367), .B2(n10821), 
        .C1(n10820), .C2(n13372), .ZN(P2_U3310) );
  INV_X1 U13463 ( .A(n10823), .ZN(n10825) );
  NAND2_X1 U13464 ( .A1(n10825), .A2(n10824), .ZN(n10826) );
  AND2_X1 U13465 ( .A1(n12908), .A2(n13194), .ZN(n10828) );
  NAND2_X1 U13466 ( .A1(n10829), .A2(n10828), .ZN(n10831) );
  OAI21_X1 U13467 ( .B1(n10829), .B2(n10828), .A(n10831), .ZN(n10933) );
  INV_X1 U13468 ( .A(n12908), .ZN(n11193) );
  NOR2_X1 U13469 ( .A1(n12860), .A2(n11193), .ZN(n10830) );
  AOI22_X1 U13470 ( .A1(n10931), .A2(n12871), .B1(n10830), .B2(n10829), .ZN(
        n10839) );
  XNOR2_X1 U13471 ( .A(n11376), .B(n6911), .ZN(n11039) );
  NAND2_X1 U13472 ( .A1(n12907), .A2(n13194), .ZN(n11040) );
  XNOR2_X1 U13473 ( .A(n11039), .B(n11040), .ZN(n10833) );
  INV_X1 U13474 ( .A(n10833), .ZN(n10838) );
  INV_X1 U13475 ( .A(n10831), .ZN(n10832) );
  NAND2_X1 U13476 ( .A1(n11049), .A2(n12871), .ZN(n10837) );
  AOI22_X1 U13477 ( .A1(n12847), .A2(n12908), .B1(n12848), .B2(n12906), .ZN(
        n10834) );
  NAND2_X1 U13478 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n14905)
         );
  OAI211_X1 U13479 ( .C1(n11203), .C2(n12877), .A(n10834), .B(n14905), .ZN(
        n10835) );
  AOI21_X1 U13480 ( .B1(n11376), .B2(n12900), .A(n10835), .ZN(n10836) );
  OAI211_X1 U13481 ( .C1(n10839), .C2(n10838), .A(n10837), .B(n10836), .ZN(
        P2_U3208) );
  INV_X1 U13482 ( .A(n13792), .ZN(n10840) );
  NOR2_X1 U13483 ( .A1(n11836), .A2(n10840), .ZN(n10841) );
  AOI21_X1 U13484 ( .B1(n13607), .B2(n11827), .A(n10841), .ZN(n10971) );
  NAND2_X1 U13485 ( .A1(n13607), .A2(n11826), .ZN(n10843) );
  NAND2_X1 U13486 ( .A1(n11827), .A2(n13792), .ZN(n10842) );
  NAND2_X1 U13487 ( .A1(n10843), .A2(n10842), .ZN(n10844) );
  XNOR2_X1 U13488 ( .A(n10844), .B(n11838), .ZN(n10970) );
  XOR2_X1 U13489 ( .A(n10971), .B(n10970), .Z(n10849) );
  AOI21_X1 U13490 ( .B1(n10849), .B2(n10848), .A(n11005), .ZN(n10856) );
  INV_X1 U13491 ( .A(n15385), .ZN(n13481) );
  OAI22_X1 U13492 ( .A1(n15388), .A2(n10851), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10850), .ZN(n10852) );
  AOI21_X1 U13493 ( .B1(n13481), .B2(n10853), .A(n10852), .ZN(n10855) );
  NAND2_X1 U13494 ( .A1(n14562), .A2(n13607), .ZN(n10854) );
  OAI211_X1 U13495 ( .C1(n10856), .C2(n15379), .A(n10855), .B(n10854), .ZN(
        P1_U3221) );
  INV_X1 U13496 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n10866) );
  INV_X1 U13497 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12454) );
  NAND2_X1 U13498 ( .A1(n8638), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n10859) );
  INV_X1 U13499 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n10857) );
  OR2_X1 U13500 ( .A1(n8639), .A2(n10857), .ZN(n10858) );
  OAI211_X1 U13501 ( .C1(n12454), .C2(n10860), .A(n10859), .B(n10858), .ZN(
        n10861) );
  INV_X1 U13502 ( .A(n10861), .ZN(n10862) );
  INV_X1 U13503 ( .A(n12450), .ZN(n10864) );
  NAND2_X1 U13504 ( .A1(n10864), .A2(n12285), .ZN(n10865) );
  OAI21_X1 U13505 ( .B1(n12285), .B2(n10866), .A(n10865), .ZN(P3_U3522) );
  NAND2_X1 U13506 ( .A1(n10872), .A2(n12911), .ZN(n10867) );
  INV_X1 U13507 ( .A(n10877), .ZN(n10879) );
  OR2_X1 U13508 ( .A1(n10870), .A2(n10879), .ZN(n10871) );
  AND2_X1 U13509 ( .A1(n10872), .A2(n10917), .ZN(n10873) );
  NAND2_X1 U13510 ( .A1(n15010), .A2(n12911), .ZN(n10875) );
  NAND2_X1 U13511 ( .A1(n10876), .A2(n10869), .ZN(n10915) );
  INV_X1 U13512 ( .A(n12910), .ZN(n10881) );
  NAND2_X1 U13513 ( .A1(n15018), .A2(n10881), .ZN(n10878) );
  NAND3_X1 U13514 ( .A1(n10915), .A2(n10879), .A3(n10878), .ZN(n10880) );
  AOI21_X1 U13515 ( .B1(n10897), .B2(n10880), .A(n13137), .ZN(n10883) );
  OAI22_X1 U13516 ( .A1(n10881), .A2(n13139), .B1(n11193), .B2(n13141), .ZN(
        n10882) );
  AOI211_X1 U13517 ( .C1(n11088), .C2(n11212), .A(n10883), .B(n10882), .ZN(
        n11092) );
  INV_X1 U13518 ( .A(n11089), .ZN(n10884) );
  NOR2_X1 U13519 ( .A1(n10922), .A2(n15018), .ZN(n10921) );
  NAND2_X1 U13520 ( .A1(n10884), .A2(n10921), .ZN(n10903) );
  OR2_X1 U13521 ( .A1(n10884), .A2(n10921), .ZN(n10885) );
  AND2_X1 U13522 ( .A1(n10903), .A2(n10885), .ZN(n11090) );
  NAND2_X1 U13523 ( .A1(n11090), .A2(n13131), .ZN(n10890) );
  OAI22_X1 U13524 ( .A1(n13219), .A2(n10887), .B1(n10886), .B2(n13217), .ZN(
        n10888) );
  AOI21_X1 U13525 ( .B1(n11089), .B2(n13234), .A(n10888), .ZN(n10889) );
  NAND2_X1 U13526 ( .A1(n10890), .A2(n10889), .ZN(n10891) );
  AOI21_X1 U13527 ( .B1(n11088), .B2(n10908), .A(n10891), .ZN(n10892) );
  OAI21_X1 U13528 ( .B1(n11092), .B2(n13212), .A(n10892), .ZN(P2_U3256) );
  XNOR2_X1 U13529 ( .A(n11195), .B(n10895), .ZN(n15034) );
  INV_X1 U13530 ( .A(n12909), .ZN(n10916) );
  NAND2_X1 U13531 ( .A1(n11089), .A2(n10916), .ZN(n10896) );
  INV_X1 U13532 ( .A(n10895), .ZN(n11194) );
  NAND3_X1 U13533 ( .A1(n10897), .A2(n11194), .A3(n10896), .ZN(n10898) );
  NAND2_X1 U13534 ( .A1(n11190), .A2(n10898), .ZN(n10899) );
  NAND2_X1 U13535 ( .A1(n10899), .A2(n13228), .ZN(n10901) );
  AOI22_X1 U13536 ( .A1(n13225), .A2(n12909), .B1(n12907), .B2(n13223), .ZN(
        n10900) );
  NAND2_X1 U13537 ( .A1(n10901), .A2(n10900), .ZN(n10902) );
  AOI21_X1 U13538 ( .B1(n15034), .B2(n11212), .A(n10902), .ZN(n15036) );
  NAND2_X1 U13539 ( .A1(n15027), .A2(n10903), .ZN(n10904) );
  NAND2_X1 U13540 ( .A1(n11202), .A2(n10904), .ZN(n15031) );
  OAI22_X1 U13541 ( .A1(n13219), .A2(n9866), .B1(n10930), .B2(n13217), .ZN(
        n10905) );
  AOI21_X1 U13542 ( .B1(n15027), .B2(n13234), .A(n10905), .ZN(n10906) );
  OAI21_X1 U13543 ( .B1(n15031), .B2(n12989), .A(n10906), .ZN(n10907) );
  AOI21_X1 U13544 ( .B1(n15034), .B2(n10908), .A(n10907), .ZN(n10909) );
  OAI21_X1 U13545 ( .B1(n15036), .B2(n13212), .A(n10909), .ZN(P2_U3255) );
  OAI21_X1 U13546 ( .B1(n10911), .B2(n10912), .A(n10910), .ZN(n15022) );
  INV_X1 U13547 ( .A(n15022), .ZN(n10920) );
  NAND2_X1 U13548 ( .A1(n10913), .A2(n10912), .ZN(n10914) );
  AOI21_X1 U13549 ( .B1(n10915), .B2(n10914), .A(n13137), .ZN(n10919) );
  OAI22_X1 U13550 ( .A1(n10917), .A2(n13139), .B1(n10916), .B2(n13141), .ZN(
        n10918) );
  AOI211_X1 U13551 ( .C1(n10920), .C2(n11212), .A(n10919), .B(n10918), .ZN(
        n15021) );
  MUX2_X1 U13552 ( .A(n9878), .B(n15021), .S(n13219), .Z(n10927) );
  AOI211_X1 U13553 ( .C1(n15018), .C2(n10922), .A(n15030), .B(n10921), .ZN(
        n15017) );
  INV_X1 U13554 ( .A(n15018), .ZN(n10924) );
  OAI22_X1 U13555 ( .A1(n10924), .A2(n13147), .B1(n10923), .B2(n13217), .ZN(
        n10925) );
  AOI21_X1 U13556 ( .B1(n15017), .B2(n13175), .A(n10925), .ZN(n10926) );
  OAI211_X1 U13557 ( .C1(n15022), .C2(n13072), .A(n10927), .B(n10926), .ZN(
        P2_U3257) );
  AOI22_X1 U13558 ( .A1(n12847), .A2(n12909), .B1(n12848), .B2(n12907), .ZN(
        n10929) );
  OAI211_X1 U13559 ( .C1(n10930), .C2(n12877), .A(n10929), .B(n10928), .ZN(
        n10935) );
  AOI211_X1 U13560 ( .C1(n10933), .C2(n10932), .A(n12902), .B(n10931), .ZN(
        n10934) );
  AOI211_X1 U13561 ( .C1(n15027), .C2(n12900), .A(n10935), .B(n10934), .ZN(
        n10936) );
  INV_X1 U13562 ( .A(n10936), .ZN(P2_U3189) );
  NOR2_X1 U13563 ( .A1(n15053), .A2(n10938), .ZN(n10939) );
  AOI22_X1 U13564 ( .A1(n11072), .A2(P3_REG1_REG_8__SCAN_IN), .B1(n10942), 
        .B2(n11081), .ZN(n10940) );
  AOI21_X1 U13565 ( .B1(n10941), .B2(n10940), .A(n11067), .ZN(n10964) );
  INV_X1 U13566 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n10955) );
  MUX2_X1 U13567 ( .A(n10943), .B(n10942), .S(n6446), .Z(n11073) );
  XNOR2_X1 U13568 ( .A(n11073), .B(n11081), .ZN(n10951) );
  MUX2_X1 U13569 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n6446), .Z(n10945) );
  OR2_X1 U13570 ( .A1(n10945), .A2(n10944), .ZN(n10949) );
  XNOR2_X1 U13571 ( .A(n10945), .B(n15053), .ZN(n15051) );
  OR2_X1 U13572 ( .A1(n10946), .A2(n10956), .ZN(n10948) );
  NAND2_X1 U13573 ( .A1(n10948), .A2(n10947), .ZN(n15050) );
  NAND2_X1 U13574 ( .A1(n10949), .A2(n15049), .ZN(n10950) );
  NAND2_X1 U13575 ( .A1(n10951), .A2(n10950), .ZN(n11074) );
  OAI21_X1 U13576 ( .B1(n10951), .B2(n10950), .A(n11074), .ZN(n10952) );
  NAND2_X1 U13577 ( .A1(n15100), .A2(n10952), .ZN(n10954) );
  AND2_X1 U13578 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n11915) );
  INV_X1 U13579 ( .A(n11915), .ZN(n10953) );
  OAI211_X1 U13580 ( .C1(n15065), .C2(n10955), .A(n10954), .B(n10953), .ZN(
        n10962) );
  XNOR2_X1 U13581 ( .A(n15053), .B(n10957), .ZN(n15054) );
  AOI22_X1 U13582 ( .A1(n11072), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n10943), 
        .B2(n11081), .ZN(n10958) );
  AOI21_X1 U13583 ( .B1(n10959), .B2(n10958), .A(n11080), .ZN(n10960) );
  NOR2_X1 U13584 ( .A1(n10960), .A2(n15081), .ZN(n10961) );
  AOI211_X1 U13585 ( .C1(n15084), .C2(n11072), .A(n10962), .B(n10961), .ZN(
        n10963) );
  OAI21_X1 U13586 ( .B1(n10964), .B2(n15097), .A(n10963), .ZN(P3_U3190) );
  NAND2_X1 U13587 ( .A1(n14693), .A2(n11826), .ZN(n10966) );
  NAND2_X1 U13588 ( .A1(n11827), .A2(n13791), .ZN(n10965) );
  NAND2_X1 U13589 ( .A1(n10966), .A2(n10965), .ZN(n10967) );
  XNOR2_X1 U13590 ( .A(n10967), .B(n11838), .ZN(n11008) );
  NAND2_X1 U13591 ( .A1(n14693), .A2(n11827), .ZN(n10969) );
  NAND2_X1 U13592 ( .A1(n11831), .A2(n13791), .ZN(n10968) );
  NAND2_X1 U13593 ( .A1(n10969), .A2(n10968), .ZN(n10973) );
  INV_X1 U13594 ( .A(n10970), .ZN(n10972) );
  NAND2_X1 U13595 ( .A1(n10972), .A2(n10971), .ZN(n11006) );
  OAI21_X1 U13596 ( .B1(n11008), .B2(n10973), .A(n11006), .ZN(n10974) );
  INV_X1 U13597 ( .A(n10973), .ZN(n11007) );
  NAND2_X1 U13598 ( .A1(n13618), .A2(n11826), .ZN(n10976) );
  OR2_X1 U13599 ( .A1(n11344), .A2(n11837), .ZN(n10975) );
  NAND2_X1 U13600 ( .A1(n10976), .A2(n10975), .ZN(n10977) );
  XNOR2_X1 U13601 ( .A(n10977), .B(n11838), .ZN(n11465) );
  NAND2_X1 U13602 ( .A1(n13618), .A2(n11827), .ZN(n10979) );
  NAND2_X1 U13603 ( .A1(n13790), .A2(n11831), .ZN(n10978) );
  NAND2_X1 U13604 ( .A1(n10979), .A2(n10978), .ZN(n11464) );
  INV_X1 U13605 ( .A(n11464), .ZN(n11466) );
  XNOR2_X1 U13606 ( .A(n11465), .B(n11466), .ZN(n10980) );
  XNOR2_X1 U13607 ( .A(n11463), .B(n10980), .ZN(n10984) );
  OR2_X1 U13608 ( .A1(n11471), .A2(n13487), .ZN(n11055) );
  NAND2_X1 U13609 ( .A1(n13791), .A2(n13478), .ZN(n11057) );
  AND2_X1 U13610 ( .A1(n11055), .A2(n11057), .ZN(n11101) );
  NAND2_X1 U13611 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n13874)
         );
  OAI21_X1 U13612 ( .B1(n15388), .B2(n11101), .A(n13874), .ZN(n10982) );
  NOR2_X1 U13613 ( .A1(n15385), .A2(n11056), .ZN(n10981) );
  AOI211_X1 U13614 ( .C1(n13618), .C2(n14562), .A(n10982), .B(n10981), .ZN(
        n10983) );
  OAI21_X1 U13615 ( .B1(n10984), .B2(n15379), .A(n10983), .ZN(P1_U3217) );
  NAND2_X1 U13616 ( .A1(n10989), .A2(n10988), .ZN(n10990) );
  INV_X1 U13617 ( .A(n10990), .ZN(n10991) );
  XNOR2_X1 U13618 ( .A(n10992), .B(n11993), .ZN(n11960) );
  NOR2_X1 U13619 ( .A1(n11959), .A2(n11128), .ZN(n10994) );
  XNOR2_X1 U13620 ( .A(n11622), .B(n10998), .ZN(n11132) );
  XNOR2_X1 U13621 ( .A(n11132), .B(n12284), .ZN(n10993) );
  NAND2_X1 U13622 ( .A1(n10994), .A2(n10993), .ZN(n11875) );
  OAI211_X1 U13623 ( .C1(n10994), .C2(n10993), .A(n11875), .B(n12041), .ZN(
        n11000) );
  INV_X1 U13624 ( .A(n12283), .ZN(n11134) );
  OAI22_X1 U13625 ( .A1(n12052), .A2(n10995), .B1(n11134), .B2(n12065), .ZN(
        n10996) );
  AOI211_X1 U13626 ( .C1(n12036), .C2(n10998), .A(n10997), .B(n10996), .ZN(
        n10999) );
  OAI211_X1 U13627 ( .C1(n11113), .C2(n12028), .A(n11000), .B(n10999), .ZN(
        P3_U3179) );
  INV_X1 U13628 ( .A(n11001), .ZN(n11004) );
  OAI222_X1 U13629 ( .A1(n14434), .A2(n11004), .B1(n11873), .B2(n11003), .C1(
        P3_U3151), .C2(n11002), .ZN(P3_U3270) );
  NAND2_X1 U13630 ( .A1(n14693), .A2(n14758), .ZN(n14801) );
  NAND2_X1 U13631 ( .A1(n7495), .A2(n11006), .ZN(n11010) );
  XNOR2_X1 U13632 ( .A(n11008), .B(n11007), .ZN(n11009) );
  XNOR2_X1 U13633 ( .A(n11010), .B(n11009), .ZN(n11011) );
  NAND2_X1 U13634 ( .A1(n11011), .A2(n14564), .ZN(n11017) );
  INV_X1 U13635 ( .A(n14689), .ZN(n11015) );
  OR2_X1 U13636 ( .A1(n11344), .A2(n13487), .ZN(n11013) );
  NAND2_X1 U13637 ( .A1(n13792), .A2(n13478), .ZN(n11012) );
  AND2_X1 U13638 ( .A1(n11013), .A2(n11012), .ZN(n14802) );
  OAI22_X1 U13639 ( .A1(n15388), .A2(n14802), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15259), .ZN(n11014) );
  AOI21_X1 U13640 ( .B1(n13481), .B2(n11015), .A(n11014), .ZN(n11016) );
  OAI211_X1 U13641 ( .C1(n11018), .C2(n14801), .A(n11017), .B(n11016), .ZN(
        P1_U3231) );
  XNOR2_X1 U13642 ( .A(n11019), .B(n11021), .ZN(n11026) );
  OR2_X1 U13643 ( .A1(n11020), .A2(n12162), .ZN(n11155) );
  OAI21_X1 U13644 ( .B1(n11022), .B2(n11021), .A(n11155), .ZN(n11023) );
  NAND2_X1 U13645 ( .A1(n11023), .A2(n15149), .ZN(n11025) );
  AOI22_X1 U13646 ( .A1(n15142), .A2(n12283), .B1(n12281), .B2(n15145), .ZN(
        n11024) );
  OAI211_X1 U13647 ( .C1(n15153), .C2(n11026), .A(n11025), .B(n11024), .ZN(
        n15192) );
  INV_X1 U13648 ( .A(n15192), .ZN(n11032) );
  INV_X1 U13649 ( .A(n11026), .ZN(n15194) );
  INV_X1 U13650 ( .A(n15156), .ZN(n11175) );
  NOR2_X1 U13651 ( .A1(n11027), .A2(n15138), .ZN(n15193) );
  INV_X1 U13652 ( .A(n11028), .ZN(n11917) );
  AOI22_X1 U13653 ( .A1(n15118), .A2(n15193), .B1(n15136), .B2(n11917), .ZN(
        n11029) );
  OAI21_X1 U13654 ( .B1(n10943), .B2(n15159), .A(n11029), .ZN(n11030) );
  AOI21_X1 U13655 ( .B1(n15194), .B2(n11175), .A(n11030), .ZN(n11031) );
  OAI21_X1 U13656 ( .B1(n11032), .B2(n14498), .A(n11031), .ZN(P3_U3225) );
  INV_X1 U13657 ( .A(n11033), .ZN(n11035) );
  OAI222_X1 U13658 ( .A1(n14318), .A2(n11034), .B1(n14312), .B2(n11035), .C1(
        P1_U3086), .C2(n13914), .ZN(P1_U3337) );
  INV_X1 U13659 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n15269) );
  INV_X1 U13660 ( .A(n12969), .ZN(n14980) );
  OAI222_X1 U13661 ( .A1(n13372), .A2(n15269), .B1(n13367), .B2(n11035), .C1(
        P2_U3088), .C2(n14980), .ZN(P2_U3309) );
  INV_X1 U13662 ( .A(n11036), .ZN(n11038) );
  INV_X1 U13663 ( .A(SI_24_), .ZN(n11037) );
  OAI222_X1 U13664 ( .A1(P3_U3151), .A2(n9084), .B1(n14434), .B2(n11038), .C1(
        n11037), .C2(n11873), .ZN(P3_U3271) );
  INV_X1 U13665 ( .A(n11039), .ZN(n11046) );
  INV_X1 U13666 ( .A(n11040), .ZN(n11041) );
  NOR2_X1 U13667 ( .A1(n11046), .A2(n11041), .ZN(n11042) );
  XNOR2_X1 U13668 ( .A(n11361), .B(n11592), .ZN(n11180) );
  NAND2_X1 U13669 ( .A1(n12906), .A2(n13194), .ZN(n11178) );
  XNOR2_X1 U13670 ( .A(n11180), .B(n11178), .ZN(n11047) );
  NAND2_X1 U13671 ( .A1(n13226), .A2(n13223), .ZN(n11044) );
  NAND2_X1 U13672 ( .A1(n12907), .A2(n13225), .ZN(n11043) );
  NAND2_X1 U13673 ( .A1(n11044), .A2(n11043), .ZN(n11217) );
  AOI22_X1 U13674 ( .A1(n12880), .A2(n11217), .B1(P2_REG3_REG_12__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11045) );
  OAI21_X1 U13675 ( .B1(n11224), .B2(n12877), .A(n11045), .ZN(n11051) );
  AOI22_X1 U13676 ( .A1(n11046), .A2(n12871), .B1(n12893), .B2(n12907), .ZN(
        n11048) );
  NOR3_X1 U13677 ( .A1(n11049), .A2(n11048), .A3(n11047), .ZN(n11050) );
  AOI211_X1 U13678 ( .C1(n11361), .C2(n12900), .A(n11051), .B(n11050), .ZN(
        n11052) );
  OAI21_X1 U13679 ( .B1(n11179), .B2(n12902), .A(n11052), .ZN(P2_U3196) );
  OAI21_X1 U13680 ( .B1(n11054), .B2(n13529), .A(n11053), .ZN(n11104) );
  INV_X1 U13681 ( .A(n11104), .ZN(n11066) );
  OAI211_X1 U13682 ( .C1(n7148), .C2(n7147), .A(n6470), .B(n14715), .ZN(n11100) );
  AOI21_X1 U13683 ( .B1(n11100), .B2(n11055), .A(n14696), .ZN(n11061) );
  OAI22_X1 U13684 ( .A1(n14710), .A2(n11057), .B1(n11056), .B2(n14708), .ZN(
        n11058) );
  AOI21_X1 U13685 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n14710), .A(n11058), 
        .ZN(n11059) );
  OAI21_X1 U13686 ( .B1(n7148), .B2(n14739), .A(n11059), .ZN(n11060) );
  NOR2_X1 U13687 ( .A1(n11061), .A2(n11060), .ZN(n11065) );
  NAND2_X1 U13688 ( .A1(n11063), .A2(n13529), .ZN(n11099) );
  NAND3_X1 U13689 ( .A1(n11062), .A2(n11099), .A3(n14118), .ZN(n11064) );
  OAI211_X1 U13690 ( .C1(n11066), .C2(n14461), .A(n11065), .B(n11064), .ZN(
        P1_U3283) );
  INV_X1 U13691 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15217) );
  AOI21_X1 U13692 ( .B1(n15217), .B2(n11068), .A(n11401), .ZN(n11087) );
  MUX2_X1 U13693 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n6446), .Z(n11070) );
  NOR2_X1 U13694 ( .A1(n11070), .A2(n11069), .ZN(n11405) );
  INV_X1 U13695 ( .A(n11405), .ZN(n11071) );
  NAND2_X1 U13696 ( .A1(n11070), .A2(n11069), .ZN(n11407) );
  NAND2_X1 U13697 ( .A1(n11071), .A2(n11407), .ZN(n11076) );
  NAND2_X1 U13698 ( .A1(n11073), .A2(n11072), .ZN(n11075) );
  NAND2_X1 U13699 ( .A1(n11075), .A2(n11074), .ZN(n11406) );
  XNOR2_X1 U13700 ( .A(n11076), .B(n11406), .ZN(n11079) );
  NOR2_X1 U13701 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11077), .ZN(n12004) );
  AOI21_X1 U13702 ( .B1(n15087), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n12004), .ZN(
        n11078) );
  OAI21_X1 U13703 ( .B1(n15074), .B2(n11079), .A(n11078), .ZN(n11085) );
  AOI21_X1 U13704 ( .B1(n8760), .B2(n11082), .A(n11420), .ZN(n11083) );
  NOR2_X1 U13705 ( .A1(n11083), .A2(n15081), .ZN(n11084) );
  AOI211_X1 U13706 ( .C1(n15084), .C2(n11419), .A(n11085), .B(n11084), .ZN(
        n11086) );
  OAI21_X1 U13707 ( .B1(n11087), .B2(n15097), .A(n11086), .ZN(P3_U3191) );
  INV_X1 U13708 ( .A(n11088), .ZN(n11093) );
  AOI22_X1 U13709 ( .A1(n11090), .A2(n13291), .B1(n15019), .B2(n11089), .ZN(
        n11091) );
  OAI211_X1 U13710 ( .C1(n15023), .C2(n11093), .A(n11092), .B(n11091), .ZN(
        n11096) );
  NAND2_X1 U13711 ( .A1(n11096), .A2(n15047), .ZN(n11094) );
  OAI21_X1 U13712 ( .B1(n15047), .B2(n11095), .A(n11094), .ZN(P2_U3508) );
  INV_X1 U13713 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11098) );
  NAND2_X1 U13714 ( .A1(n11096), .A2(n15026), .ZN(n11097) );
  OAI21_X1 U13715 ( .B1(n15026), .B2(n11098), .A(n11097), .ZN(P2_U3457) );
  NAND3_X1 U13716 ( .A1(n11062), .A2(n11099), .A3(n14730), .ZN(n11102) );
  NAND3_X1 U13717 ( .A1(n11102), .A2(n11101), .A3(n11100), .ZN(n11103) );
  AOI21_X1 U13718 ( .B1(n14807), .B2(n11104), .A(n11103), .ZN(n11108) );
  AOI22_X1 U13719 ( .A1(n13618), .A2(n9609), .B1(n9605), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n11105) );
  OAI21_X1 U13720 ( .B1(n11108), .B2(n9605), .A(n11105), .ZN(P1_U3538) );
  OAI22_X1 U13721 ( .A1(n7148), .A2(n14282), .B1(n14810), .B2(n9279), .ZN(
        n11106) );
  INV_X1 U13722 ( .A(n11106), .ZN(n11107) );
  OAI21_X1 U13723 ( .B1(n11108), .B2(n14808), .A(n11107), .ZN(P1_U3489) );
  OR2_X1 U13724 ( .A1(n11109), .A2(n12092), .ZN(n11110) );
  NAND2_X1 U13725 ( .A1(n11111), .A2(n11110), .ZN(n15186) );
  OR2_X1 U13726 ( .A1(n11112), .A2(n15138), .ZN(n15183) );
  OAI22_X1 U13727 ( .A1(n11237), .A2(n15183), .B1(n11113), .B2(n15154), .ZN(
        n11122) );
  NAND2_X1 U13728 ( .A1(n11114), .A2(n12092), .ZN(n11115) );
  NAND3_X1 U13729 ( .A1(n11116), .A2(n15149), .A3(n11115), .ZN(n11120) );
  AOI22_X1 U13730 ( .A1(n15145), .A2(n12283), .B1(n11993), .B2(n15142), .ZN(
        n11119) );
  NAND2_X1 U13731 ( .A1(n15186), .A2(n11117), .ZN(n11118) );
  NAND3_X1 U13732 ( .A1(n11120), .A2(n11119), .A3(n11118), .ZN(n15184) );
  MUX2_X1 U13733 ( .A(n15184), .B(P3_REG2_REG_6__SCAN_IN), .S(n14498), .Z(
        n11121) );
  AOI211_X1 U13734 ( .C1(n11175), .C2(n15186), .A(n11122), .B(n11121), .ZN(
        n11123) );
  INV_X1 U13735 ( .A(n11123), .ZN(P3_U3227) );
  INV_X1 U13736 ( .A(n11124), .ZN(n11126) );
  OAI222_X1 U13737 ( .A1(n14318), .A2(n11125), .B1(n14312), .B2(n11126), .C1(
        n13929), .C2(P1_U3086), .ZN(P1_U3336) );
  OAI222_X1 U13738 ( .A1(n13372), .A2(n11127), .B1(n13367), .B2(n11126), .C1(
        P2_U3088), .C2(n13230), .ZN(P2_U3308) );
  INV_X1 U13739 ( .A(n12284), .ZN(n11129) );
  XNOR2_X1 U13740 ( .A(n11622), .B(n11916), .ZN(n11135) );
  XNOR2_X1 U13741 ( .A(n11135), .B(n12282), .ZN(n11131) );
  NAND2_X1 U13742 ( .A1(n11130), .A2(n11131), .ZN(n11139) );
  INV_X1 U13743 ( .A(n11131), .ZN(n11912) );
  INV_X1 U13744 ( .A(n11132), .ZN(n11133) );
  NAND2_X1 U13745 ( .A1(n11133), .A2(n12284), .ZN(n11874) );
  INV_X1 U13746 ( .A(n11876), .ZN(n11910) );
  OAI21_X1 U13747 ( .B1(n11912), .B2(n11874), .A(n11910), .ZN(n11138) );
  INV_X1 U13748 ( .A(n11135), .ZN(n11136) );
  XNOR2_X1 U13749 ( .A(n11622), .B(n11160), .ZN(n11140) );
  XNOR2_X1 U13750 ( .A(n11140), .B(n12281), .ZN(n12002) );
  INV_X1 U13751 ( .A(n11140), .ZN(n11141) );
  INV_X1 U13752 ( .A(n12281), .ZN(n11145) );
  NAND2_X1 U13753 ( .A1(n11141), .A2(n11145), .ZN(n11142) );
  AND2_X1 U13754 ( .A1(n11999), .A2(n11142), .ZN(n11144) );
  XNOR2_X1 U13755 ( .A(n11622), .B(n11147), .ZN(n11431) );
  XNOR2_X1 U13756 ( .A(n11431), .B(n12280), .ZN(n11143) );
  OAI211_X1 U13757 ( .C1(n11144), .C2(n11143), .A(n12041), .B(n11430), .ZN(
        n11149) );
  AND2_X1 U13758 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n15079) );
  OAI22_X1 U13759 ( .A1(n12052), .A2(n11145), .B1(n11435), .B2(n12065), .ZN(
        n11146) );
  AOI211_X1 U13760 ( .C1(n12036), .C2(n11147), .A(n15079), .B(n11146), .ZN(
        n11148) );
  OAI211_X1 U13761 ( .C1(n11235), .C2(n12028), .A(n11149), .B(n11148), .ZN(
        P3_U3157) );
  OAI222_X1 U13762 ( .A1(P3_U3151), .A2(n11151), .B1(n14434), .B2(n11150), 
        .C1(n15289), .C2(n11873), .ZN(P3_U3269) );
  XNOR2_X1 U13763 ( .A(n11152), .B(n12091), .ZN(n15196) );
  AND2_X1 U13764 ( .A1(n11155), .A2(n11153), .ZN(n11157) );
  NAND2_X1 U13765 ( .A1(n11155), .A2(n11154), .ZN(n11156) );
  OAI211_X1 U13766 ( .C1(n11157), .C2(n12091), .A(n11156), .B(n15149), .ZN(
        n11159) );
  AOI22_X1 U13767 ( .A1(n15142), .A2(n12282), .B1(n12280), .B2(n15145), .ZN(
        n11158) );
  OAI211_X1 U13768 ( .C1(n15153), .C2(n15196), .A(n11159), .B(n11158), .ZN(
        n15197) );
  NAND2_X1 U13769 ( .A1(n15197), .A2(n15159), .ZN(n11164) );
  NOR2_X1 U13770 ( .A1(n11160), .A2(n15138), .ZN(n15198) );
  INV_X1 U13771 ( .A(n15198), .ZN(n11161) );
  OAI22_X1 U13772 ( .A1(n11237), .A2(n11161), .B1(n12006), .B2(n15154), .ZN(
        n11162) );
  AOI21_X1 U13773 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n14498), .A(n11162), .ZN(
        n11163) );
  OAI211_X1 U13774 ( .C1(n15196), .C2(n15156), .A(n11164), .B(n11163), .ZN(
        P3_U3224) );
  XNOR2_X1 U13775 ( .A(n11166), .B(n11165), .ZN(n11172) );
  INV_X1 U13776 ( .A(n11172), .ZN(n15190) );
  OR2_X1 U13777 ( .A1(n11167), .A2(n15138), .ZN(n15187) );
  OAI22_X1 U13778 ( .A1(n11237), .A2(n15187), .B1(n11880), .B2(n15154), .ZN(
        n11174) );
  XNOR2_X1 U13779 ( .A(n11168), .B(n12156), .ZN(n11169) );
  NAND2_X1 U13780 ( .A1(n11169), .A2(n15149), .ZN(n11171) );
  AOI22_X1 U13781 ( .A1(n15142), .A2(n12284), .B1(n12282), .B2(n15145), .ZN(
        n11170) );
  OAI211_X1 U13782 ( .C1(n11172), .C2(n15153), .A(n11171), .B(n11170), .ZN(
        n15188) );
  MUX2_X1 U13783 ( .A(n15188), .B(P3_REG2_REG_7__SCAN_IN), .S(n14498), .Z(
        n11173) );
  AOI211_X1 U13784 ( .C1(n15190), .C2(n11175), .A(n11174), .B(n11173), .ZN(
        n11176) );
  INV_X1 U13785 ( .A(n11176), .ZN(P3_U3226) );
  XNOR2_X1 U13786 ( .A(n11704), .B(n11592), .ZN(n11244) );
  AND2_X1 U13787 ( .A1(n13226), .A2(n13194), .ZN(n11177) );
  NAND2_X1 U13788 ( .A1(n11244), .A2(n11177), .ZN(n11241) );
  OAI21_X1 U13789 ( .B1(n11244), .B2(n11177), .A(n11241), .ZN(n11183) );
  INV_X1 U13790 ( .A(n11178), .ZN(n11181) );
  AOI211_X1 U13791 ( .C1(n11183), .C2(n11182), .A(n12902), .B(n11243), .ZN(
        n11188) );
  INV_X1 U13792 ( .A(n11704), .ZN(n11393) );
  INV_X1 U13793 ( .A(n11184), .ZN(n11391) );
  AOI22_X1 U13794 ( .A1(n12888), .A2(n11391), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11186) );
  AOI22_X1 U13795 ( .A1(n12847), .A2(n12906), .B1(n12848), .B2(n13203), .ZN(
        n11185) );
  OAI211_X1 U13796 ( .C1(n11393), .C2(n12883), .A(n11186), .B(n11185), .ZN(
        n11187) );
  OR2_X1 U13797 ( .A1(n11188), .A2(n11187), .ZN(P2_U3206) );
  NAND2_X1 U13798 ( .A1(n15027), .A2(n11193), .ZN(n11189) );
  NAND2_X1 U13799 ( .A1(n11190), .A2(n11189), .ZN(n11192) );
  OAI21_X1 U13800 ( .B1(n11192), .B2(n11191), .A(n11215), .ZN(n11201) );
  INV_X1 U13801 ( .A(n12906), .ZN(n11360) );
  OAI22_X1 U13802 ( .A1(n11193), .A2(n13139), .B1(n11360), .B2(n13141), .ZN(
        n11200) );
  NAND2_X1 U13803 ( .A1(n11195), .A2(n11194), .ZN(n11197) );
  XNOR2_X1 U13804 ( .A(n11209), .B(n11198), .ZN(n11380) );
  NOR2_X1 U13805 ( .A1(n11380), .A2(n9771), .ZN(n11199) );
  AOI211_X1 U13806 ( .C1(n13228), .C2(n11201), .A(n11200), .B(n11199), .ZN(
        n11379) );
  AOI21_X1 U13807 ( .B1(n11376), .B2(n11202), .A(n11221), .ZN(n11377) );
  INV_X1 U13808 ( .A(n11203), .ZN(n11204) );
  AOI22_X1 U13809 ( .A1(n13212), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11204), 
        .B2(n13209), .ZN(n11205) );
  OAI21_X1 U13810 ( .B1(n7169), .B2(n13147), .A(n11205), .ZN(n11207) );
  NOR2_X1 U13811 ( .A1(n11380), .A2(n13072), .ZN(n11206) );
  AOI211_X1 U13812 ( .C1(n11377), .C2(n13131), .A(n11207), .B(n11206), .ZN(
        n11208) );
  OAI21_X1 U13813 ( .B1(n11379), .B2(n13212), .A(n11208), .ZN(P2_U3254) );
  OAI21_X1 U13814 ( .B1(n11209), .B2(n12907), .A(n11376), .ZN(n11211) );
  NAND2_X1 U13815 ( .A1(n11209), .A2(n12907), .ZN(n11210) );
  XNOR2_X1 U13816 ( .A(n11356), .B(n11216), .ZN(n14541) );
  INV_X1 U13817 ( .A(n14541), .ZN(n11228) );
  NAND2_X1 U13818 ( .A1(n14541), .A2(n11212), .ZN(n11220) );
  NAND2_X1 U13819 ( .A1(n11376), .A2(n11213), .ZN(n11214) );
  XNOR2_X1 U13820 ( .A(n11359), .B(n11216), .ZN(n11218) );
  AOI21_X1 U13821 ( .B1(n11218), .B2(n13228), .A(n11217), .ZN(n11219) );
  NAND2_X1 U13822 ( .A1(n11220), .A2(n11219), .ZN(n14546) );
  INV_X1 U13823 ( .A(n11361), .ZN(n14543) );
  OAI211_X1 U13824 ( .C1(n14543), .C2(n11221), .A(n13291), .B(n11365), .ZN(
        n14542) );
  NOR2_X1 U13825 ( .A1(n14542), .A2(n6914), .ZN(n11223) );
  OAI21_X1 U13826 ( .B1(n14546), .B2(n11223), .A(n13219), .ZN(n11227) );
  INV_X1 U13827 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11298) );
  OAI22_X1 U13828 ( .A1(n13219), .A2(n11298), .B1(n11224), .B2(n13217), .ZN(
        n11225) );
  AOI21_X1 U13829 ( .B1(n11361), .B2(n13234), .A(n11225), .ZN(n11226) );
  OAI211_X1 U13830 ( .C1(n11228), .C2(n13072), .A(n11227), .B(n11226), .ZN(
        P2_U3253) );
  OAI21_X1 U13831 ( .B1(n6585), .B2(n7225), .A(n11229), .ZN(n15200) );
  XNOR2_X1 U13832 ( .A(n11230), .B(n7225), .ZN(n11231) );
  NAND2_X1 U13833 ( .A1(n11231), .A2(n15149), .ZN(n11233) );
  AOI22_X1 U13834 ( .A1(n15145), .A2(n12279), .B1(n12281), .B2(n15142), .ZN(
        n11232) );
  OAI211_X1 U13835 ( .C1(n15153), .C2(n15200), .A(n11233), .B(n11232), .ZN(
        n15201) );
  NAND2_X1 U13836 ( .A1(n15201), .A2(n15159), .ZN(n11240) );
  NOR2_X1 U13837 ( .A1(n11234), .A2(n15138), .ZN(n15202) );
  INV_X1 U13838 ( .A(n15202), .ZN(n11236) );
  OAI22_X1 U13839 ( .A1(n11237), .A2(n11236), .B1(n11235), .B2(n15154), .ZN(
        n11238) );
  AOI21_X1 U13840 ( .B1(n14498), .B2(P3_REG2_REG_10__SCAN_IN), .A(n11238), 
        .ZN(n11239) );
  OAI211_X1 U13841 ( .C1(n15200), .C2(n15156), .A(n11240), .B(n11239), .ZN(
        P3_U3223) );
  XNOR2_X1 U13842 ( .A(n13323), .B(n6911), .ZN(n11551) );
  NAND2_X1 U13843 ( .A1(n13203), .A2(n13194), .ZN(n11550) );
  XNOR2_X1 U13844 ( .A(n11551), .B(n11550), .ZN(n11250) );
  INV_X1 U13845 ( .A(n11241), .ZN(n11242) );
  NAND3_X1 U13846 ( .A1(n11244), .A2(n12893), .A3(n13226), .ZN(n11245) );
  OAI21_X1 U13847 ( .B1(n6706), .B2(n12902), .A(n11245), .ZN(n11251) );
  INV_X1 U13848 ( .A(n13218), .ZN(n11246) );
  AOI22_X1 U13849 ( .A1(n12888), .A2(n11246), .B1(P2_REG3_REG_14__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11248) );
  AOI22_X1 U13850 ( .A1(n12848), .A2(n13224), .B1(n12847), .B2(n13226), .ZN(
        n11247) );
  OAI211_X1 U13851 ( .C1(n11730), .C2(n12883), .A(n11248), .B(n11247), .ZN(
        n11249) );
  AOI21_X1 U13852 ( .B1(n11251), .B2(n11250), .A(n11249), .ZN(n11252) );
  OAI21_X1 U13853 ( .B1(n6705), .B2(n12902), .A(n11252), .ZN(P2_U3187) );
  INV_X1 U13854 ( .A(n11253), .ZN(n11255) );
  INV_X1 U13855 ( .A(SI_27_), .ZN(n11254) );
  OAI222_X1 U13856 ( .A1(n14434), .A2(n11255), .B1(n14433), .B2(n11254), .C1(
        P3_U3151), .C2(n6446), .ZN(P3_U3268) );
  INV_X1 U13857 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n11256) );
  NAND2_X1 U13858 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13430)
         );
  OAI21_X1 U13859 ( .B1(n14677), .B2(n11256), .A(n13430), .ZN(n11264) );
  MUX2_X1 U13860 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n11257), .S(n13894), .Z(
        n13887) );
  AOI21_X1 U13861 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n11266), .A(n11258), 
        .ZN(n13888) );
  NAND2_X1 U13862 ( .A1(n13887), .A2(n13888), .ZN(n13886) );
  OAI21_X1 U13863 ( .B1(n13894), .B2(P1_REG1_REG_14__SCAN_IN), .A(n13886), 
        .ZN(n11259) );
  NAND2_X1 U13864 ( .A1(n11273), .A2(n11259), .ZN(n11260) );
  XNOR2_X1 U13865 ( .A(n14668), .B(n11259), .ZN(n14665) );
  NAND2_X1 U13866 ( .A1(n14665), .A2(n14664), .ZN(n14663) );
  NAND2_X1 U13867 ( .A1(n11260), .A2(n14663), .ZN(n11262) );
  XNOR2_X1 U13868 ( .A(n11456), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11261) );
  NOR2_X1 U13869 ( .A1(n11261), .A2(n11262), .ZN(n11455) );
  AOI211_X1 U13870 ( .C1(n11262), .C2(n11261), .A(n11455), .B(n13799), .ZN(
        n11263) );
  AOI211_X1 U13871 ( .C1(n14669), .C2(n11456), .A(n11264), .B(n11263), .ZN(
        n11280) );
  NAND2_X1 U13872 ( .A1(n13894), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11271) );
  MUX2_X1 U13873 ( .A(n9334), .B(P1_REG2_REG_14__SCAN_IN), .S(n13894), .Z(
        n11265) );
  INV_X1 U13874 ( .A(n11265), .ZN(n13892) );
  NAND2_X1 U13875 ( .A1(n11266), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11270) );
  OR2_X1 U13876 ( .A1(n11268), .A2(n11267), .ZN(n11269) );
  NAND2_X1 U13877 ( .A1(n11270), .A2(n11269), .ZN(n13893) );
  NAND2_X1 U13878 ( .A1(n13892), .A2(n13893), .ZN(n13891) );
  NAND2_X1 U13879 ( .A1(n11271), .A2(n13891), .ZN(n11272) );
  NOR2_X1 U13880 ( .A1(n14668), .A2(n11272), .ZN(n11274) );
  XOR2_X1 U13881 ( .A(n11273), .B(n11272), .Z(n14662) );
  NOR2_X1 U13882 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14662), .ZN(n14661) );
  NOR2_X1 U13883 ( .A1(n11274), .A2(n14661), .ZN(n11278) );
  NAND2_X1 U13884 ( .A1(n11456), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11450) );
  INV_X1 U13885 ( .A(n11450), .ZN(n11275) );
  AOI21_X1 U13886 ( .B1(n11536), .B2(n11276), .A(n11275), .ZN(n11277) );
  NAND2_X1 U13887 ( .A1(n11277), .A2(n11278), .ZN(n11449) );
  OAI211_X1 U13888 ( .C1(n11278), .C2(n11277), .A(n14656), .B(n11449), .ZN(
        n11279) );
  NAND2_X1 U13889 ( .A1(n11280), .A2(n11279), .ZN(P1_U3259) );
  NAND2_X1 U13890 ( .A1(n14823), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n11281) );
  NAND2_X1 U13891 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n12828)
         );
  NAND2_X1 U13892 ( .A1(n11281), .A2(n12828), .ZN(n11291) );
  INV_X1 U13893 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11285) );
  INV_X1 U13894 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11284) );
  NAND2_X1 U13895 ( .A1(n11292), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n11282) );
  NAND2_X1 U13896 ( .A1(n11283), .A2(n11282), .ZN(n14896) );
  MUX2_X1 U13897 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n11284), .S(n11295), .Z(
        n14895) );
  NAND2_X1 U13898 ( .A1(n14896), .A2(n14895), .ZN(n14894) );
  OAI21_X1 U13899 ( .B1(n14898), .B2(n11284), .A(n14894), .ZN(n14916) );
  MUX2_X1 U13900 ( .A(n11285), .B(P2_REG1_REG_12__SCAN_IN), .S(n11297), .Z(
        n14917) );
  NAND2_X1 U13901 ( .A1(n11300), .A2(n6713), .ZN(n11286) );
  OAI21_X1 U13902 ( .B1(n11300), .B2(n6713), .A(n11286), .ZN(n14926) );
  XNOR2_X1 U13903 ( .A(n14944), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n14940) );
  NOR2_X1 U13904 ( .A1(n14941), .A2(n14940), .ZN(n14939) );
  AOI21_X1 U13905 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n14944), .A(n14939), 
        .ZN(n11287) );
  XNOR2_X1 U13906 ( .A(n14970), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14961) );
  AOI21_X1 U13907 ( .B1(n14970), .B2(P2_REG1_REG_16__SCAN_IN), .A(n14959), 
        .ZN(n11289) );
  XNOR2_X1 U13908 ( .A(n12974), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n11288) );
  NOR2_X1 U13909 ( .A1(n11289), .A2(n11288), .ZN(n12973) );
  AOI211_X1 U13910 ( .C1(n11289), .C2(n11288), .A(n14960), .B(n12973), .ZN(
        n11290) );
  AOI211_X1 U13911 ( .C1(n14971), .C2(n12974), .A(n11291), .B(n11290), .ZN(
        n11316) );
  NAND2_X1 U13912 ( .A1(n11292), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n11293) );
  NAND2_X1 U13913 ( .A1(n11294), .A2(n11293), .ZN(n14900) );
  XNOR2_X1 U13914 ( .A(n11295), .B(P2_REG2_REG_11__SCAN_IN), .ZN(n14899) );
  OR2_X1 U13915 ( .A1(n11295), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n11296) );
  NAND2_X1 U13916 ( .A1(n14902), .A2(n11296), .ZN(n14913) );
  MUX2_X1 U13917 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n11298), .S(n11297), .Z(
        n14914) );
  NAND2_X1 U13918 ( .A1(n14913), .A2(n14914), .ZN(n14912) );
  NAND2_X1 U13919 ( .A1(n14909), .A2(n11298), .ZN(n11299) );
  NAND2_X1 U13920 ( .A1(n14912), .A2(n11299), .ZN(n14925) );
  NAND2_X1 U13921 ( .A1(n11300), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11301) );
  OAI21_X1 U13922 ( .B1(n11300), .B2(P2_REG2_REG_13__SCAN_IN), .A(n11301), 
        .ZN(n14924) );
  NAND2_X1 U13923 ( .A1(n14931), .A2(n11301), .ZN(n11302) );
  NOR2_X1 U13924 ( .A1(n11302), .A2(n14944), .ZN(n11303) );
  INV_X1 U13925 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n14938) );
  NOR2_X1 U13926 ( .A1(n14937), .A2(n14938), .ZN(n14936) );
  NOR2_X1 U13927 ( .A1(n11304), .A2(n14936), .ZN(n11305) );
  NOR2_X1 U13928 ( .A1(n11305), .A2(n11306), .ZN(n11307) );
  INV_X1 U13929 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n14949) );
  XNOR2_X1 U13930 ( .A(n11306), .B(n11305), .ZN(n14950) );
  NOR2_X1 U13931 ( .A1(n14949), .A2(n14950), .ZN(n14948) );
  NOR2_X1 U13932 ( .A1(n11307), .A2(n14948), .ZN(n14967) );
  INV_X1 U13933 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11308) );
  XNOR2_X1 U13934 ( .A(n11309), .B(n11308), .ZN(n14966) );
  NAND2_X1 U13935 ( .A1(n14970), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11310) );
  NAND2_X1 U13936 ( .A1(n14963), .A2(n11310), .ZN(n11314) );
  INV_X1 U13937 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13170) );
  OR2_X1 U13938 ( .A1(n12974), .A2(n13170), .ZN(n11312) );
  NAND2_X1 U13939 ( .A1(n12974), .A2(n13170), .ZN(n11311) );
  NAND2_X1 U13940 ( .A1(n11312), .A2(n11311), .ZN(n11313) );
  NAND2_X1 U13941 ( .A1(n11314), .A2(n11313), .ZN(n12968) );
  OAI211_X1 U13942 ( .C1(n11314), .C2(n11313), .A(n12968), .B(n14985), .ZN(
        n11315) );
  NAND2_X1 U13943 ( .A1(n11316), .A2(n11315), .ZN(P2_U3231) );
  OAI211_X1 U13944 ( .C1(n7146), .C2(n6598), .A(n14715), .B(n14458), .ZN(
        n14442) );
  INV_X1 U13945 ( .A(n14442), .ZN(n11323) );
  OAI211_X1 U13946 ( .C1(n11318), .C2(n7409), .A(n11317), .B(n14730), .ZN(
        n11322) );
  OR2_X1 U13947 ( .A1(n11471), .A2(n14734), .ZN(n11320) );
  OR2_X1 U13948 ( .A1(n13636), .A2(n13487), .ZN(n11319) );
  NAND2_X1 U13949 ( .A1(n11320), .A2(n11319), .ZN(n14555) );
  INV_X1 U13950 ( .A(n14555), .ZN(n11321) );
  NAND2_X1 U13951 ( .A1(n11322), .A2(n11321), .ZN(n14443) );
  AOI21_X1 U13952 ( .B1(n11323), .B2(n13929), .A(n14443), .ZN(n11330) );
  OAI21_X1 U13953 ( .B1(n11325), .B2(n13532), .A(n11324), .ZN(n14445) );
  NOR2_X1 U13954 ( .A1(n7146), .A2(n14739), .ZN(n11328) );
  OAI22_X1 U13955 ( .A1(n14691), .A2(n11326), .B1(n14557), .B2(n14708), .ZN(
        n11327) );
  AOI211_X1 U13956 ( .C1(n14445), .C2(n14042), .A(n11328), .B(n11327), .ZN(
        n11329) );
  OAI21_X1 U13957 ( .B1(n11330), .B2(n14710), .A(n11329), .ZN(P1_U3281) );
  INV_X1 U13958 ( .A(n11331), .ZN(n11332) );
  AOI21_X1 U13959 ( .B1(n12182), .B2(n11333), .A(n11332), .ZN(n14531) );
  NAND2_X1 U13960 ( .A1(n15153), .A2(n15133), .ZN(n14511) );
  NAND2_X1 U13961 ( .A1(n15159), .A2(n14511), .ZN(n12653) );
  INV_X1 U13962 ( .A(n12280), .ZN(n11432) );
  XNOR2_X1 U13963 ( .A(n11334), .B(n12182), .ZN(n11335) );
  OAI222_X1 U13964 ( .A1(n12642), .A2(n11432), .B1(n12646), .B2(n11620), .C1(
        n11335), .C2(n12582), .ZN(n14533) );
  NAND2_X1 U13965 ( .A1(n14533), .A2(n15159), .ZN(n11339) );
  OAI22_X1 U13966 ( .A1(n15159), .A2(n11336), .B1(n11440), .B2(n15154), .ZN(
        n11337) );
  AOI21_X1 U13967 ( .B1(n14499), .B2(n11436), .A(n11337), .ZN(n11338) );
  OAI211_X1 U13968 ( .C1(n14531), .C2(n12653), .A(n11339), .B(n11338), .ZN(
        P3_U3222) );
  OAI21_X1 U13969 ( .B1(n11341), .B2(n13530), .A(n11340), .ZN(n14577) );
  AOI211_X1 U13970 ( .C1(n14563), .C2(n6470), .A(n14788), .B(n6598), .ZN(
        n14570) );
  INV_X1 U13971 ( .A(n11342), .ZN(n11343) );
  AOI21_X1 U13972 ( .B1(n11343), .B2(n13530), .A(n14704), .ZN(n11348) );
  OR2_X1 U13973 ( .A1(n11344), .A2(n14734), .ZN(n11346) );
  OR2_X1 U13974 ( .A1(n11486), .A2(n13487), .ZN(n11345) );
  NAND2_X1 U13975 ( .A1(n11346), .A2(n11345), .ZN(n14567) );
  AOI21_X1 U13976 ( .B1(n11348), .B2(n11347), .A(n14567), .ZN(n14580) );
  INV_X1 U13977 ( .A(n14580), .ZN(n11349) );
  AOI211_X1 U13978 ( .C1(n14807), .C2(n14577), .A(n14570), .B(n11349), .ZN(
        n11354) );
  INV_X1 U13979 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11350) );
  OAI22_X1 U13980 ( .A1(n14575), .A2(n14282), .B1(n14810), .B2(n11350), .ZN(
        n11351) );
  INV_X1 U13981 ( .A(n11351), .ZN(n11352) );
  OAI21_X1 U13982 ( .B1(n11354), .B2(n14808), .A(n11352), .ZN(P1_U3492) );
  AOI22_X1 U13983 ( .A1(n14563), .A2(n9609), .B1(n9605), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n11353) );
  OAI21_X1 U13984 ( .B1(n11354), .B2(n9605), .A(n11353), .ZN(P1_U3539) );
  AND2_X1 U13985 ( .A1(n11361), .A2(n12906), .ZN(n11355) );
  OR2_X1 U13986 ( .A1(n11361), .A2(n12906), .ZN(n11357) );
  XNOR2_X1 U13987 ( .A(n11703), .B(n11363), .ZN(n11394) );
  OR2_X1 U13988 ( .A1(n11361), .A2(n11360), .ZN(n11358) );
  NAND2_X1 U13989 ( .A1(n11361), .A2(n11360), .ZN(n11362) );
  XNOR2_X1 U13990 ( .A(n11677), .B(n11363), .ZN(n11364) );
  AOI222_X1 U13991 ( .A1(n13228), .A2(n11364), .B1(n13203), .B2(n13223), .C1(
        n12906), .C2(n13225), .ZN(n11399) );
  AOI21_X1 U13992 ( .B1(n11704), .B2(n11365), .A(n6941), .ZN(n11397) );
  AOI22_X1 U13993 ( .A1(n11397), .A2(n13291), .B1(n15019), .B2(n11704), .ZN(
        n11366) );
  OAI211_X1 U13994 ( .C1(n13327), .C2(n11394), .A(n11399), .B(n11366), .ZN(
        n11368) );
  NAND2_X1 U13995 ( .A1(n11368), .A2(n15047), .ZN(n11367) );
  OAI21_X1 U13996 ( .B1(n15047), .B2(n6713), .A(n11367), .ZN(P2_U3512) );
  INV_X1 U13997 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11370) );
  NAND2_X1 U13998 ( .A1(n11368), .A2(n15026), .ZN(n11369) );
  OAI21_X1 U13999 ( .B1(n15026), .B2(n11370), .A(n11369), .ZN(P2_U3469) );
  INV_X1 U14000 ( .A(n11371), .ZN(n11374) );
  OAI222_X1 U14001 ( .A1(n13372), .A2(n11373), .B1(n13367), .B2(n11374), .C1(
        n11372), .C2(P2_U3088), .ZN(P2_U3307) );
  OAI222_X1 U14002 ( .A1(n14318), .A2(n11375), .B1(P1_U3086), .B2(n9590), .C1(
        n14312), .C2(n11374), .ZN(P1_U3335) );
  AOI22_X1 U14003 ( .A1(n11377), .A2(n13291), .B1(n15019), .B2(n11376), .ZN(
        n11378) );
  OAI211_X1 U14004 ( .C1(n11380), .C2(n15023), .A(n11379), .B(n11378), .ZN(
        n11382) );
  NAND2_X1 U14005 ( .A1(n11382), .A2(n15047), .ZN(n11381) );
  OAI21_X1 U14006 ( .B1(n15047), .B2(n11284), .A(n11381), .ZN(P2_U3510) );
  INV_X1 U14007 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11384) );
  NAND2_X1 U14008 ( .A1(n11382), .A2(n15026), .ZN(n11383) );
  OAI21_X1 U14009 ( .B1(n15026), .B2(n11384), .A(n11383), .ZN(P2_U3463) );
  XOR2_X1 U14010 ( .A(n12099), .B(n11385), .Z(n11386) );
  AOI222_X1 U14011 ( .A1(n15149), .A2(n11386), .B1(n12278), .B2(n15145), .C1(
        n12279), .C2(n15142), .ZN(n14527) );
  XNOR2_X1 U14012 ( .A(n11387), .B(n12099), .ZN(n14525) );
  NOR2_X1 U14013 ( .A1(n12650), .A2(n11619), .ZN(n11389) );
  OAI22_X1 U14014 ( .A1(n15159), .A2(n12301), .B1(n11942), .B2(n15154), .ZN(
        n11388) );
  AOI211_X1 U14015 ( .C1(n14525), .C2(n12635), .A(n11389), .B(n11388), .ZN(
        n11390) );
  OAI21_X1 U14016 ( .B1(n14527), .B2(n14498), .A(n11390), .ZN(P3_U3221) );
  AOI22_X1 U14017 ( .A1(n13212), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11391), 
        .B2(n13209), .ZN(n11392) );
  OAI21_X1 U14018 ( .B1(n11393), .B2(n13147), .A(n11392), .ZN(n11396) );
  NOR2_X1 U14019 ( .A1(n11394), .A2(n13236), .ZN(n11395) );
  AOI211_X1 U14020 ( .C1(n11397), .C2(n13131), .A(n11396), .B(n11395), .ZN(
        n11398) );
  OAI21_X1 U14021 ( .B1(n13212), .B2(n11399), .A(n11398), .ZN(P2_U3252) );
  NOR2_X1 U14022 ( .A1(n11419), .A2(n11400), .ZN(n11402) );
  NAND2_X1 U14023 ( .A1(n15067), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n11403) );
  OAI21_X1 U14024 ( .B1(n15067), .B2(P3_REG1_REG_10__SCAN_IN), .A(n11403), 
        .ZN(n15069) );
  AOI21_X1 U14025 ( .B1(n8798), .B2(n11404), .A(n12318), .ZN(n11429) );
  INV_X1 U14026 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n11417) );
  MUX2_X1 U14027 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n6446), .Z(n12307) );
  XNOR2_X1 U14028 ( .A(n12307), .B(n11423), .ZN(n11413) );
  INV_X1 U14029 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15220) );
  MUX2_X1 U14030 ( .A(n8777), .B(n15220), .S(n6446), .Z(n11410) );
  INV_X1 U14031 ( .A(n15067), .ZN(n11409) );
  NAND2_X1 U14032 ( .A1(n11410), .A2(n11409), .ZN(n11408) );
  INV_X1 U14033 ( .A(n11408), .ZN(n11411) );
  OAI21_X1 U14034 ( .B1(n11410), .B2(n11409), .A(n11408), .ZN(n15073) );
  AOI21_X1 U14035 ( .B1(n11413), .B2(n11412), .A(n12308), .ZN(n11414) );
  OR2_X1 U14036 ( .A1(n15074), .A2(n11414), .ZN(n11416) );
  INV_X1 U14037 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n15231) );
  NOR2_X1 U14038 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15231), .ZN(n11437) );
  INV_X1 U14039 ( .A(n11437), .ZN(n11415) );
  OAI211_X1 U14040 ( .C1(n15065), .C2(n11417), .A(n11416), .B(n11415), .ZN(
        n11427) );
  NOR2_X1 U14041 ( .A1(n11419), .A2(n11418), .ZN(n11421) );
  NAND2_X1 U14042 ( .A1(n15067), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n11422) );
  OAI21_X1 U14043 ( .B1(n15067), .B2(P3_REG2_REG_10__SCAN_IN), .A(n11422), 
        .ZN(n15063) );
  AOI21_X1 U14044 ( .B1(n11336), .B2(n11424), .A(n12299), .ZN(n11425) );
  NOR2_X1 U14045 ( .A1(n11425), .A2(n15081), .ZN(n11426) );
  AOI211_X1 U14046 ( .C1(n15084), .C2(n7166), .A(n11427), .B(n11426), .ZN(
        n11428) );
  OAI21_X1 U14047 ( .B1(n11429), .B2(n15097), .A(n11428), .ZN(P3_U3193) );
  INV_X1 U14048 ( .A(n11935), .ZN(n11433) );
  OAI21_X1 U14049 ( .B1(n11435), .B2(n11434), .A(n11433), .ZN(n11442) );
  AOI22_X1 U14050 ( .A1(n12062), .A2(n12280), .B1(n12036), .B2(n11436), .ZN(
        n11439) );
  AOI21_X1 U14051 ( .B1(n12050), .B2(n14508), .A(n11437), .ZN(n11438) );
  OAI211_X1 U14052 ( .C1(n12028), .C2(n11440), .A(n11439), .B(n11438), .ZN(
        n11441) );
  AOI21_X1 U14053 ( .B1(n11442), .B2(n12041), .A(n11441), .ZN(n11443) );
  INV_X1 U14054 ( .A(n11443), .ZN(P3_U3176) );
  INV_X1 U14055 ( .A(n11444), .ZN(n11447) );
  OAI222_X1 U14056 ( .A1(n13372), .A2(n11446), .B1(n13367), .B2(n11447), .C1(
        P2_U3088), .C2(n11445), .ZN(P2_U3306) );
  OAI222_X1 U14057 ( .A1(n14318), .A2(n11448), .B1(n14312), .B2(n11447), .C1(
        n13548), .C2(P1_U3086), .ZN(P1_U3334) );
  NAND2_X1 U14058 ( .A1(n11450), .A2(n11449), .ZN(n11453) );
  NOR2_X1 U14059 ( .A1(n13903), .A2(n14144), .ZN(n11451) );
  AOI21_X1 U14060 ( .B1(n14144), .B2(n13903), .A(n11451), .ZN(n11452) );
  NAND2_X1 U14061 ( .A1(n11452), .A2(n11453), .ZN(n13902) );
  OAI211_X1 U14062 ( .C1(n11453), .C2(n11452), .A(n14656), .B(n13902), .ZN(
        n11462) );
  INV_X1 U14063 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n11454) );
  NAND2_X1 U14064 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13442)
         );
  OAI21_X1 U14065 ( .B1(n14677), .B2(n11454), .A(n13442), .ZN(n11460) );
  AOI21_X1 U14066 ( .B1(n11456), .B2(P1_REG1_REG_16__SCAN_IN), .A(n11455), 
        .ZN(n11458) );
  XNOR2_X1 U14067 ( .A(n13906), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n11457) );
  NOR2_X1 U14068 ( .A1(n11458), .A2(n11457), .ZN(n13905) );
  AOI211_X1 U14069 ( .C1(n11458), .C2(n11457), .A(n13905), .B(n13799), .ZN(
        n11459) );
  AOI211_X1 U14070 ( .C1(n14669), .C2(n13906), .A(n11460), .B(n11459), .ZN(
        n11461) );
  NAND2_X1 U14071 ( .A1(n11462), .A2(n11461), .ZN(P1_U3260) );
  INV_X1 U14072 ( .A(n11465), .ZN(n11467) );
  NAND2_X1 U14073 ( .A1(n14563), .A2(n11826), .ZN(n11469) );
  OR2_X1 U14074 ( .A1(n11471), .A2(n11837), .ZN(n11468) );
  NAND2_X1 U14075 ( .A1(n11469), .A2(n11468), .ZN(n11470) );
  XNOR2_X1 U14076 ( .A(n11470), .B(n6473), .ZN(n11474) );
  NOR2_X1 U14077 ( .A1(n11836), .A2(n11471), .ZN(n11472) );
  AOI21_X1 U14078 ( .B1(n14563), .B2(n11827), .A(n11472), .ZN(n11473) );
  NAND2_X1 U14079 ( .A1(n11474), .A2(n11473), .ZN(n11475) );
  OAI21_X1 U14080 ( .B1(n11474), .B2(n11473), .A(n11475), .ZN(n14560) );
  INV_X1 U14081 ( .A(n11475), .ZN(n11476) );
  NOR2_X1 U14082 ( .A1(n11486), .A2(n11837), .ZN(n11477) );
  AOI21_X1 U14083 ( .B1(n14553), .B2(n11826), .A(n11477), .ZN(n11478) );
  XNOR2_X1 U14084 ( .A(n11478), .B(n11838), .ZN(n11480) );
  AOI22_X1 U14085 ( .A1(n14553), .A2(n11827), .B1(n11831), .B2(n13788), .ZN(
        n11479) );
  XNOR2_X1 U14086 ( .A(n11480), .B(n11479), .ZN(n14550) );
  NOR2_X1 U14087 ( .A1(n11836), .A2(n13636), .ZN(n11481) );
  AOI21_X1 U14088 ( .B1(n13638), .B2(n11827), .A(n11481), .ZN(n11738) );
  NOR2_X1 U14089 ( .A1(n13636), .A2(n11837), .ZN(n11482) );
  AOI21_X1 U14090 ( .B1(n13638), .B2(n11826), .A(n11482), .ZN(n11483) );
  XNOR2_X1 U14091 ( .A(n11483), .B(n11838), .ZN(n11737) );
  XOR2_X1 U14092 ( .A(n11738), .B(n11737), .Z(n11484) );
  OAI211_X1 U14093 ( .C1(n11485), .C2(n11484), .A(n11742), .B(n14564), .ZN(
        n11493) );
  INV_X1 U14094 ( .A(n14452), .ZN(n11491) );
  OR2_X1 U14095 ( .A1(n11486), .A2(n14734), .ZN(n11488) );
  NAND2_X1 U14096 ( .A1(n13786), .A2(n13479), .ZN(n11487) );
  AND2_X1 U14097 ( .A1(n11488), .A2(n11487), .ZN(n14450) );
  OAI21_X1 U14098 ( .B1(n15388), .B2(n14450), .A(n11489), .ZN(n11490) );
  AOI21_X1 U14099 ( .B1(n13481), .B2(n11491), .A(n11490), .ZN(n11492) );
  OAI211_X1 U14100 ( .C1(n6616), .C2(n15382), .A(n11493), .B(n11492), .ZN(
        P1_U3234) );
  OAI211_X1 U14101 ( .C1(n13644), .C2(n11495), .A(n11494), .B(n14730), .ZN(
        n11498) );
  OR2_X1 U14102 ( .A1(n11752), .A2(n13487), .ZN(n11497) );
  OR2_X1 U14103 ( .A1(n13636), .A2(n14734), .ZN(n11496) );
  AND2_X1 U14104 ( .A1(n11497), .A2(n11496), .ZN(n15387) );
  NAND2_X1 U14105 ( .A1(n11499), .A2(n13644), .ZN(n11500) );
  NAND2_X1 U14106 ( .A1(n11501), .A2(n11500), .ZN(n14583) );
  INV_X1 U14107 ( .A(n14583), .ZN(n11509) );
  INV_X1 U14108 ( .A(n14459), .ZN(n11502) );
  NOR2_X1 U14109 ( .A1(n15383), .A2(n11502), .ZN(n11503) );
  OR2_X1 U14110 ( .A1(n11503), .A2(n11517), .ZN(n14581) );
  NAND2_X1 U14111 ( .A1(n14710), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11504) );
  OAI21_X1 U14112 ( .B1(n14708), .B2(n15384), .A(n11504), .ZN(n11505) );
  AOI21_X1 U14113 ( .B1(n11506), .B2(n14694), .A(n11505), .ZN(n11507) );
  OAI21_X1 U14114 ( .B1(n14581), .B2(n14460), .A(n11507), .ZN(n11508) );
  AOI21_X1 U14115 ( .B1(n11509), .B2(n14578), .A(n11508), .ZN(n11510) );
  OAI21_X1 U14116 ( .B1(n14746), .B2(n14586), .A(n11510), .ZN(P1_U3279) );
  INV_X1 U14117 ( .A(n11511), .ZN(n11513) );
  OAI222_X1 U14118 ( .A1(P3_U3151), .A2(n9031), .B1(n14434), .B2(n11513), .C1(
        n11512), .C2(n11873), .ZN(P3_U3267) );
  OAI222_X1 U14119 ( .A1(n6439), .A2(P3_U3151), .B1(n11873), .B2(n11515), .C1(
        n14434), .C2(n11514), .ZN(P3_U3266) );
  XNOR2_X1 U14120 ( .A(n11516), .B(n13534), .ZN(n14246) );
  OAI211_X1 U14121 ( .C1(n11753), .C2(n11517), .A(n14715), .B(n11534), .ZN(
        n14251) );
  OR2_X1 U14122 ( .A1(n11518), .A2(n13534), .ZN(n14250) );
  NAND3_X1 U14123 ( .A1(n14250), .A2(n14249), .A3(n14118), .ZN(n11526) );
  NOR2_X1 U14124 ( .A1(n14691), .A2(n11519), .ZN(n11524) );
  OR2_X1 U14125 ( .A1(n13656), .A2(n13487), .ZN(n11521) );
  NAND2_X1 U14126 ( .A1(n13786), .A2(n13478), .ZN(n11520) );
  NAND2_X1 U14127 ( .A1(n11521), .A2(n11520), .ZN(n14247) );
  INV_X1 U14128 ( .A(n14247), .ZN(n11522) );
  OAI22_X1 U14129 ( .A1(n14710), .A2(n11522), .B1(n13497), .B2(n14708), .ZN(
        n11523) );
  AOI211_X1 U14130 ( .C1(n14248), .C2(n14694), .A(n11524), .B(n11523), .ZN(
        n11525) );
  OAI211_X1 U14131 ( .C1(n14251), .C2(n14696), .A(n11526), .B(n11525), .ZN(
        n11527) );
  AOI21_X1 U14132 ( .B1(n14578), .B2(n14246), .A(n11527), .ZN(n11528) );
  INV_X1 U14133 ( .A(n11528), .ZN(P1_U3278) );
  INV_X1 U14134 ( .A(n11529), .ZN(n11530) );
  AOI21_X1 U14135 ( .B1(n13535), .B2(n11531), .A(n11530), .ZN(n14245) );
  INV_X1 U14136 ( .A(n14118), .ZN(n14073) );
  OAI21_X1 U14137 ( .B1(n11533), .B2(n13535), .A(n11532), .ZN(n14243) );
  AOI21_X1 U14138 ( .B1(n13657), .B2(n11534), .A(n14788), .ZN(n11535) );
  NAND2_X1 U14139 ( .A1(n11535), .A2(n14143), .ZN(n14240) );
  NOR2_X1 U14140 ( .A1(n14691), .A2(n11536), .ZN(n11541) );
  OR2_X1 U14141 ( .A1(n11752), .A2(n14734), .ZN(n11538) );
  NAND2_X1 U14142 ( .A1(n13783), .A2(n13479), .ZN(n11537) );
  AND2_X1 U14143 ( .A1(n11538), .A2(n11537), .ZN(n14239) );
  INV_X1 U14144 ( .A(n13432), .ZN(n11539) );
  OAI22_X1 U14145 ( .A1(n14710), .A2(n14239), .B1(n11539), .B2(n14708), .ZN(
        n11540) );
  AOI211_X1 U14146 ( .C1(n13657), .C2(n14694), .A(n11541), .B(n11540), .ZN(
        n11542) );
  OAI21_X1 U14147 ( .B1(n14240), .B2(n14696), .A(n11542), .ZN(n11543) );
  AOI21_X1 U14148 ( .B1(n14243), .B2(n14578), .A(n11543), .ZN(n11544) );
  OAI21_X1 U14149 ( .B1(n14245), .B2(n14073), .A(n11544), .ZN(P1_U3277) );
  INV_X1 U14150 ( .A(n11545), .ZN(n13366) );
  OAI222_X1 U14151 ( .A1(n14318), .A2(n11547), .B1(n14312), .B2(n13366), .C1(
        P1_U3086), .C2(n11546), .ZN(P1_U3331) );
  INV_X1 U14152 ( .A(n11548), .ZN(n13354) );
  OAI222_X1 U14153 ( .A1(n14318), .A2(n11549), .B1(n14312), .B2(n13354), .C1(
        n13815), .C2(P1_U3086), .ZN(P1_U3327) );
  XNOR2_X1 U14154 ( .A(n13318), .B(n11592), .ZN(n11557) );
  AOI22_X1 U14155 ( .A1(n7059), .A2(n12871), .B1(n12893), .B2(n13224), .ZN(
        n11556) );
  AOI22_X1 U14156 ( .A1(n12847), .A2(n13203), .B1(n12848), .B2(n13204), .ZN(
        n11553) );
  AOI22_X1 U14157 ( .A1(n12888), .A2(n13208), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11552) );
  NAND2_X1 U14158 ( .A1(n11553), .A2(n11552), .ZN(n11554) );
  AOI21_X1 U14159 ( .B1(n13318), .B2(n12900), .A(n11554), .ZN(n11555) );
  OAI21_X1 U14160 ( .B1(n11560), .B2(n11556), .A(n11555), .ZN(P2_U3213) );
  XNOR2_X1 U14161 ( .A(n13307), .B(n11592), .ZN(n11563) );
  INV_X1 U14162 ( .A(n11563), .ZN(n11566) );
  NAND2_X1 U14163 ( .A1(n13186), .A2(n13194), .ZN(n11565) );
  AND2_X1 U14164 ( .A1(n11558), .A2(n11557), .ZN(n11559) );
  XNOR2_X1 U14165 ( .A(n13189), .B(n11592), .ZN(n12831) );
  NAND2_X1 U14166 ( .A1(n13204), .A2(n13194), .ZN(n11561) );
  XNOR2_X1 U14167 ( .A(n12831), .B(n11561), .ZN(n12821) );
  INV_X1 U14168 ( .A(n12831), .ZN(n11562) );
  NAND2_X1 U14169 ( .A1(n11562), .A2(n11561), .ZN(n11564) );
  XOR2_X1 U14170 ( .A(n11565), .B(n11563), .Z(n12835) );
  XNOR2_X1 U14171 ( .A(n13302), .B(n6911), .ZN(n12792) );
  NAND2_X1 U14172 ( .A1(n13165), .A2(n6444), .ZN(n11567) );
  NOR2_X1 U14173 ( .A1(n12792), .A2(n11567), .ZN(n11568) );
  AOI21_X1 U14174 ( .B1(n12792), .B2(n11567), .A(n11568), .ZN(n12873) );
  INV_X1 U14175 ( .A(n11568), .ZN(n11569) );
  XNOR2_X1 U14176 ( .A(n13298), .B(n11592), .ZN(n11570) );
  NAND2_X1 U14177 ( .A1(n13126), .A2(n13194), .ZN(n11571) );
  XNOR2_X1 U14178 ( .A(n11570), .B(n11571), .ZN(n12793) );
  INV_X1 U14179 ( .A(n11570), .ZN(n12852) );
  NAND2_X1 U14180 ( .A1(n12852), .A2(n11571), .ZN(n11572) );
  NAND2_X1 U14181 ( .A1(n13106), .A2(n13194), .ZN(n11573) );
  XOR2_X1 U14182 ( .A(n11573), .B(n11575), .Z(n12854) );
  INV_X1 U14183 ( .A(n11573), .ZN(n11574) );
  XNOR2_X1 U14184 ( .A(n13286), .B(n11592), .ZN(n11578) );
  NAND2_X1 U14185 ( .A1(n13127), .A2(n13194), .ZN(n11576) );
  XNOR2_X1 U14186 ( .A(n11578), .B(n11576), .ZN(n12802) );
  INV_X1 U14187 ( .A(n11576), .ZN(n11577) );
  NAND2_X1 U14188 ( .A1(n11578), .A2(n11577), .ZN(n11579) );
  XNOR2_X1 U14189 ( .A(n13280), .B(n11592), .ZN(n11581) );
  NAND2_X1 U14190 ( .A1(n11582), .A2(n11581), .ZN(n11583) );
  XNOR2_X1 U14191 ( .A(n13275), .B(n6911), .ZN(n11586) );
  NAND2_X1 U14192 ( .A1(n13087), .A2(n6444), .ZN(n12784) );
  NAND2_X1 U14193 ( .A1(n12785), .A2(n12784), .ZN(n11589) );
  XNOR2_X1 U14194 ( .A(n13269), .B(n11592), .ZN(n12811) );
  AND2_X1 U14195 ( .A1(n13074), .A2(n6444), .ZN(n11590) );
  NAND2_X1 U14196 ( .A1(n12811), .A2(n11590), .ZN(n11591) );
  OAI21_X1 U14197 ( .B1(n12811), .B2(n11590), .A(n11591), .ZN(n12840) );
  NAND2_X1 U14198 ( .A1(n12808), .A2(n11591), .ZN(n11597) );
  XNOR2_X1 U14199 ( .A(n13266), .B(n11592), .ZN(n12892) );
  AND2_X1 U14200 ( .A1(n13060), .A2(n6444), .ZN(n11593) );
  NAND2_X1 U14201 ( .A1(n12892), .A2(n11593), .ZN(n11598) );
  INV_X1 U14202 ( .A(n12892), .ZN(n11595) );
  INV_X1 U14203 ( .A(n11593), .ZN(n11594) );
  NAND2_X1 U14204 ( .A1(n11595), .A2(n11594), .ZN(n11596) );
  AND2_X1 U14205 ( .A1(n11598), .A2(n11596), .ZN(n12809) );
  NAND2_X1 U14206 ( .A1(n13012), .A2(n13194), .ZN(n11602) );
  XNOR2_X1 U14207 ( .A(n13259), .B(n11592), .ZN(n11601) );
  XOR2_X1 U14208 ( .A(n11602), .B(n11601), .Z(n12894) );
  INV_X1 U14209 ( .A(n11598), .ZN(n11599) );
  NOR2_X1 U14210 ( .A1(n12894), .A2(n11599), .ZN(n11600) );
  INV_X1 U14211 ( .A(n11601), .ZN(n11603) );
  NAND2_X1 U14212 ( .A1(n11603), .A2(n11602), .ZN(n11604) );
  XNOR2_X1 U14213 ( .A(n13255), .B(n11592), .ZN(n11606) );
  AND2_X1 U14214 ( .A1(n13027), .A2(n13194), .ZN(n11605) );
  NAND2_X1 U14215 ( .A1(n11606), .A2(n11605), .ZN(n11607) );
  OAI21_X1 U14216 ( .B1(n11606), .B2(n11605), .A(n11607), .ZN(n12777) );
  NAND2_X1 U14217 ( .A1(n13011), .A2(n13194), .ZN(n11608) );
  XNOR2_X1 U14218 ( .A(n11608), .B(n11592), .ZN(n11609) );
  XNOR2_X1 U14219 ( .A(n13250), .B(n11609), .ZN(n11610) );
  XNOR2_X1 U14220 ( .A(n11611), .B(n11610), .ZN(n11616) );
  AOI22_X1 U14221 ( .A1(n12905), .A2(n13223), .B1(n13027), .B2(n13225), .ZN(
        n13001) );
  AOI22_X1 U14222 ( .A1(n13006), .A2(n12888), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11612) );
  OAI21_X1 U14223 ( .B1(n13001), .B2(n11613), .A(n11612), .ZN(n11614) );
  AOI21_X1 U14224 ( .B1(n13250), .B2(n12900), .A(n11614), .ZN(n11615) );
  OAI21_X1 U14225 ( .B1(n11616), .B2(n12902), .A(n11615), .ZN(P2_U3192) );
  INV_X1 U14226 ( .A(n11617), .ZN(n11618) );
  OAI222_X1 U14227 ( .A1(n13372), .A2(n15239), .B1(n13367), .B2(n11618), .C1(
        n7762), .C2(P2_U3088), .ZN(P2_U3305) );
  XNOR2_X1 U14228 ( .A(n12616), .B(n11622), .ZN(n11951) );
  XNOR2_X1 U14229 ( .A(n11622), .B(n11619), .ZN(n11621) );
  XNOR2_X1 U14230 ( .A(n11621), .B(n11620), .ZN(n11933) );
  OAI21_X1 U14231 ( .B1(n11935), .B2(n11934), .A(n11933), .ZN(n11932) );
  XNOR2_X1 U14232 ( .A(n11643), .B(n14512), .ZN(n11624) );
  INV_X1 U14233 ( .A(n11624), .ZN(n11623) );
  AND2_X1 U14234 ( .A1(n11623), .A2(n12643), .ZN(n12019) );
  NAND2_X1 U14235 ( .A1(n11624), .A2(n12278), .ZN(n12020) );
  XNOR2_X1 U14236 ( .A(n12775), .B(n11622), .ZN(n11886) );
  XNOR2_X1 U14237 ( .A(n12067), .B(n11622), .ZN(n11625) );
  NAND2_X1 U14238 ( .A1(n11625), .A2(n12647), .ZN(n11626) );
  OAI21_X1 U14239 ( .B1(n11625), .B2(n12647), .A(n11626), .ZN(n12060) );
  XNOR2_X1 U14240 ( .A(n11971), .B(n11622), .ZN(n11628) );
  XNOR2_X1 U14241 ( .A(n11628), .B(n12583), .ZN(n11972) );
  XNOR2_X1 U14242 ( .A(n12040), .B(n11622), .ZN(n11631) );
  XNOR2_X1 U14243 ( .A(n11631), .B(n12596), .ZN(n12043) );
  XNOR2_X1 U14244 ( .A(n12756), .B(n11622), .ZN(n11636) );
  XNOR2_X1 U14245 ( .A(n11636), .B(n12584), .ZN(n11904) );
  NAND2_X1 U14246 ( .A1(n12043), .A2(n11904), .ZN(n11630) );
  INV_X1 U14247 ( .A(n11628), .ZN(n11629) );
  NAND2_X1 U14248 ( .A1(n11629), .A2(n12611), .ZN(n11901) );
  OR2_X1 U14249 ( .A1(n11630), .A2(n11901), .ZN(n11635) );
  INV_X1 U14250 ( .A(n11904), .ZN(n11633) );
  INV_X1 U14251 ( .A(n11631), .ZN(n11632) );
  NAND2_X1 U14252 ( .A1(n11632), .A2(n12596), .ZN(n11902) );
  OR2_X1 U14253 ( .A1(n11633), .A2(n11902), .ZN(n11634) );
  NAND2_X1 U14254 ( .A1(n11636), .A2(n12277), .ZN(n11637) );
  XNOR2_X1 U14255 ( .A(n12223), .B(n11622), .ZN(n11638) );
  XNOR2_X1 U14256 ( .A(n11638), .B(n12568), .ZN(n12013) );
  INV_X1 U14257 ( .A(n11638), .ZN(n11639) );
  NAND2_X1 U14258 ( .A1(n11639), .A2(n12568), .ZN(n11640) );
  XNOR2_X1 U14259 ( .A(n12690), .B(n11622), .ZN(n11641) );
  XNOR2_X1 U14260 ( .A(n11641), .B(n12556), .ZN(n11925) );
  NAND2_X1 U14261 ( .A1(n11641), .A2(n12556), .ZN(n11642) );
  XNOR2_X1 U14262 ( .A(n12037), .B(n11643), .ZN(n11644) );
  INV_X1 U14263 ( .A(n11644), .ZN(n11645) );
  XNOR2_X1 U14264 ( .A(n12680), .B(n11622), .ZN(n11646) );
  NAND2_X1 U14265 ( .A1(n11895), .A2(n12533), .ZN(n11650) );
  INV_X1 U14266 ( .A(n11646), .ZN(n11647) );
  OR2_X1 U14267 ( .A1(n11648), .A2(n11647), .ZN(n11649) );
  XNOR2_X1 U14268 ( .A(n12676), .B(n11622), .ZN(n11651) );
  XNOR2_X1 U14269 ( .A(n11651), .B(n12521), .ZN(n11982) );
  NAND2_X1 U14270 ( .A1(n11651), .A2(n11946), .ZN(n11652) );
  XNOR2_X1 U14271 ( .A(n12739), .B(n11622), .ZN(n11653) );
  XNOR2_X1 U14272 ( .A(n11653), .B(n12484), .ZN(n11944) );
  INV_X1 U14273 ( .A(n11653), .ZN(n11654) );
  NAND2_X1 U14274 ( .A1(n11654), .A2(n12484), .ZN(n11655) );
  XNOR2_X1 U14275 ( .A(n12735), .B(n11622), .ZN(n11656) );
  XNOR2_X1 U14276 ( .A(n11656), .B(n12497), .ZN(n12049) );
  INV_X1 U14277 ( .A(n11656), .ZN(n11657) );
  XNOR2_X1 U14278 ( .A(n12477), .B(n11622), .ZN(n11663) );
  XNOR2_X1 U14279 ( .A(n11663), .B(n7249), .ZN(n11665) );
  XNOR2_X1 U14280 ( .A(n11666), .B(n11665), .ZN(n11658) );
  NAND2_X1 U14281 ( .A1(n11658), .A2(n12041), .ZN(n11662) );
  AOI22_X1 U14282 ( .A1(n12274), .A2(n12062), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11659) );
  OAI21_X1 U14283 ( .B1(n12472), .B2(n12065), .A(n11659), .ZN(n11660) );
  AOI21_X1 U14284 ( .B1(n12476), .B2(n12071), .A(n11660), .ZN(n11661) );
  OAI211_X1 U14285 ( .C1(n12731), .C2(n12068), .A(n11662), .B(n11661), .ZN(
        P3_U3154) );
  AOI21_X1 U14286 ( .B1(n11666), .B2(n11665), .A(n11664), .ZN(n11668) );
  XNOR2_X1 U14287 ( .A(n12461), .B(n11622), .ZN(n11667) );
  XNOR2_X1 U14288 ( .A(n11668), .B(n11667), .ZN(n11674) );
  AOI22_X1 U14289 ( .A1(n7249), .A2(n12062), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11669) );
  OAI21_X1 U14290 ( .B1(n12458), .B2(n12065), .A(n11669), .ZN(n11672) );
  NOR2_X1 U14291 ( .A1(n11670), .A2(n12068), .ZN(n11671) );
  AOI211_X1 U14292 ( .C1(n12463), .C2(n12071), .A(n11672), .B(n11671), .ZN(
        n11673) );
  OAI21_X1 U14293 ( .B1(n11674), .B2(n12073), .A(n11673), .ZN(P3_U3160) );
  INV_X1 U14294 ( .A(n13074), .ZN(n13044) );
  INV_X1 U14295 ( .A(n11675), .ZN(n11676) );
  OR2_X1 U14296 ( .A1(n13318), .A2(n11680), .ZN(n11682) );
  AND2_X1 U14297 ( .A1(n13318), .A2(n11680), .ZN(n11681) );
  NAND2_X1 U14298 ( .A1(n13185), .A2(n13184), .ZN(n13183) );
  INV_X1 U14299 ( .A(n13204), .ZN(n12833) );
  OR2_X1 U14300 ( .A1(n13189), .A2(n12833), .ZN(n11683) );
  NAND2_X1 U14301 ( .A1(n13183), .A2(n11683), .ZN(n13164) );
  INV_X1 U14302 ( .A(n13186), .ZN(n11685) );
  NAND2_X1 U14303 ( .A1(n13307), .A2(n11685), .ZN(n11684) );
  NAND2_X1 U14304 ( .A1(n13164), .A2(n11684), .ZN(n11687) );
  OR2_X1 U14305 ( .A1(n13307), .A2(n11685), .ZN(n11686) );
  NAND2_X1 U14306 ( .A1(n13302), .A2(n13138), .ZN(n11688) );
  INV_X1 U14307 ( .A(n13126), .ZN(n12851) );
  AND2_X1 U14308 ( .A1(n13298), .A2(n12851), .ZN(n11689) );
  OR2_X1 U14309 ( .A1(n13286), .A2(n12865), .ZN(n11692) );
  AND2_X1 U14310 ( .A1(n13286), .A2(n12865), .ZN(n11691) );
  AOI21_X1 U14311 ( .B1(n13103), .B2(n11692), .A(n11691), .ZN(n13086) );
  NAND2_X1 U14312 ( .A1(n13091), .A2(n13086), .ZN(n13085) );
  NAND2_X1 U14313 ( .A1(n13085), .A2(n11693), .ZN(n13073) );
  NAND2_X1 U14314 ( .A1(n13275), .A2(n12866), .ZN(n11695) );
  NOR2_X1 U14315 ( .A1(n13275), .A2(n12866), .ZN(n11694) );
  INV_X1 U14316 ( .A(n13012), .ZN(n13043) );
  INV_X1 U14317 ( .A(n13259), .ZN(n13033) );
  INV_X1 U14318 ( .A(n13027), .ZN(n12891) );
  XNOR2_X1 U14319 ( .A(n11696), .B(n11725), .ZN(n11701) );
  NOR2_X1 U14320 ( .A1(n13356), .A2(n11697), .ZN(n11698) );
  NOR2_X1 U14321 ( .A1(n13141), .A2(n11698), .ZN(n12985) );
  AOI21_X2 U14322 ( .B1(n11701), .B2(n13228), .A(n11700), .ZN(n13247) );
  NOR2_X1 U14323 ( .A1(n11704), .A2(n13226), .ZN(n11702) );
  NAND2_X1 U14324 ( .A1(n11704), .A2(n13226), .ZN(n11705) );
  NAND2_X1 U14325 ( .A1(n13216), .A2(n13215), .ZN(n11707) );
  NAND2_X1 U14326 ( .A1(n13323), .A2(n13203), .ZN(n11706) );
  INV_X1 U14327 ( .A(n13199), .ZN(n13202) );
  OR2_X1 U14328 ( .A1(n13318), .A2(n13224), .ZN(n11708) );
  NAND2_X1 U14329 ( .A1(n13189), .A2(n13204), .ZN(n11711) );
  NAND2_X1 U14330 ( .A1(n13307), .A2(n13186), .ZN(n11713) );
  INV_X1 U14331 ( .A(n13154), .ZN(n13152) );
  NOR2_X1 U14332 ( .A1(n13290), .A2(n13106), .ZN(n11717) );
  INV_X1 U14333 ( .A(n13290), .ZN(n13122) );
  INV_X1 U14334 ( .A(n13112), .ZN(n13104) );
  OR2_X1 U14335 ( .A1(n13286), .A2(n13127), .ZN(n11718) );
  NAND2_X1 U14336 ( .A1(n13280), .A2(n13105), .ZN(n11719) );
  INV_X1 U14337 ( .A(n11720), .ZN(n11722) );
  AND2_X1 U14338 ( .A1(n13259), .A2(n13012), .ZN(n11723) );
  OAI22_X1 U14339 ( .A1(n11728), .A2(n13217), .B1(n11727), .B2(n13219), .ZN(
        n11729) );
  AOI21_X1 U14340 ( .B1(n13244), .B2(n13234), .A(n11729), .ZN(n11734) );
  INV_X1 U14341 ( .A(n13250), .ZN(n13003) );
  INV_X1 U14342 ( .A(n13307), .ZN(n13172) );
  INV_X1 U14343 ( .A(n13266), .ZN(n13050) );
  OR2_X2 U14344 ( .A1(n13244), .A2(n13005), .ZN(n12991) );
  NAND2_X1 U14345 ( .A1(n13244), .A2(n13005), .ZN(n11732) );
  NAND2_X1 U14346 ( .A1(n13245), .A2(n13131), .ZN(n11733) );
  OAI211_X1 U14347 ( .C1(n13248), .C2(n13236), .A(n11734), .B(n11733), .ZN(
        n11735) );
  INV_X1 U14348 ( .A(n11735), .ZN(n11736) );
  OAI21_X1 U14349 ( .B1(n13247), .B2(n13212), .A(n11736), .ZN(P2_U3236) );
  INV_X1 U14350 ( .A(n11738), .ZN(n11739) );
  NAND2_X1 U14351 ( .A1(n11740), .A2(n11739), .ZN(n11741) );
  OAI22_X1 U14352 ( .A1(n15383), .A2(n11835), .B1(n11744), .B2(n11837), .ZN(
        n11743) );
  INV_X2 U14353 ( .A(n6473), .ZN(n11838) );
  XNOR2_X1 U14354 ( .A(n11743), .B(n11838), .ZN(n11747) );
  OAI22_X1 U14355 ( .A1(n15383), .A2(n11837), .B1(n11744), .B2(n11836), .ZN(
        n11746) );
  XNOR2_X1 U14356 ( .A(n11747), .B(n11746), .ZN(n15377) );
  OAI22_X1 U14357 ( .A1(n11753), .A2(n11835), .B1(n11752), .B2(n11837), .ZN(
        n11749) );
  XOR2_X1 U14358 ( .A(n11838), .B(n11749), .Z(n11750) );
  OAI22_X1 U14359 ( .A1(n11753), .A2(n11837), .B1(n11752), .B2(n11836), .ZN(
        n13495) );
  INV_X1 U14360 ( .A(n13495), .ZN(n11754) );
  NAND2_X1 U14361 ( .A1(n13492), .A2(n11755), .ZN(n13427) );
  INV_X1 U14362 ( .A(n13657), .ZN(n14241) );
  OAI22_X1 U14363 ( .A1(n14241), .A2(n11837), .B1(n13656), .B2(n11836), .ZN(
        n11759) );
  NAND2_X1 U14364 ( .A1(n13657), .A2(n11826), .ZN(n11757) );
  OR2_X1 U14365 ( .A1(n13656), .A2(n11837), .ZN(n11756) );
  NAND2_X1 U14366 ( .A1(n11757), .A2(n11756), .ZN(n11758) );
  XNOR2_X1 U14367 ( .A(n11758), .B(n11838), .ZN(n11760) );
  XOR2_X1 U14368 ( .A(n11759), .B(n11760), .Z(n13428) );
  NAND2_X1 U14369 ( .A1(n13427), .A2(n13428), .ZN(n13426) );
  NAND2_X1 U14370 ( .A1(n13426), .A2(n11761), .ZN(n13436) );
  NAND2_X1 U14371 ( .A1(n14235), .A2(n11826), .ZN(n11763) );
  NAND2_X1 U14372 ( .A1(n13783), .A2(n11827), .ZN(n11762) );
  NAND2_X1 U14373 ( .A1(n11763), .A2(n11762), .ZN(n11764) );
  XNOR2_X1 U14374 ( .A(n11764), .B(n11838), .ZN(n11767) );
  NAND2_X1 U14375 ( .A1(n14235), .A2(n11827), .ZN(n11766) );
  NAND2_X1 U14376 ( .A1(n11831), .A2(n13783), .ZN(n11765) );
  NAND2_X1 U14377 ( .A1(n11766), .A2(n11765), .ZN(n11768) );
  NAND2_X1 U14378 ( .A1(n11767), .A2(n11768), .ZN(n13437) );
  NAND2_X1 U14379 ( .A1(n13436), .A2(n13437), .ZN(n13435) );
  INV_X1 U14380 ( .A(n11767), .ZN(n11770) );
  INV_X1 U14381 ( .A(n11768), .ZN(n11769) );
  NAND2_X1 U14382 ( .A1(n11770), .A2(n11769), .ZN(n13439) );
  NAND2_X1 U14383 ( .A1(n13435), .A2(n13439), .ZN(n13474) );
  OAI22_X1 U14384 ( .A1(n14132), .A2(n11837), .B1(n13672), .B2(n11836), .ZN(
        n11774) );
  NAND2_X1 U14385 ( .A1(n14230), .A2(n11826), .ZN(n11772) );
  NAND2_X1 U14386 ( .A1(n13782), .A2(n11827), .ZN(n11771) );
  NAND2_X1 U14387 ( .A1(n11772), .A2(n11771), .ZN(n11773) );
  XNOR2_X1 U14388 ( .A(n11773), .B(n11838), .ZN(n11775) );
  XOR2_X1 U14389 ( .A(n11774), .B(n11775), .Z(n13475) );
  AND2_X1 U14390 ( .A1(n13781), .A2(n11831), .ZN(n11777) );
  AOI21_X1 U14391 ( .B1(n14290), .B2(n11827), .A(n11777), .ZN(n11783) );
  NAND2_X1 U14392 ( .A1(n14290), .A2(n11826), .ZN(n11779) );
  NAND2_X1 U14393 ( .A1(n13781), .A2(n11827), .ZN(n11778) );
  NAND2_X1 U14394 ( .A1(n11779), .A2(n11778), .ZN(n11780) );
  XNOR2_X1 U14395 ( .A(n11780), .B(n11838), .ZN(n11782) );
  XOR2_X1 U14396 ( .A(n11783), .B(n11782), .Z(n13399) );
  INV_X1 U14397 ( .A(n11782), .ZN(n11784) );
  INV_X1 U14398 ( .A(n14215), .ZN(n13684) );
  OAI22_X1 U14399 ( .A1(n13684), .A2(n11835), .B1(n13685), .B2(n11837), .ZN(
        n11785) );
  XNOR2_X1 U14400 ( .A(n11785), .B(n11838), .ZN(n11787) );
  AND2_X1 U14401 ( .A1(n13780), .A2(n11831), .ZN(n11786) );
  AOI21_X1 U14402 ( .B1(n14215), .B2(n11827), .A(n11786), .ZN(n11788) );
  XNOR2_X1 U14403 ( .A(n11787), .B(n11788), .ZN(n13455) );
  INV_X1 U14404 ( .A(n11787), .ZN(n11789) );
  AOI22_X1 U14405 ( .A1(n14285), .A2(n11826), .B1(n11827), .B2(n13779), .ZN(
        n11790) );
  XNOR2_X1 U14406 ( .A(n11790), .B(n11838), .ZN(n11792) );
  AOI22_X1 U14407 ( .A1(n14285), .A2(n11827), .B1(n11831), .B2(n13779), .ZN(
        n11793) );
  XNOR2_X1 U14408 ( .A(n11792), .B(n11793), .ZN(n13410) );
  INV_X1 U14409 ( .A(n13410), .ZN(n11791) );
  OR2_X1 U14410 ( .A1(n14281), .A2(n11837), .ZN(n11795) );
  NAND2_X1 U14411 ( .A1(n11831), .A2(n13778), .ZN(n11794) );
  NAND2_X1 U14412 ( .A1(n11795), .A2(n11794), .ZN(n11797) );
  OAI22_X1 U14413 ( .A1(n14281), .A2(n11835), .B1(n7138), .B2(n11837), .ZN(
        n11796) );
  XNOR2_X1 U14414 ( .A(n11796), .B(n11838), .ZN(n11798) );
  XOR2_X1 U14415 ( .A(n11797), .B(n11798), .Z(n13465) );
  NAND2_X1 U14416 ( .A1(n14049), .A2(n11826), .ZN(n11801) );
  NAND2_X1 U14417 ( .A1(n11827), .A2(n13777), .ZN(n11800) );
  NAND2_X1 U14418 ( .A1(n11801), .A2(n11800), .ZN(n11802) );
  XNOR2_X1 U14419 ( .A(n11802), .B(n11838), .ZN(n11805) );
  AOI22_X1 U14420 ( .A1(n14049), .A2(n11827), .B1(n11831), .B2(n13777), .ZN(
        n11803) );
  XNOR2_X1 U14421 ( .A(n11805), .B(n11803), .ZN(n13382) );
  INV_X1 U14422 ( .A(n11803), .ZN(n11804) );
  OR2_X1 U14423 ( .A1(n11805), .A2(n11804), .ZN(n11806) );
  NAND2_X1 U14424 ( .A1(n14272), .A2(n11826), .ZN(n11808) );
  NAND2_X1 U14425 ( .A1(n11827), .A2(n13776), .ZN(n11807) );
  NAND2_X1 U14426 ( .A1(n11808), .A2(n11807), .ZN(n11809) );
  XNOR2_X1 U14427 ( .A(n11809), .B(n11838), .ZN(n11812) );
  AOI22_X1 U14428 ( .A1(n14272), .A2(n11827), .B1(n11831), .B2(n13776), .ZN(
        n11810) );
  XNOR2_X1 U14429 ( .A(n11812), .B(n11810), .ZN(n13447) );
  INV_X1 U14430 ( .A(n11810), .ZN(n11811) );
  NAND2_X1 U14431 ( .A1(n14268), .A2(n11826), .ZN(n11814) );
  OR2_X1 U14432 ( .A1(n13486), .A2(n11837), .ZN(n11813) );
  NAND2_X1 U14433 ( .A1(n11814), .A2(n11813), .ZN(n11815) );
  XNOR2_X1 U14434 ( .A(n11815), .B(n11838), .ZN(n11816) );
  AOI22_X1 U14435 ( .A1(n14268), .A2(n11827), .B1(n11831), .B2(n13775), .ZN(
        n11817) );
  XNOR2_X1 U14436 ( .A(n11816), .B(n11817), .ZN(n13418) );
  INV_X1 U14437 ( .A(n11816), .ZN(n11818) );
  OAI22_X1 U14438 ( .A1(n14005), .A2(n11837), .B1(n13419), .B2(n11836), .ZN(
        n11823) );
  NAND2_X1 U14439 ( .A1(n14171), .A2(n11826), .ZN(n11820) );
  OR2_X1 U14440 ( .A1(n13419), .A2(n11837), .ZN(n11819) );
  NAND2_X1 U14441 ( .A1(n11820), .A2(n11819), .ZN(n11821) );
  XNOR2_X1 U14442 ( .A(n11821), .B(n11838), .ZN(n11822) );
  XOR2_X1 U14443 ( .A(n11823), .B(n11822), .Z(n13485) );
  INV_X1 U14444 ( .A(n11822), .ZN(n11825) );
  INV_X1 U14445 ( .A(n11823), .ZN(n11824) );
  NAND2_X1 U14446 ( .A1(n14165), .A2(n11826), .ZN(n11829) );
  NAND2_X1 U14447 ( .A1(n11827), .A2(n13773), .ZN(n11828) );
  NAND2_X1 U14448 ( .A1(n11829), .A2(n11828), .ZN(n11830) );
  XNOR2_X1 U14449 ( .A(n11830), .B(n11838), .ZN(n11832) );
  AOI22_X1 U14450 ( .A1(n14165), .A2(n11827), .B1(n11831), .B2(n13773), .ZN(
        n11833) );
  XNOR2_X1 U14451 ( .A(n11832), .B(n11833), .ZN(n13376) );
  INV_X1 U14452 ( .A(n11832), .ZN(n11834) );
  OAI22_X1 U14453 ( .A1(n14263), .A2(n11835), .B1(n13377), .B2(n11837), .ZN(
        n11841) );
  OAI22_X1 U14454 ( .A1(n14263), .A2(n11837), .B1(n13377), .B2(n11836), .ZN(
        n11839) );
  XNOR2_X1 U14455 ( .A(n11839), .B(n11838), .ZN(n11840) );
  XOR2_X1 U14456 ( .A(n11841), .B(n11840), .Z(n11842) );
  NAND2_X1 U14457 ( .A1(n13772), .A2(n13479), .ZN(n11844) );
  NAND2_X1 U14458 ( .A1(n13773), .A2(n13478), .ZN(n11843) );
  AND2_X1 U14459 ( .A1(n11844), .A2(n11843), .ZN(n14157) );
  INV_X1 U14460 ( .A(n14157), .ZN(n11845) );
  AOI22_X1 U14461 ( .A1(n14566), .A2(n11845), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11846) );
  OAI21_X1 U14462 ( .B1(n15385), .B2(n13970), .A(n11846), .ZN(n11847) );
  AOI21_X1 U14463 ( .B1(n13968), .B2(n14562), .A(n11847), .ZN(n11848) );
  OAI21_X1 U14464 ( .B1(n11849), .B2(n15379), .A(n11848), .ZN(P1_U3220) );
  INV_X1 U14465 ( .A(n13512), .ZN(n11862) );
  INV_X1 U14466 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13513) );
  OAI222_X1 U14467 ( .A1(n14312), .A2(n11862), .B1(P1_U3086), .B2(n9148), .C1(
        n13513), .C2(n14318), .ZN(P1_U3325) );
  NAND3_X1 U14468 ( .A1(n11850), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n11859) );
  NAND2_X1 U14469 ( .A1(n14304), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11851) );
  NAND2_X1 U14470 ( .A1(n11852), .A2(n11851), .ZN(n11869) );
  XNOR2_X1 U14471 ( .A(n11861), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n11868) );
  XNOR2_X1 U14472 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n11853) );
  XNOR2_X1 U14473 ( .A(n11854), .B(n11853), .ZN(n12080) );
  NAND2_X1 U14474 ( .A1(n12080), .A2(n11855), .ZN(n11858) );
  NAND2_X1 U14475 ( .A1(n11856), .A2(SI_31_), .ZN(n11857) );
  OAI211_X1 U14476 ( .C1(n11860), .C2(n11859), .A(n11858), .B(n11857), .ZN(
        P3_U3264) );
  OAI222_X1 U14477 ( .A1(n13357), .A2(n11862), .B1(P2_U3088), .B2(n7757), .C1(
        n11861), .C2(n13372), .ZN(P2_U3297) );
  NAND2_X1 U14478 ( .A1(n11863), .A2(n15136), .ZN(n12451) );
  OAI21_X1 U14479 ( .B1(n15159), .B2(n15246), .A(n12451), .ZN(n11865) );
  INV_X1 U14480 ( .A(SI_30_), .ZN(n11872) );
  XNOR2_X1 U14481 ( .A(n11869), .B(n11868), .ZN(n12075) );
  INV_X1 U14482 ( .A(n12075), .ZN(n11870) );
  OAI222_X1 U14483 ( .A1(n11873), .A2(n11872), .B1(P3_U3151), .B2(n11871), 
        .C1(n14434), .C2(n11870), .ZN(P3_U3265) );
  NAND2_X1 U14484 ( .A1(n11875), .A2(n11874), .ZN(n11911) );
  XNOR2_X1 U14485 ( .A(n11911), .B(n11876), .ZN(n11877) );
  NAND2_X1 U14486 ( .A1(n11877), .A2(n12041), .ZN(n11885) );
  NOR2_X1 U14487 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11878), .ZN(n15048) );
  AOI21_X1 U14488 ( .B1(n12036), .B2(n11879), .A(n15048), .ZN(n11884) );
  AOI22_X1 U14489 ( .A1(n12050), .A2(n12282), .B1(n12062), .B2(n12284), .ZN(
        n11883) );
  INV_X1 U14490 ( .A(n11880), .ZN(n11881) );
  NAND2_X1 U14491 ( .A1(n12071), .A2(n11881), .ZN(n11882) );
  NAND4_X1 U14492 ( .A1(n11885), .A2(n11884), .A3(n11883), .A4(n11882), .ZN(
        P3_U3153) );
  XNOR2_X1 U14493 ( .A(n11886), .B(n12025), .ZN(n11887) );
  XNOR2_X1 U14494 ( .A(n11888), .B(n11887), .ZN(n11894) );
  INV_X1 U14495 ( .A(n11889), .ZN(n12648) );
  NOR2_X1 U14496 ( .A1(n12775), .A2(n12068), .ZN(n11892) );
  AND2_X1 U14497 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12335) );
  AOI21_X1 U14498 ( .B1(n12050), .B2(n12610), .A(n12335), .ZN(n11890) );
  OAI21_X1 U14499 ( .B1(n12052), .B2(n12643), .A(n11890), .ZN(n11891) );
  AOI211_X1 U14500 ( .C1(n12648), .C2(n12071), .A(n11892), .B(n11891), .ZN(
        n11893) );
  OAI21_X1 U14501 ( .B1(n11894), .B2(n12073), .A(n11893), .ZN(P3_U3155) );
  XNOR2_X1 U14502 ( .A(n11895), .B(n12508), .ZN(n11900) );
  AOI22_X1 U14503 ( .A1(n12521), .A2(n12050), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11897) );
  NAND2_X1 U14504 ( .A1(n12071), .A2(n12524), .ZN(n11896) );
  OAI211_X1 U14505 ( .C1(n11928), .C2(n12052), .A(n11897), .B(n11896), .ZN(
        n11898) );
  AOI21_X1 U14506 ( .B1(n12680), .B2(n12036), .A(n11898), .ZN(n11899) );
  OAI21_X1 U14507 ( .B1(n11900), .B2(n12073), .A(n11899), .ZN(P3_U3156) );
  OR2_X1 U14508 ( .A1(n11973), .A2(n11972), .ZN(n11974) );
  NAND2_X1 U14509 ( .A1(n11974), .A2(n11901), .ZN(n12044) );
  NAND2_X1 U14510 ( .A1(n12044), .A2(n12043), .ZN(n12042) );
  NAND2_X1 U14511 ( .A1(n12042), .A2(n11902), .ZN(n11905) );
  OAI211_X1 U14512 ( .C1(n11905), .C2(n11904), .A(n11903), .B(n12041), .ZN(
        n11909) );
  AND2_X1 U14513 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12443) );
  AOI21_X1 U14514 ( .B1(n12050), .B2(n12568), .A(n12443), .ZN(n11906) );
  OAI21_X1 U14515 ( .B1(n12052), .B2(n11976), .A(n11906), .ZN(n11907) );
  AOI21_X1 U14516 ( .B1(n12572), .B2(n12071), .A(n11907), .ZN(n11908) );
  OAI211_X1 U14517 ( .C1(n12068), .C2(n12756), .A(n11909), .B(n11908), .ZN(
        P3_U3159) );
  MUX2_X1 U14518 ( .A(n12283), .B(n11911), .S(n11910), .Z(n11913) );
  XNOR2_X1 U14519 ( .A(n11913), .B(n11912), .ZN(n11914) );
  NAND2_X1 U14520 ( .A1(n11914), .A2(n12041), .ZN(n11921) );
  AOI21_X1 U14521 ( .B1(n12036), .B2(n11916), .A(n11915), .ZN(n11920) );
  AOI22_X1 U14522 ( .A1(n12050), .A2(n12281), .B1(n12062), .B2(n12283), .ZN(
        n11919) );
  NAND2_X1 U14523 ( .A1(n12071), .A2(n11917), .ZN(n11918) );
  NAND4_X1 U14524 ( .A1(n11921), .A2(n11920), .A3(n11919), .A4(n11918), .ZN(
        P3_U3161) );
  INV_X1 U14525 ( .A(n11922), .ZN(n11923) );
  AOI21_X1 U14526 ( .B1(n11925), .B2(n11924), .A(n11923), .ZN(n11931) );
  AOI22_X1 U14527 ( .A1(n12062), .A2(n12568), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11927) );
  NAND2_X1 U14528 ( .A1(n12071), .A2(n12547), .ZN(n11926) );
  OAI211_X1 U14529 ( .C1(n11928), .C2(n12065), .A(n11927), .B(n11926), .ZN(
        n11929) );
  AOI21_X1 U14530 ( .B1(n12690), .B2(n12036), .A(n11929), .ZN(n11930) );
  OAI21_X1 U14531 ( .B1(n11931), .B2(n12073), .A(n11930), .ZN(P3_U3163) );
  INV_X1 U14532 ( .A(n11932), .ZN(n11937) );
  NOR3_X1 U14533 ( .A1(n11935), .A2(n11934), .A3(n11933), .ZN(n11936) );
  OAI21_X1 U14534 ( .B1(n11937), .B2(n11936), .A(n12041), .ZN(n11941) );
  AND2_X1 U14535 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n15086) );
  AOI21_X1 U14536 ( .B1(n12062), .B2(n12279), .A(n15086), .ZN(n11938) );
  OAI21_X1 U14537 ( .B1(n12643), .B2(n12065), .A(n11938), .ZN(n11939) );
  AOI21_X1 U14538 ( .B1(n12036), .B2(n14524), .A(n11939), .ZN(n11940) );
  OAI211_X1 U14539 ( .C1(n11942), .C2(n12028), .A(n11941), .B(n11940), .ZN(
        P3_U3164) );
  XOR2_X1 U14540 ( .A(n11944), .B(n11943), .Z(n11950) );
  AOI22_X1 U14541 ( .A1(n12274), .A2(n12050), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11945) );
  OAI21_X1 U14542 ( .B1(n11946), .B2(n12052), .A(n11945), .ZN(n11948) );
  NOR2_X1 U14543 ( .A1(n12739), .A2(n12068), .ZN(n11947) );
  AOI211_X1 U14544 ( .C1(n12501), .C2(n12071), .A(n11948), .B(n11947), .ZN(
        n11949) );
  OAI21_X1 U14545 ( .B1(n11950), .B2(n12073), .A(n11949), .ZN(P3_U3165) );
  XNOR2_X1 U14546 ( .A(n11951), .B(n12066), .ZN(n11952) );
  XNOR2_X1 U14547 ( .A(n11953), .B(n11952), .ZN(n11958) );
  NAND2_X1 U14548 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12366)
         );
  OAI21_X1 U14549 ( .B1(n12065), .B2(n12583), .A(n12366), .ZN(n11954) );
  AOI21_X1 U14550 ( .B1(n12062), .B2(n12610), .A(n11954), .ZN(n11955) );
  OAI21_X1 U14551 ( .B1(n12617), .B2(n12028), .A(n11955), .ZN(n11956) );
  AOI21_X1 U14552 ( .B1(n12036), .B2(n12616), .A(n11956), .ZN(n11957) );
  OAI21_X1 U14553 ( .B1(n11958), .B2(n12073), .A(n11957), .ZN(P3_U3166) );
  AOI21_X1 U14554 ( .B1(n11961), .B2(n11960), .A(n11959), .ZN(n11962) );
  OR2_X1 U14555 ( .A1(n11962), .A2(n12073), .ZN(n11970) );
  INV_X1 U14556 ( .A(n11963), .ZN(n11965) );
  AOI21_X1 U14557 ( .B1(n12036), .B2(n11965), .A(n11964), .ZN(n11969) );
  AOI22_X1 U14558 ( .A1(n12050), .A2(n12284), .B1(n12062), .B2(n15108), .ZN(
        n11968) );
  NAND2_X1 U14559 ( .A1(n12071), .A2(n11966), .ZN(n11967) );
  NAND4_X1 U14560 ( .A1(n11970), .A2(n11969), .A3(n11968), .A4(n11967), .ZN(
        P3_U3167) );
  INV_X1 U14561 ( .A(n11971), .ZN(n12763) );
  AOI21_X1 U14562 ( .B1(n11973), .B2(n11972), .A(n12073), .ZN(n11975) );
  NAND2_X1 U14563 ( .A1(n11975), .A2(n11974), .ZN(n11980) );
  NAND2_X1 U14564 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12390)
         );
  OAI21_X1 U14565 ( .B1(n12065), .B2(n11976), .A(n12390), .ZN(n11978) );
  NOR2_X1 U14566 ( .A1(n12028), .A2(n12601), .ZN(n11977) );
  AOI211_X1 U14567 ( .C1(n12062), .C2(n12626), .A(n11978), .B(n11977), .ZN(
        n11979) );
  OAI211_X1 U14568 ( .C1(n12763), .C2(n12068), .A(n11980), .B(n11979), .ZN(
        P3_U3168) );
  XOR2_X1 U14569 ( .A(n11982), .B(n11981), .Z(n11987) );
  INV_X1 U14570 ( .A(n12484), .ZN(n12507) );
  AOI22_X1 U14571 ( .A1(n12507), .A2(n12050), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11983) );
  OAI21_X1 U14572 ( .B1(n12533), .B2(n12052), .A(n11983), .ZN(n11985) );
  NOR2_X1 U14573 ( .A1(n12514), .A2(n12068), .ZN(n11984) );
  AOI211_X1 U14574 ( .C1(n12512), .C2(n12071), .A(n11985), .B(n11984), .ZN(
        n11986) );
  OAI21_X1 U14575 ( .B1(n11987), .B2(n12073), .A(n11986), .ZN(P3_U3169) );
  AOI21_X1 U14576 ( .B1(n11990), .B2(n11989), .A(n11988), .ZN(n11991) );
  OR2_X1 U14577 ( .A1(n11991), .A2(n12073), .ZN(n11998) );
  AOI21_X1 U14578 ( .B1(n12036), .B2(n15174), .A(n11992), .ZN(n11997) );
  AOI22_X1 U14579 ( .A1(n12050), .A2(n11993), .B1(n12062), .B2(n15123), .ZN(
        n11996) );
  NAND2_X1 U14580 ( .A1(n12071), .A2(n11994), .ZN(n11995) );
  NAND4_X1 U14581 ( .A1(n11998), .A2(n11997), .A3(n11996), .A4(n11995), .ZN(
        P3_U3170) );
  INV_X1 U14582 ( .A(n11999), .ZN(n12000) );
  AOI21_X1 U14583 ( .B1(n12002), .B2(n12001), .A(n12000), .ZN(n12003) );
  OR2_X1 U14584 ( .A1(n12003), .A2(n12073), .ZN(n12011) );
  AOI21_X1 U14585 ( .B1(n12036), .B2(n12005), .A(n12004), .ZN(n12010) );
  AOI22_X1 U14586 ( .A1(n12050), .A2(n12280), .B1(n12062), .B2(n12282), .ZN(
        n12009) );
  INV_X1 U14587 ( .A(n12006), .ZN(n12007) );
  NAND2_X1 U14588 ( .A1(n12071), .A2(n12007), .ZN(n12008) );
  NAND4_X1 U14589 ( .A1(n12011), .A2(n12010), .A3(n12009), .A4(n12008), .ZN(
        P3_U3171) );
  OAI211_X1 U14590 ( .C1(n12014), .C2(n12013), .A(n12012), .B(n12041), .ZN(
        n12018) );
  AOI22_X1 U14591 ( .A1(n12050), .A2(n12276), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12015) );
  OAI21_X1 U14592 ( .B1(n12584), .B2(n12052), .A(n12015), .ZN(n12016) );
  AOI21_X1 U14593 ( .B1(n12562), .B2(n12071), .A(n12016), .ZN(n12017) );
  OAI211_X1 U14594 ( .C1(n12753), .C2(n12068), .A(n12018), .B(n12017), .ZN(
        P3_U3173) );
  INV_X1 U14595 ( .A(n12019), .ZN(n12021) );
  NAND2_X1 U14596 ( .A1(n12021), .A2(n12020), .ZN(n12022) );
  XNOR2_X1 U14597 ( .A(n12023), .B(n12022), .ZN(n12031) );
  NOR2_X1 U14598 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12024), .ZN(n12314) );
  NOR2_X1 U14599 ( .A1(n12065), .A2(n12025), .ZN(n12026) );
  AOI211_X1 U14600 ( .C1(n12062), .C2(n14508), .A(n12314), .B(n12026), .ZN(
        n12027) );
  OAI21_X1 U14601 ( .B1(n14513), .B2(n12028), .A(n12027), .ZN(n12029) );
  AOI21_X1 U14602 ( .B1(n12036), .B2(n14512), .A(n12029), .ZN(n12030) );
  OAI21_X1 U14603 ( .B1(n12031), .B2(n12073), .A(n12030), .ZN(P3_U3174) );
  XNOR2_X1 U14604 ( .A(n12032), .B(n12543), .ZN(n12039) );
  AOI22_X1 U14605 ( .A1(n12062), .A2(n12276), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12034) );
  NAND2_X1 U14606 ( .A1(n12071), .A2(n12536), .ZN(n12033) );
  OAI211_X1 U14607 ( .C1(n12533), .C2(n12065), .A(n12034), .B(n12033), .ZN(
        n12035) );
  AOI21_X1 U14608 ( .B1(n12037), .B2(n12036), .A(n12035), .ZN(n12038) );
  OAI21_X1 U14609 ( .B1(n12039), .B2(n12073), .A(n12038), .ZN(P3_U3175) );
  INV_X1 U14610 ( .A(n12040), .ZN(n12759) );
  OAI211_X1 U14611 ( .C1(n12044), .C2(n12043), .A(n12042), .B(n12041), .ZN(
        n12048) );
  NAND2_X1 U14612 ( .A1(n12062), .A2(n12611), .ZN(n12045) );
  NAND2_X1 U14613 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12414)
         );
  OAI211_X1 U14614 ( .C1(n12584), .C2(n12065), .A(n12045), .B(n12414), .ZN(
        n12046) );
  AOI21_X1 U14615 ( .B1(n12588), .B2(n12071), .A(n12046), .ZN(n12047) );
  OAI211_X1 U14616 ( .C1(n12759), .C2(n12068), .A(n12048), .B(n12047), .ZN(
        P3_U3178) );
  AOI22_X1 U14617 ( .A1(n7249), .A2(n12050), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12051) );
  OAI21_X1 U14618 ( .B1(n12484), .B2(n12052), .A(n12051), .ZN(n12054) );
  NOR2_X1 U14619 ( .A1(n12735), .A2(n12068), .ZN(n12053) );
  AOI211_X1 U14620 ( .C1(n12487), .C2(n12071), .A(n12054), .B(n12053), .ZN(
        n12055) );
  OAI21_X1 U14621 ( .B1(n12056), .B2(n12073), .A(n12055), .ZN(P3_U3180) );
  INV_X1 U14622 ( .A(n12057), .ZN(n12058) );
  AOI21_X1 U14623 ( .B1(n12060), .B2(n12059), .A(n12058), .ZN(n12074) );
  INV_X1 U14624 ( .A(n12061), .ZN(n12632) );
  NAND2_X1 U14625 ( .A1(n12062), .A2(n14507), .ZN(n12064) );
  NOR2_X1 U14626 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15254), .ZN(n14495) );
  INV_X1 U14627 ( .A(n14495), .ZN(n12063) );
  OAI211_X1 U14628 ( .C1(n12066), .C2(n12065), .A(n12064), .B(n12063), .ZN(
        n12070) );
  INV_X1 U14629 ( .A(n12067), .ZN(n12771) );
  NOR2_X1 U14630 ( .A1(n12771), .A2(n12068), .ZN(n12069) );
  AOI211_X1 U14631 ( .C1(n12632), .C2(n12071), .A(n12070), .B(n12069), .ZN(
        n12072) );
  OAI21_X1 U14632 ( .B1(n12074), .B2(n12073), .A(n12072), .ZN(P3_U3181) );
  NAND2_X1 U14633 ( .A1(n12075), .A2(n6443), .ZN(n12077) );
  NAND2_X1 U14634 ( .A1(n8664), .A2(SI_30_), .ZN(n12076) );
  NAND2_X1 U14635 ( .A1(n12077), .A2(n12076), .ZN(n14518) );
  NAND2_X1 U14636 ( .A1(n12080), .A2(n12079), .ZN(n12082) );
  NAND2_X1 U14637 ( .A1(n8664), .A2(SI_31_), .ZN(n12081) );
  INV_X1 U14638 ( .A(n12083), .ZN(n12084) );
  AOI21_X1 U14639 ( .B1(n12086), .B2(n14518), .A(n12084), .ZN(n12085) );
  NAND2_X1 U14640 ( .A1(n12724), .A2(n12450), .ZN(n12088) );
  OR2_X1 U14641 ( .A1(n14518), .A2(n12086), .ZN(n12087) );
  NAND2_X1 U14642 ( .A1(n12088), .A2(n12087), .ZN(n12262) );
  NAND2_X1 U14643 ( .A1(n12245), .A2(n12246), .ZN(n12486) );
  NOR2_X1 U14644 ( .A1(n12510), .A2(n12090), .ZN(n12117) );
  INV_X1 U14645 ( .A(n12545), .ZN(n12227) );
  NAND2_X1 U14646 ( .A1(n12233), .A2(n12234), .ZN(n12534) );
  INV_X1 U14647 ( .A(n12091), .ZN(n12167) );
  NAND4_X1 U14648 ( .A1(n12093), .A2(n12092), .A3(n10197), .A4(n12167), .ZN(
        n12098) );
  NAND4_X1 U14649 ( .A1(n12156), .A2(n12095), .A3(n12162), .A4(n12094), .ZN(
        n12097) );
  NOR3_X1 U14650 ( .A1(n12098), .A2(n12097), .A3(n12096), .ZN(n12100) );
  NAND4_X1 U14651 ( .A1(n12100), .A2(n12141), .A3(n7210), .A4(n12099), .ZN(
        n12101) );
  NOR4_X1 U14652 ( .A1(n12182), .A2(n12640), .A3(n12101), .A4(n14505), .ZN(
        n12102) );
  NAND4_X1 U14653 ( .A1(n12599), .A2(n12102), .A3(n12630), .A4(n12614), .ZN(
        n12103) );
  NOR4_X1 U14654 ( .A1(n12534), .A2(n8907), .A3(n6465), .A4(n12103), .ZN(
        n12104) );
  INV_X1 U14655 ( .A(n12552), .ZN(n12560) );
  NAND4_X1 U14656 ( .A1(n12117), .A2(n12227), .A3(n12104), .A4(n12560), .ZN(
        n12105) );
  NOR3_X1 U14657 ( .A1(n12486), .A2(n12105), .A3(n12493), .ZN(n12106) );
  NAND4_X1 U14658 ( .A1(n12461), .A2(n12106), .A3(n12258), .A4(n12248), .ZN(
        n12107) );
  INV_X1 U14659 ( .A(n12486), .ZN(n12243) );
  NAND2_X1 U14660 ( .A1(n12111), .A2(n12110), .ZN(n12112) );
  AND2_X1 U14661 ( .A1(n12112), .A2(n12113), .ZN(n12116) );
  OAI21_X1 U14662 ( .B1(n12510), .B2(n12114), .A(n12113), .ZN(n12115) );
  MUX2_X1 U14663 ( .A(n12116), .B(n12115), .S(n12260), .Z(n12239) );
  INV_X1 U14664 ( .A(n12117), .ZN(n12238) );
  MUX2_X1 U14665 ( .A(n12122), .B(n12118), .S(n12244), .Z(n12129) );
  INV_X1 U14666 ( .A(n12119), .ZN(n12120) );
  INV_X1 U14667 ( .A(n14437), .ZN(n12271) );
  NAND2_X1 U14668 ( .A1(n12120), .A2(n12271), .ZN(n12124) );
  NAND2_X1 U14669 ( .A1(n12120), .A2(n12127), .ZN(n12121) );
  NAND3_X1 U14670 ( .A1(n12122), .A2(n12121), .A3(n12244), .ZN(n12123) );
  OAI21_X1 U14671 ( .B1(n15148), .B2(n12124), .A(n12123), .ZN(n12125) );
  OAI21_X1 U14672 ( .B1(n12127), .B2(n12126), .A(n12125), .ZN(n12128) );
  NAND3_X1 U14673 ( .A1(n12129), .A2(n7210), .A3(n12128), .ZN(n12136) );
  NAND2_X1 U14674 ( .A1(n12138), .A2(n12130), .ZN(n12133) );
  NAND2_X1 U14675 ( .A1(n15144), .A2(n15131), .ZN(n12131) );
  NAND2_X1 U14676 ( .A1(n12137), .A2(n12131), .ZN(n12132) );
  MUX2_X1 U14677 ( .A(n12133), .B(n12132), .S(n12260), .Z(n12134) );
  INV_X1 U14678 ( .A(n12134), .ZN(n12135) );
  NAND2_X1 U14679 ( .A1(n12136), .A2(n12135), .ZN(n12140) );
  MUX2_X1 U14680 ( .A(n12138), .B(n12137), .S(n12244), .Z(n12139) );
  NAND2_X1 U14681 ( .A1(n12140), .A2(n12139), .ZN(n12142) );
  NAND2_X1 U14682 ( .A1(n12142), .A2(n12141), .ZN(n12148) );
  NAND2_X1 U14683 ( .A1(n15108), .A2(n12143), .ZN(n12144) );
  MUX2_X1 U14684 ( .A(n12145), .B(n12144), .S(n12244), .Z(n12147) );
  AOI21_X1 U14685 ( .B1(n12148), .B2(n12147), .A(n12146), .ZN(n12158) );
  NAND2_X1 U14686 ( .A1(n12154), .A2(n12149), .ZN(n12152) );
  NAND2_X1 U14687 ( .A1(n12153), .A2(n12150), .ZN(n12151) );
  MUX2_X1 U14688 ( .A(n12152), .B(n12151), .S(n12244), .Z(n12157) );
  MUX2_X1 U14689 ( .A(n12154), .B(n12153), .S(n12260), .Z(n12155) );
  OAI211_X1 U14690 ( .C1(n12158), .C2(n12157), .A(n12156), .B(n12155), .ZN(
        n12163) );
  MUX2_X1 U14691 ( .A(n12160), .B(n12159), .S(n12260), .Z(n12161) );
  NAND3_X1 U14692 ( .A1(n12163), .A2(n12162), .A3(n12161), .ZN(n12168) );
  MUX2_X1 U14693 ( .A(n12165), .B(n12164), .S(n12260), .Z(n12166) );
  NAND3_X1 U14694 ( .A1(n12168), .A2(n12167), .A3(n12166), .ZN(n12172) );
  MUX2_X1 U14695 ( .A(n12170), .B(n12169), .S(n12260), .Z(n12171) );
  NAND4_X1 U14696 ( .A1(n12172), .A2(n7225), .A3(n7566), .A4(n12171), .ZN(
        n12177) );
  OAI211_X1 U14697 ( .C1(n12182), .C2(n12174), .A(n12184), .B(n12173), .ZN(
        n12175) );
  NAND2_X1 U14698 ( .A1(n12175), .A2(n12244), .ZN(n12176) );
  NAND2_X1 U14699 ( .A1(n12177), .A2(n12176), .ZN(n12178) );
  NAND2_X1 U14700 ( .A1(n12178), .A2(n12180), .ZN(n12187) );
  NAND2_X1 U14701 ( .A1(n14529), .A2(n12279), .ZN(n12179) );
  OAI211_X1 U14702 ( .C1(n12182), .C2(n12181), .A(n12180), .B(n12179), .ZN(
        n12183) );
  NAND2_X1 U14703 ( .A1(n12183), .A2(n12260), .ZN(n12186) );
  NOR2_X1 U14704 ( .A1(n12184), .A2(n12244), .ZN(n12185) );
  AOI21_X1 U14705 ( .B1(n12187), .B2(n12186), .A(n12185), .ZN(n12191) );
  MUX2_X1 U14706 ( .A(n12189), .B(n12188), .S(n12244), .Z(n12190) );
  OAI211_X1 U14707 ( .C1(n12191), .C2(n14505), .A(n7221), .B(n12190), .ZN(
        n12195) );
  MUX2_X1 U14708 ( .A(n12193), .B(n12192), .S(n12244), .Z(n12194) );
  NAND3_X1 U14709 ( .A1(n12195), .A2(n12630), .A3(n12194), .ZN(n12199) );
  NAND2_X1 U14710 ( .A1(n12202), .A2(n12196), .ZN(n12197) );
  NAND2_X1 U14711 ( .A1(n12197), .A2(n12244), .ZN(n12198) );
  AOI21_X1 U14712 ( .B1(n12199), .B2(n12198), .A(n7001), .ZN(n12204) );
  AOI21_X1 U14713 ( .B1(n12201), .B2(n12200), .A(n12244), .ZN(n12203) );
  OAI22_X1 U14714 ( .A1(n12204), .A2(n12203), .B1(n12244), .B2(n12202), .ZN(
        n12205) );
  NAND3_X1 U14715 ( .A1(n12205), .A2(n12599), .A3(n12580), .ZN(n12217) );
  INV_X1 U14716 ( .A(n12211), .ZN(n12208) );
  OAI211_X1 U14717 ( .C1(n12208), .C2(n12207), .A(n12219), .B(n12206), .ZN(
        n12214) );
  INV_X1 U14718 ( .A(n12209), .ZN(n12210) );
  NAND2_X1 U14719 ( .A1(n12580), .A2(n12210), .ZN(n12212) );
  NAND3_X1 U14720 ( .A1(n12212), .A2(n12218), .A3(n12211), .ZN(n12213) );
  MUX2_X1 U14721 ( .A(n12214), .B(n12213), .S(n12244), .Z(n12215) );
  INV_X1 U14722 ( .A(n12215), .ZN(n12216) );
  NAND2_X1 U14723 ( .A1(n12217), .A2(n12216), .ZN(n12221) );
  MUX2_X1 U14724 ( .A(n12219), .B(n12218), .S(n12260), .Z(n12220) );
  NAND3_X1 U14725 ( .A1(n12221), .A2(n12560), .A3(n12220), .ZN(n12228) );
  NAND2_X1 U14726 ( .A1(n12223), .A2(n12222), .ZN(n12225) );
  MUX2_X1 U14727 ( .A(n12225), .B(n12224), .S(n12260), .Z(n12226) );
  NAND3_X1 U14728 ( .A1(n12228), .A2(n12227), .A3(n12226), .ZN(n12232) );
  INV_X1 U14729 ( .A(n12534), .ZN(n12530) );
  MUX2_X1 U14730 ( .A(n12230), .B(n12229), .S(n12244), .Z(n12231) );
  NAND3_X1 U14731 ( .A1(n12232), .A2(n12530), .A3(n12231), .ZN(n12236) );
  MUX2_X1 U14732 ( .A(n12234), .B(n12233), .S(n12260), .Z(n12235) );
  NAND2_X1 U14733 ( .A1(n12236), .A2(n12235), .ZN(n12237) );
  MUX2_X1 U14734 ( .A(n12507), .B(n12244), .S(n12240), .Z(n12241) );
  OAI21_X1 U14735 ( .B1(n12484), .B2(n12260), .A(n12241), .ZN(n12242) );
  OR3_X1 U14736 ( .A1(n12477), .A2(n12483), .A3(n12260), .ZN(n12249) );
  NAND2_X1 U14737 ( .A1(n12250), .A2(n12249), .ZN(n12251) );
  INV_X1 U14738 ( .A(n12252), .ZN(n12253) );
  NAND3_X1 U14739 ( .A1(n12254), .A2(n12260), .A3(n12253), .ZN(n12256) );
  NAND2_X1 U14740 ( .A1(n12256), .A2(n12255), .ZN(n12257) );
  OAI211_X1 U14741 ( .C1(n12261), .C2(n12260), .A(n12259), .B(n12258), .ZN(
        n12264) );
  AOI22_X1 U14742 ( .A1(n12265), .A2(n12264), .B1(n12263), .B2(n12262), .ZN(
        n12266) );
  NAND3_X1 U14743 ( .A1(n12269), .A2(n12268), .A3(n6446), .ZN(n12270) );
  OAI211_X1 U14744 ( .C1(n12271), .C2(n12273), .A(n12270), .B(P3_B_REG_SCAN_IN), .ZN(n12272) );
  MUX2_X1 U14745 ( .A(n7249), .B(P3_DATAO_REG_27__SCAN_IN), .S(n12275), .Z(
        P3_U3518) );
  MUX2_X1 U14746 ( .A(n12274), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12275), .Z(
        P3_U3517) );
  MUX2_X1 U14747 ( .A(n12507), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12275), .Z(
        P3_U3516) );
  MUX2_X1 U14748 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12521), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14749 ( .A(n12508), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12275), .Z(
        P3_U3514) );
  MUX2_X1 U14750 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12543), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14751 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12276), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14752 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12568), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14753 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12277), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14754 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12596), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14755 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12611), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14756 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12626), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14757 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12610), .S(n12285), .Z(
        P3_U3506) );
  MUX2_X1 U14758 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n14507), .S(n12285), .Z(
        P3_U3505) );
  MUX2_X1 U14759 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12278), .S(n12285), .Z(
        P3_U3504) );
  MUX2_X1 U14760 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n14508), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14761 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12279), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14762 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12280), .S(n12285), .Z(
        P3_U3501) );
  MUX2_X1 U14763 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12281), .S(n12285), .Z(
        P3_U3500) );
  MUX2_X1 U14764 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12282), .S(n12285), .Z(
        P3_U3499) );
  MUX2_X1 U14765 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12283), .S(n12285), .Z(
        P3_U3498) );
  MUX2_X1 U14766 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12284), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14767 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n15108), .S(n12285), .Z(
        P3_U3495) );
  MUX2_X1 U14768 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n15144), .S(n12285), .Z(
        P3_U3493) );
  MUX2_X1 U14769 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n15124), .S(n12285), .Z(
        P3_U3492) );
  OAI22_X1 U14770 ( .A1(n15097), .A2(n12287), .B1(n15074), .B2(n12286), .ZN(
        n12288) );
  AOI21_X1 U14771 ( .B1(P3_REG2_REG_0__SCAN_IN), .B2(n15089), .A(n12288), .ZN(
        n12290) );
  MUX2_X1 U14772 ( .A(n15068), .B(n12290), .S(n12289), .Z(n12297) );
  AOI22_X1 U14773 ( .A1(n15087), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n12296) );
  NAND2_X1 U14774 ( .A1(n15097), .A2(n15074), .ZN(n12294) );
  INV_X1 U14775 ( .A(n12292), .ZN(n12293) );
  OAI21_X1 U14776 ( .B1(n15089), .B2(n12294), .A(n12293), .ZN(n12295) );
  NAND3_X1 U14777 ( .A1(n12297), .A2(n12296), .A3(n12295), .ZN(P3_U3182) );
  NOR2_X1 U14778 ( .A1(n7166), .A2(n12298), .ZN(n12300) );
  INV_X1 U14779 ( .A(n15083), .ZN(n12320) );
  NAND2_X1 U14780 ( .A1(n12320), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12303) );
  NAND2_X1 U14781 ( .A1(n15083), .A2(n12301), .ZN(n12302) );
  NAND2_X1 U14782 ( .A1(n12303), .A2(n12302), .ZN(n15090) );
  AOI21_X1 U14783 ( .B1(n12306), .B2(n12304), .A(n12333), .ZN(n12327) );
  MUX2_X1 U14784 ( .A(n12306), .B(n12305), .S(n6446), .Z(n12337) );
  XNOR2_X1 U14785 ( .A(n12337), .B(n12336), .ZN(n12313) );
  INV_X1 U14786 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14528) );
  MUX2_X1 U14787 ( .A(n12301), .B(n14528), .S(n6446), .Z(n12310) );
  OR2_X1 U14788 ( .A1(n15083), .A2(n12310), .ZN(n12311) );
  INV_X1 U14789 ( .A(n12307), .ZN(n12309) );
  XNOR2_X1 U14790 ( .A(n12310), .B(n12320), .ZN(n15102) );
  NAND2_X1 U14791 ( .A1(n12311), .A2(n15099), .ZN(n12312) );
  AOI21_X1 U14792 ( .B1(n12313), .B2(n12312), .A(n12340), .ZN(n12316) );
  AOI21_X1 U14793 ( .B1(n15087), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12314), 
        .ZN(n12315) );
  OAI21_X1 U14794 ( .B1(n12316), .B2(n15074), .A(n12315), .ZN(n12325) );
  NOR2_X1 U14795 ( .A1(n7166), .A2(n12317), .ZN(n12319) );
  XNOR2_X1 U14796 ( .A(n15083), .B(n14528), .ZN(n15096) );
  NAND2_X1 U14797 ( .A1(n12320), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12321) );
  AOI21_X1 U14798 ( .B1(n12305), .B2(n12322), .A(n12329), .ZN(n12323) );
  NOR2_X1 U14799 ( .A1(n12323), .A2(n15097), .ZN(n12324) );
  AOI211_X1 U14800 ( .C1(n15084), .C2(n12336), .A(n12325), .B(n12324), .ZN(
        n12326) );
  OAI21_X1 U14801 ( .B1(n12327), .B2(n15081), .A(n12326), .ZN(P3_U3195) );
  NOR2_X1 U14802 ( .A1(n12336), .A2(n12328), .ZN(n12330) );
  NAND2_X1 U14803 ( .A1(n12344), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12357) );
  OAI21_X1 U14804 ( .B1(n12344), .B2(P3_REG1_REG_14__SCAN_IN), .A(n12357), 
        .ZN(n12338) );
  INV_X1 U14805 ( .A(n12350), .ZN(n12331) );
  AOI21_X1 U14806 ( .B1(n6594), .B2(n12338), .A(n12331), .ZN(n12349) );
  NOR2_X1 U14807 ( .A1(n12336), .A2(n12332), .ZN(n12334) );
  NAND2_X1 U14808 ( .A1(n12344), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12369) );
  OAI21_X1 U14809 ( .B1(n12344), .B2(P3_REG2_REG_14__SCAN_IN), .A(n12369), 
        .ZN(n12368) );
  XNOR2_X1 U14810 ( .A(n6591), .B(n12368), .ZN(n12347) );
  INV_X1 U14811 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14324) );
  INV_X1 U14812 ( .A(n12335), .ZN(n12343) );
  MUX2_X1 U14813 ( .A(n12368), .B(n12338), .S(n6446), .Z(n12339) );
  OAI21_X1 U14814 ( .B1(n6607), .B2(n12340), .A(n12339), .ZN(n12341) );
  NAND3_X1 U14815 ( .A1(n15100), .A2(n6474), .A3(n12341), .ZN(n12342) );
  OAI211_X1 U14816 ( .C1(n15065), .C2(n14324), .A(n12343), .B(n12342), .ZN(
        n12346) );
  NOR2_X1 U14817 ( .A1(n15068), .A2(n12344), .ZN(n12345) );
  AOI211_X1 U14818 ( .C1(n15089), .C2(n12347), .A(n12346), .B(n12345), .ZN(
        n12348) );
  OAI21_X1 U14819 ( .B1(n12349), .B2(n15097), .A(n12348), .ZN(P3_U3196) );
  NOR2_X1 U14820 ( .A1(n12370), .A2(n12351), .ZN(n12352) );
  OR2_X1 U14821 ( .A1(n12373), .A2(n12713), .ZN(n12383) );
  NAND2_X1 U14822 ( .A1(n12373), .A2(n12713), .ZN(n12353) );
  NAND2_X1 U14823 ( .A1(n12383), .A2(n12353), .ZN(n12355) );
  INV_X1 U14824 ( .A(n12384), .ZN(n12354) );
  AOI21_X1 U14825 ( .B1(n12356), .B2(n12355), .A(n12354), .ZN(n12382) );
  MUX2_X1 U14826 ( .A(n12369), .B(n12357), .S(n6446), .Z(n12358) );
  NAND2_X1 U14827 ( .A1(n6474), .A2(n12358), .ZN(n12359) );
  AND2_X1 U14828 ( .A1(n12359), .A2(n14484), .ZN(n12360) );
  MUX2_X1 U14829 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n6446), .Z(n14490) );
  NOR2_X1 U14830 ( .A1(n14489), .A2(n14490), .ZN(n14488) );
  NOR2_X1 U14831 ( .A1(n12361), .A2(n14488), .ZN(n12394) );
  MUX2_X1 U14832 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n6446), .Z(n12364) );
  INV_X1 U14833 ( .A(n12364), .ZN(n12362) );
  NAND2_X1 U14834 ( .A1(n12362), .A2(n12373), .ZN(n12393) );
  INV_X1 U14835 ( .A(n12373), .ZN(n12363) );
  NAND2_X1 U14836 ( .A1(n12364), .A2(n12363), .ZN(n12392) );
  NAND2_X1 U14837 ( .A1(n12393), .A2(n12392), .ZN(n12365) );
  XNOR2_X1 U14838 ( .A(n12394), .B(n12365), .ZN(n12380) );
  INV_X1 U14839 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14323) );
  NAND2_X1 U14840 ( .A1(n15084), .A2(n12373), .ZN(n12367) );
  OAI211_X1 U14841 ( .C1(n14323), .C2(n15065), .A(n12367), .B(n12366), .ZN(
        n12379) );
  NOR2_X1 U14842 ( .A1(n12370), .A2(n12371), .ZN(n12372) );
  OR2_X1 U14843 ( .A1(n12373), .A2(n12618), .ZN(n12386) );
  NAND2_X1 U14844 ( .A1(n12373), .A2(n12618), .ZN(n12374) );
  NAND2_X1 U14845 ( .A1(n12386), .A2(n12374), .ZN(n12375) );
  NAND2_X1 U14846 ( .A1(n12376), .A2(n12375), .ZN(n12377) );
  AOI21_X1 U14847 ( .B1(n12387), .B2(n12377), .A(n15081), .ZN(n12378) );
  AOI211_X1 U14848 ( .C1(n15100), .C2(n12380), .A(n12379), .B(n12378), .ZN(
        n12381) );
  OAI21_X1 U14849 ( .B1(n12382), .B2(n15097), .A(n12381), .ZN(P3_U3198) );
  AOI21_X1 U14850 ( .B1(n12709), .B2(n12385), .A(n12402), .ZN(n12401) );
  AOI21_X1 U14851 ( .B1(n12602), .B2(n12388), .A(n12418), .ZN(n12391) );
  NAND2_X1 U14852 ( .A1(n15087), .A2(P3_ADDR_REG_17__SCAN_IN), .ZN(n12389) );
  OAI211_X1 U14853 ( .C1(n15081), .C2(n12391), .A(n12390), .B(n12389), .ZN(
        n12399) );
  INV_X1 U14854 ( .A(n12392), .ZN(n12395) );
  MUX2_X1 U14855 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n6446), .Z(n12407) );
  XNOR2_X1 U14856 ( .A(n12407), .B(n12406), .ZN(n12396) );
  AOI211_X1 U14857 ( .C1(n12397), .C2(n12396), .A(n12408), .B(n15074), .ZN(
        n12398) );
  AOI211_X1 U14858 ( .C1(n15084), .C2(n12417), .A(n12399), .B(n12398), .ZN(
        n12400) );
  OAI21_X1 U14859 ( .B1(n12401), .B2(n15097), .A(n12400), .ZN(P3_U3199) );
  NOR2_X1 U14860 ( .A1(n12417), .A2(n6558), .ZN(n12403) );
  NAND2_X1 U14861 ( .A1(n12419), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12425) );
  OAI21_X1 U14862 ( .B1(n12419), .B2(P3_REG1_REG_18__SCAN_IN), .A(n12425), 
        .ZN(n12404) );
  NOR2_X1 U14863 ( .A1(n12405), .A2(n12404), .ZN(n12427) );
  AOI21_X1 U14864 ( .B1(n12405), .B2(n12404), .A(n12427), .ZN(n12424) );
  NAND2_X1 U14865 ( .A1(n12407), .A2(n12406), .ZN(n12410) );
  INV_X1 U14866 ( .A(n12408), .ZN(n12409) );
  NAND2_X1 U14867 ( .A1(n12410), .A2(n12409), .ZN(n12431) );
  MUX2_X1 U14868 ( .A(n12411), .B(n12705), .S(n6446), .Z(n12412) );
  NAND2_X1 U14869 ( .A1(n12413), .A2(n12412), .ZN(n12435) );
  OAI21_X1 U14870 ( .B1(n12413), .B2(n12412), .A(n12435), .ZN(n12423) );
  INV_X1 U14871 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n15272) );
  NAND2_X1 U14872 ( .A1(n15084), .A2(n12432), .ZN(n12415) );
  OAI211_X1 U14873 ( .C1(n15272), .C2(n15065), .A(n12415), .B(n12414), .ZN(
        n12422) );
  NAND2_X1 U14874 ( .A1(n12419), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12429) );
  OAI21_X1 U14875 ( .B1(n12419), .B2(P3_REG2_REG_18__SCAN_IN), .A(n12429), 
        .ZN(n12420) );
  XNOR2_X1 U14876 ( .A(n12428), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12438) );
  INV_X1 U14877 ( .A(n12425), .ZN(n12426) );
  MUX2_X1 U14878 ( .A(P3_REG2_REG_19__SCAN_IN), .B(n8920), .S(n12428), .Z(
        n12436) );
  INV_X1 U14879 ( .A(n12431), .ZN(n12433) );
  NAND2_X1 U14880 ( .A1(n12433), .A2(n12432), .ZN(n12434) );
  NAND2_X1 U14881 ( .A1(n12435), .A2(n12434), .ZN(n12441) );
  INV_X1 U14882 ( .A(n12436), .ZN(n12439) );
  MUX2_X1 U14883 ( .A(n12439), .B(n12438), .S(n6446), .Z(n12440) );
  AOI21_X1 U14884 ( .B1(n15087), .B2(P3_ADDR_REG_19__SCAN_IN), .A(n12443), 
        .ZN(n12444) );
  AOI21_X1 U14885 ( .B1(n12446), .B2(n15089), .A(n12445), .ZN(n12447) );
  OAI21_X1 U14886 ( .B1(n12448), .B2(n15097), .A(n12447), .ZN(P3_U3201) );
  NAND2_X1 U14887 ( .A1(n12724), .A2(n14499), .ZN(n12453) );
  INV_X1 U14888 ( .A(n12451), .ZN(n12452) );
  OAI21_X1 U14889 ( .B1(n14517), .B2(n12452), .A(n15159), .ZN(n14500) );
  OAI211_X1 U14890 ( .C1(n15159), .C2(n12454), .A(n12453), .B(n14500), .ZN(
        P3_U3202) );
  NAND2_X1 U14891 ( .A1(n7249), .A2(n15142), .ZN(n12459) );
  OAI21_X1 U14892 ( .B1(n7632), .B2(n12460), .A(n7637), .ZN(n12657) );
  XNOR2_X1 U14893 ( .A(n12462), .B(n12461), .ZN(n12658) );
  AOI22_X1 U14894 ( .A1(n12463), .A2(n15136), .B1(n14498), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12465) );
  NAND2_X1 U14895 ( .A1(n12659), .A2(n14499), .ZN(n12464) );
  OAI211_X1 U14896 ( .C1(n12658), .C2(n12653), .A(n12465), .B(n12464), .ZN(
        n12466) );
  AOI21_X1 U14897 ( .B1(n12657), .B2(n15159), .A(n12466), .ZN(n12467) );
  INV_X1 U14898 ( .A(n12467), .ZN(P3_U3205) );
  XNOR2_X1 U14899 ( .A(n12468), .B(n12471), .ZN(n12664) );
  OAI21_X1 U14900 ( .B1(n12471), .B2(n12470), .A(n12469), .ZN(n12474) );
  OAI22_X1 U14901 ( .A1(n12472), .A2(n12646), .B1(n12497), .B2(n12642), .ZN(
        n12473) );
  AOI21_X1 U14902 ( .B1(n12474), .B2(n15149), .A(n12473), .ZN(n12475) );
  AOI22_X1 U14903 ( .A1(n12476), .A2(n15136), .B1(n14498), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12479) );
  NAND2_X1 U14904 ( .A1(n12477), .A2(n14499), .ZN(n12478) );
  OAI211_X1 U14905 ( .C1(n12664), .C2(n15156), .A(n12479), .B(n12478), .ZN(
        n12480) );
  AOI21_X1 U14906 ( .B1(n12665), .B2(n15159), .A(n12480), .ZN(n12481) );
  INV_X1 U14907 ( .A(n12481), .ZN(P3_U3206) );
  INV_X1 U14908 ( .A(n12668), .ZN(n12491) );
  XOR2_X1 U14909 ( .A(n12486), .B(n12485), .Z(n12669) );
  AOI22_X1 U14910 ( .A1(n12487), .A2(n15136), .B1(n14498), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12488) );
  OAI21_X1 U14911 ( .B1(n12735), .B2(n12650), .A(n12488), .ZN(n12489) );
  AOI21_X1 U14912 ( .B1(n12669), .B2(n12635), .A(n12489), .ZN(n12490) );
  OAI21_X1 U14913 ( .B1(n12491), .B2(n14498), .A(n12490), .ZN(P3_U3207) );
  OAI211_X1 U14914 ( .C1(n12494), .C2(n12493), .A(n12492), .B(n15149), .ZN(
        n12496) );
  NAND2_X1 U14915 ( .A1(n12521), .A2(n15142), .ZN(n12495) );
  OAI211_X1 U14916 ( .C1(n12497), .C2(n12646), .A(n12496), .B(n12495), .ZN(
        n12672) );
  INV_X1 U14917 ( .A(n12672), .ZN(n12505) );
  OAI21_X1 U14918 ( .B1(n12500), .B2(n12499), .A(n12498), .ZN(n12673) );
  AOI22_X1 U14919 ( .A1(n14498), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n12501), 
        .B2(n15136), .ZN(n12502) );
  OAI21_X1 U14920 ( .B1(n12739), .B2(n12650), .A(n12502), .ZN(n12503) );
  AOI21_X1 U14921 ( .B1(n12673), .B2(n12635), .A(n12503), .ZN(n12504) );
  OAI21_X1 U14922 ( .B1(n12505), .B2(n14498), .A(n12504), .ZN(P3_U3208) );
  XNOR2_X1 U14923 ( .A(n12506), .B(n12510), .ZN(n12509) );
  AOI222_X1 U14924 ( .A1(n15149), .A2(n12509), .B1(n12508), .B2(n15142), .C1(
        n12507), .C2(n15145), .ZN(n12679) );
  XNOR2_X1 U14925 ( .A(n12511), .B(n12510), .ZN(n12677) );
  AOI22_X1 U14926 ( .A1(n14498), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15136), 
        .B2(n12512), .ZN(n12513) );
  OAI21_X1 U14927 ( .B1(n12514), .B2(n12650), .A(n12513), .ZN(n12515) );
  AOI21_X1 U14928 ( .B1(n12677), .B2(n12635), .A(n12515), .ZN(n12516) );
  OAI21_X1 U14929 ( .B1(n12679), .B2(n14498), .A(n12516), .ZN(P3_U3209) );
  XNOR2_X1 U14930 ( .A(n12517), .B(n12518), .ZN(n12681) );
  XNOR2_X1 U14931 ( .A(n12519), .B(n12518), .ZN(n12520) );
  NAND2_X1 U14932 ( .A1(n12520), .A2(n15149), .ZN(n12523) );
  AOI22_X1 U14933 ( .A1(n12521), .A2(n15145), .B1(n15142), .B2(n12543), .ZN(
        n12522) );
  OAI211_X1 U14934 ( .C1(n15153), .C2(n12681), .A(n12523), .B(n12522), .ZN(
        n12682) );
  NAND2_X1 U14935 ( .A1(n12682), .A2(n15159), .ZN(n12529) );
  INV_X1 U14936 ( .A(n12524), .ZN(n12525) );
  OAI22_X1 U14937 ( .A1(n15159), .A2(n12526), .B1(n12525), .B2(n15154), .ZN(
        n12527) );
  AOI21_X1 U14938 ( .B1(n12680), .B2(n14499), .A(n12527), .ZN(n12528) );
  OAI211_X1 U14939 ( .C1(n12681), .C2(n15156), .A(n12529), .B(n12528), .ZN(
        P3_U3210) );
  XNOR2_X1 U14940 ( .A(n12531), .B(n12530), .ZN(n12532) );
  OAI222_X1 U14941 ( .A1(n12646), .A2(n12533), .B1(n12642), .B2(n12556), .C1(
        n12582), .C2(n12532), .ZN(n12686) );
  INV_X1 U14942 ( .A(n12686), .ZN(n12540) );
  XNOR2_X1 U14943 ( .A(n12535), .B(n12534), .ZN(n12687) );
  AOI22_X1 U14944 ( .A1(n14498), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15136), 
        .B2(n12536), .ZN(n12537) );
  OAI21_X1 U14945 ( .B1(n12748), .B2(n12650), .A(n12537), .ZN(n12538) );
  AOI21_X1 U14946 ( .B1(n12687), .B2(n12635), .A(n12538), .ZN(n12539) );
  OAI21_X1 U14947 ( .B1(n12540), .B2(n14498), .A(n12539), .ZN(P3_U3211) );
  OAI21_X1 U14948 ( .B1(n12542), .B2(n12545), .A(n12541), .ZN(n12544) );
  AOI222_X1 U14949 ( .A1(n15149), .A2(n12544), .B1(n12543), .B2(n15145), .C1(
        n12568), .C2(n15142), .ZN(n12693) );
  XNOR2_X1 U14950 ( .A(n12546), .B(n12545), .ZN(n12691) );
  INV_X1 U14951 ( .A(n12690), .ZN(n12549) );
  AOI22_X1 U14952 ( .A1(n14498), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15136), 
        .B2(n12547), .ZN(n12548) );
  OAI21_X1 U14953 ( .B1(n12549), .B2(n12650), .A(n12548), .ZN(n12550) );
  AOI21_X1 U14954 ( .B1(n12691), .B2(n12635), .A(n12550), .ZN(n12551) );
  OAI21_X1 U14955 ( .B1(n12693), .B2(n14498), .A(n12551), .ZN(P3_U3212) );
  NOR2_X1 U14956 ( .A1(n12553), .A2(n12552), .ZN(n12554) );
  OAI22_X1 U14957 ( .A1(n12556), .A2(n12646), .B1(n12584), .B2(n12642), .ZN(
        n12557) );
  INV_X1 U14958 ( .A(n12557), .ZN(n12558) );
  NAND2_X1 U14959 ( .A1(n12559), .A2(n12558), .ZN(n12696) );
  INV_X1 U14960 ( .A(n12696), .ZN(n12566) );
  XNOR2_X1 U14961 ( .A(n12561), .B(n12560), .ZN(n12694) );
  AOI22_X1 U14962 ( .A1(n14498), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15136), 
        .B2(n12562), .ZN(n12563) );
  OAI21_X1 U14963 ( .B1(n12753), .B2(n12650), .A(n12563), .ZN(n12564) );
  AOI21_X1 U14964 ( .B1(n12694), .B2(n12635), .A(n12564), .ZN(n12565) );
  OAI21_X1 U14965 ( .B1(n12566), .B2(n14498), .A(n12565), .ZN(P3_U3213) );
  OAI211_X1 U14966 ( .C1(n6597), .C2(n6465), .A(n15149), .B(n12567), .ZN(
        n12570) );
  AOI22_X1 U14967 ( .A1(n12568), .A2(n15145), .B1(n15142), .B2(n12596), .ZN(
        n12569) );
  NAND2_X1 U14968 ( .A1(n12570), .A2(n12569), .ZN(n12699) );
  INV_X1 U14969 ( .A(n12699), .ZN(n12576) );
  XNOR2_X1 U14970 ( .A(n12571), .B(n6465), .ZN(n12700) );
  AOI22_X1 U14971 ( .A1(n14498), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15136), 
        .B2(n12572), .ZN(n12573) );
  OAI21_X1 U14972 ( .B1(n12756), .B2(n12650), .A(n12573), .ZN(n12574) );
  AOI21_X1 U14973 ( .B1(n12700), .B2(n12635), .A(n12574), .ZN(n12575) );
  OAI21_X1 U14974 ( .B1(n12576), .B2(n14498), .A(n12575), .ZN(P3_U3214) );
  INV_X1 U14975 ( .A(n12577), .ZN(n12578) );
  AOI21_X1 U14976 ( .B1(n12580), .B2(n12579), .A(n12578), .ZN(n12581) );
  OAI222_X1 U14977 ( .A1(n12646), .A2(n12584), .B1(n12642), .B2(n12583), .C1(
        n12582), .C2(n12581), .ZN(n12703) );
  INV_X1 U14978 ( .A(n12703), .ZN(n12592) );
  INV_X1 U14979 ( .A(n12585), .ZN(n12586) );
  AOI21_X1 U14980 ( .B1(n8907), .B2(n12587), .A(n12586), .ZN(n12704) );
  AOI22_X1 U14981 ( .A1(n14498), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15136), 
        .B2(n12588), .ZN(n12589) );
  OAI21_X1 U14982 ( .B1(n12759), .B2(n12650), .A(n12589), .ZN(n12590) );
  AOI21_X1 U14983 ( .B1(n12704), .B2(n12635), .A(n12590), .ZN(n12591) );
  OAI21_X1 U14984 ( .B1(n12592), .B2(n14498), .A(n12591), .ZN(P3_U3215) );
  OAI211_X1 U14985 ( .C1(n12595), .C2(n12594), .A(n12593), .B(n15149), .ZN(
        n12598) );
  AOI22_X1 U14986 ( .A1(n15142), .A2(n12626), .B1(n12596), .B2(n15145), .ZN(
        n12597) );
  NAND2_X1 U14987 ( .A1(n12598), .A2(n12597), .ZN(n12707) );
  INV_X1 U14988 ( .A(n12707), .ZN(n12606) );
  XNOR2_X1 U14989 ( .A(n12600), .B(n12599), .ZN(n12708) );
  NOR2_X1 U14990 ( .A1(n12763), .A2(n12650), .ZN(n12604) );
  OAI22_X1 U14991 ( .A1(n15159), .A2(n12602), .B1(n12601), .B2(n15154), .ZN(
        n12603) );
  AOI211_X1 U14992 ( .C1(n12708), .C2(n12635), .A(n12604), .B(n12603), .ZN(
        n12605) );
  OAI21_X1 U14993 ( .B1(n12606), .B2(n14498), .A(n12605), .ZN(P3_U3216) );
  OAI211_X1 U14994 ( .C1(n12609), .C2(n12608), .A(n12607), .B(n15149), .ZN(
        n12613) );
  AOI22_X1 U14995 ( .A1(n12611), .A2(n15145), .B1(n15142), .B2(n12610), .ZN(
        n12612) );
  NAND2_X1 U14996 ( .A1(n12613), .A2(n12612), .ZN(n12711) );
  INV_X1 U14997 ( .A(n12711), .ZN(n12622) );
  XNOR2_X1 U14998 ( .A(n12615), .B(n12614), .ZN(n12712) );
  INV_X1 U14999 ( .A(n12616), .ZN(n12767) );
  NOR2_X1 U15000 ( .A1(n12767), .A2(n12650), .ZN(n12620) );
  OAI22_X1 U15001 ( .A1(n15159), .A2(n12618), .B1(n12617), .B2(n15154), .ZN(
        n12619) );
  AOI211_X1 U15002 ( .C1(n12712), .C2(n12635), .A(n12620), .B(n12619), .ZN(
        n12621) );
  OAI21_X1 U15003 ( .B1(n12622), .B2(n14498), .A(n12621), .ZN(P3_U3217) );
  OAI211_X1 U15004 ( .C1(n12625), .C2(n12624), .A(n12623), .B(n15149), .ZN(
        n12628) );
  AOI22_X1 U15005 ( .A1(n12626), .A2(n15145), .B1(n15142), .B2(n14507), .ZN(
        n12627) );
  NAND2_X1 U15006 ( .A1(n12628), .A2(n12627), .ZN(n12715) );
  INV_X1 U15007 ( .A(n12715), .ZN(n12637) );
  OAI21_X1 U15008 ( .B1(n12631), .B2(n12630), .A(n12629), .ZN(n12716) );
  AOI22_X1 U15009 ( .A1(n14498), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15136), 
        .B2(n12632), .ZN(n12633) );
  OAI21_X1 U15010 ( .B1(n12650), .B2(n12771), .A(n12633), .ZN(n12634) );
  AOI21_X1 U15011 ( .B1(n12716), .B2(n12635), .A(n12634), .ZN(n12636) );
  OAI21_X1 U15012 ( .B1(n12637), .B2(n14498), .A(n12636), .ZN(P3_U3218) );
  XNOR2_X1 U15013 ( .A(n12638), .B(n12640), .ZN(n12719) );
  INV_X1 U15014 ( .A(n12719), .ZN(n12654) );
  OAI211_X1 U15015 ( .C1(n12641), .C2(n12640), .A(n12639), .B(n15149), .ZN(
        n12645) );
  OR2_X1 U15016 ( .A1(n12643), .A2(n12642), .ZN(n12644) );
  OAI211_X1 U15017 ( .C1(n12647), .C2(n12646), .A(n12645), .B(n12644), .ZN(
        n12718) );
  AOI22_X1 U15018 ( .A1(n14498), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15136), 
        .B2(n12648), .ZN(n12649) );
  OAI21_X1 U15019 ( .B1(n12650), .B2(n12775), .A(n12649), .ZN(n12651) );
  AOI21_X1 U15020 ( .B1(n12718), .B2(n15159), .A(n12651), .ZN(n12652) );
  OAI21_X1 U15021 ( .B1(n12654), .B2(n12653), .A(n12652), .ZN(P3_U3219) );
  NAND2_X1 U15022 ( .A1(n12724), .A2(n6842), .ZN(n12656) );
  NAND2_X1 U15023 ( .A1(n14517), .A2(n15222), .ZN(n12655) );
  OAI211_X1 U15024 ( .C1(n15222), .C2(n10857), .A(n12656), .B(n12655), .ZN(
        P3_U3490) );
  NAND2_X1 U15025 ( .A1(n12659), .A2(n15173), .ZN(n12660) );
  MUX2_X1 U15026 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n12728), .S(n15222), .Z(
        P3_U3487) );
  INV_X1 U15027 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12667) );
  INV_X1 U15028 ( .A(n12664), .ZN(n12666) );
  INV_X1 U15029 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12670) );
  AOI21_X1 U15030 ( .B1(n12669), .B2(n9066), .A(n12668), .ZN(n12732) );
  MUX2_X1 U15031 ( .A(n12670), .B(n12732), .S(n15222), .Z(n12671) );
  INV_X1 U15032 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12674) );
  AOI21_X1 U15033 ( .B1(n9066), .B2(n12673), .A(n12672), .ZN(n12736) );
  MUX2_X1 U15034 ( .A(n12674), .B(n12736), .S(n15222), .Z(n12675) );
  OAI21_X1 U15035 ( .B1(n12739), .B2(n12722), .A(n12675), .ZN(P3_U3484) );
  AOI22_X1 U15036 ( .A1(n12677), .A2(n9066), .B1(n15173), .B2(n12676), .ZN(
        n12678) );
  NAND2_X1 U15037 ( .A1(n12679), .A2(n12678), .ZN(n12740) );
  MUX2_X1 U15038 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n12740), .S(n15222), .Z(
        P3_U3483) );
  INV_X1 U15039 ( .A(n12680), .ZN(n12744) );
  INV_X1 U15040 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12684) );
  INV_X1 U15041 ( .A(n12681), .ZN(n12683) );
  AOI21_X1 U15042 ( .B1(n15203), .B2(n12683), .A(n12682), .ZN(n12741) );
  MUX2_X1 U15043 ( .A(n12684), .B(n12741), .S(n15222), .Z(n12685) );
  OAI21_X1 U15044 ( .B1(n12744), .B2(n12722), .A(n12685), .ZN(P3_U3482) );
  INV_X1 U15045 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12688) );
  AOI21_X1 U15046 ( .B1(n9066), .B2(n12687), .A(n12686), .ZN(n12745) );
  MUX2_X1 U15047 ( .A(n12688), .B(n12745), .S(n15222), .Z(n12689) );
  OAI21_X1 U15048 ( .B1(n12748), .B2(n12722), .A(n12689), .ZN(P3_U3481) );
  AOI22_X1 U15049 ( .A1(n12691), .A2(n9066), .B1(n15173), .B2(n12690), .ZN(
        n12692) );
  NAND2_X1 U15050 ( .A1(n12693), .A2(n12692), .ZN(n12749) );
  MUX2_X1 U15051 ( .A(P3_REG1_REG_21__SCAN_IN), .B(n12749), .S(n15222), .Z(
        P3_U3480) );
  INV_X1 U15052 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12697) );
  AND2_X1 U15053 ( .A1(n12694), .A2(n9066), .ZN(n12695) );
  NOR2_X1 U15054 ( .A1(n12696), .A2(n12695), .ZN(n12750) );
  MUX2_X1 U15055 ( .A(n12697), .B(n12750), .S(n15222), .Z(n12698) );
  OAI21_X1 U15056 ( .B1(n12753), .B2(n12722), .A(n12698), .ZN(P3_U3479) );
  INV_X1 U15057 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12701) );
  AOI21_X1 U15058 ( .B1(n9066), .B2(n12700), .A(n12699), .ZN(n12754) );
  MUX2_X1 U15059 ( .A(n12701), .B(n12754), .S(n15222), .Z(n12702) );
  OAI21_X1 U15060 ( .B1(n12722), .B2(n12756), .A(n12702), .ZN(P3_U3478) );
  AOI21_X1 U15061 ( .B1(n12704), .B2(n9066), .A(n12703), .ZN(n12757) );
  MUX2_X1 U15062 ( .A(n12705), .B(n12757), .S(n15222), .Z(n12706) );
  OAI21_X1 U15063 ( .B1(n12759), .B2(n12722), .A(n12706), .ZN(P3_U3477) );
  AOI21_X1 U15064 ( .B1(n12708), .B2(n9066), .A(n12707), .ZN(n12760) );
  MUX2_X1 U15065 ( .A(n12709), .B(n12760), .S(n15222), .Z(n12710) );
  OAI21_X1 U15066 ( .B1(n12763), .B2(n12722), .A(n12710), .ZN(P3_U3476) );
  AOI21_X1 U15067 ( .B1(n12712), .B2(n9066), .A(n12711), .ZN(n12764) );
  MUX2_X1 U15068 ( .A(n12713), .B(n12764), .S(n15222), .Z(n12714) );
  OAI21_X1 U15069 ( .B1(n12767), .B2(n12722), .A(n12714), .ZN(P3_U3475) );
  AOI21_X1 U15070 ( .B1(n9066), .B2(n12716), .A(n12715), .ZN(n12768) );
  MUX2_X1 U15071 ( .A(n14487), .B(n12768), .S(n15222), .Z(n12717) );
  OAI21_X1 U15072 ( .B1(n12771), .B2(n12722), .A(n12717), .ZN(P3_U3474) );
  INV_X1 U15073 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12720) );
  AOI21_X1 U15074 ( .B1(n9066), .B2(n12719), .A(n12718), .ZN(n12772) );
  MUX2_X1 U15075 ( .A(n12720), .B(n12772), .S(n15222), .Z(n12721) );
  OAI21_X1 U15076 ( .B1(n12722), .B2(n12775), .A(n12721), .ZN(P3_U3473) );
  INV_X1 U15077 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12727) );
  INV_X1 U15078 ( .A(n12776), .ZN(n12723) );
  NAND2_X1 U15079 ( .A1(n12724), .A2(n12723), .ZN(n12726) );
  NAND2_X1 U15080 ( .A1(n14517), .A2(n15206), .ZN(n12725) );
  OAI211_X1 U15081 ( .C1(n12727), .C2(n15206), .A(n12726), .B(n12725), .ZN(
        P3_U3458) );
  MUX2_X1 U15082 ( .A(P3_REG0_REG_28__SCAN_IN), .B(n12728), .S(n15206), .Z(
        P3_U3455) );
  INV_X1 U15083 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12730) );
  INV_X1 U15084 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12733) );
  MUX2_X1 U15085 ( .A(n12733), .B(n12732), .S(n15206), .Z(n12734) );
  INV_X1 U15086 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12737) );
  MUX2_X1 U15087 ( .A(n12737), .B(n12736), .S(n15206), .Z(n12738) );
  OAI21_X1 U15088 ( .B1(n12739), .B2(n12776), .A(n12738), .ZN(P3_U3452) );
  MUX2_X1 U15089 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n12740), .S(n15206), .Z(
        P3_U3451) );
  INV_X1 U15090 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12742) );
  MUX2_X1 U15091 ( .A(n12742), .B(n12741), .S(n15206), .Z(n12743) );
  OAI21_X1 U15092 ( .B1(n12744), .B2(n12776), .A(n12743), .ZN(P3_U3450) );
  INV_X1 U15093 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12746) );
  MUX2_X1 U15094 ( .A(n12746), .B(n12745), .S(n15206), .Z(n12747) );
  OAI21_X1 U15095 ( .B1(n12748), .B2(n12776), .A(n12747), .ZN(P3_U3449) );
  MUX2_X1 U15096 ( .A(P3_REG0_REG_21__SCAN_IN), .B(n12749), .S(n15206), .Z(
        P3_U3448) );
  INV_X1 U15097 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12751) );
  MUX2_X1 U15098 ( .A(n12751), .B(n12750), .S(n15206), .Z(n12752) );
  OAI21_X1 U15099 ( .B1(n12753), .B2(n12776), .A(n12752), .ZN(P3_U3447) );
  MUX2_X1 U15100 ( .A(n15280), .B(n12754), .S(n15206), .Z(n12755) );
  OAI21_X1 U15101 ( .B1(n12776), .B2(n12756), .A(n12755), .ZN(P3_U3446) );
  MUX2_X1 U15102 ( .A(n15282), .B(n12757), .S(n15206), .Z(n12758) );
  OAI21_X1 U15103 ( .B1(n12759), .B2(n12776), .A(n12758), .ZN(P3_U3444) );
  INV_X1 U15104 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12761) );
  MUX2_X1 U15105 ( .A(n12761), .B(n12760), .S(n15206), .Z(n12762) );
  OAI21_X1 U15106 ( .B1(n12763), .B2(n12776), .A(n12762), .ZN(P3_U3441) );
  INV_X1 U15107 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12765) );
  MUX2_X1 U15108 ( .A(n12765), .B(n12764), .S(n15206), .Z(n12766) );
  OAI21_X1 U15109 ( .B1(n12767), .B2(n12776), .A(n12766), .ZN(P3_U3438) );
  INV_X1 U15110 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12769) );
  MUX2_X1 U15111 ( .A(n12769), .B(n12768), .S(n15206), .Z(n12770) );
  OAI21_X1 U15112 ( .B1(n12771), .B2(n12776), .A(n12770), .ZN(P3_U3435) );
  MUX2_X1 U15113 ( .A(n12773), .B(n12772), .S(n15206), .Z(n12774) );
  OAI21_X1 U15114 ( .B1(n12776), .B2(n12775), .A(n12774), .ZN(P3_U3432) );
  INV_X1 U15115 ( .A(n12780), .ZN(n13019) );
  AOI22_X1 U15116 ( .A1(n13019), .A2(n12888), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12781) );
  OAI21_X1 U15117 ( .B1(n13043), .B2(n12896), .A(n12781), .ZN(n12782) );
  AOI21_X1 U15118 ( .B1(n12848), .B2(n13011), .A(n12782), .ZN(n12783) );
  NAND2_X1 U15119 ( .A1(n13087), .A2(n12893), .ZN(n12787) );
  NAND2_X1 U15120 ( .A1(n12784), .A2(n12871), .ZN(n12786) );
  MUX2_X1 U15121 ( .A(n12787), .B(n12786), .S(n12785), .Z(n12791) );
  AOI22_X1 U15122 ( .A1(n13078), .A2(n12888), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12790) );
  AOI22_X1 U15123 ( .A1(n13074), .A2(n12848), .B1(n12847), .B2(n13105), .ZN(
        n12789) );
  NAND2_X1 U15124 ( .A1(n13275), .A2(n12900), .ZN(n12788) );
  NAND4_X1 U15125 ( .A1(n12791), .A2(n12790), .A3(n12789), .A4(n12788), .ZN(
        P2_U3188) );
  OAI21_X1 U15126 ( .B1(n12793), .B2(n12872), .A(n12855), .ZN(n12799) );
  NOR3_X1 U15127 ( .A1(n12793), .A2(n12792), .A3(n12860), .ZN(n12794) );
  OAI21_X1 U15128 ( .B1(n12794), .B2(n12847), .A(n13165), .ZN(n12797) );
  NAND2_X1 U15129 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n12983)
         );
  OAI21_X1 U15130 ( .B1(n12877), .B2(n13144), .A(n12983), .ZN(n12795) );
  AOI21_X1 U15131 ( .B1(n12848), .B2(n13106), .A(n12795), .ZN(n12796) );
  OAI211_X1 U15132 ( .C1(n7027), .C2(n12883), .A(n12797), .B(n12796), .ZN(
        n12798) );
  AOI21_X1 U15133 ( .B1(n12799), .B2(n12871), .A(n12798), .ZN(n12800) );
  INV_X1 U15134 ( .A(n12800), .ZN(P2_U3191) );
  OAI211_X1 U15135 ( .C1(n12803), .C2(n12802), .A(n12801), .B(n12871), .ZN(
        n12807) );
  AOI22_X1 U15136 ( .A1(n13109), .A2(n12888), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12806) );
  AOI22_X1 U15137 ( .A1(n13105), .A2(n12848), .B1(n12847), .B2(n13106), .ZN(
        n12805) );
  NAND2_X1 U15138 ( .A1(n13286), .A2(n12900), .ZN(n12804) );
  NAND4_X1 U15139 ( .A1(n12807), .A2(n12806), .A3(n12805), .A4(n12804), .ZN(
        P2_U3195) );
  INV_X1 U15140 ( .A(n12809), .ZN(n12810) );
  AOI21_X1 U15141 ( .B1(n12808), .B2(n12810), .A(n12902), .ZN(n12815) );
  INV_X1 U15142 ( .A(n12811), .ZN(n12812) );
  NOR3_X1 U15143 ( .A1(n12812), .A2(n13044), .A3(n12860), .ZN(n12814) );
  OAI21_X1 U15144 ( .B1(n12815), .B2(n12814), .A(n12813), .ZN(n12820) );
  OAI22_X1 U15145 ( .A1(n13044), .A2(n12896), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12816), .ZN(n12818) );
  NOR2_X1 U15146 ( .A1(n13043), .A2(n12890), .ZN(n12817) );
  AOI211_X1 U15147 ( .C1(n12888), .C2(n13047), .A(n12818), .B(n12817), .ZN(
        n12819) );
  OAI211_X1 U15148 ( .C1(n13050), .C2(n12883), .A(n12820), .B(n12819), .ZN(
        P2_U3197) );
  OAI21_X1 U15149 ( .B1(n6595), .B2(n12821), .A(n12836), .ZN(n12825) );
  INV_X1 U15150 ( .A(n13189), .ZN(n13311) );
  AOI22_X1 U15151 ( .A1(n12888), .A2(n13192), .B1(P2_REG3_REG_16__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12823) );
  AOI22_X1 U15152 ( .A1(n12847), .A2(n13224), .B1(n12848), .B2(n13186), .ZN(
        n12822) );
  OAI211_X1 U15153 ( .C1(n13311), .C2(n12883), .A(n12823), .B(n12822), .ZN(
        n12824) );
  AOI21_X1 U15154 ( .B1(n12825), .B2(n12871), .A(n12824), .ZN(n12826) );
  INV_X1 U15155 ( .A(n12826), .ZN(P2_U3198) );
  INV_X1 U15156 ( .A(n12827), .ZN(n12839) );
  AOI22_X1 U15157 ( .A1(n12848), .A2(n13165), .B1(n12847), .B2(n13204), .ZN(
        n12829) );
  OAI211_X1 U15158 ( .C1(n12877), .C2(n13169), .A(n12829), .B(n12828), .ZN(
        n12830) );
  AOI21_X1 U15159 ( .B1(n13307), .B2(n12900), .A(n12830), .ZN(n12838) );
  NAND2_X1 U15160 ( .A1(n12831), .A2(n12871), .ZN(n12832) );
  OAI21_X1 U15161 ( .B1(n12833), .B2(n12860), .A(n12832), .ZN(n12834) );
  NAND3_X1 U15162 ( .A1(n12836), .A2(n12835), .A3(n12834), .ZN(n12837) );
  OAI211_X1 U15163 ( .C1(n12839), .C2(n12902), .A(n12838), .B(n12837), .ZN(
        P2_U3200) );
  INV_X1 U15164 ( .A(n13269), .ZN(n13068) );
  NAND2_X1 U15165 ( .A1(n12841), .A2(n12808), .ZN(n12845) );
  OAI22_X1 U15166 ( .A1(n13065), .A2(n12877), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15315), .ZN(n12843) );
  NOR2_X1 U15167 ( .A1(n12866), .A2(n12896), .ZN(n12842) );
  AOI211_X1 U15168 ( .C1(n12848), .C2(n13060), .A(n12843), .B(n12842), .ZN(
        n12844) );
  OAI211_X1 U15169 ( .C1(n13068), .C2(n12883), .A(n12845), .B(n12844), .ZN(
        P2_U3201) );
  INV_X1 U15170 ( .A(n12846), .ZN(n13120) );
  AOI22_X1 U15171 ( .A1(n12888), .A2(n13120), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12850) );
  AOI22_X1 U15172 ( .A1(n13127), .A2(n12848), .B1(n12847), .B2(n13126), .ZN(
        n12849) );
  OAI211_X1 U15173 ( .C1(n13122), .C2(n12883), .A(n12850), .B(n12849), .ZN(
        n12857) );
  OAI22_X1 U15174 ( .A1(n12852), .A2(n12902), .B1(n12851), .B2(n12860), .ZN(
        n12853) );
  AND3_X1 U15175 ( .A1(n12855), .A2(n12854), .A3(n12853), .ZN(n12856) );
  AOI211_X1 U15176 ( .C1(n12871), .C2(n12858), .A(n12857), .B(n12856), .ZN(
        n12859) );
  INV_X1 U15177 ( .A(n12859), .ZN(P2_U3205) );
  OAI22_X1 U15178 ( .A1(n12862), .A2(n12902), .B1(n12861), .B2(n12860), .ZN(
        n12864) );
  NAND2_X1 U15179 ( .A1(n12864), .A2(n12863), .ZN(n12870) );
  NOR2_X1 U15180 ( .A1(n13095), .A2(n12877), .ZN(n12868) );
  OAI22_X1 U15181 ( .A1(n12866), .A2(n12890), .B1(n12865), .B2(n12896), .ZN(
        n12867) );
  AOI211_X1 U15182 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(P2_U3088), .A(n12868), 
        .B(n12867), .ZN(n12869) );
  OAI211_X1 U15183 ( .C1(n7175), .C2(n12883), .A(n12870), .B(n12869), .ZN(
        P2_U3207) );
  INV_X1 U15184 ( .A(n13302), .ZN(n12884) );
  OAI211_X1 U15185 ( .C1(n12874), .C2(n12873), .A(n12872), .B(n12871), .ZN(
        n12882) );
  NAND2_X1 U15186 ( .A1(n13126), .A2(n13223), .ZN(n12876) );
  NAND2_X1 U15187 ( .A1(n13186), .A2(n13225), .ZN(n12875) );
  NAND2_X1 U15188 ( .A1(n12876), .A2(n12875), .ZN(n13155) );
  NAND2_X1 U15189 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14986)
         );
  INV_X1 U15190 ( .A(n14986), .ZN(n12879) );
  NOR2_X1 U15191 ( .A1(n12877), .A2(n13160), .ZN(n12878) );
  AOI211_X1 U15192 ( .C1(n12880), .C2(n13155), .A(n12879), .B(n12878), .ZN(
        n12881) );
  OAI211_X1 U15193 ( .C1(n12884), .C2(n12883), .A(n12882), .B(n12881), .ZN(
        P2_U3210) );
  INV_X1 U15194 ( .A(n12813), .ZN(n12887) );
  INV_X1 U15195 ( .A(n12885), .ZN(n12886) );
  AOI21_X1 U15196 ( .B1(n12894), .B2(n12887), .A(n12886), .ZN(n12903) );
  AOI22_X1 U15197 ( .A1(n13031), .A2(n12888), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12889) );
  OAI21_X1 U15198 ( .B1(n12891), .B2(n12890), .A(n12889), .ZN(n12899) );
  NAND3_X1 U15199 ( .A1(n12894), .A2(n12893), .A3(n12892), .ZN(n12897) );
  AOI21_X1 U15200 ( .B1(n12897), .B2(n12896), .A(n12895), .ZN(n12898) );
  AOI211_X1 U15201 ( .C1(n13259), .C2(n12900), .A(n12899), .B(n12898), .ZN(
        n12901) );
  OAI21_X1 U15202 ( .B1(n12903), .B2(n12902), .A(n12901), .ZN(P2_U3212) );
  INV_X2 U15203 ( .A(P2_U3947), .ZN(n12917) );
  MUX2_X1 U15204 ( .A(n12986), .B(P2_DATAO_REG_31__SCAN_IN), .S(n12917), .Z(
        P2_U3562) );
  MUX2_X1 U15205 ( .A(n12904), .B(P2_DATAO_REG_30__SCAN_IN), .S(n12917), .Z(
        P2_U3561) );
  MUX2_X1 U15206 ( .A(n12905), .B(P2_DATAO_REG_29__SCAN_IN), .S(n12917), .Z(
        P2_U3560) );
  MUX2_X1 U15207 ( .A(n13011), .B(P2_DATAO_REG_28__SCAN_IN), .S(n12917), .Z(
        P2_U3559) );
  MUX2_X1 U15208 ( .A(n13027), .B(P2_DATAO_REG_27__SCAN_IN), .S(n12917), .Z(
        P2_U3558) );
  MUX2_X1 U15209 ( .A(n13012), .B(P2_DATAO_REG_26__SCAN_IN), .S(n12917), .Z(
        P2_U3557) );
  MUX2_X1 U15210 ( .A(n13060), .B(P2_DATAO_REG_25__SCAN_IN), .S(n12917), .Z(
        P2_U3556) );
  MUX2_X1 U15211 ( .A(n13074), .B(P2_DATAO_REG_24__SCAN_IN), .S(n12917), .Z(
        P2_U3555) );
  MUX2_X1 U15212 ( .A(n13087), .B(P2_DATAO_REG_23__SCAN_IN), .S(n12917), .Z(
        P2_U3554) );
  MUX2_X1 U15213 ( .A(n13105), .B(P2_DATAO_REG_22__SCAN_IN), .S(n12917), .Z(
        P2_U3553) );
  MUX2_X1 U15214 ( .A(n13127), .B(P2_DATAO_REG_21__SCAN_IN), .S(n12917), .Z(
        P2_U3552) );
  MUX2_X1 U15215 ( .A(n13106), .B(P2_DATAO_REG_20__SCAN_IN), .S(n12917), .Z(
        P2_U3551) );
  MUX2_X1 U15216 ( .A(n13126), .B(P2_DATAO_REG_19__SCAN_IN), .S(n12917), .Z(
        P2_U3550) );
  MUX2_X1 U15217 ( .A(n13165), .B(P2_DATAO_REG_18__SCAN_IN), .S(n12917), .Z(
        P2_U3549) );
  MUX2_X1 U15218 ( .A(n13186), .B(P2_DATAO_REG_17__SCAN_IN), .S(n12917), .Z(
        P2_U3548) );
  MUX2_X1 U15219 ( .A(n13204), .B(P2_DATAO_REG_16__SCAN_IN), .S(n12917), .Z(
        P2_U3547) );
  MUX2_X1 U15220 ( .A(n13224), .B(P2_DATAO_REG_15__SCAN_IN), .S(n12917), .Z(
        P2_U3546) );
  MUX2_X1 U15221 ( .A(n13203), .B(P2_DATAO_REG_14__SCAN_IN), .S(n12917), .Z(
        P2_U3545) );
  MUX2_X1 U15222 ( .A(n13226), .B(P2_DATAO_REG_13__SCAN_IN), .S(n12917), .Z(
        P2_U3544) );
  MUX2_X1 U15223 ( .A(n12906), .B(P2_DATAO_REG_12__SCAN_IN), .S(n12917), .Z(
        P2_U3543) );
  MUX2_X1 U15224 ( .A(n12907), .B(P2_DATAO_REG_11__SCAN_IN), .S(n12917), .Z(
        P2_U3542) );
  MUX2_X1 U15225 ( .A(n12908), .B(P2_DATAO_REG_10__SCAN_IN), .S(n12917), .Z(
        P2_U3541) );
  MUX2_X1 U15226 ( .A(n12909), .B(P2_DATAO_REG_9__SCAN_IN), .S(n12917), .Z(
        P2_U3540) );
  MUX2_X1 U15227 ( .A(n12910), .B(P2_DATAO_REG_8__SCAN_IN), .S(n12917), .Z(
        P2_U3539) );
  MUX2_X1 U15228 ( .A(n12911), .B(P2_DATAO_REG_7__SCAN_IN), .S(n12917), .Z(
        P2_U3538) );
  MUX2_X1 U15229 ( .A(n12912), .B(P2_DATAO_REG_6__SCAN_IN), .S(n12917), .Z(
        P2_U3537) );
  MUX2_X1 U15230 ( .A(n12913), .B(P2_DATAO_REG_5__SCAN_IN), .S(n12917), .Z(
        P2_U3536) );
  MUX2_X1 U15231 ( .A(n12914), .B(P2_DATAO_REG_4__SCAN_IN), .S(n12917), .Z(
        P2_U3535) );
  MUX2_X1 U15232 ( .A(n12915), .B(P2_DATAO_REG_3__SCAN_IN), .S(n12917), .Z(
        P2_U3534) );
  MUX2_X1 U15233 ( .A(n12916), .B(P2_DATAO_REG_2__SCAN_IN), .S(n12917), .Z(
        P2_U3533) );
  MUX2_X1 U15234 ( .A(n9755), .B(P2_DATAO_REG_1__SCAN_IN), .S(n12917), .Z(
        P2_U3532) );
  OAI211_X1 U15235 ( .C1(n12920), .C2(n12919), .A(n14985), .B(n12918), .ZN(
        n12929) );
  OAI211_X1 U15236 ( .C1(n12923), .C2(n12922), .A(n14977), .B(n12921), .ZN(
        n12928) );
  AOI22_X1 U15237 ( .A1(n14823), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n12927) );
  INV_X1 U15238 ( .A(n12924), .ZN(n12925) );
  NAND2_X1 U15239 ( .A1(n14971), .A2(n12925), .ZN(n12926) );
  NAND4_X1 U15240 ( .A1(n12929), .A2(n12928), .A3(n12927), .A4(n12926), .ZN(
        P2_U3216) );
  INV_X1 U15241 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n12931) );
  OAI21_X1 U15242 ( .B1(n14988), .B2(n12931), .A(n12930), .ZN(n12932) );
  AOI21_X1 U15243 ( .B1(n12933), .B2(n14971), .A(n12932), .ZN(n12942) );
  OAI211_X1 U15244 ( .C1(n12936), .C2(n12935), .A(n14977), .B(n12934), .ZN(
        n12941) );
  OAI211_X1 U15245 ( .C1(n12939), .C2(n12938), .A(n14985), .B(n12937), .ZN(
        n12940) );
  NAND3_X1 U15246 ( .A1(n12942), .A2(n12941), .A3(n12940), .ZN(P2_U3219) );
  INV_X1 U15247 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n14385) );
  NAND2_X1 U15248 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n12943) );
  OAI21_X1 U15249 ( .B1(n14988), .B2(n14385), .A(n12943), .ZN(n12944) );
  AOI21_X1 U15250 ( .B1(n12945), .B2(n14971), .A(n12944), .ZN(n12954) );
  OAI211_X1 U15251 ( .C1(n12948), .C2(n12947), .A(n14985), .B(n12946), .ZN(
        n12953) );
  OAI211_X1 U15252 ( .C1(n12951), .C2(n12950), .A(n14977), .B(n12949), .ZN(
        n12952) );
  NAND3_X1 U15253 ( .A1(n12954), .A2(n12953), .A3(n12952), .ZN(P2_U3220) );
  INV_X1 U15254 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14392) );
  NAND2_X1 U15255 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n12955) );
  OAI21_X1 U15256 ( .B1(n14988), .B2(n14392), .A(n12955), .ZN(n12956) );
  AOI21_X1 U15257 ( .B1(n12957), .B2(n14971), .A(n12956), .ZN(n12966) );
  OAI211_X1 U15258 ( .C1(n12960), .C2(n12959), .A(n12958), .B(n14985), .ZN(
        n12965) );
  OAI211_X1 U15259 ( .C1(n12963), .C2(n12962), .A(n14977), .B(n12961), .ZN(
        n12964) );
  NAND3_X1 U15260 ( .A1(n12966), .A2(n12965), .A3(n12964), .ZN(P2_U3221) );
  NAND2_X1 U15261 ( .A1(n12974), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n12967) );
  NAND2_X1 U15262 ( .A1(n12968), .A2(n12967), .ZN(n12970) );
  XOR2_X1 U15263 ( .A(n12969), .B(n12970), .Z(n14976) );
  INV_X1 U15264 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n15242) );
  NAND2_X1 U15265 ( .A1(n14976), .A2(n15242), .ZN(n14975) );
  OR2_X1 U15266 ( .A1(n12970), .A2(n12969), .ZN(n12971) );
  NAND2_X1 U15267 ( .A1(n14975), .A2(n12971), .ZN(n12972) );
  XNOR2_X1 U15268 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n12972), .ZN(n12980) );
  INV_X1 U15269 ( .A(n12980), .ZN(n12978) );
  AOI21_X1 U15270 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n12974), .A(n12973), 
        .ZN(n12975) );
  NOR2_X1 U15271 ( .A1(n12975), .A2(n14980), .ZN(n12976) );
  OAI21_X1 U15272 ( .B1(n12979), .B2(n14960), .A(n14979), .ZN(n12977) );
  AOI21_X1 U15273 ( .B1(n12978), .B2(n14985), .A(n12977), .ZN(n12982) );
  AOI22_X1 U15274 ( .A1(n12980), .A2(n14985), .B1(n14977), .B2(n12979), .ZN(
        n12981) );
  MUX2_X1 U15275 ( .A(n12982), .B(n12981), .S(n13230), .Z(n12984) );
  OAI211_X1 U15276 ( .C1(n7652), .C2(n14988), .A(n12984), .B(n12983), .ZN(
        P2_U3233) );
  XOR2_X1 U15277 ( .A(n13237), .B(n12990), .Z(n13239) );
  NAND2_X1 U15278 ( .A1(n12986), .A2(n12985), .ZN(n13241) );
  NOR2_X1 U15279 ( .A1(n13212), .A2(n13241), .ZN(n12993) );
  AOI21_X1 U15280 ( .B1(n13212), .B2(P2_REG2_REG_31__SCAN_IN), .A(n12993), 
        .ZN(n12988) );
  NAND2_X1 U15281 ( .A1(n13237), .A2(n13234), .ZN(n12987) );
  OAI211_X1 U15282 ( .C1(n13239), .C2(n12989), .A(n12988), .B(n12987), .ZN(
        P2_U3234) );
  INV_X1 U15283 ( .A(n12992), .ZN(n13243) );
  AOI21_X1 U15284 ( .B1(n12992), .B2(n12991), .A(n12990), .ZN(n13240) );
  NAND2_X1 U15285 ( .A1(n13240), .A2(n13131), .ZN(n12995) );
  AOI21_X1 U15286 ( .B1(n13212), .B2(P2_REG2_REG_30__SCAN_IN), .A(n12993), 
        .ZN(n12994) );
  OAI211_X1 U15287 ( .C1(n13243), .C2(n13147), .A(n12995), .B(n12994), .ZN(
        P2_U3235) );
  OAI21_X1 U15288 ( .B1(n12997), .B2(n7282), .A(n12996), .ZN(n13253) );
  OAI211_X1 U15289 ( .C1(n13000), .C2(n12999), .A(n12998), .B(n13228), .ZN(
        n13002) );
  OR2_X1 U15290 ( .A1(n13003), .A2(n13018), .ZN(n13004) );
  AND3_X1 U15291 ( .A1(n13005), .A2(n13291), .A3(n13004), .ZN(n13249) );
  AOI22_X1 U15292 ( .A1(n13249), .A2(n13230), .B1(n13209), .B2(n13006), .ZN(
        n13007) );
  AOI21_X1 U15293 ( .B1(n13252), .B2(n13007), .A(n13212), .ZN(n13008) );
  INV_X1 U15294 ( .A(n13008), .ZN(n13010) );
  AOI22_X1 U15295 ( .A1(n13250), .A2(n13234), .B1(n13212), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n13009) );
  OAI211_X1 U15296 ( .C1(n13236), .C2(n13253), .A(n13010), .B(n13009), .ZN(
        P2_U3237) );
  INV_X1 U15297 ( .A(n13258), .ZN(n13024) );
  NAND2_X1 U15298 ( .A1(n13255), .A2(n13029), .ZN(n13016) );
  NAND2_X1 U15299 ( .A1(n13016), .A2(n13291), .ZN(n13017) );
  NOR2_X1 U15300 ( .A1(n13018), .A2(n13017), .ZN(n13254) );
  NAND2_X1 U15301 ( .A1(n13254), .A2(n13175), .ZN(n13021) );
  AOI22_X1 U15302 ( .A1(n13019), .A2(n13209), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n13212), .ZN(n13020) );
  OAI211_X1 U15303 ( .C1(n6945), .C2(n13147), .A(n13021), .B(n13020), .ZN(
        n13022) );
  AOI21_X1 U15304 ( .B1(n13024), .B2(n13023), .A(n13022), .ZN(n13025) );
  OAI21_X1 U15305 ( .B1(n13257), .B2(n13212), .A(n13025), .ZN(P2_U3238) );
  AOI222_X1 U15306 ( .A1(n13228), .A2(n13028), .B1(n13027), .B2(n13223), .C1(
        n13060), .C2(n13225), .ZN(n13262) );
  INV_X1 U15307 ( .A(n13029), .ZN(n13030) );
  AOI21_X1 U15308 ( .B1(n13259), .B2(n13046), .A(n13030), .ZN(n13260) );
  AOI22_X1 U15309 ( .A1(n13031), .A2(n13209), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n13212), .ZN(n13032) );
  OAI21_X1 U15310 ( .B1(n13033), .B2(n13147), .A(n13032), .ZN(n13036) );
  XOR2_X1 U15311 ( .A(n13035), .B(n13034), .Z(n13263) );
  OAI21_X1 U15312 ( .B1(n13262), .B2(n13212), .A(n13037), .ZN(P2_U3239) );
  XNOR2_X1 U15313 ( .A(n13038), .B(n13040), .ZN(n13268) );
  AOI21_X1 U15314 ( .B1(n13041), .B2(n13040), .A(n13039), .ZN(n13042) );
  OAI222_X1 U15315 ( .A1(n13139), .A2(n13044), .B1(n13141), .B2(n13043), .C1(
        n13137), .C2(n13042), .ZN(n13264) );
  OR2_X1 U15316 ( .A1(n13064), .A2(n13050), .ZN(n13045) );
  AND3_X1 U15317 ( .A1(n13046), .A2(n13291), .A3(n13045), .ZN(n13265) );
  NAND2_X1 U15318 ( .A1(n13265), .A2(n13175), .ZN(n13049) );
  AOI22_X1 U15319 ( .A1(n13047), .A2(n13209), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n13212), .ZN(n13048) );
  OAI211_X1 U15320 ( .C1(n13050), .C2(n13147), .A(n13049), .B(n13048), .ZN(
        n13051) );
  AOI21_X1 U15321 ( .B1(n13264), .B2(n13219), .A(n13051), .ZN(n13052) );
  OAI21_X1 U15322 ( .B1(n13268), .B2(n13236), .A(n13052), .ZN(P2_U3240) );
  NAND2_X1 U15323 ( .A1(n13053), .A2(n13056), .ZN(n13054) );
  NAND2_X1 U15324 ( .A1(n13055), .A2(n13054), .ZN(n13272) );
  NOR2_X1 U15325 ( .A1(n13057), .A2(n13056), .ZN(n13059) );
  OAI21_X1 U15326 ( .B1(n13059), .B2(n13058), .A(n13228), .ZN(n13062) );
  AOI22_X1 U15327 ( .A1(n13060), .A2(n13223), .B1(n13225), .B2(n13087), .ZN(
        n13061) );
  OAI211_X1 U15328 ( .C1(n13272), .C2(n9771), .A(n13062), .B(n13061), .ZN(
        n13274) );
  NAND2_X1 U15329 ( .A1(n13274), .A2(n13219), .ZN(n13071) );
  AND2_X1 U15330 ( .A1(n13076), .A2(n13269), .ZN(n13063) );
  NOR2_X1 U15331 ( .A1(n13064), .A2(n13063), .ZN(n13270) );
  INV_X1 U15332 ( .A(n13065), .ZN(n13066) );
  AOI22_X1 U15333 ( .A1(n13066), .A2(n13209), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n13212), .ZN(n13067) );
  OAI21_X1 U15334 ( .B1(n13068), .B2(n13147), .A(n13067), .ZN(n13069) );
  AOI21_X1 U15335 ( .B1(n13270), .B2(n13131), .A(n13069), .ZN(n13070) );
  OAI211_X1 U15336 ( .C1(n13272), .C2(n13072), .A(n13071), .B(n13070), .ZN(
        P2_U3241) );
  XOR2_X1 U15337 ( .A(n13073), .B(n13081), .Z(n13075) );
  AOI222_X1 U15338 ( .A1(n13228), .A2(n13075), .B1(n13074), .B2(n13223), .C1(
        n13105), .C2(n13225), .ZN(n13278) );
  INV_X1 U15339 ( .A(n13076), .ZN(n13077) );
  AOI21_X1 U15340 ( .B1(n13275), .B2(n13098), .A(n13077), .ZN(n13276) );
  AOI22_X1 U15341 ( .A1(n13078), .A2(n13209), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n13212), .ZN(n13079) );
  OAI21_X1 U15342 ( .B1(n7173), .B2(n13147), .A(n13079), .ZN(n13083) );
  XOR2_X1 U15343 ( .A(n13081), .B(n13080), .Z(n13279) );
  NOR2_X1 U15344 ( .A1(n13279), .A2(n13236), .ZN(n13082) );
  AOI211_X1 U15345 ( .C1(n13276), .C2(n13131), .A(n13083), .B(n13082), .ZN(
        n13084) );
  OAI21_X1 U15346 ( .B1(n13212), .B2(n13278), .A(n13084), .ZN(P2_U3242) );
  OAI211_X1 U15347 ( .C1(n13091), .C2(n13086), .A(n13085), .B(n13228), .ZN(
        n13089) );
  AOI22_X1 U15348 ( .A1(n13087), .A2(n13223), .B1(n13225), .B2(n13127), .ZN(
        n13088) );
  NAND2_X1 U15349 ( .A1(n13091), .A2(n13090), .ZN(n13092) );
  NAND2_X1 U15350 ( .A1(n13093), .A2(n13092), .ZN(n13284) );
  INV_X1 U15351 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13094) );
  OAI22_X1 U15352 ( .A1(n13095), .A2(n13217), .B1(n13094), .B2(n13219), .ZN(
        n13096) );
  AOI21_X1 U15353 ( .B1(n13280), .B2(n13234), .A(n13096), .ZN(n13100) );
  NAND2_X1 U15354 ( .A1(n13280), .A2(n13108), .ZN(n13097) );
  AND2_X1 U15355 ( .A1(n13098), .A2(n13097), .ZN(n13281) );
  NAND2_X1 U15356 ( .A1(n13281), .A2(n13131), .ZN(n13099) );
  OAI211_X1 U15357 ( .C1(n13284), .C2(n13236), .A(n13100), .B(n13099), .ZN(
        n13101) );
  INV_X1 U15358 ( .A(n13101), .ZN(n13102) );
  OAI21_X1 U15359 ( .B1(n13212), .B2(n13283), .A(n13102), .ZN(P2_U3243) );
  XNOR2_X1 U15360 ( .A(n13104), .B(n13103), .ZN(n13107) );
  AOI222_X1 U15361 ( .A1(n13228), .A2(n13107), .B1(n13106), .B2(n13225), .C1(
        n13105), .C2(n13223), .ZN(n13288) );
  AOI211_X1 U15362 ( .C1(n13286), .C2(n13118), .A(n15030), .B(n7176), .ZN(
        n13285) );
  INV_X1 U15363 ( .A(n13286), .ZN(n13111) );
  AOI22_X1 U15364 ( .A1(n13109), .A2(n13209), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n13212), .ZN(n13110) );
  OAI21_X1 U15365 ( .B1(n13111), .B2(n13147), .A(n13110), .ZN(n13115) );
  XNOR2_X1 U15366 ( .A(n13113), .B(n13112), .ZN(n13289) );
  NOR2_X1 U15367 ( .A1(n13289), .A2(n13236), .ZN(n13114) );
  AOI211_X1 U15368 ( .C1(n13285), .C2(n13175), .A(n13115), .B(n13114), .ZN(
        n13116) );
  OAI21_X1 U15369 ( .B1(n13212), .B2(n13288), .A(n13116), .ZN(P2_U3244) );
  XOR2_X1 U15370 ( .A(n13117), .B(n13123), .Z(n13295) );
  INV_X1 U15371 ( .A(n13118), .ZN(n13119) );
  AOI21_X1 U15372 ( .B1(n13290), .B2(n13142), .A(n13119), .ZN(n13292) );
  AOI22_X1 U15373 ( .A1(n13120), .A2(n13209), .B1(P2_REG2_REG_20__SCAN_IN), 
        .B2(n13212), .ZN(n13121) );
  OAI21_X1 U15374 ( .B1(n13122), .B2(n13147), .A(n13121), .ZN(n13130) );
  INV_X1 U15375 ( .A(n13123), .ZN(n13125) );
  OAI21_X1 U15376 ( .B1(n13125), .B2(n6538), .A(n13124), .ZN(n13128) );
  AOI222_X1 U15377 ( .A1(n13228), .A2(n13128), .B1(n13127), .B2(n13223), .C1(
        n13126), .C2(n13225), .ZN(n13294) );
  NOR2_X1 U15378 ( .A1(n13294), .A2(n13212), .ZN(n13129) );
  AOI211_X1 U15379 ( .C1(n13292), .C2(n13131), .A(n13130), .B(n13129), .ZN(
        n13132) );
  OAI21_X1 U15380 ( .B1(n13295), .B2(n13236), .A(n13132), .ZN(P2_U3245) );
  XNOR2_X1 U15381 ( .A(n13133), .B(n13135), .ZN(n13300) );
  XOR2_X1 U15382 ( .A(n13135), .B(n13134), .Z(n13136) );
  OAI222_X1 U15383 ( .A1(n13141), .A2(n13140), .B1(n13139), .B2(n13138), .C1(
        n13137), .C2(n13136), .ZN(n13296) );
  NAND2_X1 U15384 ( .A1(n13296), .A2(n13219), .ZN(n13150) );
  INV_X1 U15385 ( .A(n13142), .ZN(n13143) );
  AOI211_X1 U15386 ( .C1(n13298), .C2(n13157), .A(n15030), .B(n13143), .ZN(
        n13297) );
  INV_X1 U15387 ( .A(n13144), .ZN(n13145) );
  AOI22_X1 U15388 ( .A1(n13145), .A2(n13209), .B1(n13212), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n13146) );
  OAI21_X1 U15389 ( .B1(n7027), .B2(n13147), .A(n13146), .ZN(n13148) );
  AOI21_X1 U15390 ( .B1(n13297), .B2(n13175), .A(n13148), .ZN(n13149) );
  OAI211_X1 U15391 ( .C1(n13236), .C2(n13300), .A(n13150), .B(n13149), .ZN(
        P2_U3246) );
  AOI21_X1 U15392 ( .B1(n13152), .B2(n13151), .A(n6587), .ZN(n13305) );
  AOI22_X1 U15393 ( .A1(n13302), .A2(n13234), .B1(n13212), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n13163) );
  XNOR2_X1 U15394 ( .A(n13154), .B(n13153), .ZN(n13156) );
  AOI21_X1 U15395 ( .B1(n13156), .B2(n13228), .A(n13155), .ZN(n13304) );
  AOI21_X1 U15396 ( .B1(n13174), .B2(n13302), .A(n15030), .ZN(n13158) );
  AND2_X1 U15397 ( .A1(n13158), .A2(n13157), .ZN(n13301) );
  NAND2_X1 U15398 ( .A1(n13301), .A2(n13230), .ZN(n13159) );
  OAI211_X1 U15399 ( .C1(n13217), .C2(n13160), .A(n13304), .B(n13159), .ZN(
        n13161) );
  NAND2_X1 U15400 ( .A1(n13161), .A2(n13219), .ZN(n13162) );
  OAI211_X1 U15401 ( .C1(n13305), .C2(n13236), .A(n13163), .B(n13162), .ZN(
        P2_U3247) );
  XNOR2_X1 U15402 ( .A(n13164), .B(n13167), .ZN(n13166) );
  AOI222_X1 U15403 ( .A1(n13228), .A2(n13166), .B1(n13204), .B2(n13225), .C1(
        n13165), .C2(n13223), .ZN(n13309) );
  XNOR2_X1 U15404 ( .A(n13168), .B(n13167), .ZN(n13310) );
  OAI22_X1 U15405 ( .A1(n13219), .A2(n13170), .B1(n13169), .B2(n13217), .ZN(
        n13171) );
  AOI21_X1 U15406 ( .B1(n13307), .B2(n13234), .A(n13171), .ZN(n13177) );
  OR2_X1 U15407 ( .A1(n13172), .A2(n13190), .ZN(n13173) );
  AND3_X1 U15408 ( .A1(n13174), .A2(n13173), .A3(n13291), .ZN(n13306) );
  NAND2_X1 U15409 ( .A1(n13306), .A2(n13175), .ZN(n13176) );
  OAI211_X1 U15410 ( .C1(n13310), .C2(n13236), .A(n13177), .B(n13176), .ZN(
        n13178) );
  INV_X1 U15411 ( .A(n13178), .ZN(n13179) );
  OAI21_X1 U15412 ( .B1(n13309), .B2(n13212), .A(n13179), .ZN(P2_U3248) );
  INV_X1 U15413 ( .A(n13180), .ZN(n13181) );
  AOI21_X1 U15414 ( .B1(n13184), .B2(n13182), .A(n13181), .ZN(n13315) );
  INV_X1 U15415 ( .A(n13315), .ZN(n13198) );
  AOI22_X1 U15416 ( .A1(n13189), .A2(n13234), .B1(P2_REG2_REG_16__SCAN_IN), 
        .B2(n13212), .ZN(n13197) );
  OAI211_X1 U15417 ( .C1(n13185), .C2(n13184), .A(n13183), .B(n13228), .ZN(
        n13188) );
  AOI22_X1 U15418 ( .A1(n13186), .A2(n13223), .B1(n13225), .B2(n13224), .ZN(
        n13187) );
  NAND2_X1 U15419 ( .A1(n13188), .A2(n13187), .ZN(n13314) );
  AND2_X1 U15420 ( .A1(n13189), .A2(n13206), .ZN(n13191) );
  OR2_X1 U15421 ( .A1(n13191), .A2(n13190), .ZN(n13312) );
  INV_X1 U15422 ( .A(n13192), .ZN(n13193) );
  OAI22_X1 U15423 ( .A1(n13312), .A2(n13194), .B1(n13193), .B2(n13217), .ZN(
        n13195) );
  OAI21_X1 U15424 ( .B1(n13314), .B2(n13195), .A(n13219), .ZN(n13196) );
  OAI211_X1 U15425 ( .C1(n13198), .C2(n13236), .A(n13197), .B(n13196), .ZN(
        P2_U3249) );
  XNOR2_X1 U15426 ( .A(n13200), .B(n13199), .ZN(n13321) );
  XNOR2_X1 U15427 ( .A(n13202), .B(n13201), .ZN(n13205) );
  AOI222_X1 U15428 ( .A1(n13228), .A2(n13205), .B1(n13204), .B2(n13223), .C1(
        n13203), .C2(n13225), .ZN(n13320) );
  AOI21_X1 U15429 ( .B1(n13229), .B2(n13318), .A(n15030), .ZN(n13207) );
  AND2_X1 U15430 ( .A1(n13207), .A2(n13206), .ZN(n13317) );
  AOI22_X1 U15431 ( .A1(n13317), .A2(n13230), .B1(n13209), .B2(n13208), .ZN(
        n13210) );
  AOI21_X1 U15432 ( .B1(n13320), .B2(n13210), .A(n13212), .ZN(n13211) );
  INV_X1 U15433 ( .A(n13211), .ZN(n13214) );
  AOI22_X1 U15434 ( .A1(n13318), .A2(n13234), .B1(n13212), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n13213) );
  OAI211_X1 U15435 ( .C1(n13321), .C2(n13236), .A(n13214), .B(n13213), .ZN(
        P2_U3250) );
  XNOR2_X1 U15436 ( .A(n13216), .B(n13215), .ZN(n13326) );
  OAI22_X1 U15437 ( .A1(n13219), .A2(n14938), .B1(n13218), .B2(n13217), .ZN(
        n13233) );
  OAI21_X1 U15438 ( .B1(n13222), .B2(n13221), .A(n13220), .ZN(n13227) );
  AOI222_X1 U15439 ( .A1(n13228), .A2(n13227), .B1(n13226), .B2(n13225), .C1(
        n13224), .C2(n13223), .ZN(n13324) );
  AOI211_X1 U15440 ( .C1(n13323), .C2(n6944), .A(n15030), .B(n6942), .ZN(
        n13322) );
  NAND2_X1 U15441 ( .A1(n13322), .A2(n13230), .ZN(n13231) );
  AOI21_X1 U15442 ( .B1(n13324), .B2(n13231), .A(n13212), .ZN(n13232) );
  AOI211_X1 U15443 ( .C1(n13234), .C2(n13323), .A(n13233), .B(n13232), .ZN(
        n13235) );
  OAI21_X1 U15444 ( .B1(n13236), .B2(n13326), .A(n13235), .ZN(P2_U3251) );
  NAND2_X1 U15445 ( .A1(n13237), .A2(n15019), .ZN(n13238) );
  OAI211_X1 U15446 ( .C1(n13239), .C2(n15030), .A(n13241), .B(n13238), .ZN(
        n13328) );
  MUX2_X1 U15447 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13328), .S(n15047), .Z(
        P2_U3530) );
  INV_X1 U15448 ( .A(n15019), .ZN(n15028) );
  NAND2_X1 U15449 ( .A1(n13240), .A2(n13291), .ZN(n13242) );
  OAI211_X1 U15450 ( .C1(n13243), .C2(n15028), .A(n13242), .B(n13241), .ZN(
        n13329) );
  MUX2_X1 U15451 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13329), .S(n15047), .Z(
        P2_U3529) );
  AOI22_X1 U15452 ( .A1(n13245), .A2(n13291), .B1(n15019), .B2(n13244), .ZN(
        n13246) );
  OAI211_X1 U15453 ( .C1(n13248), .C2(n13327), .A(n13247), .B(n13246), .ZN(
        n13330) );
  MUX2_X1 U15454 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13330), .S(n15047), .Z(
        P2_U3528) );
  AOI21_X1 U15455 ( .B1(n15019), .B2(n13250), .A(n13249), .ZN(n13251) );
  OAI211_X1 U15456 ( .C1(n13327), .C2(n13253), .A(n13252), .B(n13251), .ZN(
        n13331) );
  MUX2_X1 U15457 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13331), .S(n15047), .Z(
        P2_U3527) );
  AOI21_X1 U15458 ( .B1(n15019), .B2(n13255), .A(n13254), .ZN(n13256) );
  OAI211_X1 U15459 ( .C1(n13327), .C2(n13258), .A(n13257), .B(n13256), .ZN(
        n13332) );
  MUX2_X1 U15460 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13332), .S(n15047), .Z(
        P2_U3526) );
  AOI22_X1 U15461 ( .A1(n13260), .A2(n13291), .B1(n15019), .B2(n13259), .ZN(
        n13261) );
  MUX2_X1 U15462 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13333), .S(n15047), .Z(
        P2_U3525) );
  AOI211_X1 U15463 ( .C1(n15019), .C2(n13266), .A(n13265), .B(n13264), .ZN(
        n13267) );
  OAI21_X1 U15464 ( .B1(n13327), .B2(n13268), .A(n13267), .ZN(n13334) );
  MUX2_X1 U15465 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13334), .S(n15047), .Z(
        P2_U3524) );
  AOI22_X1 U15466 ( .A1(n13270), .A2(n13291), .B1(n15019), .B2(n13269), .ZN(
        n13271) );
  OAI21_X1 U15467 ( .B1(n13272), .B2(n15023), .A(n13271), .ZN(n13273) );
  OR2_X1 U15468 ( .A1(n13274), .A2(n13273), .ZN(n13335) );
  MUX2_X1 U15469 ( .A(n13335), .B(P2_REG1_REG_24__SCAN_IN), .S(n15045), .Z(
        P2_U3523) );
  AOI22_X1 U15470 ( .A1(n13276), .A2(n13291), .B1(n15019), .B2(n13275), .ZN(
        n13277) );
  OAI211_X1 U15471 ( .C1(n13327), .C2(n13279), .A(n13278), .B(n13277), .ZN(
        n13336) );
  MUX2_X1 U15472 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13336), .S(n15047), .Z(
        P2_U3522) );
  AOI22_X1 U15473 ( .A1(n13281), .A2(n13291), .B1(n15019), .B2(n13280), .ZN(
        n13282) );
  OAI211_X1 U15474 ( .C1(n13284), .C2(n13327), .A(n13283), .B(n13282), .ZN(
        n13337) );
  MUX2_X1 U15475 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13337), .S(n15047), .Z(
        P2_U3521) );
  AOI21_X1 U15476 ( .B1(n15019), .B2(n13286), .A(n13285), .ZN(n13287) );
  OAI211_X1 U15477 ( .C1(n13327), .C2(n13289), .A(n13288), .B(n13287), .ZN(
        n13338) );
  MUX2_X1 U15478 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13338), .S(n15047), .Z(
        P2_U3520) );
  AOI22_X1 U15479 ( .A1(n13292), .A2(n13291), .B1(n15019), .B2(n13290), .ZN(
        n13293) );
  OAI211_X1 U15480 ( .C1(n13327), .C2(n13295), .A(n13294), .B(n13293), .ZN(
        n13339) );
  MUX2_X1 U15481 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13339), .S(n15047), .Z(
        P2_U3519) );
  AOI211_X1 U15482 ( .C1(n15019), .C2(n13298), .A(n13297), .B(n13296), .ZN(
        n13299) );
  OAI21_X1 U15483 ( .B1(n13327), .B2(n13300), .A(n13299), .ZN(n13340) );
  MUX2_X1 U15484 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13340), .S(n15047), .Z(
        P2_U3518) );
  AOI21_X1 U15485 ( .B1(n15019), .B2(n13302), .A(n13301), .ZN(n13303) );
  OAI211_X1 U15486 ( .C1(n13305), .C2(n13327), .A(n13304), .B(n13303), .ZN(
        n13341) );
  MUX2_X1 U15487 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13341), .S(n15047), .Z(
        P2_U3517) );
  AOI21_X1 U15488 ( .B1(n15019), .B2(n13307), .A(n13306), .ZN(n13308) );
  OAI211_X1 U15489 ( .C1(n13327), .C2(n13310), .A(n13309), .B(n13308), .ZN(
        n13342) );
  MUX2_X1 U15490 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13342), .S(n15047), .Z(
        P2_U3516) );
  INV_X1 U15491 ( .A(n13327), .ZN(n15014) );
  OAI22_X1 U15492 ( .A1(n13312), .A2(n15030), .B1(n13311), .B2(n15028), .ZN(
        n13313) );
  AOI211_X1 U15493 ( .C1(n13315), .C2(n15014), .A(n13314), .B(n13313), .ZN(
        n13316) );
  INV_X1 U15494 ( .A(n13316), .ZN(n13343) );
  MUX2_X1 U15495 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13343), .S(n15047), .Z(
        P2_U3515) );
  AOI21_X1 U15496 ( .B1(n15019), .B2(n13318), .A(n13317), .ZN(n13319) );
  OAI211_X1 U15497 ( .C1(n13327), .C2(n13321), .A(n13320), .B(n13319), .ZN(
        n13344) );
  MUX2_X1 U15498 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13344), .S(n15047), .Z(
        P2_U3514) );
  AOI21_X1 U15499 ( .B1(n15019), .B2(n13323), .A(n13322), .ZN(n13325) );
  OAI211_X1 U15500 ( .C1(n13327), .C2(n13326), .A(n13325), .B(n13324), .ZN(
        n13345) );
  MUX2_X1 U15501 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13345), .S(n15047), .Z(
        P2_U3513) );
  MUX2_X1 U15502 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13328), .S(n15026), .Z(
        P2_U3498) );
  MUX2_X1 U15503 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13329), .S(n15026), .Z(
        P2_U3497) );
  MUX2_X1 U15504 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13330), .S(n15026), .Z(
        P2_U3496) );
  MUX2_X1 U15505 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13331), .S(n15026), .Z(
        P2_U3495) );
  MUX2_X1 U15506 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13332), .S(n15026), .Z(
        P2_U3494) );
  MUX2_X1 U15507 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13333), .S(n15026), .Z(
        P2_U3493) );
  MUX2_X1 U15508 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13334), .S(n15026), .Z(
        P2_U3492) );
  MUX2_X1 U15509 ( .A(n13335), .B(P2_REG0_REG_24__SCAN_IN), .S(n15037), .Z(
        P2_U3491) );
  MUX2_X1 U15510 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13336), .S(n15026), .Z(
        P2_U3490) );
  MUX2_X1 U15511 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13337), .S(n15026), .Z(
        P2_U3489) );
  MUX2_X1 U15512 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13338), .S(n15026), .Z(
        P2_U3488) );
  MUX2_X1 U15513 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13339), .S(n15026), .Z(
        P2_U3487) );
  MUX2_X1 U15514 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13340), .S(n15026), .Z(
        P2_U3486) );
  MUX2_X1 U15515 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13341), .S(n15026), .Z(
        P2_U3484) );
  MUX2_X1 U15516 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13342), .S(n15026), .Z(
        P2_U3481) );
  MUX2_X1 U15517 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13343), .S(n15026), .Z(
        P2_U3478) );
  MUX2_X1 U15518 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13344), .S(n15026), .Z(
        P2_U3475) );
  MUX2_X1 U15519 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13345), .S(n15026), .Z(
        P2_U3472) );
  INV_X1 U15520 ( .A(n13501), .ZN(n13348) );
  NOR4_X1 U15521 ( .A1(n7317), .A2(P2_IR_REG_30__SCAN_IN), .A3(n7710), .A4(
        P2_U3088), .ZN(n13346) );
  AOI21_X1 U15522 ( .B1(n13352), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13346), 
        .ZN(n13347) );
  OAI21_X1 U15523 ( .B1(n13348), .B2(n13357), .A(n13347), .ZN(P2_U3296) );
  INV_X1 U15524 ( .A(n13349), .ZN(n14303) );
  OAI222_X1 U15525 ( .A1(P2_U3088), .A2(n7279), .B1(n13367), .B2(n14303), .C1(
        n13350), .C2(n13372), .ZN(P2_U3298) );
  AOI21_X1 U15526 ( .B1(n13352), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13351), 
        .ZN(n13353) );
  OAI21_X1 U15527 ( .B1(n13354), .B2(n13357), .A(n13353), .ZN(P2_U3299) );
  INV_X1 U15528 ( .A(n13355), .ZN(n14305) );
  OAI222_X1 U15529 ( .A1(n13372), .A2(n13358), .B1(n13357), .B2(n14305), .C1(
        n13356), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U15530 ( .A(n13359), .ZN(n14308) );
  OAI222_X1 U15531 ( .A1(n13361), .A2(P2_U3088), .B1(n13367), .B2(n14308), 
        .C1(n13360), .C2(n13372), .ZN(P2_U3301) );
  INV_X1 U15532 ( .A(n13362), .ZN(n14311) );
  OAI222_X1 U15533 ( .A1(n13372), .A2(n13364), .B1(n13367), .B2(n14311), .C1(
        n13363), .C2(P2_U3088), .ZN(P2_U3302) );
  OAI222_X1 U15534 ( .A1(n13372), .A2(n13368), .B1(n13367), .B2(n13366), .C1(
        n13365), .C2(P2_U3088), .ZN(P2_U3303) );
  NAND2_X1 U15535 ( .A1(n14315), .A2(n13369), .ZN(n13371) );
  OAI211_X1 U15536 ( .C1(n13373), .C2(n13372), .A(n13371), .B(n13370), .ZN(
        P2_U3304) );
  INV_X1 U15537 ( .A(n13374), .ZN(n13375) );
  MUX2_X1 U15538 ( .A(n13375), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI22_X1 U15539 ( .A1(n13419), .A2(n14734), .B1(n13377), .B2(n13487), .ZN(
        n13983) );
  AOI22_X1 U15540 ( .A1(n14566), .A2(n13983), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13378) );
  OAI21_X1 U15541 ( .B1(n15385), .B2(n13987), .A(n13378), .ZN(n13379) );
  AOI21_X1 U15542 ( .B1(n14165), .B2(n14562), .A(n13379), .ZN(n13380) );
  XOR2_X1 U15543 ( .A(n13381), .B(n13382), .Z(n13387) );
  OAI22_X1 U15544 ( .A1(n7138), .A2(n14734), .B1(n13383), .B2(n13487), .ZN(
        n14046) );
  AOI22_X1 U15545 ( .A1(n14566), .A2(n14046), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13384) );
  OAI21_X1 U15546 ( .B1(n15385), .B2(n14050), .A(n13384), .ZN(n13385) );
  AOI21_X1 U15547 ( .B1(n14049), .B2(n14562), .A(n13385), .ZN(n13386) );
  OAI21_X1 U15548 ( .B1(n13387), .B2(n15379), .A(n13386), .ZN(P1_U3216) );
  AND2_X1 U15549 ( .A1(n13389), .A2(n13388), .ZN(n13392) );
  OAI211_X1 U15550 ( .C1(n13392), .C2(n13391), .A(n14564), .B(n13390), .ZN(
        n13398) );
  AOI22_X1 U15551 ( .A1(n14566), .A2(n13393), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13397) );
  NAND2_X1 U15552 ( .A1(n13481), .A2(n10601), .ZN(n13396) );
  NAND2_X1 U15553 ( .A1(n14562), .A2(n13394), .ZN(n13395) );
  NAND4_X1 U15554 ( .A1(n13398), .A2(n13397), .A3(n13396), .A4(n13395), .ZN(
        P1_U3218) );
  AOI21_X1 U15555 ( .B1(n13400), .B2(n13399), .A(n15379), .ZN(n13402) );
  NAND2_X1 U15556 ( .A1(n13402), .A2(n13401), .ZN(n13408) );
  NAND2_X1 U15557 ( .A1(n13780), .A2(n13479), .ZN(n13404) );
  NAND2_X1 U15558 ( .A1(n13782), .A2(n13478), .ZN(n13403) );
  NAND2_X1 U15559 ( .A1(n13404), .A2(n13403), .ZN(n14111) );
  NOR2_X1 U15560 ( .A1(n13405), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13932) );
  NOR2_X1 U15561 ( .A1(n15385), .A2(n14112), .ZN(n13406) );
  AOI211_X1 U15562 ( .C1(n14566), .C2(n14111), .A(n13932), .B(n13406), .ZN(
        n13407) );
  OAI211_X1 U15563 ( .C1(n14113), .C2(n15382), .A(n13408), .B(n13407), .ZN(
        P1_U3219) );
  AOI21_X1 U15564 ( .B1(n13410), .B2(n13409), .A(n6524), .ZN(n13416) );
  NAND2_X1 U15565 ( .A1(n13780), .A2(n13478), .ZN(n13412) );
  NAND2_X1 U15566 ( .A1(n13778), .A2(n13479), .ZN(n13411) );
  NAND2_X1 U15567 ( .A1(n13412), .A2(n13411), .ZN(n14081) );
  AOI22_X1 U15568 ( .A1(n14081), .A2(n14566), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13413) );
  OAI21_X1 U15569 ( .B1(n15385), .B2(n14084), .A(n13413), .ZN(n13414) );
  AOI21_X1 U15570 ( .B1(n14285), .B2(n14562), .A(n13414), .ZN(n13415) );
  OAI21_X1 U15571 ( .B1(n13416), .B2(n15379), .A(n13415), .ZN(P1_U3223) );
  XOR2_X1 U15572 ( .A(n13418), .B(n13417), .Z(n13425) );
  NOR2_X1 U15573 ( .A1(n15385), .A2(n14018), .ZN(n13423) );
  OR2_X1 U15574 ( .A1(n13419), .A2(n13487), .ZN(n13421) );
  NAND2_X1 U15575 ( .A1(n13776), .A2(n13478), .ZN(n13420) );
  AND2_X1 U15576 ( .A1(n13421), .A2(n13420), .ZN(n14176) );
  OAI22_X1 U15577 ( .A1(n15388), .A2(n14176), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15244), .ZN(n13422) );
  AOI211_X1 U15578 ( .C1(n14268), .C2(n14562), .A(n13423), .B(n13422), .ZN(
        n13424) );
  OAI21_X1 U15579 ( .B1(n13425), .B2(n15379), .A(n13424), .ZN(P1_U3225) );
  OAI21_X1 U15580 ( .B1(n13428), .B2(n13427), .A(n13426), .ZN(n13429) );
  NAND2_X1 U15581 ( .A1(n13429), .A2(n14564), .ZN(n13434) );
  OAI21_X1 U15582 ( .B1(n15388), .B2(n14239), .A(n13430), .ZN(n13431) );
  AOI21_X1 U15583 ( .B1(n13481), .B2(n13432), .A(n13431), .ZN(n13433) );
  OAI211_X1 U15584 ( .C1(n14241), .C2(n15382), .A(n13434), .B(n13433), .ZN(
        P1_U3226) );
  INV_X1 U15585 ( .A(n13435), .ZN(n13440) );
  AOI21_X1 U15586 ( .B1(n13437), .B2(n13439), .A(n13436), .ZN(n13438) );
  AOI21_X1 U15587 ( .B1(n13440), .B2(n13439), .A(n13438), .ZN(n13445) );
  OAI22_X1 U15588 ( .A1(n13672), .A2(n13487), .B1(n13656), .B2(n14734), .ZN(
        n14138) );
  NAND2_X1 U15589 ( .A1(n14566), .A2(n14138), .ZN(n13441) );
  OAI211_X1 U15590 ( .C1(n15385), .C2(n14140), .A(n13442), .B(n13441), .ZN(
        n13443) );
  AOI21_X1 U15591 ( .B1(n14235), .B2(n14562), .A(n13443), .ZN(n13444) );
  OAI21_X1 U15592 ( .B1(n13445), .B2(n15379), .A(n13444), .ZN(P1_U3228) );
  XOR2_X1 U15593 ( .A(n13447), .B(n13446), .Z(n13453) );
  OR2_X1 U15594 ( .A1(n13486), .A2(n13487), .ZN(n13449) );
  NAND2_X1 U15595 ( .A1(n13777), .A2(n13478), .ZN(n13448) );
  NAND2_X1 U15596 ( .A1(n13449), .A2(n13448), .ZN(n14028) );
  AOI22_X1 U15597 ( .A1(n14566), .A2(n14028), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13450) );
  OAI21_X1 U15598 ( .B1(n15385), .B2(n14037), .A(n13450), .ZN(n13451) );
  AOI21_X1 U15599 ( .B1(n14272), .B2(n14562), .A(n13451), .ZN(n13452) );
  OAI21_X1 U15600 ( .B1(n13453), .B2(n15379), .A(n13452), .ZN(P1_U3229) );
  OAI211_X1 U15601 ( .C1(n13456), .C2(n13455), .A(n13454), .B(n14564), .ZN(
        n13462) );
  INV_X1 U15602 ( .A(n13457), .ZN(n14096) );
  AND2_X1 U15603 ( .A1(n13781), .A2(n13478), .ZN(n13458) );
  AOI21_X1 U15604 ( .B1(n13779), .B2(n13479), .A(n13458), .ZN(n14092) );
  OAI22_X1 U15605 ( .A1(n14092), .A2(n15388), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13459), .ZN(n13460) );
  AOI21_X1 U15606 ( .B1(n13481), .B2(n14096), .A(n13460), .ZN(n13461) );
  OAI211_X1 U15607 ( .C1(n13684), .C2(n15382), .A(n13462), .B(n13461), .ZN(
        P1_U3233) );
  OAI21_X1 U15608 ( .B1(n13465), .B2(n13464), .A(n13463), .ZN(n13466) );
  NAND2_X1 U15609 ( .A1(n13466), .A2(n14564), .ZN(n13472) );
  INV_X1 U15610 ( .A(n14067), .ZN(n13470) );
  AND2_X1 U15611 ( .A1(n13777), .A2(n13479), .ZN(n13467) );
  AOI21_X1 U15612 ( .B1(n13779), .B2(n13478), .A(n13467), .ZN(n14196) );
  INV_X1 U15613 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13468) );
  OAI22_X1 U15614 ( .A1(n14196), .A2(n15388), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13468), .ZN(n13469) );
  AOI21_X1 U15615 ( .B1(n13481), .B2(n13470), .A(n13469), .ZN(n13471) );
  OAI211_X1 U15616 ( .C1(n15382), .C2(n14281), .A(n13472), .B(n13471), .ZN(
        P1_U3235) );
  OAI21_X1 U15617 ( .B1(n13475), .B2(n13474), .A(n13473), .ZN(n13476) );
  NAND2_X1 U15618 ( .A1(n13476), .A2(n14564), .ZN(n13483) );
  INV_X1 U15619 ( .A(n13477), .ZN(n14129) );
  AOI22_X1 U15620 ( .A1(n13781), .A2(n13479), .B1(n13478), .B2(n13783), .ZN(
        n14124) );
  NAND2_X1 U15621 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13899)
         );
  OAI21_X1 U15622 ( .B1(n15388), .B2(n14124), .A(n13899), .ZN(n13480) );
  AOI21_X1 U15623 ( .B1(n13481), .B2(n14129), .A(n13480), .ZN(n13482) );
  OAI211_X1 U15624 ( .C1(n14132), .C2(n15382), .A(n13483), .B(n13482), .ZN(
        P1_U3238) );
  OAI22_X1 U15625 ( .A1(n13488), .A2(n13487), .B1(n13486), .B2(n14734), .ZN(
        n13999) );
  AOI22_X1 U15626 ( .A1(n14566), .A2(n13999), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13489) );
  OAI21_X1 U15627 ( .B1(n15385), .B2(n14002), .A(n13489), .ZN(n13490) );
  AOI21_X1 U15628 ( .B1(n14171), .B2(n14562), .A(n13490), .ZN(n13491) );
  INV_X1 U15629 ( .A(n13492), .ZN(n13493) );
  AOI21_X1 U15630 ( .B1(n13495), .B2(n13494), .A(n13493), .ZN(n13500) );
  NAND2_X1 U15631 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14675)
         );
  NAND2_X1 U15632 ( .A1(n14566), .A2(n14247), .ZN(n13496) );
  OAI211_X1 U15633 ( .C1(n15385), .C2(n13497), .A(n14675), .B(n13496), .ZN(
        n13498) );
  AOI21_X1 U15634 ( .B1(n14248), .B2(n14562), .A(n13498), .ZN(n13499) );
  OAI21_X1 U15635 ( .B1(n13500), .B2(n15379), .A(n13499), .ZN(P1_U3241) );
  INV_X1 U15636 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14297) );
  OR2_X1 U15637 ( .A1(n13514), .A2(n14297), .ZN(n13502) );
  NAND2_X1 U15638 ( .A1(n13503), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n13509) );
  INV_X1 U15639 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n13504) );
  OR2_X1 U15640 ( .A1(n13505), .A2(n13504), .ZN(n13508) );
  INV_X1 U15641 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n15227) );
  OR2_X1 U15642 ( .A1(n13506), .A2(n15227), .ZN(n13507) );
  AND3_X1 U15643 ( .A1(n13509), .A2(n13508), .A3(n13507), .ZN(n13939) );
  XNOR2_X1 U15644 ( .A(n13936), .B(n13770), .ZN(n13758) );
  INV_X1 U15645 ( .A(n13758), .ZN(n13546) );
  INV_X1 U15646 ( .A(n13510), .ZN(n13545) );
  NAND2_X1 U15647 ( .A1(n13512), .A2(n13511), .ZN(n13516) );
  OR2_X1 U15648 ( .A1(n13514), .A2(n13513), .ZN(n13515) );
  XOR2_X1 U15649 ( .A(n13771), .B(n14155), .Z(n13544) );
  INV_X1 U15650 ( .A(n13967), .ZN(n13975) );
  INV_X1 U15651 ( .A(n14054), .ZN(n13541) );
  INV_X1 U15652 ( .A(n14724), .ZN(n13518) );
  NAND4_X1 U15653 ( .A1(n13576), .A2(n13518), .A3(n13569), .A4(n13517), .ZN(
        n13521) );
  NOR3_X1 U15654 ( .A1(n13521), .A2(n13520), .A3(n13519), .ZN(n13524) );
  AND4_X1 U15655 ( .A1(n13525), .A2(n13524), .A3(n13523), .A4(n13522), .ZN(
        n13526) );
  NAND2_X1 U15656 ( .A1(n13527), .A2(n13526), .ZN(n13528) );
  OR3_X1 U15657 ( .A1(n13530), .A2(n13529), .A3(n13528), .ZN(n13531) );
  NOR2_X1 U15658 ( .A1(n13532), .A2(n13531), .ZN(n13533) );
  AND4_X1 U15659 ( .A1(n13534), .A2(n13644), .A3(n13533), .A4(n14448), .ZN(
        n13536) );
  NAND4_X1 U15660 ( .A1(n14122), .A2(n13536), .A3(n7420), .A4(n14136), .ZN(
        n13537) );
  NOR2_X1 U15661 ( .A1(n13537), .A2(n7450), .ZN(n13538) );
  NAND4_X1 U15662 ( .A1(n13539), .A2(n14098), .A3(n13538), .A4(n14078), .ZN(
        n13540) );
  NOR4_X1 U15663 ( .A1(n14024), .A2(n14014), .A3(n13541), .A4(n13540), .ZN(
        n13542) );
  NAND4_X1 U15664 ( .A1(n13975), .A2(n13998), .A3(n13542), .A4(n13980), .ZN(
        n13543) );
  NOR4_X1 U15665 ( .A1(n13546), .A2(n13545), .A3(n13544), .A4(n13543), .ZN(
        n13547) );
  XNOR2_X1 U15666 ( .A(n13547), .B(n13929), .ZN(n13764) );
  NAND2_X1 U15667 ( .A1(n13548), .A2(n13550), .ZN(n13558) );
  INV_X1 U15668 ( .A(n13558), .ZN(n13763) );
  NAND2_X1 U15669 ( .A1(n13725), .A2(n13549), .ZN(n13728) );
  NAND2_X1 U15670 ( .A1(n13551), .A2(n13550), .ZN(n13552) );
  AND2_X4 U15671 ( .A1(n13728), .A2(n13552), .ZN(n13734) );
  NAND2_X1 U15672 ( .A1(n13936), .A2(n13734), .ZN(n13755) );
  AND2_X1 U15673 ( .A1(n13553), .A2(n9590), .ZN(n13554) );
  OR2_X1 U15674 ( .A1(n13555), .A2(n13554), .ZN(n13557) );
  NAND2_X1 U15675 ( .A1(n13557), .A2(n13556), .ZN(n13757) );
  NAND2_X1 U15676 ( .A1(n13757), .A2(n13558), .ZN(n13750) );
  AOI21_X1 U15677 ( .B1(n13751), .B2(n13770), .A(n13750), .ZN(n13559) );
  OAI21_X1 U15678 ( .B1(n13770), .B2(n13755), .A(n13559), .ZN(n13762) );
  NAND2_X1 U15679 ( .A1(n14729), .A2(n13564), .ZN(n13561) );
  NAND2_X1 U15680 ( .A1(n13561), .A2(n13560), .ZN(n13563) );
  OAI211_X1 U15681 ( .C1(n13564), .C2(n14729), .A(n13563), .B(n13562), .ZN(
        n13571) );
  OAI21_X1 U15682 ( .B1(n13565), .B2(n14728), .A(n13734), .ZN(n13568) );
  AOI21_X1 U15683 ( .B1(n13565), .B2(n14728), .A(n14751), .ZN(n13567) );
  OAI22_X1 U15684 ( .A1(n13568), .A2(n13567), .B1(n13566), .B2(n13734), .ZN(
        n13570) );
  OAI211_X1 U15685 ( .C1(n13734), .C2(n13571), .A(n13570), .B(n13569), .ZN(
        n13575) );
  MUX2_X1 U15686 ( .A(n13573), .B(n13572), .S(n13734), .Z(n13574) );
  NAND2_X1 U15687 ( .A1(n13575), .A2(n13574), .ZN(n13577) );
  NAND2_X1 U15688 ( .A1(n13577), .A2(n13576), .ZN(n13582) );
  NAND2_X1 U15689 ( .A1(n13797), .A2(n13578), .ZN(n13580) );
  NAND2_X1 U15690 ( .A1(n13582), .A2(n13581), .ZN(n13587) );
  MUX2_X1 U15691 ( .A(n13796), .B(n13583), .S(n13732), .Z(n13586) );
  NAND2_X1 U15692 ( .A1(n13587), .A2(n13586), .ZN(n13585) );
  MUX2_X1 U15693 ( .A(n13583), .B(n13796), .S(n13732), .Z(n13584) );
  NAND2_X1 U15694 ( .A1(n13585), .A2(n13584), .ZN(n13589) );
  MUX2_X1 U15695 ( .A(n13590), .B(n13795), .S(n13732), .Z(n13592) );
  MUX2_X1 U15696 ( .A(n13795), .B(n13590), .S(n13732), .Z(n13591) );
  INV_X1 U15697 ( .A(n13593), .ZN(n13794) );
  MUX2_X1 U15698 ( .A(n13794), .B(n13594), .S(n13732), .Z(n13598) );
  NAND2_X1 U15699 ( .A1(n13597), .A2(n13598), .ZN(n13596) );
  MUX2_X1 U15700 ( .A(n13594), .B(n13794), .S(n13732), .Z(n13595) );
  NAND2_X1 U15701 ( .A1(n13596), .A2(n13595), .ZN(n13602) );
  INV_X1 U15702 ( .A(n13597), .ZN(n13600) );
  INV_X1 U15703 ( .A(n13598), .ZN(n13599) );
  NAND2_X1 U15704 ( .A1(n13600), .A2(n13599), .ZN(n13601) );
  MUX2_X1 U15705 ( .A(n13603), .B(n13793), .S(n13732), .Z(n13605) );
  MUX2_X1 U15706 ( .A(n13603), .B(n13793), .S(n13734), .Z(n13604) );
  INV_X1 U15707 ( .A(n13605), .ZN(n13606) );
  MUX2_X1 U15708 ( .A(n13607), .B(n13792), .S(n13734), .Z(n13611) );
  MUX2_X1 U15709 ( .A(n13607), .B(n13792), .S(n13732), .Z(n13608) );
  NAND2_X1 U15710 ( .A1(n13609), .A2(n13608), .ZN(n13615) );
  INV_X1 U15711 ( .A(n13610), .ZN(n13613) );
  INV_X1 U15712 ( .A(n13611), .ZN(n13612) );
  NAND2_X1 U15713 ( .A1(n13613), .A2(n13612), .ZN(n13614) );
  MUX2_X1 U15714 ( .A(n13791), .B(n14693), .S(n13734), .Z(n13617) );
  MUX2_X1 U15715 ( .A(n13791), .B(n14693), .S(n13732), .Z(n13616) );
  MUX2_X1 U15716 ( .A(n13790), .B(n13618), .S(n13732), .Z(n13622) );
  MUX2_X1 U15717 ( .A(n13618), .B(n13790), .S(n13732), .Z(n13619) );
  NAND2_X1 U15718 ( .A1(n13620), .A2(n13619), .ZN(n13626) );
  INV_X1 U15719 ( .A(n13621), .ZN(n13624) );
  INV_X1 U15720 ( .A(n13622), .ZN(n13623) );
  NAND2_X1 U15721 ( .A1(n13624), .A2(n13623), .ZN(n13625) );
  MUX2_X1 U15722 ( .A(n13789), .B(n14563), .S(n13734), .Z(n13628) );
  MUX2_X1 U15723 ( .A(n13789), .B(n14563), .S(n13732), .Z(n13627) );
  INV_X1 U15724 ( .A(n13628), .ZN(n13629) );
  MUX2_X1 U15725 ( .A(n13788), .B(n14553), .S(n13732), .Z(n13632) );
  NAND2_X1 U15726 ( .A1(n13633), .A2(n13632), .ZN(n13631) );
  MUX2_X1 U15727 ( .A(n13788), .B(n14553), .S(n13734), .Z(n13630) );
  NAND2_X1 U15728 ( .A1(n13631), .A2(n13630), .ZN(n13635) );
  NAND2_X1 U15729 ( .A1(n13635), .A2(n13634), .ZN(n13641) );
  MUX2_X1 U15730 ( .A(n13787), .B(n13638), .S(n13734), .Z(n13642) );
  NAND2_X1 U15731 ( .A1(n13636), .A2(n13734), .ZN(n13637) );
  OAI21_X1 U15732 ( .B1(n13638), .B2(n13734), .A(n13637), .ZN(n13643) );
  NAND2_X1 U15733 ( .A1(n13641), .A2(n13640), .ZN(n13651) );
  NAND2_X1 U15734 ( .A1(n13652), .A2(n13645), .ZN(n13646) );
  NAND2_X1 U15735 ( .A1(n13646), .A2(n13734), .ZN(n13650) );
  NAND2_X1 U15736 ( .A1(n13653), .A2(n13647), .ZN(n13648) );
  NAND2_X1 U15737 ( .A1(n13648), .A2(n13732), .ZN(n13649) );
  MUX2_X1 U15738 ( .A(n13653), .B(n13652), .S(n13732), .Z(n13654) );
  NAND2_X1 U15739 ( .A1(n13655), .A2(n13654), .ZN(n13660) );
  MUX2_X1 U15740 ( .A(n13656), .B(n14241), .S(n13734), .Z(n13659) );
  MUX2_X1 U15741 ( .A(n13784), .B(n13657), .S(n13732), .Z(n13658) );
  NAND2_X1 U15742 ( .A1(n13660), .A2(n13659), .ZN(n13661) );
  NAND2_X1 U15743 ( .A1(n13662), .A2(n13661), .ZN(n13671) );
  INV_X1 U15744 ( .A(n13663), .ZN(n13668) );
  NAND2_X1 U15745 ( .A1(n13665), .A2(n13664), .ZN(n13670) );
  MUX2_X1 U15746 ( .A(n13783), .B(n14235), .S(n13734), .Z(n13666) );
  INV_X1 U15747 ( .A(n13666), .ZN(n13667) );
  OR2_X1 U15748 ( .A1(n14290), .A2(n13669), .ZN(n13681) );
  AND2_X1 U15749 ( .A1(n13681), .A2(n13680), .ZN(n13678) );
  NAND3_X1 U15750 ( .A1(n13671), .A2(n6491), .A3(n13670), .ZN(n13677) );
  AND2_X1 U15751 ( .A1(n13782), .A2(n13734), .ZN(n13675) );
  NAND2_X1 U15752 ( .A1(n13672), .A2(n13732), .ZN(n13673) );
  NAND2_X1 U15753 ( .A1(n14230), .A2(n13673), .ZN(n13674) );
  OAI21_X1 U15754 ( .B1(n14230), .B2(n13675), .A(n13674), .ZN(n13676) );
  NAND4_X1 U15755 ( .A1(n13679), .A2(n13678), .A3(n13677), .A4(n13676), .ZN(
        n13683) );
  MUX2_X1 U15756 ( .A(n13681), .B(n13680), .S(n13734), .Z(n13682) );
  MUX2_X1 U15757 ( .A(n13685), .B(n13684), .S(n13732), .Z(n13688) );
  MUX2_X1 U15758 ( .A(n13780), .B(n14215), .S(n13734), .Z(n13686) );
  NAND2_X1 U15759 ( .A1(n13690), .A2(n13689), .ZN(n13692) );
  MUX2_X1 U15760 ( .A(n13779), .B(n14285), .S(n13734), .Z(n13691) );
  MUX2_X1 U15761 ( .A(n13779), .B(n14285), .S(n13732), .Z(n13693) );
  MUX2_X1 U15762 ( .A(n7138), .B(n14281), .S(n13732), .Z(n13698) );
  MUX2_X1 U15763 ( .A(n7138), .B(n14281), .S(n13734), .Z(n13696) );
  INV_X1 U15764 ( .A(n13696), .ZN(n13697) );
  MUX2_X1 U15765 ( .A(n13777), .B(n14049), .S(n13734), .Z(n13700) );
  MUX2_X1 U15766 ( .A(n13777), .B(n14049), .S(n13732), .Z(n13699) );
  INV_X1 U15767 ( .A(n13700), .ZN(n13701) );
  MUX2_X1 U15768 ( .A(n13776), .B(n14272), .S(n13732), .Z(n13703) );
  MUX2_X1 U15769 ( .A(n13776), .B(n14272), .S(n13734), .Z(n13702) );
  INV_X1 U15770 ( .A(n13703), .ZN(n13704) );
  MUX2_X1 U15771 ( .A(n13775), .B(n14268), .S(n13734), .Z(n13708) );
  MUX2_X1 U15772 ( .A(n13775), .B(n14268), .S(n13732), .Z(n13705) );
  NAND2_X1 U15773 ( .A1(n13706), .A2(n13705), .ZN(n13712) );
  INV_X1 U15774 ( .A(n13707), .ZN(n13710) );
  INV_X1 U15775 ( .A(n13708), .ZN(n13709) );
  NAND2_X1 U15776 ( .A1(n13710), .A2(n13709), .ZN(n13711) );
  MUX2_X1 U15777 ( .A(n13774), .B(n14171), .S(n13732), .Z(n13714) );
  MUX2_X1 U15778 ( .A(n13774), .B(n14171), .S(n13734), .Z(n13713) );
  MUX2_X1 U15779 ( .A(n13773), .B(n14165), .S(n13734), .Z(n13719) );
  NAND2_X1 U15780 ( .A1(n13718), .A2(n13719), .ZN(n13717) );
  MUX2_X1 U15781 ( .A(n13773), .B(n14165), .S(n13732), .Z(n13716) );
  INV_X1 U15782 ( .A(n13719), .ZN(n13720) );
  MUX2_X1 U15783 ( .A(n9506), .B(n13968), .S(n13732), .Z(n13723) );
  MUX2_X1 U15784 ( .A(n9506), .B(n13968), .S(n13734), .Z(n13722) );
  OR2_X1 U15785 ( .A1(n13732), .A2(n13939), .ZN(n13726) );
  INV_X1 U15786 ( .A(n13771), .ZN(n13724) );
  AOI21_X1 U15787 ( .B1(n13726), .B2(n13725), .A(n13724), .ZN(n13727) );
  AOI21_X1 U15788 ( .B1(n14155), .B2(n13732), .A(n13727), .ZN(n13743) );
  INV_X1 U15789 ( .A(n13728), .ZN(n13729) );
  OR2_X1 U15790 ( .A1(n13729), .A2(n13770), .ZN(n13730) );
  AND2_X1 U15791 ( .A1(n13730), .A2(n13771), .ZN(n13731) );
  MUX2_X1 U15792 ( .A(n13731), .B(n14155), .S(n13734), .Z(n13741) );
  INV_X1 U15793 ( .A(n13772), .ZN(n13733) );
  MUX2_X1 U15794 ( .A(n13733), .B(n13957), .S(n13732), .Z(n13738) );
  MUX2_X1 U15795 ( .A(n13772), .B(n13735), .S(n13734), .Z(n13737) );
  AOI22_X1 U15796 ( .A1(n13743), .A2(n13741), .B1(n13738), .B2(n13737), .ZN(
        n13736) );
  INV_X1 U15797 ( .A(n13737), .ZN(n13740) );
  INV_X1 U15798 ( .A(n13738), .ZN(n13739) );
  NAND2_X1 U15799 ( .A1(n13740), .A2(n13739), .ZN(n13742) );
  NAND2_X1 U15800 ( .A1(n13743), .A2(n13742), .ZN(n13747) );
  INV_X1 U15801 ( .A(n13741), .ZN(n13746) );
  INV_X1 U15802 ( .A(n13742), .ZN(n13745) );
  INV_X1 U15803 ( .A(n13743), .ZN(n13744) );
  AOI22_X1 U15804 ( .A1(n13747), .A2(n13746), .B1(n13745), .B2(n13744), .ZN(
        n13748) );
  NAND2_X1 U15805 ( .A1(n13749), .A2(n13748), .ZN(n13761) );
  NOR3_X1 U15806 ( .A1(n14257), .A2(n13770), .A3(n13750), .ZN(n13756) );
  NOR3_X1 U15807 ( .A1(n13755), .A2(n13770), .A3(n13757), .ZN(n13754) );
  NOR3_X1 U15808 ( .A1(n13752), .A2(n13939), .A3(n13936), .ZN(n13753) );
  NAND3_X1 U15809 ( .A1(n13761), .A2(n7592), .A3(n13758), .ZN(n13759) );
  NOR4_X1 U15810 ( .A1(n13766), .A2(n14734), .A3(n13765), .A4(n14617), .ZN(
        n13768) );
  OAI21_X1 U15811 ( .B1(n14316), .B2(n14320), .A(P1_B_REG_SCAN_IN), .ZN(n13767) );
  OAI22_X1 U15812 ( .A1(n13769), .A2(n14316), .B1(n13768), .B2(n13767), .ZN(
        P1_U3242) );
  MUX2_X1 U15813 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13770), .S(n13814), .Z(
        P1_U3591) );
  MUX2_X1 U15814 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13771), .S(n13814), .Z(
        P1_U3590) );
  MUX2_X1 U15815 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13772), .S(n13814), .Z(
        P1_U3589) );
  MUX2_X1 U15816 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9506), .S(n13814), .Z(
        P1_U3588) );
  MUX2_X1 U15817 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13773), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15818 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13774), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15819 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13775), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15820 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13776), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15821 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13777), .S(n13814), .Z(
        P1_U3583) );
  MUX2_X1 U15822 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13778), .S(n13814), .Z(
        P1_U3582) );
  MUX2_X1 U15823 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13779), .S(n13814), .Z(
        P1_U3581) );
  MUX2_X1 U15824 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13780), .S(n13814), .Z(
        P1_U3580) );
  MUX2_X1 U15825 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13781), .S(n13814), .Z(
        P1_U3579) );
  MUX2_X1 U15826 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13782), .S(n13814), .Z(
        P1_U3578) );
  MUX2_X1 U15827 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13783), .S(n13814), .Z(
        P1_U3577) );
  MUX2_X1 U15828 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13784), .S(n13814), .Z(
        P1_U3576) );
  MUX2_X1 U15829 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13785), .S(n13814), .Z(
        P1_U3575) );
  MUX2_X1 U15830 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13786), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15831 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13787), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15832 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13788), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15833 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13789), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15834 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13790), .S(n13814), .Z(
        P1_U3570) );
  MUX2_X1 U15835 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13791), .S(n13814), .Z(
        P1_U3569) );
  MUX2_X1 U15836 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13792), .S(n13814), .Z(
        P1_U3568) );
  MUX2_X1 U15837 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13793), .S(n13814), .Z(
        P1_U3567) );
  MUX2_X1 U15838 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13794), .S(n13814), .Z(
        P1_U3566) );
  MUX2_X1 U15839 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13795), .S(n13814), .Z(
        P1_U3565) );
  MUX2_X1 U15840 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13796), .S(n13814), .Z(
        P1_U3564) );
  MUX2_X1 U15841 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13797), .S(n13814), .Z(
        P1_U3563) );
  MUX2_X1 U15842 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13798), .S(n13814), .Z(
        P1_U3562) );
  MUX2_X1 U15843 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14728), .S(n13814), .Z(
        P1_U3561) );
  MUX2_X1 U15844 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14729), .S(n13814), .Z(
        P1_U3560) );
  OAI211_X1 U15845 ( .C1(n13802), .C2(n13801), .A(n14666), .B(n13800), .ZN(
        n13809) );
  NAND2_X1 U15846 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13811) );
  OAI211_X1 U15847 ( .C1(n9811), .C2(n13804), .A(n14656), .B(n13803), .ZN(
        n13808) );
  AOI22_X1 U15848 ( .A1(n14624), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n13807) );
  NAND2_X1 U15849 ( .A1(n14669), .A2(n13805), .ZN(n13806) );
  NAND4_X1 U15850 ( .A1(n13809), .A2(n13808), .A3(n13807), .A4(n13806), .ZN(
        P1_U3244) );
  MUX2_X1 U15851 ( .A(n13812), .B(n13811), .S(n13810), .Z(n13816) );
  NOR2_X1 U15852 ( .A1(n14617), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n13813) );
  OR2_X1 U15853 ( .A1(n13815), .A2(n13813), .ZN(n14615) );
  INV_X1 U15854 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14619) );
  NAND2_X1 U15855 ( .A1(n14615), .A2(n14619), .ZN(n14622) );
  OAI211_X1 U15856 ( .C1(n13816), .C2(n13815), .A(n13814), .B(n14622), .ZN(
        n14640) );
  NAND2_X1 U15857 ( .A1(n14624), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n13818) );
  NAND2_X1 U15858 ( .A1(P1_U3086), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n13817) );
  OAI211_X1 U15859 ( .C1(n13924), .C2(n13819), .A(n13818), .B(n13817), .ZN(
        n13820) );
  INV_X1 U15860 ( .A(n13820), .ZN(n13828) );
  OAI211_X1 U15861 ( .C1(n13823), .C2(n13822), .A(n14666), .B(n13821), .ZN(
        n13827) );
  OAI211_X1 U15862 ( .C1(n13825), .C2(n13824), .A(n14656), .B(n13837), .ZN(
        n13826) );
  NAND4_X1 U15863 ( .A1(n14640), .A2(n13828), .A3(n13827), .A4(n13826), .ZN(
        P1_U3245) );
  NOR2_X1 U15864 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10601), .ZN(n13830) );
  NOR2_X1 U15865 ( .A1(n13924), .A2(n13834), .ZN(n13829) );
  AOI211_X1 U15866 ( .C1(n14624), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n13830), .B(
        n13829), .ZN(n13841) );
  OAI211_X1 U15867 ( .C1(n13833), .C2(n13832), .A(n14666), .B(n13831), .ZN(
        n13840) );
  MUX2_X1 U15868 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9813), .S(n13834), .Z(
        n13835) );
  NAND3_X1 U15869 ( .A1(n13837), .A2(n13836), .A3(n13835), .ZN(n13838) );
  NAND3_X1 U15870 ( .A1(n14656), .A2(n14629), .A3(n13838), .ZN(n13839) );
  NAND3_X1 U15871 ( .A1(n13841), .A2(n13840), .A3(n13839), .ZN(P1_U3246) );
  NOR2_X1 U15872 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13842), .ZN(n13845) );
  NOR2_X1 U15873 ( .A1(n13924), .A2(n13843), .ZN(n13844) );
  AOI211_X1 U15874 ( .C1(n14624), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n13845), .B(
        n13844), .ZN(n13855) );
  OAI211_X1 U15875 ( .C1(n13848), .C2(n13847), .A(n14666), .B(n13846), .ZN(
        n13854) );
  OR3_X1 U15876 ( .A1(n13851), .A2(n13850), .A3(n13849), .ZN(n13852) );
  NAND3_X1 U15877 ( .A1(n14656), .A2(n13865), .A3(n13852), .ZN(n13853) );
  NAND3_X1 U15878 ( .A1(n13855), .A2(n13854), .A3(n13853), .ZN(P1_U3249) );
  NOR2_X1 U15879 ( .A1(n13924), .A2(n13856), .ZN(n13857) );
  AOI211_X1 U15880 ( .C1(n14624), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n13858), .B(
        n13857), .ZN(n13870) );
  OAI211_X1 U15881 ( .C1(n13861), .C2(n13860), .A(n14666), .B(n13859), .ZN(
        n13869) );
  INV_X1 U15882 ( .A(n13862), .ZN(n13867) );
  NAND3_X1 U15883 ( .A1(n13865), .A2(n13864), .A3(n13863), .ZN(n13866) );
  NAND3_X1 U15884 ( .A1(n14656), .A2(n13867), .A3(n13866), .ZN(n13868) );
  NAND3_X1 U15885 ( .A1(n13870), .A2(n13869), .A3(n13868), .ZN(P1_U3250) );
  OAI211_X1 U15886 ( .C1(n13873), .C2(n13872), .A(n13871), .B(n14666), .ZN(
        n13885) );
  INV_X1 U15887 ( .A(n13874), .ZN(n13877) );
  NOR2_X1 U15888 ( .A1(n13924), .A2(n13875), .ZN(n13876) );
  AOI211_X1 U15889 ( .C1(n14624), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n13877), 
        .B(n13876), .ZN(n13884) );
  OR3_X1 U15890 ( .A1(n13880), .A2(n13879), .A3(n13878), .ZN(n13881) );
  NAND3_X1 U15891 ( .A1(n13882), .A2(n14656), .A3(n13881), .ZN(n13883) );
  NAND3_X1 U15892 ( .A1(n13885), .A2(n13884), .A3(n13883), .ZN(P1_U3253) );
  OAI21_X1 U15893 ( .B1(n13888), .B2(n13887), .A(n13886), .ZN(n13889) );
  NAND2_X1 U15894 ( .A1(n13889), .A2(n14666), .ZN(n13898) );
  INV_X1 U15895 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n15386) );
  NOR2_X1 U15896 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n15386), .ZN(n13890) );
  AOI21_X1 U15897 ( .B1(n14624), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n13890), 
        .ZN(n13897) );
  OAI211_X1 U15898 ( .C1(n13893), .C2(n13892), .A(n14656), .B(n13891), .ZN(
        n13896) );
  NAND2_X1 U15899 ( .A1(n14669), .A2(n13894), .ZN(n13895) );
  NAND4_X1 U15900 ( .A1(n13898), .A2(n13897), .A3(n13896), .A4(n13895), .ZN(
        P1_U3257) );
  INV_X1 U15901 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n13900) );
  OAI21_X1 U15902 ( .B1(n14677), .B2(n13900), .A(n13899), .ZN(n13901) );
  AOI21_X1 U15903 ( .B1(n13920), .B2(n14669), .A(n13901), .ZN(n13913) );
  OAI21_X1 U15904 ( .B1(n14144), .B2(n13903), .A(n13902), .ZN(n13919) );
  XNOR2_X1 U15905 ( .A(n13914), .B(n13919), .ZN(n13904) );
  NAND2_X1 U15906 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n13904), .ZN(n13921) );
  OAI211_X1 U15907 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n13904), .A(n14656), 
        .B(n13921), .ZN(n13912) );
  AOI21_X1 U15908 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n13906), .A(n13905), 
        .ZN(n13915) );
  XNOR2_X1 U15909 ( .A(n13914), .B(n13915), .ZN(n13907) );
  INV_X1 U15910 ( .A(n13907), .ZN(n13910) );
  NOR2_X1 U15911 ( .A1(n13908), .A2(n13907), .ZN(n13917) );
  INV_X1 U15912 ( .A(n13917), .ZN(n13909) );
  OAI211_X1 U15913 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n13910), .A(n14666), 
        .B(n13909), .ZN(n13911) );
  NAND3_X1 U15914 ( .A1(n13913), .A2(n13912), .A3(n13911), .ZN(P1_U3261) );
  NOR2_X1 U15915 ( .A1(n13915), .A2(n13914), .ZN(n13916) );
  NOR2_X1 U15916 ( .A1(n13917), .A2(n13916), .ZN(n13918) );
  XNOR2_X1 U15917 ( .A(n13918), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n13928) );
  INV_X1 U15918 ( .A(n13928), .ZN(n13926) );
  NAND2_X1 U15919 ( .A1(n13920), .A2(n13919), .ZN(n13922) );
  NAND2_X1 U15920 ( .A1(n13922), .A2(n13921), .ZN(n13923) );
  XOR2_X1 U15921 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n13923), .Z(n13927) );
  OAI21_X1 U15922 ( .B1(n13927), .B2(n14672), .A(n13924), .ZN(n13925) );
  AOI21_X1 U15923 ( .B1(n13926), .B2(n14666), .A(n13925), .ZN(n13931) );
  AOI22_X1 U15924 ( .A1(n13928), .A2(n14666), .B1(n14656), .B2(n13927), .ZN(
        n13930) );
  MUX2_X1 U15925 ( .A(n13931), .B(n13930), .S(n13929), .Z(n13934) );
  INV_X1 U15926 ( .A(n13932), .ZN(n13933) );
  OAI211_X1 U15927 ( .C1(n13935), .C2(n14677), .A(n13934), .B(n13933), .ZN(
        P1_U3262) );
  XNOR2_X1 U15928 ( .A(n13944), .B(n13936), .ZN(n14150) );
  NAND2_X1 U15929 ( .A1(n14150), .A2(n13986), .ZN(n13941) );
  INV_X1 U15930 ( .A(n13937), .ZN(n13938) );
  NOR2_X1 U15931 ( .A1(n13939), .A2(n13938), .ZN(n14149) );
  INV_X1 U15932 ( .A(n14149), .ZN(n14153) );
  NOR2_X1 U15933 ( .A1(n14746), .A2(n14153), .ZN(n13946) );
  AOI21_X1 U15934 ( .B1(n14710), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13946), 
        .ZN(n13940) );
  OAI211_X1 U15935 ( .C1(n14257), .C2(n14739), .A(n13941), .B(n13940), .ZN(
        P1_U3263) );
  AND2_X1 U15936 ( .A1(n14155), .A2(n13942), .ZN(n13943) );
  INV_X1 U15937 ( .A(n14155), .ZN(n14260) );
  NOR2_X1 U15938 ( .A1(n14260), .A2(n14739), .ZN(n13945) );
  AOI211_X1 U15939 ( .C1(n14710), .C2(P1_REG2_REG_30__SCAN_IN), .A(n13946), 
        .B(n13945), .ZN(n13947) );
  OAI21_X1 U15940 ( .B1(n14696), .B2(n6488), .A(n13947), .ZN(P1_U3264) );
  INV_X1 U15941 ( .A(n13948), .ZN(n13965) );
  NOR2_X1 U15942 ( .A1(n13950), .A2(n13949), .ZN(n13953) );
  INV_X1 U15943 ( .A(n13951), .ZN(n13952) );
  AOI22_X1 U15944 ( .A1(n13954), .A2(n13953), .B1(n13952), .B2(n14737), .ZN(
        n13955) );
  OAI21_X1 U15945 ( .B1(n14746), .B2(n13956), .A(n13955), .ZN(n13959) );
  NOR2_X1 U15946 ( .A1(n13957), .A2(n14739), .ZN(n13958) );
  AOI211_X1 U15947 ( .C1(n14710), .C2(P1_REG2_REG_29__SCAN_IN), .A(n13959), 
        .B(n13958), .ZN(n13960) );
  OAI21_X1 U15948 ( .B1(n13961), .B2(n14696), .A(n13960), .ZN(n13962) );
  AOI21_X1 U15949 ( .B1(n14118), .B2(n13963), .A(n13962), .ZN(n13964) );
  OAI21_X1 U15950 ( .B1(n13965), .B2(n14461), .A(n13964), .ZN(P1_U3356) );
  AOI21_X1 U15951 ( .B1(n13968), .B2(n13984), .A(n14788), .ZN(n13969) );
  NAND2_X1 U15952 ( .A1(n13969), .A2(n6479), .ZN(n14158) );
  INV_X1 U15953 ( .A(n14158), .ZN(n13974) );
  OAI22_X1 U15954 ( .A1(n14710), .A2(n14157), .B1(n13970), .B2(n14708), .ZN(
        n13971) );
  AOI21_X1 U15955 ( .B1(P1_REG2_REG_28__SCAN_IN), .B2(n14710), .A(n13971), 
        .ZN(n13972) );
  OAI21_X1 U15956 ( .B1(n14263), .B2(n14739), .A(n13972), .ZN(n13973) );
  AOI21_X1 U15957 ( .B1(n13974), .B2(n14742), .A(n13973), .ZN(n13978) );
  XNOR2_X1 U15958 ( .A(n13976), .B(n13975), .ZN(n14159) );
  NAND2_X1 U15959 ( .A1(n14159), .A2(n14118), .ZN(n13977) );
  OAI211_X1 U15960 ( .C1(n14162), .C2(n14461), .A(n13978), .B(n13977), .ZN(
        P1_U3265) );
  XNOR2_X1 U15961 ( .A(n13979), .B(n13980), .ZN(n14164) );
  NAND3_X1 U15962 ( .A1(n13996), .A2(n9554), .A3(n13981), .ZN(n13982) );
  INV_X1 U15963 ( .A(n14165), .ZN(n13991) );
  INV_X1 U15964 ( .A(n13984), .ZN(n13985) );
  AOI21_X1 U15965 ( .B1(n14165), .B2(n14006), .A(n13985), .ZN(n14166) );
  NAND2_X1 U15966 ( .A1(n14166), .A2(n13986), .ZN(n13990) );
  INV_X1 U15967 ( .A(n13987), .ZN(n13988) );
  AOI22_X1 U15968 ( .A1(n14710), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13988), 
        .B2(n14737), .ZN(n13989) );
  OAI211_X1 U15969 ( .C1(n13991), .C2(n14739), .A(n13990), .B(n13989), .ZN(
        n13992) );
  AOI21_X1 U15970 ( .B1(n14164), .B2(n14743), .A(n13992), .ZN(n13993) );
  OAI21_X1 U15971 ( .B1(n14168), .B2(n14710), .A(n13993), .ZN(P1_U3266) );
  XNOR2_X1 U15972 ( .A(n13995), .B(n13994), .ZN(n14174) );
  OAI21_X1 U15973 ( .B1(n13998), .B2(n13997), .A(n13996), .ZN(n14000) );
  AOI21_X1 U15974 ( .B1(n14000), .B2(n14730), .A(n13999), .ZN(n14173) );
  NAND2_X1 U15975 ( .A1(n14710), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n14001) );
  OAI21_X1 U15976 ( .B1(n14708), .B2(n14002), .A(n14001), .ZN(n14003) );
  AOI21_X1 U15977 ( .B1(n14171), .B2(n14694), .A(n14003), .ZN(n14009) );
  OR2_X1 U15978 ( .A1(n14005), .A2(n14004), .ZN(n14007) );
  AND3_X1 U15979 ( .A1(n14007), .A2(n14006), .A3(n14715), .ZN(n14170) );
  NAND2_X1 U15980 ( .A1(n14170), .A2(n14742), .ZN(n14008) );
  OAI211_X1 U15981 ( .C1(n14173), .C2(n14710), .A(n14009), .B(n14008), .ZN(
        n14010) );
  INV_X1 U15982 ( .A(n14010), .ZN(n14011) );
  OAI21_X1 U15983 ( .B1(n14461), .B2(n14174), .A(n14011), .ZN(P1_U3267) );
  OAI21_X1 U15984 ( .B1(n14013), .B2(n14014), .A(n14012), .ZN(n14175) );
  NAND2_X1 U15985 ( .A1(n14015), .A2(n14014), .ZN(n14016) );
  NAND2_X1 U15986 ( .A1(n14017), .A2(n14016), .ZN(n14179) );
  XNOR2_X1 U15987 ( .A(n14035), .B(n14268), .ZN(n14177) );
  OAI22_X1 U15988 ( .A1(n14710), .A2(n14176), .B1(n14018), .B2(n14708), .ZN(
        n14019) );
  AOI21_X1 U15989 ( .B1(P1_REG2_REG_25__SCAN_IN), .B2(n14710), .A(n14019), 
        .ZN(n14021) );
  NAND2_X1 U15990 ( .A1(n14268), .A2(n14694), .ZN(n14020) );
  OAI211_X1 U15991 ( .C1(n14177), .C2(n14460), .A(n14021), .B(n14020), .ZN(
        n14022) );
  AOI21_X1 U15992 ( .B1(n14179), .B2(n14118), .A(n14022), .ZN(n14023) );
  OAI21_X1 U15993 ( .B1(n14175), .B2(n14461), .A(n14023), .ZN(P1_U3268) );
  NAND2_X1 U15994 ( .A1(n14025), .A2(n14024), .ZN(n14026) );
  NAND3_X1 U15995 ( .A1(n14027), .A2(n14730), .A3(n14026), .ZN(n14030) );
  INV_X1 U15996 ( .A(n14028), .ZN(n14029) );
  AND2_X1 U15997 ( .A1(n14030), .A2(n14029), .ZN(n14187) );
  NAND2_X1 U15998 ( .A1(n14031), .A2(n14032), .ZN(n14033) );
  NAND2_X1 U15999 ( .A1(n14034), .A2(n14033), .ZN(n14184) );
  AOI21_X1 U16000 ( .B1(n14048), .B2(n14272), .A(n14788), .ZN(n14036) );
  NAND2_X1 U16001 ( .A1(n14036), .A2(n14035), .ZN(n14185) );
  INV_X1 U16002 ( .A(n14037), .ZN(n14038) );
  AOI22_X1 U16003 ( .A1(n14746), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14038), 
        .B2(n14737), .ZN(n14040) );
  NAND2_X1 U16004 ( .A1(n14272), .A2(n14694), .ZN(n14039) );
  OAI211_X1 U16005 ( .C1(n14185), .C2(n14696), .A(n14040), .B(n14039), .ZN(
        n14041) );
  AOI21_X1 U16006 ( .B1(n14184), .B2(n14042), .A(n14041), .ZN(n14043) );
  OAI21_X1 U16007 ( .B1(n14187), .B2(n14710), .A(n14043), .ZN(P1_U3269) );
  OAI21_X1 U16008 ( .B1(n14045), .B2(n14054), .A(n14044), .ZN(n14047) );
  AOI21_X1 U16009 ( .B1(n14047), .B2(n14730), .A(n14046), .ZN(n14190) );
  AOI211_X1 U16010 ( .C1(n14049), .C2(n14066), .A(n14788), .B(n7159), .ZN(
        n14192) );
  INV_X1 U16011 ( .A(n14049), .ZN(n14277) );
  NOR2_X1 U16012 ( .A1(n14277), .A2(n14739), .ZN(n14053) );
  OAI22_X1 U16013 ( .A1(n14691), .A2(n14051), .B1(n14050), .B2(n14708), .ZN(
        n14052) );
  AOI211_X1 U16014 ( .C1(n14192), .C2(n14742), .A(n14053), .B(n14052), .ZN(
        n14059) );
  NAND2_X1 U16015 ( .A1(n14055), .A2(n14054), .ZN(n14056) );
  AND2_X1 U16016 ( .A1(n14057), .A2(n14056), .ZN(n14193) );
  NAND2_X1 U16017 ( .A1(n14193), .A2(n14578), .ZN(n14058) );
  OAI211_X1 U16018 ( .C1(n14746), .C2(n14190), .A(n14059), .B(n14058), .ZN(
        P1_U3270) );
  XNOR2_X1 U16019 ( .A(n14060), .B(n14061), .ZN(n14200) );
  OR2_X1 U16020 ( .A1(n14062), .A2(n14061), .ZN(n14063) );
  NAND2_X1 U16021 ( .A1(n14064), .A2(n14063), .ZN(n14199) );
  OR2_X1 U16022 ( .A1(n14281), .A2(n14077), .ZN(n14065) );
  NAND2_X1 U16023 ( .A1(n14066), .A2(n14065), .ZN(n14197) );
  OAI22_X1 U16024 ( .A1(n14196), .A2(n14710), .B1(n14067), .B2(n14708), .ZN(
        n14069) );
  NOR2_X1 U16025 ( .A1(n14281), .A2(n14739), .ZN(n14068) );
  AOI211_X1 U16026 ( .C1(n14710), .C2(P1_REG2_REG_22__SCAN_IN), .A(n14069), 
        .B(n14068), .ZN(n14070) );
  OAI21_X1 U16027 ( .B1(n14460), .B2(n14197), .A(n14070), .ZN(n14071) );
  AOI21_X1 U16028 ( .B1(n14578), .B2(n14199), .A(n14071), .ZN(n14072) );
  OAI21_X1 U16029 ( .B1(n14200), .B2(n14073), .A(n14072), .ZN(P1_U3271) );
  XNOR2_X1 U16030 ( .A(n14074), .B(n14078), .ZN(n14206) );
  INV_X1 U16031 ( .A(n14206), .ZN(n14089) );
  NAND2_X1 U16032 ( .A1(n14285), .A2(n14094), .ZN(n14075) );
  NAND2_X1 U16033 ( .A1(n14075), .A2(n14715), .ZN(n14076) );
  OR2_X1 U16034 ( .A1(n14077), .A2(n14076), .ZN(n14208) );
  XNOR2_X1 U16035 ( .A(n14079), .B(n7443), .ZN(n14080) );
  NAND2_X1 U16036 ( .A1(n14080), .A2(n14730), .ZN(n14210) );
  INV_X1 U16037 ( .A(n14081), .ZN(n14207) );
  OAI211_X1 U16038 ( .C1(n14082), .C2(n14208), .A(n14210), .B(n14207), .ZN(
        n14083) );
  NAND2_X1 U16039 ( .A1(n14083), .A2(n14691), .ZN(n14088) );
  INV_X1 U16040 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14085) );
  OAI22_X1 U16041 ( .A1(n14691), .A2(n14085), .B1(n14084), .B2(n14708), .ZN(
        n14086) );
  AOI21_X1 U16042 ( .B1(n14285), .B2(n14694), .A(n14086), .ZN(n14087) );
  OAI211_X1 U16043 ( .C1(n14089), .C2(n14461), .A(n14088), .B(n14087), .ZN(
        P1_U3272) );
  OAI211_X1 U16044 ( .C1(n14098), .C2(n14091), .A(n14090), .B(n14730), .ZN(
        n14093) );
  INV_X1 U16045 ( .A(n14094), .ZN(n14095) );
  AOI211_X1 U16046 ( .C1(n14215), .C2(n14110), .A(n14788), .B(n14095), .ZN(
        n14214) );
  AOI22_X1 U16047 ( .A1(n14710), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14096), 
        .B2(n14737), .ZN(n14097) );
  OAI21_X1 U16048 ( .B1(n13684), .B2(n14739), .A(n14097), .ZN(n14103) );
  NAND2_X1 U16049 ( .A1(n14099), .A2(n14098), .ZN(n14100) );
  NAND2_X1 U16050 ( .A1(n14101), .A2(n14100), .ZN(n14218) );
  NOR2_X1 U16051 ( .A1(n14218), .A2(n14461), .ZN(n14102) );
  AOI211_X1 U16052 ( .C1(n14214), .C2(n14742), .A(n14103), .B(n14102), .ZN(
        n14104) );
  OAI21_X1 U16053 ( .B1(n14746), .B2(n14216), .A(n14104), .ZN(P1_U3273) );
  XNOR2_X1 U16054 ( .A(n14106), .B(n14105), .ZN(n14223) );
  INV_X1 U16055 ( .A(n14223), .ZN(n14120) );
  NAND2_X1 U16056 ( .A1(n14107), .A2(n7450), .ZN(n14108) );
  NAND2_X1 U16057 ( .A1(n14109), .A2(n14108), .ZN(n14222) );
  OAI211_X1 U16058 ( .C1(n14127), .C2(n14113), .A(n14715), .B(n14110), .ZN(
        n14220) );
  INV_X1 U16059 ( .A(n14111), .ZN(n14219) );
  OAI22_X1 U16060 ( .A1(n14219), .A2(n14710), .B1(n14112), .B2(n14708), .ZN(
        n14115) );
  NOR2_X1 U16061 ( .A1(n14113), .A2(n14739), .ZN(n14114) );
  AOI211_X1 U16062 ( .C1(n14710), .C2(P1_REG2_REG_19__SCAN_IN), .A(n14115), 
        .B(n14114), .ZN(n14116) );
  OAI21_X1 U16063 ( .B1(n14696), .B2(n14220), .A(n14116), .ZN(n14117) );
  AOI21_X1 U16064 ( .B1(n14222), .B2(n14118), .A(n14117), .ZN(n14119) );
  OAI21_X1 U16065 ( .B1(n14120), .B2(n14461), .A(n14119), .ZN(P1_U3274) );
  XNOR2_X1 U16066 ( .A(n14121), .B(n14122), .ZN(n14228) );
  XNOR2_X1 U16067 ( .A(n14123), .B(n14122), .ZN(n14125) );
  OAI21_X1 U16068 ( .B1(n14125), .B2(n14704), .A(n14124), .ZN(n14126) );
  AOI21_X1 U16069 ( .B1(n14793), .B2(n14228), .A(n14126), .ZN(n14232) );
  INV_X1 U16070 ( .A(n14142), .ZN(n14128) );
  AOI211_X1 U16071 ( .C1(n14230), .C2(n14128), .A(n14788), .B(n14127), .ZN(
        n14229) );
  NAND2_X1 U16072 ( .A1(n14229), .A2(n14742), .ZN(n14131) );
  AOI22_X1 U16073 ( .A1(n14710), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14129), 
        .B2(n14737), .ZN(n14130) );
  OAI211_X1 U16074 ( .C1(n14132), .C2(n14739), .A(n14131), .B(n14130), .ZN(
        n14133) );
  AOI21_X1 U16075 ( .B1(n14743), .B2(n14228), .A(n14133), .ZN(n14134) );
  OAI21_X1 U16076 ( .B1(n14232), .B2(n14710), .A(n14134), .ZN(P1_U3275) );
  XNOR2_X1 U16077 ( .A(n14135), .B(n14136), .ZN(n14238) );
  XNOR2_X1 U16078 ( .A(n14137), .B(n14136), .ZN(n14139) );
  AOI21_X1 U16079 ( .B1(n14139), .B2(n14730), .A(n14138), .ZN(n14236) );
  OAI21_X1 U16080 ( .B1(n14140), .B2(n14708), .A(n14236), .ZN(n14141) );
  NAND2_X1 U16081 ( .A1(n14141), .A2(n14691), .ZN(n14148) );
  AOI211_X1 U16082 ( .C1(n14235), .C2(n14143), .A(n14788), .B(n14142), .ZN(
        n14234) );
  INV_X1 U16083 ( .A(n14235), .ZN(n14145) );
  OAI22_X1 U16084 ( .A1(n14145), .A2(n14739), .B1(n14144), .B2(n14691), .ZN(
        n14146) );
  AOI21_X1 U16085 ( .B1(n14234), .B2(n14742), .A(n14146), .ZN(n14147) );
  OAI211_X1 U16086 ( .C1(n14238), .C2(n14461), .A(n14148), .B(n14147), .ZN(
        P1_U3276) );
  INV_X1 U16087 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14151) );
  AOI21_X1 U16088 ( .B1(n14150), .B2(n14715), .A(n14149), .ZN(n14255) );
  MUX2_X1 U16089 ( .A(n14151), .B(n14255), .S(n14822), .Z(n14152) );
  OAI21_X1 U16090 ( .B1(n14257), .B2(n14205), .A(n14152), .ZN(P1_U3559) );
  AOI21_X1 U16091 ( .B1(n9609), .B2(n14155), .A(n14154), .ZN(n14156) );
  INV_X1 U16092 ( .A(n14156), .ZN(P1_U3558) );
  AND2_X1 U16093 ( .A1(n14158), .A2(n14157), .ZN(n14161) );
  NAND2_X1 U16094 ( .A1(n14159), .A2(n14730), .ZN(n14160) );
  OAI211_X1 U16095 ( .C1(n14162), .C2(n14762), .A(n14161), .B(n14160), .ZN(
        n14261) );
  OAI21_X1 U16096 ( .B1(n14263), .B2(n14205), .A(n14163), .ZN(P1_U3556) );
  INV_X1 U16097 ( .A(n14164), .ZN(n14169) );
  AOI22_X1 U16098 ( .A1(n14166), .A2(n14715), .B1(n14758), .B2(n14165), .ZN(
        n14167) );
  OAI211_X1 U16099 ( .C1(n14169), .C2(n14789), .A(n14168), .B(n14167), .ZN(
        n14264) );
  MUX2_X1 U16100 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14264), .S(n14822), .Z(
        P1_U3555) );
  AOI21_X1 U16101 ( .B1(n14758), .B2(n14171), .A(n14170), .ZN(n14172) );
  OAI211_X1 U16102 ( .C1(n14174), .C2(n14762), .A(n14173), .B(n14172), .ZN(
        n14265) );
  MUX2_X1 U16103 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14265), .S(n14822), .Z(
        P1_U3554) );
  OR2_X1 U16104 ( .A1(n14175), .A2(n14762), .ZN(n14181) );
  OAI21_X1 U16105 ( .B1(n14177), .B2(n14788), .A(n14176), .ZN(n14178) );
  AOI21_X1 U16106 ( .B1(n14179), .B2(n14730), .A(n14178), .ZN(n14180) );
  NAND2_X1 U16107 ( .A1(n14181), .A2(n14180), .ZN(n14266) );
  MUX2_X1 U16108 ( .A(n14266), .B(P1_REG1_REG_25__SCAN_IN), .S(n9605), .Z(
        n14182) );
  AOI21_X1 U16109 ( .B1(n9609), .B2(n14268), .A(n14182), .ZN(n14183) );
  INV_X1 U16110 ( .A(n14183), .ZN(P1_U3553) );
  NAND2_X1 U16111 ( .A1(n14184), .A2(n14807), .ZN(n14186) );
  NAND3_X1 U16112 ( .A1(n14187), .A2(n14186), .A3(n14185), .ZN(n14270) );
  MUX2_X1 U16113 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14270), .S(n14822), .Z(
        n14188) );
  AOI21_X1 U16114 ( .B1(n9609), .B2(n14272), .A(n14188), .ZN(n14189) );
  INV_X1 U16115 ( .A(n14189), .ZN(P1_U3552) );
  INV_X1 U16116 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n14194) );
  INV_X1 U16117 ( .A(n14190), .ZN(n14191) );
  AOI211_X1 U16118 ( .C1(n14193), .C2(n14807), .A(n14192), .B(n14191), .ZN(
        n14274) );
  MUX2_X1 U16119 ( .A(n14194), .B(n14274), .S(n14822), .Z(n14195) );
  OAI21_X1 U16120 ( .B1(n14277), .B2(n14205), .A(n14195), .ZN(P1_U3551) );
  OAI21_X1 U16121 ( .B1(n14197), .B2(n14788), .A(n14196), .ZN(n14198) );
  AOI21_X1 U16122 ( .B1(n14199), .B2(n14807), .A(n14198), .ZN(n14202) );
  OR2_X1 U16123 ( .A1(n14200), .A2(n14704), .ZN(n14201) );
  NAND2_X1 U16124 ( .A1(n14202), .A2(n14201), .ZN(n14278) );
  MUX2_X1 U16125 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14278), .S(n14822), .Z(
        n14203) );
  INV_X1 U16126 ( .A(n14203), .ZN(n14204) );
  OAI21_X1 U16127 ( .B1(n14205), .B2(n14281), .A(n14204), .ZN(P1_U3550) );
  NAND2_X1 U16128 ( .A1(n14206), .A2(n14807), .ZN(n14211) );
  AND2_X1 U16129 ( .A1(n14208), .A2(n14207), .ZN(n14209) );
  NAND3_X1 U16130 ( .A1(n14211), .A2(n14210), .A3(n14209), .ZN(n14283) );
  MUX2_X1 U16131 ( .A(n14283), .B(P1_REG1_REG_21__SCAN_IN), .S(n9605), .Z(
        n14212) );
  AOI21_X1 U16132 ( .B1(n9609), .B2(n14285), .A(n14212), .ZN(n14213) );
  INV_X1 U16133 ( .A(n14213), .ZN(P1_U3549) );
  AOI21_X1 U16134 ( .B1(n14758), .B2(n14215), .A(n14214), .ZN(n14217) );
  OAI211_X1 U16135 ( .C1(n14762), .C2(n14218), .A(n14217), .B(n14216), .ZN(
        n14287) );
  MUX2_X1 U16136 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14287), .S(n14822), .Z(
        P1_U3548) );
  NAND2_X1 U16137 ( .A1(n14220), .A2(n14219), .ZN(n14221) );
  AOI21_X1 U16138 ( .B1(n14222), .B2(n14730), .A(n14221), .ZN(n14225) );
  NAND2_X1 U16139 ( .A1(n14223), .A2(n14807), .ZN(n14224) );
  NAND2_X1 U16140 ( .A1(n14225), .A2(n14224), .ZN(n14288) );
  MUX2_X1 U16141 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14288), .S(n14822), .Z(
        n14226) );
  AOI21_X1 U16142 ( .B1(n9609), .B2(n14290), .A(n14226), .ZN(n14227) );
  INV_X1 U16143 ( .A(n14227), .ZN(P1_U3547) );
  INV_X1 U16144 ( .A(n14228), .ZN(n14233) );
  AOI21_X1 U16145 ( .B1(n14758), .B2(n14230), .A(n14229), .ZN(n14231) );
  OAI211_X1 U16146 ( .C1(n14789), .C2(n14233), .A(n14232), .B(n14231), .ZN(
        n14292) );
  MUX2_X1 U16147 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14292), .S(n14822), .Z(
        P1_U3546) );
  AOI21_X1 U16148 ( .B1(n14758), .B2(n14235), .A(n14234), .ZN(n14237) );
  OAI211_X1 U16149 ( .C1(n14762), .C2(n14238), .A(n14237), .B(n14236), .ZN(
        n14293) );
  MUX2_X1 U16150 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14293), .S(n14822), .Z(
        P1_U3545) );
  OAI211_X1 U16151 ( .C1(n14241), .C2(n14796), .A(n14240), .B(n14239), .ZN(
        n14242) );
  AOI21_X1 U16152 ( .B1(n14243), .B2(n14807), .A(n14242), .ZN(n14244) );
  OAI21_X1 U16153 ( .B1(n14245), .B2(n14704), .A(n14244), .ZN(n14294) );
  MUX2_X1 U16154 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14294), .S(n14822), .Z(
        P1_U3544) );
  NAND2_X1 U16155 ( .A1(n14246), .A2(n14807), .ZN(n14254) );
  AOI21_X1 U16156 ( .B1(n14248), .B2(n14758), .A(n14247), .ZN(n14253) );
  NAND3_X1 U16157 ( .A1(n14250), .A2(n14249), .A3(n14730), .ZN(n14252) );
  NAND4_X1 U16158 ( .A1(n14254), .A2(n14253), .A3(n14252), .A4(n14251), .ZN(
        n14295) );
  MUX2_X1 U16159 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n14295), .S(n14822), .Z(
        P1_U3543) );
  MUX2_X1 U16160 ( .A(n15227), .B(n14255), .S(n14810), .Z(n14256) );
  OAI21_X1 U16161 ( .B1(n14257), .B2(n14282), .A(n14256), .ZN(P1_U3527) );
  OAI21_X1 U16162 ( .B1(n14263), .B2(n14282), .A(n14262), .ZN(P1_U3524) );
  MUX2_X1 U16163 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14264), .S(n14810), .Z(
        P1_U3523) );
  MUX2_X1 U16164 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14265), .S(n14810), .Z(
        P1_U3522) );
  MUX2_X1 U16165 ( .A(n14266), .B(P1_REG0_REG_25__SCAN_IN), .S(n14808), .Z(
        n14267) );
  AOI21_X1 U16166 ( .B1(n9614), .B2(n14268), .A(n14267), .ZN(n14269) );
  INV_X1 U16167 ( .A(n14269), .ZN(P1_U3521) );
  MUX2_X1 U16168 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14270), .S(n14810), .Z(
        n14271) );
  AOI21_X1 U16169 ( .B1(n9614), .B2(n14272), .A(n14271), .ZN(n14273) );
  INV_X1 U16170 ( .A(n14273), .ZN(P1_U3520) );
  MUX2_X1 U16171 ( .A(n14275), .B(n14274), .S(n14810), .Z(n14276) );
  OAI21_X1 U16172 ( .B1(n14277), .B2(n14282), .A(n14276), .ZN(P1_U3519) );
  MUX2_X1 U16173 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14278), .S(n14810), .Z(
        n14279) );
  INV_X1 U16174 ( .A(n14279), .ZN(n14280) );
  OAI21_X1 U16175 ( .B1(n14282), .B2(n14281), .A(n14280), .ZN(P1_U3518) );
  MUX2_X1 U16176 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14283), .S(n14810), .Z(
        n14284) );
  AOI21_X1 U16177 ( .B1(n9614), .B2(n14285), .A(n14284), .ZN(n14286) );
  INV_X1 U16178 ( .A(n14286), .ZN(P1_U3517) );
  MUX2_X1 U16179 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14287), .S(n14810), .Z(
        P1_U3516) );
  MUX2_X1 U16180 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14288), .S(n14810), .Z(
        n14289) );
  AOI21_X1 U16181 ( .B1(n9614), .B2(n14290), .A(n14289), .ZN(n14291) );
  INV_X1 U16182 ( .A(n14291), .ZN(P1_U3515) );
  MUX2_X1 U16183 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14292), .S(n14810), .Z(
        P1_U3513) );
  MUX2_X1 U16184 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14293), .S(n14810), .Z(
        P1_U3510) );
  MUX2_X1 U16185 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14294), .S(n14810), .Z(
        P1_U3507) );
  MUX2_X1 U16186 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n14295), .S(n14810), .Z(
        P1_U3504) );
  NAND3_X1 U16187 ( .A1(n14296), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n14298) );
  OAI22_X1 U16188 ( .A1(n14299), .A2(n14298), .B1(n14297), .B2(n14318), .ZN(
        n14300) );
  AOI21_X1 U16189 ( .B1(n13501), .B2(n14314), .A(n14300), .ZN(n14301) );
  INV_X1 U16190 ( .A(n14301), .ZN(P1_U3324) );
  OAI222_X1 U16191 ( .A1(n14318), .A2(n14304), .B1(n14312), .B2(n14303), .C1(
        n14302), .C2(P1_U3086), .ZN(P1_U3326) );
  OAI222_X1 U16192 ( .A1(n14318), .A2(n14306), .B1(P1_U3086), .B2(n14617), 
        .C1(n14312), .C2(n14305), .ZN(P1_U3328) );
  OAI222_X1 U16193 ( .A1(P1_U3086), .A2(n14309), .B1(n14312), .B2(n14308), 
        .C1(n14307), .C2(n14318), .ZN(P1_U3329) );
  OAI222_X1 U16194 ( .A1(n14318), .A2(n14313), .B1(n14312), .B2(n14311), .C1(
        P1_U3086), .C2(n14310), .ZN(P1_U3330) );
  NAND2_X1 U16195 ( .A1(n14315), .A2(n14314), .ZN(n14317) );
  OAI211_X1 U16196 ( .C1(n14319), .C2(n14318), .A(n14317), .B(n14316), .ZN(
        P1_U3332) );
  MUX2_X1 U16197 ( .A(n14321), .B(n14320), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U16198 ( .A(n14322), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NOR2_X1 U16199 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14323), .ZN(n14355) );
  INV_X1 U16200 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14483) );
  INV_X1 U16201 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14678) );
  NOR2_X1 U16202 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14678), .ZN(n14354) );
  NOR2_X1 U16203 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n14324), .ZN(n14353) );
  INV_X1 U16204 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14351) );
  XNOR2_X1 U16205 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(n14660), .ZN(n14363) );
  INV_X1 U16206 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14348) );
  XNOR2_X1 U16207 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n14403) );
  INV_X1 U16208 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14344) );
  XNOR2_X1 U16209 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(n14344), .ZN(n14367) );
  INV_X1 U16210 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14342) );
  XNOR2_X1 U16211 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n14394) );
  INV_X1 U16212 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14336) );
  XNOR2_X1 U16213 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n14371) );
  NAND2_X1 U16214 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14326), .ZN(n14328) );
  NAND2_X1 U16215 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14329), .ZN(n14331) );
  NAND2_X1 U16216 ( .A1(n14368), .A2(n14644), .ZN(n14330) );
  NAND2_X1 U16217 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14332), .ZN(n14334) );
  NAND2_X1 U16218 ( .A1(n14381), .A2(n9805), .ZN(n14333) );
  INV_X1 U16219 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n14337) );
  NAND2_X1 U16220 ( .A1(n14338), .A2(n14337), .ZN(n14340) );
  XNOR2_X1 U16221 ( .A(n14338), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n14390) );
  NAND2_X1 U16222 ( .A1(n14390), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14339) );
  NAND2_X1 U16223 ( .A1(n14340), .A2(n14339), .ZN(n14395) );
  NAND2_X1 U16224 ( .A1(n14394), .A2(n14395), .ZN(n14341) );
  NOR2_X1 U16225 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14364), .ZN(n14346) );
  NAND2_X1 U16226 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14364), .ZN(n14345) );
  NAND2_X1 U16227 ( .A1(n14403), .A2(n14402), .ZN(n14347) );
  AND2_X1 U16228 ( .A1(n14351), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14350) );
  INV_X1 U16229 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14352) );
  OAI22_X1 U16230 ( .A1(n14353), .A2(n14410), .B1(P3_ADDR_REG_14__SCAN_IN), 
        .B2(n14352), .ZN(n14358) );
  OAI22_X1 U16231 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14483), .B1(n14354), 
        .B2(n14358), .ZN(n14413) );
  OAI22_X1 U16232 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n11256), .B1(n14355), 
        .B2(n14413), .ZN(n14416) );
  INV_X1 U16233 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14418) );
  NAND2_X1 U16234 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14418), .ZN(n14356) );
  OAI21_X1 U16235 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(n14418), .A(n14356), 
        .ZN(n14357) );
  XOR2_X1 U16236 ( .A(n14416), .B(n14357), .Z(n14467) );
  XNOR2_X1 U16237 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n14359) );
  XNOR2_X1 U16238 ( .A(n14359), .B(n14358), .ZN(n14608) );
  XNOR2_X1 U16239 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n14361) );
  XOR2_X1 U16240 ( .A(n14361), .B(n14360), .Z(n14408) );
  XOR2_X1 U16241 ( .A(n14363), .B(n14362), .Z(n14404) );
  XNOR2_X1 U16242 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n14365) );
  XNOR2_X1 U16243 ( .A(n14365), .B(n14364), .ZN(n14440) );
  XOR2_X1 U16244 ( .A(n14367), .B(n14366), .Z(n14399) );
  INV_X1 U16245 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14865) );
  XNOR2_X1 U16246 ( .A(n14370), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n15405) );
  XOR2_X1 U16247 ( .A(n14372), .B(n14371), .Z(n14424) );
  INV_X1 U16248 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n14378) );
  NOR2_X1 U16249 ( .A1(n14377), .A2(n14378), .ZN(n14379) );
  AOI21_X1 U16250 ( .B1(n14375), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n14374), .ZN(
        n14376) );
  INV_X1 U16251 ( .A(n14376), .ZN(n15400) );
  NAND2_X1 U16252 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15400), .ZN(n15410) );
  NOR2_X1 U16253 ( .A1(n15410), .A2(n15409), .ZN(n15408) );
  NAND2_X1 U16254 ( .A1(n14424), .A2(n14423), .ZN(n14422) );
  NAND2_X1 U16255 ( .A1(n14382), .A2(n14383), .ZN(n14384) );
  NOR2_X1 U16256 ( .A1(n14386), .A2(n14385), .ZN(n14389) );
  XNOR2_X1 U16257 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n14388) );
  XOR2_X1 U16258 ( .A(n14388), .B(n14387), .Z(n14427) );
  NOR2_X1 U16259 ( .A1(n14391), .A2(n14392), .ZN(n14393) );
  XNOR2_X1 U16260 ( .A(n14390), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15403) );
  NOR2_X1 U16261 ( .A1(n15403), .A2(n15402), .ZN(n15401) );
  XNOR2_X1 U16262 ( .A(n14395), .B(n14394), .ZN(n14397) );
  NAND2_X1 U16263 ( .A1(n14396), .A2(n14397), .ZN(n14398) );
  INV_X1 U16264 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14878) );
  NOR2_X1 U16265 ( .A1(n14399), .A2(n14400), .ZN(n14401) );
  INV_X1 U16266 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14893) );
  XNOR2_X1 U16267 ( .A(n14403), .B(n14402), .ZN(n14595) );
  NAND2_X1 U16268 ( .A1(n14404), .A2(n14405), .ZN(n14406) );
  INV_X1 U16269 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14923) );
  INV_X1 U16270 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14935) );
  XOR2_X1 U16271 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n14409) );
  XOR2_X1 U16272 ( .A(n14410), .B(n14409), .Z(n14411) );
  INV_X1 U16273 ( .A(n14604), .ZN(n14605) );
  INV_X1 U16274 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14947) );
  NAND2_X1 U16275 ( .A1(n14608), .A2(n14609), .ZN(n14607) );
  XNOR2_X1 U16276 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(P3_ADDR_REG_16__SCAN_IN), 
        .ZN(n14414) );
  XOR2_X1 U16277 ( .A(n14414), .B(n14413), .Z(n14612) );
  NAND2_X1 U16278 ( .A1(n14467), .A2(n14468), .ZN(n14466) );
  OR2_X1 U16279 ( .A1(n14418), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n14417) );
  AOI22_X1 U16280 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14418), .B1(n14417), 
        .B2(n14416), .ZN(n14471) );
  NAND2_X1 U16281 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n15272), .ZN(n14419) );
  OAI21_X1 U16282 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15272), .A(n14419), 
        .ZN(n14470) );
  XNOR2_X1 U16283 ( .A(n14471), .B(n14470), .ZN(n14474) );
  AOI21_X1 U16284 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14420) );
  OAI21_X1 U16285 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14420), 
        .ZN(U28) );
  AOI21_X1 U16286 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14421) );
  OAI21_X1 U16287 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14421), 
        .ZN(U29) );
  OAI21_X1 U16288 ( .B1(n14424), .B2(n14423), .A(n14422), .ZN(n14425) );
  XNOR2_X1 U16289 ( .A(n14425), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16290 ( .B1(n14428), .B2(n14427), .A(n14426), .ZN(SUB_1596_U57) );
  OAI21_X1 U16291 ( .B1(n14430), .B2(n14878), .A(n14429), .ZN(SUB_1596_U55) );
  AOI21_X1 U16292 ( .B1(n14893), .B2(n14432), .A(n14431), .ZN(SUB_1596_U54) );
  OAI22_X1 U16293 ( .A1(n14435), .A2(n14434), .B1(SI_22_), .B2(n14433), .ZN(
        n14436) );
  AOI21_X1 U16294 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n14437), .A(n14436), .ZN(
        P3_U3273) );
  AOI21_X1 U16295 ( .B1(n14440), .B2(n14439), .A(n14438), .ZN(n14441) );
  XOR2_X1 U16296 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14441), .Z(SUB_1596_U70)
         );
  OAI21_X1 U16297 ( .B1(n7146), .B2(n14796), .A(n14442), .ZN(n14444) );
  AOI211_X1 U16298 ( .C1(n14807), .C2(n14445), .A(n14444), .B(n14443), .ZN(
        n14446) );
  AOI22_X1 U16299 ( .A1(n14810), .A2(n14446), .B1(n9305), .B2(n14808), .ZN(
        P1_U3495) );
  AOI22_X1 U16300 ( .A1(n14822), .A2(n14446), .B1(n10729), .B2(n9605), .ZN(
        P1_U3540) );
  OAI211_X1 U16301 ( .C1(n14449), .C2(n14448), .A(n14447), .B(n14730), .ZN(
        n14451) );
  NAND2_X1 U16302 ( .A1(n14451), .A2(n14450), .ZN(n14588) );
  OAI22_X1 U16303 ( .A1(n6616), .A2(n14453), .B1(n14708), .B2(n14452), .ZN(
        n14454) );
  NOR2_X1 U16304 ( .A1(n14588), .A2(n14454), .ZN(n14465) );
  OAI21_X1 U16305 ( .B1(n14457), .B2(n14456), .A(n14455), .ZN(n14590) );
  INV_X1 U16306 ( .A(n14590), .ZN(n14462) );
  OAI21_X1 U16307 ( .B1(n6616), .B2(n6617), .A(n14459), .ZN(n14587) );
  OAI22_X1 U16308 ( .A1(n14462), .A2(n14461), .B1(n14460), .B2(n14587), .ZN(
        n14463) );
  AOI21_X1 U16309 ( .B1(n14746), .B2(P1_REG2_REG_13__SCAN_IN), .A(n14463), 
        .ZN(n14464) );
  OAI21_X1 U16310 ( .B1(n14465), .B2(n14746), .A(n14464), .ZN(P1_U3280) );
  OAI21_X1 U16311 ( .B1(n14468), .B2(n14467), .A(n14466), .ZN(n14469) );
  XNOR2_X1 U16312 ( .A(n14469), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  NOR2_X1 U16313 ( .A1(n14471), .A2(n14470), .ZN(n14472) );
  AOI21_X1 U16314 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n15272), .A(n14472), 
        .ZN(n14479) );
  XNOR2_X1 U16315 ( .A(n14476), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n14477) );
  XNOR2_X1 U16316 ( .A(n14477), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n14478) );
  AOI21_X1 U16317 ( .B1(n14482), .B2(n14481), .A(n14480), .ZN(n14497) );
  OAI22_X1 U16318 ( .A1(n15068), .A2(n14484), .B1(n14483), .B2(n15065), .ZN(
        n14494) );
  AOI21_X1 U16319 ( .B1(n14487), .B2(n14486), .A(n14485), .ZN(n14492) );
  AOI21_X1 U16320 ( .B1(n14490), .B2(n14489), .A(n14488), .ZN(n14491) );
  OAI22_X1 U16321 ( .A1(n14492), .A2(n15097), .B1(n14491), .B2(n15074), .ZN(
        n14493) );
  NOR3_X1 U16322 ( .A1(n14495), .A2(n14494), .A3(n14493), .ZN(n14496) );
  OAI21_X1 U16323 ( .B1(n14497), .B2(n15081), .A(n14496), .ZN(P3_U3197) );
  AOI22_X1 U16324 ( .A1(n14518), .A2(n14499), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n14498), .ZN(n14501) );
  NAND2_X1 U16325 ( .A1(n14501), .A2(n14500), .ZN(P3_U3203) );
  INV_X1 U16326 ( .A(n14505), .ZN(n14502) );
  XNOR2_X1 U16327 ( .A(n14503), .B(n14502), .ZN(n14520) );
  OAI211_X1 U16328 ( .C1(n14506), .C2(n14505), .A(n14504), .B(n15149), .ZN(
        n14510) );
  AOI22_X1 U16329 ( .A1(n15142), .A2(n14508), .B1(n14507), .B2(n15145), .ZN(
        n14509) );
  NAND2_X1 U16330 ( .A1(n14510), .A2(n14509), .ZN(n14523) );
  AOI21_X1 U16331 ( .B1(n14520), .B2(n14511), .A(n14523), .ZN(n14516) );
  AND2_X1 U16332 ( .A1(n14512), .A2(n15173), .ZN(n14521) );
  INV_X1 U16333 ( .A(n14513), .ZN(n14514) );
  AOI22_X1 U16334 ( .A1(n15118), .A2(n14521), .B1(n15136), .B2(n14514), .ZN(
        n14515) );
  OAI221_X1 U16335 ( .B1(n14498), .B2(n14516), .C1(n15159), .C2(n12306), .A(
        n14515), .ZN(P3_U3220) );
  AOI21_X1 U16336 ( .B1(n14518), .B2(n15173), .A(n14517), .ZN(n14535) );
  INV_X1 U16337 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14519) );
  AOI22_X1 U16338 ( .A1(n15222), .A2(n14535), .B1(n14519), .B2(n15219), .ZN(
        P3_U3489) );
  AND2_X1 U16339 ( .A1(n14520), .A2(n9066), .ZN(n14522) );
  NOR3_X1 U16340 ( .A1(n14523), .A2(n14522), .A3(n14521), .ZN(n14537) );
  AOI22_X1 U16341 ( .A1(n15222), .A2(n14537), .B1(n12305), .B2(n15219), .ZN(
        P3_U3472) );
  AOI22_X1 U16342 ( .A1(n14525), .A2(n9066), .B1(n15173), .B2(n14524), .ZN(
        n14526) );
  AND2_X1 U16343 ( .A1(n14527), .A2(n14526), .ZN(n14538) );
  AOI22_X1 U16344 ( .A1(n15222), .A2(n14538), .B1(n14528), .B2(n15219), .ZN(
        P3_U3471) );
  OAI22_X1 U16345 ( .A1(n14531), .A2(n14530), .B1(n14529), .B2(n15138), .ZN(
        n14532) );
  NOR2_X1 U16346 ( .A1(n14533), .A2(n14532), .ZN(n14540) );
  AOI22_X1 U16347 ( .A1(n15222), .A2(n14540), .B1(n8798), .B2(n15219), .ZN(
        P3_U3470) );
  AOI22_X1 U16348 ( .A1(n15206), .A2(n14535), .B1(n14534), .B2(n15205), .ZN(
        P3_U3457) );
  INV_X1 U16349 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14536) );
  AOI22_X1 U16350 ( .A1(n15206), .A2(n14537), .B1(n14536), .B2(n15205), .ZN(
        P3_U3429) );
  AOI22_X1 U16351 ( .A1(n15206), .A2(n14538), .B1(n8818), .B2(n15205), .ZN(
        P3_U3426) );
  INV_X1 U16352 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14539) );
  AOI22_X1 U16353 ( .A1(n15206), .A2(n14540), .B1(n14539), .B2(n15205), .ZN(
        P3_U3423) );
  AND2_X1 U16354 ( .A1(n14541), .A2(n15033), .ZN(n14545) );
  OAI21_X1 U16355 ( .B1(n14543), .B2(n15028), .A(n14542), .ZN(n14544) );
  NOR3_X1 U16356 ( .A1(n14546), .A2(n14545), .A3(n14544), .ZN(n14548) );
  AOI22_X1 U16357 ( .A1(n15047), .A2(n14548), .B1(n11285), .B2(n15045), .ZN(
        P2_U3511) );
  INV_X1 U16358 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14547) );
  AOI22_X1 U16359 ( .A1(n15026), .A2(n14548), .B1(n14547), .B2(n15037), .ZN(
        P2_U3466) );
  AOI21_X1 U16360 ( .B1(n14551), .B2(n14550), .A(n14549), .ZN(n14552) );
  INV_X1 U16361 ( .A(n14552), .ZN(n14554) );
  AOI222_X1 U16362 ( .A1(n14555), .A2(n14566), .B1(n14554), .B2(n14564), .C1(
        n14553), .C2(n14562), .ZN(n14556) );
  NAND2_X1 U16363 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n14658)
         );
  OAI211_X1 U16364 ( .C1(n15385), .C2(n14557), .A(n14556), .B(n14658), .ZN(
        P1_U3224) );
  AOI21_X1 U16365 ( .B1(n14560), .B2(n14559), .A(n14558), .ZN(n14561) );
  INV_X1 U16366 ( .A(n14561), .ZN(n14565) );
  AOI222_X1 U16367 ( .A1(n14567), .A2(n14566), .B1(n14565), .B2(n14564), .C1(
        n14563), .C2(n14562), .ZN(n14569) );
  OAI211_X1 U16368 ( .C1(n15385), .C2(n14571), .A(n14569), .B(n14568), .ZN(
        P1_U3236) );
  NAND2_X1 U16369 ( .A1(n14570), .A2(n14742), .ZN(n14574) );
  INV_X1 U16370 ( .A(n14571), .ZN(n14572) );
  AOI22_X1 U16371 ( .A1(n14746), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n14572), 
        .B2(n14737), .ZN(n14573) );
  OAI211_X1 U16372 ( .C1(n14575), .C2(n14739), .A(n14574), .B(n14573), .ZN(
        n14576) );
  AOI21_X1 U16373 ( .B1(n14578), .B2(n14577), .A(n14576), .ZN(n14579) );
  OAI21_X1 U16374 ( .B1(n14746), .B2(n14580), .A(n14579), .ZN(P1_U3282) );
  OAI22_X1 U16375 ( .A1(n14581), .A2(n14788), .B1(n15383), .B2(n14796), .ZN(
        n14582) );
  INV_X1 U16376 ( .A(n14582), .ZN(n14585) );
  OR2_X1 U16377 ( .A1(n14583), .A2(n14762), .ZN(n14584) );
  AOI22_X1 U16378 ( .A1(n14822), .A2(n14592), .B1(n11257), .B2(n9605), .ZN(
        P1_U3542) );
  OAI22_X1 U16379 ( .A1(n14587), .A2(n14788), .B1(n6616), .B2(n14796), .ZN(
        n14589) );
  AOI211_X1 U16380 ( .C1(n14807), .C2(n14590), .A(n14589), .B(n14588), .ZN(
        n14593) );
  AOI22_X1 U16381 ( .A1(n14822), .A2(n14593), .B1(n10727), .B2(n9605), .ZN(
        P1_U3541) );
  INV_X1 U16382 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14591) );
  AOI22_X1 U16383 ( .A1(n14810), .A2(n14592), .B1(n14591), .B2(n14808), .ZN(
        P1_U3501) );
  AOI22_X1 U16384 ( .A1(n14810), .A2(n14593), .B1(n9322), .B2(n14808), .ZN(
        P1_U3498) );
  AOI21_X1 U16385 ( .B1(n14596), .B2(n14595), .A(n14594), .ZN(n14597) );
  XOR2_X1 U16386 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n14597), .Z(SUB_1596_U69)
         );
  OAI21_X1 U16387 ( .B1(n14599), .B2(n14923), .A(n14598), .ZN(SUB_1596_U68) );
  OAI222_X1 U16388 ( .A1(n14935), .A2(n14602), .B1(n14935), .B2(n6783), .C1(
        n14601), .C2(n14600), .ZN(SUB_1596_U67) );
  OAI222_X1 U16389 ( .A1(n14947), .A2(n14606), .B1(n14947), .B2(n14605), .C1(
        n14604), .C2(n14603), .ZN(SUB_1596_U66) );
  OAI21_X1 U16390 ( .B1(n14609), .B2(n14608), .A(n14607), .ZN(n14610) );
  XNOR2_X1 U16391 ( .A(n14610), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  OAI21_X1 U16392 ( .B1(n14613), .B2(n14612), .A(n14611), .ZN(n14614) );
  XNOR2_X1 U16393 ( .A(n14614), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  INV_X1 U16394 ( .A(n14615), .ZN(n14618) );
  NAND2_X1 U16395 ( .A1(n14617), .A2(n14616), .ZN(n14620) );
  NAND2_X1 U16396 ( .A1(n14618), .A2(n14620), .ZN(n14621) );
  MUX2_X1 U16397 ( .A(n14621), .B(n14620), .S(n14619), .Z(n14623) );
  NAND2_X1 U16398 ( .A1(n14623), .A2(n14622), .ZN(n14626) );
  AOI22_X1 U16399 ( .A1(n14624), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14625) );
  OAI21_X1 U16400 ( .B1(n14627), .B2(n14626), .A(n14625), .ZN(P1_U3243) );
  MUX2_X1 U16401 ( .A(n9808), .B(P1_REG2_REG_4__SCAN_IN), .S(n14633), .Z(
        n14630) );
  NAND3_X1 U16402 ( .A1(n14630), .A2(n14629), .A3(n14628), .ZN(n14631) );
  NAND3_X1 U16403 ( .A1(n14656), .A2(n14632), .A3(n14631), .ZN(n14639) );
  NAND2_X1 U16404 ( .A1(n14669), .A2(n14633), .ZN(n14638) );
  OAI211_X1 U16405 ( .C1(n14636), .C2(n14635), .A(n14666), .B(n14634), .ZN(
        n14637) );
  AND4_X1 U16406 ( .A1(n14640), .A2(n14639), .A3(n14638), .A4(n14637), .ZN(
        n14643) );
  NAND2_X1 U16407 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n14642) );
  OAI211_X1 U16408 ( .C1(n14677), .C2(n14644), .A(n14643), .B(n14642), .ZN(
        P1_U3247) );
  OAI21_X1 U16409 ( .B1(n14647), .B2(n14646), .A(n14645), .ZN(n14657) );
  MUX2_X1 U16410 ( .A(n10729), .B(P1_REG1_REG_12__SCAN_IN), .S(n14655), .Z(
        n14650) );
  INV_X1 U16411 ( .A(n14648), .ZN(n14649) );
  NAND2_X1 U16412 ( .A1(n14650), .A2(n14649), .ZN(n14652) );
  OAI21_X1 U16413 ( .B1(n14653), .B2(n14652), .A(n14651), .ZN(n14654) );
  AOI222_X1 U16414 ( .A1(n14657), .A2(n14656), .B1(n14655), .B2(n14669), .C1(
        n14654), .C2(n14666), .ZN(n14659) );
  OAI211_X1 U16415 ( .C1(n14660), .C2(n14677), .A(n14659), .B(n14658), .ZN(
        P1_U3255) );
  AOI21_X1 U16416 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14662), .A(n14661), 
        .ZN(n14673) );
  OAI21_X1 U16417 ( .B1(n14665), .B2(n14664), .A(n14663), .ZN(n14667) );
  NAND2_X1 U16418 ( .A1(n14667), .A2(n14666), .ZN(n14671) );
  NAND2_X1 U16419 ( .A1(n14669), .A2(n14668), .ZN(n14670) );
  OAI211_X1 U16420 ( .C1(n14673), .C2(n14672), .A(n14671), .B(n14670), .ZN(
        n14674) );
  INV_X1 U16421 ( .A(n14674), .ZN(n14676) );
  OAI211_X1 U16422 ( .C1(n14678), .C2(n14677), .A(n14676), .B(n14675), .ZN(
        P1_U3258) );
  OAI21_X1 U16423 ( .B1(n14680), .B2(n14681), .A(n14679), .ZN(n14806) );
  INV_X1 U16424 ( .A(n14802), .ZN(n14685) );
  NAND2_X1 U16425 ( .A1(n14682), .A2(n14681), .ZN(n14683) );
  AOI21_X1 U16426 ( .B1(n14684), .B2(n14683), .A(n14704), .ZN(n14804) );
  AOI211_X1 U16427 ( .C1(n14793), .C2(n14806), .A(n14685), .B(n14804), .ZN(
        n14699) );
  AOI21_X1 U16428 ( .B1(n14686), .B2(n14693), .A(n14788), .ZN(n14688) );
  NAND2_X1 U16429 ( .A1(n14688), .A2(n14687), .ZN(n14803) );
  OAI22_X1 U16430 ( .A1(n14691), .A2(n14690), .B1(n14689), .B2(n14708), .ZN(
        n14692) );
  AOI21_X1 U16431 ( .B1(n14694), .B2(n14693), .A(n14692), .ZN(n14695) );
  OAI21_X1 U16432 ( .B1(n14803), .B2(n14696), .A(n14695), .ZN(n14697) );
  AOI21_X1 U16433 ( .B1(n14806), .B2(n14743), .A(n14697), .ZN(n14698) );
  OAI21_X1 U16434 ( .B1(n14746), .B2(n14699), .A(n14698), .ZN(P1_U3284) );
  XNOR2_X1 U16435 ( .A(n14700), .B(n14701), .ZN(n14783) );
  XNOR2_X1 U16436 ( .A(n14702), .B(n14701), .ZN(n14705) );
  OAI21_X1 U16437 ( .B1(n14705), .B2(n14704), .A(n14703), .ZN(n14706) );
  AOI21_X1 U16438 ( .B1(n14783), .B2(n14793), .A(n14706), .ZN(n14780) );
  NOR2_X1 U16439 ( .A1(n14708), .A2(n14707), .ZN(n14709) );
  AOI21_X1 U16440 ( .B1(n14710), .B2(P1_REG2_REG_6__SCAN_IN), .A(n14709), .ZN(
        n14711) );
  OAI21_X1 U16441 ( .B1(n14739), .B2(n14779), .A(n14711), .ZN(n14712) );
  INV_X1 U16442 ( .A(n14712), .ZN(n14720) );
  INV_X1 U16443 ( .A(n14713), .ZN(n14717) );
  INV_X1 U16444 ( .A(n14714), .ZN(n14716) );
  OAI211_X1 U16445 ( .C1(n14779), .C2(n14717), .A(n14716), .B(n14715), .ZN(
        n14778) );
  INV_X1 U16446 ( .A(n14778), .ZN(n14718) );
  AOI22_X1 U16447 ( .A1(n14783), .A2(n14743), .B1(n14742), .B2(n14718), .ZN(
        n14719) );
  OAI211_X1 U16448 ( .C1(n14746), .C2(n14780), .A(n14720), .B(n14719), .ZN(
        P1_U3287) );
  XNOR2_X1 U16449 ( .A(n14724), .B(n14721), .ZN(n14755) );
  INV_X1 U16450 ( .A(n14722), .ZN(n14736) );
  OAI21_X1 U16451 ( .B1(n14724), .B2(n14723), .A(n14730), .ZN(n14733) );
  OR2_X1 U16452 ( .A1(n14751), .A2(n14725), .ZN(n14727) );
  NAND2_X1 U16453 ( .A1(n14727), .A2(n14726), .ZN(n14741) );
  XNOR2_X1 U16454 ( .A(n14741), .B(n14728), .ZN(n14731) );
  AOI21_X1 U16455 ( .B1(n14731), .B2(n14730), .A(n14729), .ZN(n14732) );
  AOI21_X1 U16456 ( .B1(n14734), .B2(n14733), .A(n14732), .ZN(n14735) );
  AOI211_X1 U16457 ( .C1(n14793), .C2(n14755), .A(n14736), .B(n14735), .ZN(
        n14752) );
  AOI22_X1 U16458 ( .A1(n14710), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n14737), .ZN(n14738) );
  OAI21_X1 U16459 ( .B1(n14739), .B2(n14751), .A(n14738), .ZN(n14740) );
  INV_X1 U16460 ( .A(n14740), .ZN(n14745) );
  NOR2_X1 U16461 ( .A1(n14741), .A2(n14788), .ZN(n14749) );
  AOI22_X1 U16462 ( .A1(n14743), .A2(n14755), .B1(n14742), .B2(n14749), .ZN(
        n14744) );
  OAI211_X1 U16463 ( .C1(n14746), .C2(n14752), .A(n14745), .B(n14744), .ZN(
        P1_U3292) );
  AND2_X1 U16464 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14748), .ZN(P1_U3294) );
  AND2_X1 U16465 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14748), .ZN(P1_U3295) );
  AND2_X1 U16466 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14748), .ZN(P1_U3296) );
  AND2_X1 U16467 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14748), .ZN(P1_U3297) );
  AND2_X1 U16468 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14748), .ZN(P1_U3298) );
  AND2_X1 U16469 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14748), .ZN(P1_U3299) );
  AND2_X1 U16470 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14748), .ZN(P1_U3300) );
  AND2_X1 U16471 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14748), .ZN(P1_U3301) );
  AND2_X1 U16472 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14748), .ZN(P1_U3302) );
  AND2_X1 U16473 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14748), .ZN(P1_U3303) );
  AND2_X1 U16474 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14748), .ZN(P1_U3304) );
  AND2_X1 U16475 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14748), .ZN(P1_U3305) );
  AND2_X1 U16476 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14748), .ZN(P1_U3306) );
  INV_X1 U16477 ( .A(n14748), .ZN(n14747) );
  INV_X1 U16478 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15256) );
  NOR2_X1 U16479 ( .A1(n14747), .A2(n15256), .ZN(P1_U3307) );
  AND2_X1 U16480 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14748), .ZN(P1_U3308) );
  AND2_X1 U16481 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14748), .ZN(P1_U3309) );
  INV_X1 U16482 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n15290) );
  NOR2_X1 U16483 ( .A1(n14747), .A2(n15290), .ZN(P1_U3310) );
  AND2_X1 U16484 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14748), .ZN(P1_U3311) );
  AND2_X1 U16485 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14748), .ZN(P1_U3312) );
  AND2_X1 U16486 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14748), .ZN(P1_U3313) );
  AND2_X1 U16487 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14748), .ZN(P1_U3314) );
  AND2_X1 U16488 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14748), .ZN(P1_U3315) );
  AND2_X1 U16489 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14748), .ZN(P1_U3316) );
  AND2_X1 U16490 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14748), .ZN(P1_U3317) );
  INV_X1 U16491 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15316) );
  NOR2_X1 U16492 ( .A1(n14747), .A2(n15316), .ZN(P1_U3318) );
  AND2_X1 U16493 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14748), .ZN(P1_U3319) );
  AND2_X1 U16494 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14748), .ZN(P1_U3320) );
  AND2_X1 U16495 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14748), .ZN(P1_U3321) );
  AND2_X1 U16496 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14748), .ZN(P1_U3322) );
  AND2_X1 U16497 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14748), .ZN(P1_U3323) );
  INV_X1 U16498 ( .A(n14749), .ZN(n14750) );
  OAI21_X1 U16499 ( .B1(n14751), .B2(n14796), .A(n14750), .ZN(n14754) );
  INV_X1 U16500 ( .A(n14752), .ZN(n14753) );
  AOI211_X1 U16501 ( .C1(n14784), .C2(n14755), .A(n14754), .B(n14753), .ZN(
        n14812) );
  AOI22_X1 U16502 ( .A1(n14810), .A2(n14812), .B1(n9145), .B2(n14808), .ZN(
        P1_U3462) );
  AOI21_X1 U16503 ( .B1(n14758), .B2(n14757), .A(n14756), .ZN(n14760) );
  OAI211_X1 U16504 ( .C1(n14762), .C2(n14761), .A(n14760), .B(n14759), .ZN(
        n14763) );
  INV_X1 U16505 ( .A(n14763), .ZN(n14814) );
  AOI22_X1 U16506 ( .A1(n14810), .A2(n14814), .B1(n9175), .B2(n14808), .ZN(
        P1_U3465) );
  INV_X1 U16507 ( .A(n14764), .ZN(n14770) );
  INV_X1 U16508 ( .A(n14765), .ZN(n14767) );
  NAND3_X1 U16509 ( .A1(n14768), .A2(n14767), .A3(n14766), .ZN(n14769) );
  AOI21_X1 U16510 ( .B1(n14770), .B2(n14807), .A(n14769), .ZN(n14815) );
  AOI22_X1 U16511 ( .A1(n14810), .A2(n14815), .B1(n9194), .B2(n14808), .ZN(
        P1_U3471) );
  INV_X1 U16512 ( .A(n14771), .ZN(n14773) );
  NAND4_X1 U16513 ( .A1(n14775), .A2(n14774), .A3(n14773), .A4(n14772), .ZN(
        n14776) );
  AOI21_X1 U16514 ( .B1(n14777), .B2(n14807), .A(n14776), .ZN(n14816) );
  AOI22_X1 U16515 ( .A1(n14810), .A2(n14816), .B1(n9215), .B2(n14808), .ZN(
        P1_U3474) );
  OAI21_X1 U16516 ( .B1(n14779), .B2(n14796), .A(n14778), .ZN(n14782) );
  INV_X1 U16517 ( .A(n14780), .ZN(n14781) );
  AOI211_X1 U16518 ( .C1(n14784), .C2(n14783), .A(n14782), .B(n14781), .ZN(
        n14818) );
  AOI22_X1 U16519 ( .A1(n14810), .A2(n14818), .B1(n9226), .B2(n14808), .ZN(
        P1_U3477) );
  INV_X1 U16520 ( .A(n14790), .ZN(n14794) );
  OAI211_X1 U16521 ( .C1(n14788), .C2(n14787), .A(n14786), .B(n14785), .ZN(
        n14792) );
  NOR2_X1 U16522 ( .A1(n14790), .A2(n14789), .ZN(n14791) );
  AOI211_X1 U16523 ( .C1(n14794), .C2(n14793), .A(n14792), .B(n14791), .ZN(
        n14819) );
  AOI22_X1 U16524 ( .A1(n14810), .A2(n14819), .B1(n9238), .B2(n14808), .ZN(
        P1_U3480) );
  OAI21_X1 U16525 ( .B1(n14797), .B2(n14796), .A(n14795), .ZN(n14799) );
  AOI211_X1 U16526 ( .C1(n14800), .C2(n14807), .A(n14799), .B(n14798), .ZN(
        n14820) );
  AOI22_X1 U16527 ( .A1(n14810), .A2(n14820), .B1(n9251), .B2(n14808), .ZN(
        P1_U3483) );
  NAND3_X1 U16528 ( .A1(n14803), .A2(n14802), .A3(n14801), .ZN(n14805) );
  AOI211_X1 U16529 ( .C1(n14807), .C2(n14806), .A(n14805), .B(n14804), .ZN(
        n14821) );
  INV_X1 U16530 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14809) );
  AOI22_X1 U16531 ( .A1(n14810), .A2(n14821), .B1(n14809), .B2(n14808), .ZN(
        P1_U3486) );
  AOI22_X1 U16532 ( .A1(n14822), .A2(n14812), .B1(n14811), .B2(n9605), .ZN(
        P1_U3529) );
  AOI22_X1 U16533 ( .A1(n14822), .A2(n14814), .B1(n14813), .B2(n9605), .ZN(
        P1_U3530) );
  AOI22_X1 U16534 ( .A1(n14822), .A2(n14815), .B1(n9795), .B2(n9605), .ZN(
        P1_U3532) );
  AOI22_X1 U16535 ( .A1(n14822), .A2(n14816), .B1(n9828), .B2(n9605), .ZN(
        P1_U3533) );
  AOI22_X1 U16536 ( .A1(n14822), .A2(n14818), .B1(n14817), .B2(n9605), .ZN(
        P1_U3534) );
  AOI22_X1 U16537 ( .A1(n14822), .A2(n14819), .B1(n9829), .B2(n9605), .ZN(
        P1_U3535) );
  AOI22_X1 U16538 ( .A1(n14822), .A2(n14820), .B1(n9850), .B2(n9605), .ZN(
        P1_U3536) );
  AOI22_X1 U16539 ( .A1(n14822), .A2(n14821), .B1(n10139), .B2(n9605), .ZN(
        P1_U3537) );
  NOR2_X1 U16540 ( .A1(n14823), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16541 ( .A1(n14823), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n14838) );
  OAI21_X1 U16542 ( .B1(n14826), .B2(n14825), .A(n14824), .ZN(n14835) );
  NAND2_X1 U16543 ( .A1(n14971), .A2(n14827), .ZN(n14834) );
  INV_X1 U16544 ( .A(n14828), .ZN(n14830) );
  NAND2_X1 U16545 ( .A1(n14830), .A2(n14829), .ZN(n14831) );
  NAND3_X1 U16546 ( .A1(n14985), .A2(n14832), .A3(n14831), .ZN(n14833) );
  OAI211_X1 U16547 ( .C1(n14960), .C2(n14835), .A(n14834), .B(n14833), .ZN(
        n14836) );
  INV_X1 U16548 ( .A(n14836), .ZN(n14837) );
  NAND2_X1 U16549 ( .A1(n14838), .A2(n14837), .ZN(P2_U3215) );
  OAI21_X1 U16550 ( .B1(n14841), .B2(n14840), .A(n14839), .ZN(n14848) );
  OAI211_X1 U16551 ( .C1(n14844), .C2(n14843), .A(n14985), .B(n14842), .ZN(
        n14847) );
  NAND2_X1 U16552 ( .A1(n14971), .A2(n14845), .ZN(n14846) );
  OAI211_X1 U16553 ( .C1(n14960), .C2(n14848), .A(n14847), .B(n14846), .ZN(
        n14849) );
  INV_X1 U16554 ( .A(n14849), .ZN(n14851) );
  NAND2_X1 U16555 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n14850) );
  OAI211_X1 U16556 ( .C1(n14988), .C2(n6918), .A(n14851), .B(n14850), .ZN(
        P2_U3217) );
  OAI21_X1 U16557 ( .B1(n14854), .B2(n14853), .A(n14852), .ZN(n14861) );
  OAI211_X1 U16558 ( .C1(n14857), .C2(n14856), .A(n14985), .B(n14855), .ZN(
        n14860) );
  NAND2_X1 U16559 ( .A1(n14971), .A2(n14858), .ZN(n14859) );
  OAI211_X1 U16560 ( .C1(n14960), .C2(n14861), .A(n14860), .B(n14859), .ZN(
        n14862) );
  INV_X1 U16561 ( .A(n14862), .ZN(n14864) );
  OAI211_X1 U16562 ( .C1(n14988), .C2(n14865), .A(n14864), .B(n14863), .ZN(
        P2_U3218) );
  OAI211_X1 U16563 ( .C1(n14868), .C2(n14867), .A(n14866), .B(n14977), .ZN(
        n14873) );
  OAI211_X1 U16564 ( .C1(n14871), .C2(n14870), .A(n14869), .B(n14985), .ZN(
        n14872) );
  OAI211_X1 U16565 ( .C1(n14979), .C2(n14874), .A(n14873), .B(n14872), .ZN(
        n14875) );
  INV_X1 U16566 ( .A(n14875), .ZN(n14877) );
  OAI211_X1 U16567 ( .C1(n14878), .C2(n14988), .A(n14877), .B(n14876), .ZN(
        P2_U3222) );
  NAND2_X1 U16568 ( .A1(n14880), .A2(n14879), .ZN(n14881) );
  AOI21_X1 U16569 ( .B1(n14882), .B2(n14881), .A(n14960), .ZN(n14890) );
  NAND2_X1 U16570 ( .A1(n14884), .A2(n14883), .ZN(n14885) );
  AOI21_X1 U16571 ( .B1(n14886), .B2(n14885), .A(n14965), .ZN(n14889) );
  NOR2_X1 U16572 ( .A1(n14979), .A2(n14887), .ZN(n14888) );
  NOR3_X1 U16573 ( .A1(n14890), .A2(n14889), .A3(n14888), .ZN(n14892) );
  OAI211_X1 U16574 ( .C1(n14893), .C2(n14988), .A(n14892), .B(n14891), .ZN(
        P2_U3223) );
  INV_X1 U16575 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14907) );
  OAI211_X1 U16576 ( .C1(n14896), .C2(n14895), .A(n14894), .B(n14977), .ZN(
        n14897) );
  OAI21_X1 U16577 ( .B1(n14979), .B2(n14898), .A(n14897), .ZN(n14904) );
  NAND2_X1 U16578 ( .A1(n14900), .A2(n14899), .ZN(n14901) );
  AOI21_X1 U16579 ( .B1(n14902), .B2(n14901), .A(n14965), .ZN(n14903) );
  NOR2_X1 U16580 ( .A1(n14904), .A2(n14903), .ZN(n14906) );
  OAI211_X1 U16581 ( .C1(n14907), .C2(n14988), .A(n14906), .B(n14905), .ZN(
        P2_U3225) );
  INV_X1 U16582 ( .A(n14908), .ZN(n14910) );
  OAI21_X1 U16583 ( .B1(n14910), .B2(n14909), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n14911) );
  OAI21_X1 U16584 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n14911), .ZN(n14922) );
  OAI21_X1 U16585 ( .B1(n14914), .B2(n14913), .A(n14912), .ZN(n14920) );
  AOI21_X1 U16586 ( .B1(n14917), .B2(n14916), .A(n14915), .ZN(n14918) );
  NOR2_X1 U16587 ( .A1(n14918), .A2(n14960), .ZN(n14919) );
  AOI21_X1 U16588 ( .B1(n14985), .B2(n14920), .A(n14919), .ZN(n14921) );
  OAI211_X1 U16589 ( .C1(n14923), .C2(n14988), .A(n14922), .B(n14921), .ZN(
        P2_U3226) );
  AOI21_X1 U16590 ( .B1(n14925), .B2(n14924), .A(n14965), .ZN(n14932) );
  OAI21_X1 U16591 ( .B1(n14927), .B2(n14926), .A(n14977), .ZN(n14929) );
  OAI22_X1 U16592 ( .A1(n14929), .A2(n14928), .B1(n6714), .B2(n14979), .ZN(
        n14930) );
  AOI21_X1 U16593 ( .B1(n14932), .B2(n14931), .A(n14930), .ZN(n14934) );
  NAND2_X1 U16594 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n14933)
         );
  OAI211_X1 U16595 ( .C1(n14935), .C2(n14988), .A(n14934), .B(n14933), .ZN(
        P2_U3227) );
  AOI211_X1 U16596 ( .C1(n14938), .C2(n14937), .A(n14965), .B(n14936), .ZN(
        n14943) );
  AOI211_X1 U16597 ( .C1(n14941), .C2(n14940), .A(n14960), .B(n14939), .ZN(
        n14942) );
  AOI211_X1 U16598 ( .C1(n14971), .C2(n14944), .A(n14943), .B(n14942), .ZN(
        n14946) );
  NAND2_X1 U16599 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14945)
         );
  OAI211_X1 U16600 ( .C1(n14947), .C2(n14988), .A(n14946), .B(n14945), .ZN(
        P2_U3228) );
  AOI211_X1 U16601 ( .C1(n14950), .C2(n14949), .A(n14948), .B(n14965), .ZN(
        n14955) );
  AOI211_X1 U16602 ( .C1(n14953), .C2(n14952), .A(n14951), .B(n14960), .ZN(
        n14954) );
  AOI211_X1 U16603 ( .C1(n14971), .C2(n14956), .A(n14955), .B(n14954), .ZN(
        n14958) );
  NAND2_X1 U16604 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n14957)
         );
  OAI211_X1 U16605 ( .C1(n6774), .C2(n14988), .A(n14958), .B(n14957), .ZN(
        P2_U3229) );
  INV_X1 U16606 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14974) );
  AOI211_X1 U16607 ( .C1(n14962), .C2(n14961), .A(n14960), .B(n14959), .ZN(
        n14969) );
  INV_X1 U16608 ( .A(n14963), .ZN(n14964) );
  AOI211_X1 U16609 ( .C1(n14967), .C2(n14966), .A(n14965), .B(n14964), .ZN(
        n14968) );
  AOI211_X1 U16610 ( .C1(n14971), .C2(n14970), .A(n14969), .B(n14968), .ZN(
        n14973) );
  NAND2_X1 U16611 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n14972)
         );
  OAI211_X1 U16612 ( .C1(n14974), .C2(n14988), .A(n14973), .B(n14972), .ZN(
        P2_U3230) );
  INV_X1 U16613 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n14989) );
  OAI21_X1 U16614 ( .B1(n14976), .B2(n15242), .A(n14975), .ZN(n14984) );
  OAI21_X1 U16615 ( .B1(n14978), .B2(P2_REG1_REG_18__SCAN_IN), .A(n14977), 
        .ZN(n14982) );
  OAI22_X1 U16616 ( .A1(n14982), .A2(n14981), .B1(n14980), .B2(n14979), .ZN(
        n14983) );
  AOI21_X1 U16617 ( .B1(n14985), .B2(n14984), .A(n14983), .ZN(n14987) );
  OAI211_X1 U16618 ( .C1(n14989), .C2(n14988), .A(n14987), .B(n14986), .ZN(
        P2_U3232) );
  INV_X1 U16619 ( .A(n14991), .ZN(n14992) );
  AND2_X1 U16620 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14992), .ZN(P2_U3266) );
  AND2_X1 U16621 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14992), .ZN(P2_U3267) );
  AND2_X1 U16622 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14992), .ZN(P2_U3268) );
  INV_X1 U16623 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15287) );
  NOR2_X1 U16624 ( .A1(n14991), .A2(n15287), .ZN(P2_U3269) );
  AND2_X1 U16625 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14992), .ZN(P2_U3270) );
  AND2_X1 U16626 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14992), .ZN(P2_U3271) );
  AND2_X1 U16627 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14992), .ZN(P2_U3272) );
  AND2_X1 U16628 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14992), .ZN(P2_U3273) );
  AND2_X1 U16629 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14992), .ZN(P2_U3274) );
  AND2_X1 U16630 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14992), .ZN(P2_U3275) );
  AND2_X1 U16631 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14992), .ZN(P2_U3276) );
  AND2_X1 U16632 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14992), .ZN(P2_U3277) );
  AND2_X1 U16633 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14992), .ZN(P2_U3278) );
  AND2_X1 U16634 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14992), .ZN(P2_U3279) );
  AND2_X1 U16635 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14992), .ZN(P2_U3280) );
  AND2_X1 U16636 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14992), .ZN(P2_U3281) );
  AND2_X1 U16637 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14992), .ZN(P2_U3282) );
  AND2_X1 U16638 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14992), .ZN(P2_U3283) );
  AND2_X1 U16639 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14992), .ZN(P2_U3284) );
  AND2_X1 U16640 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14992), .ZN(P2_U3285) );
  AND2_X1 U16641 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14992), .ZN(P2_U3286) );
  AND2_X1 U16642 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14992), .ZN(P2_U3287) );
  AND2_X1 U16643 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14992), .ZN(P2_U3288) );
  AND2_X1 U16644 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14992), .ZN(P2_U3289) );
  AND2_X1 U16645 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14992), .ZN(P2_U3290) );
  INV_X1 U16646 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15303) );
  NOR2_X1 U16647 ( .A1(n14991), .A2(n15303), .ZN(P2_U3291) );
  AND2_X1 U16648 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14992), .ZN(P2_U3292) );
  AND2_X1 U16649 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14992), .ZN(P2_U3293) );
  AND2_X1 U16650 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14992), .ZN(P2_U3294) );
  AND2_X1 U16651 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14992), .ZN(P2_U3295) );
  AOI22_X1 U16652 ( .A1(n14998), .A2(n14994), .B1(n14993), .B2(n14995), .ZN(
        P2_U3416) );
  AOI22_X1 U16653 ( .A1(n14998), .A2(n14997), .B1(n14996), .B2(n14995), .ZN(
        P2_U3417) );
  INV_X1 U16654 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14999) );
  AOI22_X1 U16655 ( .A1(n15026), .A2(n15000), .B1(n14999), .B2(n15037), .ZN(
        P2_U3430) );
  INV_X1 U16656 ( .A(n15001), .ZN(n15002) );
  OAI22_X1 U16657 ( .A1(n15003), .A2(n15030), .B1(n15002), .B2(n15028), .ZN(
        n15004) );
  AOI21_X1 U16658 ( .B1(n15005), .B2(n15033), .A(n15004), .ZN(n15006) );
  AND2_X1 U16659 ( .A1(n15007), .A2(n15006), .ZN(n15040) );
  INV_X1 U16660 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15008) );
  AOI22_X1 U16661 ( .A1(n15026), .A2(n15040), .B1(n15008), .B2(n15037), .ZN(
        P2_U3448) );
  INV_X1 U16662 ( .A(n15009), .ZN(n15015) );
  OAI22_X1 U16663 ( .A1(n15011), .A2(n15030), .B1(n15010), .B2(n15028), .ZN(
        n15013) );
  AOI211_X1 U16664 ( .C1(n15015), .C2(n15014), .A(n15013), .B(n15012), .ZN(
        n15042) );
  INV_X1 U16665 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15016) );
  AOI22_X1 U16666 ( .A1(n15026), .A2(n15042), .B1(n15016), .B2(n15037), .ZN(
        P2_U3451) );
  AOI21_X1 U16667 ( .B1(n15019), .B2(n15018), .A(n15017), .ZN(n15020) );
  OAI211_X1 U16668 ( .C1(n15023), .C2(n15022), .A(n15021), .B(n15020), .ZN(
        n15024) );
  INV_X1 U16669 ( .A(n15024), .ZN(n15044) );
  INV_X1 U16670 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15025) );
  AOI22_X1 U16671 ( .A1(n15026), .A2(n15044), .B1(n15025), .B2(n15037), .ZN(
        P2_U3454) );
  INV_X1 U16672 ( .A(n15027), .ZN(n15029) );
  OAI22_X1 U16673 ( .A1(n15031), .A2(n15030), .B1(n15029), .B2(n15028), .ZN(
        n15032) );
  AOI21_X1 U16674 ( .B1(n15034), .B2(n15033), .A(n15032), .ZN(n15035) );
  AND2_X1 U16675 ( .A1(n15036), .A2(n15035), .ZN(n15046) );
  INV_X1 U16676 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15038) );
  AOI22_X1 U16677 ( .A1(n15026), .A2(n15046), .B1(n15038), .B2(n15037), .ZN(
        P2_U3460) );
  AOI22_X1 U16678 ( .A1(n15047), .A2(n15040), .B1(n15039), .B2(n15045), .ZN(
        P2_U3505) );
  AOI22_X1 U16679 ( .A1(n15047), .A2(n15042), .B1(n15041), .B2(n15045), .ZN(
        P2_U3506) );
  AOI22_X1 U16680 ( .A1(n15047), .A2(n15044), .B1(n15043), .B2(n15045), .ZN(
        P2_U3507) );
  AOI22_X1 U16681 ( .A1(n15047), .A2(n15046), .B1(n9884), .B2(n15045), .ZN(
        P2_U3509) );
  NOR2_X1 U16682 ( .A1(P3_U3897), .A2(n15087), .ZN(P3_U3150) );
  AOI21_X1 U16683 ( .B1(P3_ADDR_REG_7__SCAN_IN), .B2(n15087), .A(n15048), .ZN(
        n15062) );
  OAI21_X1 U16684 ( .B1(n15051), .B2(n15050), .A(n15049), .ZN(n15052) );
  AOI22_X1 U16685 ( .A1(n15084), .A2(n15053), .B1(n15100), .B2(n15052), .ZN(
        n15061) );
  OAI221_X1 U16686 ( .B1(n15055), .B2(n8730), .C1(n15055), .C2(n15054), .A(
        n15089), .ZN(n15060) );
  AOI21_X1 U16687 ( .B1(n15057), .B2(n8727), .A(n15056), .ZN(n15058) );
  OR2_X1 U16688 ( .A1(n15058), .A2(n15097), .ZN(n15059) );
  NAND4_X1 U16689 ( .A1(n15062), .A2(n15061), .A3(n15060), .A4(n15059), .ZN(
        P3_U3189) );
  AOI21_X1 U16690 ( .B1(n15064), .B2(n15063), .A(n6599), .ZN(n15082) );
  INV_X1 U16691 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n15066) );
  OAI22_X1 U16692 ( .A1(n15068), .A2(n15067), .B1(n15066), .B2(n15065), .ZN(
        n15078) );
  AOI21_X1 U16693 ( .B1(n15070), .B2(n15069), .A(n6600), .ZN(n15076) );
  AOI21_X1 U16694 ( .B1(n15073), .B2(n15072), .A(n15071), .ZN(n15075) );
  OAI22_X1 U16695 ( .A1(n15076), .A2(n15097), .B1(n15075), .B2(n15074), .ZN(
        n15077) );
  NOR3_X1 U16696 ( .A1(n15079), .A2(n15078), .A3(n15077), .ZN(n15080) );
  OAI21_X1 U16697 ( .B1(n15082), .B2(n15081), .A(n15080), .ZN(P3_U3192) );
  AND2_X1 U16698 ( .A1(n15084), .A2(n15083), .ZN(n15085) );
  AOI211_X1 U16699 ( .C1(P3_ADDR_REG_12__SCAN_IN), .C2(n15087), .A(n15086), 
        .B(n15085), .ZN(n15106) );
  INV_X1 U16700 ( .A(n15088), .ZN(n15092) );
  OAI221_X1 U16701 ( .B1(n15092), .B2(n15091), .C1(n15092), .C2(n15090), .A(
        n15089), .ZN(n15105) );
  INV_X1 U16702 ( .A(n15093), .ZN(n15094) );
  AOI21_X1 U16703 ( .B1(n15096), .B2(n15095), .A(n15094), .ZN(n15098) );
  OR2_X1 U16704 ( .A1(n15098), .A2(n15097), .ZN(n15104) );
  OAI211_X1 U16705 ( .C1(n15102), .C2(n15101), .A(n15100), .B(n15099), .ZN(
        n15103) );
  NAND4_X1 U16706 ( .A1(n15106), .A2(n15105), .A3(n15104), .A4(n15103), .ZN(
        P3_U3194) );
  XNOR2_X1 U16707 ( .A(n15107), .B(n15110), .ZN(n15114) );
  INV_X1 U16708 ( .A(n15114), .ZN(n15171) );
  AOI22_X1 U16709 ( .A1(n15142), .A2(n15144), .B1(n15108), .B2(n15145), .ZN(
        n15113) );
  OAI211_X1 U16710 ( .C1(n15111), .C2(n15110), .A(n15149), .B(n15109), .ZN(
        n15112) );
  OAI211_X1 U16711 ( .C1(n15114), .C2(n15153), .A(n15113), .B(n15112), .ZN(
        n15169) );
  AOI21_X1 U16712 ( .B1(n15115), .B2(n15171), .A(n15169), .ZN(n15120) );
  NOR2_X1 U16713 ( .A1(n15116), .A2(n15138), .ZN(n15170) );
  AOI22_X1 U16714 ( .A1(n15118), .A2(n15170), .B1(n15136), .B2(n15117), .ZN(
        n15119) );
  OAI221_X1 U16715 ( .B1(n14498), .B2(n15120), .C1(n15159), .C2(n10475), .A(
        n15119), .ZN(P3_U3230) );
  OAI21_X1 U16716 ( .B1(n15122), .B2(n7210), .A(n15121), .ZN(n15167) );
  INV_X1 U16717 ( .A(n15167), .ZN(n15134) );
  AOI22_X1 U16718 ( .A1(n15142), .A2(n15124), .B1(n15123), .B2(n15145), .ZN(
        n15130) );
  OAI21_X1 U16719 ( .B1(n15127), .B2(n15126), .A(n15125), .ZN(n15128) );
  NAND2_X1 U16720 ( .A1(n15128), .A2(n15149), .ZN(n15129) );
  OAI211_X1 U16721 ( .C1(n15134), .C2(n15153), .A(n15130), .B(n15129), .ZN(
        n15165) );
  NOR2_X1 U16722 ( .A1(n15131), .A2(n15138), .ZN(n15166) );
  INV_X1 U16723 ( .A(n15166), .ZN(n15132) );
  OAI22_X1 U16724 ( .A1(n15134), .A2(n15133), .B1(n15140), .B2(n15132), .ZN(
        n15135) );
  AOI211_X1 U16725 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15136), .A(n15165), .B(
        n15135), .ZN(n15137) );
  AOI22_X1 U16726 ( .A1(n14498), .A2(n10469), .B1(n15137), .B2(n15159), .ZN(
        P3_U3231) );
  NOR2_X1 U16727 ( .A1(n15139), .A2(n15138), .ZN(n15163) );
  XNOR2_X1 U16728 ( .A(n15148), .B(n15141), .ZN(n15161) );
  AOI22_X1 U16729 ( .A1(n15145), .A2(n15144), .B1(n15143), .B2(n15142), .ZN(
        n15152) );
  OAI21_X1 U16730 ( .B1(n15148), .B2(n15147), .A(n15146), .ZN(n15150) );
  NAND2_X1 U16731 ( .A1(n15150), .A2(n15149), .ZN(n15151) );
  OAI211_X1 U16732 ( .C1(n15161), .C2(n15153), .A(n15152), .B(n15151), .ZN(
        n15162) );
  AOI21_X1 U16733 ( .B1(n15163), .B2(n6677), .A(n15162), .ZN(n15160) );
  OAI22_X1 U16734 ( .A1(n15156), .A2(n15161), .B1(n15155), .B2(n15154), .ZN(
        n15157) );
  INV_X1 U16735 ( .A(n15157), .ZN(n15158) );
  OAI221_X1 U16736 ( .B1(n14498), .B2(n15160), .C1(n15159), .C2(n10413), .A(
        n15158), .ZN(P3_U3232) );
  INV_X1 U16737 ( .A(n15161), .ZN(n15164) );
  AOI211_X1 U16738 ( .C1(n15203), .C2(n15164), .A(n15163), .B(n15162), .ZN(
        n15207) );
  AOI22_X1 U16739 ( .A1(n15206), .A2(n15207), .B1(n7218), .B2(n15205), .ZN(
        P3_U3393) );
  AOI211_X1 U16740 ( .C1(n15203), .C2(n15167), .A(n15166), .B(n15165), .ZN(
        n15208) );
  INV_X1 U16741 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15168) );
  AOI22_X1 U16742 ( .A1(n15206), .A2(n15208), .B1(n15168), .B2(n15205), .ZN(
        P3_U3396) );
  AOI211_X1 U16743 ( .C1(n15171), .C2(n15203), .A(n15170), .B(n15169), .ZN(
        n15209) );
  INV_X1 U16744 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15172) );
  AOI22_X1 U16745 ( .A1(n15206), .A2(n15209), .B1(n15172), .B2(n15205), .ZN(
        P3_U3399) );
  AOI22_X1 U16746 ( .A1(n15175), .A2(n15203), .B1(n15174), .B2(n15173), .ZN(
        n15176) );
  AND2_X1 U16747 ( .A1(n15177), .A2(n15176), .ZN(n15211) );
  AOI22_X1 U16748 ( .A1(n15206), .A2(n15211), .B1(n8679), .B2(n15205), .ZN(
        P3_U3402) );
  INV_X1 U16749 ( .A(n15178), .ZN(n15181) );
  AOI211_X1 U16750 ( .C1(n15181), .C2(n15203), .A(n15180), .B(n15179), .ZN(
        n15212) );
  INV_X1 U16751 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15182) );
  AOI22_X1 U16752 ( .A1(n15206), .A2(n15212), .B1(n15182), .B2(n15205), .ZN(
        P3_U3405) );
  INV_X1 U16753 ( .A(n15183), .ZN(n15185) );
  AOI211_X1 U16754 ( .C1(n15203), .C2(n15186), .A(n15185), .B(n15184), .ZN(
        n15214) );
  AOI22_X1 U16755 ( .A1(n15206), .A2(n15214), .B1(n8707), .B2(n15205), .ZN(
        P3_U3408) );
  INV_X1 U16756 ( .A(n15187), .ZN(n15189) );
  AOI211_X1 U16757 ( .C1(n15190), .C2(n15203), .A(n15189), .B(n15188), .ZN(
        n15215) );
  INV_X1 U16758 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15191) );
  AOI22_X1 U16759 ( .A1(n15206), .A2(n15215), .B1(n15191), .B2(n15205), .ZN(
        P3_U3411) );
  AOI211_X1 U16760 ( .C1(n15194), .C2(n15203), .A(n15193), .B(n15192), .ZN(
        n15216) );
  INV_X1 U16761 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15195) );
  AOI22_X1 U16762 ( .A1(n15206), .A2(n15216), .B1(n15195), .B2(n15205), .ZN(
        P3_U3414) );
  INV_X1 U16763 ( .A(n15196), .ZN(n15199) );
  AOI211_X1 U16764 ( .C1(n15199), .C2(n15203), .A(n15198), .B(n15197), .ZN(
        n15218) );
  AOI22_X1 U16765 ( .A1(n15206), .A2(n15218), .B1(n8757), .B2(n15205), .ZN(
        P3_U3417) );
  INV_X1 U16766 ( .A(n15200), .ZN(n15204) );
  AOI211_X1 U16767 ( .C1(n15204), .C2(n15203), .A(n15202), .B(n15201), .ZN(
        n15221) );
  AOI22_X1 U16768 ( .A1(n15206), .A2(n15221), .B1(n8774), .B2(n15205), .ZN(
        P3_U3420) );
  AOI22_X1 U16769 ( .A1(n15222), .A2(n15207), .B1(n10412), .B2(n15219), .ZN(
        P3_U3460) );
  AOI22_X1 U16770 ( .A1(n15222), .A2(n15208), .B1(n10468), .B2(n15219), .ZN(
        P3_U3461) );
  AOI22_X1 U16771 ( .A1(n15222), .A2(n15209), .B1(n10474), .B2(n15219), .ZN(
        P3_U3462) );
  AOI22_X1 U16772 ( .A1(n15222), .A2(n15211), .B1(n15210), .B2(n15219), .ZN(
        P3_U3463) );
  AOI22_X1 U16773 ( .A1(n15222), .A2(n15212), .B1(n10613), .B2(n15219), .ZN(
        P3_U3464) );
  AOI22_X1 U16774 ( .A1(n15222), .A2(n15214), .B1(n15213), .B2(n15219), .ZN(
        P3_U3465) );
  AOI22_X1 U16775 ( .A1(n15222), .A2(n15215), .B1(n8727), .B2(n15219), .ZN(
        P3_U3466) );
  AOI22_X1 U16776 ( .A1(n15222), .A2(n15216), .B1(n10942), .B2(n15219), .ZN(
        P3_U3467) );
  AOI22_X1 U16777 ( .A1(n15222), .A2(n15218), .B1(n15217), .B2(n15219), .ZN(
        P3_U3468) );
  AOI22_X1 U16778 ( .A1(n15222), .A2(n15221), .B1(n15220), .B2(n15219), .ZN(
        P3_U3469) );
  OAI22_X1 U16779 ( .A1(n15225), .A2(keyinput22), .B1(n15224), .B2(keyinput19), 
        .ZN(n15223) );
  AOI221_X1 U16780 ( .B1(n15225), .B2(keyinput22), .C1(keyinput19), .C2(n15224), .A(n15223), .ZN(n15237) );
  OAI22_X1 U16781 ( .A1(n15228), .A2(keyinput2), .B1(n15227), .B2(keyinput57), 
        .ZN(n15226) );
  AOI221_X1 U16782 ( .B1(n15228), .B2(keyinput2), .C1(keyinput57), .C2(n15227), 
        .A(n15226), .ZN(n15236) );
  INV_X1 U16783 ( .A(keyinput13), .ZN(n15230) );
  OAI22_X1 U16784 ( .A1(n15231), .A2(keyinput20), .B1(n15230), .B2(
        P3_ADDR_REG_10__SCAN_IN), .ZN(n15229) );
  AOI221_X1 U16785 ( .B1(n15231), .B2(keyinput20), .C1(P3_ADDR_REG_10__SCAN_IN), .C2(n15230), .A(n15229), .ZN(n15235) );
  INV_X1 U16786 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n15233) );
  OAI22_X1 U16787 ( .A1(n15233), .A2(keyinput58), .B1(n8818), .B2(keyinput12), 
        .ZN(n15232) );
  AOI221_X1 U16788 ( .B1(n15233), .B2(keyinput58), .C1(keyinput12), .C2(n8818), 
        .A(n15232), .ZN(n15234) );
  NAND4_X1 U16789 ( .A1(n15237), .A2(n15236), .A3(n15235), .A4(n15234), .ZN(
        n15376) );
  OAI22_X1 U16790 ( .A1(n15239), .A2(keyinput11), .B1(n10140), .B2(keyinput33), 
        .ZN(n15238) );
  AOI221_X1 U16791 ( .B1(n15239), .B2(keyinput11), .C1(keyinput33), .C2(n10140), .A(n15238), .ZN(n15252) );
  INV_X1 U16792 ( .A(keyinput41), .ZN(n15241) );
  OAI22_X1 U16793 ( .A1(n15242), .A2(keyinput16), .B1(n15241), .B2(
        P3_DATAO_REG_31__SCAN_IN), .ZN(n15240) );
  AOI221_X1 U16794 ( .B1(n15242), .B2(keyinput16), .C1(
        P3_DATAO_REG_31__SCAN_IN), .C2(n15241), .A(n15240), .ZN(n15251) );
  OAI22_X1 U16795 ( .A1(n15245), .A2(keyinput52), .B1(n15244), .B2(keyinput44), 
        .ZN(n15243) );
  AOI221_X1 U16796 ( .B1(n15245), .B2(keyinput52), .C1(keyinput44), .C2(n15244), .A(n15243), .ZN(n15250) );
  XOR2_X1 U16797 ( .A(P3_IR_REG_8__SCAN_IN), .B(keyinput15), .Z(n15248) );
  XNOR2_X1 U16798 ( .A(n15246), .B(keyinput45), .ZN(n15247) );
  NOR2_X1 U16799 ( .A1(n15248), .A2(n15247), .ZN(n15249) );
  NAND4_X1 U16800 ( .A1(n15252), .A2(n15251), .A3(n15250), .A4(n15249), .ZN(
        n15375) );
  AOI22_X1 U16801 ( .A1(n15254), .A2(keyinput10), .B1(keyinput50), .B2(n10475), 
        .ZN(n15253) );
  OAI221_X1 U16802 ( .B1(n15254), .B2(keyinput10), .C1(n10475), .C2(keyinput50), .A(n15253), .ZN(n15266) );
  AOI22_X1 U16803 ( .A1(n15257), .A2(keyinput25), .B1(keyinput51), .B2(n15256), 
        .ZN(n15255) );
  OAI221_X1 U16804 ( .B1(n15257), .B2(keyinput25), .C1(n15256), .C2(keyinput51), .A(n15255), .ZN(n15265) );
  AOI22_X1 U16805 ( .A1(n15260), .A2(keyinput7), .B1(keyinput59), .B2(n15259), 
        .ZN(n15258) );
  OAI221_X1 U16806 ( .B1(n15260), .B2(keyinput7), .C1(n15259), .C2(keyinput59), 
        .A(n15258), .ZN(n15264) );
  XOR2_X1 U16807 ( .A(n11727), .B(keyinput60), .Z(n15262) );
  XNOR2_X1 U16808 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput4), .ZN(n15261) );
  NAND2_X1 U16809 ( .A1(n15262), .A2(n15261), .ZN(n15263) );
  NOR4_X1 U16810 ( .A1(n15266), .A2(n15265), .A3(n15264), .A4(n15263), .ZN(
        n15313) );
  AOI22_X1 U16811 ( .A1(n11298), .A2(keyinput35), .B1(keyinput30), .B2(n10850), 
        .ZN(n15267) );
  OAI221_X1 U16812 ( .B1(n11298), .B2(keyinput35), .C1(n10850), .C2(keyinput30), .A(n15267), .ZN(n15277) );
  INV_X1 U16813 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n15270) );
  AOI22_X1 U16814 ( .A1(n15270), .A2(keyinput48), .B1(n15269), .B2(keyinput61), 
        .ZN(n15268) );
  OAI221_X1 U16815 ( .B1(n15270), .B2(keyinput48), .C1(n15269), .C2(keyinput61), .A(n15268), .ZN(n15276) );
  AOI22_X1 U16816 ( .A1(n11257), .A2(keyinput26), .B1(keyinput55), .B2(n15272), 
        .ZN(n15271) );
  OAI221_X1 U16817 ( .B1(n11257), .B2(keyinput26), .C1(n15272), .C2(keyinput55), .A(n15271), .ZN(n15275) );
  INV_X1 U16818 ( .A(keyinput18), .ZN(n15340) );
  AOI22_X1 U16819 ( .A1(n8679), .A2(keyinput43), .B1(P3_DATAO_REG_3__SCAN_IN), 
        .B2(n15340), .ZN(n15273) );
  OAI221_X1 U16820 ( .B1(n8679), .B2(keyinput43), .C1(n15340), .C2(
        P3_DATAO_REG_3__SCAN_IN), .A(n15273), .ZN(n15274) );
  NOR4_X1 U16821 ( .A1(n15277), .A2(n15276), .A3(n15275), .A4(n15274), .ZN(
        n15312) );
  INV_X1 U16822 ( .A(keyinput24), .ZN(n15279) );
  AOI22_X1 U16823 ( .A1(n15280), .A2(keyinput47), .B1(P3_DATAO_REG_5__SCAN_IN), 
        .B2(n15279), .ZN(n15278) );
  OAI221_X1 U16824 ( .B1(n15280), .B2(keyinput47), .C1(n15279), .C2(
        P3_DATAO_REG_5__SCAN_IN), .A(n15278), .ZN(n15285) );
  AOI22_X1 U16825 ( .A1(n15283), .A2(keyinput40), .B1(keyinput6), .B2(n15282), 
        .ZN(n15281) );
  OAI221_X1 U16826 ( .B1(n15283), .B2(keyinput40), .C1(n15282), .C2(keyinput6), 
        .A(n15281), .ZN(n15284) );
  NOR2_X1 U16827 ( .A1(n15285), .A2(n15284), .ZN(n15295) );
  INV_X1 U16828 ( .A(keyinput8), .ZN(n15286) );
  XNOR2_X1 U16829 ( .A(n15287), .B(n15286), .ZN(n15294) );
  AOI22_X1 U16830 ( .A1(n15290), .A2(keyinput53), .B1(n15289), .B2(keyinput23), 
        .ZN(n15288) );
  OAI221_X1 U16831 ( .B1(n15290), .B2(keyinput53), .C1(n15289), .C2(keyinput23), .A(n15288), .ZN(n15291) );
  INV_X1 U16832 ( .A(n15291), .ZN(n15293) );
  XNOR2_X1 U16833 ( .A(P2_REG1_REG_0__SCAN_IN), .B(keyinput34), .ZN(n15292) );
  AND4_X1 U16834 ( .A1(n15295), .A2(n15294), .A3(n15293), .A4(n15292), .ZN(
        n15311) );
  AOI22_X1 U16835 ( .A1(n15298), .A2(keyinput27), .B1(keyinput14), .B2(n15297), 
        .ZN(n15296) );
  OAI221_X1 U16836 ( .B1(n15298), .B2(keyinput27), .C1(n15297), .C2(keyinput14), .A(n15296), .ZN(n15309) );
  INV_X1 U16837 ( .A(keyinput32), .ZN(n15300) );
  AOI22_X1 U16838 ( .A1(n10087), .A2(keyinput49), .B1(P3_DATAO_REG_0__SCAN_IN), 
        .B2(n15300), .ZN(n15299) );
  OAI221_X1 U16839 ( .B1(n10087), .B2(keyinput49), .C1(n15300), .C2(
        P3_DATAO_REG_0__SCAN_IN), .A(n15299), .ZN(n15308) );
  AOI22_X1 U16840 ( .A1(n15303), .A2(keyinput56), .B1(keyinput17), .B2(n15302), 
        .ZN(n15301) );
  OAI221_X1 U16841 ( .B1(n15303), .B2(keyinput56), .C1(n15302), .C2(keyinput17), .A(n15301), .ZN(n15307) );
  XNOR2_X1 U16842 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(keyinput42), .ZN(n15305)
         );
  XNOR2_X1 U16843 ( .A(keyinput38), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n15304)
         );
  NAND2_X1 U16844 ( .A1(n15305), .A2(n15304), .ZN(n15306) );
  NOR4_X1 U16845 ( .A1(n15309), .A2(n15308), .A3(n15307), .A4(n15306), .ZN(
        n15310) );
  NAND4_X1 U16846 ( .A1(n15313), .A2(n15312), .A3(n15311), .A4(n15310), .ZN(
        n15374) );
  AOI22_X1 U16847 ( .A1(n15316), .A2(keyinput1), .B1(n15315), .B2(keyinput21), 
        .ZN(n15314) );
  OAI221_X1 U16848 ( .B1(n15316), .B2(keyinput1), .C1(n15315), .C2(keyinput21), 
        .A(n15314), .ZN(n15326) );
  AOI22_X1 U16849 ( .A1(n15319), .A2(keyinput36), .B1(keyinput46), .B2(n15318), 
        .ZN(n15317) );
  OAI221_X1 U16850 ( .B1(n15319), .B2(keyinput36), .C1(n15318), .C2(keyinput46), .A(n15317), .ZN(n15325) );
  XNOR2_X1 U16851 ( .A(P1_REG1_REG_21__SCAN_IN), .B(keyinput31), .ZN(n15323)
         );
  XNOR2_X1 U16852 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput5), .ZN(n15322) );
  XNOR2_X1 U16853 ( .A(P2_IR_REG_27__SCAN_IN), .B(keyinput0), .ZN(n15321) );
  XNOR2_X1 U16854 ( .A(keyinput28), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n15320)
         );
  NAND4_X1 U16855 ( .A1(n15323), .A2(n15322), .A3(n15321), .A4(n15320), .ZN(
        n15324) );
  NOR3_X1 U16856 ( .A1(n15326), .A2(n15325), .A3(n15324), .ZN(n15372) );
  INV_X1 U16857 ( .A(keyinput63), .ZN(n15328) );
  AOI22_X1 U16858 ( .A1(n15329), .A2(keyinput39), .B1(P1_ADDR_REG_1__SCAN_IN), 
        .B2(n15328), .ZN(n15327) );
  OAI221_X1 U16859 ( .B1(n15329), .B2(keyinput39), .C1(n15328), .C2(
        P1_ADDR_REG_1__SCAN_IN), .A(n15327), .ZN(n15339) );
  INV_X1 U16860 ( .A(keyinput37), .ZN(n15331) );
  AOI22_X1 U16861 ( .A1(n15332), .A2(keyinput29), .B1(P2_ADDR_REG_18__SCAN_IN), 
        .B2(n15331), .ZN(n15330) );
  OAI221_X1 U16862 ( .B1(n15332), .B2(keyinput29), .C1(n15331), .C2(
        P2_ADDR_REG_18__SCAN_IN), .A(n15330), .ZN(n15338) );
  XNOR2_X1 U16863 ( .A(SI_7_), .B(keyinput62), .ZN(n15336) );
  XNOR2_X1 U16864 ( .A(P2_B_REG_SCAN_IN), .B(keyinput3), .ZN(n15335) );
  XNOR2_X1 U16865 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput9), .ZN(n15334) );
  XNOR2_X1 U16866 ( .A(SI_0_), .B(keyinput54), .ZN(n15333) );
  NAND4_X1 U16867 ( .A1(n15336), .A2(n15335), .A3(n15334), .A4(n15333), .ZN(
        n15337) );
  NOR3_X1 U16868 ( .A1(n15339), .A2(n15338), .A3(n15337), .ZN(n15371) );
  NAND2_X1 U16869 ( .A1(keyinput60), .A2(keyinput7), .ZN(n15346) );
  NOR2_X1 U16870 ( .A1(keyinput30), .A2(keyinput48), .ZN(n15344) );
  NAND3_X1 U16871 ( .A1(keyinput25), .A2(keyinput51), .A3(keyinput10), .ZN(
        n15342) );
  NAND3_X1 U16872 ( .A1(keyinput55), .A2(keyinput26), .A3(n15340), .ZN(n15341)
         );
  NOR4_X1 U16873 ( .A1(keyinput50), .A2(keyinput43), .A3(n15342), .A4(n15341), 
        .ZN(n15343) );
  NAND4_X1 U16874 ( .A1(keyinput35), .A2(keyinput61), .A3(n15344), .A4(n15343), 
        .ZN(n15345) );
  NOR4_X1 U16875 ( .A1(keyinput4), .A2(keyinput59), .A3(n15346), .A4(n15345), 
        .ZN(n15369) );
  NAND2_X1 U16876 ( .A1(keyinput6), .A2(keyinput23), .ZN(n15352) );
  NOR2_X1 U16877 ( .A1(keyinput32), .A2(keyinput56), .ZN(n15350) );
  NAND3_X1 U16878 ( .A1(keyinput8), .A2(keyinput34), .A3(keyinput47), .ZN(
        n15348) );
  NAND3_X1 U16879 ( .A1(keyinput38), .A2(keyinput42), .A3(keyinput14), .ZN(
        n15347) );
  NOR4_X1 U16880 ( .A1(keyinput24), .A2(keyinput27), .A3(n15348), .A4(n15347), 
        .ZN(n15349) );
  NAND4_X1 U16881 ( .A1(keyinput49), .A2(keyinput17), .A3(n15350), .A4(n15349), 
        .ZN(n15351) );
  NOR4_X1 U16882 ( .A1(keyinput40), .A2(keyinput53), .A3(n15352), .A4(n15351), 
        .ZN(n15368) );
  NAND2_X1 U16883 ( .A1(keyinput52), .A2(keyinput33), .ZN(n15358) );
  NOR2_X1 U16884 ( .A1(keyinput57), .A2(keyinput22), .ZN(n15356) );
  NAND3_X1 U16885 ( .A1(keyinput15), .A2(keyinput45), .A3(keyinput16), .ZN(
        n15354) );
  NAND3_X1 U16886 ( .A1(keyinput12), .A2(keyinput13), .A3(keyinput20), .ZN(
        n15353) );
  NOR4_X1 U16887 ( .A1(keyinput41), .A2(keyinput58), .A3(n15354), .A4(n15353), 
        .ZN(n15355) );
  NAND4_X1 U16888 ( .A1(keyinput2), .A2(keyinput19), .A3(n15356), .A4(n15355), 
        .ZN(n15357) );
  NOR4_X1 U16889 ( .A1(keyinput44), .A2(keyinput11), .A3(n15358), .A4(n15357), 
        .ZN(n15367) );
  NAND2_X1 U16890 ( .A1(keyinput54), .A2(keyinput3), .ZN(n15365) );
  NOR2_X1 U16891 ( .A1(keyinput31), .A2(keyinput36), .ZN(n15363) );
  NAND3_X1 U16892 ( .A1(keyinput29), .A2(keyinput37), .A3(keyinput63), .ZN(
        n15361) );
  INV_X1 U16893 ( .A(keyinput1), .ZN(n15359) );
  NAND3_X1 U16894 ( .A1(keyinput0), .A2(keyinput21), .A3(n15359), .ZN(n15360)
         );
  NOR4_X1 U16895 ( .A1(keyinput39), .A2(keyinput28), .A3(n15361), .A4(n15360), 
        .ZN(n15362) );
  NAND4_X1 U16896 ( .A1(keyinput5), .A2(keyinput46), .A3(n15363), .A4(n15362), 
        .ZN(n15364) );
  NOR4_X1 U16897 ( .A1(keyinput9), .A2(keyinput62), .A3(n15365), .A4(n15364), 
        .ZN(n15366) );
  NAND4_X1 U16898 ( .A1(n15369), .A2(n15368), .A3(n15367), .A4(n15366), .ZN(
        n15370) );
  NAND3_X1 U16899 ( .A1(n15372), .A2(n15371), .A3(n15370), .ZN(n15373) );
  NOR4_X1 U16900 ( .A1(n15376), .A2(n15375), .A3(n15374), .A4(n15373), .ZN(
        n15394) );
  NAND2_X1 U16901 ( .A1(n15378), .A2(n15377), .ZN(n15380) );
  AOI21_X1 U16902 ( .B1(n15381), .B2(n15380), .A(n15379), .ZN(n15392) );
  NOR2_X1 U16903 ( .A1(n15383), .A2(n15382), .ZN(n15391) );
  NOR2_X1 U16904 ( .A1(n15385), .A2(n15384), .ZN(n15390) );
  OAI22_X1 U16905 ( .A1(n15388), .A2(n15387), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15386), .ZN(n15389) );
  NOR4_X1 U16906 ( .A1(n15392), .A2(n15391), .A3(n15390), .A4(n15389), .ZN(
        n15393) );
  XNOR2_X1 U16907 ( .A(n15394), .B(n15393), .ZN(P1_U3215) );
  AOI21_X1 U16908 ( .B1(n15397), .B2(n15396), .A(n15395), .ZN(SUB_1596_U59) );
  OAI21_X1 U16909 ( .B1(n15399), .B2(n12931), .A(n15398), .ZN(SUB_1596_U58) );
  XOR2_X1 U16910 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15400), .Z(SUB_1596_U53) );
  AOI21_X1 U16911 ( .B1(n15403), .B2(n15402), .A(n15401), .ZN(SUB_1596_U56) );
  OAI21_X1 U16912 ( .B1(n15406), .B2(n15405), .A(n15404), .ZN(n15407) );
  XNOR2_X1 U16913 ( .A(n15407), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  AOI21_X1 U16914 ( .B1(n15410), .B2(n15409), .A(n15408), .ZN(SUB_1596_U5) );
  BUF_X1 U7194 ( .A(n8395), .Z(n6442) );
  INV_X1 U7256 ( .A(n8615), .ZN(n11871) );
  CLKBUF_X1 U7191 ( .A(n8395), .Z(n6441) );
  XNOR2_X1 U7427 ( .A(n7744), .B(P2_IR_REG_29__SCAN_IN), .ZN(n7758) );
  CLKBUF_X1 U7196 ( .A(n11584), .Z(n6911) );
  INV_X1 U7212 ( .A(n13505), .ZN(n9512) );
  CLKBUF_X1 U7224 ( .A(n8169), .Z(n8356) );
  CLKBUF_X1 U7335 ( .A(n8459), .Z(n6445) );
  CLKBUF_X1 U7461 ( .A(n9567), .Z(n13815) );
endmodule

