

module b20_C_AntiSAT_k_256_3 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, ADD_1068_U4, ADD_1068_U55, 
        ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, 
        ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, 
        ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, 
        ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, 
        P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, 
        P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, 
        P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, 
        P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, 
        P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, 
        P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, 
        P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, 
        P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, 
        P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, 
        P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, 
        P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, 
        P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447;

  INV_X4 U4999 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  BUF_X2 U5000 ( .A(n6124), .Z(n8255) );
  BUF_X1 U5001 ( .A(n7534), .Z(n7560) );
  CLKBUF_X1 U5002 ( .A(n5237), .Z(n6067) );
  OAI21_X1 U5003 ( .B1(n5964), .B2(n4735), .A(n4731), .ZN(n6417) );
  AND2_X1 U5004 ( .A1(n5149), .A2(n5150), .ZN(n5237) );
  CLKBUF_X3 U5005 ( .A(n5256), .Z(n5903) );
  INV_X1 U5006 ( .A(n6486), .ZN(n7900) );
  OR2_X1 U5007 ( .A1(n9303), .A2(n8908), .ZN(n9869) );
  INV_X1 U5008 ( .A(n5304), .ZN(n8738) );
  OAI22_X1 U5009 ( .A1(n7879), .A2(n7878), .B1(n7877), .B2(n8413), .ZN(n8097)
         );
  NAND2_X1 U5010 ( .A1(n7760), .A2(n7739), .ZN(n7700) );
  INV_X1 U5011 ( .A(n5289), .ZN(n6072) );
  NAND2_X1 U5012 ( .A1(n6904), .A2(n9086), .ZN(n6163) );
  INV_X1 U5013 ( .A(n7035), .ZN(n7671) );
  NOR3_X1 U5014 ( .A1(n9719), .A2(n9718), .A3(n9717), .ZN(n9720) );
  OR2_X1 U5015 ( .A1(n5145), .A2(n5599), .ZN(n5147) );
  AOI22_X1 U5016 ( .A1(n9187), .A2(n10203), .B1(n10194), .B2(n9222), .ZN(n9739) );
  XNOR2_X1 U5017 ( .A(n5147), .B(n5146), .ZN(n5149) );
  OAI21_X2 U5018 ( .B1(n6365), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6364), .ZN(
        n9826) );
  XNOR2_X2 U5019 ( .A(n7903), .B(n7901), .ZN(n7953) );
  OAI21_X2 U5020 ( .B1(n8043), .B2(n8039), .A(n8040), .ZN(n7903) );
  OAI21_X2 U5021 ( .B1(n5095), .B2(n7222), .A(n5094), .ZN(n8701) );
  AOI21_X2 U5022 ( .B1(n9291), .B2(n9290), .A(n8982), .ZN(n9277) );
  AND2_X1 U5023 ( .A1(n5018), .A2(n5017), .ZN(n6907) );
  XNOR2_X2 U5024 ( .A(n6299), .B(n6298), .ZN(n7942) );
  NAND2_X2 U5025 ( .A1(n8564), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6299) );
  OAI21_X1 U5026 ( .B1(n8347), .B2(n7487), .A(n7812), .ZN(n8334) );
  AOI21_X1 U5027 ( .B1(n8387), .B2(n4939), .A(n4508), .ZN(n8359) );
  INV_X2 U5028 ( .A(n6486), .ZN(n6644) );
  OR2_X1 U5029 ( .A1(n7437), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n4496) );
  NAND4_X2 U5030 ( .A1(n6505), .A2(n6504), .A3(n6503), .A4(n6502), .ZN(n8115)
         );
  NAND4_X1 U5031 ( .A1(n6661), .A2(n6660), .A3(n6659), .A4(n6658), .ZN(n8114)
         );
  NAND4_X1 U5032 ( .A1(n6516), .A2(n6515), .A3(n6514), .A4(n6513), .ZN(n10287)
         );
  CLKBUF_X2 U5033 ( .A(n6500), .Z(n7679) );
  INV_X1 U5034 ( .A(n6718), .ZN(n10138) );
  CLKBUF_X2 U5035 ( .A(n6499), .Z(n7078) );
  NOR2_X1 U5036 ( .A1(n10121), .A2(n7413), .ZN(n6820) );
  INV_X4 U5037 ( .A(n6766), .ZN(n4494) );
  NAND2_X1 U5038 ( .A1(n7865), .A2(n8261), .ZN(n6469) );
  CLKBUF_X2 U5039 ( .A(n6494), .Z(n7659) );
  INV_X4 U5040 ( .A(n5201), .ZN(n7631) );
  NOR2_X1 U5041 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5127) );
  NOR2_X1 U5042 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5965) );
  INV_X1 U5043 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6511) );
  INV_X1 U5044 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10295) );
  OAI21_X1 U5045 ( .B1(n7649), .B2(n10384), .A(n7651), .ZN(n7654) );
  OAI21_X1 U5046 ( .B1(n7649), .B2(n10369), .A(n5118), .ZN(n7648) );
  NAND2_X1 U5047 ( .A1(n7934), .A2(n7646), .ZN(n7649) );
  AND2_X1 U5048 ( .A1(n4509), .A2(n4722), .ZN(n7934) );
  AOI21_X1 U5049 ( .B1(n8859), .B2(n4647), .A(n4646), .ZN(n4645) );
  AND2_X1 U5050 ( .A1(n7644), .A2(n7643), .ZN(n4509) );
  OAI21_X1 U5051 ( .B1(n8280), .B2(n4918), .A(n4916), .ZN(n7675) );
  XNOR2_X1 U5052 ( .A(n9147), .B(n9146), .ZN(n9150) );
  NAND2_X1 U5053 ( .A1(n4608), .A2(n4607), .ZN(n5084) );
  NAND2_X1 U5054 ( .A1(n4941), .A2(n4940), .ZN(n7541) );
  NAND2_X1 U5055 ( .A1(n7908), .A2(n7907), .ZN(n7996) );
  NAND2_X1 U5056 ( .A1(n8334), .A2(n7819), .ZN(n4934) );
  OAI21_X1 U5057 ( .B1(n8334), .B2(n4505), .A(n4502), .ZN(n4941) );
  NAND2_X1 U5058 ( .A1(n4786), .A2(n4788), .ZN(n9209) );
  NAND2_X1 U5059 ( .A1(n4507), .A2(n7808), .ZN(n8347) );
  NAND2_X1 U5060 ( .A1(n9178), .A2(n9179), .ZN(n9177) );
  AND2_X1 U5061 ( .A1(n4881), .A2(n4499), .ZN(n4879) );
  NAND2_X1 U5062 ( .A1(n8359), .A2(n7811), .ZN(n4507) );
  INV_X1 U5063 ( .A(n4883), .ZN(n4499) );
  AND2_X1 U5064 ( .A1(n7627), .A2(n7582), .ZN(n4883) );
  OR2_X1 U5065 ( .A1(n7929), .A2(n8278), .ZN(n7627) );
  AND2_X1 U5066 ( .A1(n7540), .A2(n7831), .ZN(n4940) );
  AND2_X1 U5067 ( .A1(n4822), .A2(n4824), .ZN(n9276) );
  AND2_X1 U5068 ( .A1(n4672), .A2(n4503), .ZN(n4502) );
  INV_X1 U5069 ( .A(n4674), .ZN(n4505) );
  NAND2_X1 U5070 ( .A1(n4674), .A2(n4504), .ZN(n4503) );
  NAND2_X1 U5071 ( .A1(n4580), .A2(n4523), .ZN(n4508) );
  INV_X1 U5072 ( .A(n8289), .ZN(n8085) );
  AOI21_X1 U5073 ( .B1(n7604), .B2(n7692), .A(n7716), .ZN(n7281) );
  NAND2_X1 U5074 ( .A1(n4498), .A2(n7552), .ZN(n8289) );
  OAI21_X1 U5075 ( .B1(n9064), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9063), .ZN(
        n9065) );
  INV_X1 U5076 ( .A(n7819), .ZN(n4504) );
  NAND2_X1 U5077 ( .A1(n7145), .A2(n4942), .ZN(n7264) );
  NAND2_X1 U5078 ( .A1(n8281), .A2(n7558), .ZN(n4498) );
  NAND2_X1 U5079 ( .A1(n7096), .A2(n7760), .ZN(n7098) );
  NAND2_X1 U5080 ( .A1(n7096), .A2(n4506), .ZN(n7145) );
  AOI21_X1 U5081 ( .B1(n5048), .B2(n5051), .A(n8064), .ZN(n5046) );
  NAND2_X1 U5082 ( .A1(n7556), .A2(n7546), .ZN(n8281) );
  NAND2_X1 U5083 ( .A1(n4929), .A2(n4927), .ZN(n7095) );
  NAND2_X1 U5084 ( .A1(n6916), .A2(n7695), .ZN(n4929) );
  NAND2_X1 U5085 ( .A1(n6865), .A2(n7748), .ZN(n6916) );
  INV_X1 U5086 ( .A(n7522), .ZN(n7521) );
  NAND2_X1 U5087 ( .A1(n6783), .A2(n7696), .ZN(n6865) );
  OR2_X1 U5088 ( .A1(n7511), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n7522) );
  AND2_X1 U5089 ( .A1(n6969), .A2(n8952), .ZN(n6970) );
  OR2_X1 U5090 ( .A1(n7503), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n7511) );
  NAND2_X1 U5091 ( .A1(n7493), .A2(n7492), .ZN(n7503) );
  OAI22_X1 U5092 ( .A1(n6907), .A2(n6906), .B1(n6905), .B2(n8114), .ZN(n6908)
         );
  AND2_X1 U5093 ( .A1(n7097), .A2(n7760), .ZN(n4506) );
  NAND2_X1 U5094 ( .A1(n5431), .A2(n5430), .ZN(n10209) );
  NAND2_X1 U5095 ( .A1(n5479), .A2(n5478), .ZN(n10219) );
  INV_X2 U5096 ( .A(n9309), .ZN(n4495) );
  NAND2_X1 U5097 ( .A1(n7724), .A2(n7729), .ZN(n6750) );
  NAND2_X1 U5098 ( .A1(n8754), .A2(n8873), .ZN(n6740) );
  NAND2_X1 U5099 ( .A1(n6611), .A2(n7726), .ZN(n6614) );
  OR2_X1 U5100 ( .A1(n4512), .A2(n6618), .ZN(n7724) );
  OR2_X1 U5101 ( .A1(n8114), .A2(n10325), .ZN(n7748) );
  NAND2_X1 U5102 ( .A1(n6534), .A2(n6615), .ZN(n6611) );
  NAND2_X1 U5103 ( .A1(n6490), .A2(n4511), .ZN(n4512) );
  AND3_X1 U5104 ( .A1(n6871), .A2(n6870), .A3(n6869), .ZN(n10330) );
  NAND2_X1 U5105 ( .A1(n4497), .A2(n8007), .ZN(n7437) );
  INV_X1 U5106 ( .A(n6535), .ZN(n6534) );
  INV_X1 U5107 ( .A(n4497), .ZN(n7427) );
  NAND4_X1 U5108 ( .A1(n6307), .A2(n4540), .A3(n6306), .A4(n6305), .ZN(n6535)
         );
  NOR2_X1 U5109 ( .A1(n7374), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n4497) );
  AND2_X1 U5110 ( .A1(n6488), .A2(n6489), .ZN(n4511) );
  INV_X1 U5111 ( .A(n7560), .ZN(n7526) );
  AND3_X1 U5112 ( .A1(n6485), .A2(n6484), .A3(n6483), .ZN(n6618) );
  INV_X1 U5113 ( .A(n7327), .ZN(n7326) );
  INV_X1 U5114 ( .A(n6501), .ZN(n6766) );
  NAND2_X1 U5115 ( .A1(n6303), .A2(n7933), .ZN(n6500) );
  INV_X1 U5116 ( .A(n4500), .ZN(n7283) );
  NAND2_X1 U5117 ( .A1(n4500), .A2(n7282), .ZN(n7327) );
  AND2_X2 U5118 ( .A1(n5834), .A2(n5183), .ZN(n9005) );
  NAND4_X1 U5119 ( .A1(n5154), .A2(n5153), .A3(n5152), .A4(n5151), .ZN(n10121)
         );
  OR2_X1 U5120 ( .A1(n7942), .A2(n7933), .ZN(n6499) );
  CLKBUF_X1 U5121 ( .A(n5833), .Z(n6167) );
  CLKBUF_X1 U5122 ( .A(n6492), .Z(n7035) );
  NAND2_X1 U5123 ( .A1(n6278), .A2(n6277), .ZN(n7865) );
  NOR2_X1 U5124 ( .A1(n7274), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n4500) );
  XNOR2_X1 U5125 ( .A(n5156), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5833) );
  XNOR2_X1 U5126 ( .A(n6302), .B(n6301), .ZN(n7933) );
  XNOR2_X1 U5127 ( .A(n6282), .B(n6281), .ZN(n8261) );
  NAND2_X1 U5128 ( .A1(n5155), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5156) );
  AOI21_X1 U5129 ( .B1(n5964), .B2(n4546), .A(n4732), .ZN(n4731) );
  XNOR2_X1 U5130 ( .A(n5187), .B(n5186), .ZN(n9086) );
  OR2_X1 U5131 ( .A1(n6300), .A2(n6279), .ZN(n6302) );
  XNOR2_X1 U5132 ( .A(n5991), .B(n5990), .ZN(n6295) );
  AND2_X4 U5133 ( .A1(n9813), .A2(n5149), .ZN(n5241) );
  XNOR2_X1 U5134 ( .A(n5994), .B(n5993), .ZN(n6124) );
  NOR2_X1 U5135 ( .A1(n6297), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U5136 ( .A1(n5144), .A2(n5143), .ZN(n9813) );
  NAND2_X1 U5137 ( .A1(n5992), .A2(n5993), .ZN(n6297) );
  NAND2_X1 U5138 ( .A1(n4501), .A2(n6879), .ZN(n6931) );
  NOR2_X1 U5139 ( .A1(n6040), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n6062) );
  NOR2_X1 U5140 ( .A1(n4937), .A2(n6040), .ZN(n5992) );
  AND2_X1 U5141 ( .A1(n4789), .A2(n4793), .ZN(n5140) );
  INV_X1 U5142 ( .A(n6880), .ZN(n4501) );
  NAND2_X1 U5143 ( .A1(n6014), .A2(n6019), .ZN(n6482) );
  NOR2_X1 U5144 ( .A1(n4790), .A2(n5109), .ZN(n4789) );
  OR2_X1 U5145 ( .A1(n6764), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6880) );
  NAND2_X1 U5146 ( .A1(n5970), .A2(n5971), .ZN(n5065) );
  NOR2_X1 U5148 ( .A1(n5056), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5055) );
  NOR2_X2 U5149 ( .A1(n5082), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U5150 ( .A1(n6275), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n4735) );
  AND3_X1 U5151 ( .A1(n5965), .A2(n6281), .A3(n4745), .ZN(n5971) );
  AND4_X1 U5152 ( .A1(n5968), .A2(n5969), .A3(n5967), .A4(n5966), .ZN(n5970)
         );
  NAND4_X1 U5153 ( .A1(n5563), .A2(n5132), .A3(n5473), .A4(n5131), .ZN(n5133)
         );
  NAND2_X1 U5154 ( .A1(n5218), .A2(n5127), .ZN(n5279) );
  NAND2_X1 U5155 ( .A1(n6511), .A2(n10295), .ZN(n6655) );
  NAND2_X1 U5156 ( .A1(n5128), .A2(n5083), .ZN(n5082) );
  INV_X1 U5157 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5139) );
  INV_X1 U5158 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5168) );
  INV_X1 U5159 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5563) );
  INV_X1 U5160 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5566) );
  INV_X1 U5161 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5498) );
  INV_X1 U5162 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5128) );
  INV_X1 U5163 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5473) );
  INV_X1 U5164 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5083) );
  INV_X1 U5165 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5474) );
  INV_X1 U5166 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5181) );
  INV_X4 U5167 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5168 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5980) );
  INV_X1 U5169 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5132) );
  INV_X1 U5170 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5131) );
  NOR2_X1 U5171 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5957) );
  INV_X1 U5172 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5966) );
  NOR2_X1 U5173 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5969) );
  INV_X1 U5174 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6281) );
  NOR2_X1 U5175 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5958) );
  NOR2_X1 U5176 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4932) );
  NOR2_X1 U5177 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5967) );
  NOR2_X1 U5178 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5067) );
  NAND2_X1 U5179 ( .A1(n6654), .A2(n6653), .ZN(n6764) );
  NAND3_X1 U5180 ( .A1(n5970), .A2(n5971), .A3(n5067), .ZN(n5066) );
  NAND2_X1 U5181 ( .A1(n4510), .A2(n7733), .ZN(n6782) );
  NAND2_X1 U5182 ( .A1(n6749), .A2(n7743), .ZN(n4510) );
  XNOR2_X1 U5183 ( .A(n4510), .B(n6781), .ZN(n10319) );
  OAI21_X2 U5184 ( .B1(n7373), .B2(n7372), .A(n7371), .ZN(n7879) );
  AOI21_X2 U5185 ( .B1(n7318), .B2(n7317), .A(n5113), .ZN(n7373) );
  NOR2_X2 U5186 ( .A1(n6908), .A2(n6909), .ZN(n7009) );
  AND2_X4 U5187 ( .A1(n5148), .A2(n5150), .ZN(n5238) );
  OR2_X1 U5188 ( .A1(n8537), .A2(n7887), .ZN(n7803) );
  AND2_X1 U5189 ( .A1(n5014), .A2(n5012), .ZN(n5126) );
  INV_X1 U5190 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4821) );
  NAND2_X1 U5191 ( .A1(n4706), .A2(n5785), .ZN(n5805) );
  NAND2_X1 U5192 ( .A1(n4690), .A2(n5619), .ZN(n5644) );
  NAND2_X1 U5193 ( .A1(n5618), .A2(n5617), .ZN(n4690) );
  AOI21_X1 U5194 ( .B1(n4919), .B2(n4917), .A(n4553), .ZN(n4916) );
  INV_X1 U5195 ( .A(n7839), .ZN(n4917) );
  NAND2_X1 U5196 ( .A1(n6476), .A2(n7631), .ZN(n6494) );
  XNOR2_X1 U5197 ( .A(n7929), .B(n8278), .ZN(n7920) );
  NOR2_X1 U5198 ( .A1(n4537), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n4858) );
  INV_X1 U5199 ( .A(n5066), .ZN(n4859) );
  AOI21_X1 U5200 ( .B1(n4525), .B2(n4513), .A(n4593), .ZN(n4824) );
  OR2_X1 U5201 ( .A1(n9305), .A2(n4825), .ZN(n4822) );
  NOR2_X1 U5202 ( .A1(n8500), .A2(n7915), .ZN(n7834) );
  OR2_X1 U5203 ( .A1(n9730), .A2(n9193), .ZN(n8897) );
  AOI21_X1 U5204 ( .B1(n5899), .B2(n4588), .A(n5009), .ZN(n5011) );
  OAI21_X1 U5205 ( .B1(n5914), .B2(n5010), .A(n7630), .ZN(n5009) );
  AND2_X1 U5206 ( .A1(n4518), .A2(n4718), .ZN(n4717) );
  NAND2_X1 U5207 ( .A1(n5643), .A2(n5642), .ZN(n4718) );
  AND2_X1 U5208 ( .A1(n4994), .A2(n5688), .ZN(n4993) );
  NAND2_X1 U5209 ( .A1(n5668), .A2(n5667), .ZN(n4994) );
  NAND2_X1 U5210 ( .A1(n5033), .A2(n5037), .ZN(n5029) );
  OAI21_X1 U5211 ( .B1(n5035), .B2(n5034), .A(n7297), .ZN(n5033) );
  OR2_X1 U5212 ( .A1(n5034), .A2(n5031), .ZN(n5030) );
  INV_X1 U5213 ( .A(n5037), .ZN(n5031) );
  OR2_X1 U5214 ( .A1(n6845), .A2(n6844), .ZN(n6846) );
  OAI21_X1 U5215 ( .B1(n7635), .B2(n4879), .A(n4878), .ZN(n4877) );
  NAND2_X1 U5216 ( .A1(n7635), .A2(n4881), .ZN(n4878) );
  NAND2_X1 U5217 ( .A1(n4870), .A2(n4548), .ZN(n4869) );
  NAND2_X1 U5218 ( .A1(n4539), .A2(n7339), .ZN(n4870) );
  OR2_X1 U5219 ( .A1(n6527), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n6624) );
  AND2_X1 U5220 ( .A1(n6062), .A2(n5961), .ZN(n6078) );
  INV_X1 U5221 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5961) );
  INV_X1 U5222 ( .A(n5559), .ZN(n5773) );
  NOR2_X1 U5223 ( .A1(n8596), .A2(n8595), .ZN(n5088) );
  OR2_X1 U5224 ( .A1(n9160), .A2(n9715), .ZN(n8895) );
  OR2_X1 U5225 ( .A1(n5873), .A2(n9616), .ZN(n5924) );
  NOR2_X1 U5226 ( .A1(n9117), .A2(n4812), .ZN(n4811) );
  INV_X1 U5227 ( .A(n4813), .ZN(n4812) );
  AND2_X1 U5228 ( .A1(n9892), .A2(n9108), .ZN(n8908) );
  INV_X1 U5229 ( .A(n9813), .ZN(n5150) );
  NAND2_X1 U5230 ( .A1(n5807), .A2(n5806), .ZN(n5891) );
  NAND2_X1 U5231 ( .A1(n5755), .A2(n5754), .ZN(n5784) );
  INV_X1 U5232 ( .A(n5729), .ZN(n4711) );
  OAI21_X1 U5233 ( .B1(n5644), .B2(n5643), .A(n5642), .ZN(n5669) );
  NAND2_X1 U5234 ( .A1(n4719), .A2(n5003), .ZN(n5618) );
  AOI21_X1 U5235 ( .B1(n5007), .B2(n5005), .A(n5004), .ZN(n5003) );
  NAND2_X1 U5236 ( .A1(n5539), .A2(n4551), .ZN(n4719) );
  INV_X1 U5237 ( .A(n5592), .ZN(n5004) );
  AND2_X1 U5238 ( .A1(n5619), .A2(n5598), .ZN(n5617) );
  NAND2_X1 U5239 ( .A1(n4678), .A2(n4677), .ZN(n5520) );
  AOI21_X1 U5240 ( .B1(n4679), .B2(n4682), .A(n5516), .ZN(n4677) );
  INV_X1 U5241 ( .A(n4686), .ZN(n4685) );
  OAI21_X1 U5242 ( .B1(n5471), .B2(n4687), .A(n5472), .ZN(n4686) );
  NAND2_X1 U5243 ( .A1(n5419), .A2(n5422), .ZN(n4687) );
  NAND2_X1 U5244 ( .A1(n5417), .A2(n5416), .ZN(n5443) );
  NAND2_X1 U5245 ( .A1(n5406), .A2(n5121), .ZN(n5417) );
  AND2_X1 U5246 ( .A1(n6647), .A2(n5016), .ZN(n5015) );
  INV_X1 U5247 ( .A(n6650), .ZN(n5016) );
  NAND2_X1 U5248 ( .A1(n7964), .A2(n8029), .ZN(n7895) );
  OAI21_X1 U5249 ( .B1(n7675), .B2(n7674), .A(n4694), .ZN(n4693) );
  NOR2_X1 U5250 ( .A1(n7686), .A2(n4695), .ZN(n4694) );
  NOR2_X1 U5251 ( .A1(n8490), .A2(n8496), .ZN(n4695) );
  INV_X1 U5252 ( .A(n4692), .ZN(n4691) );
  OAI21_X1 U5253 ( .B1(n7685), .B2(n8273), .A(n6417), .ZN(n4692) );
  XNOR2_X1 U5254 ( .A(n6482), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n6188) );
  INV_X1 U5255 ( .A(n4862), .ZN(n4861) );
  OAI21_X1 U5256 ( .B1(n4863), .B2(n8373), .A(n7575), .ZN(n4862) );
  NAND2_X1 U5257 ( .A1(n4885), .A2(n4884), .ZN(n8388) );
  AOI21_X1 U5258 ( .B1(n4519), .B2(n4891), .A(n4552), .ZN(n4884) );
  AND2_X1 U5259 ( .A1(n6055), .A2(n5043), .ZN(n5041) );
  NAND2_X1 U5260 ( .A1(n4906), .A2(n4915), .ZN(n4903) );
  NAND2_X1 U5261 ( .A1(n4909), .A2(n4915), .ZN(n4904) );
  OR2_X1 U5262 ( .A1(n8523), .A2(n8346), .ZN(n7820) );
  NAND2_X1 U5263 ( .A1(n7479), .A2(n7478), .ZN(n7896) );
  NAND2_X1 U5264 ( .A1(n6533), .A2(n6532), .ZN(n10289) );
  AND2_X1 U5265 ( .A1(n7857), .A2(n6543), .ZN(n10285) );
  INV_X1 U5266 ( .A(n7659), .ZN(n7456) );
  INV_X1 U5267 ( .A(n6476), .ZN(n7454) );
  OR2_X1 U5268 ( .A1(n10365), .A2(n7609), .ZN(n7717) );
  NAND2_X1 U5269 ( .A1(n4936), .A2(n4935), .ZN(n5983) );
  INV_X1 U5270 ( .A(n6040), .ZN(n4936) );
  NOR2_X1 U5271 ( .A1(n5066), .A2(n4537), .ZN(n4935) );
  INV_X1 U5272 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5990) );
  INV_X1 U5273 ( .A(n9741), .ZN(n9123) );
  NOR2_X1 U5274 ( .A1(n8678), .A2(n5093), .ZN(n5092) );
  NOR2_X1 U5275 ( .A1(n4516), .A2(n7397), .ZN(n5093) );
  AND2_X1 U5276 ( .A1(n5579), .A2(n5578), .ZN(n5586) );
  OR3_X1 U5277 ( .A1(n6181), .A2(n5836), .A3(P1_U3086), .ZN(n6037) );
  NOR2_X1 U5278 ( .A1(n8936), .A2(n4527), .ZN(n4647) );
  INV_X1 U5279 ( .A(n5237), .ZN(n5928) );
  INV_X1 U5280 ( .A(n5238), .ZN(n5943) );
  INV_X1 U5281 ( .A(n5240), .ZN(n5289) );
  NAND2_X1 U5282 ( .A1(n9935), .A2(n9936), .ZN(n9934) );
  AND2_X1 U5283 ( .A1(n4775), .A2(n9234), .ZN(n4771) );
  NOR2_X1 U5284 ( .A1(n9110), .A2(n4829), .ZN(n4828) );
  INV_X1 U5285 ( .A(n4831), .ZN(n4829) );
  OR2_X1 U5286 ( .A1(n5606), .A2(n5605), .ZN(n5627) );
  OR2_X1 U5287 ( .A1(n9892), .A2(n9898), .ZN(n4831) );
  AOI21_X1 U5288 ( .B1(n7249), .B2(n7248), .A(n7247), .ZN(n9106) );
  NOR2_X1 U5289 ( .A1(n9010), .A2(n7190), .ZN(n7247) );
  INV_X1 U5290 ( .A(n8745), .ZN(n5649) );
  INV_X1 U5291 ( .A(n5307), .ZN(n5648) );
  AND4_X1 U5292 ( .A1(n5081), .A2(n4804), .A3(n5080), .A4(n4521), .ZN(n4791)
         );
  NOR2_X1 U5293 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5108) );
  NAND2_X1 U5294 ( .A1(n5356), .A2(n5355), .ZN(n5359) );
  NAND2_X1 U5295 ( .A1(n4666), .A2(n5253), .ZN(n5273) );
  NAND2_X1 U5296 ( .A1(n8115), .A2(n6646), .ZN(n6647) );
  INV_X1 U5297 ( .A(n6645), .ZN(n6646) );
  NAND2_X1 U5298 ( .A1(n7565), .A2(n7564), .ZN(n8278) );
  NAND2_X1 U5299 ( .A1(n7599), .A2(n10386), .ZN(n7596) );
  NAND2_X1 U5300 ( .A1(n7554), .A2(n7553), .ZN(n7929) );
  OAI21_X1 U5301 ( .B1(n4660), .B2(n8860), .A(n4659), .ZN(n8796) );
  AOI21_X1 U5302 ( .B1(n8782), .B2(n4662), .A(n4661), .ZN(n4660) );
  NAND2_X1 U5303 ( .A1(n8784), .A2(n8860), .ZN(n4659) );
  NAND2_X1 U5304 ( .A1(n8795), .A2(n8783), .ZN(n4661) );
  OR2_X1 U5305 ( .A1(n4566), .A2(n7770), .ZN(n4740) );
  AND2_X1 U5306 ( .A1(n4755), .A2(n4577), .ZN(n4754) );
  OR2_X1 U5307 ( .A1(n7828), .A2(n7850), .ZN(n4755) );
  NAND2_X1 U5308 ( .A1(n4758), .A2(n4759), .ZN(n4756) );
  INV_X1 U5309 ( .A(n7821), .ZN(n4759) );
  INV_X1 U5310 ( .A(n4754), .ZN(n4749) );
  INV_X1 U5311 ( .A(n4747), .ZN(n4746) );
  OAI21_X1 U5312 ( .B1(n4754), .B2(n4750), .A(n4751), .ZN(n4747) );
  AOI21_X1 U5313 ( .B1(n4753), .B2(n7857), .A(n4752), .ZN(n4751) );
  NAND2_X1 U5314 ( .A1(n4756), .A2(n4757), .ZN(n4750) );
  NAND2_X1 U5315 ( .A1(n4654), .A2(n4653), .ZN(n8836) );
  INV_X1 U5316 ( .A(n7629), .ZN(n5010) );
  NAND2_X1 U5317 ( .A1(n6482), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4962) );
  INV_X1 U5318 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5959) );
  OAI21_X1 U5319 ( .B1(n5344), .B2(n5079), .A(n5364), .ZN(n5078) );
  NAND2_X1 U5320 ( .A1(n5078), .A2(n5076), .ZN(n5074) );
  NAND2_X1 U5321 ( .A1(n5344), .A2(n5079), .ZN(n5076) );
  NOR2_X1 U5322 ( .A1(n9149), .A2(n5013), .ZN(n5012) );
  INV_X1 U5323 ( .A(n8741), .ZN(n5013) );
  INV_X1 U5324 ( .A(n5642), .ZN(n4715) );
  NAND2_X1 U5325 ( .A1(n5443), .A2(n4679), .ZN(n4678) );
  AND2_X1 U5326 ( .A1(n8014), .A2(n5049), .ZN(n5048) );
  NAND2_X1 U5327 ( .A1(n5050), .A2(n5052), .ZN(n5049) );
  INV_X1 U5328 ( .A(n5053), .ZN(n5050) );
  INV_X1 U5329 ( .A(n5052), .ZN(n5051) );
  OR2_X1 U5330 ( .A1(n7940), .A2(n7634), .ZN(n7688) );
  NAND2_X1 U5331 ( .A1(n6592), .A2(n4614), .ZN(n6685) );
  NAND2_X1 U5332 ( .A1(n6454), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4614) );
  NAND2_X1 U5333 ( .A1(n6848), .A2(n4615), .ZN(n6995) );
  NAND2_X1 U5334 ( .A1(n6683), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4615) );
  OR2_X1 U5335 ( .A1(n7197), .A2(n7196), .ZN(n7198) );
  NOR2_X1 U5336 ( .A1(n4520), .A2(n7795), .ZN(n4939) );
  NAND2_X1 U5337 ( .A1(n8389), .A2(n7794), .ZN(n4938) );
  AND2_X1 U5338 ( .A1(n7803), .A2(n8369), .ZN(n7802) );
  OR2_X1 U5339 ( .A1(n8360), .A2(n8345), .ZN(n7811) );
  NAND2_X1 U5340 ( .A1(n7447), .A2(n7446), .ZN(n7459) );
  INV_X1 U5341 ( .A(n4496), .ZN(n7447) );
  INV_X1 U5342 ( .A(n7291), .ZN(n4873) );
  INV_X1 U5343 ( .A(n7339), .ZN(n4872) );
  NOR2_X1 U5344 ( .A1(n4869), .A2(n4867), .ZN(n4866) );
  INV_X1 U5345 ( .A(n5123), .ZN(n4867) );
  AND2_X1 U5346 ( .A1(n4563), .A2(n4515), .ZN(n4853) );
  OR2_X1 U5347 ( .A1(n8111), .A2(n10339), .ZN(n7760) );
  OR2_X1 U5348 ( .A1(n7834), .A2(n7710), .ZN(n7829) );
  NAND2_X1 U5349 ( .A1(n8511), .A2(n8328), .ZN(n4915) );
  NOR2_X1 U5350 ( .A1(n4895), .A2(n4894), .ZN(n4893) );
  AND2_X1 U5351 ( .A1(n7569), .A2(n7568), .ZN(n4895) );
  INV_X1 U5352 ( .A(n7690), .ZN(n4894) );
  OR2_X1 U5353 ( .A1(n8546), .A2(n8391), .ZN(n7789) );
  OR2_X1 U5354 ( .A1(n8558), .A2(n8089), .ZN(n7777) );
  NOR2_X1 U5355 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4968) );
  INV_X1 U5356 ( .A(n5687), .ZN(n5099) );
  NAND2_X1 U5357 ( .A1(n6575), .A2(n6576), .ZN(n5265) );
  NOR2_X1 U5358 ( .A1(n5666), .A2(n5106), .ZN(n5105) );
  INV_X1 U5359 ( .A(n5638), .ZN(n5106) );
  NAND2_X1 U5360 ( .A1(n8626), .A2(n5706), .ZN(n5726) );
  NAND2_X1 U5361 ( .A1(n8596), .A2(n8595), .ZN(n5089) );
  INV_X1 U5362 ( .A(n5088), .ZN(n5087) );
  INV_X1 U5363 ( .A(n5996), .ZN(n5836) );
  NOR2_X1 U5364 ( .A1(n5157), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n5179) );
  OR2_X1 U5365 ( .A1(n9131), .A2(n9722), .ZN(n8896) );
  AOI21_X1 U5366 ( .B1(n9127), .B2(n4837), .A(n9126), .ZN(n4836) );
  INV_X1 U5367 ( .A(n9124), .ZN(n4837) );
  NAND2_X1 U5368 ( .A1(n9121), .A2(n9122), .ZN(n4833) );
  NAND2_X1 U5369 ( .A1(n9127), .A2(n4839), .ZN(n4838) );
  INV_X1 U5370 ( .A(n9125), .ZN(n4839) );
  AND2_X1 U5371 ( .A1(n9202), .A2(n8837), .ZN(n8865) );
  NOR2_X1 U5372 ( .A1(n9117), .A2(n4816), .ZN(n4809) );
  NOR2_X1 U5373 ( .A1(n4779), .A2(n9253), .ZN(n4778) );
  INV_X1 U5374 ( .A(n9137), .ZN(n4779) );
  NOR2_X1 U5375 ( .A1(n9285), .A2(n9272), .ZN(n4797) );
  NOR2_X1 U5376 ( .A1(n9911), .A2(n10240), .ZN(n4803) );
  AND2_X1 U5377 ( .A1(n4846), .A2(n4844), .ZN(n4843) );
  INV_X1 U5378 ( .A(n8885), .ZN(n4844) );
  INV_X1 U5379 ( .A(n4848), .ZN(n4841) );
  NAND2_X1 U5380 ( .A1(n7175), .A2(n10216), .ZN(n4851) );
  NOR2_X1 U5381 ( .A1(n10209), .A2(n4800), .ZN(n4799) );
  INV_X1 U5382 ( .A(n4801), .ZN(n4800) );
  NOR2_X1 U5383 ( .A1(n7393), .A2(n10183), .ZN(n4801) );
  NAND2_X1 U5384 ( .A1(n10143), .A2(n5287), .ZN(n8944) );
  NAND2_X1 U5385 ( .A1(n5833), .A2(n6904), .ZN(n5190) );
  OAI21_X1 U5386 ( .B1(n7658), .B2(SI_29_), .A(n7657), .ZN(n7662) );
  XNOR2_X1 U5387 ( .A(n7656), .B(n7655), .ZN(n7658) );
  AND2_X1 U5388 ( .A1(n5806), .A2(n5789), .ZN(n5804) );
  AND2_X1 U5389 ( .A1(n5785), .A2(n5759), .ZN(n5783) );
  AND2_X1 U5390 ( .A1(n5690), .A2(n5673), .ZN(n5688) );
  NOR2_X1 U5391 ( .A1(n5372), .A2(n5110), .ZN(n5600) );
  INV_X1 U5392 ( .A(n5133), .ZN(n4806) );
  NOR2_X1 U5393 ( .A1(n5471), .A2(n4689), .ZN(n4688) );
  INV_X1 U5394 ( .A(n5422), .ZN(n4689) );
  NAND2_X1 U5395 ( .A1(n5000), .A2(n4999), .ZN(n4998) );
  AOI21_X1 U5396 ( .B1(n5000), .B2(n4549), .A(n4997), .ZN(n4996) );
  INV_X1 U5397 ( .A(n5374), .ZN(n5002) );
  OAI211_X1 U5398 ( .C1(n4728), .C2(n4726), .A(n4724), .B(n4723), .ZN(n5303)
         );
  NAND2_X1 U5399 ( .A1(n4725), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n4724) );
  NAND2_X1 U5400 ( .A1(n4651), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4728) );
  INV_X1 U5401 ( .A(n7919), .ZN(n5059) );
  NOR2_X1 U5402 ( .A1(n7945), .A2(n5063), .ZN(n5062) );
  INV_X1 U5403 ( .A(n7917), .ZN(n5063) );
  AND2_X2 U5404 ( .A1(n6472), .A2(n6471), .ZN(n6486) );
  INV_X1 U5405 ( .A(n7975), .ZN(n5025) );
  OR2_X1 U5406 ( .A1(n8004), .A2(n8391), .ZN(n5053) );
  NAND2_X1 U5407 ( .A1(n8004), .A2(n8391), .ZN(n5052) );
  NAND2_X1 U5408 ( .A1(n7235), .A2(n8111), .ZN(n5038) );
  NOR2_X1 U5409 ( .A1(n5036), .A2(n7237), .ZN(n5035) );
  INV_X1 U5410 ( .A(n5039), .ZN(n5036) );
  AOI21_X1 U5411 ( .B1(n5029), .B2(n5030), .A(n4556), .ZN(n5026) );
  NOR2_X1 U5412 ( .A1(n5025), .A2(n5021), .ZN(n5020) );
  INV_X1 U5413 ( .A(n8031), .ZN(n5021) );
  OAI21_X1 U5414 ( .B1(n8006), .B2(n5051), .A(n5048), .ZN(n8062) );
  AND2_X1 U5415 ( .A1(n7539), .A2(n7538), .ZN(n7915) );
  AND4_X1 U5416 ( .A1(n7464), .A2(n7463), .A3(n7462), .A4(n7461), .ZN(n7887)
         );
  NAND2_X1 U5417 ( .A1(n6477), .A2(n4965), .ZN(n6131) );
  NAND2_X1 U5418 ( .A1(n4966), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4965) );
  NOR2_X1 U5419 ( .A1(n6216), .A2(n6601), .ZN(n6215) );
  OAI21_X1 U5420 ( .B1(n6187), .B2(n6188), .A(n4612), .ZN(n4611) );
  XNOR2_X1 U5421 ( .A(n4611), .B(n6498), .ZN(n6223) );
  NAND2_X1 U5422 ( .A1(n6242), .A2(n4613), .ZN(n6333) );
  NAND2_X1 U5423 ( .A1(n6640), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4613) );
  NAND2_X1 U5424 ( .A1(n6458), .A2(n6459), .ZN(n6592) );
  XNOR2_X1 U5425 ( .A(n6685), .B(n7088), .ZN(n6593) );
  NAND2_X1 U5426 ( .A1(n6688), .A2(n6689), .ZN(n6848) );
  XNOR2_X1 U5427 ( .A(n6995), .B(n7266), .ZN(n6849) );
  OR2_X1 U5428 ( .A1(n7198), .A2(n8122), .ZN(n4979) );
  XNOR2_X1 U5429 ( .A(n8172), .B(n8167), .ZN(n8149) );
  NAND2_X1 U5430 ( .A1(n8147), .A2(n4644), .ZN(n8172) );
  OR2_X1 U5431 ( .A1(n8148), .A2(n9471), .ZN(n4644) );
  NAND2_X1 U5432 ( .A1(n8149), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8174) );
  OR2_X1 U5433 ( .A1(n8146), .A2(n4973), .ZN(n4972) );
  OR2_X1 U5434 ( .A1(n8171), .A2(n8415), .ZN(n4973) );
  NAND2_X1 U5435 ( .A1(n8168), .A2(n4971), .ZN(n4970) );
  INV_X1 U5436 ( .A(n8171), .ZN(n4971) );
  INV_X1 U5437 ( .A(n4628), .ZN(n4622) );
  OAI21_X1 U5438 ( .B1(n4517), .B2(n4631), .A(n4629), .ZN(n4628) );
  NAND2_X1 U5439 ( .A1(n4630), .A2(n4641), .ZN(n4629) );
  INV_X1 U5440 ( .A(n4637), .ZN(n4630) );
  AND2_X1 U5441 ( .A1(n4877), .A2(n4579), .ZN(n4875) );
  NAND2_X1 U5442 ( .A1(n4877), .A2(n4880), .ZN(n4876) );
  NAND2_X1 U5443 ( .A1(n7843), .A2(n4881), .ZN(n4880) );
  OR2_X1 U5444 ( .A1(n7480), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n7494) );
  NAND2_X1 U5445 ( .A1(n8358), .A2(n4864), .ZN(n4863) );
  INV_X1 U5446 ( .A(n7573), .ZN(n4864) );
  AND2_X1 U5447 ( .A1(n8537), .A2(n8356), .ZN(n7573) );
  OR2_X1 U5448 ( .A1(n7459), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n7470) );
  NAND2_X1 U5449 ( .A1(n7326), .A2(n9652), .ZN(n7374) );
  AND2_X1 U5450 ( .A1(n7717), .A2(n7718), .ZN(n7693) );
  OR2_X1 U5451 ( .A1(n7157), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7274) );
  AND2_X1 U5452 ( .A1(n7090), .A2(n7089), .ZN(n7239) );
  INV_X1 U5453 ( .A(n10285), .ZN(n8426) );
  OR2_X1 U5454 ( .A1(n7850), .A2(n6543), .ZN(n8424) );
  OR2_X1 U5455 ( .A1(n7645), .A2(n10351), .ZN(n7646) );
  INV_X1 U5456 ( .A(n8283), .ZN(n8443) );
  OR2_X1 U5457 ( .A1(n8505), .A2(n7909), .ZN(n7831) );
  AOI21_X1 U5458 ( .B1(n4674), .B2(n7828), .A(n4673), .ZN(n4672) );
  INV_X1 U5459 ( .A(n7830), .ZN(n4673) );
  AOI21_X1 U5460 ( .B1(n4675), .B2(n7826), .A(n4753), .ZN(n4674) );
  INV_X1 U5461 ( .A(n4933), .ZN(n4675) );
  AND2_X1 U5462 ( .A1(n7831), .A2(n7830), .ZN(n8304) );
  INV_X1 U5463 ( .A(n8304), .ZN(n8296) );
  AND2_X1 U5464 ( .A1(n7823), .A2(n7820), .ZN(n4933) );
  NOR2_X1 U5465 ( .A1(n7579), .A2(n4913), .ZN(n4912) );
  INV_X1 U5466 ( .A(n4914), .ZN(n4913) );
  INV_X1 U5467 ( .A(n7579), .ZN(n4910) );
  AND2_X1 U5468 ( .A1(n8335), .A2(n4914), .ZN(n4911) );
  OR2_X1 U5469 ( .A1(n8523), .A2(n8327), .ZN(n4914) );
  AOI21_X1 U5470 ( .B1(n8343), .B2(n8348), .A(n7577), .ZN(n8336) );
  AND2_X1 U5471 ( .A1(n7820), .A2(n7819), .ZN(n8335) );
  AND2_X1 U5472 ( .A1(n8374), .A2(n8373), .ZN(n8375) );
  OR2_X1 U5473 ( .A1(n8061), .A2(n8392), .ZN(n8369) );
  AND2_X1 U5474 ( .A1(n8061), .A2(n8392), .ZN(n8367) );
  AOI21_X1 U5475 ( .B1(n8388), .B2(n8389), .A(n7570), .ZN(n7615) );
  INV_X1 U5476 ( .A(n4893), .ZN(n4891) );
  AOI21_X1 U5477 ( .B1(n4893), .B2(n4890), .A(n4889), .ZN(n4888) );
  INV_X1 U5478 ( .A(n7568), .ZN(n4890) );
  INV_X1 U5479 ( .A(n7691), .ZN(n4889) );
  INV_X1 U5480 ( .A(n8424), .ZN(n10286) );
  AND2_X1 U5481 ( .A1(n7691), .A2(n7690), .ZN(n8411) );
  AOI21_X1 U5482 ( .B1(n4924), .B2(n4926), .A(n4923), .ZN(n4922) );
  INV_X1 U5483 ( .A(n7773), .ZN(n4923) );
  NAND2_X1 U5484 ( .A1(n7281), .A2(n7693), .ZN(n7347) );
  AND3_X1 U5485 ( .A1(n6643), .A2(n6642), .A3(n6641), .ZN(n10321) );
  NAND2_X1 U5486 ( .A1(n6541), .A2(n7359), .ZN(n10309) );
  NAND2_X1 U5487 ( .A1(n6468), .A2(n7066), .ZN(n10356) );
  OR3_X1 U5488 ( .A1(n7865), .A2(n6417), .A3(n6532), .ZN(n7358) );
  NOR2_X1 U5489 ( .A1(n6422), .A2(n6317), .ZN(n7361) );
  INV_X1 U5490 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5979) );
  INV_X1 U5491 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5960) );
  AND2_X1 U5492 ( .A1(n6078), .A2(n4572), .ZN(n6280) );
  INV_X1 U5493 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4743) );
  NAND2_X1 U5494 ( .A1(n6078), .A2(n4744), .ZN(n6713) );
  AND2_X1 U5495 ( .A1(n6624), .A2(n6528), .ZN(n8199) );
  NAND2_X1 U5496 ( .A1(n6078), .A2(n5966), .ZN(n6151) );
  OR2_X1 U5497 ( .A1(n6019), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n6021) );
  AOI21_X1 U5498 ( .B1(n5092), .B2(n4516), .A(n4555), .ZN(n5090) );
  NAND2_X1 U5499 ( .A1(n5307), .A2(n4794), .ZN(n4795) );
  OAI21_X1 U5500 ( .B1(n6003), .B2(n5201), .A(n4559), .ZN(n4794) );
  AND2_X1 U5501 ( .A1(n6180), .A2(n5196), .ZN(n6380) );
  NAND2_X1 U5502 ( .A1(n8627), .A2(n8628), .ZN(n8626) );
  NAND2_X1 U5503 ( .A1(n5550), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5606) );
  NAND2_X1 U5504 ( .A1(n5781), .A2(n8661), .ZN(n8664) );
  OR2_X1 U5505 ( .A1(n5763), .A2(n5762), .ZN(n5818) );
  NAND2_X1 U5506 ( .A1(n6724), .A2(n5996), .ZN(n5125) );
  NAND2_X1 U5507 ( .A1(n5635), .A2(n5634), .ZN(n8713) );
  NAND2_X1 U5508 ( .A1(n4981), .A2(n8935), .ZN(n4646) );
  OAI21_X1 U5509 ( .B1(n8856), .B2(n8855), .A(n8933), .ZN(n8857) );
  NOR2_X1 U5510 ( .A1(n8743), .A2(n8752), .ZN(n8854) );
  INV_X1 U5511 ( .A(n8847), .ZN(n8853) );
  NAND2_X1 U5512 ( .A1(n5840), .A2(n5167), .ZN(n5996) );
  AND2_X1 U5513 ( .A1(n5837), .A2(n5852), .ZN(n5167) );
  NAND2_X1 U5514 ( .A1(n9934), .A2(n6091), .ZN(n4700) );
  NAND2_X1 U5515 ( .A1(n4700), .A2(n4699), .ZN(n4698) );
  INV_X1 U5516 ( .A(n9955), .ZN(n4699) );
  NOR2_X1 U5517 ( .A1(n9838), .A2(n4585), .ZN(n9853) );
  NOR2_X1 U5518 ( .A1(n9853), .A2(n9854), .ZN(n9852) );
  NAND2_X1 U5519 ( .A1(n8736), .A2(n8735), .ZN(n9095) );
  NAND2_X1 U5520 ( .A1(n4784), .A2(n4782), .ZN(n9178) );
  INV_X1 U5521 ( .A(n4783), .ZN(n4782) );
  OAI22_X1 U5522 ( .A1(n4787), .A2(n9214), .B1(n9143), .B2(n9142), .ZN(n4783)
         );
  AND2_X1 U5523 ( .A1(n5924), .A2(n5874), .ZN(n9174) );
  INV_X1 U5524 ( .A(n9127), .ZN(n9179) );
  NAND2_X1 U5525 ( .A1(n9277), .A2(n4778), .ZN(n4774) );
  AND2_X1 U5526 ( .A1(n4776), .A2(n8833), .ZN(n4775) );
  AOI21_X1 U5527 ( .B1(n4816), .B2(n4814), .A(n4590), .ZN(n4813) );
  INV_X1 U5528 ( .A(n9115), .ZN(n4814) );
  NAND2_X1 U5529 ( .A1(n4781), .A2(n8819), .ZN(n4780) );
  INV_X1 U5530 ( .A(n9277), .ZN(n4781) );
  AND2_X1 U5531 ( .A1(n8869), .A2(n8911), .ZN(n9290) );
  NAND2_X1 U5532 ( .A1(n4828), .A2(n9109), .ZN(n4827) );
  AND2_X1 U5533 ( .A1(n8870), .A2(n8909), .ZN(n9876) );
  AOI21_X1 U5534 ( .B1(n9318), .B2(n4762), .A(n4761), .ZN(n4760) );
  INV_X1 U5535 ( .A(n8906), .ZN(n4762) );
  NAND2_X1 U5536 ( .A1(n9321), .A2(n5115), .ZN(n9305) );
  OR2_X1 U5537 ( .A1(n4802), .A2(n9908), .ZN(n5115) );
  OR2_X1 U5538 ( .A1(n10209), .A2(n10216), .ZN(n8787) );
  AND2_X1 U5539 ( .A1(n8790), .A2(n8962), .ZN(n8885) );
  NAND2_X1 U5540 ( .A1(n4847), .A2(n4851), .ZN(n4846) );
  INV_X1 U5541 ( .A(n4849), .ZN(n4847) );
  AOI21_X1 U5542 ( .B1(n7103), .B2(n4852), .A(n4850), .ZN(n4849) );
  AND2_X1 U5543 ( .A1(n4851), .A2(n4852), .ZN(n4848) );
  OR2_X1 U5544 ( .A1(n7393), .A2(n9012), .ZN(n4852) );
  AOI21_X1 U5545 ( .B1(n7020), .B2(n7029), .A(n5112), .ZN(n7104) );
  NAND2_X1 U5546 ( .A1(n10057), .A2(n4801), .ZN(n7171) );
  NOR2_X1 U5547 ( .A1(n6826), .A2(n10091), .ZN(n10096) );
  NOR2_X1 U5548 ( .A1(n10244), .A2(n6167), .ZN(n6161) );
  INV_X1 U5549 ( .A(n9180), .ZN(n9715) );
  INV_X1 U5550 ( .A(n9298), .ZN(n9787) );
  NAND2_X1 U5551 ( .A1(n5603), .A2(n5602), .ZN(n9892) );
  INV_X1 U5552 ( .A(n10053), .ZN(n10179) );
  AOI21_X1 U5553 ( .B1(n5854), .B2(n5853), .A(n6059), .ZN(n6172) );
  AOI21_X1 U5554 ( .B1(n10113), .B2(n6159), .A(n6158), .ZN(n6722) );
  INV_X1 U5555 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5599) );
  XNOR2_X1 U5556 ( .A(n7662), .B(n7661), .ZN(n8739) );
  XNOR2_X1 U5557 ( .A(n7658), .B(SI_29_), .ZN(n8744) );
  NAND2_X1 U5558 ( .A1(n5899), .A2(n5898), .ZN(n5915) );
  AND2_X1 U5559 ( .A1(n4521), .A2(n5141), .ZN(n4820) );
  XNOR2_X1 U5560 ( .A(n5891), .B(n5890), .ZN(n8577) );
  NAND2_X1 U5561 ( .A1(n4710), .A2(n4708), .ZN(n5753) );
  AOI21_X1 U5562 ( .B1(n4541), .B2(n4716), .A(n4709), .ZN(n4708) );
  INV_X1 U5563 ( .A(n5728), .ZN(n4709) );
  AND2_X1 U5564 ( .A1(n5754), .A2(n5733), .ZN(n5752) );
  XNOR2_X1 U5565 ( .A(n5835), .B(P1_IR_REG_23__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U5566 ( .A1(n5834), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5835) );
  NAND2_X1 U5567 ( .A1(n4712), .A2(n4713), .ZN(n5730) );
  NAND2_X1 U5568 ( .A1(n4987), .A2(n4988), .ZN(n5710) );
  OR2_X1 U5569 ( .A1(n5669), .A2(n4991), .ZN(n4987) );
  OAI21_X1 U5570 ( .B1(n5539), .B2(n5561), .A(n5007), .ZN(n5594) );
  NAND2_X1 U5571 ( .A1(n5539), .A2(n5538), .ZN(n5562) );
  NAND2_X1 U5572 ( .A1(n4676), .A2(n4679), .ZN(n5517) );
  OR2_X1 U5573 ( .A1(n5443), .A2(n4682), .ZN(n4676) );
  XNOR2_X1 U5574 ( .A(n5401), .B(n5400), .ZN(n7036) );
  OAI21_X1 U5575 ( .B1(n5359), .B2(n5002), .A(n5000), .ZN(n5401) );
  NAND2_X1 U5576 ( .A1(n4720), .A2(n5334), .ZN(n5356) );
  INV_X1 U5577 ( .A(n5276), .ZN(n4767) );
  NAND2_X1 U5578 ( .A1(n4667), .A2(n5225), .ZN(n5250) );
  XNOR2_X1 U5579 ( .A(n5251), .B(SI_2_), .ZN(n5249) );
  AND3_X1 U5580 ( .A1(n6922), .A2(n6921), .A3(n6920), .ZN(n10334) );
  AND3_X1 U5581 ( .A1(n7498), .A2(n7497), .A3(n7496), .ZN(n8346) );
  AOI21_X1 U5582 ( .B1(n8316), .B2(n7558), .A(n7515), .ZN(n8000) );
  INV_X1 U5583 ( .A(n8094), .ZN(n8081) );
  AOI21_X1 U5584 ( .B1(n7866), .B2(n7865), .A(n4730), .ZN(n7868) );
  AOI21_X1 U5585 ( .B1(n4693), .B2(n4691), .A(n7867), .ZN(n4730) );
  INV_X1 U5586 ( .A(n7066), .ZN(n7872) );
  INV_X1 U5587 ( .A(n7915), .ZN(n8298) );
  INV_X1 U5588 ( .A(n8000), .ZN(n8328) );
  INV_X1 U5589 ( .A(n7887), .ZN(n8356) );
  INV_X1 U5590 ( .A(n8071), .ZN(n8402) );
  OR2_X1 U5591 ( .A1(n6500), .A2(n10298), .ZN(n6503) );
  OR2_X1 U5592 ( .A1(n7078), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6504) );
  AND2_X1 U5593 ( .A1(n4534), .A2(n4954), .ZN(n6982) );
  NAND2_X1 U5594 ( .A1(n7272), .A2(n7271), .ZN(n10365) );
  INV_X1 U5595 ( .A(n8420), .ZN(n10296) );
  NAND2_X1 U5596 ( .A1(n7673), .A2(n7672), .ZN(n8490) );
  AOI21_X1 U5597 ( .B1(n7591), .B2(n10289), .A(n7590), .ZN(n7599) );
  NAND2_X1 U5598 ( .A1(n7589), .A2(n7588), .ZN(n7590) );
  AOI21_X1 U5599 ( .B1(n8641), .B2(n5591), .A(n5590), .ZN(n8655) );
  OR2_X1 U5600 ( .A1(n5610), .A2(n5609), .ZN(n9898) );
  INV_X1 U5601 ( .A(n10118), .ZN(n9013) );
  INV_X1 U5602 ( .A(n9091), .ZN(n9711) );
  NAND2_X1 U5603 ( .A1(n5283), .A2(n4664), .ZN(n10078) );
  INV_X1 U5604 ( .A(n4665), .ZN(n4664) );
  OAI21_X1 U5605 ( .B1(n6639), .B2(n5304), .A(n4538), .ZN(n4665) );
  NAND2_X1 U5606 ( .A1(n5238), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5199) );
  AND2_X1 U5607 ( .A1(n5108), .A2(n4568), .ZN(n5107) );
  AOI21_X1 U5608 ( .B1(n8758), .B2(n8855), .A(n4663), .ZN(n8759) );
  AND2_X1 U5609 ( .A1(n8878), .A2(n8781), .ZN(n4662) );
  INV_X1 U5610 ( .A(n7769), .ZN(n4742) );
  AOI21_X1 U5611 ( .B1(n8796), .B2(n8786), .A(n8785), .ZN(n8789) );
  AND3_X1 U5612 ( .A1(n4741), .A2(n4740), .A3(n4571), .ZN(n7776) );
  AOI21_X1 U5613 ( .B1(n8816), .B2(n8815), .A(n8908), .ZN(n8822) );
  NAND2_X1 U5614 ( .A1(n4758), .A2(n8335), .ZN(n4757) );
  NOR2_X1 U5615 ( .A1(n7824), .A2(n7857), .ZN(n4752) );
  NAND2_X1 U5616 ( .A1(n4655), .A2(n4543), .ZN(n4654) );
  NAND2_X1 U5617 ( .A1(n4656), .A2(n4777), .ZN(n4655) );
  OR2_X1 U5618 ( .A1(n8832), .A2(n8831), .ZN(n4653) );
  NAND2_X1 U5619 ( .A1(n4749), .A2(n4756), .ZN(n4748) );
  AND2_X1 U5620 ( .A1(n7693), .A2(n7692), .ZN(n7770) );
  INV_X1 U5621 ( .A(n5593), .ZN(n5006) );
  INV_X1 U5622 ( .A(n5038), .ZN(n5034) );
  NAND2_X1 U5623 ( .A1(n7296), .A2(n8110), .ZN(n5037) );
  MUX2_X1 U5624 ( .A(n8844), .B(n8843), .S(n8855), .Z(n8849) );
  NAND2_X1 U5625 ( .A1(n5014), .A2(n4601), .ZN(n8927) );
  INV_X1 U5626 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5129) );
  INV_X1 U5627 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4805) );
  AND2_X1 U5628 ( .A1(n5561), .A2(n5006), .ZN(n5005) );
  NAND2_X1 U5629 ( .A1(n5543), .A2(n5542), .ZN(n5592) );
  INV_X1 U5630 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5418) );
  INV_X1 U5631 ( .A(n5399), .ZN(n4997) );
  INV_X1 U5632 ( .A(n5400), .ZN(n4999) );
  NAND2_X1 U5633 ( .A1(n4668), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4651) );
  NAND2_X1 U5634 ( .A1(n4652), .A2(n5168), .ZN(n4727) );
  NAND2_X1 U5635 ( .A1(n4670), .A2(n4669), .ZN(n4652) );
  NAND2_X1 U5636 ( .A1(n4958), .A2(n4957), .ZN(n6192) );
  NAND2_X1 U5637 ( .A1(n6135), .A2(n4962), .ZN(n4957) );
  OR2_X1 U5638 ( .A1(n6215), .A2(n4959), .ZN(n4958) );
  NAND2_X1 U5639 ( .A1(n4962), .A2(n6132), .ZN(n4959) );
  OR2_X1 U5640 ( .A1(n6389), .A2(n6388), .ZN(n6390) );
  NAND2_X1 U5641 ( .A1(n7202), .A2(n7203), .ZN(n8123) );
  NAND2_X1 U5642 ( .A1(n8249), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4639) );
  NAND2_X1 U5643 ( .A1(n8224), .A2(n8247), .ZN(n4637) );
  AOI21_X1 U5644 ( .B1(n4558), .B2(n7627), .A(n4882), .ZN(n4881) );
  NOR2_X1 U5645 ( .A1(n7853), .A2(n7949), .ZN(n4882) );
  NAND2_X1 U5646 ( .A1(n4721), .A2(n7920), .ZN(n4918) );
  NAND2_X1 U5647 ( .A1(n8276), .A2(n7839), .ZN(n4721) );
  INV_X1 U5648 ( .A(n4918), .ZN(n4919) );
  INV_X1 U5649 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8007) );
  INV_X1 U5650 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6879) );
  OR2_X1 U5651 ( .A1(n8443), .A2(n8289), .ZN(n7582) );
  INV_X1 U5652 ( .A(n7580), .ZN(n4899) );
  NAND2_X1 U5653 ( .A1(n4902), .A2(n7580), .ZN(n4901) );
  INV_X1 U5654 ( .A(n4904), .ZN(n4902) );
  OR2_X1 U5655 ( .A1(n7896), .A2(n7897), .ZN(n7812) );
  INV_X1 U5656 ( .A(n4925), .ZN(n4924) );
  OAI21_X1 U5657 ( .B1(n7693), .B2(n4926), .A(n7772), .ZN(n4925) );
  INV_X1 U5658 ( .A(n7717), .ZN(n4926) );
  INV_X1 U5659 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4734) );
  AOI22_X1 U5660 ( .A1(n6279), .A2(n4734), .B1(n4733), .B2(
        P2_IR_REG_31__SCAN_IN), .ZN(n4732) );
  NAND2_X1 U5661 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(n4734), .ZN(n4733) );
  AND2_X1 U5662 ( .A1(n5120), .A2(n4545), .ZN(n4744) );
  NAND2_X1 U5663 ( .A1(n5959), .A2(n5057), .ZN(n5056) );
  NOR2_X1 U5664 ( .A1(n5447), .A2(n7388), .ZN(n5432) );
  AND2_X1 U5665 ( .A1(n5549), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U5666 ( .A1(n5073), .A2(n5075), .ZN(n5388) );
  NAND2_X1 U5667 ( .A1(n5077), .A2(n5079), .ZN(n5075) );
  INV_X1 U5668 ( .A(n5078), .ZN(n5077) );
  INV_X1 U5669 ( .A(n4983), .ZN(n4982) );
  OAI21_X1 U5670 ( .B1(n8864), .B2(n8861), .A(n4984), .ZN(n4983) );
  NAND2_X1 U5671 ( .A1(n8939), .A2(n8995), .ZN(n4984) );
  INV_X1 U5672 ( .A(n8927), .ZN(n8851) );
  OR2_X1 U5673 ( .A1(n9095), .A2(n9094), .ZN(n8933) );
  AOI21_X1 U5674 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n10015), .A(n10010), .ZN(
        n7114) );
  NAND2_X1 U5675 ( .A1(n8739), .A2(n8738), .ZN(n5014) );
  NAND2_X1 U5676 ( .A1(n4788), .A2(n8898), .ZN(n4787) );
  AND2_X1 U5677 ( .A1(n8985), .A2(n9185), .ZN(n9143) );
  INV_X1 U5678 ( .A(n4787), .ZN(n4785) );
  AND2_X1 U5679 ( .A1(n9210), .A2(n8900), .ZN(n4788) );
  AND2_X1 U5680 ( .A1(n9292), .A2(n4574), .ZN(n9216) );
  NAND2_X1 U5681 ( .A1(n4826), .A2(n4513), .ZN(n4825) );
  INV_X1 U5682 ( .A(n9111), .ZN(n4826) );
  OR2_X1 U5683 ( .A1(n9330), .A2(n9908), .ZN(n8973) );
  OR2_X1 U5684 ( .A1(n10240), .A2(n9907), .ZN(n8967) );
  INV_X1 U5685 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5392) );
  OR2_X1 U5686 ( .A1(n5393), .A2(n5392), .ZN(n5447) );
  NAND2_X1 U5687 ( .A1(n8944), .A2(n8761), .ZN(n4663) );
  NAND2_X1 U5688 ( .A1(n10117), .A2(n7413), .ZN(n6826) );
  NAND2_X1 U5689 ( .A1(n6167), .A2(n9005), .ZN(n8931) );
  INV_X1 U5690 ( .A(SI_23_), .ZN(n9615) );
  AND2_X1 U5691 ( .A1(n4805), .A2(n5129), .ZN(n4804) );
  AND2_X1 U5692 ( .A1(n5914), .A2(n5897), .ZN(n5898) );
  NAND2_X1 U5693 ( .A1(n5893), .A2(n5892), .ZN(n5899) );
  AND2_X1 U5694 ( .A1(n4714), .A2(n4986), .ZN(n4713) );
  AOI21_X1 U5695 ( .B1(n4518), .B2(n4991), .A(n4596), .ZN(n4986) );
  NAND2_X1 U5696 ( .A1(n4717), .A2(n4715), .ZN(n4714) );
  INV_X1 U5697 ( .A(n4717), .ZN(n4716) );
  AOI21_X1 U5698 ( .B1(n4993), .B2(n4990), .A(n4989), .ZN(n4988) );
  INV_X1 U5699 ( .A(n5690), .ZN(n4989) );
  INV_X1 U5700 ( .A(n5667), .ZN(n4990) );
  INV_X1 U5701 ( .A(n4993), .ZN(n4991) );
  INV_X1 U5702 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9386) );
  INV_X1 U5703 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5130) );
  INV_X1 U5704 ( .A(n5008), .ZN(n5007) );
  OAI21_X1 U5705 ( .B1(n5561), .B2(n5538), .A(n5541), .ZN(n5008) );
  NAND2_X1 U5706 ( .A1(n5536), .A2(n5535), .ZN(n5539) );
  AOI21_X1 U5707 ( .B1(n4681), .B2(n4680), .A(n4595), .ZN(n4679) );
  INV_X1 U5708 ( .A(n4688), .ZN(n4680) );
  INV_X1 U5709 ( .A(n5001), .ZN(n5000) );
  OAI21_X1 U5710 ( .B1(n5002), .B2(n5358), .A(n5378), .ZN(n5001) );
  NOR2_X1 U5711 ( .A1(n4767), .A2(n4536), .ZN(n4765) );
  OR2_X1 U5712 ( .A1(n5301), .A2(n4536), .ZN(n4763) );
  OAI21_X1 U5713 ( .B1(n5201), .B2(n6004), .A(n4648), .ZN(n5224) );
  NAND2_X1 U5714 ( .A1(n5201), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4648) );
  NOR2_X2 U5715 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5218) );
  INV_X1 U5716 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4669) );
  INV_X1 U5717 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4668) );
  AND2_X1 U5718 ( .A1(n8029), .A2(n7890), .ZN(n7962) );
  NAND2_X1 U5719 ( .A1(n7895), .A2(n8031), .ZN(n7973) );
  NAND2_X1 U5720 ( .A1(n5028), .A2(n5029), .ZN(n7983) );
  OR2_X1 U5721 ( .A1(n7034), .A2(n5030), .ZN(n5028) );
  INV_X1 U5722 ( .A(n8090), .ZN(n8080) );
  OR2_X1 U5723 ( .A1(n5992), .A2(n6279), .ZN(n5994) );
  OAI21_X1 U5724 ( .B1(n7715), .B2(n6417), .A(n6531), .ZN(n7867) );
  AND2_X1 U5725 ( .A1(n7682), .A2(n7681), .ZN(n8103) );
  AND2_X1 U5726 ( .A1(n7682), .A2(n7587), .ZN(n7634) );
  INV_X1 U5727 ( .A(n7078), .ZN(n7558) );
  INV_X1 U5728 ( .A(n7679), .ZN(n7559) );
  OR2_X1 U5729 ( .A1(n6215), .A2(n6133), .ZN(n4961) );
  INV_X1 U5730 ( .A(n6135), .ZN(n4960) );
  AOI21_X1 U5731 ( .B1(n6225), .B2(n6194), .A(n6195), .ZN(n6247) );
  INV_X1 U5732 ( .A(n6778), .ZN(n6248) );
  NAND2_X1 U5733 ( .A1(n6250), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4964) );
  NAND2_X1 U5734 ( .A1(n6334), .A2(n6335), .ZN(n6336) );
  AND2_X1 U5735 ( .A1(n4963), .A2(n4964), .ZN(n6343) );
  OR2_X1 U5736 ( .A1(n6390), .A2(n6919), .ZN(n4943) );
  NAND2_X1 U5737 ( .A1(n6456), .A2(n6457), .ZN(n6458) );
  AND2_X1 U5738 ( .A1(n7088), .A2(n4946), .ZN(n4945) );
  INV_X1 U5739 ( .A(n6583), .ZN(n4947) );
  NAND2_X1 U5740 ( .A1(n6686), .A2(n6687), .ZN(n6688) );
  NAND2_X1 U5741 ( .A1(n6996), .A2(n6997), .ZN(n6998) );
  NAND2_X1 U5742 ( .A1(n6998), .A2(n6999), .ZN(n7202) );
  XNOR2_X1 U5743 ( .A(n8123), .B(n7320), .ZN(n7204) );
  NAND2_X1 U5744 ( .A1(n4533), .A2(n4979), .ZN(n4978) );
  INV_X1 U5745 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9652) );
  OR2_X1 U5746 ( .A1(n8146), .A2(n8415), .ZN(n4975) );
  AND3_X1 U5747 ( .A1(n4970), .A2(n4604), .A3(n4972), .ZN(n8221) );
  OAI21_X1 U5748 ( .B1(n8256), .B2(n4635), .A(n4634), .ZN(n4633) );
  NOR2_X1 U5749 ( .A1(n4636), .A2(n8250), .ZN(n4635) );
  NAND2_X1 U5750 ( .A1(n8256), .A2(n4639), .ZN(n4634) );
  INV_X1 U5751 ( .A(n4639), .ZN(n4636) );
  NAND2_X1 U5752 ( .A1(n8257), .A2(n4637), .ZN(n4631) );
  NAND2_X1 U5753 ( .A1(n7521), .A2(n7520), .ZN(n7532) );
  INV_X1 U5754 ( .A(n7494), .ZN(n7493) );
  NAND2_X1 U5755 ( .A1(n7469), .A2(n7468), .ZN(n7480) );
  INV_X1 U5756 ( .A(n7470), .ZN(n7469) );
  INV_X1 U5757 ( .A(n8401), .ZN(n8423) );
  NOR2_X1 U5758 ( .A1(n4873), .A2(n4872), .ZN(n4871) );
  INV_X1 U5759 ( .A(n7076), .ZN(n7075) );
  OR2_X1 U5760 ( .A1(n6931), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7076) );
  INV_X1 U5761 ( .A(n8109), .ZN(n7982) );
  INV_X1 U5762 ( .A(n7055), .ZN(n4854) );
  INV_X1 U5763 ( .A(n7749), .ZN(n4928) );
  AND2_X1 U5764 ( .A1(n4515), .A2(n6926), .ZN(n4855) );
  NOR2_X1 U5765 ( .A1(n4857), .A2(n4856), .ZN(n6928) );
  INV_X1 U5766 ( .A(n6926), .ZN(n4856) );
  INV_X1 U5767 ( .A(n6927), .ZN(n4857) );
  NAND2_X1 U5768 ( .A1(n6773), .A2(n6772), .ZN(n6875) );
  INV_X1 U5769 ( .A(n6538), .ZN(n7721) );
  NAND2_X1 U5770 ( .A1(n8105), .A2(n10286), .ZN(n7589) );
  OR2_X1 U5771 ( .A1(n8443), .A2(n8085), .ZN(n7839) );
  AND2_X1 U5772 ( .A1(n7531), .A2(n7530), .ZN(n7913) );
  AND2_X1 U5773 ( .A1(n4900), .A2(n4897), .ZN(n8288) );
  INV_X1 U5774 ( .A(n4898), .ZN(n4897) );
  OR2_X1 U5775 ( .A1(n8336), .A2(n4901), .ZN(n4900) );
  OAI21_X1 U5776 ( .B1(n4903), .B2(n4899), .A(n4514), .ZN(n4898) );
  OAI21_X1 U5777 ( .B1(n8387), .B2(n8389), .A(n7794), .ZN(n8368) );
  AND2_X1 U5778 ( .A1(n7039), .A2(n7038), .ZN(n10339) );
  OR2_X1 U5779 ( .A1(n6548), .A2(n7872), .ZN(n10351) );
  AND2_X1 U5780 ( .A1(n6294), .A2(n6315), .ZN(n7357) );
  AND2_X1 U5781 ( .A1(n6287), .A2(n6051), .ZN(n6315) );
  INV_X1 U5782 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6301) );
  CLKBUF_X1 U5783 ( .A(n6010), .Z(n6017) );
  AND2_X1 U5784 ( .A1(n4969), .A2(n4967), .ZN(n6477) );
  NAND2_X1 U5785 ( .A1(n4560), .A2(P2_IR_REG_1__SCAN_IN), .ZN(n4969) );
  NOR2_X1 U5786 ( .A1(n4930), .A2(n4968), .ZN(n4967) );
  AND2_X1 U5787 ( .A1(n8660), .A2(n5750), .ZN(n8608) );
  INV_X1 U5788 ( .A(n5102), .ZN(n5101) );
  AOI21_X1 U5789 ( .B1(n5102), .B2(n5100), .A(n5099), .ZN(n5098) );
  INV_X1 U5790 ( .A(n5105), .ZN(n5100) );
  OR2_X1 U5791 ( .A1(n5320), .A2(n5321), .ZN(n5068) );
  AND2_X1 U5792 ( .A1(n5782), .A2(n5780), .ZN(n8661) );
  NOR2_X1 U5793 ( .A1(n8672), .A2(n5103), .ZN(n5102) );
  INV_X1 U5794 ( .A(n5665), .ZN(n5103) );
  NAND2_X1 U5795 ( .A1(n8713), .A2(n5105), .ZN(n5104) );
  OR2_X1 U5796 ( .A1(n5503), .A2(n8682), .ZN(n5526) );
  OR2_X1 U5797 ( .A1(n5694), .A2(n5693), .ZN(n5719) );
  INV_X1 U5798 ( .A(n5725), .ZN(n4607) );
  INV_X1 U5799 ( .A(n5726), .ZN(n4608) );
  AOI21_X1 U5800 ( .B1(n5391), .B2(n5097), .A(n4600), .ZN(n5094) );
  CLKBUF_X1 U5801 ( .A(n6834), .Z(n6835) );
  AND2_X1 U5802 ( .A1(n5858), .A2(n5830), .ZN(n5831) );
  NAND2_X1 U5803 ( .A1(n8634), .A2(n8635), .ZN(n5832) );
  INV_X1 U5804 ( .A(n8683), .ZN(n8726) );
  OR2_X1 U5805 ( .A1(n4564), .A2(n5088), .ZN(n5085) );
  NAND2_X1 U5806 ( .A1(n5180), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U5807 ( .A1(n5182), .A2(n5181), .ZN(n5834) );
  NAND2_X1 U5808 ( .A1(n9938), .A2(n9939), .ZN(n9937) );
  NAND2_X1 U5809 ( .A1(n9953), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4697) );
  AND2_X1 U5810 ( .A1(n9950), .A2(n6108), .ZN(n9970) );
  AOI21_X1 U5811 ( .B1(n9964), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9968), .ZN(
        n9843) );
  AOI21_X1 U5812 ( .B1(n9856), .B2(P1_REG1_REG_8__SCAN_IN), .A(n9857), .ZN(
        n6112) );
  AOI21_X1 U5813 ( .B1(n9832), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9824), .ZN(
        n9985) );
  NOR2_X1 U5814 ( .A1(n9827), .A2(n4704), .ZN(n9980) );
  AND2_X1 U5815 ( .A1(n9832), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4704) );
  NOR2_X1 U5816 ( .A1(n9980), .A2(n9981), .ZN(n9979) );
  AOI21_X1 U5817 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n10003), .A(n9995), .ZN(
        n10012) );
  XNOR2_X1 U5818 ( .A(n7124), .B(n7125), .ZN(n10025) );
  NOR2_X1 U5819 ( .A1(n10007), .A2(n4701), .ZN(n7124) );
  AND2_X1 U5820 ( .A1(n10015), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4701) );
  NAND2_X1 U5821 ( .A1(n9065), .A2(n9066), .ZN(n9079) );
  NAND2_X1 U5822 ( .A1(n9079), .A2(n4609), .ZN(n10035) );
  NAND2_X1 U5823 ( .A1(n9069), .A2(n5608), .ZN(n4609) );
  AND2_X1 U5824 ( .A1(n8896), .A2(n8988), .ZN(n9128) );
  NAND2_X1 U5825 ( .A1(n8747), .A2(n8746), .ZN(n9131) );
  NOR2_X1 U5826 ( .A1(n9157), .A2(n9131), .ZN(n9130) );
  NAND2_X1 U5827 ( .A1(n5921), .A2(n5920), .ZN(n9160) );
  NAND2_X1 U5828 ( .A1(n9173), .A2(n9723), .ZN(n9157) );
  NOR2_X1 U5829 ( .A1(n4838), .A2(n4835), .ZN(n4834) );
  INV_X1 U5830 ( .A(n9122), .ZN(n4835) );
  NAND2_X1 U5831 ( .A1(n5791), .A2(n5790), .ZN(n9202) );
  OR2_X1 U5832 ( .A1(n8745), .A2(n7244), .ZN(n5790) );
  NOR2_X1 U5833 ( .A1(n9217), .A2(n9202), .ZN(n9201) );
  NOR2_X1 U5834 ( .A1(n8912), .A2(n8865), .ZN(n9210) );
  NAND2_X1 U5835 ( .A1(n4810), .A2(n4808), .ZN(n9215) );
  AOI21_X1 U5836 ( .B1(n4809), .B2(n4813), .A(n4587), .ZN(n4808) );
  NAND2_X1 U5837 ( .A1(n9292), .A2(n4797), .ZN(n9265) );
  NAND2_X1 U5838 ( .A1(n9292), .A2(n9778), .ZN(n9279) );
  AND2_X1 U5839 ( .A1(n9877), .A2(n9787), .ZN(n9292) );
  NAND2_X1 U5840 ( .A1(n5625), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5654) );
  AND2_X1 U5841 ( .A1(n9879), .A2(n9885), .ZN(n9877) );
  NOR2_X1 U5842 ( .A1(n9326), .A2(n9892), .ZN(n9879) );
  OR2_X1 U5843 ( .A1(n8871), .A2(n8908), .ZN(n9304) );
  AOI21_X1 U5844 ( .B1(n9106), .B2(n9105), .A(n9104), .ZN(n9338) );
  AND2_X1 U5845 ( .A1(n10240), .A2(n9103), .ZN(n9104) );
  NAND2_X1 U5846 ( .A1(n7250), .A2(n9102), .ZN(n9340) );
  NAND2_X1 U5847 ( .A1(n5502), .A2(n5501), .ZN(n7190) );
  OAI21_X1 U5848 ( .B1(n7104), .B2(n4842), .A(n4840), .ZN(n7249) );
  AOI21_X1 U5849 ( .B1(n4843), .B2(n4841), .A(n4554), .ZN(n4840) );
  INV_X1 U5850 ( .A(n4843), .ZN(n4842) );
  AND2_X1 U5851 ( .A1(n10057), .A2(n4529), .ZN(n7189) );
  NAND2_X1 U5852 ( .A1(n10057), .A2(n4799), .ZN(n7169) );
  AND2_X1 U5853 ( .A1(n8783), .A2(n8781), .ZN(n10054) );
  AND2_X1 U5854 ( .A1(n8950), .A2(n8777), .ZN(n10068) );
  NOR2_X1 U5855 ( .A1(n10082), .A2(n10153), .ZN(n10071) );
  OR2_X1 U5856 ( .A1(n10081), .A2(n10078), .ZN(n10082) );
  INV_X1 U5857 ( .A(n4663), .ZN(n10079) );
  NAND2_X1 U5858 ( .A1(n10096), .A2(n10138), .ZN(n10081) );
  AND2_X1 U5859 ( .A1(n8755), .A2(n8943), .ZN(n10094) );
  INV_X1 U5860 ( .A(n8875), .ZN(n6821) );
  NAND2_X1 U5861 ( .A1(n7409), .A2(n6904), .ZN(n9339) );
  INV_X1 U5862 ( .A(n9160), .ZN(n9723) );
  NAND2_X1 U5863 ( .A1(n5761), .A2(n5760), .ZN(n9750) );
  INV_X1 U5864 ( .A(n10192), .ZN(n10216) );
  INV_X1 U5865 ( .A(n9010), .ZN(n10235) );
  INV_X1 U5866 ( .A(n10166), .ZN(n10149) );
  INV_X1 U5867 ( .A(n10227), .ZN(n10241) );
  NAND2_X1 U5868 ( .A1(n7409), .A2(n6163), .ZN(n10227) );
  NAND2_X1 U5869 ( .A1(n8855), .A2(n6904), .ZN(n10244) );
  NAND2_X1 U5870 ( .A1(n10116), .A2(n10244), .ZN(n10231) );
  INV_X1 U5871 ( .A(n6037), .ZN(n6156) );
  AND2_X1 U5872 ( .A1(n7630), .A2(n5919), .ZN(n7629) );
  XNOR2_X1 U5873 ( .A(n5162), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U5874 ( .A1(n5161), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5162) );
  XNOR2_X1 U5875 ( .A(n5164), .B(P1_IR_REG_25__SCAN_IN), .ZN(n5837) );
  XNOR2_X1 U5876 ( .A(n5166), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5852) );
  NAND2_X1 U5877 ( .A1(n4992), .A2(n5667), .ZN(n5689) );
  OR2_X1 U5878 ( .A1(n5669), .A2(n5668), .ZN(n4992) );
  INV_X1 U5879 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U5880 ( .A1(n4683), .A2(n4685), .ZN(n5497) );
  NAND2_X1 U5881 ( .A1(n5443), .A2(n4688), .ZN(n4683) );
  NAND2_X1 U5882 ( .A1(n4684), .A2(n5422), .ZN(n5470) );
  OR2_X1 U5883 ( .A1(n5443), .A2(n5419), .ZN(n4684) );
  AND2_X1 U5884 ( .A1(n5081), .A2(n5080), .ZN(n5353) );
  NAND2_X1 U5885 ( .A1(n7631), .A2(n5171), .ZN(n5203) );
  NAND2_X1 U5886 ( .A1(n5064), .A2(n7917), .ZN(n7946) );
  NAND2_X1 U5887 ( .A1(n5064), .A2(n5062), .ZN(n7947) );
  AOI21_X1 U5888 ( .B1(n5062), .B2(n5060), .A(n5059), .ZN(n5058) );
  INV_X1 U5889 ( .A(n5062), .ZN(n5061) );
  INV_X1 U5890 ( .A(n8079), .ZN(n5060) );
  NAND2_X1 U5891 ( .A1(n7034), .A2(n5039), .ZN(n7238) );
  AOI21_X1 U5892 ( .B1(n6486), .B2(n6478), .A(n6538), .ZN(n6562) );
  NAND2_X1 U5893 ( .A1(n6790), .A2(n6793), .ZN(n5017) );
  NAND2_X1 U5894 ( .A1(n5047), .A2(n5052), .ZN(n8013) );
  NAND2_X1 U5895 ( .A1(n8006), .A2(n5053), .ZN(n5047) );
  NAND2_X1 U5896 ( .A1(n5032), .A2(n5038), .ZN(n7298) );
  NAND2_X1 U5897 ( .A1(n7034), .A2(n5035), .ZN(n5032) );
  NAND2_X1 U5898 ( .A1(n5019), .A2(n5023), .ZN(n8043) );
  AOI21_X1 U5899 ( .B1(n7975), .B2(n5024), .A(n4526), .ZN(n5023) );
  OR2_X1 U5900 ( .A1(n6509), .A2(n6508), .ZN(n8090) );
  INV_X1 U5901 ( .A(n8092), .ZN(n8084) );
  NAND2_X1 U5902 ( .A1(n6323), .A2(n8430), .ZN(n8101) );
  INV_X1 U5903 ( .A(n7634), .ZN(n8105) );
  AND2_X1 U5904 ( .A1(n6145), .A2(n6144), .ZN(n10283) );
  INV_X1 U5905 ( .A(n4961), .ZN(n6134) );
  OAI21_X1 U5906 ( .B1(n6223), .B2(n10373), .A(n4610), .ZN(n6189) );
  XNOR2_X1 U5907 ( .A(n6333), .B(n6248), .ZN(n6244) );
  NAND2_X1 U5908 ( .A1(n6244), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U5909 ( .A1(n4943), .A2(n6441), .ZN(n6391) );
  AND2_X1 U5910 ( .A1(n6441), .A2(n4944), .ZN(n6444) );
  NAND2_X1 U5911 ( .A1(n4948), .A2(n6669), .ZN(n6584) );
  AND2_X1 U5912 ( .A1(n6669), .A2(n4949), .ZN(n6673) );
  NOR2_X1 U5913 ( .A1(n6984), .A2(n7610), .ZN(n4953) );
  INV_X1 U5914 ( .A(n6982), .ZN(n4951) );
  INV_X1 U5915 ( .A(n4978), .ZN(n8118) );
  NAND2_X1 U5916 ( .A1(n8174), .A2(n8175), .ZN(n8176) );
  NAND2_X1 U5917 ( .A1(n4972), .A2(n4970), .ZN(n8196) );
  XNOR2_X1 U5918 ( .A(n8221), .B(n8232), .ZN(n8197) );
  AOI21_X1 U5919 ( .B1(n8226), .B2(n8225), .A(n8224), .ZN(n8248) );
  NOR2_X1 U5920 ( .A1(n8266), .A2(n4599), .ZN(n4624) );
  INV_X1 U5921 ( .A(n4633), .ZN(n4625) );
  NAND2_X1 U5922 ( .A1(n8251), .A2(n4598), .ZN(n4616) );
  AND2_X1 U5923 ( .A1(n8256), .A2(n8250), .ZN(n4632) );
  NAND2_X1 U5924 ( .A1(n8267), .A2(n4603), .ZN(n4626) );
  NAND2_X1 U5925 ( .A1(n4622), .A2(n4619), .ZN(n4618) );
  NOR2_X1 U5926 ( .A1(n8226), .A2(n4620), .ZN(n4619) );
  INV_X1 U5927 ( .A(n4631), .ZN(n4620) );
  AND2_X1 U5928 ( .A1(n4627), .A2(n8226), .ZN(n4623) );
  NAND2_X1 U5929 ( .A1(n4517), .A2(n4641), .ZN(n4627) );
  NAND2_X1 U5930 ( .A1(n7633), .A2(n7632), .ZN(n7940) );
  OR2_X1 U5931 ( .A1(n7645), .A2(n10309), .ZN(n4722) );
  AND2_X1 U5932 ( .A1(n7544), .A2(n7543), .ZN(n8283) );
  NOR2_X1 U5933 ( .A1(n8375), .A2(n7573), .ZN(n8355) );
  OR2_X1 U5934 ( .A1(n8375), .A2(n4863), .ZN(n8354) );
  NAND2_X1 U5935 ( .A1(n7436), .A2(n7435), .ZN(n8475) );
  INV_X1 U5936 ( .A(n4868), .ZN(n7340) );
  AOI21_X1 U5937 ( .B1(n7605), .B2(n7291), .A(n4539), .ZN(n4868) );
  NAND2_X1 U5938 ( .A1(n7145), .A2(n7757), .ZN(n7263) );
  INV_X1 U5939 ( .A(n8361), .ZN(n10292) );
  NAND2_X1 U5940 ( .A1(n8433), .A2(n6610), .ZN(n8420) );
  OR2_X1 U5941 ( .A1(n6552), .A2(n6322), .ZN(n8430) );
  INV_X1 U5942 ( .A(n10304), .ZN(n6478) );
  INV_X1 U5943 ( .A(n8430), .ZN(n10294) );
  AOI21_X1 U5944 ( .B1(n8739), .B2(n7671), .A(n7660), .ZN(n8496) );
  INV_X1 U5945 ( .A(n7913), .ZN(n8500) );
  NAND2_X1 U5946 ( .A1(n4941), .A2(n7831), .ZN(n8286) );
  NAND2_X1 U5947 ( .A1(n4671), .A2(n4674), .ZN(n8303) );
  OR2_X1 U5948 ( .A1(n4934), .A2(n7828), .ZN(n4671) );
  OR2_X1 U5949 ( .A1(n7659), .A2(n7517), .ZN(n7518) );
  NAND2_X1 U5950 ( .A1(n4896), .A2(n4903), .ZN(n8297) );
  OR2_X1 U5951 ( .A1(n8336), .A2(n4904), .ZN(n4896) );
  NAND2_X1 U5952 ( .A1(n4934), .A2(n4933), .ZN(n8318) );
  NAND2_X1 U5953 ( .A1(n7510), .A2(n7509), .ZN(n8511) );
  NAND2_X1 U5954 ( .A1(n4905), .A2(n4909), .ZN(n8311) );
  NAND2_X1 U5955 ( .A1(n8336), .A2(n4912), .ZN(n4905) );
  NAND2_X1 U5956 ( .A1(n7502), .A2(n7501), .ZN(n8517) );
  NAND2_X1 U5957 ( .A1(n4908), .A2(n4914), .ZN(n8326) );
  OR2_X1 U5958 ( .A1(n8336), .A2(n8335), .ZN(n4908) );
  NAND2_X1 U5959 ( .A1(n4934), .A2(n7820), .ZN(n8324) );
  NAND2_X1 U5960 ( .A1(n7491), .A2(n7490), .ZN(n8523) );
  OR2_X1 U5961 ( .A1(n10369), .A2(n10356), .ZN(n8534) );
  NAND2_X1 U5962 ( .A1(n7458), .A2(n7457), .ZN(n8537) );
  NAND2_X1 U5963 ( .A1(n7445), .A2(n7444), .ZN(n8061) );
  NAND2_X1 U5964 ( .A1(n7426), .A2(n7425), .ZN(n8546) );
  NAND2_X1 U5965 ( .A1(n4887), .A2(n4888), .ZN(n8400) );
  OR2_X1 U5966 ( .A1(n8421), .A2(n4891), .ZN(n4887) );
  NAND2_X1 U5967 ( .A1(n7420), .A2(n7419), .ZN(n8552) );
  OR2_X1 U5968 ( .A1(n8421), .A2(n7569), .ZN(n4892) );
  NAND2_X1 U5969 ( .A1(n7370), .A2(n7369), .ZN(n8558) );
  NAND2_X1 U5970 ( .A1(n7322), .A2(n7321), .ZN(n7416) );
  NAND2_X1 U5971 ( .A1(n7347), .A2(n7717), .ZN(n7415) );
  INV_X1 U5972 ( .A(n8534), .ZN(n8559) );
  NOR2_X1 U5973 ( .A1(n5984), .A2(n5992), .ZN(n6055) );
  NAND2_X1 U5974 ( .A1(n5977), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5975) );
  OR2_X1 U5975 ( .A1(n5976), .A2(n5979), .ZN(n5978) );
  INV_X1 U5976 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7500) );
  INV_X1 U5977 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7489) );
  XNOR2_X1 U5978 ( .A(n5973), .B(n5972), .ZN(n7066) );
  INV_X1 U5979 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7477) );
  INV_X1 U5980 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n9367) );
  OR2_X1 U5981 ( .A1(n6276), .A2(n6275), .ZN(n6277) );
  NAND2_X1 U5982 ( .A1(n6276), .A2(n6275), .ZN(n6278) );
  OR2_X1 U5983 ( .A1(n6280), .A2(n6279), .ZN(n6282) );
  INV_X1 U5984 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6716) );
  INV_X1 U5985 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6626) );
  INV_X1 U5986 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9499) );
  INV_X1 U5987 ( .A(n8148), .ZN(n8145) );
  INV_X1 U5988 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6080) );
  INV_X1 U5989 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6048) );
  INV_X1 U5990 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6045) );
  INV_X1 U5991 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6032) );
  INV_X1 U5992 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6918) );
  INV_X1 U5993 ( .A(n6348), .ZN(n6868) );
  INV_X1 U5994 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6775) );
  NAND2_X1 U5995 ( .A1(n4643), .A2(n4642), .ZN(n6014) );
  NAND2_X1 U5996 ( .A1(n6013), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4642) );
  OAI21_X1 U5997 ( .B1(n4930), .B2(n6279), .A(P2_IR_REG_2__SCAN_IN), .ZN(n4643) );
  INV_X1 U5998 ( .A(n6477), .ZN(n6213) );
  NAND2_X1 U5999 ( .A1(n5902), .A2(n5901), .ZN(n9730) );
  OR2_X1 U6000 ( .A1(n8745), .A2(n9815), .ZN(n5901) );
  NAND2_X1 U6001 ( .A1(n5091), .A2(n5090), .ZN(n8598) );
  NAND2_X1 U6002 ( .A1(n7396), .A2(n5092), .ZN(n5091) );
  INV_X1 U6003 ( .A(n9784), .ZN(n9889) );
  NAND2_X1 U6004 ( .A1(n8713), .A2(n5638), .ZN(n8620) );
  INV_X1 U6005 ( .A(n5095), .ZN(n7135) );
  INV_X1 U6006 ( .A(n9767), .ZN(n9241) );
  NAND2_X1 U6007 ( .A1(n5104), .A2(n5665), .ZN(n8671) );
  INV_X1 U6008 ( .A(n7190), .ZN(n10228) );
  INV_X1 U6009 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8682) );
  AOI21_X1 U6010 ( .B1(n7396), .B2(n7397), .A(n4516), .ZN(n8679) );
  INV_X1 U6011 ( .A(n9011), .ZN(n10206) );
  INV_X1 U6012 ( .A(n9871), .ZN(n9283) );
  OR2_X1 U6013 ( .A1(n5616), .A2(n5615), .ZN(n5116) );
  AND2_X1 U6014 ( .A1(n5856), .A2(n5871), .ZN(n8680) );
  INV_X1 U6015 ( .A(n9343), .ZN(n9908) );
  INV_X1 U6016 ( .A(n5586), .ZN(n8723) );
  NAND2_X1 U6017 ( .A1(n5569), .A2(n5568), .ZN(n9911) );
  INV_X1 U6018 ( .A(n8680), .ZN(n8733) );
  OAI21_X1 U6019 ( .B1(n4645), .B2(n6904), .A(n8999), .ZN(n9000) );
  NAND2_X1 U6020 ( .A1(n8998), .A2(n6904), .ZN(n8999) );
  NAND2_X1 U6021 ( .A1(n4985), .A2(n8864), .ZN(n8863) );
  NAND2_X1 U6022 ( .A1(n8859), .A2(n8858), .ZN(n4985) );
  NAND2_X1 U6023 ( .A1(n5931), .A2(n5930), .ZN(n9180) );
  NAND2_X1 U6024 ( .A1(n5880), .A2(n5879), .ZN(n9735) );
  NAND2_X1 U6025 ( .A1(n5824), .A2(n5823), .ZN(n9741) );
  OR2_X1 U6026 ( .A1(n5862), .A2(n5943), .ZN(n5824) );
  NAND2_X1 U6027 ( .A1(n5797), .A2(n5796), .ZN(n9222) );
  NAND3_X1 U6028 ( .A1(n5296), .A2(n5122), .A3(n5295), .ZN(n6632) );
  NAND4_X1 U6029 ( .A1(n5271), .A2(n5270), .A3(n5269), .A4(n5268), .ZN(n5287)
         );
  OR2_X1 U6030 ( .A1(n5289), .A2(n5267), .ZN(n5268) );
  NAND4_X1 U6031 ( .A1(n5245), .A2(n5244), .A3(n5243), .A4(n5242), .ZN(n10089)
         );
  NAND2_X1 U6032 ( .A1(n9019), .A2(n9025), .ZN(n9018) );
  INV_X1 U6033 ( .A(n4700), .ZN(n9956) );
  INV_X1 U6034 ( .A(n4698), .ZN(n9954) );
  NOR2_X1 U6035 ( .A1(n9852), .A2(n4584), .ZN(n6098) );
  NAND2_X1 U6036 ( .A1(n6098), .A2(n6099), .ZN(n6357) );
  NOR2_X1 U6037 ( .A1(n9979), .A2(n4703), .ZN(n6360) );
  AND2_X1 U6038 ( .A1(n9978), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4703) );
  NAND2_X1 U6039 ( .A1(n6360), .A2(n6361), .ZN(n7119) );
  NOR2_X1 U6040 ( .A1(n10009), .A2(n10008), .ZN(n10007) );
  NOR2_X1 U6041 ( .A1(n9998), .A2(n4702), .ZN(n10009) );
  AND2_X1 U6042 ( .A1(n10003), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4702) );
  NOR2_X1 U6043 ( .A1(n9059), .A2(n4602), .ZN(n9060) );
  NAND2_X1 U6044 ( .A1(n9060), .A2(n9061), .ZN(n9075) );
  NOR2_X1 U6045 ( .A1(n10039), .A2(n10038), .ZN(n10037) );
  NAND2_X1 U6046 ( .A1(n9075), .A2(n4696), .ZN(n10039) );
  NAND2_X1 U6047 ( .A1(n9069), .A2(n9308), .ZN(n4696) );
  INV_X1 U6048 ( .A(n9009), .ZN(n9722) );
  OAI21_X1 U6049 ( .B1(n9188), .B2(n9125), .A(n9124), .ZN(n9172) );
  INV_X1 U6050 ( .A(n9735), .ZN(n9193) );
  NAND2_X1 U6051 ( .A1(n5813), .A2(n5812), .ZN(n9736) );
  NOR2_X1 U6052 ( .A1(n4773), .A2(n4772), .ZN(n9235) );
  INV_X1 U6053 ( .A(n4775), .ZN(n4772) );
  INV_X1 U6054 ( .A(n4774), .ZN(n4773) );
  OAI21_X1 U6055 ( .B1(n9259), .B2(n4815), .A(n4813), .ZN(n9232) );
  NAND2_X1 U6056 ( .A1(n4780), .A2(n9137), .ZN(n9252) );
  AND2_X1 U6057 ( .A1(n4817), .A2(n4818), .ZN(n9247) );
  NAND2_X1 U6058 ( .A1(n9259), .A2(n9115), .ZN(n4817) );
  NAND2_X1 U6059 ( .A1(n5692), .A2(n5691), .ZN(n9272) );
  NAND2_X1 U6060 ( .A1(n5651), .A2(n5650), .ZN(n9298) );
  NAND2_X1 U6061 ( .A1(n4823), .A2(n4513), .ZN(n9289) );
  NAND2_X1 U6062 ( .A1(n9305), .A2(n4828), .ZN(n4823) );
  NAND2_X1 U6063 ( .A1(n5624), .A2(n5623), .ZN(n9874) );
  NAND2_X1 U6064 ( .A1(n4830), .A2(n4831), .ZN(n9875) );
  OR2_X1 U6065 ( .A1(n9305), .A2(n9109), .ZN(n4830) );
  NAND2_X1 U6066 ( .A1(n4845), .A2(n4846), .ZN(n7182) );
  NAND2_X1 U6067 ( .A1(n7104), .A2(n4848), .ZN(n4845) );
  OAI21_X1 U6068 ( .B1(n7104), .B2(n7103), .A(n4852), .ZN(n7168) );
  AND2_X1 U6069 ( .A1(n10057), .A2(n6971), .ZN(n6972) );
  OR2_X1 U6070 ( .A1(n4495), .A2(n10234), .ZN(n9348) );
  NAND2_X1 U6071 ( .A1(n4770), .A2(n4769), .ZN(n10053) );
  AND2_X1 U6072 ( .A1(n5383), .A2(n4573), .ZN(n4769) );
  NAND2_X1 U6073 ( .A1(n7036), .A2(n8738), .ZN(n4770) );
  OR2_X1 U6074 ( .A1(n4495), .A2(n8995), .ZN(n9327) );
  INV_X1 U6075 ( .A(n9353), .ZN(n9301) );
  OR2_X1 U6076 ( .A1(n4495), .A2(n6727), .ZN(n9341) );
  OR2_X1 U6077 ( .A1(n8745), .A2(n6006), .ZN(n5227) );
  INV_X1 U6078 ( .A(n9322), .ZN(n10102) );
  AND4_X1 U6079 ( .A1(n5217), .A2(n5216), .A3(n5215), .A4(n5214), .ZN(n10118)
         );
  OR2_X1 U6080 ( .A1(n4495), .A2(n6726), .ZN(n9322) );
  NAND2_X1 U6081 ( .A1(n6161), .A2(n6156), .ZN(n9306) );
  INV_X1 U6082 ( .A(n9327), .ZN(n10101) );
  INV_X1 U6083 ( .A(n9341), .ZN(n10090) );
  INV_X1 U6084 ( .A(n9192), .ZN(n9344) );
  AND2_X2 U6085 ( .A1(n6722), .A2(n6162), .ZN(n10251) );
  AND2_X1 U6086 ( .A1(n9821), .A2(n7221), .ZN(n6059) );
  NAND2_X1 U6087 ( .A1(n6156), .A2(n6057), .ZN(n10113) );
  XNOR2_X1 U6088 ( .A(n7670), .B(n7669), .ZN(n9807) );
  MUX2_X1 U6089 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5142), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5143) );
  XNOR2_X1 U6090 ( .A(n4707), .B(n7629), .ZN(n8569) );
  NAND2_X1 U6091 ( .A1(n5915), .A2(n5914), .ZN(n4707) );
  NAND2_X1 U6092 ( .A1(n4819), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5177) );
  INV_X1 U6093 ( .A(n5837), .ZN(n7246) );
  INV_X1 U6094 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7070) );
  INV_X1 U6095 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9604) );
  INV_X1 U6096 ( .A(n9005), .ZN(n7068) );
  INV_X1 U6097 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6902) );
  INV_X1 U6098 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6817) );
  INV_X1 U6099 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6637) );
  INV_X1 U6100 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6529) );
  INV_X1 U6101 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6065) );
  INV_X1 U6102 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6033) );
  INV_X1 U6103 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U6104 ( .A1(n5359), .A2(n5358), .ZN(n5375) );
  INV_X1 U6105 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6008) );
  OAI21_X1 U6106 ( .B1(n5277), .B2(n4768), .A(n4766), .ZN(n5331) );
  NAND2_X1 U6107 ( .A1(n5277), .A2(n5276), .ZN(n5302) );
  OAI21_X1 U6108 ( .B1(n5220), .B2(n5219), .A(n5246), .ZN(n6100) );
  XNOR2_X1 U6109 ( .A(n4705), .B(n5204), .ZN(n6101) );
  NAND2_X1 U6110 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4705) );
  NAND2_X1 U6111 ( .A1(n6648), .A2(n6647), .ZN(n6649) );
  NAND2_X1 U6112 ( .A1(n7596), .A2(n7595), .ZN(n7598) );
  NAND2_X1 U6113 ( .A1(n10384), .A2(n9638), .ZN(n7595) );
  MUX2_X1 U6114 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9793), .S(n10274), .Z(n9712) );
  NAND2_X1 U6115 ( .A1(n6417), .A2(n7872), .ZN(n7850) );
  AND2_X1 U6116 ( .A1(n4557), .A2(n4827), .ZN(n4513) );
  OR2_X1 U6117 ( .A1(n8505), .A2(n8312), .ZN(n4514) );
  INV_X1 U6118 ( .A(n7850), .ZN(n7857) );
  NAND2_X1 U6119 ( .A1(n7759), .A2(n7094), .ZN(n4515) );
  AND2_X2 U6120 ( .A1(n7942), .A2(n7933), .ZN(n7534) );
  AND2_X1 U6121 ( .A1(n5493), .A2(n5492), .ZN(n4516) );
  AND2_X1 U6122 ( .A1(n8225), .A2(n8247), .ZN(n4517) );
  AND4_X1 U6123 ( .A1(n7432), .A2(n7431), .A3(n7430), .A4(n7429), .ZN(n8391)
         );
  INV_X1 U6124 ( .A(n4682), .ZN(n4681) );
  NAND2_X1 U6125 ( .A1(n4685), .A2(n5494), .ZN(n4682) );
  AND2_X1 U6126 ( .A1(n4988), .A2(n5707), .ZN(n4518) );
  AND2_X1 U6127 ( .A1(n4888), .A2(n4886), .ZN(n4519) );
  OR2_X1 U6128 ( .A1(n8367), .A2(n7798), .ZN(n4520) );
  AND2_X1 U6129 ( .A1(n5139), .A2(n4821), .ZN(n4521) );
  OR2_X1 U6130 ( .A1(n8116), .A2(n6615), .ZN(n4522) );
  OR2_X1 U6131 ( .A1(n7798), .A2(n7802), .ZN(n4523) );
  NAND2_X1 U6132 ( .A1(n7529), .A2(n7528), .ZN(n8312) );
  OR2_X1 U6133 ( .A1(n6040), .A2(n5066), .ZN(n4524) );
  NOR2_X1 U6134 ( .A1(n9111), .A2(n4828), .ZN(n4525) );
  NOR2_X1 U6135 ( .A1(n7898), .A2(n7576), .ZN(n4526) );
  NAND2_X1 U6136 ( .A1(n8858), .A2(n8862), .ZN(n4527) );
  AND2_X1 U6137 ( .A1(n4797), .A2(n4796), .ZN(n4528) );
  AND2_X1 U6138 ( .A1(n4799), .A2(n4798), .ZN(n4529) );
  OR2_X1 U6139 ( .A1(n5315), .A2(n5318), .ZN(n4530) );
  NAND2_X1 U6140 ( .A1(n5548), .A2(n5547), .ZN(n9330) );
  INV_X1 U6141 ( .A(n9330), .ZN(n4802) );
  AND2_X1 U6142 ( .A1(n5095), .A2(n5390), .ZN(n4531) );
  AND2_X1 U6143 ( .A1(n8117), .A2(n4978), .ZN(n4532) );
  INV_X1 U6144 ( .A(n6984), .ZN(n4955) );
  AND2_X1 U6145 ( .A1(n8117), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4533) );
  AND2_X1 U6146 ( .A1(n6980), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4534) );
  INV_X1 U6147 ( .A(n8381), .ZN(n8433) );
  AND2_X1 U6148 ( .A1(n4980), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4535) );
  NAND2_X2 U6149 ( .A1(n5905), .A2(n5559), .ZN(n5256) );
  INV_X1 U6150 ( .A(n6417), .ZN(n6468) );
  AND2_X1 U6151 ( .A1(n5303), .A2(SI_4_), .ZN(n4536) );
  NAND2_X1 U6152 ( .A1(n5128), .A2(n5081), .ZN(n5281) );
  AND2_X1 U6153 ( .A1(n9813), .A2(n5148), .ZN(n5240) );
  NAND3_X1 U6154 ( .A1(n5980), .A2(n5988), .A3(n5979), .ZN(n4537) );
  NOR2_X1 U6155 ( .A1(n5279), .A2(n5082), .ZN(n5298) );
  OR2_X1 U6156 ( .A1(n5307), .A2(n6106), .ZN(n4538) );
  INV_X1 U6157 ( .A(n8325), .ZN(n4758) );
  NOR2_X1 U6158 ( .A1(n8050), .A2(n8108), .ZN(n4539) );
  OR2_X1 U6159 ( .A1(n6501), .A2(n6559), .ZN(n4540) );
  AND2_X1 U6160 ( .A1(n4713), .A2(n4711), .ZN(n4541) );
  XNOR2_X1 U6161 ( .A(n8443), .B(n8085), .ZN(n8276) );
  INV_X1 U6162 ( .A(n8276), .ZN(n4920) );
  NOR2_X1 U6163 ( .A1(n8085), .A2(n8283), .ZN(n4542) );
  NAND2_X1 U6164 ( .A1(n5675), .A2(n5674), .ZN(n9285) );
  OR2_X1 U6165 ( .A1(n8916), .A2(n8855), .ZN(n4543) );
  INV_X1 U6166 ( .A(n8907), .ZN(n4761) );
  NAND2_X1 U6167 ( .A1(n5716), .A2(n5715), .ZN(n9763) );
  INV_X1 U6168 ( .A(n9763), .ZN(n4796) );
  OR3_X1 U6169 ( .A1(n8852), .A2(n8851), .A3(n8850), .ZN(n4544) );
  AND2_X1 U6170 ( .A1(n5966), .A2(n4745), .ZN(n4545) );
  AND2_X1 U6171 ( .A1(n5160), .A2(n5107), .ZN(n5145) );
  NAND2_X1 U6172 ( .A1(n5726), .A2(n5725), .ZN(n8607) );
  AND2_X1 U6173 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4734), .ZN(n4546) );
  AND2_X1 U6174 ( .A1(n4698), .A2(n4697), .ZN(n4547) );
  OR2_X1 U6175 ( .A1(n10365), .A2(n8107), .ZN(n4548) );
  AOI21_X1 U6176 ( .B1(n5301), .B2(n4767), .A(n4536), .ZN(n4766) );
  OR2_X1 U6177 ( .A1(n9750), .A2(n9206), .ZN(n8900) );
  NAND2_X1 U6178 ( .A1(n5524), .A2(n5523), .ZN(n10240) );
  NAND2_X1 U6179 ( .A1(n4792), .A2(n5139), .ZN(n5163) );
  NAND2_X1 U6180 ( .A1(n5735), .A2(n5734), .ZN(n9243) );
  AND2_X1 U6181 ( .A1(n5002), .A2(n4999), .ZN(n4549) );
  AND2_X1 U6182 ( .A1(n4796), .A2(n9241), .ZN(n4550) );
  INV_X1 U6183 ( .A(n4930), .ZN(n5997) );
  AND2_X1 U6184 ( .A1(n7789), .A2(n7788), .ZN(n8399) );
  INV_X1 U6185 ( .A(n8399), .ZN(n4886) );
  XNOR2_X1 U6186 ( .A(n7675), .B(n7635), .ZN(n7645) );
  AND2_X1 U6187 ( .A1(n5007), .A2(n5006), .ZN(n4551) );
  INV_X1 U6188 ( .A(n4816), .ZN(n4815) );
  NOR2_X1 U6189 ( .A1(n4550), .A2(n9114), .ZN(n4816) );
  OR2_X1 U6190 ( .A1(n8511), .A2(n8000), .ZN(n7827) );
  INV_X1 U6191 ( .A(n7827), .ZN(n4753) );
  AND2_X1 U6192 ( .A1(n8546), .A2(n8412), .ZN(n4552) );
  NOR2_X1 U6193 ( .A1(n7949), .A2(n7929), .ZN(n4553) );
  INV_X1 U6194 ( .A(n6893), .ZN(n5079) );
  INV_X1 U6195 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4966) );
  INV_X1 U6196 ( .A(n4909), .ZN(n4907) );
  AOI21_X1 U6197 ( .B1(n4911), .B2(n4910), .A(n4561), .ZN(n4909) );
  NOR2_X1 U6198 ( .A1(n10219), .A2(n9011), .ZN(n4554) );
  INV_X1 U6199 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5176) );
  AOI21_X1 U6200 ( .B1(n7973), .B2(n7974), .A(n5025), .ZN(n5022) );
  NOR2_X1 U6201 ( .A1(n5515), .A2(n5514), .ZN(n4555) );
  OR2_X1 U6202 ( .A1(n7310), .A2(n7309), .ZN(n4556) );
  INV_X1 U6203 ( .A(n10117), .ZN(n6382) );
  AND2_X1 U6204 ( .A1(n4562), .A2(n4795), .ZN(n10117) );
  OR2_X1 U6205 ( .A1(n9885), .A2(n9889), .ZN(n4557) );
  AND2_X1 U6206 ( .A1(n4542), .A2(n7582), .ZN(n4558) );
  NAND2_X1 U6207 ( .A1(n5201), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4559) );
  AND2_X1 U6208 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4560) );
  NOR2_X1 U6209 ( .A1(n7578), .A2(n8046), .ZN(n4561) );
  OAI21_X1 U6210 ( .B1(n4907), .B2(n4912), .A(n8319), .ZN(n4906) );
  INV_X1 U6211 ( .A(n6498), .ZN(n6231) );
  OR2_X1 U6212 ( .A1(n5307), .A2(n6101), .ZN(n4562) );
  AND2_X1 U6213 ( .A1(n7700), .A2(n6926), .ZN(n4563) );
  AND2_X1 U6214 ( .A1(n5090), .A2(n5089), .ZN(n4564) );
  AND2_X1 U6215 ( .A1(n5092), .A2(n5087), .ZN(n4565) );
  OR2_X1 U6216 ( .A1(n7771), .A2(n7850), .ZN(n4566) );
  INV_X1 U6217 ( .A(n7222), .ZN(n5097) );
  NAND2_X1 U6218 ( .A1(n8050), .A2(n8108), .ZN(n4567) );
  NOR2_X1 U6219 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n4568) );
  AND2_X1 U6220 ( .A1(n4803), .A2(n4802), .ZN(n4569) );
  NAND2_X1 U6221 ( .A1(n7519), .A2(n7518), .ZN(n8505) );
  AND2_X1 U6222 ( .A1(n4780), .A2(n4778), .ZN(n4570) );
  NAND2_X1 U6223 ( .A1(n7771), .A2(n7850), .ZN(n4571) );
  AND2_X1 U6224 ( .A1(n4744), .A2(n4743), .ZN(n4572) );
  OR2_X1 U6225 ( .A1(n5307), .A2(n6035), .ZN(n4573) );
  AND2_X1 U6226 ( .A1(n4528), .A2(n9757), .ZN(n4574) );
  AND2_X1 U6227 ( .A1(n4966), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4575) );
  AND2_X1 U6228 ( .A1(n4975), .A2(n4974), .ZN(n4576) );
  INV_X1 U6229 ( .A(n5138), .ZN(n5109) );
  OR2_X1 U6230 ( .A1(n7825), .A2(n7857), .ZN(n4577) );
  OAI21_X1 U6231 ( .B1(n4838), .B2(n4833), .A(n4836), .ZN(n4832) );
  OR2_X1 U6232 ( .A1(n4871), .A2(n4869), .ZN(n4578) );
  INV_X1 U6233 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6234 ( .A1(n7635), .A2(n4883), .ZN(n4579) );
  OR2_X1 U6235 ( .A1(n4520), .A2(n4938), .ZN(n4580) );
  INV_X1 U6236 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n4745) );
  INV_X1 U6237 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n4931) );
  AND2_X1 U6238 ( .A1(n7250), .A2(n4803), .ZN(n4581) );
  AND2_X1 U6239 ( .A1(n9292), .A2(n4528), .ZN(n4582) );
  OR2_X1 U6240 ( .A1(n6017), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n4583) );
  AND2_X1 U6241 ( .A1(n9856), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4584) );
  INV_X1 U6242 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4726) );
  AND2_X1 U6243 ( .A1(n9837), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4585) );
  NAND2_X1 U6244 ( .A1(n9334), .A2(n8906), .ZN(n9317) );
  NAND2_X1 U6245 ( .A1(n4892), .A2(n7568), .ZN(n8410) );
  INV_X1 U6246 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5057) );
  INV_X1 U6247 ( .A(n7974), .ZN(n5024) );
  OR3_X1 U6248 ( .A1(n6040), .A2(P2_IR_REG_10__SCAN_IN), .A3(n5065), .ZN(n4586) );
  INV_X1 U6249 ( .A(n5241), .ZN(n5877) );
  NAND2_X1 U6250 ( .A1(n7290), .A2(n5123), .ZN(n7605) );
  AND2_X1 U6251 ( .A1(n9757), .A2(n9116), .ZN(n4587) );
  AND2_X1 U6252 ( .A1(n5898), .A2(n7629), .ZN(n4588) );
  AND2_X1 U6253 ( .A1(n5104), .A2(n5102), .ZN(n4589) );
  AND2_X1 U6254 ( .A1(n9763), .A2(n9767), .ZN(n4590) );
  OR2_X1 U6255 ( .A1(n5134), .A2(n5133), .ZN(n4591) );
  AND2_X1 U6256 ( .A1(n4951), .A2(n6980), .ZN(n4592) );
  AND2_X1 U6257 ( .A1(n9787), .A2(n9283), .ZN(n4593) );
  NAND2_X1 U6258 ( .A1(n6078), .A2(n4545), .ZN(n4594) );
  AND2_X1 U6259 ( .A1(n5496), .A2(SI_12_), .ZN(n4595) );
  AND2_X1 U6260 ( .A1(n5709), .A2(SI_21_), .ZN(n4596) );
  INV_X1 U6261 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6275) );
  INV_X1 U6262 ( .A(n7088), .ZN(n6684) );
  INV_X1 U6263 ( .A(n6582), .ZN(n4946) );
  OR2_X1 U6264 ( .A1(n5372), .A2(n4591), .ZN(n4597) );
  INV_X1 U6265 ( .A(n9114), .ZN(n4818) );
  INV_X1 U6266 ( .A(n10299), .ZN(n8381) );
  NAND2_X1 U6267 ( .A1(n7467), .A2(n7466), .ZN(n8360) );
  NAND2_X1 U6268 ( .A1(n5044), .A2(n6055), .ZN(n6271) );
  AND2_X1 U6269 ( .A1(n7068), .A2(n8995), .ZN(n8855) );
  NAND2_X1 U6270 ( .A1(n5385), .A2(n5386), .ZN(n5390) );
  NAND2_X1 U6271 ( .A1(n5265), .A2(n5264), .ZN(n6629) );
  AND2_X1 U6272 ( .A1(n8267), .A2(n4632), .ZN(n4598) );
  AND2_X1 U6273 ( .A1(n8267), .A2(n4625), .ZN(n4599) );
  XNOR2_X1 U6274 ( .A(n5975), .B(n5980), .ZN(n6027) );
  NAND2_X1 U6275 ( .A1(n6835), .A2(n5344), .ZN(n6892) );
  NAND2_X1 U6276 ( .A1(n7056), .A2(n7055), .ZN(n7083) );
  AND2_X1 U6277 ( .A1(n5415), .A2(n5414), .ZN(n4600) );
  NAND2_X1 U6278 ( .A1(n6927), .A2(n4855), .ZN(n7056) );
  AND2_X1 U6279 ( .A1(n4530), .A2(n5070), .ZN(n6800) );
  NAND2_X1 U6280 ( .A1(n4929), .A2(n7749), .ZN(n6923) );
  AND2_X1 U6281 ( .A1(n5012), .A2(n8742), .ZN(n4601) );
  INV_X1 U6282 ( .A(n8121), .ZN(n4980) );
  INV_X1 U6283 ( .A(n8112), .ZN(n5040) );
  CLKBUF_X1 U6284 ( .A(n6535), .Z(n8116) );
  XNOR2_X1 U6285 ( .A(n5177), .B(n5176), .ZN(n9924) );
  AND2_X1 U6286 ( .A1(n6321), .A2(n6320), .ZN(n8096) );
  INV_X1 U6287 ( .A(n8096), .ZN(n8066) );
  AOI22_X1 U6288 ( .A1(n8875), .A2(n6819), .B1(n6731), .B2(n10117), .ZN(n10093) );
  AND2_X1 U6289 ( .A1(n9064), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4602) );
  INV_X1 U6290 ( .A(n10219), .ZN(n4798) );
  NOR2_X1 U6291 ( .A1(n8256), .A2(n4636), .ZN(n4603) );
  INV_X1 U6292 ( .A(n8257), .ZN(n4641) );
  NAND2_X1 U6293 ( .A1(n8195), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4604) );
  INV_X1 U6294 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5146) );
  INV_X1 U6295 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5988) );
  AND2_X1 U6296 ( .A1(n4961), .A2(n4960), .ZN(n4605) );
  INV_X1 U6297 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4670) );
  INV_X1 U6298 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5043) );
  INV_X1 U6299 ( .A(n9223), .ZN(n4786) );
  INV_X1 U6300 ( .A(n6735), .ZN(n8873) );
  OAI21_X1 U6301 ( .B1(n9334), .B2(n9319), .A(n4760), .ZN(n9303) );
  NAND2_X1 U6302 ( .A1(n7011), .A2(n7010), .ZN(n7034) );
  NAND2_X1 U6303 ( .A1(n4859), .A2(n4858), .ZN(n4937) );
  NOR2_X1 U6304 ( .A1(n8097), .A2(n8098), .ZN(n8095) );
  XNOR2_X1 U6305 ( .A(n6479), .B(n8116), .ZN(n6561) );
  INV_X1 U6306 ( .A(n5982), .ZN(n5984) );
  NAND2_X1 U6307 ( .A1(n6507), .A2(n6506), .ZN(n6648) );
  NAND2_X1 U6308 ( .A1(n5044), .A2(n5041), .ZN(n6273) );
  NAND3_X1 U6309 ( .A1(n4606), .A2(n7947), .A3(n8066), .ZN(n7952) );
  NAND2_X1 U6310 ( .A1(n7946), .A2(n7945), .ZN(n4606) );
  NAND2_X1 U6311 ( .A1(n7033), .A2(n5040), .ZN(n5039) );
  INV_X1 U6312 ( .A(n6041), .ZN(n4729) );
  NAND2_X1 U6313 ( .A1(n6027), .A2(n5042), .ZN(n5044) );
  NAND2_X1 U6314 ( .A1(n5974), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5976) );
  NAND2_X1 U6315 ( .A1(n4524), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U6316 ( .A1(n5027), .A2(n5026), .ZN(n7318) );
  NAND2_X1 U6317 ( .A1(n6434), .A2(n6435), .ZN(n5236) );
  XNOR2_X1 U6318 ( .A(n5233), .B(n5232), .ZN(n6435) );
  NAND2_X1 U6319 ( .A1(n5086), .A2(n5085), .ZN(n8641) );
  NOR2_X1 U6320 ( .A1(n9084), .A2(n10032), .ZN(n9082) );
  XNOR2_X1 U6321 ( .A(n9081), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9084) );
  NAND2_X1 U6322 ( .A1(n4611), .A2(n6498), .ZN(n4610) );
  OR2_X1 U6323 ( .A1(n6186), .A2(n10371), .ZN(n4612) );
  OAI211_X1 U6324 ( .C1(n8251), .C2(n4626), .A(n4624), .B(n4616), .ZN(n4617)
         );
  INV_X1 U6325 ( .A(n4617), .ZN(n4638) );
  NAND3_X1 U6326 ( .A1(n4621), .A2(n4618), .A3(n8227), .ZN(n4640) );
  NAND2_X1 U6327 ( .A1(n4623), .A2(n4622), .ZN(n4621) );
  NAND2_X1 U6328 ( .A1(n4640), .A2(n4638), .ZN(P2_U3201) );
  AND2_X2 U6329 ( .A1(n4650), .A2(n4649), .ZN(n5201) );
  NAND3_X1 U6330 ( .A1(n4668), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4649) );
  NAND3_X1 U6331 ( .A1(n4670), .A2(n5168), .A3(n4669), .ZN(n4650) );
  NAND3_X1 U6332 ( .A1(n4658), .A2(n8827), .A3(n4657), .ZN(n4656) );
  NAND3_X1 U6333 ( .A1(n8825), .A2(n8855), .A3(n8824), .ZN(n4657) );
  NAND3_X1 U6334 ( .A1(n8820), .A2(n8819), .A3(n8860), .ZN(n4658) );
  NAND2_X1 U6335 ( .A1(n5250), .A2(n5249), .ZN(n4666) );
  NAND2_X1 U6336 ( .A1(n5222), .A2(n5223), .ZN(n4667) );
  MUX2_X1 U6337 ( .A(n6824), .B(P1_REG2_REG_1__SCAN_IN), .S(n6101), .Z(n9019)
         );
  NAND2_X1 U6338 ( .A1(n5805), .A2(n5804), .ZN(n5807) );
  NAND2_X1 U6339 ( .A1(n5784), .A2(n5783), .ZN(n4706) );
  OR2_X1 U6340 ( .A1(n5644), .A2(n4716), .ZN(n4712) );
  NAND2_X1 U6341 ( .A1(n5644), .A2(n4541), .ZN(n4710) );
  NAND3_X1 U6342 ( .A1(n4763), .A2(n5330), .A3(n4764), .ZN(n4720) );
  INV_X1 U6343 ( .A(n4727), .ZN(n4725) );
  NAND3_X1 U6344 ( .A1(n4727), .A2(n4728), .A3(P2_DATAO_REG_4__SCAN_IN), .ZN(
        n4723) );
  NAND2_X2 U6345 ( .A1(n4729), .A2(n5960), .ZN(n6040) );
  NAND2_X1 U6346 ( .A1(n5964), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6276) );
  NAND2_X1 U6347 ( .A1(n4736), .A2(n7770), .ZN(n4741) );
  NAND2_X1 U6348 ( .A1(n4737), .A2(n7768), .ZN(n4736) );
  NAND3_X1 U6349 ( .A1(n4739), .A2(n4738), .A3(n4742), .ZN(n4737) );
  NAND2_X1 U6350 ( .A1(n7754), .A2(n7857), .ZN(n4738) );
  NAND2_X1 U6351 ( .A1(n7755), .A2(n7850), .ZN(n4739) );
  OAI21_X1 U6352 ( .B1(n4748), .B2(n7818), .A(n4746), .ZN(n7833) );
  MUX2_X1 U6353 ( .A(n6006), .B(n6480), .S(n5201), .Z(n5251) );
  NAND2_X1 U6354 ( .A1(n5202), .A2(n5203), .ZN(n5222) );
  NAND2_X1 U6355 ( .A1(n5277), .A2(n4765), .ZN(n4764) );
  INV_X1 U6356 ( .A(n5301), .ZN(n4768) );
  NAND2_X1 U6357 ( .A1(n4771), .A2(n4774), .ZN(n9233) );
  INV_X1 U6358 ( .A(n9253), .ZN(n4777) );
  NAND3_X1 U6359 ( .A1(n9137), .A2(n9138), .A3(n4777), .ZN(n4776) );
  NAND2_X1 U6360 ( .A1(n9224), .A2(n4785), .ZN(n4784) );
  NOR2_X2 U6361 ( .A1(n9224), .A2(n9225), .ZN(n9223) );
  NOR2_X1 U6362 ( .A1(n9223), .A2(n9141), .ZN(n9211) );
  INV_X2 U6363 ( .A(n5279), .ZN(n5081) );
  NAND3_X1 U6364 ( .A1(n5081), .A2(n4804), .A3(n5080), .ZN(n4790) );
  AND3_X2 U6365 ( .A1(n4793), .A2(n4791), .A3(n5138), .ZN(n5160) );
  CLKBUF_X1 U6366 ( .A(n5140), .Z(n4792) );
  INV_X1 U6367 ( .A(n4792), .ZN(n5165) );
  NOR2_X1 U6368 ( .A1(n5133), .A2(n5134), .ZN(n4793) );
  NAND2_X1 U6369 ( .A1(n5307), .A2(n7631), .ZN(n5304) );
  NAND2_X2 U6370 ( .A1(n5872), .A2(n9924), .ZN(n5307) );
  NAND2_X2 U6371 ( .A1(n5307), .A2(n5201), .ZN(n8745) );
  NAND2_X1 U6372 ( .A1(n7250), .A2(n4569), .ZN(n9326) );
  XNOR2_X1 U6373 ( .A(n6717), .B(n10117), .ZN(n8875) );
  NAND3_X1 U6374 ( .A1(n4807), .A2(n4805), .A3(n4806), .ZN(n5110) );
  INV_X1 U6375 ( .A(n5134), .ZN(n4807) );
  NAND2_X1 U6376 ( .A1(n9259), .A2(n4811), .ZN(n4810) );
  NAND2_X1 U6377 ( .A1(n5140), .A2(n4820), .ZN(n4819) );
  AOI21_X1 U6378 ( .B1(n9200), .B2(n4834), .A(n4832), .ZN(n9156) );
  OAI21_X1 U6379 ( .B1(n9200), .B2(n9121), .A(n9122), .ZN(n9188) );
  INV_X1 U6380 ( .A(n8881), .ZN(n4850) );
  INV_X1 U6381 ( .A(n7942), .ZN(n6303) );
  NAND2_X1 U6382 ( .A1(n6304), .A2(n7942), .ZN(n6501) );
  AOI22_X1 U6383 ( .A1(n6927), .A2(n4853), .B1(n4854), .B2(n7700), .ZN(n7086)
         );
  OR2_X1 U6384 ( .A1(n8374), .A2(n4863), .ZN(n4860) );
  NAND2_X1 U6385 ( .A1(n4860), .A2(n4861), .ZN(n8343) );
  NAND2_X1 U6386 ( .A1(n4865), .A2(n4578), .ZN(n7343) );
  NAND2_X1 U6387 ( .A1(n7290), .A2(n4866), .ZN(n4865) );
  NAND2_X1 U6388 ( .A1(n7583), .A2(n4875), .ZN(n4874) );
  OAI21_X1 U6389 ( .B1(n7583), .B2(n4542), .A(n7582), .ZN(n7628) );
  OAI211_X1 U6390 ( .C1(n7583), .C2(n4876), .A(n10289), .B(n4874), .ZN(n7644)
         );
  NAND2_X1 U6391 ( .A1(n8421), .A2(n4519), .ZN(n4885) );
  OAI21_X1 U6392 ( .B1(n8280), .B2(n8276), .A(n7839), .ZN(n7636) );
  NAND2_X1 U6393 ( .A1(n4921), .A2(n4922), .ZN(n8428) );
  NAND2_X1 U6394 ( .A1(n7281), .A2(n4924), .ZN(n4921) );
  NOR2_X1 U6395 ( .A1(n4515), .A2(n4928), .ZN(n4927) );
  CLKBUF_X1 U6396 ( .A(n4932), .Z(n4930) );
  NAND3_X1 U6397 ( .A1(n4932), .A2(n5958), .A3(n5957), .ZN(n6010) );
  NAND2_X1 U6398 ( .A1(n4930), .A2(n6013), .ZN(n6019) );
  OR2_X1 U6399 ( .A1(n5997), .A2(n4931), .ZN(n6129) );
  OR2_X1 U6400 ( .A1(n5997), .A2(n6432), .ZN(n6132) );
  NAND2_X1 U6401 ( .A1(n4575), .A2(n5997), .ZN(n6127) );
  AND2_X1 U6402 ( .A1(n7766), .A2(n7757), .ZN(n4942) );
  NAND3_X1 U6403 ( .A1(n4943), .A2(P2_REG2_REG_7__SCAN_IN), .A3(n6441), .ZN(
        n4944) );
  NAND2_X1 U6404 ( .A1(n6390), .A2(n6919), .ZN(n6441) );
  INV_X1 U6405 ( .A(n4944), .ZN(n6442) );
  OAI21_X1 U6406 ( .B1(n6583), .B2(n6582), .A(n6684), .ZN(n6669) );
  NAND2_X1 U6407 ( .A1(n4947), .A2(n4945), .ZN(n4948) );
  NAND3_X1 U6408 ( .A1(n4948), .A2(P2_REG2_REG_9__SCAN_IN), .A3(n6669), .ZN(
        n4949) );
  INV_X1 U6409 ( .A(n4949), .ZN(n6670) );
  NAND2_X1 U6410 ( .A1(n6981), .A2(n4955), .ZN(n4950) );
  NAND2_X1 U6411 ( .A1(n4950), .A2(n4952), .ZN(n7197) );
  NAND3_X1 U6412 ( .A1(n4954), .A2(n6980), .A3(n4953), .ZN(n4952) );
  NAND2_X1 U6413 ( .A1(n4954), .A2(n6980), .ZN(n6847) );
  NAND2_X1 U6414 ( .A1(n4956), .A2(n7266), .ZN(n4954) );
  INV_X1 U6415 ( .A(n6846), .ZN(n4956) );
  INV_X1 U6416 ( .A(n6338), .ZN(n4963) );
  NOR2_X1 U6417 ( .A1(n6338), .A2(n4964), .ZN(n6339) );
  NAND2_X1 U6418 ( .A1(n4963), .A2(n6250), .ZN(n6251) );
  INV_X1 U6419 ( .A(n4975), .ZN(n8169) );
  INV_X1 U6420 ( .A(n8168), .ZN(n4974) );
  NAND2_X1 U6421 ( .A1(n8119), .A2(n4980), .ZN(n4977) );
  NAND2_X1 U6422 ( .A1(n4977), .A2(n4976), .ZN(n8144) );
  NAND3_X1 U6423 ( .A1(n4979), .A2(n8117), .A3(n4535), .ZN(n4976) );
  NAND2_X1 U6424 ( .A1(n4979), .A2(n8117), .ZN(n7200) );
  OR2_X1 U6425 ( .A1(n8936), .A2(n4982), .ZN(n4981) );
  MUX2_X1 U6426 ( .A(n6775), .B(n6008), .S(n7631), .Z(n5332) );
  MUX2_X1 U6427 ( .A(n6918), .B(n6024), .S(n7631), .Z(n5376) );
  MUX2_X1 U6428 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7631), .Z(n5537) );
  MUX2_X1 U6429 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n7631), .Z(n5540) );
  MUX2_X1 U6430 ( .A(n9499), .B(n6529), .S(n7631), .Z(n5543) );
  MUX2_X1 U6431 ( .A(n6626), .B(n6637), .S(n7631), .Z(n5596) );
  MUX2_X1 U6432 ( .A(n6716), .B(n5620), .S(n7631), .Z(n5640) );
  MUX2_X1 U6433 ( .A(n6816), .B(n6817), .S(n7631), .Z(n5645) );
  MUX2_X1 U6434 ( .A(n9367), .B(n6902), .S(n7631), .Z(n5671) );
  MUX2_X1 U6435 ( .A(n7477), .B(n6961), .S(n7631), .Z(n5708) );
  MUX2_X1 U6436 ( .A(n7489), .B(n9604), .S(n7631), .Z(n5712) );
  MUX2_X1 U6437 ( .A(n7500), .B(n7070), .S(n7631), .Z(n5731) );
  MUX2_X1 U6438 ( .A(n7508), .B(n7219), .S(n7631), .Z(n5757) );
  MUX2_X1 U6439 ( .A(n7517), .B(n7244), .S(n7631), .Z(n5787) );
  MUX2_X1 U6440 ( .A(n8579), .B(n9818), .S(n7631), .Z(n5809) );
  MUX2_X1 U6441 ( .A(n7542), .B(n9815), .S(n7631), .Z(n5895) );
  INV_X1 U6442 ( .A(n5359), .ZN(n4995) );
  OAI21_X1 U6443 ( .B1(n4995), .B2(n4998), .A(n4996), .ZN(n5406) );
  INV_X1 U6444 ( .A(n5011), .ZN(n7656) );
  NAND2_X1 U6445 ( .A1(n5014), .A2(n8741), .ZN(n9091) );
  NAND2_X1 U6446 ( .A1(n6648), .A2(n5015), .ZN(n5018) );
  INV_X1 U6447 ( .A(n5018), .ZN(n6789) );
  NAND2_X1 U6448 ( .A1(n7895), .A2(n5020), .ZN(n5019) );
  NAND2_X1 U6449 ( .A1(n7034), .A2(n5029), .ZN(n5027) );
  XNOR2_X1 U6450 ( .A(n6026), .B(P2_B_REG_SCAN_IN), .ZN(n5042) );
  NAND2_X1 U6451 ( .A1(n8006), .A2(n5048), .ZN(n5045) );
  NAND2_X1 U6452 ( .A1(n5045), .A2(n5046), .ZN(n7886) );
  INV_X1 U6453 ( .A(n6010), .ZN(n5054) );
  NAND2_X1 U6454 ( .A1(n5054), .A2(n5055), .ZN(n6041) );
  NOR3_X1 U6455 ( .A1(n6010), .A2(P2_IR_REG_7__SCAN_IN), .A3(
        P2_IR_REG_6__SCAN_IN), .ZN(n6030) );
  OAI21_X1 U6456 ( .B1(n8078), .B2(n5061), .A(n5058), .ZN(n7922) );
  NAND2_X1 U6457 ( .A1(n8078), .A2(n8079), .ZN(n5064) );
  AND2_X2 U6458 ( .A1(n6800), .A2(n6799), .ZN(n6802) );
  AND2_X1 U6459 ( .A1(n5069), .A2(n5068), .ZN(n6799) );
  NAND3_X1 U6460 ( .A1(n5265), .A2(n5071), .A3(n5264), .ZN(n5069) );
  NAND3_X1 U6461 ( .A1(n5265), .A2(n5264), .A3(n5072), .ZN(n5070) );
  NOR2_X1 U6462 ( .A1(n6630), .A2(n5321), .ZN(n5071) );
  NOR2_X1 U6463 ( .A1(n6630), .A2(n5315), .ZN(n5072) );
  NAND2_X1 U6464 ( .A1(n6834), .A2(n5074), .ZN(n5073) );
  NAND3_X1 U6465 ( .A1(n5084), .A2(n5727), .A3(n8607), .ZN(n8606) );
  NAND2_X1 U6466 ( .A1(n5084), .A2(n8607), .ZN(n8691) );
  NAND2_X1 U6467 ( .A1(n7396), .A2(n4565), .ZN(n5086) );
  NAND3_X1 U6468 ( .A1(n5390), .A2(n5096), .A3(n5389), .ZN(n5095) );
  NAND2_X1 U6469 ( .A1(n5390), .A2(n5389), .ZN(n7137) );
  INV_X1 U6470 ( .A(n7136), .ZN(n5096) );
  OAI21_X2 U6471 ( .B1(n8713), .B2(n5101), .A(n5098), .ZN(n8627) );
  NAND2_X1 U6472 ( .A1(n5160), .A2(n5108), .ZN(n5173) );
  OR2_X1 U6473 ( .A1(n6500), .A2(n6432), .ZN(n6311) );
  OR2_X1 U6474 ( .A1(n6500), .A2(n6601), .ZN(n6307) );
  OR2_X1 U6475 ( .A1(n6499), .A2(n6563), .ZN(n6305) );
  NAND2_X1 U6476 ( .A1(n6476), .A2(n5201), .ZN(n6492) );
  OAI21_X1 U6477 ( .B1(n5859), .B2(n5858), .A(n5857), .ZN(n5889) );
  NAND2_X2 U6478 ( .A1(n6295), .A2(n6124), .ZN(n6476) );
  NAND2_X1 U6479 ( .A1(n5940), .A2(n5117), .ZN(n5956) );
  NAND2_X1 U6480 ( .A1(n5240), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5217) );
  XNOR2_X1 U6481 ( .A(n5207), .B(n5532), .ZN(n5210) );
  NAND2_X2 U6482 ( .A1(n7912), .A2(n7911), .ZN(n8078) );
  INV_X1 U6483 ( .A(n6547), .ZN(n6615) );
  NAND2_X1 U6484 ( .A1(n5173), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5175) );
  OAI21_X1 U6485 ( .B1(n5173), .B2(P1_IR_REG_28__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5142) );
  AND2_X1 U6486 ( .A1(n8586), .A2(n8680), .ZN(n5857) );
  AND2_X1 U6487 ( .A1(n7363), .A2(n7362), .ZN(n10369) );
  AND2_X1 U6488 ( .A1(n6315), .A2(n6271), .ZN(n6050) );
  AND3_X2 U6489 ( .A1(n6558), .A2(n6557), .A3(n6556), .ZN(n10386) );
  AND2_X1 U6490 ( .A1(n7534), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5111) );
  INV_X1 U6491 ( .A(n6536), .ZN(n6313) );
  AND2_X1 U6492 ( .A1(n6975), .A2(n6971), .ZN(n5112) );
  AND2_X1 U6493 ( .A1(n7316), .A2(n8107), .ZN(n5113) );
  OR2_X1 U6494 ( .A1(n9723), .A2(n9715), .ZN(n5114) );
  INV_X1 U6495 ( .A(n8345), .ZN(n8378) );
  AND4_X1 U6496 ( .A1(n7475), .A2(n7474), .A3(n7473), .A4(n7472), .ZN(n8345)
         );
  INV_X1 U6497 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6279) );
  AND3_X1 U6498 ( .A1(n5939), .A2(n8680), .A3(n5938), .ZN(n5117) );
  OR2_X1 U6499 ( .A1(n10367), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5118) );
  AND2_X1 U6500 ( .A1(n6192), .A2(n6231), .ZN(n5119) );
  AND2_X1 U6501 ( .A1(n5965), .A2(n5963), .ZN(n5120) );
  AND4_X1 U6502 ( .A1(n7486), .A2(n7485), .A3(n7484), .A4(n7483), .ZN(n7897)
         );
  AND2_X1 U6503 ( .A1(n5416), .A2(n5405), .ZN(n5121) );
  NOR2_X1 U6504 ( .A1(n8855), .A2(n8927), .ZN(n8743) );
  INV_X1 U6505 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n6298) );
  AND2_X1 U6506 ( .A1(n5294), .A2(n5293), .ZN(n5122) );
  OR2_X1 U6507 ( .A1(n7305), .A2(n8109), .ZN(n5123) );
  NAND2_X1 U6508 ( .A1(n6723), .A2(n9306), .ZN(n9309) );
  AND3_X1 U6509 ( .A1(n5942), .A2(n5941), .A3(n8680), .ZN(n5124) );
  INV_X1 U6510 ( .A(n7896), .ZN(n8530) );
  NAND2_X1 U6511 ( .A1(n7688), .A2(n7684), .ZN(n7843) );
  NAND2_X1 U6512 ( .A1(n8760), .A2(n8759), .ZN(n8774) );
  INV_X1 U6513 ( .A(n9094), .ZN(n8742) );
  NOR2_X1 U6514 ( .A1(n8928), .A2(n8749), .ZN(n8750) );
  AND4_X1 U6515 ( .A1(n5137), .A2(n5136), .A3(n5135), .A4(n5181), .ZN(n5138)
         );
  INV_X1 U6516 ( .A(n7897), .ZN(n7576) );
  AND2_X1 U6517 ( .A1(n10078), .A2(n5580), .ZN(n5288) );
  AND2_X1 U6518 ( .A1(n7026), .A2(n8783), .ZN(n8768) );
  INV_X1 U6519 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5178) );
  NOR2_X1 U6520 ( .A1(n7308), .A2(n7982), .ZN(n7309) );
  INV_X1 U6521 ( .A(n7933), .ZN(n6304) );
  INV_X1 U6522 ( .A(n7843), .ZN(n7635) );
  NAND2_X1 U6523 ( .A1(n7574), .A2(n8345), .ZN(n7575) );
  INV_X1 U6524 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7282) );
  INV_X1 U6525 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6653) );
  NOR2_X1 U6526 ( .A1(n7896), .A2(n7576), .ZN(n7577) );
  OR2_X1 U6527 ( .A1(n8113), .A2(n10330), .ZN(n7749) );
  INV_X1 U6528 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5993) );
  INV_X1 U6529 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6411) );
  NAND2_X1 U6530 ( .A1(n6632), .A2(n5580), .ZN(n5309) );
  INV_X1 U6531 ( .A(n8857), .ZN(n8858) );
  INV_X1 U6532 ( .A(n5526), .ZN(n5525) );
  INV_X1 U6533 ( .A(SI_19_), .ZN(n9668) );
  AND2_X1 U6534 ( .A1(n7007), .A2(n8113), .ZN(n7008) );
  NAND2_X1 U6535 ( .A1(n7075), .A2(n7074), .ZN(n7157) );
  NAND2_X1 U6536 ( .A1(n7694), .A2(n6538), .ZN(n6612) );
  INV_X1 U6537 ( .A(n8312), .ZN(n7909) );
  INV_X1 U6538 ( .A(n8261), .ZN(n7455) );
  AOI21_X1 U6539 ( .B1(n6875), .B2(n6874), .A(n6873), .ZN(n6877) );
  OR2_X1 U6540 ( .A1(n7850), .A2(n6469), .ZN(n7359) );
  INV_X1 U6541 ( .A(n8716), .ZN(n5634) );
  INV_X1 U6542 ( .A(n5386), .ZN(n5387) );
  OAI21_X1 U6543 ( .B1(n5466), .B2(n8704), .A(n5465), .ZN(n5467) );
  INV_X1 U6544 ( .A(n8692), .ZN(n5727) );
  OR2_X1 U6545 ( .A1(n5676), .A2(n9461), .ZN(n5694) );
  NAND2_X1 U6546 ( .A1(n5525), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5571) );
  INV_X1 U6547 ( .A(n9128), .ZN(n9146) );
  INV_X1 U6548 ( .A(n5627), .ZN(n5625) );
  INV_X1 U6549 ( .A(n5190), .ZN(n6724) );
  INV_X1 U6550 ( .A(n10194), .ZN(n10234) );
  INV_X1 U6551 ( .A(n9285), .ZN(n9778) );
  INV_X1 U6552 ( .A(n10091), .ZN(n10095) );
  INV_X1 U6553 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5174) );
  NAND2_X1 U6554 ( .A1(n5596), .A2(n5595), .ZN(n5619) );
  OR2_X1 U6555 ( .A1(n5521), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5522) );
  OR2_X1 U6556 ( .A1(n5427), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5476) );
  OR2_X1 U6557 ( .A1(n7545), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n7556) );
  AOI21_X1 U6558 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8145), .A(n8144), .ZN(
        n8166) );
  OR2_X1 U6559 ( .A1(n7532), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n7545) );
  INV_X1 U6560 ( .A(n8377), .ZN(n8392) );
  OR2_X1 U6561 ( .A1(n10356), .A2(n6548), .ZN(n6552) );
  AND2_X1 U6562 ( .A1(n6316), .A2(n6315), .ZN(n6423) );
  OR3_X1 U6563 ( .A1(n8376), .A2(n8375), .A3(n10301), .ZN(n8380) );
  INV_X1 U6564 ( .A(n8107), .ZN(n7609) );
  AND2_X1 U6565 ( .A1(n7748), .A2(n7744), .ZN(n7696) );
  INV_X1 U6566 ( .A(n10289), .ZN(n10301) );
  INV_X1 U6567 ( .A(n5467), .ZN(n5468) );
  OR2_X1 U6568 ( .A1(n5589), .A2(n5588), .ZN(n5590) );
  INV_X1 U6569 ( .A(n5462), .ZN(n8702) );
  INV_X1 U6570 ( .A(n8693), .ZN(n8729) );
  INV_X1 U6571 ( .A(n8933), .ZN(n8992) );
  INV_X1 U6572 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7388) );
  OR2_X1 U6573 ( .A1(n9933), .A2(n9024), .ZN(n10032) );
  AND3_X1 U6574 ( .A1(n6075), .A2(n6074), .A3(n6073), .ZN(n9149) );
  INV_X1 U6575 ( .A(n9754), .ZN(n9206) );
  INV_X1 U6576 ( .A(n9103), .ZN(n9907) );
  INV_X1 U6577 ( .A(n9897), .ZN(n10237) );
  OR2_X1 U6578 ( .A1(n10053), .A2(n10184), .ZN(n6965) );
  INV_X1 U6579 ( .A(n8931), .ZN(n5882) );
  INV_X1 U6580 ( .A(n9736), .ZN(n9195) );
  INV_X1 U6581 ( .A(n9874), .ZN(n9885) );
  OR3_X1 U6582 ( .A1(n7259), .A2(n7258), .A3(n10222), .ZN(n10242) );
  AND2_X1 U6583 ( .A1(n8953), .A2(n8956), .ZN(n7103) );
  INV_X1 U6584 ( .A(n7409), .ZN(n6169) );
  AND2_X1 U6585 ( .A1(n5892), .A2(n5811), .ZN(n5890) );
  INV_X1 U6586 ( .A(SI_6_), .ZN(n9498) );
  NAND2_X1 U6587 ( .A1(n5986), .A2(n5985), .ZN(n6287) );
  AND2_X1 U6588 ( .A1(n6296), .A2(n6508), .ZN(n8092) );
  AND2_X1 U6589 ( .A1(n6293), .A2(n6292), .ZN(n8094) );
  AND4_X1 U6590 ( .A1(n7442), .A2(n7441), .A3(n7440), .A4(n7439), .ZN(n8071)
         );
  AND2_X1 U6591 ( .A1(n6141), .A2(n6142), .ZN(n10280) );
  INV_X1 U6592 ( .A(n10283), .ZN(n8202) );
  INV_X1 U6593 ( .A(n8264), .ZN(n10279) );
  AND2_X1 U6594 ( .A1(n10280), .A2(n8255), .ZN(n8267) );
  OR2_X1 U6595 ( .A1(n10356), .A2(n6283), .ZN(n8308) );
  INV_X1 U6596 ( .A(n8470), .ZN(n8486) );
  AND3_X1 U6597 ( .A1(n6424), .A2(n6423), .A3(n6422), .ZN(n6557) );
  INV_X1 U6598 ( .A(n7829), .ZN(n8287) );
  AND2_X1 U6599 ( .A1(n8380), .A2(n8379), .ZN(n8536) );
  NAND2_X1 U6600 ( .A1(n10309), .A2(n10351), .ZN(n10345) );
  INV_X1 U6601 ( .A(n10356), .ZN(n10366) );
  INV_X1 U6602 ( .A(n5952), .ZN(n5953) );
  INV_X1 U6603 ( .A(n8696), .ZN(n8725) );
  NAND2_X1 U6604 ( .A1(n9306), .A2(n5861), .ZN(n8731) );
  OR2_X1 U6605 ( .A1(n9161), .A2(n5943), .ZN(n5931) );
  INV_X1 U6606 ( .A(n10032), .ZN(n9988) );
  INV_X1 U6607 ( .A(n9086), .ZN(n8995) );
  AND2_X1 U6608 ( .A1(n8861), .A2(n8737), .ZN(n10222) );
  OAI21_X1 U6609 ( .B1(n10055), .B2(n10054), .A(n6965), .ZN(n7020) );
  INV_X1 U6610 ( .A(n10236), .ZN(n10191) );
  INV_X1 U6611 ( .A(n9339), .ZN(n10097) );
  NOR2_X1 U6612 ( .A1(n6173), .A2(n6720), .ZN(n6174) );
  INV_X1 U6613 ( .A(n10231), .ZN(n10198) );
  INV_X1 U6614 ( .A(n10222), .ZN(n10203) );
  NAND2_X1 U6615 ( .A1(n5839), .A2(n5840), .ZN(n6057) );
  NOR2_X1 U6616 ( .A1(n6287), .A2(n7071), .ZN(n6143) );
  INV_X1 U6617 ( .A(n8101), .ZN(n8076) );
  INV_X1 U6618 ( .A(n8103), .ZN(n8270) );
  INV_X1 U6619 ( .A(n8346), .ZN(n8327) );
  INV_X1 U6620 ( .A(n8391), .ZN(n8412) );
  INV_X1 U6621 ( .A(P2_U3893), .ZN(n8236) );
  OR2_X1 U6622 ( .A1(P2_U3150), .A2(n6143), .ZN(n8204) );
  OR2_X1 U6623 ( .A1(n6136), .A2(n8255), .ZN(n8268) );
  NAND2_X1 U6624 ( .A1(n6430), .A2(n8430), .ZN(n10299) );
  OR2_X1 U6625 ( .A1(n6430), .A2(n8308), .ZN(n8361) );
  INV_X1 U6626 ( .A(n10386), .ZN(n10384) );
  OR2_X1 U6627 ( .A1(n10369), .A2(n10361), .ZN(n8555) );
  INV_X2 U6628 ( .A(n10369), .ZN(n10367) );
  INV_X1 U6629 ( .A(n6050), .ZN(n6036) );
  INV_X1 U6630 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7517) );
  INV_X1 U6631 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6816) );
  INV_X1 U6632 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6064) );
  INV_X1 U6633 ( .A(n9243), .ZN(n9757) );
  NOR2_X1 U6634 ( .A1(n5124), .A2(n5953), .ZN(n5954) );
  INV_X1 U6635 ( .A(n9750), .ZN(n9221) );
  INV_X1 U6636 ( .A(n8731), .ZN(n8689) );
  AND2_X1 U6637 ( .A1(n6183), .A2(n9007), .ZN(n8696) );
  AND3_X1 U6638 ( .A1(n6070), .A2(n6069), .A3(n6068), .ZN(n9094) );
  NAND2_X1 U6639 ( .A1(n5770), .A2(n5769), .ZN(n9754) );
  INV_X1 U6640 ( .A(n9945), .ZN(n10046) );
  OR2_X1 U6641 ( .A1(n4495), .A2(n10222), .ZN(n9353) );
  INV_X1 U6642 ( .A(n10274), .ZN(n10272) );
  AND2_X2 U6643 ( .A1(n6722), .A2(n6174), .ZN(n10274) );
  INV_X1 U6644 ( .A(n10251), .ZN(n10249) );
  INV_X1 U6645 ( .A(n10113), .ZN(n10115) );
  INV_X1 U6646 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7244) );
  INV_X1 U6647 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6961) );
  INV_X1 U6648 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6121) );
  INV_X1 U6649 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6039) );
  AND2_X1 U6650 ( .A1(n6143), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3893) );
  NAND2_X1 U6651 ( .A1(n5889), .A2(n5888), .ZN(P1_U3240) );
  NAND4_X1 U6652 ( .A1(n5498), .A2(n5130), .A3(n5474), .A4(n5566), .ZN(n5134)
         );
  NOR2_X1 U6653 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5137) );
  NOR2_X1 U6654 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5136) );
  NOR2_X1 U6655 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5135) );
  INV_X1 U6656 ( .A(n5145), .ZN(n5144) );
  INV_X1 U6657 ( .A(n5149), .ZN(n5148) );
  NAND2_X1 U6658 ( .A1(n5240), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U6659 ( .A1(n5238), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5153) );
  NAND2_X1 U6660 ( .A1(n5237), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U6661 ( .A1(n5241), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5151) );
  NAND2_X1 U6662 ( .A1(n5600), .A2(n9386), .ZN(n5621) );
  NOR2_X2 U6663 ( .A1(n5621), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U6664 ( .A1(n5184), .A2(n5186), .ZN(n5157) );
  INV_X1 U6665 ( .A(n5179), .ZN(n5155) );
  NAND2_X1 U6666 ( .A1(n5157), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5159) );
  INV_X1 U6667 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5158) );
  XNOR2_X2 U6668 ( .A(n5159), .B(n5158), .ZN(n6904) );
  INV_X1 U6669 ( .A(n5160), .ZN(n5161) );
  NAND2_X1 U6670 ( .A1(n5163), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5164) );
  NAND2_X1 U6671 ( .A1(n5165), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5166) );
  INV_X2 U6672 ( .A(n5125), .ZN(n5829) );
  INV_X1 U6673 ( .A(SI_0_), .ZN(n5170) );
  INV_X1 U6674 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5169) );
  OAI21_X1 U6675 ( .B1(n5201), .B2(n5170), .A(n5169), .ZN(n5172) );
  AND2_X1 U6676 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5171) );
  AND2_X1 U6677 ( .A1(n5172), .A2(n5203), .ZN(n9823) );
  XNOR2_X2 U6678 ( .A(n5175), .B(n5174), .ZN(n5872) );
  MUX2_X1 U6679 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9823), .S(n5307), .Z(n6827) );
  NAND2_X1 U6680 ( .A1(n5179), .A2(n5178), .ZN(n5180) );
  OR2_X1 U6681 ( .A1(n5182), .A2(n5181), .ZN(n5183) );
  INV_X1 U6682 ( .A(n5184), .ZN(n5185) );
  NAND2_X1 U6683 ( .A1(n5185), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U6684 ( .A1(n9005), .A2(n9086), .ZN(n6164) );
  NAND2_X1 U6685 ( .A1(n5190), .A2(n6163), .ZN(n5188) );
  NAND2_X1 U6686 ( .A1(n6164), .A2(n5188), .ZN(n5189) );
  NAND2_X2 U6687 ( .A1(n5189), .A2(n5996), .ZN(n5905) );
  NAND3_X1 U6688 ( .A1(n6164), .A2(n5996), .A3(n5190), .ZN(n5559) );
  AND2_X1 U6689 ( .A1(n6827), .A2(n5256), .ZN(n5191) );
  AOI21_X1 U6690 ( .B1(n10121), .B2(n5829), .A(n5191), .ZN(n5195) );
  NAND2_X1 U6691 ( .A1(n5836), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6692 ( .A1(n5195), .A2(n5192), .ZN(n6178) );
  INV_X4 U6693 ( .A(n5905), .ZN(n5935) );
  NAND2_X1 U6694 ( .A1(n10121), .A2(n5935), .ZN(n5194) );
  AOI22_X1 U6695 ( .A1(n6827), .A2(n5829), .B1(n5836), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5193) );
  NAND2_X1 U6696 ( .A1(n5194), .A2(n5193), .ZN(n6177) );
  NAND2_X1 U6697 ( .A1(n6178), .A2(n6177), .ZN(n6180) );
  NAND2_X1 U6698 ( .A1(n5195), .A2(n5773), .ZN(n5196) );
  NAND2_X1 U6699 ( .A1(n5237), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U6700 ( .A1(n5241), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6701 ( .A1(n5240), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5197) );
  NAND4_X2 U6702 ( .A1(n5200), .A2(n5199), .A3(n5198), .A4(n5197), .ZN(n6717)
         );
  NAND2_X1 U6703 ( .A1(n6717), .A2(n5829), .ZN(n5206) );
  XNOR2_X1 U6704 ( .A(n5224), .B(SI_1_), .ZN(n5221) );
  NAND3_X1 U6705 ( .A1(n5201), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n5202) );
  XNOR2_X1 U6706 ( .A(n5221), .B(n5222), .ZN(n6473) );
  INV_X1 U6707 ( .A(n6473), .ZN(n6003) );
  INV_X1 U6708 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6004) );
  INV_X1 U6709 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5204) );
  NAND2_X1 U6710 ( .A1(n6382), .A2(n5256), .ZN(n5205) );
  NAND2_X1 U6711 ( .A1(n5206), .A2(n5205), .ZN(n5207) );
  BUF_X1 U6712 ( .A(n5559), .Z(n5532) );
  AND2_X1 U6713 ( .A1(n6717), .A2(n5935), .ZN(n5209) );
  AND2_X1 U6714 ( .A1(n6382), .A2(n5829), .ZN(n5208) );
  NOR2_X1 U6715 ( .A1(n5209), .A2(n5208), .ZN(n5211) );
  XNOR2_X1 U6716 ( .A(n5210), .B(n5211), .ZN(n6378) );
  NAND2_X1 U6717 ( .A1(n6380), .A2(n6378), .ZN(n6379) );
  INV_X1 U6718 ( .A(n5210), .ZN(n5212) );
  NAND2_X1 U6719 ( .A1(n5212), .A2(n5211), .ZN(n5213) );
  NAND2_X1 U6720 ( .A1(n6379), .A2(n5213), .ZN(n6434) );
  NAND2_X1 U6721 ( .A1(n5238), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U6722 ( .A1(n5237), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5215) );
  NAND2_X1 U6723 ( .A1(n5241), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U6724 ( .A1(n9013), .A2(n5829), .ZN(n5229) );
  OR2_X1 U6725 ( .A1(n5218), .A2(n5599), .ZN(n5220) );
  INV_X1 U6726 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5219) );
  NAND2_X1 U6727 ( .A1(n5220), .A2(n5219), .ZN(n5246) );
  INV_X1 U6728 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6006) );
  INV_X1 U6729 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6480) );
  INV_X1 U6730 ( .A(n5221), .ZN(n5223) );
  NAND2_X1 U6731 ( .A1(n5224), .A2(SI_1_), .ZN(n5225) );
  XNOR2_X1 U6732 ( .A(n5249), .B(n5250), .ZN(n6481) );
  OR2_X1 U6733 ( .A1(n5304), .A2(n6481), .ZN(n5226) );
  OAI211_X2 U6734 ( .C1(n5307), .C2(n6100), .A(n5227), .B(n5226), .ZN(n10091)
         );
  NAND2_X1 U6735 ( .A1(n10091), .A2(n5256), .ZN(n5228) );
  NAND2_X1 U6736 ( .A1(n5229), .A2(n5228), .ZN(n5230) );
  BUF_X1 U6737 ( .A(n5559), .Z(n5511) );
  XNOR2_X1 U6738 ( .A(n5230), .B(n5511), .ZN(n5232) );
  AND2_X1 U6739 ( .A1(n10091), .A2(n5829), .ZN(n5231) );
  AOI21_X1 U6740 ( .B1(n9013), .B2(n5935), .A(n5231), .ZN(n5233) );
  INV_X1 U6741 ( .A(n5232), .ZN(n5234) );
  NAND2_X1 U6742 ( .A1(n5234), .A2(n5233), .ZN(n5235) );
  NAND2_X1 U6743 ( .A1(n5236), .A2(n5235), .ZN(n6575) );
  NAND2_X1 U6744 ( .A1(n5237), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5245) );
  INV_X1 U6745 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6746 ( .A1(n5238), .A2(n5239), .ZN(n5244) );
  NAND2_X1 U6747 ( .A1(n5240), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U6748 ( .A1(n5241), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5242) );
  NAND2_X1 U6749 ( .A1(n10089), .A2(n5580), .ZN(n5258) );
  NAND2_X1 U6750 ( .A1(n5246), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5248) );
  INV_X1 U6751 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5247) );
  XNOR2_X1 U6752 ( .A(n5248), .B(n5247), .ZN(n6104) );
  INV_X1 U6753 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6005) );
  OR2_X1 U6754 ( .A1(n8745), .A2(n6005), .ZN(n5255) );
  INV_X1 U6755 ( .A(n5251), .ZN(n5252) );
  NAND2_X1 U6756 ( .A1(n5252), .A2(SI_2_), .ZN(n5253) );
  INV_X1 U6757 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6495) );
  MUX2_X1 U6758 ( .A(n6495), .B(n6005), .S(n7631), .Z(n5274) );
  XNOR2_X1 U6759 ( .A(n5274), .B(SI_3_), .ZN(n5272) );
  XNOR2_X1 U6760 ( .A(n5273), .B(n5272), .ZN(n6493) );
  OR2_X1 U6761 ( .A1(n5304), .A2(n6493), .ZN(n5254) );
  OAI211_X1 U6762 ( .C1(n5307), .C2(n6104), .A(n5255), .B(n5254), .ZN(n6718)
         );
  NAND2_X1 U6763 ( .A1(n6718), .A2(n5903), .ZN(n5257) );
  NAND2_X1 U6764 ( .A1(n5258), .A2(n5257), .ZN(n5259) );
  XNOR2_X1 U6765 ( .A(n5259), .B(n5532), .ZN(n5261) );
  AND2_X1 U6766 ( .A1(n6718), .A2(n5829), .ZN(n5260) );
  AOI21_X1 U6767 ( .B1(n10089), .B2(n5935), .A(n5260), .ZN(n5262) );
  XNOR2_X1 U6768 ( .A(n5261), .B(n5262), .ZN(n6576) );
  INV_X1 U6769 ( .A(n5261), .ZN(n5263) );
  NAND2_X1 U6770 ( .A1(n5263), .A2(n5262), .ZN(n5264) );
  NAND2_X1 U6771 ( .A1(n5241), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6772 ( .A1(n5237), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5270) );
  INV_X1 U6773 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5266) );
  XNOR2_X1 U6774 ( .A(n5266), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n10077) );
  NAND2_X1 U6775 ( .A1(n5238), .A2(n10077), .ZN(n5269) );
  INV_X1 U6776 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5267) );
  NAND2_X1 U6777 ( .A1(n5287), .A2(n5580), .ZN(n5285) );
  INV_X1 U6778 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6007) );
  OR2_X1 U6779 ( .A1(n8745), .A2(n6007), .ZN(n5283) );
  NAND2_X1 U6780 ( .A1(n5273), .A2(n5272), .ZN(n5277) );
  INV_X1 U6781 ( .A(n5274), .ZN(n5275) );
  NAND2_X1 U6782 ( .A1(n5275), .A2(SI_3_), .ZN(n5276) );
  INV_X1 U6783 ( .A(SI_4_), .ZN(n5278) );
  XNOR2_X1 U6784 ( .A(n5303), .B(n5278), .ZN(n5301) );
  XNOR2_X1 U6785 ( .A(n5302), .B(n5301), .ZN(n6639) );
  NAND2_X1 U6786 ( .A1(n5279), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5280) );
  MUX2_X1 U6787 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5280), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5282) );
  NAND2_X1 U6788 ( .A1(n5282), .A2(n5281), .ZN(n6106) );
  NAND2_X1 U6789 ( .A1(n10078), .A2(n5903), .ZN(n5284) );
  NAND2_X1 U6790 ( .A1(n5285), .A2(n5284), .ZN(n5286) );
  XNOR2_X1 U6791 ( .A(n5286), .B(n5773), .ZN(n5311) );
  AOI21_X1 U6792 ( .B1(n5287), .B2(n5935), .A(n5288), .ZN(n5312) );
  XNOR2_X1 U6793 ( .A(n5311), .B(n5312), .ZN(n6630) );
  NAND2_X1 U6794 ( .A1(n5240), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5296) );
  NAND3_X1 U6795 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5323) );
  INV_X1 U6796 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6797 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5290) );
  NAND2_X1 U6798 ( .A1(n5291), .A2(n5290), .ZN(n5292) );
  AND2_X1 U6799 ( .A1(n5323), .A2(n5292), .ZN(n6813) );
  NAND2_X1 U6800 ( .A1(n5238), .A2(n6813), .ZN(n5294) );
  NAND2_X1 U6801 ( .A1(n5237), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6802 ( .A1(n5241), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5295) );
  NAND2_X1 U6803 ( .A1(n5281), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5297) );
  MUX2_X1 U6804 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5297), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5300) );
  INV_X1 U6805 ( .A(n5298), .ZN(n5299) );
  AND2_X1 U6806 ( .A1(n5300), .A2(n5299), .ZN(n9953) );
  INV_X1 U6807 ( .A(n9953), .ZN(n6092) );
  XNOR2_X1 U6808 ( .A(n5332), .B(SI_5_), .ZN(n5330) );
  XNOR2_X1 U6809 ( .A(n5331), .B(n5330), .ZN(n6774) );
  OR2_X1 U6810 ( .A1(n5304), .A2(n6774), .ZN(n5306) );
  OR2_X1 U6811 ( .A1(n8745), .A2(n6008), .ZN(n5305) );
  OAI211_X1 U6812 ( .C1(n5307), .C2(n6092), .A(n5306), .B(n5305), .ZN(n10153)
         );
  NAND2_X1 U6813 ( .A1(n10153), .A2(n5903), .ZN(n5308) );
  NAND2_X1 U6814 ( .A1(n5309), .A2(n5308), .ZN(n5310) );
  XNOR2_X1 U6815 ( .A(n5310), .B(n5532), .ZN(n6804) );
  INV_X1 U6816 ( .A(n6804), .ZN(n5315) );
  INV_X1 U6817 ( .A(n5311), .ZN(n5314) );
  INV_X1 U6818 ( .A(n5312), .ZN(n5313) );
  NAND2_X1 U6819 ( .A1(n5314), .A2(n5313), .ZN(n5318) );
  NAND2_X1 U6820 ( .A1(n6632), .A2(n5935), .ZN(n5317) );
  NAND2_X1 U6821 ( .A1(n10153), .A2(n5580), .ZN(n5316) );
  NAND2_X1 U6822 ( .A1(n5317), .A2(n5316), .ZN(n6808) );
  INV_X1 U6823 ( .A(n6808), .ZN(n5321) );
  INV_X1 U6824 ( .A(n5318), .ZN(n5319) );
  NOR2_X1 U6825 ( .A1(n6804), .A2(n5319), .ZN(n5320) );
  NAND2_X1 U6826 ( .A1(n5241), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5328) );
  NAND2_X1 U6827 ( .A1(n6067), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5327) );
  INV_X1 U6828 ( .A(n5323), .ZN(n5322) );
  NAND2_X1 U6829 ( .A1(n5322), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5347) );
  INV_X1 U6830 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9601) );
  NAND2_X1 U6831 ( .A1(n5323), .A2(n9601), .ZN(n5324) );
  AND2_X1 U6832 ( .A1(n5347), .A2(n5324), .ZN(n10066) );
  NAND2_X1 U6833 ( .A1(n5238), .A2(n10066), .ZN(n5326) );
  NAND2_X1 U6834 ( .A1(n6072), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5325) );
  NAND4_X1 U6835 ( .A1(n5328), .A2(n5327), .A3(n5326), .A4(n5325), .ZN(n10166)
         );
  NAND2_X1 U6836 ( .A1(n10166), .A2(n5580), .ZN(n5338) );
  OR2_X1 U6837 ( .A1(n5298), .A2(n5599), .ZN(n5329) );
  XNOR2_X1 U6838 ( .A(n5329), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9964) );
  INV_X1 U6839 ( .A(n9964), .ZN(n6094) );
  INV_X1 U6840 ( .A(n5332), .ZN(n5333) );
  NAND2_X1 U6841 ( .A1(n5333), .A2(SI_5_), .ZN(n5334) );
  MUX2_X1 U6842 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7631), .Z(n5357) );
  XNOR2_X1 U6843 ( .A(n5357), .B(n9498), .ZN(n5355) );
  XNOR2_X1 U6844 ( .A(n5356), .B(n5355), .ZN(n6866) );
  OR2_X1 U6845 ( .A1(n5304), .A2(n6866), .ZN(n5336) );
  INV_X1 U6846 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6009) );
  OR2_X1 U6847 ( .A1(n8745), .A2(n6009), .ZN(n5335) );
  OAI211_X1 U6848 ( .C1(n5307), .C2(n6094), .A(n5336), .B(n5335), .ZN(n10067)
         );
  NAND2_X1 U6849 ( .A1(n10067), .A2(n5903), .ZN(n5337) );
  NAND2_X1 U6850 ( .A1(n5338), .A2(n5337), .ZN(n5339) );
  XNOR2_X1 U6851 ( .A(n5339), .B(n5511), .ZN(n5341) );
  AND2_X1 U6852 ( .A1(n10067), .A2(n5580), .ZN(n5340) );
  AOI21_X1 U6853 ( .B1(n10166), .B2(n5935), .A(n5340), .ZN(n5342) );
  XNOR2_X1 U6854 ( .A(n5341), .B(n5342), .ZN(n6836) );
  NAND2_X1 U6855 ( .A1(n6802), .A2(n6836), .ZN(n6834) );
  INV_X1 U6856 ( .A(n5341), .ZN(n5343) );
  NAND2_X1 U6857 ( .A1(n5343), .A2(n5342), .ZN(n5344) );
  NAND2_X1 U6858 ( .A1(n5241), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U6859 ( .A1(n6067), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5351) );
  INV_X1 U6860 ( .A(n5347), .ZN(n5345) );
  NAND2_X1 U6861 ( .A1(n5345), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5366) );
  INV_X1 U6862 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6863 ( .A1(n5347), .A2(n5346), .ZN(n5348) );
  AND2_X1 U6864 ( .A1(n5366), .A2(n5348), .ZN(n6953) );
  NAND2_X1 U6865 ( .A1(n5238), .A2(n6953), .ZN(n5350) );
  NAND2_X1 U6866 ( .A1(n6072), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5349) );
  NAND4_X1 U6867 ( .A1(n5352), .A2(n5351), .A3(n5350), .A4(n5349), .ZN(n10065)
         );
  OR2_X1 U6868 ( .A1(n5353), .A2(n5599), .ZN(n5354) );
  XNOR2_X1 U6869 ( .A(n5354), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9837) );
  INV_X1 U6870 ( .A(n9837), .ZN(n6025) );
  NAND2_X1 U6871 ( .A1(n5357), .A2(SI_6_), .ZN(n5358) );
  XNOR2_X1 U6872 ( .A(n5376), .B(SI_7_), .ZN(n5374) );
  XNOR2_X1 U6873 ( .A(n5375), .B(n5374), .ZN(n6917) );
  OR2_X1 U6874 ( .A1(n5304), .A2(n6917), .ZN(n5361) );
  OR2_X1 U6875 ( .A1(n8745), .A2(n6024), .ZN(n5360) );
  OAI211_X1 U6876 ( .C1(n5307), .C2(n6025), .A(n5361), .B(n5360), .ZN(n6951)
         );
  AND2_X1 U6877 ( .A1(n6951), .A2(n5829), .ZN(n5362) );
  AOI21_X1 U6878 ( .B1(n10065), .B2(n5935), .A(n5362), .ZN(n6893) );
  AOI22_X1 U6879 ( .A1(n10065), .A2(n5580), .B1(n6951), .B2(n5903), .ZN(n5363)
         );
  XNOR2_X1 U6880 ( .A(n5363), .B(n5532), .ZN(n6894) );
  INV_X1 U6881 ( .A(n6894), .ZN(n5364) );
  INV_X1 U6882 ( .A(n5388), .ZN(n5385) );
  NAND2_X1 U6883 ( .A1(n6067), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5371) );
  NAND2_X1 U6884 ( .A1(n6072), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5370) );
  INV_X1 U6885 ( .A(n5366), .ZN(n5365) );
  NAND2_X1 U6886 ( .A1(n5365), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5393) );
  INV_X1 U6887 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7138) );
  NAND2_X1 U6888 ( .A1(n5366), .A2(n7138), .ZN(n5367) );
  AND2_X1 U6889 ( .A1(n5393), .A2(n5367), .ZN(n10052) );
  NAND2_X1 U6890 ( .A1(n5238), .A2(n10052), .ZN(n5369) );
  NAND2_X1 U6891 ( .A1(n5241), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5368) );
  NAND4_X1 U6892 ( .A1(n5371), .A2(n5370), .A3(n5369), .A4(n5368), .ZN(n10184)
         );
  NAND2_X1 U6893 ( .A1(n5372), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5373) );
  XNOR2_X1 U6894 ( .A(n5373), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9856) );
  INV_X1 U6895 ( .A(n9856), .ZN(n6035) );
  INV_X1 U6896 ( .A(n5376), .ZN(n5377) );
  NAND2_X1 U6897 ( .A1(n5377), .A2(SI_7_), .ZN(n5378) );
  MUX2_X1 U6898 ( .A(n6032), .B(n6033), .S(n7631), .Z(n5380) );
  INV_X1 U6899 ( .A(SI_8_), .ZN(n5379) );
  NAND2_X1 U6900 ( .A1(n5380), .A2(n5379), .ZN(n5399) );
  INV_X1 U6901 ( .A(n5380), .ZN(n5381) );
  NAND2_X1 U6902 ( .A1(n5381), .A2(SI_8_), .ZN(n5382) );
  NAND2_X1 U6903 ( .A1(n5399), .A2(n5382), .ZN(n5400) );
  OR2_X1 U6904 ( .A1(n8745), .A2(n6033), .ZN(n5383) );
  AOI22_X1 U6905 ( .A1(n10184), .A2(n5829), .B1(n10053), .B2(n5903), .ZN(n5384) );
  XNOR2_X1 U6906 ( .A(n5384), .B(n5511), .ZN(n5386) );
  NAND2_X1 U6907 ( .A1(n5388), .A2(n5387), .ZN(n5389) );
  INV_X1 U6908 ( .A(n10184), .ZN(n7022) );
  OAI22_X1 U6909 ( .A1(n7022), .A2(n5905), .B1(n10179), .B2(n5125), .ZN(n7136)
         );
  INV_X1 U6910 ( .A(n5390), .ZN(n5391) );
  NAND2_X1 U6911 ( .A1(n5241), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U6912 ( .A1(n6067), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6913 ( .A1(n5393), .A2(n5392), .ZN(n5394) );
  AND2_X1 U6914 ( .A1(n5447), .A2(n5394), .ZN(n7224) );
  NAND2_X1 U6915 ( .A1(n5238), .A2(n7224), .ZN(n5396) );
  NAND2_X1 U6916 ( .A1(n6072), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5395) );
  NAND4_X1 U6917 ( .A1(n5398), .A2(n5397), .A3(n5396), .A4(n5395), .ZN(n10193)
         );
  INV_X2 U6918 ( .A(n5125), .ZN(n5580) );
  NAND2_X1 U6919 ( .A1(n10193), .A2(n5580), .ZN(n5412) );
  MUX2_X1 U6920 ( .A(n6045), .B(n6039), .S(n7631), .Z(n5403) );
  INV_X1 U6921 ( .A(SI_9_), .ZN(n5402) );
  NAND2_X1 U6922 ( .A1(n5403), .A2(n5402), .ZN(n5416) );
  INV_X1 U6923 ( .A(n5403), .ZN(n5404) );
  NAND2_X1 U6924 ( .A1(n5404), .A2(SI_9_), .ZN(n5405) );
  OR2_X1 U6925 ( .A1(n5406), .A2(n5121), .ZN(n5407) );
  NAND2_X1 U6926 ( .A1(n5417), .A2(n5407), .ZN(n7087) );
  NAND2_X1 U6927 ( .A1(n7087), .A2(n8738), .ZN(n5410) );
  OR2_X1 U6928 ( .A1(n5372), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U6929 ( .A1(n5427), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5408) );
  XNOR2_X1 U6930 ( .A(n5408), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6365) );
  AOI22_X1 U6931 ( .A1(n5649), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5648), .B2(
        n6365), .ZN(n5409) );
  NAND2_X1 U6932 ( .A1(n5410), .A2(n5409), .ZN(n10183) );
  NAND2_X1 U6933 ( .A1(n10183), .A2(n5903), .ZN(n5411) );
  NAND2_X1 U6934 ( .A1(n5412), .A2(n5411), .ZN(n5413) );
  XNOR2_X1 U6935 ( .A(n5413), .B(n5773), .ZN(n5415) );
  AOI22_X1 U6936 ( .A1(n10193), .A2(n5935), .B1(n5580), .B2(n10183), .ZN(n5414) );
  NOR2_X1 U6937 ( .A1(n5415), .A2(n5414), .ZN(n7222) );
  MUX2_X1 U6938 ( .A(n6048), .B(n5418), .S(n7631), .Z(n5420) );
  XNOR2_X1 U6939 ( .A(n5420), .B(SI_10_), .ZN(n5442) );
  INV_X1 U6940 ( .A(n5442), .ZN(n5419) );
  INV_X1 U6941 ( .A(n5420), .ZN(n5421) );
  NAND2_X1 U6942 ( .A1(n5421), .A2(SI_10_), .ZN(n5422) );
  MUX2_X1 U6943 ( .A(n6064), .B(n6065), .S(n7631), .Z(n5424) );
  INV_X1 U6944 ( .A(SI_11_), .ZN(n5423) );
  NAND2_X1 U6945 ( .A1(n5424), .A2(n5423), .ZN(n5472) );
  INV_X1 U6946 ( .A(n5424), .ZN(n5425) );
  NAND2_X1 U6947 ( .A1(n5425), .A2(SI_11_), .ZN(n5426) );
  NAND2_X1 U6948 ( .A1(n5472), .A2(n5426), .ZN(n5471) );
  XNOR2_X1 U6949 ( .A(n5470), .B(n5471), .ZN(n7265) );
  NAND2_X1 U6950 ( .A1(n7265), .A2(n8738), .ZN(n5431) );
  NAND2_X1 U6951 ( .A1(n5476), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U6952 ( .A1(n5444), .A2(n5474), .ZN(n5428) );
  NAND2_X1 U6953 ( .A1(n5428), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5429) );
  XNOR2_X1 U6954 ( .A(n5429), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9978) );
  AOI22_X1 U6955 ( .A1(n5649), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5648), .B2(
        n9978), .ZN(n5430) );
  NAND2_X1 U6956 ( .A1(n10209), .A2(n5903), .ZN(n5440) );
  NAND2_X1 U6957 ( .A1(n5241), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5438) );
  NAND2_X1 U6958 ( .A1(n6067), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U6959 ( .A1(n5432), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5482) );
  INV_X1 U6960 ( .A(n5432), .ZN(n5449) );
  INV_X1 U6961 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U6962 ( .A1(n5449), .A2(n5433), .ZN(n5434) );
  AND2_X1 U6963 ( .A1(n5482), .A2(n5434), .ZN(n8707) );
  NAND2_X1 U6964 ( .A1(n5238), .A2(n8707), .ZN(n5436) );
  NAND2_X1 U6965 ( .A1(n6072), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5435) );
  NAND4_X1 U6966 ( .A1(n5438), .A2(n5437), .A3(n5436), .A4(n5435), .ZN(n10192)
         );
  NAND2_X1 U6967 ( .A1(n10192), .A2(n5580), .ZN(n5439) );
  NAND2_X1 U6968 ( .A1(n5440), .A2(n5439), .ZN(n5441) );
  XNOR2_X1 U6969 ( .A(n5441), .B(n5773), .ZN(n5463) );
  AOI22_X1 U6970 ( .A1(n10209), .A2(n5580), .B1(n5935), .B2(n10192), .ZN(n8703) );
  XNOR2_X1 U6971 ( .A(n5443), .B(n5442), .ZN(n7146) );
  NAND2_X1 U6972 ( .A1(n7146), .A2(n8738), .ZN(n5446) );
  XNOR2_X1 U6973 ( .A(n5444), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9832) );
  AOI22_X1 U6974 ( .A1(n5649), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5648), .B2(
        n9832), .ZN(n5445) );
  NAND2_X1 U6975 ( .A1(n5446), .A2(n5445), .ZN(n7393) );
  NAND2_X1 U6976 ( .A1(n7393), .A2(n5903), .ZN(n5455) );
  NAND2_X1 U6977 ( .A1(n6067), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U6978 ( .A1(n6072), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U6979 ( .A1(n5447), .A2(n7388), .ZN(n5448) );
  AND2_X1 U6980 ( .A1(n5449), .A2(n5448), .ZN(n7387) );
  NAND2_X1 U6981 ( .A1(n5238), .A2(n7387), .ZN(n5451) );
  NAND2_X1 U6982 ( .A1(n5241), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5450) );
  NAND4_X1 U6983 ( .A1(n5453), .A2(n5452), .A3(n5451), .A4(n5450), .ZN(n9012)
         );
  NAND2_X1 U6984 ( .A1(n9012), .A2(n5580), .ZN(n5454) );
  NAND2_X1 U6985 ( .A1(n5455), .A2(n5454), .ZN(n5456) );
  XNOR2_X1 U6986 ( .A(n5456), .B(n5532), .ZN(n5462) );
  NAND2_X1 U6987 ( .A1(n7393), .A2(n5580), .ZN(n5458) );
  NAND2_X1 U6988 ( .A1(n9012), .A2(n5935), .ZN(n5457) );
  NAND2_X1 U6989 ( .A1(n5458), .A2(n5457), .ZN(n7385) );
  NAND2_X1 U6990 ( .A1(n5462), .A2(n7385), .ZN(n5459) );
  OAI21_X1 U6991 ( .B1(n5463), .B2(n8703), .A(n5459), .ZN(n5460) );
  INV_X1 U6992 ( .A(n5460), .ZN(n5461) );
  NAND2_X1 U6993 ( .A1(n8701), .A2(n5461), .ZN(n5469) );
  INV_X1 U6994 ( .A(n7385), .ZN(n5464) );
  AOI21_X1 U6995 ( .B1(n8702), .B2(n5464), .A(n8703), .ZN(n5466) );
  INV_X1 U6996 ( .A(n5463), .ZN(n8704) );
  NAND3_X1 U6997 ( .A1(n8703), .A2(n5464), .A3(n8702), .ZN(n5465) );
  NAND2_X1 U6998 ( .A1(n5469), .A2(n5468), .ZN(n7396) );
  MUX2_X1 U6999 ( .A(n6080), .B(n6121), .S(n7631), .Z(n5495) );
  XNOR2_X1 U7000 ( .A(n5495), .B(SI_12_), .ZN(n5494) );
  XNOR2_X1 U7001 ( .A(n5497), .B(n5494), .ZN(n7269) );
  NAND2_X1 U7002 ( .A1(n7269), .A2(n8738), .ZN(n5479) );
  NAND2_X1 U7003 ( .A1(n5474), .A2(n5473), .ZN(n5475) );
  NOR2_X1 U7004 ( .A1(n5476), .A2(n5475), .ZN(n5499) );
  OR2_X1 U7005 ( .A1(n5499), .A2(n5599), .ZN(n5477) );
  XNOR2_X1 U7006 ( .A(n5477), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7120) );
  AOI22_X1 U7007 ( .A1(n5649), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5648), .B2(
        n7120), .ZN(n5478) );
  NAND2_X1 U7008 ( .A1(n10219), .A2(n5903), .ZN(n5489) );
  NAND2_X1 U7009 ( .A1(n5241), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U7010 ( .A1(n6067), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5486) );
  INV_X1 U7011 ( .A(n5482), .ZN(n5480) );
  NAND2_X1 U7012 ( .A1(n5480), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5503) );
  INV_X1 U7013 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5481) );
  NAND2_X1 U7014 ( .A1(n5482), .A2(n5481), .ZN(n5483) );
  AND2_X1 U7015 ( .A1(n5503), .A2(n5483), .ZN(n7401) );
  NAND2_X1 U7016 ( .A1(n5238), .A2(n7401), .ZN(n5485) );
  NAND2_X1 U7017 ( .A1(n6072), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5484) );
  NAND4_X1 U7018 ( .A1(n5487), .A2(n5486), .A3(n5485), .A4(n5484), .ZN(n9011)
         );
  NAND2_X1 U7019 ( .A1(n9011), .A2(n5580), .ZN(n5488) );
  NAND2_X1 U7020 ( .A1(n5489), .A2(n5488), .ZN(n5490) );
  XNOR2_X1 U7021 ( .A(n5490), .B(n5511), .ZN(n5491) );
  AOI22_X1 U7022 ( .A1(n10219), .A2(n5580), .B1(n5935), .B2(n9011), .ZN(n5492)
         );
  XNOR2_X1 U7023 ( .A(n5491), .B(n5492), .ZN(n7397) );
  INV_X1 U7024 ( .A(n5491), .ZN(n5493) );
  INV_X1 U7025 ( .A(n5495), .ZN(n5496) );
  MUX2_X1 U7026 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7631), .Z(n5518) );
  XNOR2_X1 U7027 ( .A(n5518), .B(SI_13_), .ZN(n5516) );
  XNOR2_X1 U7028 ( .A(n5517), .B(n5516), .ZN(n7319) );
  NAND2_X1 U7029 ( .A1(n7319), .A2(n8738), .ZN(n5502) );
  NAND2_X1 U7030 ( .A1(n5499), .A2(n5498), .ZN(n5521) );
  NAND2_X1 U7031 ( .A1(n5521), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5500) );
  XNOR2_X1 U7032 ( .A(n5500), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10003) );
  AOI22_X1 U7033 ( .A1(n5649), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5648), .B2(
        n10003), .ZN(n5501) );
  NAND2_X1 U7034 ( .A1(n5241), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U7035 ( .A1(n5237), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U7036 ( .A1(n5503), .A2(n8682), .ZN(n5504) );
  AND2_X1 U7037 ( .A1(n5526), .A2(n5504), .ZN(n8686) );
  NAND2_X1 U7038 ( .A1(n5238), .A2(n8686), .ZN(n5506) );
  NAND2_X1 U7039 ( .A1(n6072), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5505) );
  NAND4_X1 U7040 ( .A1(n5508), .A2(n5507), .A3(n5506), .A4(n5505), .ZN(n9010)
         );
  AOI22_X1 U7041 ( .A1(n7190), .A2(n5580), .B1(n5935), .B2(n9010), .ZN(n5513)
         );
  NAND2_X1 U7042 ( .A1(n7190), .A2(n5903), .ZN(n5510) );
  NAND2_X1 U7043 ( .A1(n9010), .A2(n5580), .ZN(n5509) );
  NAND2_X1 U7044 ( .A1(n5510), .A2(n5509), .ZN(n5512) );
  XNOR2_X1 U7045 ( .A(n5512), .B(n5511), .ZN(n5515) );
  XOR2_X1 U7046 ( .A(n5513), .B(n5515), .Z(n8678) );
  INV_X1 U7047 ( .A(n5513), .ZN(n5514) );
  NAND2_X1 U7048 ( .A1(n5518), .A2(SI_13_), .ZN(n5519) );
  NAND2_X1 U7049 ( .A1(n5520), .A2(n5519), .ZN(n5536) );
  XNOR2_X1 U7050 ( .A(n5537), .B(SI_14_), .ZN(n5534) );
  XNOR2_X1 U7051 ( .A(n5536), .B(n5534), .ZN(n7368) );
  NAND2_X1 U7052 ( .A1(n7368), .A2(n8738), .ZN(n5524) );
  NAND2_X1 U7053 ( .A1(n5522), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5564) );
  XNOR2_X1 U7054 ( .A(n5564), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10015) );
  AOI22_X1 U7055 ( .A1(n5649), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5648), .B2(
        n10015), .ZN(n5523) );
  NAND2_X1 U7056 ( .A1(n5241), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U7057 ( .A1(n5237), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5530) );
  INV_X1 U7058 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8600) );
  NAND2_X1 U7059 ( .A1(n5526), .A2(n8600), .ZN(n5527) );
  AND2_X1 U7060 ( .A1(n5571), .A2(n5527), .ZN(n8599) );
  NAND2_X1 U7061 ( .A1(n5238), .A2(n8599), .ZN(n5529) );
  NAND2_X1 U7062 ( .A1(n6072), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5528) );
  NAND4_X1 U7063 ( .A1(n5531), .A2(n5530), .A3(n5529), .A4(n5528), .ZN(n9103)
         );
  AOI22_X1 U7064 ( .A1(n10240), .A2(n5903), .B1(n5829), .B2(n9103), .ZN(n5533)
         );
  XNOR2_X1 U7065 ( .A(n5533), .B(n5532), .ZN(n8596) );
  AOI22_X1 U7066 ( .A1(n10240), .A2(n5580), .B1(n5935), .B2(n9103), .ZN(n8595)
         );
  INV_X1 U7067 ( .A(n5534), .ZN(n5535) );
  NAND2_X1 U7068 ( .A1(n5537), .A2(SI_14_), .ZN(n5538) );
  XNOR2_X1 U7069 ( .A(n5540), .B(SI_15_), .ZN(n5561) );
  NAND2_X1 U7070 ( .A1(n5540), .A2(SI_15_), .ZN(n5541) );
  INV_X1 U7071 ( .A(SI_16_), .ZN(n5542) );
  INV_X1 U7072 ( .A(n5543), .ZN(n5544) );
  NAND2_X1 U7073 ( .A1(n5544), .A2(SI_16_), .ZN(n5545) );
  NAND2_X1 U7074 ( .A1(n5592), .A2(n5545), .ZN(n5593) );
  XNOR2_X1 U7075 ( .A(n5594), .B(n5593), .ZN(n7424) );
  NAND2_X1 U7076 ( .A1(n7424), .A2(n8738), .ZN(n5548) );
  NAND2_X1 U7077 ( .A1(n4597), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5546) );
  XNOR2_X1 U7078 ( .A(n5546), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9064) );
  AOI22_X1 U7079 ( .A1(n5649), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5648), .B2(
        n9064), .ZN(n5547) );
  NAND2_X1 U7080 ( .A1(n9330), .A2(n5903), .ZN(n5558) );
  NAND2_X1 U7081 ( .A1(n5241), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U7082 ( .A1(n6067), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5555) );
  INV_X1 U7083 ( .A(n5571), .ZN(n5549) );
  INV_X1 U7084 ( .A(n5550), .ZN(n5573) );
  INV_X1 U7085 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U7086 ( .A1(n5573), .A2(n5551), .ZN(n5552) );
  AND2_X1 U7087 ( .A1(n5606), .A2(n5552), .ZN(n9323) );
  NAND2_X1 U7088 ( .A1(n5238), .A2(n9323), .ZN(n5554) );
  NAND2_X1 U7089 ( .A1(n6072), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5553) );
  NAND4_X1 U7090 ( .A1(n5556), .A2(n5555), .A3(n5554), .A4(n5553), .ZN(n9343)
         );
  NAND2_X1 U7091 ( .A1(n9343), .A2(n5580), .ZN(n5557) );
  NAND2_X1 U7092 ( .A1(n5558), .A2(n5557), .ZN(n5560) );
  XNOR2_X1 U7093 ( .A(n5560), .B(n5511), .ZN(n8644) );
  AOI22_X1 U7094 ( .A1(n9330), .A2(n5580), .B1(n5935), .B2(n9343), .ZN(n8643)
         );
  INV_X1 U7095 ( .A(n8643), .ZN(n5585) );
  XNOR2_X1 U7096 ( .A(n5562), .B(n5561), .ZN(n7418) );
  NAND2_X1 U7097 ( .A1(n7418), .A2(n8738), .ZN(n5569) );
  NAND2_X1 U7098 ( .A1(n5564), .A2(n5563), .ZN(n5565) );
  NAND2_X1 U7099 ( .A1(n5565), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5567) );
  XNOR2_X1 U7100 ( .A(n5567), .B(n5566), .ZN(n7125) );
  INV_X1 U7101 ( .A(n7125), .ZN(n10028) );
  AOI22_X1 U7102 ( .A1(n5649), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5648), .B2(
        n10028), .ZN(n5568) );
  NAND2_X1 U7103 ( .A1(n9911), .A2(n5580), .ZN(n5579) );
  NAND2_X1 U7104 ( .A1(n6067), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5577) );
  NAND2_X1 U7105 ( .A1(n5241), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5576) );
  INV_X1 U7106 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U7107 ( .A1(n5571), .A2(n5570), .ZN(n5572) );
  AND2_X1 U7108 ( .A1(n5573), .A2(n5572), .ZN(n9345) );
  NAND2_X1 U7109 ( .A1(n5238), .A2(n9345), .ZN(n5575) );
  NAND2_X1 U7110 ( .A1(n6072), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5574) );
  NAND4_X1 U7111 ( .A1(n5577), .A2(n5576), .A3(n5575), .A4(n5574), .ZN(n9897)
         );
  NAND2_X1 U7112 ( .A1(n9897), .A2(n5935), .ZN(n5578) );
  NAND2_X1 U7113 ( .A1(n9911), .A2(n5903), .ZN(n5582) );
  NAND2_X1 U7114 ( .A1(n9897), .A2(n5580), .ZN(n5581) );
  NAND2_X1 U7115 ( .A1(n5582), .A2(n5581), .ZN(n5583) );
  XNOR2_X1 U7116 ( .A(n5583), .B(n5773), .ZN(n8642) );
  INV_X1 U7117 ( .A(n8642), .ZN(n5584) );
  AOI22_X1 U7118 ( .A1(n8644), .A2(n5585), .B1(n8723), .B2(n5584), .ZN(n5591)
         );
  NOR3_X1 U7119 ( .A1(n5585), .A2(n5584), .A3(n8723), .ZN(n5589) );
  AOI21_X1 U7120 ( .B1(n8642), .B2(n5586), .A(n8643), .ZN(n5587) );
  NOR2_X1 U7121 ( .A1(n5587), .A2(n8644), .ZN(n5588) );
  INV_X1 U7122 ( .A(SI_17_), .ZN(n5595) );
  INV_X1 U7123 ( .A(n5596), .ZN(n5597) );
  NAND2_X1 U7124 ( .A1(n5597), .A2(SI_17_), .ZN(n5598) );
  XNOR2_X1 U7125 ( .A(n5618), .B(n5617), .ZN(n7434) );
  NAND2_X1 U7126 ( .A1(n7434), .A2(n8738), .ZN(n5603) );
  OR2_X1 U7127 ( .A1(n5600), .A2(n5599), .ZN(n5601) );
  XNOR2_X1 U7128 ( .A(n5601), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9080) );
  AOI22_X1 U7129 ( .A1(n5649), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5648), .B2(
        n9080), .ZN(n5602) );
  NAND2_X1 U7130 ( .A1(n9892), .A2(n5903), .ZN(n5612) );
  INV_X1 U7131 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9308) );
  INV_X1 U7132 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n5604) );
  OAI22_X1 U7133 ( .A1(n5289), .A2(n9308), .B1(n5877), .B2(n5604), .ZN(n5610)
         );
  INV_X1 U7134 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n5608) );
  INV_X1 U7135 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U7136 ( .A1(n5606), .A2(n5605), .ZN(n5607) );
  NAND2_X1 U7137 ( .A1(n5627), .A2(n5607), .ZN(n9307) );
  OAI22_X1 U7138 ( .A1(n5928), .A2(n5608), .B1(n5943), .B2(n9307), .ZN(n5609)
         );
  NAND2_X1 U7139 ( .A1(n9898), .A2(n5580), .ZN(n5611) );
  NAND2_X1 U7140 ( .A1(n5612), .A2(n5611), .ZN(n5613) );
  XNOR2_X1 U7141 ( .A(n5613), .B(n5511), .ZN(n5614) );
  AOI22_X1 U7142 ( .A1(n9892), .A2(n5580), .B1(n5935), .B2(n9898), .ZN(n5615)
         );
  XNOR2_X1 U7143 ( .A(n5614), .B(n5615), .ZN(n8654) );
  NAND2_X1 U7144 ( .A1(n8655), .A2(n8654), .ZN(n8653) );
  INV_X1 U7145 ( .A(n5614), .ZN(n5616) );
  NAND2_X1 U7146 ( .A1(n8653), .A2(n5116), .ZN(n8715) );
  INV_X1 U7147 ( .A(n8715), .ZN(n5635) );
  INV_X1 U7148 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5620) );
  XNOR2_X1 U7149 ( .A(n5640), .B(SI_18_), .ZN(n5639) );
  XNOR2_X1 U7150 ( .A(n5644), .B(n5639), .ZN(n7443) );
  NAND2_X1 U7151 ( .A1(n7443), .A2(n8738), .ZN(n5624) );
  NAND2_X1 U7152 ( .A1(n5621), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5622) );
  XNOR2_X1 U7153 ( .A(n5622), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10042) );
  AOI22_X1 U7154 ( .A1(n5649), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5648), .B2(
        n10042), .ZN(n5623) );
  NAND2_X1 U7155 ( .A1(n6067), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U7156 ( .A1(n5241), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5631) );
  INV_X1 U7157 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U7158 ( .A1(n5627), .A2(n5626), .ZN(n5628) );
  AND2_X1 U7159 ( .A1(n5654), .A2(n5628), .ZN(n9873) );
  NAND2_X1 U7160 ( .A1(n5238), .A2(n9873), .ZN(n5630) );
  NAND2_X1 U7161 ( .A1(n6072), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5629) );
  NAND4_X1 U7162 ( .A1(n5632), .A2(n5631), .A3(n5630), .A4(n5629), .ZN(n9784)
         );
  AOI22_X1 U7163 ( .A1(n9874), .A2(n5903), .B1(n5829), .B2(n9784), .ZN(n5633)
         );
  XNOR2_X1 U7164 ( .A(n5633), .B(n5511), .ZN(n5637) );
  AOI22_X1 U7165 ( .A1(n9874), .A2(n5580), .B1(n5935), .B2(n9784), .ZN(n5636)
         );
  XNOR2_X1 U7166 ( .A(n5637), .B(n5636), .ZN(n8716) );
  NAND2_X1 U7167 ( .A1(n5637), .A2(n5636), .ZN(n5638) );
  INV_X1 U7168 ( .A(n5639), .ZN(n5643) );
  INV_X1 U7169 ( .A(n5640), .ZN(n5641) );
  NAND2_X1 U7170 ( .A1(n5641), .A2(SI_18_), .ZN(n5642) );
  NAND2_X1 U7171 ( .A1(n5645), .A2(n9668), .ZN(n5667) );
  INV_X1 U7172 ( .A(n5645), .ZN(n5646) );
  NAND2_X1 U7173 ( .A1(n5646), .A2(SI_19_), .ZN(n5647) );
  NAND2_X1 U7174 ( .A1(n5667), .A2(n5647), .ZN(n5668) );
  XNOR2_X1 U7175 ( .A(n5669), .B(n5668), .ZN(n7453) );
  NAND2_X1 U7176 ( .A1(n7453), .A2(n8738), .ZN(n5651) );
  AOI22_X1 U7177 ( .A1(n5649), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8995), .B2(
        n5648), .ZN(n5650) );
  NAND2_X1 U7178 ( .A1(n9298), .A2(n5903), .ZN(n5661) );
  NAND2_X1 U7179 ( .A1(n6067), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5659) );
  NAND2_X1 U7180 ( .A1(n6072), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5658) );
  INV_X1 U7181 ( .A(n5654), .ZN(n5652) );
  NAND2_X1 U7182 ( .A1(n5652), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5676) );
  INV_X1 U7183 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U7184 ( .A1(n5654), .A2(n5653), .ZN(n5655) );
  AND2_X1 U7185 ( .A1(n5676), .A2(n5655), .ZN(n9294) );
  NAND2_X1 U7186 ( .A1(n5238), .A2(n9294), .ZN(n5657) );
  NAND2_X1 U7187 ( .A1(n5241), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5656) );
  NAND4_X1 U7188 ( .A1(n5659), .A2(n5658), .A3(n5657), .A4(n5656), .ZN(n9871)
         );
  NAND2_X1 U7189 ( .A1(n9871), .A2(n5580), .ZN(n5660) );
  NAND2_X1 U7190 ( .A1(n5661), .A2(n5660), .ZN(n5662) );
  XNOR2_X1 U7191 ( .A(n5662), .B(n5511), .ZN(n8618) );
  NAND2_X1 U7192 ( .A1(n9298), .A2(n5580), .ZN(n5664) );
  NAND2_X1 U7193 ( .A1(n9871), .A2(n5935), .ZN(n5663) );
  NAND2_X1 U7194 ( .A1(n5664), .A2(n5663), .ZN(n8617) );
  NOR2_X1 U7195 ( .A1(n8618), .A2(n8617), .ZN(n5666) );
  NAND2_X1 U7196 ( .A1(n8618), .A2(n8617), .ZN(n5665) );
  INV_X1 U7197 ( .A(SI_20_), .ZN(n5670) );
  NAND2_X1 U7198 ( .A1(n5671), .A2(n5670), .ZN(n5690) );
  INV_X1 U7199 ( .A(n5671), .ZN(n5672) );
  NAND2_X1 U7200 ( .A1(n5672), .A2(SI_20_), .ZN(n5673) );
  XNOR2_X1 U7201 ( .A(n5689), .B(n5688), .ZN(n7465) );
  NAND2_X1 U7202 ( .A1(n7465), .A2(n8738), .ZN(n5675) );
  OR2_X1 U7203 ( .A1(n8745), .A2(n6902), .ZN(n5674) );
  NAND2_X1 U7204 ( .A1(n9285), .A2(n5903), .ZN(n5683) );
  NAND2_X1 U7205 ( .A1(n6067), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5681) );
  NAND2_X1 U7206 ( .A1(n5241), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5680) );
  INV_X1 U7207 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9461) );
  NAND2_X1 U7208 ( .A1(n5676), .A2(n9461), .ZN(n5677) );
  AND2_X1 U7209 ( .A1(n5694), .A2(n5677), .ZN(n9280) );
  NAND2_X1 U7210 ( .A1(n5238), .A2(n9280), .ZN(n5679) );
  NAND2_X1 U7211 ( .A1(n6072), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5678) );
  NAND4_X1 U7212 ( .A1(n5681), .A2(n5680), .A3(n5679), .A4(n5678), .ZN(n9783)
         );
  NAND2_X1 U7213 ( .A1(n9783), .A2(n5580), .ZN(n5682) );
  NAND2_X1 U7214 ( .A1(n5683), .A2(n5682), .ZN(n5684) );
  XNOR2_X1 U7215 ( .A(n5684), .B(n5773), .ZN(n5686) );
  AOI22_X1 U7216 ( .A1(n9285), .A2(n5829), .B1(n5935), .B2(n9783), .ZN(n5685)
         );
  NAND2_X1 U7217 ( .A1(n5686), .A2(n5685), .ZN(n5687) );
  OAI21_X1 U7218 ( .B1(n5686), .B2(n5685), .A(n5687), .ZN(n8672) );
  XNOR2_X1 U7219 ( .A(n5708), .B(SI_21_), .ZN(n5707) );
  XNOR2_X1 U7220 ( .A(n5710), .B(n5707), .ZN(n7476) );
  NAND2_X1 U7221 ( .A1(n7476), .A2(n8738), .ZN(n5692) );
  OR2_X1 U7222 ( .A1(n8745), .A2(n6961), .ZN(n5691) );
  NAND2_X1 U7223 ( .A1(n9272), .A2(n5903), .ZN(n5701) );
  NAND2_X1 U7224 ( .A1(n5241), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5699) );
  NAND2_X1 U7225 ( .A1(n6067), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5698) );
  INV_X1 U7226 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5693) );
  NAND2_X1 U7227 ( .A1(n5694), .A2(n5693), .ZN(n5695) );
  AND2_X1 U7228 ( .A1(n5719), .A2(n5695), .ZN(n9267) );
  NAND2_X1 U7229 ( .A1(n5238), .A2(n9267), .ZN(n5697) );
  NAND2_X1 U7230 ( .A1(n6072), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5696) );
  NAND4_X1 U7231 ( .A1(n5699), .A2(n5698), .A3(n5697), .A4(n5696), .ZN(n9775)
         );
  NAND2_X1 U7232 ( .A1(n9775), .A2(n5580), .ZN(n5700) );
  NAND2_X1 U7233 ( .A1(n5701), .A2(n5700), .ZN(n5702) );
  XNOR2_X1 U7234 ( .A(n5702), .B(n5532), .ZN(n5703) );
  AOI22_X1 U7235 ( .A1(n9272), .A2(n5829), .B1(n5935), .B2(n9775), .ZN(n5704)
         );
  XNOR2_X1 U7236 ( .A(n5703), .B(n5704), .ZN(n8628) );
  INV_X1 U7237 ( .A(n5703), .ZN(n5705) );
  NAND2_X1 U7238 ( .A1(n5705), .A2(n5704), .ZN(n5706) );
  INV_X1 U7239 ( .A(n5708), .ZN(n5709) );
  INV_X1 U7240 ( .A(SI_22_), .ZN(n5711) );
  NAND2_X1 U7241 ( .A1(n5712), .A2(n5711), .ZN(n5728) );
  INV_X1 U7242 ( .A(n5712), .ZN(n5713) );
  NAND2_X1 U7243 ( .A1(n5713), .A2(SI_22_), .ZN(n5714) );
  NAND2_X1 U7244 ( .A1(n5728), .A2(n5714), .ZN(n5729) );
  XNOR2_X1 U7245 ( .A(n5730), .B(n5729), .ZN(n7488) );
  NAND2_X1 U7246 ( .A1(n7488), .A2(n8738), .ZN(n5716) );
  OR2_X1 U7247 ( .A1(n8745), .A2(n9604), .ZN(n5715) );
  AOI22_X1 U7248 ( .A1(n6067), .A2(P1_REG1_REG_22__SCAN_IN), .B1(n6072), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n5723) );
  INV_X1 U7249 ( .A(n5719), .ZN(n5717) );
  NAND2_X1 U7250 ( .A1(n5717), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5738) );
  INV_X1 U7251 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5718) );
  NAND2_X1 U7252 ( .A1(n5719), .A2(n5718), .ZN(n5720) );
  NAND2_X1 U7253 ( .A1(n5738), .A2(n5720), .ZN(n9248) );
  OR2_X1 U7254 ( .A1(n9248), .A2(n5943), .ZN(n5722) );
  NAND2_X1 U7255 ( .A1(n5241), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5721) );
  NAND3_X1 U7256 ( .A1(n5723), .A2(n5722), .A3(n5721), .ZN(n9767) );
  AOI22_X1 U7257 ( .A1(n9763), .A2(n5903), .B1(n5580), .B2(n9767), .ZN(n5724)
         );
  XNOR2_X1 U7258 ( .A(n5724), .B(n5511), .ZN(n5725) );
  OAI22_X1 U7259 ( .A1(n4796), .A2(n5125), .B1(n9241), .B2(n5905), .ZN(n8692)
         );
  NAND2_X1 U7260 ( .A1(n8606), .A2(n8607), .ZN(n5751) );
  NAND2_X1 U7261 ( .A1(n5731), .A2(n9615), .ZN(n5754) );
  INV_X1 U7262 ( .A(n5731), .ZN(n5732) );
  NAND2_X1 U7263 ( .A1(n5732), .A2(SI_23_), .ZN(n5733) );
  XNOR2_X1 U7264 ( .A(n5753), .B(n5752), .ZN(n7499) );
  NAND2_X1 U7265 ( .A1(n7499), .A2(n8738), .ZN(n5735) );
  OR2_X1 U7266 ( .A1(n8745), .A2(n7070), .ZN(n5734) );
  NAND2_X1 U7267 ( .A1(n9243), .A2(n5903), .ZN(n5743) );
  INV_X1 U7268 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9238) );
  INV_X1 U7269 ( .A(n5738), .ZN(n5736) );
  NAND2_X1 U7270 ( .A1(n5736), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5763) );
  INV_X1 U7271 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5737) );
  NAND2_X1 U7272 ( .A1(n5738), .A2(n5737), .ZN(n5739) );
  NAND2_X1 U7273 ( .A1(n5763), .A2(n5739), .ZN(n9237) );
  OR2_X1 U7274 ( .A1(n9237), .A2(n5943), .ZN(n5741) );
  AOI22_X1 U7275 ( .A1(n6067), .A2(P1_REG1_REG_23__SCAN_IN), .B1(n5241), .B2(
        P1_REG0_REG_23__SCAN_IN), .ZN(n5740) );
  OAI211_X1 U7276 ( .C1(n5289), .C2(n9238), .A(n5741), .B(n5740), .ZN(n9251)
         );
  NAND2_X1 U7277 ( .A1(n9251), .A2(n5580), .ZN(n5742) );
  NAND2_X1 U7278 ( .A1(n5743), .A2(n5742), .ZN(n5744) );
  XNOR2_X1 U7279 ( .A(n5744), .B(n5773), .ZN(n5746) );
  AND2_X1 U7280 ( .A1(n9251), .A2(n5935), .ZN(n5745) );
  AOI21_X1 U7281 ( .B1(n9243), .B2(n5829), .A(n5745), .ZN(n5747) );
  NAND2_X1 U7282 ( .A1(n5746), .A2(n5747), .ZN(n8660) );
  INV_X1 U7283 ( .A(n5746), .ZN(n5749) );
  INV_X1 U7284 ( .A(n5747), .ZN(n5748) );
  NAND2_X1 U7285 ( .A1(n5749), .A2(n5748), .ZN(n5750) );
  NAND2_X1 U7286 ( .A1(n5751), .A2(n8608), .ZN(n8610) );
  NAND2_X1 U7287 ( .A1(n8610), .A2(n8660), .ZN(n5781) );
  NAND2_X1 U7288 ( .A1(n5753), .A2(n5752), .ZN(n5755) );
  INV_X1 U7289 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7508) );
  INV_X1 U7290 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7219) );
  INV_X1 U7291 ( .A(SI_24_), .ZN(n5756) );
  NAND2_X1 U7292 ( .A1(n5757), .A2(n5756), .ZN(n5785) );
  INV_X1 U7293 ( .A(n5757), .ZN(n5758) );
  NAND2_X1 U7294 ( .A1(n5758), .A2(SI_24_), .ZN(n5759) );
  XNOR2_X1 U7295 ( .A(n5784), .B(n5783), .ZN(n7507) );
  NAND2_X1 U7296 ( .A1(n7507), .A2(n8738), .ZN(n5761) );
  OR2_X1 U7297 ( .A1(n8745), .A2(n7219), .ZN(n5760) );
  NAND2_X1 U7298 ( .A1(n9750), .A2(n5903), .ZN(n5772) );
  INV_X1 U7299 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U7300 ( .A1(n5763), .A2(n5762), .ZN(n5764) );
  AND2_X1 U7301 ( .A1(n5818), .A2(n5764), .ZN(n9219) );
  NAND2_X1 U7302 ( .A1(n9219), .A2(n5238), .ZN(n5770) );
  INV_X1 U7303 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5767) );
  NAND2_X1 U7304 ( .A1(n5241), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5766) );
  NAND2_X1 U7305 ( .A1(n6072), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5765) );
  OAI211_X1 U7306 ( .C1(n5928), .C2(n5767), .A(n5766), .B(n5765), .ZN(n5768)
         );
  INV_X1 U7307 ( .A(n5768), .ZN(n5769) );
  NAND2_X1 U7308 ( .A1(n9754), .A2(n5580), .ZN(n5771) );
  NAND2_X1 U7309 ( .A1(n5772), .A2(n5771), .ZN(n5774) );
  XNOR2_X1 U7310 ( .A(n5774), .B(n5773), .ZN(n5776) );
  AND2_X1 U7311 ( .A1(n9754), .A2(n5935), .ZN(n5775) );
  AOI21_X1 U7312 ( .B1(n9750), .B2(n5829), .A(n5775), .ZN(n5777) );
  NAND2_X1 U7313 ( .A1(n5776), .A2(n5777), .ZN(n5782) );
  INV_X1 U7314 ( .A(n5776), .ZN(n5779) );
  INV_X1 U7315 ( .A(n5777), .ZN(n5778) );
  NAND2_X1 U7316 ( .A1(n5779), .A2(n5778), .ZN(n5780) );
  NAND2_X1 U7317 ( .A1(n8664), .A2(n5782), .ZN(n8634) );
  INV_X1 U7318 ( .A(SI_25_), .ZN(n5786) );
  NAND2_X1 U7319 ( .A1(n5787), .A2(n5786), .ZN(n5806) );
  INV_X1 U7320 ( .A(n5787), .ZN(n5788) );
  NAND2_X1 U7321 ( .A1(n5788), .A2(SI_25_), .ZN(n5789) );
  XNOR2_X1 U7322 ( .A(n5805), .B(n5804), .ZN(n7516) );
  NAND2_X1 U7323 ( .A1(n7516), .A2(n8738), .ZN(n5791) );
  NAND2_X1 U7324 ( .A1(n9202), .A2(n5903), .ZN(n5799) );
  XNOR2_X1 U7325 ( .A(n5818), .B(P1_REG3_REG_25__SCAN_IN), .ZN(n9203) );
  NAND2_X1 U7326 ( .A1(n9203), .A2(n5238), .ZN(n5797) );
  INV_X1 U7327 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7328 ( .A1(n5241), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U7329 ( .A1(n6072), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5792) );
  OAI211_X1 U7330 ( .C1(n5928), .C2(n5794), .A(n5793), .B(n5792), .ZN(n5795)
         );
  INV_X1 U7331 ( .A(n5795), .ZN(n5796) );
  NAND2_X1 U7332 ( .A1(n9222), .A2(n5580), .ZN(n5798) );
  NAND2_X1 U7333 ( .A1(n5799), .A2(n5798), .ZN(n5800) );
  XNOR2_X1 U7334 ( .A(n5800), .B(n5511), .ZN(n5801) );
  AOI22_X1 U7335 ( .A1(n9202), .A2(n5829), .B1(n5935), .B2(n9222), .ZN(n5802)
         );
  XNOR2_X1 U7336 ( .A(n5801), .B(n5802), .ZN(n8635) );
  INV_X1 U7337 ( .A(n5801), .ZN(n5803) );
  NAND2_X1 U7338 ( .A1(n5803), .A2(n5802), .ZN(n5830) );
  AND2_X1 U7339 ( .A1(n5832), .A2(n5830), .ZN(n5859) );
  INV_X1 U7340 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8579) );
  INV_X1 U7341 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9818) );
  INV_X1 U7342 ( .A(SI_26_), .ZN(n5808) );
  NAND2_X1 U7343 ( .A1(n5809), .A2(n5808), .ZN(n5892) );
  INV_X1 U7344 ( .A(n5809), .ZN(n5810) );
  NAND2_X1 U7345 ( .A1(n5810), .A2(SI_26_), .ZN(n5811) );
  NAND2_X1 U7346 ( .A1(n8577), .A2(n8738), .ZN(n5813) );
  OR2_X1 U7347 ( .A1(n8745), .A2(n9818), .ZN(n5812) );
  NAND2_X1 U7348 ( .A1(n9736), .A2(n5903), .ZN(n5826) );
  INV_X1 U7349 ( .A(n5818), .ZN(n5815) );
  AND2_X1 U7350 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n5814) );
  NAND2_X1 U7351 ( .A1(n5815), .A2(n5814), .ZN(n5873) );
  INV_X1 U7352 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5817) );
  INV_X1 U7353 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5816) );
  OAI21_X1 U7354 ( .B1(n5818), .B2(n5817), .A(n5816), .ZN(n5819) );
  NAND2_X1 U7355 ( .A1(n5873), .A2(n5819), .ZN(n5862) );
  INV_X1 U7356 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9630) );
  NAND2_X1 U7357 ( .A1(n6072), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5821) );
  NAND2_X1 U7358 ( .A1(n5241), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5820) );
  OAI211_X1 U7359 ( .C1(n5928), .C2(n9630), .A(n5821), .B(n5820), .ZN(n5822)
         );
  INV_X1 U7360 ( .A(n5822), .ZN(n5823) );
  NAND2_X1 U7361 ( .A1(n9741), .A2(n5580), .ZN(n5825) );
  NAND2_X1 U7362 ( .A1(n5826), .A2(n5825), .ZN(n5827) );
  XNOR2_X1 U7363 ( .A(n5827), .B(n5532), .ZN(n5910) );
  AND2_X1 U7364 ( .A1(n9741), .A2(n5935), .ZN(n5828) );
  AOI21_X1 U7365 ( .B1(n9736), .B2(n5580), .A(n5828), .ZN(n5908) );
  XNOR2_X1 U7366 ( .A(n5910), .B(n5908), .ZN(n5858) );
  NAND2_X1 U7367 ( .A1(n5832), .A2(n5831), .ZN(n8586) );
  INV_X1 U7368 ( .A(n6167), .ZN(n8939) );
  AND2_X1 U7369 ( .A1(n7068), .A2(n8939), .ZN(n7409) );
  NAND2_X1 U7370 ( .A1(n10227), .A2(n8931), .ZN(n5864) );
  NOR2_X1 U7371 ( .A1(n5864), .A2(n6037), .ZN(n5856) );
  NAND2_X1 U7372 ( .A1(n7246), .A2(P1_B_REG_SCAN_IN), .ZN(n5838) );
  MUX2_X1 U7373 ( .A(n5838), .B(P1_B_REG_SCAN_IN), .S(n5852), .Z(n5839) );
  INV_X1 U7374 ( .A(n5840), .ZN(n9821) );
  NAND2_X1 U7375 ( .A1(n9821), .A2(n7246), .ZN(n9805) );
  OAI21_X1 U7376 ( .B1(n6057), .B2(P1_D_REG_1__SCAN_IN), .A(n9805), .ZN(n6160)
         );
  NOR2_X1 U7377 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .ZN(
        n5844) );
  NOR4_X1 U7378 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5843) );
  NOR4_X1 U7379 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5842) );
  NOR4_X1 U7380 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5841) );
  NAND4_X1 U7381 ( .A1(n5844), .A2(n5843), .A3(n5842), .A4(n5841), .ZN(n5850)
         );
  NOR4_X1 U7382 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5848) );
  NOR4_X1 U7383 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5847) );
  NOR4_X1 U7384 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5846) );
  NOR4_X1 U7385 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5845) );
  NAND4_X1 U7386 ( .A1(n5848), .A2(n5847), .A3(n5846), .A4(n5845), .ZN(n5849)
         );
  NOR2_X1 U7387 ( .A1(n5850), .A2(n5849), .ZN(n6155) );
  NOR2_X1 U7388 ( .A1(n6057), .A2(n6155), .ZN(n5851) );
  NOR2_X1 U7389 ( .A1(n6160), .A2(n5851), .ZN(n5855) );
  INV_X1 U7390 ( .A(n6057), .ZN(n5854) );
  INV_X1 U7391 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5853) );
  INV_X1 U7392 ( .A(n5852), .ZN(n7221) );
  AND2_X1 U7393 ( .A1(n5855), .A2(n6172), .ZN(n5871) );
  NOR2_X1 U7394 ( .A1(n6169), .A2(n6904), .ZN(n5863) );
  NAND2_X1 U7395 ( .A1(n6156), .A2(n5863), .ZN(n5860) );
  INV_X1 U7396 ( .A(n5871), .ZN(n5868) );
  OR2_X1 U7397 ( .A1(n5860), .A2(n5868), .ZN(n5861) );
  INV_X1 U7398 ( .A(n5862), .ZN(n9190) );
  INV_X1 U7399 ( .A(n5863), .ZN(n6727) );
  NAND2_X1 U7400 ( .A1(n5864), .A2(n6727), .ZN(n5865) );
  NAND2_X1 U7401 ( .A1(n5868), .A2(n5865), .ZN(n5866) );
  NAND2_X1 U7402 ( .A1(n5882), .A2(n6163), .ZN(n6157) );
  NAND3_X1 U7403 ( .A1(n5866), .A2(n5996), .A3(n6157), .ZN(n5867) );
  NAND2_X1 U7404 ( .A1(n5867), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5870) );
  NOR2_X1 U7405 ( .A1(n8931), .A2(n6163), .ZN(n7408) );
  NAND3_X1 U7406 ( .A1(n5868), .A2(n6156), .A3(n7408), .ZN(n5869) );
  AND2_X1 U7407 ( .A1(n5870), .A2(n5869), .ZN(n6183) );
  NAND2_X1 U7408 ( .A1(n6181), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9007) );
  INV_X1 U7409 ( .A(n9222), .ZN(n8837) );
  NOR2_X1 U7410 ( .A1(n6037), .A2(n6163), .ZN(n9003) );
  AND2_X1 U7411 ( .A1(n9003), .A2(n5871), .ZN(n5881) );
  INV_X1 U7412 ( .A(n5872), .ZN(n9027) );
  AND2_X2 U7413 ( .A1(n5882), .A2(n9027), .ZN(n10194) );
  NAND2_X1 U7414 ( .A1(n5881), .A2(n10194), .ZN(n8683) );
  INV_X1 U7415 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9616) );
  NAND2_X1 U7416 ( .A1(n5873), .A2(n9616), .ZN(n5874) );
  NAND2_X1 U7417 ( .A1(n9174), .A2(n5238), .ZN(n5880) );
  INV_X1 U7418 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9631) );
  NAND2_X1 U7419 ( .A1(n6067), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5876) );
  NAND2_X1 U7420 ( .A1(n6072), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5875) );
  OAI211_X1 U7421 ( .C1(n5877), .C2(n9631), .A(n5876), .B(n5875), .ZN(n5878)
         );
  INV_X1 U7422 ( .A(n5878), .ZN(n5879) );
  INV_X1 U7423 ( .A(n5881), .ZN(n5883) );
  NAND2_X1 U7424 ( .A1(n5882), .A2(n5872), .ZN(n10236) );
  NOR2_X2 U7425 ( .A1(n5883), .A2(n10236), .ZN(n8693) );
  AOI22_X1 U7426 ( .A1(n9735), .A2(n8693), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n5884) );
  OAI21_X1 U7427 ( .B1(n8837), .B2(n8683), .A(n5884), .ZN(n5885) );
  AOI21_X1 U7428 ( .B1(n9190), .B2(n8725), .A(n5885), .ZN(n5886) );
  OAI21_X1 U7429 ( .B1(n9195), .B2(n8689), .A(n5886), .ZN(n5887) );
  INV_X1 U7430 ( .A(n5887), .ZN(n5888) );
  NAND2_X1 U7431 ( .A1(n5891), .A2(n5890), .ZN(n5893) );
  INV_X1 U7432 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7542) );
  INV_X1 U7433 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9815) );
  INV_X1 U7434 ( .A(SI_27_), .ZN(n5894) );
  NAND2_X1 U7435 ( .A1(n5895), .A2(n5894), .ZN(n5914) );
  INV_X1 U7436 ( .A(n5895), .ZN(n5896) );
  NAND2_X1 U7437 ( .A1(n5896), .A2(SI_27_), .ZN(n5897) );
  OR2_X1 U7438 ( .A1(n5899), .A2(n5898), .ZN(n5900) );
  NAND2_X1 U7439 ( .A1(n5915), .A2(n5900), .ZN(n8572) );
  NAND2_X1 U7440 ( .A1(n8572), .A2(n8738), .ZN(n5902) );
  AOI22_X1 U7441 ( .A1(n9730), .A2(n5903), .B1(n5829), .B2(n9735), .ZN(n5904)
         );
  XOR2_X1 U7442 ( .A(n5511), .B(n5904), .Z(n5907) );
  INV_X1 U7443 ( .A(n9730), .ZN(n9176) );
  OAI22_X1 U7444 ( .A1(n9176), .A2(n5125), .B1(n9193), .B2(n5905), .ZN(n5906)
         );
  NOR2_X1 U7445 ( .A1(n5907), .A2(n5906), .ZN(n5941) );
  AOI21_X1 U7446 ( .B1(n5907), .B2(n5906), .A(n5941), .ZN(n8584) );
  INV_X1 U7447 ( .A(n8584), .ZN(n5912) );
  INV_X1 U7448 ( .A(n5908), .ZN(n5909) );
  NAND2_X1 U7449 ( .A1(n5910), .A2(n5909), .ZN(n8585) );
  INV_X1 U7450 ( .A(n8585), .ZN(n5911) );
  NOR2_X1 U7451 ( .A1(n5912), .A2(n5911), .ZN(n5913) );
  AND2_X2 U7452 ( .A1(n8586), .A2(n5913), .ZN(n8588) );
  INV_X1 U7453 ( .A(n8588), .ZN(n5940) );
  INV_X1 U7454 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9496) );
  INV_X1 U7455 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7405) );
  MUX2_X1 U7456 ( .A(n9496), .B(n7405), .S(n7631), .Z(n5917) );
  INV_X1 U7457 ( .A(SI_28_), .ZN(n5916) );
  NAND2_X1 U7458 ( .A1(n5917), .A2(n5916), .ZN(n7630) );
  INV_X1 U7459 ( .A(n5917), .ZN(n5918) );
  NAND2_X1 U7460 ( .A1(n5918), .A2(SI_28_), .ZN(n5919) );
  NAND2_X1 U7461 ( .A1(n8569), .A2(n8738), .ZN(n5921) );
  OR2_X1 U7462 ( .A1(n8745), .A2(n7405), .ZN(n5920) );
  NAND2_X1 U7463 ( .A1(n9160), .A2(n5903), .ZN(n5933) );
  INV_X1 U7464 ( .A(n5924), .ZN(n5922) );
  NAND2_X1 U7465 ( .A1(n5922), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9132) );
  INV_X1 U7466 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U7467 ( .A1(n5924), .A2(n5923), .ZN(n5925) );
  NAND2_X1 U7468 ( .A1(n9132), .A2(n5925), .ZN(n9161) );
  INV_X1 U7469 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9624) );
  NAND2_X1 U7470 ( .A1(n5241), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U7471 ( .A1(n6072), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5926) );
  OAI211_X1 U7472 ( .C1(n5928), .C2(n9624), .A(n5927), .B(n5926), .ZN(n5929)
         );
  INV_X1 U7473 ( .A(n5929), .ZN(n5930) );
  NAND2_X1 U7474 ( .A1(n9180), .A2(n5580), .ZN(n5932) );
  NAND2_X1 U7475 ( .A1(n5933), .A2(n5932), .ZN(n5934) );
  XNOR2_X1 U7476 ( .A(n5934), .B(n5511), .ZN(n5937) );
  AOI22_X1 U7477 ( .A1(n9160), .A2(n5580), .B1(n5935), .B2(n9180), .ZN(n5936)
         );
  XNOR2_X1 U7478 ( .A(n5937), .B(n5936), .ZN(n5942) );
  INV_X1 U7479 ( .A(n5942), .ZN(n5939) );
  INV_X1 U7480 ( .A(n5941), .ZN(n5938) );
  NAND3_X1 U7481 ( .A1(n8588), .A2(n8680), .A3(n5942), .ZN(n5955) );
  AOI22_X1 U7482 ( .A1(n9735), .A2(n8726), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n5950) );
  OR2_X1 U7483 ( .A1(n9132), .A2(n5943), .ZN(n5948) );
  NAND2_X1 U7484 ( .A1(n6072), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7485 ( .A1(n6067), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7486 ( .A1(n5241), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5944) );
  AND3_X1 U7487 ( .A1(n5946), .A2(n5945), .A3(n5944), .ZN(n5947) );
  NAND2_X1 U7488 ( .A1(n5948), .A2(n5947), .ZN(n9009) );
  NAND2_X1 U7489 ( .A1(n9009), .A2(n8693), .ZN(n5949) );
  OAI211_X1 U7490 ( .C1(n8696), .C2(n9161), .A(n5950), .B(n5949), .ZN(n5951)
         );
  AOI21_X1 U7491 ( .B1(n9160), .B2(n8731), .A(n5951), .ZN(n5952) );
  NAND3_X1 U7492 ( .A1(n5956), .A2(n5955), .A3(n5954), .ZN(P1_U3220) );
  INV_X1 U7493 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7494 ( .A1(n6411), .A2(n5962), .ZN(n6524) );
  INV_X1 U7495 ( .A(n6524), .ZN(n5963) );
  NAND2_X1 U7496 ( .A1(n6280), .A2(n6281), .ZN(n5964) );
  NOR2_X1 U7497 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5968) );
  NAND2_X1 U7498 ( .A1(n4586), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5973) );
  INV_X1 U7499 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7500 ( .A1(n5987), .A2(n5988), .ZN(n5974) );
  NAND2_X1 U7501 ( .A1(n5976), .A2(n5979), .ZN(n5977) );
  INV_X1 U7502 ( .A(n6027), .ZN(n5986) );
  NAND2_X1 U7503 ( .A1(n5978), .A2(n5977), .ZN(n6026) );
  NAND2_X1 U7504 ( .A1(n5983), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5981) );
  MUX2_X1 U7505 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5981), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5982) );
  INV_X1 U7506 ( .A(n6055), .ZN(n8580) );
  NOR2_X1 U7507 ( .A1(n6026), .A2(n8580), .ZN(n5985) );
  NAND2_X1 U7508 ( .A1(n7850), .A2(n6287), .ZN(n5989) );
  XNOR2_X1 U7509 ( .A(n5987), .B(n5988), .ZN(n6286) );
  NAND2_X1 U7510 ( .A1(n5989), .A2(n6286), .ZN(n6141) );
  NAND2_X1 U7511 ( .A1(n6297), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7512 ( .A1(n6141), .A2(n6476), .ZN(n5995) );
  NAND2_X1 U7513 ( .A1(n5995), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U7514 ( .A(n6286), .ZN(n7071) );
  OR3_X2 U7515 ( .A1(n6181), .A2(P1_U3086), .A3(n5996), .ZN(n9030) );
  INV_X1 U7516 ( .A(n9030), .ZN(P1_U3973) );
  AND2_X1 U7517 ( .A1(n7631), .A2(P2_U3151), .ZN(n8574) );
  INV_X2 U7518 ( .A(n8574), .ZN(n8578) );
  INV_X1 U7519 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7520 ( .A1(n5201), .A2(P2_U3151), .ZN(n8576) );
  OAI222_X1 U7521 ( .A1(n8578), .A2(n5998), .B1(n8576), .B2(n6003), .C1(
        P2_U3151), .C2(n6213), .ZN(P2_U3294) );
  INV_X1 U7522 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U7523 ( .A1(n6021), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5999) );
  MUX2_X1 U7524 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5999), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n6002) );
  INV_X1 U7525 ( .A(n6021), .ZN(n6001) );
  INV_X1 U7526 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7527 ( .A1(n6001), .A2(n6000), .ZN(n6015) );
  NAND2_X1 U7528 ( .A1(n6002), .A2(n6015), .ZN(n6640) );
  OAI222_X1 U7529 ( .A1(n8578), .A2(n4726), .B1(n8576), .B2(n6639), .C1(
        P2_U3151), .C2(n6640), .ZN(P2_U3291) );
  NAND2_X1 U7530 ( .A1(n5201), .A2(P1_U3086), .ZN(n9817) );
  NOR2_X1 U7531 ( .A1(n5201), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9806) );
  INV_X2 U7532 ( .A(n9806), .ZN(n9820) );
  OAI222_X1 U7533 ( .A1(n9817), .A2(n6004), .B1(n9820), .B2(n6003), .C1(n6101), 
        .C2(P1_U3086), .ZN(P1_U3354) );
  OAI222_X1 U7534 ( .A1(n9817), .A2(n6005), .B1(n9820), .B2(n6493), .C1(n6104), 
        .C2(P1_U3086), .ZN(P1_U3352) );
  OAI222_X1 U7535 ( .A1(n9817), .A2(n6006), .B1(n9820), .B2(n6481), .C1(n6100), 
        .C2(P1_U3086), .ZN(P1_U3353) );
  OAI222_X1 U7536 ( .A1(n6106), .A2(P1_U3086), .B1(n9820), .B2(n6639), .C1(
        n6007), .C2(n9817), .ZN(P1_U3351) );
  OAI222_X1 U7537 ( .A1(n6092), .A2(P1_U3086), .B1(n9820), .B2(n6774), .C1(
        n6008), .C2(n9817), .ZN(P1_U3350) );
  OAI222_X1 U7538 ( .A1(n6094), .A2(P1_U3086), .B1(n9820), .B2(n6866), .C1(
        n6009), .C2(n9817), .ZN(P1_U3349) );
  INV_X1 U7539 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6867) );
  NAND2_X1 U7540 ( .A1(n6017), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6011) );
  MUX2_X1 U7541 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6011), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n6012) );
  AND2_X1 U7542 ( .A1(n6012), .A2(n4583), .ZN(n6348) );
  OAI222_X1 U7543 ( .A1(n8578), .A2(n6867), .B1(n8576), .B2(n6866), .C1(
        P2_U3151), .C2(n6868), .ZN(P2_U3289) );
  INV_X1 U7544 ( .A(n8576), .ZN(n8568) );
  INV_X1 U7545 ( .A(n8568), .ZN(n8582) );
  OAI222_X1 U7546 ( .A1(n8578), .A2(n6480), .B1(n8582), .B2(n6481), .C1(
        P2_U3151), .C2(n6482), .ZN(P2_U3293) );
  NAND2_X1 U7547 ( .A1(n6015), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6016) );
  MUX2_X1 U7548 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6016), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n6018) );
  NAND2_X1 U7549 ( .A1(n6018), .A2(n6017), .ZN(n6778) );
  OAI222_X1 U7550 ( .A1(n8578), .A2(n6775), .B1(n8582), .B2(n6774), .C1(
        P2_U3151), .C2(n6778), .ZN(P2_U3290) );
  NAND2_X1 U7551 ( .A1(n6019), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6020) );
  MUX2_X1 U7552 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6020), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n6022) );
  NAND2_X1 U7553 ( .A1(n6022), .A2(n6021), .ZN(n6498) );
  OAI222_X1 U7554 ( .A1(n8578), .A2(n6495), .B1(n8582), .B2(n6493), .C1(
        P2_U3151), .C2(n6498), .ZN(P2_U3292) );
  NAND2_X1 U7555 ( .A1(n4583), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6023) );
  XNOR2_X1 U7556 ( .A(n6023), .B(n5057), .ZN(n6919) );
  OAI222_X1 U7557 ( .A1(n8578), .A2(n6918), .B1(n8576), .B2(n6917), .C1(
        P2_U3151), .C2(n6919), .ZN(P2_U3288) );
  INV_X1 U7558 ( .A(n9817), .ZN(n6627) );
  INV_X1 U7559 ( .A(n6627), .ZN(n9814) );
  OAI222_X1 U7560 ( .A1(n6025), .A2(P1_U3086), .B1(n9820), .B2(n6917), .C1(
        n6024), .C2(n9814), .ZN(P1_U3348) );
  AND2_X1 U7561 ( .A1(n6286), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6051) );
  INV_X1 U7562 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n9600) );
  NOR2_X1 U7563 ( .A1(n6050), .A2(n9600), .ZN(P2_U3258) );
  INV_X1 U7564 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n9612) );
  NOR2_X1 U7565 ( .A1(n6050), .A2(n9612), .ZN(P2_U3243) );
  INV_X1 U7566 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n6028) );
  NOR2_X1 U7567 ( .A1(n6050), .A2(n6028), .ZN(P2_U3252) );
  INV_X1 U7568 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n9683) );
  NOR2_X1 U7569 ( .A1(n6050), .A2(n9683), .ZN(P2_U3234) );
  INV_X1 U7570 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6029) );
  NOR2_X1 U7571 ( .A1(n6050), .A2(n6029), .ZN(P2_U3235) );
  INV_X1 U7572 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n9603) );
  NOR2_X1 U7573 ( .A1(n6050), .A2(n9603), .ZN(P2_U3263) );
  INV_X1 U7574 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n9677) );
  NOR2_X1 U7575 ( .A1(n6050), .A2(n9677), .ZN(P2_U3238) );
  INV_X1 U7576 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n9641) );
  NOR2_X1 U7577 ( .A1(n6050), .A2(n9641), .ZN(P2_U3240) );
  INV_X1 U7578 ( .A(n7036), .ZN(n6034) );
  OR2_X1 U7579 ( .A1(n6030), .A2(n6279), .ZN(n6031) );
  XNOR2_X1 U7580 ( .A(n6031), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7037) );
  INV_X1 U7581 ( .A(n7037), .ZN(n6454) );
  OAI222_X1 U7582 ( .A1(n8578), .A2(n6032), .B1(n8576), .B2(n6034), .C1(
        P2_U3151), .C2(n6454), .ZN(P2_U3287) );
  OAI222_X1 U7583 ( .A1(n6035), .A2(P1_U3086), .B1(n9820), .B2(n6034), .C1(
        n6033), .C2(n9817), .ZN(P1_U3347) );
  AND2_X1 U7584 ( .A1(n6036), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U7585 ( .A1(n6036), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U7586 ( .A1(n6036), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U7587 ( .A1(n6036), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U7588 ( .A1(n6036), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U7589 ( .A1(n6036), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U7590 ( .A1(n6036), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  NAND2_X1 U7591 ( .A1(n6037), .A2(n9007), .ZN(n6082) );
  OR2_X1 U7592 ( .A1(n8931), .A2(n6181), .ZN(n6038) );
  NAND2_X1 U7593 ( .A1(n6038), .A2(n5307), .ZN(n6081) );
  AND2_X1 U7594 ( .A1(n6082), .A2(n6081), .ZN(n9945) );
  NOR2_X1 U7595 ( .A1(n9945), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U7596 ( .A(n6365), .ZN(n6117) );
  INV_X1 U7597 ( .A(n7087), .ZN(n6044) );
  OAI222_X1 U7598 ( .A1(n6117), .A2(P1_U3086), .B1(n9820), .B2(n6044), .C1(
        n6039), .C2(n9814), .ZN(P1_U3346) );
  NAND2_X1 U7599 ( .A1(n6041), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6042) );
  MUX2_X1 U7600 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6042), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n6043) );
  AND2_X1 U7601 ( .A1(n6040), .A2(n6043), .ZN(n7088) );
  OAI222_X1 U7602 ( .A1(n8578), .A2(n6045), .B1(n8576), .B2(n6044), .C1(
        P2_U3151), .C2(n6684), .ZN(P2_U3286) );
  INV_X1 U7603 ( .A(n7146), .ZN(n6049) );
  AOI22_X1 U7604 ( .A1(n9832), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n6627), .ZN(n6046) );
  OAI21_X1 U7605 ( .B1(n6049), .B2(n9820), .A(n6046), .ZN(P1_U3345) );
  NAND2_X1 U7606 ( .A1(n6040), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6047) );
  XNOR2_X1 U7607 ( .A(n6047), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7147) );
  INV_X1 U7608 ( .A(n7147), .ZN(n6683) );
  OAI222_X1 U7609 ( .A1(n8582), .A2(n6049), .B1(n6683), .B2(P2_U3151), .C1(
        n6048), .C2(n8578), .ZN(P2_U3285) );
  INV_X1 U7610 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6053) );
  AND3_X1 U7611 ( .A1(n6027), .A2(n6051), .A3(n8580), .ZN(n6052) );
  AOI21_X1 U7612 ( .B1(n6036), .B2(n6053), .A(n6052), .ZN(P2_U3377) );
  INV_X1 U7613 ( .A(n6026), .ZN(n6054) );
  NOR4_X1 U7614 ( .A1(n6055), .A2(n6054), .A3(n7071), .A4(P2_U3151), .ZN(n6056) );
  AOI21_X1 U7615 ( .B1(n6036), .B2(n5043), .A(n6056), .ZN(P2_U3376) );
  NAND2_X1 U7616 ( .A1(n10113), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6058) );
  OAI21_X1 U7617 ( .B1(n10113), .B2(n6059), .A(n6058), .ZN(P1_U3439) );
  AND2_X1 U7618 ( .A1(n6036), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U7619 ( .A1(n6036), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U7620 ( .A1(n6036), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U7621 ( .A1(n6036), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U7622 ( .A1(n6036), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U7623 ( .A1(n6036), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U7624 ( .A1(n6036), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U7625 ( .A1(n6036), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U7626 ( .A1(n6036), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U7627 ( .A1(n6036), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U7628 ( .A1(n6036), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U7629 ( .A1(n6036), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U7630 ( .A1(n6036), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U7631 ( .A1(n6036), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U7632 ( .A1(n6036), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  INV_X1 U7633 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7634 ( .A1(n10121), .A2(P1_U3973), .ZN(n6060) );
  OAI21_X1 U7635 ( .B1(P1_U3973), .B2(n6061), .A(n6060), .ZN(P1_U3554) );
  INV_X1 U7636 ( .A(n7265), .ZN(n6066) );
  OR2_X1 U7637 ( .A1(n6062), .A2(n6279), .ZN(n6063) );
  XNOR2_X1 U7638 ( .A(n6063), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7266) );
  INV_X1 U7639 ( .A(n7266), .ZN(n6994) );
  OAI222_X1 U7640 ( .A1(n8578), .A2(n6064), .B1(n8576), .B2(n6066), .C1(
        P2_U3151), .C2(n6994), .ZN(P2_U3284) );
  INV_X1 U7641 ( .A(n9978), .ZN(n6358) );
  OAI222_X1 U7642 ( .A1(n6358), .A2(P1_U3086), .B1(n9820), .B2(n6066), .C1(
        n6065), .C2(n9814), .ZN(P1_U3344) );
  NAND2_X1 U7643 ( .A1(n6067), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7644 ( .A1(n6072), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7645 ( .A1(n5241), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7646 ( .A1(n9030), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n6071) );
  OAI21_X1 U7647 ( .B1(n9094), .B2(n9030), .A(n6071), .ZN(P1_U3585) );
  INV_X1 U7648 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7943) );
  NAND2_X1 U7649 ( .A1(n6067), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7650 ( .A1(n6072), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7651 ( .A1(n5241), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6073) );
  INV_X1 U7652 ( .A(n9149), .ZN(n6076) );
  NAND2_X1 U7653 ( .A1(n6076), .A2(P1_U3973), .ZN(n6077) );
  OAI21_X1 U7654 ( .B1(n7943), .B2(P1_U3973), .A(n6077), .ZN(P1_U3584) );
  INV_X1 U7655 ( .A(n7269), .ZN(n6122) );
  OR2_X1 U7656 ( .A1(n6078), .A2(n6279), .ZN(n6079) );
  XNOR2_X1 U7657 ( .A(n6079), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7270) );
  INV_X1 U7658 ( .A(n7270), .ZN(n7201) );
  OAI222_X1 U7659 ( .A1(n8582), .A2(n6122), .B1(n7201), .B2(P2_U3151), .C1(
        n6080), .C2(n8578), .ZN(P2_U3283) );
  INV_X1 U7660 ( .A(n6081), .ZN(n6083) );
  NAND2_X1 U7661 ( .A1(n6083), .A2(n6082), .ZN(n9933) );
  OR2_X1 U7662 ( .A1(n5872), .A2(n9924), .ZN(n6084) );
  NOR2_X2 U7663 ( .A1(n9933), .A2(n6084), .ZN(n9983) );
  INV_X1 U7664 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6085) );
  AOI22_X1 U7665 ( .A1(n6365), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n6085), .B2(
        n6117), .ZN(n6099) );
  INV_X1 U7666 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6086) );
  MUX2_X1 U7667 ( .A(n6086), .B(P1_REG2_REG_2__SCAN_IN), .S(n6100), .Z(n9042)
         );
  INV_X1 U7668 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6824) );
  AND2_X1 U7669 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9025) );
  INV_X1 U7670 ( .A(n6101), .ZN(n9017) );
  NAND2_X1 U7671 ( .A1(n9017), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7672 ( .A1(n9018), .A2(n6087), .ZN(n9041) );
  NAND2_X1 U7673 ( .A1(n9042), .A2(n9041), .ZN(n9040) );
  INV_X1 U7674 ( .A(n6100), .ZN(n9036) );
  NAND2_X1 U7675 ( .A1(n9036), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7676 ( .A1(n9040), .A2(n6088), .ZN(n9054) );
  INV_X1 U7677 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6089) );
  MUX2_X1 U7678 ( .A(n6089), .B(P1_REG2_REG_3__SCAN_IN), .S(n6104), .Z(n9055)
         );
  NAND2_X1 U7679 ( .A1(n9054), .A2(n9055), .ZN(n9053) );
  INV_X1 U7680 ( .A(n6104), .ZN(n9052) );
  NAND2_X1 U7681 ( .A1(n9052), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7682 ( .A1(n9053), .A2(n6090), .ZN(n9935) );
  MUX2_X1 U7683 ( .A(n5267), .B(P1_REG2_REG_4__SCAN_IN), .S(n6106), .Z(n9936)
         );
  INV_X1 U7684 ( .A(n6106), .ZN(n9940) );
  NAND2_X1 U7685 ( .A1(n9940), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6091) );
  INV_X1 U7686 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6093) );
  AOI22_X1 U7687 ( .A1(n9953), .A2(n6093), .B1(P1_REG2_REG_5__SCAN_IN), .B2(
        n6092), .ZN(n9955) );
  INV_X1 U7688 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6095) );
  AOI22_X1 U7689 ( .A1(n9964), .A2(n6095), .B1(P1_REG2_REG_6__SCAN_IN), .B2(
        n6094), .ZN(n9966) );
  NOR2_X1 U7690 ( .A1(n4547), .A2(n9966), .ZN(n9965) );
  AOI21_X1 U7691 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n9964), .A(n9965), .ZN(
        n9839) );
  NAND2_X1 U7692 ( .A1(n9837), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6096) );
  OAI21_X1 U7693 ( .B1(n9837), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6096), .ZN(
        n9840) );
  NOR2_X1 U7694 ( .A1(n9839), .A2(n9840), .ZN(n9838) );
  NAND2_X1 U7695 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n9856), .ZN(n6097) );
  OAI21_X1 U7696 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9856), .A(n6097), .ZN(
        n9854) );
  OAI21_X1 U7697 ( .B1(n6099), .B2(n6098), .A(n6357), .ZN(n6119) );
  NOR2_X2 U7698 ( .A1(n9933), .A2(n9027), .ZN(n10043) );
  INV_X1 U7699 ( .A(n10043), .ZN(n9070) );
  INV_X1 U7700 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10265) );
  AOI22_X1 U7701 ( .A1(n6365), .A2(P1_REG1_REG_9__SCAN_IN), .B1(n10265), .B2(
        n6117), .ZN(n6113) );
  INV_X1 U7702 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10254) );
  MUX2_X1 U7703 ( .A(n10254), .B(P1_REG1_REG_2__SCAN_IN), .S(n6100), .Z(n9039)
         );
  INV_X1 U7704 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10252) );
  MUX2_X1 U7705 ( .A(n10252), .B(P1_REG1_REG_1__SCAN_IN), .S(n6101), .Z(n9016)
         );
  AND2_X1 U7706 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9015) );
  NAND2_X1 U7707 ( .A1(n9016), .A2(n9015), .ZN(n9014) );
  NAND2_X1 U7708 ( .A1(n9017), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7709 ( .A1(n9014), .A2(n6102), .ZN(n9038) );
  NAND2_X1 U7710 ( .A1(n9039), .A2(n9038), .ZN(n9037) );
  NAND2_X1 U7711 ( .A1(n9036), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7712 ( .A1(n9037), .A2(n6103), .ZN(n9047) );
  INV_X1 U7713 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10256) );
  MUX2_X1 U7714 ( .A(n10256), .B(P1_REG1_REG_3__SCAN_IN), .S(n6104), .Z(n9048)
         );
  NAND2_X1 U7715 ( .A1(n9047), .A2(n9048), .ZN(n9046) );
  NAND2_X1 U7716 ( .A1(n9052), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7717 ( .A1(n9046), .A2(n6105), .ZN(n9938) );
  INV_X1 U7718 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10258) );
  MUX2_X1 U7719 ( .A(n10258), .B(P1_REG1_REG_4__SCAN_IN), .S(n6106), .Z(n9939)
         );
  NAND2_X1 U7720 ( .A1(n9940), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7721 ( .A1(n9937), .A2(n6107), .ZN(n9951) );
  INV_X1 U7722 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10260) );
  MUX2_X1 U7723 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10260), .S(n9953), .Z(n9952)
         );
  NAND2_X1 U7724 ( .A1(n9951), .A2(n9952), .ZN(n9950) );
  NAND2_X1 U7725 ( .A1(n9953), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6108) );
  INV_X1 U7726 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6109) );
  MUX2_X1 U7727 ( .A(n6109), .B(P1_REG1_REG_6__SCAN_IN), .S(n9964), .Z(n9969)
         );
  NOR2_X1 U7728 ( .A1(n9970), .A2(n9969), .ZN(n9968) );
  INV_X1 U7729 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6110) );
  MUX2_X1 U7730 ( .A(n6110), .B(P1_REG1_REG_7__SCAN_IN), .S(n9837), .Z(n9844)
         );
  NOR2_X1 U7731 ( .A1(n9843), .A2(n9844), .ZN(n9842) );
  AOI21_X1 U7732 ( .B1(n9837), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9842), .ZN(
        n9858) );
  INV_X1 U7733 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6111) );
  MUX2_X1 U7734 ( .A(n6111), .B(P1_REG1_REG_8__SCAN_IN), .S(n9856), .Z(n9859)
         );
  NOR2_X1 U7735 ( .A1(n9858), .A2(n9859), .ZN(n9857) );
  NAND2_X1 U7736 ( .A1(n6113), .A2(n6112), .ZN(n6364) );
  OAI21_X1 U7737 ( .B1(n6113), .B2(n6112), .A(n6364), .ZN(n6114) );
  INV_X1 U7738 ( .A(n9924), .ZN(n9024) );
  NAND2_X1 U7739 ( .A1(n6114), .A2(n9988), .ZN(n6116) );
  AND2_X1 U7740 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7225) );
  AOI21_X1 U7741 ( .B1(n9945), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7225), .ZN(
        n6115) );
  OAI211_X1 U7742 ( .C1(n9070), .C2(n6117), .A(n6116), .B(n6115), .ZN(n6118)
         );
  AOI21_X1 U7743 ( .B1(n9983), .B2(n6119), .A(n6118), .ZN(n6120) );
  INV_X1 U7744 ( .A(n6120), .ZN(P1_U3252) );
  INV_X1 U7745 ( .A(n7120), .ZN(n6370) );
  OAI222_X1 U7746 ( .A1(P1_U3086), .A2(n6370), .B1(n9820), .B2(n6122), .C1(
        n6121), .C2(n9814), .ZN(P1_U3343) );
  INV_X1 U7747 ( .A(n7319), .ZN(n6153) );
  AOI22_X1 U7748 ( .A1(n10003), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n6627), .ZN(n6123) );
  OAI21_X1 U7749 ( .B1(n6153), .B2(n9820), .A(n6123), .ZN(P1_U3342) );
  NAND2_X1 U7750 ( .A1(P2_U3893), .A2(n6295), .ZN(n8264) );
  MUX2_X1 U7751 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8255), .Z(n6125) );
  XNOR2_X1 U7752 ( .A(n6125), .B(n6213), .ZN(n6212) );
  INV_X1 U7753 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6432) );
  MUX2_X1 U7754 ( .A(n6432), .B(n4931), .S(n8255), .Z(n10276) );
  AND2_X1 U7755 ( .A1(n10276), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10278) );
  INV_X1 U7756 ( .A(n6125), .ZN(n6126) );
  OAI22_X1 U7757 ( .A1(n6212), .A2(n10278), .B1(n6477), .B2(n6126), .ZN(n6203)
         );
  MUX2_X1 U7758 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8255), .Z(n6201) );
  XOR2_X1 U7759 ( .A(n6482), .B(n6201), .Z(n6202) );
  XNOR2_X1 U7760 ( .A(n6203), .B(n6202), .ZN(n6150) );
  OR2_X1 U7761 ( .A1(n6295), .A2(P2_U3151), .ZN(n8570) );
  INV_X1 U7762 ( .A(n8570), .ZN(n6142) );
  INV_X1 U7763 ( .A(n8267), .ZN(n8246) );
  NAND2_X1 U7764 ( .A1(n6213), .A2(n6129), .ZN(n6128) );
  NAND2_X1 U7765 ( .A1(n6128), .A2(n6127), .ZN(n6214) );
  INV_X1 U7766 ( .A(n6129), .ZN(n6130) );
  AOI21_X1 U7767 ( .B1(n6214), .B2(P2_REG1_REG_1__SCAN_IN), .A(n6130), .ZN(
        n6187) );
  XOR2_X1 U7768 ( .A(n6188), .B(n6187), .Z(n6138) );
  XNOR2_X1 U7769 ( .A(n6482), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7770 ( .A1(n6131), .A2(n6132), .ZN(n6216) );
  INV_X1 U7771 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6601) );
  INV_X1 U7772 ( .A(n6132), .ZN(n6133) );
  AOI21_X1 U7773 ( .B1(n6135), .B2(n6134), .A(n4605), .ZN(n6137) );
  INV_X1 U7774 ( .A(n10280), .ZN(n6136) );
  OAI22_X1 U7775 ( .A1(n8246), .A2(n6138), .B1(n6137), .B2(n8268), .ZN(n6148)
         );
  INV_X1 U7776 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6139) );
  NOR2_X1 U7777 ( .A1(n8204), .A2(n6139), .ZN(n6147) );
  NOR2_X1 U7778 ( .A1(n8255), .A2(P2_U3151), .ZN(n8573) );
  AND2_X1 U7779 ( .A1(n8573), .A2(n6295), .ZN(n6140) );
  NAND2_X1 U7780 ( .A1(n6141), .A2(n6140), .ZN(n6145) );
  NAND2_X1 U7781 ( .A1(n6143), .A2(n6142), .ZN(n6144) );
  OAI22_X1 U7782 ( .A1(n10283), .A2(n6482), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6619), .ZN(n6146) );
  NOR3_X1 U7783 ( .A1(n6148), .A2(n6147), .A3(n6146), .ZN(n6149) );
  OAI21_X1 U7784 ( .B1(n8264), .B2(n6150), .A(n6149), .ZN(P2_U3184) );
  INV_X1 U7785 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U7786 ( .A1(n6151), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6152) );
  XNOR2_X1 U7787 ( .A(n6152), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7320) );
  INV_X1 U7788 ( .A(n7320), .ZN(n8122) );
  OAI222_X1 U7789 ( .A1(n8578), .A2(n6154), .B1(n8576), .B2(n6153), .C1(
        P2_U3151), .C2(n8122), .ZN(P2_U3282) );
  NAND2_X1 U7790 ( .A1(n6156), .A2(n6155), .ZN(n6159) );
  INV_X1 U7791 ( .A(n6157), .ZN(n6158) );
  INV_X1 U7792 ( .A(n6160), .ZN(n6721) );
  OR2_X1 U7793 ( .A1(n6161), .A2(n6721), .ZN(n6173) );
  NOR2_X1 U7794 ( .A1(n6173), .A2(n6172), .ZN(n6162) );
  INV_X1 U7795 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6171) );
  INV_X1 U7796 ( .A(n6827), .ZN(n7413) );
  AND2_X1 U7797 ( .A1(n10121), .A2(n7413), .ZN(n8940) );
  NOR2_X1 U7798 ( .A1(n6820), .A2(n8940), .ZN(n8872) );
  NAND2_X1 U7799 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  NAND2_X1 U7800 ( .A1(n6169), .A2(n6165), .ZN(n6166) );
  OR2_X1 U7801 ( .A1(n6166), .A2(n7408), .ZN(n10116) );
  NAND2_X1 U7802 ( .A1(n9005), .A2(n8995), .ZN(n8861) );
  INV_X1 U7803 ( .A(n6904), .ZN(n8997) );
  NAND2_X1 U7804 ( .A1(n6167), .A2(n8997), .ZN(n8737) );
  NOR2_X1 U7805 ( .A1(n10231), .A2(n10203), .ZN(n6168) );
  INV_X1 U7806 ( .A(n6717), .ZN(n6731) );
  OAI222_X1 U7807 ( .A1(n7413), .A2(n6169), .B1(n8872), .B2(n6168), .C1(n10236), .C2(n6731), .ZN(n6175) );
  NAND2_X1 U7808 ( .A1(n6175), .A2(n10251), .ZN(n6170) );
  OAI21_X1 U7809 ( .B1(n10251), .B2(n6171), .A(n6170), .ZN(P1_U3453) );
  INV_X1 U7810 ( .A(n6172), .ZN(n6720) );
  INV_X1 U7811 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9923) );
  NAND2_X1 U7812 ( .A1(n6175), .A2(n10274), .ZN(n6176) );
  OAI21_X1 U7813 ( .B1(n10274), .B2(n9923), .A(n6176), .ZN(P1_U3522) );
  OR2_X1 U7814 ( .A1(n6178), .A2(n6177), .ZN(n6179) );
  NAND2_X1 U7815 ( .A1(n6180), .A2(n6179), .ZN(n9026) );
  INV_X1 U7816 ( .A(n6181), .ZN(n6182) );
  NAND3_X1 U7817 ( .A1(n6183), .A2(P1_STATE_REG_SCAN_IN), .A3(n6182), .ZN(
        n6438) );
  OAI22_X1 U7818 ( .A1(n8729), .A2(n6731), .B1(n8689), .B2(n7413), .ZN(n6184)
         );
  AOI21_X1 U7819 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n6438), .A(n6184), .ZN(
        n6185) );
  OAI21_X1 U7820 ( .B1(n9026), .B2(n8733), .A(n6185), .ZN(P1_U3232) );
  INV_X1 U7821 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6211) );
  INV_X1 U7822 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6510) );
  MUX2_X1 U7823 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6510), .S(n6640), .Z(n6190)
         );
  INV_X1 U7824 ( .A(n6482), .ZN(n6186) );
  INV_X1 U7825 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10371) );
  NAND2_X1 U7826 ( .A1(n6189), .A2(n6190), .ZN(n6242) );
  OAI21_X1 U7827 ( .B1(n6190), .B2(n6189), .A(n6242), .ZN(n6200) );
  NOR2_X1 U7828 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6511), .ZN(n6662) );
  INV_X1 U7829 ( .A(n6662), .ZN(n6191) );
  OAI21_X1 U7830 ( .B1(n10283), .B2(n6640), .A(n6191), .ZN(n6199) );
  NOR2_X1 U7831 ( .A1(n6192), .A2(n6231), .ZN(n6193) );
  NOR2_X1 U7832 ( .A1(n6193), .A2(n5119), .ZN(n6224) );
  NAND2_X1 U7833 ( .A1(n6224), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6225) );
  INV_X1 U7834 ( .A(n6193), .ZN(n6194) );
  XNOR2_X1 U7835 ( .A(n6640), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n6195) );
  INV_X1 U7836 ( .A(n6247), .ZN(n6197) );
  NAND3_X1 U7837 ( .A1(n6225), .A2(n6195), .A3(n6194), .ZN(n6196) );
  AOI21_X1 U7838 ( .B1(n6197), .B2(n6196), .A(n8268), .ZN(n6198) );
  AOI211_X1 U7839 ( .C1(n8267), .C2(n6200), .A(n6199), .B(n6198), .ZN(n6210)
         );
  AOI22_X1 U7840 ( .A1(n6203), .A2(n6202), .B1(n6201), .B2(n6482), .ZN(n6234)
         );
  MUX2_X1 U7841 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8255), .Z(n6204) );
  XOR2_X1 U7842 ( .A(n6498), .B(n6204), .Z(n6233) );
  NAND2_X1 U7843 ( .A1(n6234), .A2(n6233), .ZN(n6232) );
  INV_X1 U7844 ( .A(n6204), .ZN(n6205) );
  NAND2_X1 U7845 ( .A1(n6205), .A2(n6231), .ZN(n6206) );
  AND2_X1 U7846 ( .A1(n6232), .A2(n6206), .ZN(n6208) );
  MUX2_X1 U7847 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8255), .Z(n6239) );
  INV_X1 U7848 ( .A(n6640), .ZN(n6243) );
  XNOR2_X1 U7849 ( .A(n6239), .B(n6243), .ZN(n6207) );
  NAND3_X1 U7850 ( .A1(n6232), .A2(n6206), .A3(n6207), .ZN(n6240) );
  OAI211_X1 U7851 ( .C1(n6208), .C2(n6207), .A(n10279), .B(n6240), .ZN(n6209)
         );
  OAI211_X1 U7852 ( .C1(n8204), .C2(n6211), .A(n6210), .B(n6209), .ZN(P2_U3186) );
  XNOR2_X1 U7853 ( .A(n6212), .B(n10278), .ZN(n6222) );
  INV_X1 U7854 ( .A(n8204), .ZN(n10275) );
  INV_X1 U7855 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6563) );
  OAI22_X1 U7856 ( .A1(n10283), .A2(n6213), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6563), .ZN(n6220) );
  INV_X1 U7857 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6559) );
  XNOR2_X1 U7858 ( .A(n6214), .B(n6559), .ZN(n6218) );
  AOI21_X1 U7859 ( .B1(n6601), .B2(n6216), .A(n6215), .ZN(n6217) );
  OAI22_X1 U7860 ( .A1(n8246), .A2(n6218), .B1(n6217), .B2(n8268), .ZN(n6219)
         );
  AOI211_X1 U7861 ( .C1(n10275), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n6220), .B(
        n6219), .ZN(n6221) );
  OAI21_X1 U7862 ( .B1(n8264), .B2(n6222), .A(n6221), .ZN(P2_U3183) );
  INV_X1 U7863 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6238) );
  NOR2_X1 U7864 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10295), .ZN(n6517) );
  XNOR2_X1 U7865 ( .A(n6223), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n6229) );
  INV_X1 U7866 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10298) );
  INV_X1 U7867 ( .A(n6224), .ZN(n6227) );
  INV_X1 U7868 ( .A(n6225), .ZN(n6226) );
  AOI21_X1 U7869 ( .B1(n10298), .B2(n6227), .A(n6226), .ZN(n6228) );
  OAI22_X1 U7870 ( .A1(n8246), .A2(n6229), .B1(n6228), .B2(n8268), .ZN(n6230)
         );
  AOI211_X1 U7871 ( .C1(n6231), .C2(n8202), .A(n6517), .B(n6230), .ZN(n6237)
         );
  OAI21_X1 U7872 ( .B1(n6234), .B2(n6233), .A(n6232), .ZN(n6235) );
  NAND2_X1 U7873 ( .A1(n6235), .A2(n10279), .ZN(n6236) );
  OAI211_X1 U7874 ( .C1(n6238), .C2(n8204), .A(n6237), .B(n6236), .ZN(P2_U3185) );
  INV_X1 U7875 ( .A(n6239), .ZN(n6241) );
  OAI21_X1 U7876 ( .B1(n6243), .B2(n6241), .A(n6240), .ZN(n6329) );
  INV_X1 U7877 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6657) );
  INV_X1 U7878 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6652) );
  MUX2_X1 U7879 ( .A(n6657), .B(n6652), .S(n8255), .Z(n6326) );
  XNOR2_X1 U7880 ( .A(n6326), .B(n6778), .ZN(n6328) );
  XNOR2_X1 U7881 ( .A(n6329), .B(n6328), .ZN(n6257) );
  OAI21_X1 U7882 ( .B1(n6244), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6334), .ZN(
        n6255) );
  INV_X1 U7883 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6246) );
  NOR2_X1 U7884 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6653), .ZN(n6791) );
  AOI21_X1 U7885 ( .B1(n8202), .B2(n6248), .A(n6791), .ZN(n6245) );
  OAI21_X1 U7886 ( .B1(n6246), .B2(n8204), .A(n6245), .ZN(n6254) );
  AOI21_X1 U7887 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n6640), .A(n6247), .ZN(
        n6249) );
  NOR2_X1 U7888 ( .A1(n6249), .A2(n6248), .ZN(n6338) );
  NAND2_X1 U7889 ( .A1(n6249), .A2(n6248), .ZN(n6250) );
  AOI21_X1 U7890 ( .B1(n6251), .B2(n6657), .A(n6339), .ZN(n6252) );
  NOR2_X1 U7891 ( .A1(n6252), .A2(n8268), .ZN(n6253) );
  AOI211_X1 U7892 ( .C1(n8267), .C2(n6255), .A(n6254), .B(n6253), .ZN(n6256)
         );
  OAI21_X1 U7893 ( .B1(n8264), .B2(n6257), .A(n6256), .ZN(P2_U3187) );
  OR2_X1 U7894 ( .A1(n6271), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U7895 ( .A1(n6027), .A2(n8580), .ZN(n6258) );
  NAND2_X1 U7896 ( .A1(n6259), .A2(n6258), .ZN(n6554) );
  NOR2_X1 U7897 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6263) );
  NOR4_X1 U7898 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6262) );
  NOR4_X1 U7899 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6261) );
  NOR4_X1 U7900 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n6260) );
  NAND4_X1 U7901 ( .A1(n6263), .A2(n6262), .A3(n6261), .A4(n6260), .ZN(n6269)
         );
  NOR4_X1 U7902 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6267) );
  NOR4_X1 U7903 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6266) );
  NOR4_X1 U7904 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n6265) );
  NOR4_X1 U7905 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6264) );
  NAND4_X1 U7906 ( .A1(n6267), .A2(n6266), .A3(n6265), .A4(n6264), .ZN(n6268)
         );
  NOR2_X1 U7907 ( .A1(n6269), .A2(n6268), .ZN(n6270) );
  OR2_X1 U7908 ( .A1(n6271), .A2(n6270), .ZN(n6316) );
  NAND2_X1 U7909 ( .A1(n6554), .A2(n6316), .ZN(n6274) );
  NAND2_X1 U7910 ( .A1(n8580), .A2(n6026), .ZN(n6272) );
  AND2_X2 U7911 ( .A1(n6273), .A2(n6272), .ZN(n6467) );
  NOR2_X1 U7912 ( .A1(n6274), .A2(n6467), .ZN(n6294) );
  NAND2_X1 U7913 ( .A1(n7455), .A2(n7872), .ZN(n6532) );
  INV_X1 U7914 ( .A(n6316), .ZN(n6284) );
  INV_X1 U7915 ( .A(n6554), .ZN(n6420) );
  NAND2_X1 U7916 ( .A1(n6467), .A2(n6420), .ZN(n6422) );
  NAND3_X1 U7917 ( .A1(n7358), .A2(n7850), .A3(n10356), .ZN(n6318) );
  NAND2_X1 U7918 ( .A1(n7865), .A2(n7455), .ZN(n6548) );
  INV_X1 U7919 ( .A(n6548), .ZN(n6283) );
  NAND2_X1 U7920 ( .A1(n6318), .A2(n8308), .ZN(n7356) );
  OAI21_X1 U7921 ( .B1(n6284), .B2(n6422), .A(n7356), .ZN(n6289) );
  INV_X1 U7922 ( .A(n6469), .ZN(n6285) );
  OR2_X1 U7923 ( .A1(n7850), .A2(n6285), .ZN(n6424) );
  AND3_X1 U7924 ( .A1(n6424), .A2(n6287), .A3(n6286), .ZN(n6288) );
  OAI211_X1 U7925 ( .C1(n6294), .C2(n7358), .A(n6289), .B(n6288), .ZN(n6290)
         );
  NAND2_X1 U7926 ( .A1(n6290), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6293) );
  INV_X1 U7927 ( .A(n6315), .ZN(n6322) );
  NOR2_X1 U7928 ( .A1(n7359), .A2(n6322), .ZN(n7870) );
  INV_X1 U7929 ( .A(n6294), .ZN(n6291) );
  NAND2_X1 U7930 ( .A1(n7870), .A2(n6291), .ZN(n6292) );
  NOR2_X1 U7931 ( .A1(n8081), .A2(P2_U3151), .ZN(n6570) );
  INV_X1 U7932 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6427) );
  INV_X1 U7933 ( .A(n7359), .ZN(n6428) );
  NAND2_X1 U7934 ( .A1(n7357), .A2(n6428), .ZN(n6509) );
  INV_X1 U7935 ( .A(n6509), .ZN(n6296) );
  INV_X1 U7936 ( .A(n6295), .ZN(n7869) );
  XNOR2_X1 U7937 ( .A(n7869), .B(n8255), .ZN(n6543) );
  INV_X1 U7938 ( .A(n6543), .ZN(n6508) );
  NAND2_X1 U7939 ( .A1(n6300), .A2(n6301), .ZN(n8564) );
  NAND2_X1 U7940 ( .A1(n7534), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6306) );
  OR2_X1 U7941 ( .A1(n6499), .A2(n6427), .ZN(n6310) );
  OR2_X1 U7942 ( .A1(n6501), .A2(n4931), .ZN(n6309) );
  NAND2_X1 U7943 ( .A1(n7534), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6308) );
  NAND4_X1 U7944 ( .A1(n6311), .A2(n6310), .A3(n6309), .A4(n6308), .ZN(n6536)
         );
  NAND2_X1 U7945 ( .A1(n5201), .A2(SI_0_), .ZN(n6312) );
  XNOR2_X1 U7946 ( .A(n6312), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8583) );
  MUX2_X1 U7947 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8583), .S(n6476), .Z(n10304)
         );
  AND2_X1 U7948 ( .A1(n6313), .A2(n10304), .ZN(n6538) );
  NAND2_X1 U7949 ( .A1(n6536), .A2(n6478), .ZN(n7720) );
  AND2_X1 U7950 ( .A1(n7721), .A2(n7720), .ZN(n10300) );
  INV_X1 U7951 ( .A(n7358), .ZN(n6314) );
  NAND2_X1 U7952 ( .A1(n7357), .A2(n6314), .ZN(n6321) );
  INV_X1 U7953 ( .A(n6423), .ZN(n6317) );
  INV_X1 U7954 ( .A(n6318), .ZN(n6319) );
  NAND2_X1 U7955 ( .A1(n7361), .A2(n6319), .ZN(n6320) );
  NAND2_X1 U7956 ( .A1(n7361), .A2(n10366), .ZN(n6323) );
  OAI22_X1 U7957 ( .A1(n10300), .A2(n8096), .B1(n8076), .B2(n6478), .ZN(n6324)
         );
  AOI21_X1 U7958 ( .B1(n8092), .B2(n8116), .A(n6324), .ZN(n6325) );
  OAI21_X1 U7959 ( .B1(n6570), .B2(n6427), .A(n6325), .ZN(P2_U3172) );
  INV_X1 U7960 ( .A(n6326), .ZN(n6327) );
  AOI22_X1 U7961 ( .A1(n6329), .A2(n6328), .B1(n6327), .B2(n6778), .ZN(n6332)
         );
  MUX2_X1 U7962 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8255), .Z(n6330) );
  NOR2_X1 U7963 ( .A1(n6330), .A2(n6868), .ZN(n6392) );
  AOI21_X1 U7964 ( .B1(n6330), .B2(n6868), .A(n6392), .ZN(n6331) );
  NAND2_X1 U7965 ( .A1(n6332), .A2(n6331), .ZN(n6398) );
  OAI21_X1 U7966 ( .B1(n6332), .B2(n6331), .A(n6398), .ZN(n6353) );
  INV_X1 U7967 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6351) );
  INV_X1 U7968 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10377) );
  AOI22_X1 U7969 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(n6868), .B1(n6348), .B2(
        n10377), .ZN(n6337) );
  NAND2_X1 U7970 ( .A1(n6333), .A2(n6778), .ZN(n6335) );
  NAND2_X1 U7971 ( .A1(n6337), .A2(n6336), .ZN(n6400) );
  OAI21_X1 U7972 ( .B1(n6337), .B2(n6336), .A(n6400), .ZN(n6346) );
  INV_X1 U7973 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6340) );
  NOR2_X1 U7974 ( .A1(n6348), .A2(n6340), .ZN(n6388) );
  INV_X1 U7975 ( .A(n6388), .ZN(n6341) );
  OAI21_X1 U7976 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n6868), .A(n6341), .ZN(
        n6342) );
  NOR2_X1 U7977 ( .A1(n6343), .A2(n6342), .ZN(n6389) );
  AOI21_X1 U7978 ( .B1(n6343), .B2(n6342), .A(n6389), .ZN(n6344) );
  NOR2_X1 U7979 ( .A1(n6344), .A2(n8268), .ZN(n6345) );
  AOI21_X1 U7980 ( .B1(n6346), .B2(n8267), .A(n6345), .ZN(n6350) );
  NAND2_X1 U7981 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3151), .ZN(n6911) );
  INV_X1 U7982 ( .A(n6911), .ZN(n6347) );
  AOI21_X1 U7983 ( .B1(n8202), .B2(n6348), .A(n6347), .ZN(n6349) );
  OAI211_X1 U7984 ( .C1(n6351), .C2(n8204), .A(n6350), .B(n6349), .ZN(n6352)
         );
  AOI21_X1 U7985 ( .B1(n6353), .B2(n10279), .A(n6352), .ZN(n6354) );
  INV_X1 U7986 ( .A(n6354), .ZN(P2_U3188) );
  INV_X1 U7987 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6355) );
  AOI22_X1 U7988 ( .A1(n7120), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n6355), .B2(
        n6370), .ZN(n6361) );
  NAND2_X1 U7989 ( .A1(n9832), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6356) );
  OAI21_X1 U7990 ( .B1(n9832), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6356), .ZN(
        n9828) );
  OAI21_X1 U7991 ( .B1(n6365), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6357), .ZN(
        n9829) );
  NOR2_X1 U7992 ( .A1(n9828), .A2(n9829), .ZN(n9827) );
  INV_X1 U7993 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6359) );
  AOI22_X1 U7994 ( .A1(n9978), .A2(n6359), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n6358), .ZN(n9981) );
  OAI21_X1 U7995 ( .B1(n6361), .B2(n6360), .A(n7119), .ZN(n6362) );
  NAND2_X1 U7996 ( .A1(n6362), .A2(n9983), .ZN(n6374) );
  INV_X1 U7997 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6363) );
  MUX2_X1 U7998 ( .A(n6363), .B(P1_REG1_REG_10__SCAN_IN), .S(n9832), .Z(n9825)
         );
  NOR2_X1 U7999 ( .A1(n9825), .A2(n9826), .ZN(n9824) );
  INV_X1 U8000 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6366) );
  MUX2_X1 U8001 ( .A(n6366), .B(P1_REG1_REG_11__SCAN_IN), .S(n9978), .Z(n9986)
         );
  NOR2_X1 U8002 ( .A1(n9985), .A2(n9986), .ZN(n9984) );
  AOI21_X1 U8003 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9978), .A(n9984), .ZN(
        n6368) );
  INV_X1 U8004 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10269) );
  AOI22_X1 U8005 ( .A1(n7120), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n10269), .B2(
        n6370), .ZN(n6367) );
  NAND2_X1 U8006 ( .A1(n6368), .A2(n6367), .ZN(n7111) );
  OAI21_X1 U8007 ( .B1(n6368), .B2(n6367), .A(n7111), .ZN(n6372) );
  NAND2_X1 U8008 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7399) );
  NAND2_X1 U8009 ( .A1(n9945), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6369) );
  OAI211_X1 U8010 ( .C1(n9070), .C2(n6370), .A(n7399), .B(n6369), .ZN(n6371)
         );
  AOI21_X1 U8011 ( .B1(n6372), .B2(n9988), .A(n6371), .ZN(n6373) );
  NAND2_X1 U8012 ( .A1(n6374), .A2(n6373), .ZN(P1_U3255) );
  INV_X1 U8013 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6375) );
  INV_X1 U8014 ( .A(n7368), .ZN(n6377) );
  NAND2_X1 U8015 ( .A1(n4594), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6526) );
  XNOR2_X1 U8016 ( .A(n6526), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8148) );
  OAI222_X1 U8017 ( .A1(n8578), .A2(n6375), .B1(n8576), .B2(n6377), .C1(
        P2_U3151), .C2(n8145), .ZN(P2_U3281) );
  INV_X1 U8018 ( .A(n10015), .ZN(n7122) );
  INV_X1 U8019 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6376) );
  OAI222_X1 U8020 ( .A1(n7122), .A2(P1_U3086), .B1(n9820), .B2(n6377), .C1(
        n6376), .C2(n9814), .ZN(P1_U3341) );
  INV_X1 U8021 ( .A(n6438), .ZN(n6387) );
  INV_X1 U8022 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6823) );
  OAI21_X1 U8023 ( .B1(n6378), .B2(n6380), .A(n6379), .ZN(n6381) );
  NAND2_X1 U8024 ( .A1(n6381), .A2(n8680), .ZN(n6386) );
  INV_X1 U8025 ( .A(n10121), .ZN(n6383) );
  OAI22_X1 U8026 ( .A1(n6383), .A2(n8683), .B1(n8689), .B2(n10117), .ZN(n6384)
         );
  AOI21_X1 U8027 ( .B1(n8693), .B2(n9013), .A(n6384), .ZN(n6385) );
  OAI211_X1 U8028 ( .C1(n6387), .C2(n6823), .A(n6386), .B(n6385), .ZN(P1_U3222) );
  INV_X1 U8029 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6939) );
  AOI21_X1 U8030 ( .B1(n6391), .B2(n6939), .A(n6442), .ZN(n6410) );
  INV_X1 U8031 ( .A(n6392), .ZN(n6397) );
  INV_X1 U8032 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6878) );
  MUX2_X1 U8033 ( .A(n6939), .B(n6878), .S(n8255), .Z(n6393) );
  INV_X1 U8034 ( .A(n6919), .ZN(n6403) );
  NAND2_X1 U8035 ( .A1(n6393), .A2(n6403), .ZN(n6445) );
  INV_X1 U8036 ( .A(n6393), .ZN(n6394) );
  NAND2_X1 U8037 ( .A1(n6394), .A2(n6919), .ZN(n6395) );
  NAND2_X1 U8038 ( .A1(n6445), .A2(n6395), .ZN(n6396) );
  AOI21_X1 U8039 ( .B1(n6398), .B2(n6397), .A(n6396), .ZN(n6451) );
  AND3_X1 U8040 ( .A1(n6398), .A2(n6397), .A3(n6396), .ZN(n6399) );
  OAI21_X1 U8041 ( .B1(n6451), .B2(n6399), .A(n10279), .ZN(n6409) );
  NAND2_X1 U8042 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(n6868), .ZN(n6401) );
  NAND2_X1 U8043 ( .A1(n6401), .A2(n6400), .ZN(n6455) );
  XNOR2_X1 U8044 ( .A(n6455), .B(n6403), .ZN(n6402) );
  NAND2_X1 U8045 ( .A1(P2_REG1_REG_7__SCAN_IN), .A2(n6402), .ZN(n6456) );
  OAI21_X1 U8046 ( .B1(n6402), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6456), .ZN(
        n6407) );
  INV_X1 U8047 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6405) );
  NOR2_X1 U8048 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6879), .ZN(n7014) );
  AOI21_X1 U8049 ( .B1(n8202), .B2(n6403), .A(n7014), .ZN(n6404) );
  OAI21_X1 U8050 ( .B1(n6405), .B2(n8204), .A(n6404), .ZN(n6406) );
  AOI21_X1 U8051 ( .B1(n8267), .B2(n6407), .A(n6406), .ZN(n6408) );
  OAI211_X1 U8052 ( .C1(n6410), .C2(n8268), .A(n6409), .B(n6408), .ZN(P2_U3189) );
  INV_X1 U8053 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6414) );
  INV_X1 U8054 ( .A(n7418), .ZN(n6416) );
  NAND2_X1 U8055 ( .A1(n6526), .A2(n6411), .ZN(n6412) );
  NAND2_X1 U8056 ( .A1(n6412), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6413) );
  XNOR2_X1 U8057 ( .A(n6413), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8167) );
  INV_X1 U8058 ( .A(n8167), .ZN(n8173) );
  OAI222_X1 U8059 ( .A1(n8578), .A2(n6414), .B1(n8576), .B2(n6416), .C1(
        P2_U3151), .C2(n8173), .ZN(P2_U3280) );
  INV_X1 U8060 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6415) );
  OAI222_X1 U8061 ( .A1(n7125), .A2(P1_U3086), .B1(n9820), .B2(n6416), .C1(
        n6415), .C2(n9814), .ZN(P1_U3340) );
  NAND2_X1 U8062 ( .A1(n6417), .A2(n7865), .ZN(n6470) );
  NAND2_X1 U8063 ( .A1(n6470), .A2(n7066), .ZN(n6418) );
  NAND2_X1 U8064 ( .A1(n6418), .A2(n8261), .ZN(n6540) );
  OR2_X1 U8065 ( .A1(n6540), .A2(n7865), .ZN(n6419) );
  NAND2_X1 U8066 ( .A1(n6419), .A2(n7850), .ZN(n6555) );
  OR2_X1 U8067 ( .A1(n6555), .A2(n6420), .ZN(n6426) );
  INV_X1 U8068 ( .A(n6467), .ZN(n6421) );
  NAND2_X1 U8069 ( .A1(n6555), .A2(n6421), .ZN(n6425) );
  NAND3_X1 U8070 ( .A1(n6426), .A2(n6425), .A3(n6557), .ZN(n6430) );
  NOR2_X1 U8071 ( .A1(n6534), .A2(n8424), .ZN(n10303) );
  NOR3_X1 U8072 ( .A1(n10300), .A2(n6428), .A3(n10366), .ZN(n6429) );
  AOI211_X1 U8073 ( .C1(n10294), .C2(P2_REG3_REG_0__SCAN_IN), .A(n10303), .B(
        n6429), .ZN(n6431) );
  MUX2_X1 U8074 ( .A(n6432), .B(n6431), .S(n10299), .Z(n6433) );
  OAI21_X1 U8075 ( .B1(n8361), .B2(n6478), .A(n6433), .ZN(P2_U3233) );
  XOR2_X1 U8076 ( .A(n6435), .B(n6434), .Z(n6440) );
  INV_X1 U8077 ( .A(n10089), .ZN(n6719) );
  AOI22_X1 U8078 ( .A1(n8726), .A2(n6717), .B1(n10091), .B2(n8731), .ZN(n6436)
         );
  OAI21_X1 U8079 ( .B1(n6719), .B2(n8729), .A(n6436), .ZN(n6437) );
  AOI21_X1 U8080 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n6438), .A(n6437), .ZN(
        n6439) );
  OAI21_X1 U8081 ( .B1(n6440), .B2(n8733), .A(n6439), .ZN(P1_U3237) );
  INV_X1 U8082 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7060) );
  AOI22_X1 U8083 ( .A1(n7037), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n7060), .B2(
        n6454), .ZN(n6443) );
  NOR2_X1 U8084 ( .A1(n6444), .A2(n6443), .ZN(n6583) );
  AOI21_X1 U8085 ( .B1(n6444), .B2(n6443), .A(n6583), .ZN(n6466) );
  INV_X1 U8086 ( .A(n6445), .ZN(n6450) );
  INV_X1 U8087 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6930) );
  MUX2_X1 U8088 ( .A(n7060), .B(n6930), .S(n8255), .Z(n6446) );
  NAND2_X1 U8089 ( .A1(n6446), .A2(n7037), .ZN(n6589) );
  INV_X1 U8090 ( .A(n6446), .ZN(n6447) );
  NAND2_X1 U8091 ( .A1(n6447), .A2(n6454), .ZN(n6448) );
  AND2_X1 U8092 ( .A1(n6589), .A2(n6448), .ZN(n6449) );
  OAI21_X1 U8093 ( .B1(n6451), .B2(n6450), .A(n6449), .ZN(n6590) );
  INV_X1 U8094 ( .A(n6590), .ZN(n6453) );
  NOR3_X1 U8095 ( .A1(n6451), .A2(n6450), .A3(n6449), .ZN(n6452) );
  OAI21_X1 U8096 ( .B1(n6453), .B2(n6452), .A(n10279), .ZN(n6465) );
  AOI22_X1 U8097 ( .A1(n7037), .A2(n6930), .B1(P2_REG1_REG_8__SCAN_IN), .B2(
        n6454), .ZN(n6459) );
  NAND2_X1 U8098 ( .A1(n6455), .A2(n6919), .ZN(n6457) );
  OAI21_X1 U8099 ( .B1(n6459), .B2(n6458), .A(n6592), .ZN(n6463) );
  INV_X1 U8100 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n9665) );
  NAND2_X1 U8101 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3151), .ZN(n7047) );
  INV_X1 U8102 ( .A(n7047), .ZN(n6460) );
  AOI21_X1 U8103 ( .B1(n8202), .B2(n7037), .A(n6460), .ZN(n6461) );
  OAI21_X1 U8104 ( .B1(n9665), .B2(n8204), .A(n6461), .ZN(n6462) );
  AOI21_X1 U8105 ( .B1(n6463), .B2(n8267), .A(n6462), .ZN(n6464) );
  OAI211_X1 U8106 ( .C1(n6466), .C2(n8268), .A(n6465), .B(n6464), .ZN(P2_U3190) );
  INV_X1 U8107 ( .A(n7865), .ZN(n6531) );
  NAND3_X1 U8108 ( .A1(n6468), .A2(n6531), .A3(n6467), .ZN(n6472) );
  AND2_X1 U8109 ( .A1(n6470), .A2(n6469), .ZN(n6471) );
  OR2_X1 U8110 ( .A1(n6492), .A2(n6473), .ZN(n6475) );
  OR2_X1 U8111 ( .A1(n6494), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6474) );
  OAI211_X1 U8112 ( .C1(n6477), .C2(n6476), .A(n6475), .B(n6474), .ZN(n6547)
         );
  XNOR2_X1 U8113 ( .A(n6486), .B(n6615), .ZN(n6479) );
  OAI22_X1 U8114 ( .A1(n6561), .A2(n6562), .B1(n8116), .B2(n6479), .ZN(n6569)
         );
  OR2_X1 U8115 ( .A1(n6494), .A2(n6480), .ZN(n6485) );
  OR2_X1 U8116 ( .A1(n6492), .A2(n6481), .ZN(n6484) );
  OR2_X1 U8117 ( .A1(n6476), .A2(n6482), .ZN(n6483) );
  INV_X1 U8118 ( .A(n6618), .ZN(n10312) );
  XNOR2_X1 U8119 ( .A(n10312), .B(n6644), .ZN(n6491) );
  NOR2_X1 U8120 ( .A1(n6501), .A2(n10371), .ZN(n6487) );
  NOR2_X1 U8121 ( .A1(n6487), .A2(n5111), .ZN(n6490) );
  INV_X1 U8122 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6619) );
  OR2_X1 U8123 ( .A1(n6499), .A2(n6619), .ZN(n6489) );
  INV_X1 U8124 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6622) );
  OR2_X1 U8125 ( .A1(n6500), .A2(n6622), .ZN(n6488) );
  XNOR2_X1 U8126 ( .A(n6491), .B(n4512), .ZN(n6568) );
  INV_X1 U8127 ( .A(n4512), .ZN(n6520) );
  AOI22_X1 U8128 ( .A1(n6569), .A2(n6568), .B1(n6520), .B2(n6491), .ZN(n6507)
         );
  OR2_X1 U8129 ( .A1(n7035), .A2(n6493), .ZN(n6497) );
  OR2_X1 U8130 ( .A1(n7659), .A2(n6495), .ZN(n6496) );
  OAI211_X1 U8131 ( .C1(n6476), .C2(n6498), .A(n6497), .B(n6496), .ZN(n10293)
         );
  XNOR2_X1 U8132 ( .A(n6644), .B(n10293), .ZN(n6645) );
  NAND2_X1 U8133 ( .A1(n7560), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6505) );
  OR2_X1 U8134 ( .A1(n4494), .A2(n10373), .ZN(n6502) );
  INV_X1 U8135 ( .A(n8115), .ZN(n6665) );
  XNOR2_X1 U8136 ( .A(n6645), .B(n8115), .ZN(n6506) );
  OAI211_X1 U8137 ( .C1(n6507), .C2(n6506), .A(n6648), .B(n8066), .ZN(n6523)
         );
  NAND2_X1 U8138 ( .A1(n7534), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6516) );
  OR2_X1 U8139 ( .A1(n4494), .A2(n6510), .ZN(n6515) );
  NAND2_X1 U8140 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6512) );
  AND2_X1 U8141 ( .A1(n6655), .A2(n6512), .ZN(n6651) );
  OR2_X1 U8142 ( .A1(n7078), .A2(n6651), .ZN(n6514) );
  INV_X1 U8143 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6759) );
  OR2_X1 U8144 ( .A1(n7679), .A2(n6759), .ZN(n6513) );
  NAND2_X1 U8145 ( .A1(n8092), .A2(n10287), .ZN(n6519) );
  AOI21_X1 U8146 ( .B1(n8101), .B2(n10293), .A(n6517), .ZN(n6518) );
  OAI211_X1 U8147 ( .C1(n6520), .C2(n8090), .A(n6519), .B(n6518), .ZN(n6521)
         );
  AOI21_X1 U8148 ( .B1(n10295), .B2(n8081), .A(n6521), .ZN(n6522) );
  NAND2_X1 U8149 ( .A1(n6523), .A2(n6522), .ZN(P2_U3158) );
  INV_X1 U8150 ( .A(n7424), .ZN(n6530) );
  NAND2_X1 U8151 ( .A1(n6524), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6525) );
  NAND2_X1 U8152 ( .A1(n6526), .A2(n6525), .ZN(n6527) );
  NAND2_X1 U8153 ( .A1(n6527), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n6528) );
  INV_X1 U8154 ( .A(n8199), .ZN(n8195) );
  OAI222_X1 U8155 ( .A1(n8578), .A2(n9499), .B1(n8576), .B2(n6530), .C1(
        P2_U3151), .C2(n8195), .ZN(P2_U3279) );
  INV_X1 U8156 ( .A(n9064), .ZN(n7127) );
  OAI222_X1 U8157 ( .A1(n7127), .A2(P1_U3086), .B1(n9820), .B2(n6530), .C1(
        n6529), .C2(n9814), .ZN(P1_U3339) );
  NAND2_X1 U8158 ( .A1(n6417), .A2(n6531), .ZN(n6533) );
  NAND2_X1 U8159 ( .A1(n6535), .A2(n6547), .ZN(n7726) );
  INV_X1 U8160 ( .A(n6614), .ZN(n7694) );
  NAND2_X1 U8161 ( .A1(n6536), .A2(n10304), .ZN(n6613) );
  INV_X1 U8162 ( .A(n6613), .ZN(n6537) );
  XNOR2_X1 U8163 ( .A(n6614), .B(n6537), .ZN(n6546) );
  NAND2_X1 U8164 ( .A1(n6614), .A2(n7721), .ZN(n6539) );
  NAND2_X1 U8165 ( .A1(n6612), .A2(n6539), .ZN(n6604) );
  INV_X1 U8166 ( .A(n6540), .ZN(n6541) );
  INV_X1 U8167 ( .A(n10309), .ZN(n6542) );
  NAND2_X1 U8168 ( .A1(n6604), .A2(n6542), .ZN(n6545) );
  AOI22_X1 U8169 ( .A1(n10286), .A2(n4512), .B1(n6536), .B2(n10285), .ZN(n6544) );
  OAI211_X1 U8170 ( .C1(n10301), .C2(n6546), .A(n6545), .B(n6544), .ZN(n6600)
         );
  INV_X1 U8171 ( .A(n10351), .ZN(n6549) );
  NAND2_X1 U8172 ( .A1(n6604), .A2(n6549), .ZN(n6550) );
  OAI21_X1 U8173 ( .B1(n10356), .B2(n6547), .A(n6550), .ZN(n6551) );
  NOR2_X1 U8174 ( .A1(n6600), .A2(n6551), .ZN(n10306) );
  AND2_X1 U8175 ( .A1(n6552), .A2(n6467), .ZN(n6553) );
  OR2_X1 U8176 ( .A1(n6555), .A2(n6553), .ZN(n6558) );
  NAND2_X1 U8177 ( .A1(n6555), .A2(n6554), .ZN(n6556) );
  MUX2_X1 U8178 ( .A(n6559), .B(n10306), .S(n10386), .Z(n6560) );
  INV_X1 U8179 ( .A(n6560), .ZN(P2_U3460) );
  XOR2_X1 U8180 ( .A(n6561), .B(n6562), .Z(n6567) );
  OAI22_X1 U8181 ( .A1(n8076), .A2(n6547), .B1(n8090), .B2(n6313), .ZN(n6565)
         );
  NOR2_X1 U8182 ( .A1(n6570), .A2(n6563), .ZN(n6564) );
  AOI211_X1 U8183 ( .C1(n8092), .C2(n4512), .A(n6565), .B(n6564), .ZN(n6566)
         );
  OAI21_X1 U8184 ( .B1(n8096), .B2(n6567), .A(n6566), .ZN(P2_U3162) );
  XOR2_X1 U8185 ( .A(n6569), .B(n6568), .Z(n6574) );
  OAI22_X1 U8186 ( .A1(n6618), .A2(n8076), .B1(n8090), .B2(n6534), .ZN(n6572)
         );
  NOR2_X1 U8187 ( .A1(n6570), .A2(n6619), .ZN(n6571) );
  AOI211_X1 U8188 ( .C1(n8092), .C2(n8115), .A(n6572), .B(n6571), .ZN(n6573)
         );
  OAI21_X1 U8189 ( .B1(n8096), .B2(n6574), .A(n6573), .ZN(P2_U3177) );
  XNOR2_X1 U8190 ( .A(n6575), .B(n6576), .ZN(n6577) );
  NAND2_X1 U8191 ( .A1(n6577), .A2(n8680), .ZN(n6581) );
  NAND2_X1 U8192 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9049) );
  INV_X1 U8193 ( .A(n9049), .ZN(n6579) );
  INV_X1 U8194 ( .A(n5287), .ZN(n10150) );
  OAI22_X1 U8195 ( .A1(n8729), .A2(n10150), .B1(n10118), .B2(n8683), .ZN(n6578) );
  AOI211_X1 U8196 ( .C1(n6718), .C2(n8731), .A(n6579), .B(n6578), .ZN(n6580)
         );
  OAI211_X1 U8197 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8696), .A(n6581), .B(
        n6580), .ZN(P1_U3218) );
  NOR2_X1 U8198 ( .A1(n7037), .A2(n7060), .ZN(n6582) );
  INV_X1 U8199 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7092) );
  AOI21_X1 U8200 ( .B1(n6584), .B2(n7092), .A(n6670), .ZN(n6599) );
  INV_X1 U8201 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7041) );
  MUX2_X1 U8202 ( .A(n7092), .B(n7041), .S(n8255), .Z(n6585) );
  NAND2_X1 U8203 ( .A1(n6585), .A2(n7088), .ZN(n6674) );
  INV_X1 U8204 ( .A(n6585), .ZN(n6586) );
  NAND2_X1 U8205 ( .A1(n6586), .A2(n6684), .ZN(n6587) );
  NAND2_X1 U8206 ( .A1(n6674), .A2(n6587), .ZN(n6588) );
  AOI21_X1 U8207 ( .B1(n6590), .B2(n6589), .A(n6588), .ZN(n6680) );
  AND3_X1 U8208 ( .A1(n6590), .A2(n6589), .A3(n6588), .ZN(n6591) );
  OAI21_X1 U8209 ( .B1(n6680), .B2(n6591), .A(n10279), .ZN(n6598) );
  NAND2_X1 U8210 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n6593), .ZN(n6686) );
  OAI21_X1 U8211 ( .B1(n6593), .B2(P2_REG1_REG_9__SCAN_IN), .A(n6686), .ZN(
        n6596) );
  INV_X1 U8212 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n6704) );
  INV_X1 U8213 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7042) );
  NOR2_X1 U8214 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7042), .ZN(n7231) );
  AOI21_X1 U8215 ( .B1(n8202), .B2(n7088), .A(n7231), .ZN(n6594) );
  OAI21_X1 U8216 ( .B1(n6704), .B2(n8204), .A(n6594), .ZN(n6595) );
  AOI21_X1 U8217 ( .B1(n6596), .B2(n8267), .A(n6595), .ZN(n6597) );
  OAI211_X1 U8218 ( .C1(n6599), .C2(n8268), .A(n6598), .B(n6597), .ZN(P2_U3191) );
  INV_X1 U8219 ( .A(n6600), .ZN(n6607) );
  NOR2_X1 U8220 ( .A1(n6470), .A2(n8261), .ZN(n6608) );
  NAND2_X1 U8221 ( .A1(n8433), .A2(n6608), .ZN(n7937) );
  INV_X1 U8222 ( .A(n7937), .ZN(n6605) );
  NOR2_X1 U8223 ( .A1(n8433), .A2(n6601), .ZN(n6603) );
  OAI22_X1 U8224 ( .A1(n8361), .A2(n6547), .B1(n6563), .B2(n8430), .ZN(n6602)
         );
  AOI211_X1 U8225 ( .C1(n6605), .C2(n6604), .A(n6603), .B(n6602), .ZN(n6606)
         );
  OAI21_X1 U8226 ( .B1(n8381), .B2(n6607), .A(n6606), .ZN(P2_U3232) );
  INV_X1 U8227 ( .A(n6608), .ZN(n6609) );
  NAND2_X1 U8228 ( .A1(n10309), .A2(n6609), .ZN(n6610) );
  NAND2_X1 U8229 ( .A1(n4512), .A2(n6618), .ZN(n7729) );
  NAND2_X1 U8230 ( .A1(n6612), .A2(n6611), .ZN(n6747) );
  XNOR2_X1 U8231 ( .A(n6750), .B(n6747), .ZN(n10308) );
  INV_X1 U8232 ( .A(n6750), .ZN(n6746) );
  NAND2_X1 U8233 ( .A1(n6614), .A2(n6613), .ZN(n6616) );
  NAND2_X1 U8234 ( .A1(n6616), .A2(n4522), .ZN(n6751) );
  XNOR2_X1 U8235 ( .A(n6746), .B(n6751), .ZN(n6617) );
  OAI222_X1 U8236 ( .A1(n8424), .A2(n6665), .B1(n8426), .B2(n6534), .C1(n10301), .C2(n6617), .ZN(n10310) );
  OAI22_X1 U8237 ( .A1(n8430), .A2(n6619), .B1(n6618), .B2(n8308), .ZN(n6620)
         );
  NOR2_X1 U8238 ( .A1(n10310), .A2(n6620), .ZN(n6621) );
  MUX2_X1 U8239 ( .A(n6622), .B(n6621), .S(n10299), .Z(n6623) );
  OAI21_X1 U8240 ( .B1(n8420), .B2(n10308), .A(n6623), .ZN(P2_U3231) );
  INV_X1 U8241 ( .A(n7434), .ZN(n6638) );
  NAND2_X1 U8242 ( .A1(n6624), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6625) );
  XNOR2_X1 U8243 ( .A(n6625), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8232) );
  INV_X1 U8244 ( .A(n8232), .ZN(n8217) );
  OAI222_X1 U8245 ( .A1(n8582), .A2(n6638), .B1(n8217), .B2(P2_U3151), .C1(
        n6626), .C2(n8578), .ZN(P2_U3278) );
  INV_X1 U8246 ( .A(n7443), .ZN(n6715) );
  AOI22_X1 U8247 ( .A1(n10042), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n6627), .ZN(n6628) );
  OAI21_X1 U8248 ( .B1(n6715), .B2(n9820), .A(n6628), .ZN(P1_U3337) );
  INV_X1 U8249 ( .A(n10077), .ZN(n6636) );
  AOI21_X1 U8250 ( .B1(n6629), .B2(n6630), .A(n8733), .ZN(n6631) );
  OR2_X1 U8251 ( .A1(n6629), .A2(n6630), .ZN(n6803) );
  NAND2_X1 U8252 ( .A1(n6631), .A2(n6803), .ZN(n6635) );
  AND2_X1 U8253 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9944) );
  INV_X1 U8254 ( .A(n6632), .ZN(n6943) );
  OAI22_X1 U8255 ( .A1(n8729), .A2(n6943), .B1(n6719), .B2(n8683), .ZN(n6633)
         );
  AOI211_X1 U8256 ( .C1(n10078), .C2(n8731), .A(n9944), .B(n6633), .ZN(n6634)
         );
  OAI211_X1 U8257 ( .C1(n8696), .C2(n6636), .A(n6635), .B(n6634), .ZN(P1_U3230) );
  INV_X1 U8258 ( .A(n9080), .ZN(n9069) );
  OAI222_X1 U8259 ( .A1(P1_U3086), .A2(n9069), .B1(n9820), .B2(n6638), .C1(
        n6637), .C2(n9814), .ZN(P1_U3338) );
  OR2_X1 U8260 ( .A1(n7035), .A2(n6639), .ZN(n6643) );
  OR2_X1 U8261 ( .A1(n7659), .A2(n4726), .ZN(n6642) );
  OR2_X1 U8262 ( .A1(n6476), .A2(n6640), .ZN(n6641) );
  XNOR2_X1 U8263 ( .A(n6644), .B(n10321), .ZN(n6788) );
  XNOR2_X1 U8264 ( .A(n6788), .B(n10287), .ZN(n6650) );
  AOI21_X1 U8265 ( .B1(n6650), .B2(n6649), .A(n6789), .ZN(n6668) );
  INV_X1 U8266 ( .A(n6651), .ZN(n6760) );
  NAND2_X1 U8267 ( .A1(n7560), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6661) );
  OR2_X1 U8268 ( .A1(n4494), .A2(n6652), .ZN(n6660) );
  INV_X1 U8269 ( .A(n6655), .ZN(n6654) );
  NAND2_X1 U8270 ( .A1(n6655), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6656) );
  AND2_X1 U8271 ( .A1(n6764), .A2(n6656), .ZN(n6794) );
  OR2_X1 U8272 ( .A1(n7078), .A2(n6794), .ZN(n6659) );
  OR2_X1 U8273 ( .A1(n7679), .A2(n6657), .ZN(n6658) );
  NAND2_X1 U8274 ( .A1(n8092), .A2(n8114), .ZN(n6664) );
  INV_X1 U8275 ( .A(n10321), .ZN(n6771) );
  AOI21_X1 U8276 ( .B1(n8101), .B2(n6771), .A(n6662), .ZN(n6663) );
  OAI211_X1 U8277 ( .C1(n6665), .C2(n8090), .A(n6664), .B(n6663), .ZN(n6666)
         );
  AOI21_X1 U8278 ( .B1(n6760), .B2(n8081), .A(n6666), .ZN(n6667) );
  OAI21_X1 U8279 ( .B1(n6668), .B2(n8096), .A(n6667), .ZN(P2_U3170) );
  INV_X1 U8280 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6671) );
  AOI22_X1 U8281 ( .A1(n7147), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n6671), .B2(
        n6683), .ZN(n6672) );
  NOR2_X1 U8282 ( .A1(n6673), .A2(n6672), .ZN(n6845) );
  AOI21_X1 U8283 ( .B1(n6673), .B2(n6672), .A(n6845), .ZN(n6696) );
  INV_X1 U8284 ( .A(n6674), .ZN(n6679) );
  INV_X1 U8285 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7073) );
  MUX2_X1 U8286 ( .A(n6671), .B(n7073), .S(n8255), .Z(n6675) );
  NAND2_X1 U8287 ( .A1(n6675), .A2(n7147), .ZN(n6856) );
  INV_X1 U8288 ( .A(n6675), .ZN(n6676) );
  NAND2_X1 U8289 ( .A1(n6676), .A2(n6683), .ZN(n6677) );
  AND2_X1 U8290 ( .A1(n6856), .A2(n6677), .ZN(n6678) );
  OAI21_X1 U8291 ( .B1(n6680), .B2(n6679), .A(n6678), .ZN(n6857) );
  INV_X1 U8292 ( .A(n6857), .ZN(n6682) );
  NOR3_X1 U8293 ( .A1(n6680), .A2(n6679), .A3(n6678), .ZN(n6681) );
  OAI21_X1 U8294 ( .B1(n6682), .B2(n6681), .A(n10279), .ZN(n6695) );
  AOI22_X1 U8295 ( .A1(n7147), .A2(n7073), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n6683), .ZN(n6689) );
  NAND2_X1 U8296 ( .A1(n6685), .A2(n6684), .ZN(n6687) );
  OAI21_X1 U8297 ( .B1(n6689), .B2(n6688), .A(n6848), .ZN(n6693) );
  INV_X1 U8298 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n6703) );
  INV_X1 U8299 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6690) );
  NOR2_X1 U8300 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6690), .ZN(n7300) );
  AOI21_X1 U8301 ( .B1(n8202), .B2(n7147), .A(n7300), .ZN(n6691) );
  OAI21_X1 U8302 ( .B1(n6703), .B2(n8204), .A(n6691), .ZN(n6692) );
  AOI21_X1 U8303 ( .B1(n6693), .B2(n8267), .A(n6692), .ZN(n6694) );
  OAI211_X1 U8304 ( .C1(n6696), .C2(n8268), .A(n6695), .B(n6694), .ZN(P2_U3192) );
  INV_X1 U8305 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10399) );
  INV_X1 U8306 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10047) );
  NOR2_X1 U8307 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n6697) );
  AOI21_X1 U8308 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n6697), .ZN(n10402) );
  NOR2_X1 U8309 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n6698) );
  AOI21_X1 U8310 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n6698), .ZN(n10405) );
  NOR2_X1 U8311 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n6699) );
  AOI21_X1 U8312 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n6699), .ZN(n10408) );
  INV_X1 U8313 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10019) );
  INV_X1 U8314 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n9357) );
  AOI22_X1 U8315 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .B1(n10019), .B2(n9357), .ZN(n10411) );
  NOR2_X1 U8316 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n6700) );
  AOI21_X1 U8317 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n6700), .ZN(n10414) );
  NOR2_X1 U8318 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n6701) );
  AOI21_X1 U8319 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n6701), .ZN(n10417) );
  NOR2_X1 U8320 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n6702) );
  AOI21_X1 U8321 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n6702), .ZN(n10420) );
  INV_X1 U8322 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9836) );
  AOI22_X1 U8323 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .B1(n6703), .B2(n9836), .ZN(n10423) );
  INV_X1 U8324 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9640) );
  AOI22_X1 U8325 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(P2_ADDR_REG_9__SCAN_IN), 
        .B1(n6704), .B2(n9640), .ZN(n10438) );
  INV_X1 U8326 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9867) );
  AOI22_X1 U8327 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(P2_ADDR_REG_8__SCAN_IN), 
        .B1(n9665), .B2(n9867), .ZN(n10429) );
  NOR2_X1 U8328 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n6705) );
  AOI21_X1 U8329 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n6705), .ZN(n10435) );
  NOR2_X1 U8330 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n6706) );
  AOI21_X1 U8331 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n6706), .ZN(n10426) );
  NOR2_X1 U8332 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n6707) );
  AOI21_X1 U8333 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n6707), .ZN(n10432) );
  INV_X1 U8334 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10394) );
  INV_X1 U8335 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10393) );
  NOR2_X1 U8336 ( .A1(n10394), .A2(n10393), .ZN(n10392) );
  NOR2_X1 U8337 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10392), .ZN(n10388) );
  INV_X1 U8338 ( .A(n10388), .ZN(n10389) );
  INV_X1 U8339 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10391) );
  NAND3_X1 U8340 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_1__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10390) );
  NAND2_X1 U8341 ( .A1(n10391), .A2(n10390), .ZN(n10387) );
  NAND2_X1 U8342 ( .A1(n10389), .A2(n10387), .ZN(n10441) );
  NAND2_X1 U8343 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n6708) );
  OAI21_X1 U8344 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n6708), .ZN(n10440) );
  NOR2_X1 U8345 ( .A1(n10441), .A2(n10440), .ZN(n10439) );
  AOI21_X1 U8346 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10439), .ZN(n10444) );
  NAND2_X1 U8347 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n6709) );
  OAI21_X1 U8348 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n6709), .ZN(n10443) );
  NOR2_X1 U8349 ( .A1(n10444), .A2(n10443), .ZN(n10442) );
  AOI21_X1 U8350 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10442), .ZN(n10447) );
  INV_X1 U8351 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9676) );
  AOI22_X1 U8352 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .B1(n9676), .B2(n6211), .ZN(n10446) );
  NAND2_X1 U8353 ( .A1(n10447), .A2(n10446), .ZN(n10445) );
  OAI21_X1 U8354 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n10445), .ZN(n10431) );
  NAND2_X1 U8355 ( .A1(n10432), .A2(n10431), .ZN(n10430) );
  OAI21_X1 U8356 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10430), .ZN(n10425) );
  NAND2_X1 U8357 ( .A1(n10426), .A2(n10425), .ZN(n10424) );
  OAI21_X1 U8358 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10424), .ZN(n10434) );
  NAND2_X1 U8359 ( .A1(n10435), .A2(n10434), .ZN(n10433) );
  OAI21_X1 U8360 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10433), .ZN(n10428) );
  NAND2_X1 U8361 ( .A1(n10429), .A2(n10428), .ZN(n10427) );
  OAI21_X1 U8362 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n10427), .ZN(n10437) );
  NAND2_X1 U8363 ( .A1(n10438), .A2(n10437), .ZN(n10436) );
  OAI21_X1 U8364 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n10436), .ZN(n10422) );
  NAND2_X1 U8365 ( .A1(n10423), .A2(n10422), .ZN(n10421) );
  OAI21_X1 U8366 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10421), .ZN(n10419) );
  NAND2_X1 U8367 ( .A1(n10420), .A2(n10419), .ZN(n10418) );
  OAI21_X1 U8368 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10418), .ZN(n10416) );
  NAND2_X1 U8369 ( .A1(n10417), .A2(n10416), .ZN(n10415) );
  OAI21_X1 U8370 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10415), .ZN(n10413) );
  NAND2_X1 U8371 ( .A1(n10414), .A2(n10413), .ZN(n10412) );
  OAI21_X1 U8372 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10412), .ZN(n10410) );
  NAND2_X1 U8373 ( .A1(n10411), .A2(n10410), .ZN(n10409) );
  OAI21_X1 U8374 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10409), .ZN(n10407) );
  NAND2_X1 U8375 ( .A1(n10408), .A2(n10407), .ZN(n10406) );
  OAI21_X1 U8376 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10406), .ZN(n10404) );
  NAND2_X1 U8377 ( .A1(n10405), .A2(n10404), .ZN(n10403) );
  OAI21_X1 U8378 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10403), .ZN(n10401) );
  NAND2_X1 U8379 ( .A1(n10402), .A2(n10401), .ZN(n10400) );
  OAI21_X1 U8380 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10400), .ZN(n6710) );
  OR2_X1 U8381 ( .A1(n10047), .A2(n6710), .ZN(n10398) );
  NAND2_X1 U8382 ( .A1(n10399), .A2(n10398), .ZN(n10395) );
  NAND2_X1 U8383 ( .A1(n10047), .A2(n6710), .ZN(n10397) );
  NAND2_X1 U8384 ( .A1(n10395), .A2(n10397), .ZN(n6712) );
  XNOR2_X1 U8385 ( .A(n5168), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n6711) );
  XNOR2_X1 U8386 ( .A(n6712), .B(n6711), .ZN(ADD_1068_U4) );
  NAND2_X1 U8387 ( .A1(n6713), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6714) );
  XNOR2_X1 U8388 ( .A(n6714), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8253) );
  INV_X1 U8389 ( .A(n8253), .ZN(n8249) );
  OAI222_X1 U8390 ( .A1(n8578), .A2(n6716), .B1(n8249), .B2(P2_U3151), .C1(
        n8582), .C2(n6715), .ZN(P2_U3277) );
  NAND2_X1 U8391 ( .A1(n10121), .A2(n6827), .ZN(n6819) );
  NAND2_X1 U8392 ( .A1(n10118), .A2(n10091), .ZN(n8755) );
  NAND2_X1 U8393 ( .A1(n9013), .A2(n10095), .ZN(n8943) );
  OAI22_X1 U8394 ( .A1(n10093), .A2(n10094), .B1(n10091), .B2(n9013), .ZN(
        n6739) );
  NAND2_X1 U8395 ( .A1(n6719), .A2(n6718), .ZN(n8753) );
  NAND2_X1 U8396 ( .A1(n10089), .A2(n10138), .ZN(n8762) );
  NAND2_X1 U8397 ( .A1(n8753), .A2(n8762), .ZN(n6735) );
  AOI22_X1 U8398 ( .A1(n6739), .A2(n6735), .B1(n6719), .B2(n10138), .ZN(n10080) );
  NAND2_X1 U8399 ( .A1(n10150), .A2(n10078), .ZN(n8761) );
  INV_X1 U8400 ( .A(n10078), .ZN(n10143) );
  OAI22_X1 U8401 ( .A1(n10080), .A2(n10079), .B1(n10078), .B2(n5287), .ZN(
        n6945) );
  NAND2_X1 U8402 ( .A1(n6943), .A2(n10153), .ZN(n8775) );
  INV_X1 U8403 ( .A(n10153), .ZN(n6944) );
  NAND2_X1 U8404 ( .A1(n6632), .A2(n6944), .ZN(n8772) );
  NAND2_X1 U8405 ( .A1(n8775), .A2(n8772), .ZN(n8874) );
  INV_X1 U8406 ( .A(n8874), .ZN(n6946) );
  XNOR2_X1 U8407 ( .A(n6945), .B(n6946), .ZN(n10155) );
  NAND3_X1 U8408 ( .A1(n6722), .A2(n6721), .A3(n6720), .ZN(n6723) );
  NAND2_X1 U8409 ( .A1(n6724), .A2(n8995), .ZN(n6725) );
  AND2_X1 U8410 ( .A1(n10116), .A2(n6725), .ZN(n6726) );
  AOI211_X1 U8411 ( .C1(n10153), .C2(n10082), .A(n9339), .B(n10071), .ZN(
        n10151) );
  INV_X2 U8412 ( .A(n9306), .ZN(n10092) );
  AOI22_X1 U8413 ( .A1(n4495), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n6813), .B2(
        n10092), .ZN(n6728) );
  OAI21_X1 U8414 ( .B1(n9341), .B2(n6944), .A(n6728), .ZN(n6730) );
  OR2_X1 U8415 ( .A1(n4495), .A2(n10236), .ZN(n9192) );
  OAI22_X1 U8416 ( .A1(n10149), .A2(n9192), .B1(n9348), .B2(n10150), .ZN(n6729) );
  AOI211_X1 U8417 ( .C1(n10151), .C2(n10101), .A(n6730), .B(n6729), .ZN(n6738)
         );
  NAND2_X1 U8418 ( .A1(n6821), .A2(n6820), .ZN(n6733) );
  NAND2_X1 U8419 ( .A1(n6731), .A2(n6382), .ZN(n6732) );
  NAND2_X1 U8420 ( .A1(n6733), .A2(n6732), .ZN(n10087) );
  NAND2_X1 U8421 ( .A1(n10087), .A2(n8943), .ZN(n6734) );
  NAND2_X1 U8422 ( .A1(n6734), .A2(n8755), .ZN(n8754) );
  NAND2_X1 U8423 ( .A1(n6740), .A2(n8753), .ZN(n10075) );
  NAND2_X1 U8424 ( .A1(n10075), .A2(n8944), .ZN(n6736) );
  NAND2_X1 U8425 ( .A1(n6736), .A2(n8761), .ZN(n6947) );
  XNOR2_X1 U8426 ( .A(n6947), .B(n6946), .ZN(n10157) );
  NAND2_X1 U8427 ( .A1(n10157), .A2(n9301), .ZN(n6737) );
  OAI211_X1 U8428 ( .C1(n10155), .C2(n9322), .A(n6738), .B(n6737), .ZN(
        P1_U3288) );
  XNOR2_X1 U8429 ( .A(n6739), .B(n8873), .ZN(n10134) );
  OAI21_X1 U8430 ( .B1(n8873), .B2(n8754), .A(n6740), .ZN(n6741) );
  AOI222_X1 U8431 ( .A1(n10203), .A2(n6741), .B1(n5287), .B2(n10191), .C1(
        n9013), .C2(n10194), .ZN(n10137) );
  MUX2_X1 U8432 ( .A(n6089), .B(n10137), .S(n9309), .Z(n6745) );
  OR2_X1 U8433 ( .A1(n10096), .A2(n10138), .ZN(n6742) );
  AND3_X1 U8434 ( .A1(n6742), .A2(n10081), .A3(n10097), .ZN(n10135) );
  OAI22_X1 U8435 ( .A1(n9341), .A2(n10138), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9306), .ZN(n6743) );
  AOI21_X1 U8436 ( .B1(n10101), .B2(n10135), .A(n6743), .ZN(n6744) );
  OAI211_X1 U8437 ( .C1(n10134), .C2(n9322), .A(n6745), .B(n6744), .ZN(
        P1_U3290) );
  OR2_X1 U8438 ( .A1(n10287), .A2(n10321), .ZN(n7736) );
  NAND2_X1 U8439 ( .A1(n10287), .A2(n10321), .ZN(n7745) );
  NAND2_X1 U8440 ( .A1(n7736), .A2(n7745), .ZN(n6781) );
  NAND2_X1 U8441 ( .A1(n6747), .A2(n6746), .ZN(n6748) );
  NAND2_X1 U8442 ( .A1(n6748), .A2(n7724), .ZN(n10291) );
  XNOR2_X1 U8443 ( .A(n8115), .B(n10293), .ZN(n10290) );
  NAND2_X1 U8444 ( .A1(n10291), .A2(n10290), .ZN(n6749) );
  INV_X1 U8445 ( .A(n10293), .ZN(n10315) );
  OR2_X1 U8446 ( .A1(n8115), .A2(n10315), .ZN(n7743) );
  NAND2_X1 U8447 ( .A1(n6751), .A2(n6750), .ZN(n6753) );
  OR2_X1 U8448 ( .A1(n4512), .A2(n10312), .ZN(n6752) );
  NAND2_X1 U8449 ( .A1(n6753), .A2(n6752), .ZN(n10284) );
  NOR2_X1 U8450 ( .A1(n8115), .A2(n10293), .ZN(n6755) );
  NAND2_X1 U8451 ( .A1(n8115), .A2(n10293), .ZN(n6754) );
  OAI21_X1 U8452 ( .B1(n10284), .B2(n6755), .A(n6754), .ZN(n6756) );
  INV_X1 U8453 ( .A(n6756), .ZN(n6757) );
  NAND2_X1 U8454 ( .A1(n6757), .A2(n6781), .ZN(n6773) );
  OAI21_X1 U8455 ( .B1(n6757), .B2(n6781), .A(n6773), .ZN(n6758) );
  AOI222_X1 U8456 ( .A1(n10289), .A2(n6758), .B1(n8115), .B2(n10285), .C1(
        n8114), .C2(n10286), .ZN(n10320) );
  MUX2_X1 U8457 ( .A(n6759), .B(n10320), .S(n10299), .Z(n6762) );
  AOI22_X1 U8458 ( .A1(n10292), .A2(n6771), .B1(n10294), .B2(n6760), .ZN(n6761) );
  OAI211_X1 U8459 ( .C1(n8420), .C2(n10319), .A(n6762), .B(n6761), .ZN(
        P2_U3229) );
  NAND2_X1 U8460 ( .A1(n7559), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6770) );
  INV_X1 U8461 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6763) );
  OR2_X1 U8462 ( .A1(n7526), .A2(n6763), .ZN(n6769) );
  NAND2_X1 U8463 ( .A1(n6764), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6765) );
  AND2_X1 U8464 ( .A1(n6880), .A2(n6765), .ZN(n6912) );
  OR2_X1 U8465 ( .A1(n7078), .A2(n6912), .ZN(n6768) );
  OR2_X1 U8466 ( .A1(n4494), .A2(n10377), .ZN(n6767) );
  NAND4_X1 U8467 ( .A1(n6770), .A2(n6769), .A3(n6768), .A4(n6767), .ZN(n8113)
         );
  INV_X1 U8468 ( .A(n8113), .ZN(n6780) );
  INV_X1 U8469 ( .A(n10287), .ZN(n6793) );
  OR2_X1 U8470 ( .A1(n10287), .A2(n6771), .ZN(n6772) );
  OR2_X1 U8471 ( .A1(n7035), .A2(n6774), .ZN(n6777) );
  OR2_X1 U8472 ( .A1(n7659), .A2(n6775), .ZN(n6776) );
  OAI211_X1 U8473 ( .C1(n6476), .C2(n6778), .A(n6777), .B(n6776), .ZN(n6872)
         );
  INV_X1 U8474 ( .A(n6872), .ZN(n10325) );
  NAND2_X1 U8475 ( .A1(n8114), .A2(n10325), .ZN(n7744) );
  XNOR2_X1 U8476 ( .A(n6875), .B(n7696), .ZN(n6779) );
  OAI222_X1 U8477 ( .A1(n8424), .A2(n6780), .B1(n8426), .B2(n6793), .C1(n10301), .C2(n6779), .ZN(n10326) );
  INV_X1 U8478 ( .A(n10326), .ZN(n6787) );
  INV_X1 U8479 ( .A(n6781), .ZN(n7733) );
  NAND2_X1 U8480 ( .A1(n6782), .A2(n7736), .ZN(n6783) );
  OAI21_X1 U8481 ( .B1(n6783), .B2(n7696), .A(n6865), .ZN(n10328) );
  NOR2_X1 U8482 ( .A1(n10299), .A2(n6657), .ZN(n6785) );
  OAI22_X1 U8483 ( .A1(n8361), .A2(n10325), .B1(n6794), .B2(n8430), .ZN(n6784)
         );
  AOI211_X1 U8484 ( .C1(n10328), .C2(n10296), .A(n6785), .B(n6784), .ZN(n6786)
         );
  OAI21_X1 U8485 ( .B1(n6787), .B2(n8381), .A(n6786), .ZN(P2_U3228) );
  XNOR2_X1 U8486 ( .A(n7900), .B(n10325), .ZN(n6905) );
  XNOR2_X1 U8487 ( .A(n6905), .B(n8114), .ZN(n6906) );
  INV_X1 U8488 ( .A(n6788), .ZN(n6790) );
  XOR2_X1 U8489 ( .A(n6906), .B(n6907), .Z(n6798) );
  AOI21_X1 U8490 ( .B1(n8101), .B2(n6872), .A(n6791), .ZN(n6792) );
  OAI21_X1 U8491 ( .B1(n8090), .B2(n6793), .A(n6792), .ZN(n6796) );
  NOR2_X1 U8492 ( .A1(n8094), .A2(n6794), .ZN(n6795) );
  AOI211_X1 U8493 ( .C1(n8092), .C2(n8113), .A(n6796), .B(n6795), .ZN(n6797)
         );
  OAI21_X1 U8494 ( .B1(n6798), .B2(n8096), .A(n6797), .ZN(P2_U3167) );
  INV_X1 U8495 ( .A(n6799), .ZN(n6801) );
  NAND2_X1 U8496 ( .A1(n6801), .A2(n6800), .ZN(n6807) );
  NAND2_X1 U8497 ( .A1(n6803), .A2(n5318), .ZN(n6805) );
  OR2_X1 U8498 ( .A1(n6805), .A2(n6804), .ZN(n6806) );
  AOI22_X1 U8499 ( .A1(n6808), .A2(n6807), .B1(n6802), .B2(n6806), .ZN(n6815)
         );
  AOI22_X1 U8500 ( .A1(n8726), .A2(n5287), .B1(n8693), .B2(n10166), .ZN(n6811)
         );
  NAND2_X1 U8501 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9961) );
  INV_X1 U8502 ( .A(n9961), .ZN(n6809) );
  AOI21_X1 U8503 ( .B1(n8731), .B2(n10153), .A(n6809), .ZN(n6810) );
  NAND2_X1 U8504 ( .A1(n6811), .A2(n6810), .ZN(n6812) );
  AOI21_X1 U8505 ( .B1(n6813), .B2(n8725), .A(n6812), .ZN(n6814) );
  OAI21_X1 U8506 ( .B1(n6815), .B2(n8733), .A(n6814), .ZN(P1_U3227) );
  INV_X1 U8507 ( .A(n7453), .ZN(n6818) );
  OAI222_X1 U8508 ( .A1(n8578), .A2(n6816), .B1(n8576), .B2(n6818), .C1(n8261), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  OAI222_X1 U8509 ( .A1(n9086), .A2(P1_U3086), .B1(n9820), .B2(n6818), .C1(
        n6817), .C2(n9814), .ZN(P1_U3336) );
  XNOR2_X1 U8510 ( .A(n6821), .B(n6819), .ZN(n10124) );
  XNOR2_X1 U8511 ( .A(n6821), .B(n6820), .ZN(n6822) );
  NAND2_X1 U8512 ( .A1(n6822), .A2(n10203), .ZN(n10122) );
  INV_X1 U8513 ( .A(n10122), .ZN(n6832) );
  OAI22_X1 U8514 ( .A1(n9309), .A2(n6824), .B1(n6823), .B2(n9306), .ZN(n6825)
         );
  AOI21_X1 U8515 ( .B1(n10090), .B2(n6382), .A(n6825), .ZN(n6830) );
  INV_X1 U8516 ( .A(n6826), .ZN(n10099) );
  AOI211_X1 U8517 ( .C1(n6827), .C2(n6382), .A(n9339), .B(n10099), .ZN(n10119)
         );
  INV_X1 U8518 ( .A(n9348), .ZN(n6828) );
  AOI22_X1 U8519 ( .A1(n10119), .A2(n10101), .B1(n6828), .B2(n10121), .ZN(
        n6829) );
  OAI211_X1 U8520 ( .C1(n10118), .C2(n9192), .A(n6830), .B(n6829), .ZN(n6831)
         );
  AOI21_X1 U8521 ( .B1(n6832), .B2(n9309), .A(n6831), .ZN(n6833) );
  OAI21_X1 U8522 ( .B1(n9322), .B2(n10124), .A(n6833), .ZN(P1_U3292) );
  INV_X1 U8523 ( .A(n10066), .ZN(n6843) );
  OAI21_X1 U8524 ( .B1(n6836), .B2(n6802), .A(n6835), .ZN(n6837) );
  NAND2_X1 U8525 ( .A1(n6837), .A2(n8680), .ZN(n6842) );
  INV_X1 U8526 ( .A(n10065), .ZN(n6963) );
  NAND2_X1 U8527 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9975) );
  INV_X1 U8528 ( .A(n9975), .ZN(n6838) );
  AOI21_X1 U8529 ( .B1(n8726), .B2(n6632), .A(n6838), .ZN(n6839) );
  OAI21_X1 U8530 ( .B1(n6963), .B2(n8729), .A(n6839), .ZN(n6840) );
  AOI21_X1 U8531 ( .B1(n10067), .B2(n8731), .A(n6840), .ZN(n6841) );
  OAI211_X1 U8532 ( .C1(n8696), .C2(n6843), .A(n6842), .B(n6841), .ZN(P1_U3239) );
  NOR2_X1 U8533 ( .A1(n7147), .A2(n6671), .ZN(n6844) );
  NAND2_X1 U8534 ( .A1(n6846), .A2(n6994), .ZN(n6980) );
  INV_X1 U8535 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7610) );
  AOI21_X1 U8536 ( .B1(n6847), .B2(n7610), .A(n6982), .ZN(n6864) );
  NAND2_X1 U8537 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n6849), .ZN(n6996) );
  OAI21_X1 U8538 ( .B1(n6849), .B2(P2_REG1_REG_11__SCAN_IN), .A(n6996), .ZN(
        n6862) );
  INV_X1 U8539 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n6851) );
  AND2_X1 U8540 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8054) );
  AOI21_X1 U8541 ( .B1(n8202), .B2(n7266), .A(n8054), .ZN(n6850) );
  OAI21_X1 U8542 ( .B1(n6851), .B2(n8204), .A(n6850), .ZN(n6861) );
  INV_X1 U8543 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7155) );
  MUX2_X1 U8544 ( .A(n7610), .B(n7155), .S(n8255), .Z(n6852) );
  NAND2_X1 U8545 ( .A1(n6852), .A2(n7266), .ZN(n6985) );
  INV_X1 U8546 ( .A(n6852), .ZN(n6853) );
  NAND2_X1 U8547 ( .A1(n6853), .A2(n6994), .ZN(n6854) );
  NAND2_X1 U8548 ( .A1(n6985), .A2(n6854), .ZN(n6855) );
  AOI21_X1 U8549 ( .B1(n6857), .B2(n6856), .A(n6855), .ZN(n6991) );
  INV_X1 U8550 ( .A(n6991), .ZN(n6859) );
  NAND3_X1 U8551 ( .A1(n6857), .A2(n6856), .A3(n6855), .ZN(n6858) );
  AOI21_X1 U8552 ( .B1(n6859), .B2(n6858), .A(n8264), .ZN(n6860) );
  AOI211_X1 U8553 ( .C1(n8267), .C2(n6862), .A(n6861), .B(n6860), .ZN(n6863)
         );
  OAI21_X1 U8554 ( .B1(n6864), .B2(n8268), .A(n6863), .ZN(P2_U3193) );
  OR2_X1 U8555 ( .A1(n7035), .A2(n6866), .ZN(n6871) );
  OR2_X1 U8556 ( .A1(n7659), .A2(n6867), .ZN(n6870) );
  OR2_X1 U8557 ( .A1(n6476), .A2(n6868), .ZN(n6869) );
  NAND2_X1 U8558 ( .A1(n8113), .A2(n10330), .ZN(n7751) );
  NAND2_X1 U8559 ( .A1(n7749), .A2(n7751), .ZN(n6876) );
  INV_X1 U8560 ( .A(n6876), .ZN(n7695) );
  XNOR2_X1 U8561 ( .A(n6916), .B(n7695), .ZN(n10333) );
  INV_X1 U8562 ( .A(n10333), .ZN(n6891) );
  NAND2_X1 U8563 ( .A1(n8114), .A2(n6872), .ZN(n6874) );
  NOR2_X1 U8564 ( .A1(n8114), .A2(n6872), .ZN(n6873) );
  NAND2_X1 U8565 ( .A1(n6877), .A2(n6876), .ZN(n6927) );
  OAI211_X1 U8566 ( .C1(n6877), .C2(n6876), .A(n6927), .B(n10289), .ZN(n6887)
         );
  NAND2_X1 U8567 ( .A1(n7560), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6885) );
  OR2_X1 U8568 ( .A1(n4494), .A2(n6878), .ZN(n6884) );
  NAND2_X1 U8569 ( .A1(n6880), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6881) );
  AND2_X1 U8570 ( .A1(n6931), .A2(n6881), .ZN(n7013) );
  OR2_X1 U8571 ( .A1(n7078), .A2(n7013), .ZN(n6883) );
  OR2_X1 U8572 ( .A1(n7679), .A2(n6939), .ZN(n6882) );
  NAND4_X1 U8573 ( .A1(n6885), .A2(n6884), .A3(n6883), .A4(n6882), .ZN(n8112)
         );
  AOI22_X1 U8574 ( .A1(n10285), .A2(n8114), .B1(n8112), .B2(n10286), .ZN(n6886) );
  NAND2_X1 U8575 ( .A1(n6887), .A2(n6886), .ZN(n10331) );
  NOR2_X1 U8576 ( .A1(n8433), .A2(n6340), .ZN(n6889) );
  OAI22_X1 U8577 ( .A1(n8361), .A2(n10330), .B1(n6912), .B2(n8430), .ZN(n6888)
         );
  AOI211_X1 U8578 ( .C1(n10331), .C2(n10299), .A(n6889), .B(n6888), .ZN(n6890)
         );
  OAI21_X1 U8579 ( .B1(n8420), .B2(n6891), .A(n6890), .ZN(P2_U3227) );
  XNOR2_X1 U8580 ( .A(n6894), .B(n6893), .ZN(n6895) );
  XNOR2_X1 U8581 ( .A(n6892), .B(n6895), .ZN(n6901) );
  NAND2_X1 U8582 ( .A1(n8725), .A2(n6953), .ZN(n6898) );
  NAND2_X1 U8583 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9849) );
  INV_X1 U8584 ( .A(n9849), .ZN(n6896) );
  AOI21_X1 U8585 ( .B1(n8726), .B2(n10166), .A(n6896), .ZN(n6897) );
  OAI211_X1 U8586 ( .C1(n7022), .C2(n8729), .A(n6898), .B(n6897), .ZN(n6899)
         );
  AOI21_X1 U8587 ( .B1(n6951), .B2(n8731), .A(n6899), .ZN(n6900) );
  OAI21_X1 U8588 ( .B1(n6901), .B2(n8733), .A(n6900), .ZN(P1_U3213) );
  INV_X1 U8589 ( .A(n7465), .ZN(n6903) );
  OAI222_X1 U8590 ( .A1(n8582), .A2(n6903), .B1(P2_U3151), .B2(n7865), .C1(
        n9367), .C2(n8578), .ZN(P2_U3275) );
  OAI222_X1 U8591 ( .A1(P1_U3086), .A2(n6904), .B1(n9820), .B2(n6903), .C1(
        n6902), .C2(n9814), .ZN(P1_U3335) );
  XNOR2_X1 U8592 ( .A(n7900), .B(n10330), .ZN(n7007) );
  XNOR2_X1 U8593 ( .A(n7007), .B(n8113), .ZN(n6909) );
  AOI211_X1 U8594 ( .C1(n6909), .C2(n6908), .A(n8096), .B(n7009), .ZN(n6915)
         );
  OAI22_X1 U8595 ( .A1(n8084), .A2(n5040), .B1(n10330), .B2(n8076), .ZN(n6914)
         );
  NAND2_X1 U8596 ( .A1(n8080), .A2(n8114), .ZN(n6910) );
  OAI211_X1 U8597 ( .C1(n8094), .C2(n6912), .A(n6911), .B(n6910), .ZN(n6913)
         );
  OR3_X1 U8598 ( .A1(n6915), .A2(n6914), .A3(n6913), .ZN(P2_U3179) );
  OR2_X1 U8599 ( .A1(n7035), .A2(n6917), .ZN(n6922) );
  OR2_X1 U8600 ( .A1(n7659), .A2(n6918), .ZN(n6921) );
  OR2_X1 U8601 ( .A1(n6476), .A2(n6919), .ZN(n6920) );
  OR2_X1 U8602 ( .A1(n8112), .A2(n10334), .ZN(n7759) );
  NAND2_X1 U8603 ( .A1(n8112), .A2(n10334), .ZN(n7094) );
  NAND2_X1 U8604 ( .A1(n6923), .A2(n4515), .ZN(n6924) );
  NAND2_X1 U8605 ( .A1(n7095), .A2(n6924), .ZN(n10335) );
  INV_X1 U8606 ( .A(n10330), .ZN(n6925) );
  NAND2_X1 U8607 ( .A1(n8113), .A2(n6925), .ZN(n6926) );
  OAI21_X1 U8608 ( .B1(n6928), .B2(n4515), .A(n7056), .ZN(n6929) );
  NAND2_X1 U8609 ( .A1(n6929), .A2(n10289), .ZN(n6938) );
  NAND2_X1 U8610 ( .A1(n7560), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6936) );
  OR2_X1 U8611 ( .A1(n4494), .A2(n6930), .ZN(n6935) );
  NAND2_X1 U8612 ( .A1(n6931), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6932) );
  AND2_X1 U8613 ( .A1(n7076), .A2(n6932), .ZN(n7059) );
  OR2_X1 U8614 ( .A1(n7078), .A2(n7059), .ZN(n6934) );
  OR2_X1 U8615 ( .A1(n7679), .A2(n7060), .ZN(n6933) );
  NAND4_X1 U8616 ( .A1(n6936), .A2(n6935), .A3(n6934), .A4(n6933), .ZN(n8111)
         );
  AOI22_X1 U8617 ( .A1(n10285), .A2(n8113), .B1(n8111), .B2(n10286), .ZN(n6937) );
  OAI211_X1 U8618 ( .C1(n10335), .C2(n10309), .A(n6938), .B(n6937), .ZN(n10337) );
  NAND2_X1 U8619 ( .A1(n10337), .A2(n8433), .ZN(n6942) );
  INV_X1 U8620 ( .A(n10334), .ZN(n7054) );
  OAI22_X1 U8621 ( .A1(n8433), .A2(n6939), .B1(n7013), .B2(n8430), .ZN(n6940)
         );
  AOI21_X1 U8622 ( .B1(n10292), .B2(n7054), .A(n6940), .ZN(n6941) );
  OAI211_X1 U8623 ( .C1(n10335), .C2(n7937), .A(n6942), .B(n6941), .ZN(
        P2_U3226) );
  INV_X1 U8624 ( .A(n7476), .ZN(n6962) );
  OAI222_X1 U8625 ( .A1(n8582), .A2(n6962), .B1(P2_U3151), .B2(n6468), .C1(
        n7477), .C2(n8578), .ZN(P2_U3274) );
  AOI22_X1 U8626 ( .A1(n6945), .A2(n8874), .B1(n6944), .B2(n6943), .ZN(n10069)
         );
  NAND2_X1 U8627 ( .A1(n10149), .A2(n10067), .ZN(n8950) );
  INV_X1 U8628 ( .A(n10067), .ZN(n10160) );
  NAND2_X1 U8629 ( .A1(n10166), .A2(n10160), .ZN(n8777) );
  OAI22_X1 U8630 ( .A1(n10069), .A2(n10068), .B1(n10166), .B2(n10067), .ZN(
        n6964) );
  NAND2_X1 U8631 ( .A1(n6963), .A2(n6951), .ZN(n7026) );
  INV_X1 U8632 ( .A(n6951), .ZN(n10169) );
  NAND2_X1 U8633 ( .A1(n10065), .A2(n10169), .ZN(n8878) );
  NAND2_X1 U8634 ( .A1(n7026), .A2(n8878), .ZN(n8769) );
  INV_X1 U8635 ( .A(n8769), .ZN(n8779) );
  XNOR2_X1 U8636 ( .A(n6964), .B(n8779), .ZN(n10173) );
  NAND2_X1 U8637 ( .A1(n6947), .A2(n6946), .ZN(n6948) );
  NAND2_X1 U8638 ( .A1(n6948), .A2(n8775), .ZN(n10063) );
  INV_X1 U8639 ( .A(n8950), .ZN(n8765) );
  OAI21_X1 U8640 ( .B1(n10063), .B2(n8765), .A(n8777), .ZN(n6949) );
  NOR2_X1 U8641 ( .A1(n6949), .A2(n8769), .ZN(n7028) );
  AOI21_X1 U8642 ( .B1(n8769), .B2(n6949), .A(n7028), .ZN(n6950) );
  NOR2_X1 U8643 ( .A1(n6950), .A2(n10222), .ZN(n10171) );
  NAND2_X1 U8644 ( .A1(n10071), .A2(n10160), .ZN(n10070) );
  AOI21_X1 U8645 ( .B1(n10070), .B2(n6951), .A(n9339), .ZN(n6952) );
  OR2_X1 U8646 ( .A1(n10070), .A2(n6951), .ZN(n10056) );
  NAND2_X1 U8647 ( .A1(n6952), .A2(n10056), .ZN(n10168) );
  OR2_X1 U8648 ( .A1(n9192), .A2(n7022), .ZN(n6955) );
  AOI22_X1 U8649 ( .A1(n4495), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n6953), .B2(
        n10092), .ZN(n6954) );
  OAI211_X1 U8650 ( .C1(n9348), .C2(n10149), .A(n6955), .B(n6954), .ZN(n6957)
         );
  NOR2_X1 U8651 ( .A1(n9341), .A2(n10169), .ZN(n6956) );
  NOR2_X1 U8652 ( .A1(n6957), .A2(n6956), .ZN(n6958) );
  OAI21_X1 U8653 ( .B1(n10168), .B2(n9327), .A(n6958), .ZN(n6959) );
  AOI21_X1 U8654 ( .B1(n10171), .B2(n9309), .A(n6959), .ZN(n6960) );
  OAI21_X1 U8655 ( .B1(n10173), .B2(n9322), .A(n6960), .ZN(P1_U3286) );
  OAI222_X1 U8656 ( .A1(P1_U3086), .A2(n8939), .B1(n9820), .B2(n6962), .C1(
        n6961), .C2(n9814), .ZN(P1_U3334) );
  AOI22_X1 U8657 ( .A1(n6964), .A2(n8769), .B1(n10169), .B2(n6963), .ZN(n10055) );
  NAND2_X1 U8658 ( .A1(n7022), .A2(n10053), .ZN(n8783) );
  NAND2_X1 U8659 ( .A1(n10184), .A2(n10179), .ZN(n8781) );
  INV_X1 U8660 ( .A(n10193), .ZN(n6975) );
  NAND2_X1 U8661 ( .A1(n6975), .A2(n10183), .ZN(n8795) );
  INV_X1 U8662 ( .A(n10183), .ZN(n6971) );
  NAND2_X1 U8663 ( .A1(n10193), .A2(n6971), .ZN(n8786) );
  NAND2_X1 U8664 ( .A1(n8795), .A2(n8786), .ZN(n7029) );
  INV_X1 U8665 ( .A(n7393), .ZN(n10197) );
  NAND2_X1 U8666 ( .A1(n10197), .A2(n9012), .ZN(n8953) );
  INV_X1 U8667 ( .A(n9012), .ZN(n10205) );
  NAND2_X1 U8668 ( .A1(n7393), .A2(n10205), .ZN(n8956) );
  INV_X1 U8669 ( .A(n7103), .ZN(n8882) );
  XNOR2_X1 U8670 ( .A(n7104), .B(n8882), .ZN(n10199) );
  NAND2_X1 U8671 ( .A1(n8768), .A2(n8795), .ZN(n8883) );
  OR3_X1 U8672 ( .A1(n10063), .A2(n8765), .A3(n8883), .ZN(n6969) );
  NAND2_X1 U8673 ( .A1(n8781), .A2(n8786), .ZN(n6967) );
  NAND2_X1 U8674 ( .A1(n6967), .A2(n8795), .ZN(n6966) );
  NAND2_X1 U8675 ( .A1(n8883), .A2(n6966), .ZN(n8951) );
  INV_X1 U8676 ( .A(n6967), .ZN(n8879) );
  NAND3_X1 U8677 ( .A1(n8879), .A2(n8777), .A3(n8878), .ZN(n6968) );
  NAND2_X1 U8678 ( .A1(n8951), .A2(n6968), .ZN(n8952) );
  NAND2_X2 U8679 ( .A1(n6970), .A2(n7103), .ZN(n7176) );
  OAI21_X1 U8680 ( .B1(n6970), .B2(n7103), .A(n7176), .ZN(n10202) );
  NOR2_X4 U8681 ( .A1(n10056), .A2(n10053), .ZN(n10057) );
  OAI211_X1 U8682 ( .C1(n6972), .C2(n10197), .A(n10097), .B(n7171), .ZN(n10196) );
  NAND2_X1 U8683 ( .A1(n9344), .A2(n10192), .ZN(n6974) );
  AOI22_X1 U8684 ( .A1(n4495), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7387), .B2(
        n10092), .ZN(n6973) );
  OAI211_X1 U8685 ( .C1(n6975), .C2(n9348), .A(n6974), .B(n6973), .ZN(n6976)
         );
  AOI21_X1 U8686 ( .B1(n10090), .B2(n7393), .A(n6976), .ZN(n6977) );
  OAI21_X1 U8687 ( .B1(n10196), .B2(n9327), .A(n6977), .ZN(n6978) );
  AOI21_X1 U8688 ( .B1(n10202), .B2(n9301), .A(n6978), .ZN(n6979) );
  OAI21_X1 U8689 ( .B1(n10199), .B2(n9322), .A(n6979), .ZN(P1_U3283) );
  INV_X1 U8690 ( .A(n6980), .ZN(n6981) );
  INV_X1 U8691 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7276) );
  NOR2_X1 U8692 ( .A1(n7270), .A2(n7276), .ZN(n7196) );
  INV_X1 U8693 ( .A(n7196), .ZN(n6983) );
  OAI21_X1 U8694 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7201), .A(n6983), .ZN(
        n6984) );
  AOI21_X1 U8695 ( .B1(n4592), .B2(n6984), .A(n7197), .ZN(n7006) );
  INV_X1 U8696 ( .A(n6985), .ZN(n6990) );
  INV_X1 U8697 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7273) );
  MUX2_X1 U8698 ( .A(n7276), .B(n7273), .S(n8255), .Z(n6986) );
  NAND2_X1 U8699 ( .A1(n6986), .A2(n7270), .ZN(n7210) );
  INV_X1 U8700 ( .A(n6986), .ZN(n6987) );
  NAND2_X1 U8701 ( .A1(n6987), .A2(n7201), .ZN(n6988) );
  AND2_X1 U8702 ( .A1(n7210), .A2(n6988), .ZN(n6989) );
  OAI21_X1 U8703 ( .B1(n6991), .B2(n6990), .A(n6989), .ZN(n7211) );
  INV_X1 U8704 ( .A(n7211), .ZN(n6993) );
  NOR3_X1 U8705 ( .A1(n6991), .A2(n6990), .A3(n6989), .ZN(n6992) );
  OAI21_X1 U8706 ( .B1(n6993), .B2(n6992), .A(n10279), .ZN(n7005) );
  AOI22_X1 U8707 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n7201), .B1(n7270), .B2(
        n7273), .ZN(n6999) );
  NAND2_X1 U8708 ( .A1(n6995), .A2(n6994), .ZN(n6997) );
  OAI21_X1 U8709 ( .B1(n6999), .B2(n6998), .A(n7202), .ZN(n7003) );
  INV_X1 U8710 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n9679) );
  INV_X1 U8711 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7000) );
  NOR2_X1 U8712 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7000), .ZN(n7990) );
  AOI21_X1 U8713 ( .B1(n8202), .B2(n7270), .A(n7990), .ZN(n7001) );
  OAI21_X1 U8714 ( .B1(n9679), .B2(n8204), .A(n7001), .ZN(n7002) );
  AOI21_X1 U8715 ( .B1(n7003), .B2(n8267), .A(n7002), .ZN(n7004) );
  OAI211_X1 U8716 ( .C1(n7006), .C2(n8268), .A(n7005), .B(n7004), .ZN(P2_U3194) );
  NOR2_X1 U8717 ( .A1(n7009), .A2(n7008), .ZN(n7011) );
  XNOR2_X1 U8718 ( .A(n7900), .B(n7054), .ZN(n7033) );
  XNOR2_X1 U8719 ( .A(n7033), .B(n8112), .ZN(n7010) );
  OAI21_X1 U8720 ( .B1(n7011), .B2(n7010), .A(n7034), .ZN(n7012) );
  NAND2_X1 U8721 ( .A1(n7012), .A2(n8066), .ZN(n7019) );
  INV_X1 U8722 ( .A(n7013), .ZN(n7017) );
  INV_X1 U8723 ( .A(n8111), .ZN(n7236) );
  AOI21_X1 U8724 ( .B1(n8080), .B2(n8113), .A(n7014), .ZN(n7015) );
  OAI21_X1 U8725 ( .B1(n8084), .B2(n7236), .A(n7015), .ZN(n7016) );
  AOI21_X1 U8726 ( .B1(n7017), .B2(n8081), .A(n7016), .ZN(n7018) );
  OAI211_X1 U8727 ( .C1(n10334), .C2(n8076), .A(n7019), .B(n7018), .ZN(
        P2_U3153) );
  XOR2_X1 U8728 ( .A(n7029), .B(n7020), .Z(n10187) );
  AOI22_X1 U8729 ( .A1(n4495), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7224), .B2(
        n10092), .ZN(n7021) );
  OAI21_X1 U8730 ( .B1(n9348), .B2(n7022), .A(n7021), .ZN(n7025) );
  XNOR2_X1 U8731 ( .A(n10057), .B(n10183), .ZN(n7023) );
  AOI22_X1 U8732 ( .A1(n7023), .A2(n10097), .B1(n10191), .B2(n9012), .ZN(
        n10186) );
  NOR2_X1 U8733 ( .A1(n10186), .A2(n9327), .ZN(n7024) );
  AOI211_X1 U8734 ( .C1(n10090), .C2(n10183), .A(n7025), .B(n7024), .ZN(n7032)
         );
  INV_X1 U8735 ( .A(n7026), .ZN(n7027) );
  NOR2_X1 U8736 ( .A1(n7028), .A2(n7027), .ZN(n10049) );
  NAND2_X1 U8737 ( .A1(n10049), .A2(n10054), .ZN(n10048) );
  NAND2_X1 U8738 ( .A1(n10048), .A2(n8781), .ZN(n7030) );
  XNOR2_X1 U8739 ( .A(n7030), .B(n7029), .ZN(n10189) );
  NAND2_X1 U8740 ( .A1(n10189), .A2(n9301), .ZN(n7031) );
  OAI211_X1 U8741 ( .C1(n10187), .C2(n9322), .A(n7032), .B(n7031), .ZN(
        P1_U3284) );
  NAND2_X1 U8742 ( .A1(n7036), .A2(n7671), .ZN(n7039) );
  AOI22_X1 U8743 ( .A1(n7456), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7454), .B2(
        n7037), .ZN(n7038) );
  XNOR2_X1 U8744 ( .A(n7900), .B(n10339), .ZN(n7235) );
  XNOR2_X1 U8745 ( .A(n7235), .B(n8111), .ZN(n7040) );
  XNOR2_X1 U8746 ( .A(n7238), .B(n7040), .ZN(n7052) );
  INV_X1 U8747 ( .A(n10339), .ZN(n7084) );
  NAND2_X1 U8748 ( .A1(n7560), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7046) );
  OR2_X1 U8749 ( .A1(n4494), .A2(n7041), .ZN(n7045) );
  XNOR2_X1 U8750 ( .A(n7076), .B(n7042), .ZN(n7234) );
  OR2_X1 U8751 ( .A1(n7078), .A2(n7234), .ZN(n7044) );
  OR2_X1 U8752 ( .A1(n7679), .A2(n7092), .ZN(n7043) );
  NAND4_X1 U8753 ( .A1(n7046), .A2(n7045), .A3(n7044), .A4(n7043), .ZN(n8110)
         );
  NAND2_X1 U8754 ( .A1(n8092), .A2(n8110), .ZN(n7048) );
  OAI211_X1 U8755 ( .C1(n5040), .C2(n8090), .A(n7048), .B(n7047), .ZN(n7050)
         );
  NOR2_X1 U8756 ( .A1(n8094), .A2(n7059), .ZN(n7049) );
  AOI211_X1 U8757 ( .C1(n7084), .C2(n8101), .A(n7050), .B(n7049), .ZN(n7051)
         );
  OAI21_X1 U8758 ( .B1(n7052), .B2(n8096), .A(n7051), .ZN(P2_U3161) );
  NAND2_X1 U8759 ( .A1(n7095), .A2(n7094), .ZN(n7053) );
  NAND2_X1 U8760 ( .A1(n8111), .A2(n10339), .ZN(n7739) );
  XNOR2_X1 U8761 ( .A(n7053), .B(n7700), .ZN(n10342) );
  INV_X1 U8762 ( .A(n10342), .ZN(n7065) );
  INV_X1 U8763 ( .A(n8110), .ZN(n7058) );
  OR2_X1 U8764 ( .A1(n8112), .A2(n7054), .ZN(n7055) );
  XOR2_X1 U8765 ( .A(n7083), .B(n7700), .Z(n7057) );
  OAI222_X1 U8766 ( .A1(n8426), .A2(n5040), .B1(n8424), .B2(n7058), .C1(n10301), .C2(n7057), .ZN(n10340) );
  NAND2_X1 U8767 ( .A1(n10340), .A2(n8433), .ZN(n7064) );
  OAI22_X1 U8768 ( .A1(n10299), .A2(n7060), .B1(n7059), .B2(n8430), .ZN(n7062)
         );
  NOR2_X1 U8769 ( .A1(n8361), .A2(n10339), .ZN(n7061) );
  NOR2_X1 U8770 ( .A1(n7062), .A2(n7061), .ZN(n7063) );
  OAI211_X1 U8771 ( .C1(n7065), .C2(n8420), .A(n7064), .B(n7063), .ZN(P2_U3225) );
  INV_X1 U8772 ( .A(n7488), .ZN(n7067) );
  OAI222_X1 U8773 ( .A1(n8578), .A2(n7489), .B1(n8582), .B2(n7067), .C1(n7066), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U8774 ( .A1(n7068), .A2(P1_U3086), .B1(n9820), .B2(n7067), .C1(
        n9604), .C2(n9814), .ZN(P1_U3333) );
  NAND2_X1 U8775 ( .A1(n7499), .A2(n9806), .ZN(n7069) );
  OAI211_X1 U8776 ( .C1(n7070), .C2(n9817), .A(n7069), .B(n9007), .ZN(P1_U3332) );
  NAND2_X1 U8777 ( .A1(n7499), .A2(n8568), .ZN(n7072) );
  NAND2_X1 U8778 ( .A1(n7071), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7874) );
  OAI211_X1 U8779 ( .C1(n7500), .C2(n8578), .A(n7072), .B(n7874), .ZN(P2_U3272) );
  NAND2_X1 U8780 ( .A1(n7560), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7082) );
  OR2_X1 U8781 ( .A1(n4494), .A2(n7073), .ZN(n7081) );
  NOR2_X1 U8782 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n7074) );
  OAI21_X1 U8783 ( .B1(n7076), .B2(P2_REG3_REG_9__SCAN_IN), .A(
        P2_REG3_REG_10__SCAN_IN), .ZN(n7077) );
  AND2_X1 U8784 ( .A1(n7157), .A2(n7077), .ZN(n7303) );
  OR2_X1 U8785 ( .A1(n7078), .A2(n7303), .ZN(n7080) );
  OR2_X1 U8786 ( .A1(n7679), .A2(n6671), .ZN(n7079) );
  NAND4_X1 U8787 ( .A1(n7082), .A2(n7081), .A3(n7080), .A4(n7079), .ZN(n8109)
         );
  OR2_X1 U8788 ( .A1(n8111), .A2(n7084), .ZN(n7085) );
  NAND2_X1 U8789 ( .A1(n7086), .A2(n7085), .ZN(n7151) );
  NAND2_X1 U8790 ( .A1(n7087), .A2(n7671), .ZN(n7090) );
  AOI22_X1 U8791 ( .A1(n7456), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7454), .B2(
        n7088), .ZN(n7089) );
  OR2_X1 U8792 ( .A1(n7239), .A2(n8110), .ZN(n7761) );
  NAND2_X1 U8793 ( .A1(n7239), .A2(n8110), .ZN(n7757) );
  NAND2_X1 U8794 ( .A1(n7761), .A2(n7757), .ZN(n7698) );
  XOR2_X1 U8795 ( .A(n7151), .B(n7698), .Z(n7091) );
  OAI222_X1 U8796 ( .A1(n8426), .A2(n7236), .B1(n8424), .B2(n7982), .C1(n10301), .C2(n7091), .ZN(n10346) );
  INV_X1 U8797 ( .A(n10346), .ZN(n7101) );
  INV_X1 U8798 ( .A(n7239), .ZN(n10348) );
  OAI22_X1 U8799 ( .A1(n10299), .A2(n7092), .B1(n7234), .B2(n8430), .ZN(n7093)
         );
  AOI21_X1 U8800 ( .B1(n10292), .B2(n10348), .A(n7093), .ZN(n7100) );
  AND2_X1 U8801 ( .A1(n7094), .A2(n7739), .ZN(n7758) );
  NAND2_X1 U8802 ( .A1(n7095), .A2(n7758), .ZN(n7096) );
  INV_X1 U8803 ( .A(n7698), .ZN(n7097) );
  NAND2_X1 U8804 ( .A1(n7098), .A2(n7698), .ZN(n10344) );
  NAND3_X1 U8805 ( .A1(n7145), .A2(n10344), .A3(n10296), .ZN(n7099) );
  OAI211_X1 U8806 ( .C1(n7101), .C2(n8381), .A(n7100), .B(n7099), .ZN(P2_U3224) );
  NAND2_X1 U8807 ( .A1(n10209), .A2(n10216), .ZN(n8957) );
  AND2_X1 U8808 ( .A1(n8957), .A2(n8956), .ZN(n8797) );
  NAND2_X1 U8809 ( .A1(n7176), .A2(n8797), .ZN(n7183) );
  NAND2_X1 U8810 ( .A1(n7183), .A2(n8787), .ZN(n7102) );
  OR2_X1 U8811 ( .A1(n10219), .A2(n10206), .ZN(n8790) );
  NAND2_X1 U8812 ( .A1(n10219), .A2(n10206), .ZN(n8962) );
  XNOR2_X1 U8813 ( .A(n7102), .B(n8885), .ZN(n10221) );
  NAND2_X1 U8814 ( .A1(n8787), .A2(n8957), .ZN(n8881) );
  INV_X1 U8815 ( .A(n10209), .ZN(n7175) );
  XNOR2_X1 U8816 ( .A(n7182), .B(n8885), .ZN(n10224) );
  NAND2_X1 U8817 ( .A1(n10224), .A2(n10102), .ZN(n7110) );
  AOI211_X1 U8818 ( .C1(n10219), .C2(n7169), .A(n9339), .B(n7189), .ZN(n10217)
         );
  AOI22_X1 U8819 ( .A1(n4495), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7401), .B2(
        n10092), .ZN(n7105) );
  OAI21_X1 U8820 ( .B1(n9348), .B2(n10216), .A(n7105), .ZN(n7106) );
  AOI21_X1 U8821 ( .B1(n9344), .B2(n9010), .A(n7106), .ZN(n7107) );
  OAI21_X1 U8822 ( .B1(n4798), .B2(n9341), .A(n7107), .ZN(n7108) );
  AOI21_X1 U8823 ( .B1(n10217), .B2(n10101), .A(n7108), .ZN(n7109) );
  OAI211_X1 U8824 ( .C1(n10221), .C2(n9353), .A(n7110), .B(n7109), .ZN(
        P1_U3281) );
  INV_X1 U8825 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9906) );
  AOI22_X1 U8826 ( .A1(n9064), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9906), .B2(
        n7127), .ZN(n7117) );
  OAI21_X1 U8827 ( .B1(n7120), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7111), .ZN(
        n9996) );
  INV_X1 U8828 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7112) );
  MUX2_X1 U8829 ( .A(n7112), .B(P1_REG1_REG_13__SCAN_IN), .S(n10003), .Z(n9997) );
  NOR2_X1 U8830 ( .A1(n9996), .A2(n9997), .ZN(n9995) );
  INV_X1 U8831 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7113) );
  MUX2_X1 U8832 ( .A(n7113), .B(P1_REG1_REG_14__SCAN_IN), .S(n10015), .Z(
        n10011) );
  NOR2_X1 U8833 ( .A1(n10012), .A2(n10011), .ZN(n10010) );
  NOR2_X1 U8834 ( .A1(n7114), .A2(n7125), .ZN(n7115) );
  INV_X1 U8835 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10021) );
  XNOR2_X1 U8836 ( .A(n7125), .B(n7114), .ZN(n10022) );
  NOR2_X1 U8837 ( .A1(n10021), .A2(n10022), .ZN(n10020) );
  NOR2_X1 U8838 ( .A1(n7115), .A2(n10020), .ZN(n7116) );
  NAND2_X1 U8839 ( .A1(n7117), .A2(n7116), .ZN(n9063) );
  OAI21_X1 U8840 ( .B1(n7117), .B2(n7116), .A(n9063), .ZN(n7133) );
  NAND2_X1 U8841 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8648) );
  NAND2_X1 U8842 ( .A1(n9945), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7118) );
  OAI211_X1 U8843 ( .C1(n9070), .C2(n7127), .A(n8648), .B(n7118), .ZN(n7132)
         );
  OAI21_X1 U8844 ( .B1(n7120), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7119), .ZN(
        n10000) );
  INV_X1 U8845 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7121) );
  MUX2_X1 U8846 ( .A(n7121), .B(P1_REG2_REG_13__SCAN_IN), .S(n10003), .Z(n9999) );
  NOR2_X1 U8847 ( .A1(n10000), .A2(n9999), .ZN(n9998) );
  INV_X1 U8848 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7123) );
  AOI22_X1 U8849 ( .A1(n10015), .A2(n7123), .B1(P1_REG2_REG_14__SCAN_IN), .B2(
        n7122), .ZN(n10008) );
  NOR2_X1 U8850 ( .A1(n7124), .A2(n7125), .ZN(n7126) );
  INV_X1 U8851 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10024) );
  NOR2_X1 U8852 ( .A1(n10024), .A2(n10025), .ZN(n10023) );
  NOR2_X1 U8853 ( .A1(n7126), .A2(n10023), .ZN(n7130) );
  INV_X1 U8854 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7128) );
  AOI22_X1 U8855 ( .A1(n9064), .A2(n7128), .B1(P1_REG2_REG_16__SCAN_IN), .B2(
        n7127), .ZN(n7129) );
  NOR2_X1 U8856 ( .A1(n7130), .A2(n7129), .ZN(n9059) );
  INV_X1 U8857 ( .A(n9983), .ZN(n10036) );
  AOI211_X1 U8858 ( .C1(n7130), .C2(n7129), .A(n9059), .B(n10036), .ZN(n7131)
         );
  AOI211_X1 U8859 ( .C1(n9988), .C2(n7133), .A(n7132), .B(n7131), .ZN(n7134)
         );
  INV_X1 U8860 ( .A(n7134), .ZN(P1_U3259) );
  AOI21_X1 U8861 ( .B1(n7137), .B2(n7136), .A(n7135), .ZN(n7144) );
  INV_X1 U8862 ( .A(n10052), .ZN(n7141) );
  NOR2_X1 U8863 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7138), .ZN(n9864) );
  AOI21_X1 U8864 ( .B1(n8726), .B2(n10065), .A(n9864), .ZN(n7140) );
  NAND2_X1 U8865 ( .A1(n8693), .A2(n10193), .ZN(n7139) );
  OAI211_X1 U8866 ( .C1(n8696), .C2(n7141), .A(n7140), .B(n7139), .ZN(n7142)
         );
  AOI21_X1 U8867 ( .B1(n10053), .B2(n8731), .A(n7142), .ZN(n7143) );
  OAI21_X1 U8868 ( .B1(n7144), .B2(n8733), .A(n7143), .ZN(P1_U3221) );
  NAND2_X1 U8869 ( .A1(n7146), .A2(n7671), .ZN(n7149) );
  AOI22_X1 U8870 ( .A1(n7456), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7454), .B2(
        n7147), .ZN(n7148) );
  NAND2_X1 U8871 ( .A1(n7149), .A2(n7148), .ZN(n7305) );
  INV_X1 U8872 ( .A(n7305), .ZN(n10350) );
  AND2_X1 U8873 ( .A1(n10350), .A2(n8109), .ZN(n7756) );
  NAND2_X1 U8874 ( .A1(n7305), .A2(n7982), .ZN(n7767) );
  INV_X1 U8875 ( .A(n7767), .ZN(n7150) );
  NOR2_X1 U8876 ( .A1(n7756), .A2(n7150), .ZN(n7703) );
  XNOR2_X1 U8877 ( .A(n7263), .B(n7703), .ZN(n10352) );
  NAND2_X1 U8878 ( .A1(n7151), .A2(n7698), .ZN(n7153) );
  OR2_X1 U8879 ( .A1(n8110), .A2(n10348), .ZN(n7152) );
  NAND2_X1 U8880 ( .A1(n7153), .A2(n7152), .ZN(n7289) );
  XOR2_X1 U8881 ( .A(n7289), .B(n7703), .Z(n7154) );
  NAND2_X1 U8882 ( .A1(n7154), .A2(n10289), .ZN(n7164) );
  OR2_X1 U8883 ( .A1(n4494), .A2(n7155), .ZN(n7162) );
  INV_X1 U8884 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7156) );
  OR2_X1 U8885 ( .A1(n7526), .A2(n7156), .ZN(n7161) );
  NAND2_X1 U8886 ( .A1(n7157), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7158) );
  AND2_X1 U8887 ( .A1(n7274), .A2(n7158), .ZN(n8057) );
  OR2_X1 U8888 ( .A1(n7078), .A2(n8057), .ZN(n7160) );
  OR2_X1 U8889 ( .A1(n7679), .A2(n7610), .ZN(n7159) );
  NAND4_X1 U8890 ( .A1(n7162), .A2(n7161), .A3(n7160), .A4(n7159), .ZN(n8108)
         );
  AOI22_X1 U8891 ( .A1(n10285), .A2(n8110), .B1(n8108), .B2(n10286), .ZN(n7163) );
  OAI211_X1 U8892 ( .C1(n10352), .C2(n10309), .A(n7164), .B(n7163), .ZN(n10354) );
  NAND2_X1 U8893 ( .A1(n10354), .A2(n10299), .ZN(n7167) );
  OAI22_X1 U8894 ( .A1(n10299), .A2(n6671), .B1(n7303), .B2(n8430), .ZN(n7165)
         );
  AOI21_X1 U8895 ( .B1(n10292), .B2(n7305), .A(n7165), .ZN(n7166) );
  OAI211_X1 U8896 ( .C1(n10352), .C2(n7937), .A(n7167), .B(n7166), .ZN(
        P2_U3223) );
  XOR2_X1 U8897 ( .A(n8881), .B(n7168), .Z(n10212) );
  INV_X1 U8898 ( .A(n7169), .ZN(n7170) );
  AOI211_X1 U8899 ( .C1(n10209), .C2(n7171), .A(n9339), .B(n7170), .ZN(n10207)
         );
  AOI22_X1 U8900 ( .A1(n4495), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8707), .B2(
        n10092), .ZN(n7172) );
  OAI21_X1 U8901 ( .B1(n9348), .B2(n10205), .A(n7172), .ZN(n7173) );
  AOI21_X1 U8902 ( .B1(n9344), .B2(n9011), .A(n7173), .ZN(n7174) );
  OAI21_X1 U8903 ( .B1(n7175), .B2(n9341), .A(n7174), .ZN(n7180) );
  NAND2_X1 U8904 ( .A1(n7176), .A2(n8956), .ZN(n7177) );
  XNOR2_X1 U8905 ( .A(n7177), .B(n4850), .ZN(n7178) );
  NAND2_X1 U8906 ( .A1(n7178), .A2(n10203), .ZN(n10210) );
  NOR2_X1 U8907 ( .A1(n10210), .A2(n4495), .ZN(n7179) );
  AOI211_X1 U8908 ( .C1(n10207), .C2(n10101), .A(n7180), .B(n7179), .ZN(n7181)
         );
  OAI21_X1 U8909 ( .B1(n10212), .B2(n9322), .A(n7181), .ZN(P1_U3282) );
  OR2_X1 U8910 ( .A1(n7190), .A2(n10235), .ZN(n8966) );
  NAND2_X1 U8911 ( .A1(n7190), .A2(n10235), .ZN(n8963) );
  NAND2_X1 U8912 ( .A1(n8966), .A2(n8963), .ZN(n7248) );
  XNOR2_X1 U8913 ( .A(n7249), .B(n7248), .ZN(n10232) );
  INV_X1 U8914 ( .A(n10232), .ZN(n7195) );
  INV_X1 U8915 ( .A(n7248), .ZN(n8886) );
  AND2_X1 U8916 ( .A1(n8790), .A2(n8787), .ZN(n8961) );
  NAND2_X1 U8917 ( .A1(n7183), .A2(n8961), .ZN(n7184) );
  NAND2_X1 U8918 ( .A1(n7184), .A2(n8962), .ZN(n7185) );
  NAND2_X2 U8919 ( .A1(n7185), .A2(n8886), .ZN(n7257) );
  OAI21_X1 U8920 ( .B1(n8886), .B2(n7185), .A(n7257), .ZN(n7186) );
  NAND2_X1 U8921 ( .A1(n7186), .A2(n10203), .ZN(n7188) );
  AOI22_X1 U8922 ( .A1(n10194), .A2(n9011), .B1(n9103), .B2(n10191), .ZN(n7187) );
  NAND2_X1 U8923 ( .A1(n7188), .A2(n7187), .ZN(n10230) );
  AND2_X2 U8924 ( .A1(n7189), .A2(n10228), .ZN(n7250) );
  INV_X1 U8925 ( .A(n7250), .ZN(n7252) );
  OAI211_X1 U8926 ( .C1(n10228), .C2(n7189), .A(n7252), .B(n10097), .ZN(n10226) );
  AOI22_X1 U8927 ( .A1(n4495), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8686), .B2(
        n10092), .ZN(n7192) );
  NAND2_X1 U8928 ( .A1(n7190), .A2(n10090), .ZN(n7191) );
  OAI211_X1 U8929 ( .C1(n10226), .C2(n9327), .A(n7192), .B(n7191), .ZN(n7193)
         );
  AOI21_X1 U8930 ( .B1(n10230), .B2(n9309), .A(n7193), .ZN(n7194) );
  OAI21_X1 U8931 ( .B1(n7195), .B2(n9322), .A(n7194), .ZN(P1_U3280) );
  NAND2_X1 U8932 ( .A1(n7198), .A2(n8122), .ZN(n8117) );
  INV_X1 U8933 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7199) );
  AOI21_X1 U8934 ( .B1(n7200), .B2(n7199), .A(n8118), .ZN(n7218) );
  NAND2_X1 U8935 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n7201), .ZN(n7203) );
  NAND2_X1 U8936 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n7204), .ZN(n8124) );
  OAI21_X1 U8937 ( .B1(n7204), .B2(P2_REG1_REG_13__SCAN_IN), .A(n8124), .ZN(
        n7216) );
  INV_X1 U8938 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n9666) );
  AND2_X1 U8939 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7334) );
  AOI21_X1 U8940 ( .B1(n8202), .B2(n7320), .A(n7334), .ZN(n7205) );
  OAI21_X1 U8941 ( .B1(n9666), .B2(n8204), .A(n7205), .ZN(n7215) );
  INV_X1 U8942 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7353) );
  MUX2_X1 U8943 ( .A(n7199), .B(n7353), .S(n8255), .Z(n7206) );
  NAND2_X1 U8944 ( .A1(n7206), .A2(n7320), .ZN(n8132) );
  INV_X1 U8945 ( .A(n7206), .ZN(n7207) );
  NAND2_X1 U8946 ( .A1(n7207), .A2(n8122), .ZN(n7208) );
  NAND2_X1 U8947 ( .A1(n8132), .A2(n7208), .ZN(n7209) );
  AOI21_X1 U8948 ( .B1(n7211), .B2(n7210), .A(n7209), .ZN(n8138) );
  INV_X1 U8949 ( .A(n8138), .ZN(n7213) );
  NAND3_X1 U8950 ( .A1(n7211), .A2(n7210), .A3(n7209), .ZN(n7212) );
  AOI21_X1 U8951 ( .B1(n7213), .B2(n7212), .A(n8264), .ZN(n7214) );
  AOI211_X1 U8952 ( .C1(n8267), .C2(n7216), .A(n7215), .B(n7214), .ZN(n7217)
         );
  OAI21_X1 U8953 ( .B1(n7218), .B2(n8268), .A(n7217), .ZN(P2_U3195) );
  INV_X1 U8954 ( .A(n7507), .ZN(n7220) );
  OAI222_X1 U8955 ( .A1(n8582), .A2(n7220), .B1(P2_U3151), .B2(n6026), .C1(
        n7508), .C2(n8578), .ZN(P2_U3271) );
  OAI222_X1 U8956 ( .A1(P1_U3086), .A2(n7221), .B1(n9820), .B2(n7220), .C1(
        n7219), .C2(n9814), .ZN(P1_U3331) );
  NOR2_X1 U8957 ( .A1(n7222), .A2(n4600), .ZN(n7223) );
  XNOR2_X1 U8958 ( .A(n4531), .B(n7223), .ZN(n7230) );
  NAND2_X1 U8959 ( .A1(n8725), .A2(n7224), .ZN(n7227) );
  AOI21_X1 U8960 ( .B1(n8726), .B2(n10184), .A(n7225), .ZN(n7226) );
  OAI211_X1 U8961 ( .C1(n10205), .C2(n8729), .A(n7227), .B(n7226), .ZN(n7228)
         );
  AOI21_X1 U8962 ( .B1(n10183), .B2(n8731), .A(n7228), .ZN(n7229) );
  OAI21_X1 U8963 ( .B1(n7230), .B2(n8733), .A(n7229), .ZN(P1_U3231) );
  INV_X1 U8964 ( .A(n7516), .ZN(n7245) );
  OAI222_X1 U8965 ( .A1(n8582), .A2(n7245), .B1(P2_U3151), .B2(n6027), .C1(
        n7517), .C2(n8578), .ZN(P2_U3270) );
  AOI21_X1 U8966 ( .B1(n8080), .B2(n8111), .A(n7231), .ZN(n7233) );
  NAND2_X1 U8967 ( .A1(n8092), .A2(n8109), .ZN(n7232) );
  OAI211_X1 U8968 ( .C1(n8094), .C2(n7234), .A(n7233), .B(n7232), .ZN(n7242)
         );
  NOR2_X1 U8969 ( .A1(n7235), .A2(n8111), .ZN(n7237) );
  XNOR2_X1 U8970 ( .A(n7239), .B(n7900), .ZN(n7296) );
  XOR2_X1 U8971 ( .A(n8110), .B(n7296), .Z(n7297) );
  XNOR2_X1 U8972 ( .A(n7298), .B(n7297), .ZN(n7240) );
  NOR2_X1 U8973 ( .A1(n7240), .A2(n8096), .ZN(n7241) );
  AOI211_X1 U8974 ( .C1(n10348), .C2(n8101), .A(n7242), .B(n7241), .ZN(n7243)
         );
  INV_X1 U8975 ( .A(n7243), .ZN(P2_U3171) );
  OAI222_X1 U8976 ( .A1(P1_U3086), .A2(n7246), .B1(n9820), .B2(n7245), .C1(
        n7244), .C2(n9814), .ZN(P1_U3330) );
  NAND2_X1 U8977 ( .A1(n10240), .A2(n9907), .ZN(n8806) );
  NAND2_X1 U8978 ( .A1(n8967), .A2(n8806), .ZN(n7256) );
  XNOR2_X1 U8979 ( .A(n9106), .B(n7256), .ZN(n10245) );
  INV_X1 U8980 ( .A(n10240), .ZN(n9102) );
  INV_X1 U8981 ( .A(n9340), .ZN(n7251) );
  AOI211_X1 U8982 ( .C1(n10240), .C2(n7252), .A(n9339), .B(n7251), .ZN(n10238)
         );
  AOI22_X1 U8983 ( .A1(n4495), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8599), .B2(
        n10092), .ZN(n7253) );
  OAI21_X1 U8984 ( .B1(n9348), .B2(n10235), .A(n7253), .ZN(n7254) );
  AOI21_X1 U8985 ( .B1(n9344), .B2(n9897), .A(n7254), .ZN(n7255) );
  OAI21_X1 U8986 ( .B1(n9102), .B2(n9341), .A(n7255), .ZN(n7261) );
  INV_X1 U8987 ( .A(n8963), .ZN(n8959) );
  NOR2_X1 U8988 ( .A1(n7256), .A2(n8959), .ZN(n8802) );
  NAND2_X1 U8989 ( .A1(n7257), .A2(n8802), .ZN(n8905) );
  INV_X1 U8990 ( .A(n8905), .ZN(n7259) );
  INV_X1 U8991 ( .A(n7256), .ZN(n8887) );
  AOI21_X1 U8992 ( .B1(n7257), .B2(n8963), .A(n8887), .ZN(n7258) );
  NOR2_X1 U8993 ( .A1(n10242), .A2(n4495), .ZN(n7260) );
  AOI211_X1 U8994 ( .C1(n10238), .C2(n10101), .A(n7261), .B(n7260), .ZN(n7262)
         );
  OAI21_X1 U8995 ( .B1(n10245), .B2(n9322), .A(n7262), .ZN(P1_U3279) );
  NAND2_X1 U8996 ( .A1(n7264), .A2(n7767), .ZN(n7604) );
  NAND2_X1 U8997 ( .A1(n7265), .A2(n7671), .ZN(n7268) );
  AOI22_X1 U8998 ( .A1(n7456), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n7454), .B2(
        n7266), .ZN(n7267) );
  NAND2_X1 U8999 ( .A1(n7268), .A2(n7267), .ZN(n8050) );
  XNOR2_X1 U9000 ( .A(n8050), .B(n8108), .ZN(n7692) );
  INV_X1 U9001 ( .A(n8108), .ZN(n7988) );
  AND2_X1 U9002 ( .A1(n8050), .A2(n7988), .ZN(n7716) );
  NAND2_X1 U9003 ( .A1(n7269), .A2(n7671), .ZN(n7272) );
  AOI22_X1 U9004 ( .A1(n7456), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7454), .B2(
        n7270), .ZN(n7271) );
  NAND2_X1 U9005 ( .A1(n7560), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7280) );
  OR2_X1 U9006 ( .A1(n4494), .A2(n7273), .ZN(n7279) );
  NAND2_X1 U9007 ( .A1(n7274), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7275) );
  AND2_X1 U9008 ( .A1(n7283), .A2(n7275), .ZN(n7992) );
  OR2_X1 U9009 ( .A1(n7078), .A2(n7992), .ZN(n7278) );
  OR2_X1 U9010 ( .A1(n7679), .A2(n7276), .ZN(n7277) );
  NAND4_X1 U9011 ( .A1(n7280), .A2(n7279), .A3(n7278), .A4(n7277), .ZN(n8107)
         );
  NAND2_X1 U9012 ( .A1(n10365), .A2(n7609), .ZN(n7718) );
  OAI21_X1 U9013 ( .B1(n7281), .B2(n7693), .A(n7347), .ZN(n10362) );
  INV_X1 U9014 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9636) );
  OR2_X1 U9015 ( .A1(n7526), .A2(n9636), .ZN(n7288) );
  OR2_X1 U9016 ( .A1(n4494), .A2(n7353), .ZN(n7287) );
  NAND2_X1 U9017 ( .A1(n7283), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7284) );
  AND2_X1 U9018 ( .A1(n7327), .A2(n7284), .ZN(n7348) );
  OR2_X1 U9019 ( .A1(n7078), .A2(n7348), .ZN(n7286) );
  OR2_X1 U9020 ( .A1(n7679), .A2(n7199), .ZN(n7285) );
  NAND4_X1 U9021 ( .A1(n7288), .A2(n7287), .A3(n7286), .A4(n7285), .ZN(n8106)
         );
  INV_X1 U9022 ( .A(n8106), .ZN(n8425) );
  INV_X1 U9023 ( .A(n7289), .ZN(n7290) );
  NAND2_X1 U9024 ( .A1(n7305), .A2(n8109), .ZN(n7606) );
  AND2_X1 U9025 ( .A1(n4567), .A2(n7606), .ZN(n7291) );
  XNOR2_X1 U9026 ( .A(n7340), .B(n7693), .ZN(n7292) );
  OAI222_X1 U9027 ( .A1(n8424), .A2(n8425), .B1(n8426), .B2(n7988), .C1(n10301), .C2(n7292), .ZN(n10363) );
  NAND2_X1 U9028 ( .A1(n10363), .A2(n10299), .ZN(n7295) );
  OAI22_X1 U9029 ( .A1(n8433), .A2(n7276), .B1(n7992), .B2(n8430), .ZN(n7293)
         );
  AOI21_X1 U9030 ( .B1(n10292), .B2(n10365), .A(n7293), .ZN(n7294) );
  OAI211_X1 U9031 ( .C1(n8420), .C2(n10362), .A(n7295), .B(n7294), .ZN(
        P2_U3221) );
  XNOR2_X1 U9032 ( .A(n7305), .B(n7900), .ZN(n7308) );
  INV_X1 U9033 ( .A(n7308), .ZN(n7311) );
  XNOR2_X1 U9034 ( .A(n7983), .B(n7982), .ZN(n7299) );
  NOR2_X1 U9035 ( .A1(n7299), .A2(n7311), .ZN(n7981) );
  AOI21_X1 U9036 ( .B1(n7311), .B2(n7299), .A(n7981), .ZN(n7307) );
  AOI21_X1 U9037 ( .B1(n8080), .B2(n8110), .A(n7300), .ZN(n7302) );
  NAND2_X1 U9038 ( .A1(n8092), .A2(n8108), .ZN(n7301) );
  OAI211_X1 U9039 ( .C1(n7303), .C2(n8094), .A(n7302), .B(n7301), .ZN(n7304)
         );
  AOI21_X1 U9040 ( .B1(n7305), .B2(n8101), .A(n7304), .ZN(n7306) );
  OAI21_X1 U9041 ( .B1(n7307), .B2(n8096), .A(n7306), .ZN(P2_U3157) );
  XNOR2_X1 U9042 ( .A(n8050), .B(n6486), .ZN(n7984) );
  NAND2_X1 U9043 ( .A1(n7984), .A2(n8108), .ZN(n7985) );
  INV_X1 U9044 ( .A(n7985), .ZN(n7310) );
  INV_X1 U9045 ( .A(n7984), .ZN(n7314) );
  OAI21_X1 U9046 ( .B1(n7311), .B2(n8109), .A(n8108), .ZN(n7313) );
  NOR3_X1 U9047 ( .A1(n7311), .A2(n8109), .A3(n8108), .ZN(n7312) );
  XNOR2_X1 U9048 ( .A(n10365), .B(n7900), .ZN(n7315) );
  XNOR2_X1 U9049 ( .A(n7315), .B(n7609), .ZN(n7987) );
  AOI211_X1 U9050 ( .C1(n7314), .C2(n7313), .A(n7312), .B(n7987), .ZN(n7317)
         );
  INV_X1 U9051 ( .A(n7315), .ZN(n7316) );
  NAND2_X1 U9052 ( .A1(n7319), .A2(n7671), .ZN(n7322) );
  AOI22_X1 U9053 ( .A1(n7456), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7454), .B2(
        n7320), .ZN(n7321) );
  XNOR2_X1 U9054 ( .A(n7416), .B(n6486), .ZN(n7323) );
  NOR2_X1 U9055 ( .A1(n7323), .A2(n8106), .ZN(n7372) );
  INV_X1 U9056 ( .A(n7372), .ZN(n7324) );
  NAND2_X1 U9057 ( .A1(n7323), .A2(n8106), .ZN(n7371) );
  NAND2_X1 U9058 ( .A1(n7324), .A2(n7371), .ZN(n7325) );
  XNOR2_X1 U9059 ( .A(n7373), .B(n7325), .ZN(n7338) );
  INV_X1 U9060 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9623) );
  OR2_X1 U9061 ( .A1(n7526), .A2(n9623), .ZN(n7332) );
  INV_X1 U9062 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8432) );
  OR2_X1 U9063 ( .A1(n7679), .A2(n8432), .ZN(n7331) );
  NAND2_X1 U9064 ( .A1(n7327), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7328) );
  AND2_X1 U9065 ( .A1(n7374), .A2(n7328), .ZN(n8431) );
  OR2_X1 U9066 ( .A1(n7078), .A2(n8431), .ZN(n7330) );
  INV_X1 U9067 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9471) );
  OR2_X1 U9068 ( .A1(n4494), .A2(n9471), .ZN(n7329) );
  NAND4_X1 U9069 ( .A1(n7332), .A2(n7331), .A3(n7330), .A4(n7329), .ZN(n8413)
         );
  NOR2_X1 U9070 ( .A1(n8090), .A2(n7609), .ZN(n7333) );
  AOI211_X1 U9071 ( .C1(n8092), .C2(n8413), .A(n7334), .B(n7333), .ZN(n7335)
         );
  OAI21_X1 U9072 ( .B1(n7348), .B2(n8094), .A(n7335), .ZN(n7336) );
  AOI21_X1 U9073 ( .B1(n7416), .B2(n8101), .A(n7336), .ZN(n7337) );
  OAI21_X1 U9074 ( .B1(n7338), .B2(n8096), .A(n7337), .ZN(P2_U3174) );
  INV_X1 U9075 ( .A(n8308), .ZN(n8427) );
  NAND2_X1 U9076 ( .A1(n10365), .A2(n8107), .ZN(n7339) );
  OR2_X1 U9077 ( .A1(n7416), .A2(n8106), .ZN(n7342) );
  NAND2_X1 U9078 ( .A1(n7343), .A2(n7342), .ZN(n7567) );
  NAND2_X1 U9079 ( .A1(n7416), .A2(n8106), .ZN(n7566) );
  INV_X1 U9080 ( .A(n7566), .ZN(n7341) );
  NOR2_X1 U9081 ( .A1(n7567), .A2(n7341), .ZN(n7346) );
  NAND2_X1 U9082 ( .A1(n7342), .A2(n7566), .ZN(n7701) );
  INV_X1 U9083 ( .A(n7701), .ZN(n7775) );
  OAI21_X1 U9084 ( .B1(n7343), .B2(n7775), .A(n10289), .ZN(n7345) );
  AOI22_X1 U9085 ( .A1(n10286), .A2(n8413), .B1(n8107), .B2(n10285), .ZN(n7344) );
  OAI21_X1 U9086 ( .B1(n7346), .B2(n7345), .A(n7344), .ZN(n7352) );
  AOI21_X1 U9087 ( .B1(n8427), .B2(n7416), .A(n7352), .ZN(n7351) );
  XNOR2_X1 U9088 ( .A(n7415), .B(n7775), .ZN(n7365) );
  OAI22_X1 U9089 ( .A1(n8433), .A2(n7199), .B1(n7348), .B2(n8430), .ZN(n7349)
         );
  AOI21_X1 U9090 ( .B1(n7365), .B2(n10296), .A(n7349), .ZN(n7350) );
  OAI21_X1 U9091 ( .B1(n7351), .B2(n8381), .A(n7350), .ZN(P2_U3220) );
  INV_X1 U9092 ( .A(n7352), .ZN(n7364) );
  MUX2_X1 U9093 ( .A(n7353), .B(n7364), .S(n10386), .Z(n7355) );
  NAND2_X1 U9094 ( .A1(n10386), .A2(n10345), .ZN(n8484) );
  INV_X1 U9095 ( .A(n8484), .ZN(n8487) );
  NAND2_X1 U9096 ( .A1(n10386), .A2(n10366), .ZN(n8470) );
  AOI22_X1 U9097 ( .A1(n7365), .A2(n8487), .B1(n8486), .B2(n7416), .ZN(n7354)
         );
  NAND2_X1 U9098 ( .A1(n7355), .A2(n7354), .ZN(P2_U3472) );
  NAND2_X1 U9099 ( .A1(n7357), .A2(n7356), .ZN(n7363) );
  NAND2_X1 U9100 ( .A1(n7359), .A2(n7358), .ZN(n7360) );
  NAND2_X1 U9101 ( .A1(n7361), .A2(n7360), .ZN(n7362) );
  MUX2_X1 U9102 ( .A(n9636), .B(n7364), .S(n10367), .Z(n7367) );
  INV_X1 U9103 ( .A(n10345), .ZN(n10361) );
  INV_X1 U9104 ( .A(n8555), .ZN(n8560) );
  AOI22_X1 U9105 ( .A1(n7365), .A2(n8560), .B1(n8559), .B2(n7416), .ZN(n7366)
         );
  NAND2_X1 U9106 ( .A1(n7367), .A2(n7366), .ZN(P2_U3429) );
  NAND2_X1 U9107 ( .A1(n7368), .A2(n7671), .ZN(n7370) );
  AOI22_X1 U9108 ( .A1(n7456), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7454), .B2(
        n8148), .ZN(n7369) );
  XNOR2_X1 U9109 ( .A(n8558), .B(n7900), .ZN(n7876) );
  INV_X1 U9110 ( .A(n8413), .ZN(n8089) );
  XNOR2_X1 U9111 ( .A(n7876), .B(n8089), .ZN(n7878) );
  XOR2_X1 U9112 ( .A(n7878), .B(n7879), .Z(n7384) );
  NAND2_X1 U9113 ( .A1(n7560), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7379) );
  INV_X1 U9114 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8481) );
  OR2_X1 U9115 ( .A1(n4494), .A2(n8481), .ZN(n7378) );
  NAND2_X1 U9116 ( .A1(n7374), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7375) );
  AND2_X1 U9117 ( .A1(n7427), .A2(n7375), .ZN(n8416) );
  OR2_X1 U9118 ( .A1(n7078), .A2(n8416), .ZN(n7377) );
  INV_X1 U9119 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8415) );
  OR2_X1 U9120 ( .A1(n7679), .A2(n8415), .ZN(n7376) );
  NAND4_X1 U9121 ( .A1(n7379), .A2(n7378), .A3(n7377), .A4(n7376), .ZN(n8401)
         );
  OAI22_X1 U9122 ( .A1(n8084), .A2(n8423), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9652), .ZN(n7380) );
  AOI21_X1 U9123 ( .B1(n8080), .B2(n8106), .A(n7380), .ZN(n7381) );
  OAI21_X1 U9124 ( .B1(n8431), .B2(n8094), .A(n7381), .ZN(n7382) );
  AOI21_X1 U9125 ( .B1(n8558), .B2(n8101), .A(n7382), .ZN(n7383) );
  OAI21_X1 U9126 ( .B1(n7384), .B2(n8096), .A(n7383), .ZN(P2_U3155) );
  XNOR2_X1 U9127 ( .A(n8701), .B(n8702), .ZN(n7386) );
  NOR2_X1 U9128 ( .A1(n7386), .A2(n7385), .ZN(n8700) );
  AOI21_X1 U9129 ( .B1(n7386), .B2(n7385), .A(n8700), .ZN(n7395) );
  INV_X1 U9130 ( .A(n7387), .ZN(n7391) );
  NOR2_X1 U9131 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7388), .ZN(n9833) );
  AOI21_X1 U9132 ( .B1(n8726), .B2(n10193), .A(n9833), .ZN(n7390) );
  NAND2_X1 U9133 ( .A1(n8693), .A2(n10192), .ZN(n7389) );
  OAI211_X1 U9134 ( .C1(n8696), .C2(n7391), .A(n7390), .B(n7389), .ZN(n7392)
         );
  AOI21_X1 U9135 ( .B1(n7393), .B2(n8731), .A(n7392), .ZN(n7394) );
  OAI21_X1 U9136 ( .B1(n7395), .B2(n8733), .A(n7394), .ZN(P1_U3217) );
  XOR2_X1 U9137 ( .A(n7397), .B(n7396), .Z(n7404) );
  NAND2_X1 U9138 ( .A1(n8693), .A2(n9010), .ZN(n7398) );
  OAI211_X1 U9139 ( .C1(n10216), .C2(n8683), .A(n7399), .B(n7398), .ZN(n7400)
         );
  AOI21_X1 U9140 ( .B1(n8725), .B2(n7401), .A(n7400), .ZN(n7403) );
  NAND2_X1 U9141 ( .A1(n10219), .A2(n8731), .ZN(n7402) );
  OAI211_X1 U9142 ( .C1(n7404), .C2(n8733), .A(n7403), .B(n7402), .ZN(P1_U3224) );
  INV_X1 U9143 ( .A(n8569), .ZN(n7406) );
  OAI222_X1 U9144 ( .A1(P1_U3086), .A2(n5872), .B1(n9820), .B2(n7406), .C1(
        n7405), .C2(n9817), .ZN(P1_U3327) );
  AOI21_X1 U9145 ( .B1(n10101), .B2(n10097), .A(n10090), .ZN(n7414) );
  INV_X1 U9146 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7407) );
  INV_X1 U9147 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9518) );
  OAI22_X1 U9148 ( .A1(n9309), .A2(n7407), .B1(n9518), .B2(n9306), .ZN(n7411)
         );
  NOR4_X1 U9149 ( .A1(n8872), .A2(n4495), .A3(n7409), .A4(n7408), .ZN(n7410)
         );
  AOI211_X1 U9150 ( .C1(n9344), .C2(n6717), .A(n7411), .B(n7410), .ZN(n7412)
         );
  OAI21_X1 U9151 ( .B1(n7414), .B2(n7413), .A(n7412), .ZN(P1_U3293) );
  NAND2_X1 U9152 ( .A1(n7416), .A2(n8425), .ZN(n7772) );
  OR2_X1 U9153 ( .A1(n7416), .A2(n8425), .ZN(n7773) );
  NAND2_X1 U9154 ( .A1(n8558), .A2(n8089), .ZN(n7778) );
  NAND2_X1 U9155 ( .A1(n8428), .A2(n7778), .ZN(n7417) );
  NAND2_X1 U9156 ( .A1(n7417), .A2(n7777), .ZN(n8409) );
  NAND2_X1 U9157 ( .A1(n7418), .A2(n7671), .ZN(n7420) );
  AOI22_X1 U9158 ( .A1(n7456), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7454), .B2(
        n8167), .ZN(n7419) );
  NAND2_X1 U9159 ( .A1(n8552), .A2(n8423), .ZN(n7421) );
  NAND2_X1 U9160 ( .A1(n8409), .A2(n7421), .ZN(n7423) );
  OR2_X1 U9161 ( .A1(n8552), .A2(n8423), .ZN(n7422) );
  NAND2_X1 U9162 ( .A1(n7423), .A2(n7422), .ZN(n8398) );
  NAND2_X1 U9163 ( .A1(n7424), .A2(n7671), .ZN(n7426) );
  AOI22_X1 U9164 ( .A1(n7456), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7454), .B2(
        n8199), .ZN(n7425) );
  NAND2_X1 U9165 ( .A1(n7534), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7432) );
  INV_X1 U9166 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8404) );
  OR2_X1 U9167 ( .A1(n7679), .A2(n8404), .ZN(n7431) );
  NAND2_X1 U9168 ( .A1(n7427), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7428) );
  AND2_X1 U9169 ( .A1(n7437), .A2(n7428), .ZN(n8405) );
  OR2_X1 U9170 ( .A1(n7078), .A2(n8405), .ZN(n7430) );
  INV_X1 U9171 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8478) );
  OR2_X1 U9172 ( .A1(n4494), .A2(n8478), .ZN(n7429) );
  NAND2_X1 U9173 ( .A1(n8546), .A2(n8391), .ZN(n7788) );
  NAND2_X1 U9174 ( .A1(n8398), .A2(n7788), .ZN(n7433) );
  NAND2_X1 U9175 ( .A1(n7433), .A2(n7789), .ZN(n8387) );
  NAND2_X1 U9176 ( .A1(n7434), .A2(n7671), .ZN(n7436) );
  AOI22_X1 U9177 ( .A1(n7456), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7454), .B2(
        n8232), .ZN(n7435) );
  INV_X1 U9178 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8476) );
  OR2_X1 U9179 ( .A1(n4494), .A2(n8476), .ZN(n7442) );
  INV_X1 U9180 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9691) );
  OR2_X1 U9181 ( .A1(n7526), .A2(n9691), .ZN(n7441) );
  NAND2_X1 U9182 ( .A1(n7437), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7438) );
  AND2_X1 U9183 ( .A1(n4496), .A2(n7438), .ZN(n8393) );
  OR2_X1 U9184 ( .A1(n7078), .A2(n8393), .ZN(n7440) );
  INV_X1 U9185 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8394) );
  OR2_X1 U9186 ( .A1(n7679), .A2(n8394), .ZN(n7439) );
  OR2_X1 U9187 ( .A1(n8475), .A2(n8071), .ZN(n7793) );
  NAND2_X1 U9188 ( .A1(n8475), .A2(n8071), .ZN(n7794) );
  NAND2_X1 U9189 ( .A1(n7793), .A2(n7794), .ZN(n8389) );
  NAND2_X1 U9190 ( .A1(n7443), .A2(n7671), .ZN(n7445) );
  AOI22_X1 U9191 ( .A1(n7456), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7454), .B2(
        n8253), .ZN(n7444) );
  NAND2_X1 U9192 ( .A1(n6766), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7452) );
  INV_X1 U9193 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9654) );
  OR2_X1 U9194 ( .A1(n7526), .A2(n9654), .ZN(n7451) );
  INV_X1 U9195 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7446) );
  NAND2_X1 U9196 ( .A1(n4496), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7448) );
  AND2_X1 U9197 ( .A1(n7459), .A2(n7448), .ZN(n7623) );
  OR2_X1 U9198 ( .A1(n7078), .A2(n7623), .ZN(n7450) );
  INV_X1 U9199 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8222) );
  OR2_X1 U9200 ( .A1(n7679), .A2(n8222), .ZN(n7449) );
  NAND4_X1 U9201 ( .A1(n7452), .A2(n7451), .A3(n7450), .A4(n7449), .ZN(n8377)
         );
  NAND2_X1 U9202 ( .A1(n7453), .A2(n7671), .ZN(n7458) );
  AOI22_X1 U9203 ( .A1(n7456), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7455), .B2(
        n7454), .ZN(n7457) );
  NAND2_X1 U9204 ( .A1(n7560), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n7464) );
  INV_X1 U9205 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8471) );
  OR2_X1 U9206 ( .A1(n4494), .A2(n8471), .ZN(n7463) );
  NAND2_X1 U9207 ( .A1(n7459), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n7460) );
  AND2_X1 U9208 ( .A1(n7470), .A2(n7460), .ZN(n7967) );
  OR2_X1 U9209 ( .A1(n7078), .A2(n7967), .ZN(n7462) );
  INV_X1 U9210 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8382) );
  OR2_X1 U9211 ( .A1(n7679), .A2(n8382), .ZN(n7461) );
  NAND2_X1 U9212 ( .A1(n8537), .A2(n7887), .ZN(n7809) );
  INV_X1 U9213 ( .A(n7809), .ZN(n7798) );
  NAND2_X1 U9214 ( .A1(n7465), .A2(n7671), .ZN(n7467) );
  OR2_X1 U9215 ( .A1(n7659), .A2(n9367), .ZN(n7466) );
  NAND2_X1 U9216 ( .A1(n6766), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n7475) );
  INV_X1 U9217 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7468) );
  NAND2_X1 U9218 ( .A1(n7470), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n7471) );
  AND2_X1 U9219 ( .A1(n7480), .A2(n7471), .ZN(n8362) );
  OR2_X1 U9220 ( .A1(n8362), .A2(n7078), .ZN(n7474) );
  INV_X1 U9221 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8532) );
  OR2_X1 U9222 ( .A1(n7526), .A2(n8532), .ZN(n7473) );
  INV_X1 U9223 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8363) );
  OR2_X1 U9224 ( .A1(n7679), .A2(n8363), .ZN(n7472) );
  NAND2_X1 U9225 ( .A1(n8360), .A2(n8345), .ZN(n7808) );
  NAND2_X1 U9226 ( .A1(n7476), .A2(n7671), .ZN(n7479) );
  OR2_X1 U9227 ( .A1(n7659), .A2(n7477), .ZN(n7478) );
  NAND2_X1 U9228 ( .A1(n7480), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n7481) );
  NAND2_X1 U9229 ( .A1(n7494), .A2(n7481), .ZN(n8349) );
  NAND2_X1 U9230 ( .A1(n8349), .A2(n7558), .ZN(n7486) );
  NAND2_X1 U9231 ( .A1(n6766), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n7485) );
  NAND2_X1 U9232 ( .A1(n7560), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7484) );
  INV_X1 U9233 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n7482) );
  OR2_X1 U9234 ( .A1(n7679), .A2(n7482), .ZN(n7483) );
  NAND2_X1 U9235 ( .A1(n7896), .A2(n7897), .ZN(n7814) );
  INV_X1 U9236 ( .A(n7814), .ZN(n7487) );
  NAND2_X1 U9237 ( .A1(n7488), .A2(n7671), .ZN(n7491) );
  OR2_X1 U9238 ( .A1(n7659), .A2(n7489), .ZN(n7490) );
  INV_X1 U9239 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n7492) );
  NAND2_X1 U9240 ( .A1(n7494), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n7495) );
  NAND2_X1 U9241 ( .A1(n7503), .A2(n7495), .ZN(n8340) );
  NAND2_X1 U9242 ( .A1(n8340), .A2(n7558), .ZN(n7498) );
  AOI22_X1 U9243 ( .A1(n6766), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n7560), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n7497) );
  INV_X1 U9244 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8339) );
  OR2_X1 U9245 ( .A1(n7679), .A2(n8339), .ZN(n7496) );
  NAND2_X1 U9246 ( .A1(n8523), .A2(n8346), .ZN(n7819) );
  NAND2_X1 U9247 ( .A1(n7499), .A2(n7671), .ZN(n7502) );
  OR2_X1 U9248 ( .A1(n7659), .A2(n7500), .ZN(n7501) );
  INV_X1 U9249 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8455) );
  NAND2_X1 U9250 ( .A1(n7503), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n7504) );
  NAND2_X1 U9251 ( .A1(n7511), .A2(n7504), .ZN(n8331) );
  NAND2_X1 U9252 ( .A1(n8331), .A2(n7558), .ZN(n7506) );
  AOI22_X1 U9253 ( .A1(n7559), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n7534), .B2(
        P2_REG0_REG_23__SCAN_IN), .ZN(n7505) );
  OAI211_X1 U9254 ( .C1(n4494), .C2(n8455), .A(n7506), .B(n7505), .ZN(n8337)
         );
  INV_X1 U9255 ( .A(n8337), .ZN(n8046) );
  NOR2_X1 U9256 ( .A1(n8517), .A2(n8046), .ZN(n7822) );
  NAND2_X1 U9257 ( .A1(n7507), .A2(n7671), .ZN(n7510) );
  OR2_X1 U9258 ( .A1(n7659), .A2(n7508), .ZN(n7509) );
  NAND2_X1 U9259 ( .A1(n7511), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n7512) );
  NAND2_X1 U9260 ( .A1(n7522), .A2(n7512), .ZN(n8316) );
  INV_X1 U9261 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9690) );
  NAND2_X1 U9262 ( .A1(n7560), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n7514) );
  NAND2_X1 U9263 ( .A1(n7559), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n7513) );
  OAI211_X1 U9264 ( .C1(n4494), .C2(n9690), .A(n7514), .B(n7513), .ZN(n7515)
         );
  NAND2_X1 U9265 ( .A1(n8511), .A2(n8000), .ZN(n7824) );
  NAND2_X1 U9266 ( .A1(n8517), .A2(n8046), .ZN(n8317) );
  AND2_X1 U9267 ( .A1(n7824), .A2(n8317), .ZN(n7826) );
  NAND2_X1 U9268 ( .A1(n7516), .A2(n7671), .ZN(n7519) );
  INV_X1 U9269 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n7520) );
  NAND2_X1 U9270 ( .A1(n7522), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n7523) );
  NAND2_X1 U9271 ( .A1(n7532), .A2(n7523), .ZN(n8302) );
  NAND2_X1 U9272 ( .A1(n8302), .A2(n7558), .ZN(n7529) );
  INV_X1 U9273 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9457) );
  NAND2_X1 U9274 ( .A1(n6766), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n7525) );
  NAND2_X1 U9275 ( .A1(n7559), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n7524) );
  OAI211_X1 U9276 ( .C1(n7526), .C2(n9457), .A(n7525), .B(n7524), .ZN(n7527)
         );
  INV_X1 U9277 ( .A(n7527), .ZN(n7528) );
  NAND2_X1 U9278 ( .A1(n8505), .A2(n7909), .ZN(n7830) );
  NAND2_X1 U9279 ( .A1(n8577), .A2(n7671), .ZN(n7531) );
  OR2_X1 U9280 ( .A1(n7659), .A2(n8579), .ZN(n7530) );
  NAND2_X1 U9281 ( .A1(n7532), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n7533) );
  NAND2_X1 U9282 ( .A1(n7545), .A2(n7533), .ZN(n8292) );
  NAND2_X1 U9283 ( .A1(n8292), .A2(n7558), .ZN(n7539) );
  INV_X1 U9284 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8291) );
  NAND2_X1 U9285 ( .A1(n6766), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n7536) );
  NAND2_X1 U9286 ( .A1(n7534), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n7535) );
  OAI211_X1 U9287 ( .C1(n8291), .C2(n7679), .A(n7536), .B(n7535), .ZN(n7537)
         );
  INV_X1 U9288 ( .A(n7537), .ZN(n7538) );
  INV_X1 U9289 ( .A(n7834), .ZN(n7540) );
  NAND2_X1 U9290 ( .A1(n8500), .A2(n7915), .ZN(n7835) );
  NAND2_X1 U9291 ( .A1(n7541), .A2(n7835), .ZN(n8280) );
  NAND2_X1 U9292 ( .A1(n8572), .A2(n7671), .ZN(n7544) );
  OR2_X1 U9293 ( .A1(n7659), .A2(n7542), .ZN(n7543) );
  NAND2_X1 U9294 ( .A1(n7545), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n7546) );
  INV_X1 U9295 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n7550) );
  NAND2_X1 U9296 ( .A1(n7560), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7549) );
  INV_X1 U9297 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n7547) );
  OR2_X1 U9298 ( .A1(n4494), .A2(n7547), .ZN(n7548) );
  OAI211_X1 U9299 ( .C1(n7550), .C2(n7679), .A(n7549), .B(n7548), .ZN(n7551)
         );
  INV_X1 U9300 ( .A(n7551), .ZN(n7552) );
  NAND2_X1 U9301 ( .A1(n8569), .A2(n7671), .ZN(n7554) );
  OR2_X1 U9302 ( .A1(n7659), .A2(n9496), .ZN(n7553) );
  INV_X1 U9303 ( .A(n7556), .ZN(n7555) );
  INV_X1 U9304 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7924) );
  NAND2_X1 U9305 ( .A1(n7555), .A2(n7924), .ZN(n7935) );
  NAND2_X1 U9306 ( .A1(n7556), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n7557) );
  NAND2_X1 U9307 ( .A1(n7935), .A2(n7557), .ZN(n7923) );
  NAND2_X1 U9308 ( .A1(n7923), .A2(n7558), .ZN(n7565) );
  INV_X1 U9309 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9638) );
  NAND2_X1 U9310 ( .A1(n7559), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n7562) );
  NAND2_X1 U9311 ( .A1(n7560), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7561) );
  OAI211_X1 U9312 ( .C1(n4494), .C2(n9638), .A(n7562), .B(n7561), .ZN(n7563)
         );
  INV_X1 U9313 ( .A(n7563), .ZN(n7564) );
  XNOR2_X1 U9314 ( .A(n7636), .B(n7920), .ZN(n7603) );
  INV_X1 U9315 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n7592) );
  NAND2_X1 U9316 ( .A1(n7567), .A2(n7566), .ZN(n8421) );
  AND2_X1 U9317 ( .A1(n8558), .A2(n8413), .ZN(n7569) );
  OR2_X1 U9318 ( .A1(n8558), .A2(n8413), .ZN(n7568) );
  NAND2_X1 U9319 ( .A1(n8552), .A2(n8401), .ZN(n7690) );
  OR2_X1 U9320 ( .A1(n8552), .A2(n8401), .ZN(n7691) );
  AND2_X1 U9321 ( .A1(n8475), .A2(n8402), .ZN(n7570) );
  NAND2_X1 U9322 ( .A1(n8061), .A2(n8377), .ZN(n7572) );
  NOR2_X1 U9323 ( .A1(n8061), .A2(n8377), .ZN(n7571) );
  AOI21_X1 U9324 ( .B1(n7615), .B2(n7572), .A(n7571), .ZN(n8374) );
  NAND2_X1 U9325 ( .A1(n7803), .A2(n7809), .ZN(n8373) );
  NAND2_X1 U9326 ( .A1(n7811), .A2(n7808), .ZN(n8358) );
  INV_X1 U9327 ( .A(n8360), .ZN(n7574) );
  NAND2_X1 U9328 ( .A1(n7812), .A2(n7814), .ZN(n8348) );
  NOR2_X1 U9329 ( .A1(n8517), .A2(n8337), .ZN(n7579) );
  INV_X1 U9330 ( .A(n8517), .ZN(n7578) );
  NAND2_X1 U9331 ( .A1(n7827), .A2(n7824), .ZN(n8319) );
  NAND2_X1 U9332 ( .A1(n8505), .A2(n8312), .ZN(n7580) );
  INV_X1 U9333 ( .A(n8505), .ZN(n8295) );
  NAND2_X1 U9334 ( .A1(n7913), .A2(n7915), .ZN(n7581) );
  AOI22_X1 U9335 ( .A1(n8288), .A2(n7581), .B1(n8500), .B2(n8298), .ZN(n8277)
         );
  INV_X1 U9336 ( .A(n8277), .ZN(n7583) );
  XOR2_X1 U9337 ( .A(n7920), .B(n7628), .Z(n7591) );
  OR2_X1 U9338 ( .A1(n7935), .A2(n7078), .ZN(n7682) );
  INV_X1 U9339 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n7936) );
  NAND2_X1 U9340 ( .A1(n7534), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7585) );
  NAND2_X1 U9341 ( .A1(n6766), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7584) );
  OAI211_X1 U9342 ( .C1(n7679), .C2(n7936), .A(n7585), .B(n7584), .ZN(n7586)
         );
  INV_X1 U9343 ( .A(n7586), .ZN(n7587) );
  NAND2_X1 U9344 ( .A1(n8289), .A2(n10285), .ZN(n7588) );
  MUX2_X1 U9345 ( .A(n7592), .B(n7599), .S(n10367), .Z(n7594) );
  NAND2_X1 U9346 ( .A1(n7929), .A2(n8559), .ZN(n7593) );
  OAI211_X1 U9347 ( .C1(n7603), .C2(n8555), .A(n7594), .B(n7593), .ZN(P2_U3455) );
  NAND2_X1 U9348 ( .A1(n7929), .A2(n8486), .ZN(n7597) );
  OAI211_X1 U9349 ( .C1(n7603), .C2(n8484), .A(n7598), .B(n7597), .ZN(P2_U3487) );
  INV_X1 U9350 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n7600) );
  MUX2_X1 U9351 ( .A(n7600), .B(n7599), .S(n10299), .Z(n7602) );
  AOI22_X1 U9352 ( .A1(n7929), .A2(n10292), .B1(n10294), .B2(n7923), .ZN(n7601) );
  OAI211_X1 U9353 ( .C1(n7603), .C2(n8420), .A(n7602), .B(n7601), .ZN(P2_U3205) );
  XOR2_X1 U9354 ( .A(n7692), .B(n7604), .Z(n10358) );
  NAND2_X1 U9355 ( .A1(n7605), .A2(n7606), .ZN(n7607) );
  XOR2_X1 U9356 ( .A(n7692), .B(n7607), .Z(n7608) );
  OAI222_X1 U9357 ( .A1(n8424), .A2(n7609), .B1(n8426), .B2(n7982), .C1(n10301), .C2(n7608), .ZN(n10360) );
  NAND2_X1 U9358 ( .A1(n10360), .A2(n10299), .ZN(n7613) );
  OAI22_X1 U9359 ( .A1(n8433), .A2(n7610), .B1(n8057), .B2(n8430), .ZN(n7611)
         );
  AOI21_X1 U9360 ( .B1(n10292), .B2(n8050), .A(n7611), .ZN(n7612) );
  OAI211_X1 U9361 ( .C1(n10358), .C2(n8420), .A(n7613), .B(n7612), .ZN(
        P2_U3222) );
  INV_X1 U9362 ( .A(n8369), .ZN(n7614) );
  NOR2_X1 U9363 ( .A1(n7614), .A2(n8367), .ZN(n7706) );
  XOR2_X1 U9364 ( .A(n7706), .B(n8368), .Z(n7626) );
  XOR2_X1 U9365 ( .A(n7706), .B(n7615), .Z(n7616) );
  AOI222_X1 U9366 ( .A1(n10289), .A2(n7616), .B1(n8356), .B2(n10286), .C1(
        n8402), .C2(n10285), .ZN(n7622) );
  MUX2_X1 U9367 ( .A(n9654), .B(n7622), .S(n10367), .Z(n7618) );
  NAND2_X1 U9368 ( .A1(n8061), .A2(n8559), .ZN(n7617) );
  OAI211_X1 U9369 ( .C1(n7626), .C2(n8555), .A(n7618), .B(n7617), .ZN(P2_U3444) );
  INV_X1 U9370 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7619) );
  MUX2_X1 U9371 ( .A(n7619), .B(n7622), .S(n10386), .Z(n7621) );
  NAND2_X1 U9372 ( .A1(n8061), .A2(n8486), .ZN(n7620) );
  OAI211_X1 U9373 ( .C1(n8484), .C2(n7626), .A(n7621), .B(n7620), .ZN(P2_U3477) );
  MUX2_X1 U9374 ( .A(n8222), .B(n7622), .S(n10299), .Z(n7625) );
  INV_X1 U9375 ( .A(n7623), .ZN(n8073) );
  AOI22_X1 U9376 ( .A1(n8061), .A2(n10292), .B1(n10294), .B2(n8073), .ZN(n7624) );
  OAI211_X1 U9377 ( .C1(n7626), .C2(n8420), .A(n7625), .B(n7624), .ZN(P2_U3215) );
  INV_X1 U9378 ( .A(n8278), .ZN(n7949) );
  INV_X1 U9379 ( .A(n7929), .ZN(n7853) );
  INV_X1 U9380 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7932) );
  INV_X1 U9381 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9811) );
  MUX2_X1 U9382 ( .A(n7932), .B(n9811), .S(n7631), .Z(n7655) );
  NAND2_X1 U9383 ( .A1(n8744), .A2(n7671), .ZN(n7633) );
  OR2_X1 U9384 ( .A1(n7659), .A2(n7932), .ZN(n7632) );
  NAND2_X1 U9385 ( .A1(n7940), .A2(n7634), .ZN(n7684) );
  INV_X1 U9386 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n7639) );
  NAND2_X1 U9387 ( .A1(n6766), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7638) );
  NAND2_X1 U9388 ( .A1(n7534), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7637) );
  OAI211_X1 U9389 ( .C1(n7639), .C2(n7679), .A(n7638), .B(n7637), .ZN(n7640)
         );
  INV_X1 U9390 ( .A(n7640), .ZN(n7641) );
  NAND2_X1 U9391 ( .A1(n7682), .A2(n7641), .ZN(n8104) );
  AND2_X1 U9392 ( .A1(n6476), .A2(P2_B_REG_SCAN_IN), .ZN(n7642) );
  NOR2_X1 U9393 ( .A1(n8424), .A2(n7642), .ZN(n8269) );
  AOI22_X1 U9394 ( .A1(n8278), .A2(n10285), .B1(n8104), .B2(n8269), .ZN(n7643)
         );
  INV_X1 U9395 ( .A(n7940), .ZN(n7652) );
  OR2_X1 U9396 ( .A1(n7652), .A2(n8534), .ZN(n7647) );
  NAND2_X1 U9397 ( .A1(n7648), .A2(n7647), .ZN(P2_U3456) );
  INV_X1 U9398 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7650) );
  NAND2_X1 U9399 ( .A1(n10384), .A2(n7650), .ZN(n7651) );
  OR2_X1 U9400 ( .A1(n7652), .A2(n8470), .ZN(n7653) );
  NAND2_X1 U9401 ( .A1(n7654), .A2(n7653), .ZN(P2_U3488) );
  INV_X1 U9402 ( .A(n7688), .ZN(n7674) );
  NAND2_X1 U9403 ( .A1(n7656), .A2(n7655), .ZN(n7657) );
  INV_X1 U9404 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8740) );
  MUX2_X1 U9405 ( .A(n8740), .B(n7943), .S(n5201), .Z(n7664) );
  XNOR2_X1 U9406 ( .A(n7664), .B(SI_30_), .ZN(n7661) );
  NOR2_X1 U9407 ( .A1(n7659), .A2(n7943), .ZN(n7660) );
  NAND2_X1 U9408 ( .A1(n7662), .A2(n7661), .ZN(n7666) );
  INV_X1 U9409 ( .A(SI_30_), .ZN(n7663) );
  NAND2_X1 U9410 ( .A1(n7664), .A2(n7663), .ZN(n7665) );
  NAND2_X1 U9411 ( .A1(n7666), .A2(n7665), .ZN(n7670) );
  MUX2_X1 U9412 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n5201), .Z(n7668) );
  INV_X1 U9413 ( .A(SI_31_), .ZN(n7667) );
  XNOR2_X1 U9414 ( .A(n7668), .B(n7667), .ZN(n7669) );
  NAND2_X1 U9415 ( .A1(n9807), .A2(n7671), .ZN(n7673) );
  INV_X1 U9416 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8567) );
  OR2_X1 U9417 ( .A1(n7659), .A2(n8567), .ZN(n7672) );
  INV_X1 U9418 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9462) );
  NAND2_X1 U9419 ( .A1(n7534), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7678) );
  INV_X1 U9420 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7676) );
  OR2_X1 U9421 ( .A1(n4494), .A2(n7676), .ZN(n7677) );
  OAI211_X1 U9422 ( .C1(n9462), .C2(n7679), .A(n7678), .B(n7677), .ZN(n7680)
         );
  INV_X1 U9423 ( .A(n7680), .ZN(n7681) );
  OR2_X1 U9424 ( .A1(n8490), .A2(n8103), .ZN(n7859) );
  INV_X1 U9425 ( .A(n8496), .ZN(n8439) );
  INV_X1 U9426 ( .A(n8104), .ZN(n7683) );
  NAND2_X1 U9427 ( .A1(n8439), .A2(n7683), .ZN(n7847) );
  AND2_X1 U9428 ( .A1(n7847), .A2(n7684), .ZN(n7842) );
  NAND2_X1 U9429 ( .A1(n7859), .A2(n7842), .ZN(n7686) );
  INV_X1 U9430 ( .A(n8490), .ZN(n8273) );
  AND2_X1 U9431 ( .A1(n8496), .A2(n8104), .ZN(n7687) );
  NOR2_X1 U9432 ( .A1(n7687), .A2(n8103), .ZN(n7685) );
  INV_X1 U9433 ( .A(n7686), .ZN(n7714) );
  INV_X1 U9434 ( .A(n7687), .ZN(n7849) );
  AND2_X1 U9435 ( .A1(n7849), .A2(n7688), .ZN(n7851) );
  INV_X1 U9436 ( .A(n7920), .ZN(n7712) );
  INV_X1 U9437 ( .A(n8317), .ZN(n7689) );
  OR2_X1 U9438 ( .A1(n7822), .A2(n7689), .ZN(n8325) );
  INV_X1 U9439 ( .A(n8319), .ZN(n8310) );
  INV_X1 U9440 ( .A(n8335), .ZN(n7708) );
  INV_X1 U9441 ( .A(n8373), .ZN(n8371) );
  INV_X1 U9442 ( .A(n8389), .ZN(n8386) );
  NAND2_X1 U9443 ( .A1(n7777), .A2(n7778), .ZN(n8429) );
  AND4_X1 U9444 ( .A1(n7733), .A2(n6746), .A3(n7694), .A4(n10300), .ZN(n7697)
         );
  NAND4_X1 U9445 ( .A1(n7697), .A2(n7696), .A3(n7695), .A4(n10290), .ZN(n7699)
         );
  NOR4_X1 U9446 ( .A1(n4515), .A2(n7700), .A3(n7699), .A4(n7698), .ZN(n7702)
         );
  NAND4_X1 U9447 ( .A1(n7770), .A2(n7703), .A3(n7702), .A4(n7701), .ZN(n7704)
         );
  NOR4_X1 U9448 ( .A1(n4886), .A2(n8411), .A3(n8429), .A4(n7704), .ZN(n7705)
         );
  NAND4_X1 U9449 ( .A1(n8371), .A2(n8386), .A3(n7706), .A4(n7705), .ZN(n7707)
         );
  NOR4_X1 U9450 ( .A1(n7708), .A2(n8348), .A3(n8358), .A4(n7707), .ZN(n7709)
         );
  NAND4_X1 U9451 ( .A1(n8304), .A2(n4758), .A3(n8310), .A4(n7709), .ZN(n7711)
         );
  INV_X1 U9452 ( .A(n7835), .ZN(n7710) );
  NOR4_X1 U9453 ( .A1(n7712), .A2(n8276), .A3(n7711), .A4(n7829), .ZN(n7713)
         );
  NAND2_X1 U9454 ( .A1(n8490), .A2(n8103), .ZN(n7863) );
  NAND4_X1 U9455 ( .A1(n7714), .A2(n7851), .A3(n7713), .A4(n7863), .ZN(n7715)
         );
  NAND2_X1 U9456 ( .A1(n7717), .A2(n7716), .ZN(n7719) );
  NAND2_X1 U9457 ( .A1(n7719), .A2(n7718), .ZN(n7771) );
  INV_X1 U9458 ( .A(n6611), .ZN(n7723) );
  INV_X1 U9459 ( .A(n7720), .ZN(n7728) );
  AOI21_X1 U9460 ( .B1(n7721), .B2(n6468), .A(n7728), .ZN(n7722) );
  OAI211_X1 U9461 ( .C1(n7723), .C2(n7722), .A(n6746), .B(n7726), .ZN(n7725)
         );
  NAND3_X1 U9462 ( .A1(n7725), .A2(n7724), .A3(n7743), .ZN(n7732) );
  INV_X1 U9463 ( .A(n7726), .ZN(n7727) );
  OAI211_X1 U9464 ( .C1(n7728), .C2(n7727), .A(n6746), .B(n6611), .ZN(n7730)
         );
  NAND2_X1 U9465 ( .A1(n8115), .A2(n10315), .ZN(n7735) );
  NAND3_X1 U9466 ( .A1(n7730), .A2(n7735), .A3(n7729), .ZN(n7731) );
  MUX2_X1 U9467 ( .A(n7732), .B(n7731), .S(n7857), .Z(n7734) );
  NAND2_X1 U9468 ( .A1(n7734), .A2(n7733), .ZN(n7747) );
  INV_X1 U9469 ( .A(n7735), .ZN(n7737) );
  OAI211_X1 U9470 ( .C1(n7747), .C2(n7737), .A(n7748), .B(n7736), .ZN(n7738)
         );
  NAND3_X1 U9471 ( .A1(n7738), .A2(n7744), .A3(n7751), .ZN(n7742) );
  NAND2_X1 U9472 ( .A1(n7761), .A2(n7760), .ZN(n7741) );
  NAND2_X1 U9473 ( .A1(n7757), .A2(n7739), .ZN(n7740) );
  MUX2_X1 U9474 ( .A(n7741), .B(n7740), .S(n7857), .Z(n7763) );
  NOR2_X1 U9475 ( .A1(n7763), .A2(n4515), .ZN(n7752) );
  AND3_X1 U9476 ( .A1(n7742), .A2(n7752), .A3(n7749), .ZN(n7755) );
  INV_X1 U9477 ( .A(n7743), .ZN(n7746) );
  OAI211_X1 U9478 ( .C1(n7747), .C2(n7746), .A(n7745), .B(n7744), .ZN(n7750)
         );
  NAND3_X1 U9479 ( .A1(n7750), .A2(n7749), .A3(n7748), .ZN(n7753) );
  AND3_X1 U9480 ( .A1(n7753), .A2(n7752), .A3(n7751), .ZN(n7754) );
  INV_X1 U9481 ( .A(n7756), .ZN(n7766) );
  OAI211_X1 U9482 ( .C1(n7763), .C2(n7758), .A(n7766), .B(n7757), .ZN(n7765)
         );
  AND2_X1 U9483 ( .A1(n7760), .A2(n7759), .ZN(n7762) );
  OAI211_X1 U9484 ( .C1(n7763), .C2(n7762), .A(n7761), .B(n7767), .ZN(n7764)
         );
  MUX2_X1 U9485 ( .A(n7765), .B(n7764), .S(n7857), .Z(n7769) );
  MUX2_X1 U9486 ( .A(n7767), .B(n7766), .S(n7857), .Z(n7768) );
  MUX2_X1 U9487 ( .A(n7773), .B(n7772), .S(n7850), .Z(n7774) );
  OAI21_X1 U9488 ( .B1(n7776), .B2(n7775), .A(n7774), .ZN(n7783) );
  INV_X1 U9489 ( .A(n8429), .ZN(n7782) );
  INV_X1 U9490 ( .A(n7777), .ZN(n7780) );
  INV_X1 U9491 ( .A(n7778), .ZN(n7779) );
  MUX2_X1 U9492 ( .A(n7780), .B(n7779), .S(n7850), .Z(n7781) );
  AOI211_X1 U9493 ( .C1(n7783), .C2(n7782), .A(n8411), .B(n7781), .ZN(n7792)
         );
  NAND2_X1 U9494 ( .A1(n8552), .A2(n7857), .ZN(n7786) );
  INV_X1 U9495 ( .A(n8552), .ZN(n7784) );
  NAND2_X1 U9496 ( .A1(n7784), .A2(n7850), .ZN(n7785) );
  MUX2_X1 U9497 ( .A(n7786), .B(n7785), .S(n8401), .Z(n7787) );
  NAND2_X1 U9498 ( .A1(n8399), .A2(n7787), .ZN(n7791) );
  MUX2_X1 U9499 ( .A(n7789), .B(n7788), .S(n7850), .Z(n7790) );
  OAI211_X1 U9500 ( .C1(n7792), .C2(n7791), .A(n8386), .B(n7790), .ZN(n7800)
         );
  AND2_X1 U9501 ( .A1(n8369), .A2(n7793), .ZN(n7797) );
  INV_X1 U9502 ( .A(n7794), .ZN(n7795) );
  NOR2_X1 U9503 ( .A1(n8367), .A2(n7795), .ZN(n7796) );
  MUX2_X1 U9504 ( .A(n7797), .B(n7796), .S(n7857), .Z(n7799) );
  AOI21_X1 U9505 ( .B1(n7800), .B2(n7799), .A(n7798), .ZN(n7806) );
  INV_X1 U9506 ( .A(n8367), .ZN(n7801) );
  MUX2_X1 U9507 ( .A(n7802), .B(n7801), .S(n7850), .Z(n7805) );
  AOI21_X1 U9508 ( .B1(n7811), .B2(n7803), .A(n7857), .ZN(n7804) );
  AOI21_X1 U9509 ( .B1(n7806), .B2(n7805), .A(n7804), .ZN(n7810) );
  NAND2_X1 U9510 ( .A1(n7814), .A2(n7808), .ZN(n7807) );
  OAI21_X1 U9511 ( .B1(n7810), .B2(n7807), .A(n7812), .ZN(n7817) );
  NAND3_X1 U9512 ( .A1(n7810), .A2(n7809), .A3(n7808), .ZN(n7813) );
  NAND3_X1 U9513 ( .A1(n7813), .A2(n7812), .A3(n7811), .ZN(n7815) );
  NAND2_X1 U9514 ( .A1(n7815), .A2(n7814), .ZN(n7816) );
  MUX2_X1 U9515 ( .A(n7817), .B(n7816), .S(n7857), .Z(n7818) );
  MUX2_X1 U9516 ( .A(n7820), .B(n7819), .S(n7857), .Z(n7821) );
  INV_X1 U9517 ( .A(n7822), .ZN(n7823) );
  NAND2_X1 U9518 ( .A1(n7827), .A2(n7823), .ZN(n7825) );
  INV_X1 U9519 ( .A(n7826), .ZN(n7828) );
  MUX2_X1 U9520 ( .A(n7831), .B(n7830), .S(n7857), .Z(n7832) );
  OAI211_X1 U9521 ( .C1(n7833), .C2(n8296), .A(n8287), .B(n7832), .ZN(n7837)
         );
  MUX2_X1 U9522 ( .A(n7835), .B(n7540), .S(n7857), .Z(n7836) );
  NAND3_X1 U9523 ( .A1(n7837), .A2(n4920), .A3(n7836), .ZN(n7841) );
  NAND2_X1 U9524 ( .A1(n8443), .A2(n8085), .ZN(n7838) );
  MUX2_X1 U9525 ( .A(n7839), .B(n7838), .S(n7857), .Z(n7840) );
  NAND2_X1 U9526 ( .A1(n7841), .A2(n7840), .ZN(n7845) );
  MUX2_X1 U9527 ( .A(n7949), .B(n7853), .S(n7850), .Z(n7844) );
  AOI21_X1 U9528 ( .B1(n7845), .B2(n7844), .A(n7843), .ZN(n7854) );
  INV_X1 U9529 ( .A(n7842), .ZN(n7846) );
  NOR3_X1 U9530 ( .A1(n7845), .A2(n7844), .A3(n7843), .ZN(n7855) );
  AOI211_X1 U9531 ( .C1(n7854), .C2(n7949), .A(n7846), .B(n7855), .ZN(n7862)
         );
  INV_X1 U9532 ( .A(n7847), .ZN(n7848) );
  AOI21_X1 U9533 ( .B1(n7850), .B2(n7849), .A(n7848), .ZN(n7861) );
  INV_X1 U9534 ( .A(n7851), .ZN(n7852) );
  AOI21_X1 U9535 ( .B1(n7854), .B2(n7853), .A(n7852), .ZN(n7858) );
  INV_X1 U9536 ( .A(n7855), .ZN(n7856) );
  NAND3_X1 U9537 ( .A1(n7858), .A2(n7857), .A3(n7856), .ZN(n7860) );
  OAI211_X1 U9538 ( .C1(n7862), .C2(n7861), .A(n7860), .B(n7859), .ZN(n7864)
         );
  NAND2_X1 U9539 ( .A1(n7864), .A2(n7863), .ZN(n7866) );
  XNOR2_X1 U9540 ( .A(n7868), .B(n7455), .ZN(n7875) );
  NAND3_X1 U9541 ( .A1(n7870), .A2(n7869), .A3(n8255), .ZN(n7871) );
  OAI211_X1 U9542 ( .C1(n7872), .C2(n7874), .A(n7871), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7873) );
  OAI21_X1 U9543 ( .B1(n7875), .B2(n7874), .A(n7873), .ZN(P2_U3296) );
  INV_X1 U9544 ( .A(n7876), .ZN(n7877) );
  XNOR2_X1 U9545 ( .A(n8552), .B(n7900), .ZN(n7880) );
  XNOR2_X1 U9546 ( .A(n7880), .B(n8423), .ZN(n8098) );
  NOR2_X1 U9547 ( .A1(n7880), .A2(n8423), .ZN(n7881) );
  NOR2_X2 U9548 ( .A1(n8095), .A2(n7881), .ZN(n8006) );
  XNOR2_X1 U9549 ( .A(n8546), .B(n7900), .ZN(n8004) );
  XNOR2_X1 U9550 ( .A(n8475), .B(n6486), .ZN(n7882) );
  NOR2_X1 U9551 ( .A1(n7882), .A2(n8402), .ZN(n8064) );
  AOI21_X1 U9552 ( .B1(n7882), .B2(n8402), .A(n8064), .ZN(n8014) );
  XNOR2_X1 U9553 ( .A(n8061), .B(n7900), .ZN(n7883) );
  NAND2_X1 U9554 ( .A1(n7883), .A2(n8392), .ZN(n7961) );
  INV_X1 U9555 ( .A(n7883), .ZN(n7884) );
  NAND2_X1 U9556 ( .A1(n7884), .A2(n8377), .ZN(n7885) );
  AND2_X1 U9557 ( .A1(n7961), .A2(n7885), .ZN(n8063) );
  NAND2_X1 U9558 ( .A1(n7886), .A2(n8063), .ZN(n7960) );
  NAND2_X1 U9559 ( .A1(n7960), .A2(n7961), .ZN(n7891) );
  XNOR2_X1 U9560 ( .A(n8537), .B(n7900), .ZN(n7888) );
  NAND2_X1 U9561 ( .A1(n7888), .A2(n7887), .ZN(n8029) );
  INV_X1 U9562 ( .A(n7888), .ZN(n7889) );
  NAND2_X1 U9563 ( .A1(n7889), .A2(n8356), .ZN(n7890) );
  NAND2_X1 U9564 ( .A1(n7891), .A2(n7962), .ZN(n7964) );
  XNOR2_X1 U9565 ( .A(n8360), .B(n7900), .ZN(n7892) );
  NAND2_X1 U9566 ( .A1(n7892), .A2(n8345), .ZN(n7974) );
  INV_X1 U9567 ( .A(n7892), .ZN(n7893) );
  NAND2_X1 U9568 ( .A1(n7893), .A2(n8378), .ZN(n7894) );
  AND2_X1 U9569 ( .A1(n7974), .A2(n7894), .ZN(n8031) );
  XNOR2_X1 U9570 ( .A(n7896), .B(n6486), .ZN(n7898) );
  XNOR2_X1 U9571 ( .A(n7898), .B(n7897), .ZN(n7975) );
  XNOR2_X1 U9572 ( .A(n8523), .B(n6486), .ZN(n7899) );
  NOR2_X1 U9573 ( .A1(n7899), .A2(n8327), .ZN(n8039) );
  NAND2_X1 U9574 ( .A1(n7899), .A2(n8327), .ZN(n8040) );
  XNOR2_X1 U9575 ( .A(n8517), .B(n7900), .ZN(n7901) );
  NAND2_X1 U9576 ( .A1(n7953), .A2(n8046), .ZN(n7905) );
  INV_X1 U9577 ( .A(n7901), .ZN(n7902) );
  OR2_X1 U9578 ( .A1(n7903), .A2(n7902), .ZN(n7904) );
  NAND2_X1 U9579 ( .A1(n7905), .A2(n7904), .ZN(n8022) );
  XNOR2_X1 U9580 ( .A(n8511), .B(n7900), .ZN(n7906) );
  XNOR2_X1 U9581 ( .A(n7906), .B(n8328), .ZN(n8023) );
  NAND2_X1 U9582 ( .A1(n8022), .A2(n8023), .ZN(n7908) );
  NAND2_X1 U9583 ( .A1(n7906), .A2(n8000), .ZN(n7907) );
  XNOR2_X1 U9584 ( .A(n8505), .B(n6644), .ZN(n7910) );
  XNOR2_X1 U9585 ( .A(n7910), .B(n8312), .ZN(n7997) );
  NAND2_X1 U9586 ( .A1(n7996), .A2(n7997), .ZN(n7912) );
  NAND2_X1 U9587 ( .A1(n7910), .A2(n7909), .ZN(n7911) );
  XNOR2_X1 U9588 ( .A(n7913), .B(n7900), .ZN(n7914) );
  XNOR2_X1 U9589 ( .A(n7914), .B(n7915), .ZN(n8079) );
  INV_X1 U9590 ( .A(n7914), .ZN(n7916) );
  NAND2_X1 U9591 ( .A1(n7916), .A2(n7915), .ZN(n7917) );
  XNOR2_X1 U9592 ( .A(n8283), .B(n7900), .ZN(n7918) );
  NAND2_X1 U9593 ( .A1(n7918), .A2(n8289), .ZN(n7919) );
  OAI21_X1 U9594 ( .B1(n7918), .B2(n8289), .A(n7919), .ZN(n7945) );
  XNOR2_X1 U9595 ( .A(n7920), .B(n6644), .ZN(n7921) );
  XNOR2_X1 U9596 ( .A(n7922), .B(n7921), .ZN(n7931) );
  INV_X1 U9597 ( .A(n7923), .ZN(n7927) );
  OAI22_X1 U9598 ( .A1(n8085), .A2(n8090), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7924), .ZN(n7925) );
  AOI21_X1 U9599 ( .B1(n8105), .B2(n8092), .A(n7925), .ZN(n7926) );
  OAI21_X1 U9600 ( .B1(n7927), .B2(n8094), .A(n7926), .ZN(n7928) );
  AOI21_X1 U9601 ( .B1(n7929), .B2(n8101), .A(n7928), .ZN(n7930) );
  OAI21_X1 U9602 ( .B1(n7931), .B2(n8096), .A(n7930), .ZN(P2_U3160) );
  INV_X1 U9603 ( .A(n8744), .ZN(n9812) );
  OAI222_X1 U9604 ( .A1(n8576), .A2(n9812), .B1(n7933), .B2(P2_U3151), .C1(
        n7932), .C2(n8578), .ZN(P2_U3266) );
  INV_X1 U9605 ( .A(n8739), .ZN(n7944) );
  OAI222_X1 U9606 ( .A1(P1_U3086), .A2(n5149), .B1(n9820), .B2(n7944), .C1(
        n8740), .C2(n9817), .ZN(P1_U3325) );
  OR2_X1 U9607 ( .A1(n7935), .A2(n8430), .ZN(n8271) );
  OAI21_X1 U9608 ( .B1(n10299), .B2(n7936), .A(n8271), .ZN(n7939) );
  NOR2_X1 U9609 ( .A1(n7645), .A2(n7937), .ZN(n7938) );
  AOI211_X1 U9610 ( .C1(n10292), .C2(n7940), .A(n7939), .B(n7938), .ZN(n7941)
         );
  OAI21_X1 U9611 ( .B1(n7934), .B2(n8381), .A(n7941), .ZN(P2_U3204) );
  OAI222_X1 U9612 ( .A1(n8576), .A2(n7944), .B1(n8578), .B2(n7943), .C1(
        P2_U3151), .C2(n7942), .ZN(P2_U3265) );
  AOI22_X1 U9613 ( .A1(n8298), .A2(n8080), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7948) );
  OAI21_X1 U9614 ( .B1(n7949), .B2(n8084), .A(n7948), .ZN(n7950) );
  AOI21_X1 U9615 ( .B1(n8281), .B2(n8081), .A(n7950), .ZN(n7951) );
  OAI211_X1 U9616 ( .C1(n8283), .C2(n8076), .A(n7952), .B(n7951), .ZN(P2_U3154) );
  XNOR2_X1 U9617 ( .A(n7953), .B(n8337), .ZN(n7959) );
  INV_X1 U9618 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7954) );
  OAI22_X1 U9619 ( .A1(n8090), .A2(n8346), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7954), .ZN(n7956) );
  NOR2_X1 U9620 ( .A1(n8084), .A2(n8000), .ZN(n7955) );
  AOI211_X1 U9621 ( .C1(n8331), .C2(n8081), .A(n7956), .B(n7955), .ZN(n7958)
         );
  NAND2_X1 U9622 ( .A1(n8517), .A2(n8101), .ZN(n7957) );
  OAI211_X1 U9623 ( .C1(n7959), .C2(n8096), .A(n7958), .B(n7957), .ZN(P2_U3156) );
  INV_X1 U9624 ( .A(n8537), .ZN(n7972) );
  INV_X1 U9625 ( .A(n7960), .ZN(n8067) );
  INV_X1 U9626 ( .A(n7961), .ZN(n7963) );
  NOR3_X1 U9627 ( .A1(n8067), .A2(n7963), .A3(n7962), .ZN(n7966) );
  INV_X1 U9628 ( .A(n7964), .ZN(n7965) );
  OAI21_X1 U9629 ( .B1(n7966), .B2(n7965), .A(n8066), .ZN(n7971) );
  INV_X1 U9630 ( .A(n7967), .ZN(n8383) );
  NAND2_X1 U9631 ( .A1(n8092), .A2(n8378), .ZN(n7968) );
  NAND2_X1 U9632 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8260) );
  OAI211_X1 U9633 ( .C1(n8392), .C2(n8090), .A(n7968), .B(n8260), .ZN(n7969)
         );
  AOI21_X1 U9634 ( .B1(n8383), .B2(n8081), .A(n7969), .ZN(n7970) );
  OAI211_X1 U9635 ( .C1(n7972), .C2(n8076), .A(n7971), .B(n7970), .ZN(P2_U3159) );
  INV_X1 U9636 ( .A(n7973), .ZN(n8032) );
  NOR3_X1 U9637 ( .A1(n8032), .A2(n5024), .A3(n7975), .ZN(n7976) );
  OAI21_X1 U9638 ( .B1(n7976), .B2(n5022), .A(n8066), .ZN(n7980) );
  AOI22_X1 U9639 ( .A1(n8080), .A2(n8378), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n7977) );
  OAI21_X1 U9640 ( .B1(n8346), .B2(n8084), .A(n7977), .ZN(n7978) );
  AOI21_X1 U9641 ( .B1(n8081), .B2(n8349), .A(n7978), .ZN(n7979) );
  OAI211_X1 U9642 ( .C1(n8530), .C2(n8076), .A(n7980), .B(n7979), .ZN(P2_U3163) );
  AOI21_X1 U9643 ( .B1(n7983), .B2(n7982), .A(n7981), .ZN(n8053) );
  XNOR2_X1 U9644 ( .A(n7984), .B(n7988), .ZN(n8052) );
  NAND2_X1 U9645 ( .A1(n8053), .A2(n8052), .ZN(n8051) );
  NAND2_X1 U9646 ( .A1(n8051), .A2(n7985), .ZN(n7986) );
  XOR2_X1 U9647 ( .A(n7987), .B(n7986), .Z(n7995) );
  NOR2_X1 U9648 ( .A1(n8090), .A2(n7988), .ZN(n7989) );
  AOI211_X1 U9649 ( .C1(n8092), .C2(n8106), .A(n7990), .B(n7989), .ZN(n7991)
         );
  OAI21_X1 U9650 ( .B1(n7992), .B2(n8094), .A(n7991), .ZN(n7993) );
  AOI21_X1 U9651 ( .B1(n10365), .B2(n8101), .A(n7993), .ZN(n7994) );
  OAI21_X1 U9652 ( .B1(n7995), .B2(n8096), .A(n7994), .ZN(P2_U3164) );
  XOR2_X1 U9653 ( .A(n7997), .B(n7996), .Z(n8003) );
  AOI22_X1 U9654 ( .A1(n8298), .A2(n8092), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n7999) );
  NAND2_X1 U9655 ( .A1(n8081), .A2(n8302), .ZN(n7998) );
  OAI211_X1 U9656 ( .C1(n8000), .C2(n8090), .A(n7999), .B(n7998), .ZN(n8001)
         );
  AOI21_X1 U9657 ( .B1(n8505), .B2(n8101), .A(n8001), .ZN(n8002) );
  OAI21_X1 U9658 ( .B1(n8003), .B2(n8096), .A(n8002), .ZN(P2_U3165) );
  XNOR2_X1 U9659 ( .A(n8004), .B(n8391), .ZN(n8005) );
  XNOR2_X1 U9660 ( .A(n8006), .B(n8005), .ZN(n8012) );
  NOR2_X1 U9661 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8007), .ZN(n8187) );
  NOR2_X1 U9662 ( .A1(n8090), .A2(n8423), .ZN(n8008) );
  AOI211_X1 U9663 ( .C1(n8092), .C2(n8402), .A(n8187), .B(n8008), .ZN(n8009)
         );
  OAI21_X1 U9664 ( .B1(n8405), .B2(n8094), .A(n8009), .ZN(n8010) );
  AOI21_X1 U9665 ( .B1(n8546), .B2(n8101), .A(n8010), .ZN(n8011) );
  OAI21_X1 U9666 ( .B1(n8012), .B2(n8096), .A(n8011), .ZN(P2_U3166) );
  INV_X1 U9667 ( .A(n8475), .ZN(n8021) );
  OAI21_X1 U9668 ( .B1(n8014), .B2(n8013), .A(n8062), .ZN(n8015) );
  NAND2_X1 U9669 ( .A1(n8015), .A2(n8066), .ZN(n8020) );
  INV_X1 U9670 ( .A(n8393), .ZN(n8018) );
  AND2_X1 U9671 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8201) );
  AOI21_X1 U9672 ( .B1(n8092), .B2(n8377), .A(n8201), .ZN(n8016) );
  OAI21_X1 U9673 ( .B1(n8391), .B2(n8090), .A(n8016), .ZN(n8017) );
  AOI21_X1 U9674 ( .B1(n8018), .B2(n8081), .A(n8017), .ZN(n8019) );
  OAI211_X1 U9675 ( .C1(n8021), .C2(n8076), .A(n8020), .B(n8019), .ZN(P2_U3168) );
  XOR2_X1 U9676 ( .A(n8023), .B(n8022), .Z(n8028) );
  AOI22_X1 U9677 ( .A1(n8312), .A2(n8092), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8025) );
  NAND2_X1 U9678 ( .A1(n8081), .A2(n8316), .ZN(n8024) );
  OAI211_X1 U9679 ( .C1(n8046), .C2(n8090), .A(n8025), .B(n8024), .ZN(n8026)
         );
  AOI21_X1 U9680 ( .B1(n8511), .B2(n8101), .A(n8026), .ZN(n8027) );
  OAI21_X1 U9681 ( .B1(n8028), .B2(n8096), .A(n8027), .ZN(P2_U3169) );
  INV_X1 U9682 ( .A(n8029), .ZN(n8030) );
  NOR2_X1 U9683 ( .A1(n8031), .A2(n8030), .ZN(n8033) );
  AOI21_X1 U9684 ( .B1(n8033), .B2(n7964), .A(n8032), .ZN(n8038) );
  AOI22_X1 U9685 ( .A1(n8092), .A2(n7576), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8035) );
  NAND2_X1 U9686 ( .A1(n8080), .A2(n8356), .ZN(n8034) );
  OAI211_X1 U9687 ( .C1(n8362), .C2(n8094), .A(n8035), .B(n8034), .ZN(n8036)
         );
  AOI21_X1 U9688 ( .B1(n8360), .B2(n8101), .A(n8036), .ZN(n8037) );
  OAI21_X1 U9689 ( .B1(n8038), .B2(n8096), .A(n8037), .ZN(P2_U3173) );
  INV_X1 U9690 ( .A(n8039), .ZN(n8041) );
  NAND2_X1 U9691 ( .A1(n8041), .A2(n8040), .ZN(n8042) );
  XNOR2_X1 U9692 ( .A(n8043), .B(n8042), .ZN(n8049) );
  NAND2_X1 U9693 ( .A1(n8081), .A2(n8340), .ZN(n8045) );
  AOI22_X1 U9694 ( .A1(n8080), .A2(n7576), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8044) );
  OAI211_X1 U9695 ( .C1(n8046), .C2(n8084), .A(n8045), .B(n8044), .ZN(n8047)
         );
  AOI21_X1 U9696 ( .B1(n8523), .B2(n8101), .A(n8047), .ZN(n8048) );
  OAI21_X1 U9697 ( .B1(n8049), .B2(n8096), .A(n8048), .ZN(P2_U3175) );
  INV_X1 U9698 ( .A(n8050), .ZN(n10357) );
  OAI211_X1 U9699 ( .C1(n8053), .C2(n8052), .A(n8051), .B(n8066), .ZN(n8060)
         );
  AOI21_X1 U9700 ( .B1(n8080), .B2(n8109), .A(n8054), .ZN(n8056) );
  NAND2_X1 U9701 ( .A1(n8092), .A2(n8107), .ZN(n8055) );
  OAI211_X1 U9702 ( .C1(n8057), .C2(n8094), .A(n8056), .B(n8055), .ZN(n8058)
         );
  INV_X1 U9703 ( .A(n8058), .ZN(n8059) );
  OAI211_X1 U9704 ( .C1(n10357), .C2(n8076), .A(n8060), .B(n8059), .ZN(
        P2_U3176) );
  INV_X1 U9705 ( .A(n8061), .ZN(n8077) );
  INV_X1 U9706 ( .A(n8062), .ZN(n8065) );
  NOR3_X1 U9707 ( .A1(n8065), .A2(n8064), .A3(n8063), .ZN(n8068) );
  OAI21_X1 U9708 ( .B1(n8068), .B2(n8067), .A(n8066), .ZN(n8075) );
  NAND2_X1 U9709 ( .A1(n8092), .A2(n8356), .ZN(n8070) );
  AND2_X1 U9710 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8242) );
  INV_X1 U9711 ( .A(n8242), .ZN(n8069) );
  OAI211_X1 U9712 ( .C1(n8071), .C2(n8090), .A(n8070), .B(n8069), .ZN(n8072)
         );
  AOI21_X1 U9713 ( .B1(n8073), .B2(n8081), .A(n8072), .ZN(n8074) );
  OAI211_X1 U9714 ( .C1(n8077), .C2(n8076), .A(n8075), .B(n8074), .ZN(P2_U3178) );
  XOR2_X1 U9715 ( .A(n8079), .B(n8078), .Z(n8088) );
  AOI22_X1 U9716 ( .A1(n8312), .A2(n8080), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8083) );
  NAND2_X1 U9717 ( .A1(n8081), .A2(n8292), .ZN(n8082) );
  OAI211_X1 U9718 ( .C1(n8085), .C2(n8084), .A(n8083), .B(n8082), .ZN(n8086)
         );
  AOI21_X1 U9719 ( .B1(n8500), .B2(n8101), .A(n8086), .ZN(n8087) );
  OAI21_X1 U9720 ( .B1(n8088), .B2(n8096), .A(n8087), .ZN(P2_U3180) );
  AND2_X1 U9721 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8150) );
  NOR2_X1 U9722 ( .A1(n8090), .A2(n8089), .ZN(n8091) );
  AOI211_X1 U9723 ( .C1(n8092), .C2(n8412), .A(n8150), .B(n8091), .ZN(n8093)
         );
  OAI21_X1 U9724 ( .B1(n8416), .B2(n8094), .A(n8093), .ZN(n8100) );
  AOI211_X1 U9725 ( .C1(n8098), .C2(n8097), .A(n8096), .B(n8095), .ZN(n8099)
         );
  AOI211_X1 U9726 ( .C1(n8552), .C2(n8101), .A(n8100), .B(n8099), .ZN(n8102)
         );
  INV_X1 U9727 ( .A(n8102), .ZN(P2_U3181) );
  MUX2_X1 U9728 ( .A(n8270), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8236), .Z(
        P2_U3522) );
  MUX2_X1 U9729 ( .A(n8104), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8236), .Z(
        P2_U3521) );
  MUX2_X1 U9730 ( .A(n8105), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8236), .Z(
        P2_U3520) );
  MUX2_X1 U9731 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8278), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9732 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8289), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9733 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8298), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9734 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8312), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9735 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8328), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9736 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8337), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U9737 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8327), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9738 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n7576), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9739 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8378), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9740 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8356), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9741 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8377), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9742 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8402), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9743 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8412), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9744 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8401), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9745 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8413), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9746 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8106), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U9747 ( .A(n8107), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8236), .Z(
        P2_U3503) );
  MUX2_X1 U9748 ( .A(n8108), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8236), .Z(
        P2_U3502) );
  MUX2_X1 U9749 ( .A(n8109), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8236), .Z(
        P2_U3501) );
  MUX2_X1 U9750 ( .A(n8110), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8236), .Z(
        P2_U3500) );
  MUX2_X1 U9751 ( .A(n8111), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8236), .Z(
        P2_U3499) );
  MUX2_X1 U9752 ( .A(n8112), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8236), .Z(
        P2_U3498) );
  MUX2_X1 U9753 ( .A(n8113), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8236), .Z(
        P2_U3497) );
  MUX2_X1 U9754 ( .A(n8114), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8236), .Z(
        P2_U3496) );
  MUX2_X1 U9755 ( .A(n10287), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8236), .Z(
        P2_U3495) );
  MUX2_X1 U9756 ( .A(n8115), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8236), .Z(
        P2_U3494) );
  MUX2_X1 U9757 ( .A(n4512), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8236), .Z(
        P2_U3493) );
  MUX2_X1 U9758 ( .A(n8116), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8236), .Z(
        P2_U3492) );
  MUX2_X1 U9759 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n6536), .S(P2_U3893), .Z(
        P2_U3491) );
  INV_X1 U9760 ( .A(n8117), .ZN(n8119) );
  NAND2_X1 U9761 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8145), .ZN(n8120) );
  OAI21_X1 U9762 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8145), .A(n8120), .ZN(
        n8121) );
  AOI21_X1 U9763 ( .B1(n4532), .B2(n8121), .A(n8144), .ZN(n8143) );
  AOI22_X1 U9764 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8145), .B1(n8148), .B2(
        n9471), .ZN(n8127) );
  NAND2_X1 U9765 ( .A1(n8123), .A2(n8122), .ZN(n8125) );
  NAND2_X1 U9766 ( .A1(n8125), .A2(n8124), .ZN(n8126) );
  NAND2_X1 U9767 ( .A1(n8127), .A2(n8126), .ZN(n8147) );
  OAI21_X1 U9768 ( .B1(n8127), .B2(n8126), .A(n8147), .ZN(n8131) );
  NOR2_X1 U9769 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9652), .ZN(n8128) );
  AOI21_X1 U9770 ( .B1(n8202), .B2(n8148), .A(n8128), .ZN(n8129) );
  OAI21_X1 U9771 ( .B1(n9357), .B2(n8204), .A(n8129), .ZN(n8130) );
  AOI21_X1 U9772 ( .B1(n8131), .B2(n8267), .A(n8130), .ZN(n8142) );
  INV_X1 U9773 ( .A(n8132), .ZN(n8137) );
  MUX2_X1 U9774 ( .A(n8432), .B(n9471), .S(n8255), .Z(n8133) );
  NAND2_X1 U9775 ( .A1(n8133), .A2(n8148), .ZN(n8157) );
  INV_X1 U9776 ( .A(n8133), .ZN(n8134) );
  NAND2_X1 U9777 ( .A1(n8134), .A2(n8145), .ZN(n8135) );
  AND2_X1 U9778 ( .A1(n8157), .A2(n8135), .ZN(n8136) );
  OAI21_X1 U9779 ( .B1(n8138), .B2(n8137), .A(n8136), .ZN(n8158) );
  INV_X1 U9780 ( .A(n8158), .ZN(n8140) );
  NOR3_X1 U9781 ( .A1(n8138), .A2(n8137), .A3(n8136), .ZN(n8139) );
  OAI21_X1 U9782 ( .B1(n8140), .B2(n8139), .A(n10279), .ZN(n8141) );
  OAI211_X1 U9783 ( .C1(n8143), .C2(n8268), .A(n8142), .B(n8141), .ZN(P2_U3196) );
  XNOR2_X1 U9784 ( .A(n8167), .B(n8166), .ZN(n8146) );
  AOI21_X1 U9785 ( .B1(n8415), .B2(n8146), .A(n8169), .ZN(n8165) );
  OAI21_X1 U9786 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n8149), .A(n8174), .ZN(
        n8163) );
  INV_X1 U9787 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8152) );
  AOI21_X1 U9788 ( .B1(n8202), .B2(n8167), .A(n8150), .ZN(n8151) );
  OAI21_X1 U9789 ( .B1(n8152), .B2(n8204), .A(n8151), .ZN(n8162) );
  MUX2_X1 U9790 ( .A(n8415), .B(n8481), .S(n8255), .Z(n8153) );
  NAND2_X1 U9791 ( .A1(n8153), .A2(n8167), .ZN(n8178) );
  INV_X1 U9792 ( .A(n8153), .ZN(n8154) );
  NAND2_X1 U9793 ( .A1(n8154), .A2(n8173), .ZN(n8155) );
  NAND2_X1 U9794 ( .A1(n8178), .A2(n8155), .ZN(n8156) );
  AOI21_X1 U9795 ( .B1(n8158), .B2(n8157), .A(n8156), .ZN(n8184) );
  INV_X1 U9796 ( .A(n8184), .ZN(n8160) );
  NAND3_X1 U9797 ( .A1(n8158), .A2(n8157), .A3(n8156), .ZN(n8159) );
  AOI21_X1 U9798 ( .B1(n8160), .B2(n8159), .A(n8264), .ZN(n8161) );
  AOI211_X1 U9799 ( .C1(n8163), .C2(n8267), .A(n8162), .B(n8161), .ZN(n8164)
         );
  OAI21_X1 U9800 ( .B1(n8165), .B2(n8268), .A(n8164), .ZN(P2_U3197) );
  NOR2_X1 U9801 ( .A1(n8167), .A2(n8166), .ZN(n8168) );
  NAND2_X1 U9802 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8195), .ZN(n8170) );
  OAI21_X1 U9803 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8195), .A(n8170), .ZN(
        n8171) );
  AOI21_X1 U9804 ( .B1(n4576), .B2(n8171), .A(n8196), .ZN(n8194) );
  AOI22_X1 U9805 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8195), .B1(n8199), .B2(
        n8478), .ZN(n8177) );
  NAND2_X1 U9806 ( .A1(n8173), .A2(n8172), .ZN(n8175) );
  NAND2_X1 U9807 ( .A1(n8177), .A2(n8176), .ZN(n8198) );
  OAI21_X1 U9808 ( .B1(n8177), .B2(n8176), .A(n8198), .ZN(n8192) );
  INV_X1 U9809 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8190) );
  INV_X1 U9810 ( .A(n8178), .ZN(n8183) );
  MUX2_X1 U9811 ( .A(n8404), .B(n8478), .S(n8255), .Z(n8179) );
  NAND2_X1 U9812 ( .A1(n8179), .A2(n8199), .ZN(n8206) );
  INV_X1 U9813 ( .A(n8179), .ZN(n8180) );
  NAND2_X1 U9814 ( .A1(n8180), .A2(n8195), .ZN(n8181) );
  AND2_X1 U9815 ( .A1(n8206), .A2(n8181), .ZN(n8182) );
  OAI21_X1 U9816 ( .B1(n8184), .B2(n8183), .A(n8182), .ZN(n8208) );
  INV_X1 U9817 ( .A(n8208), .ZN(n8186) );
  NOR3_X1 U9818 ( .A1(n8184), .A2(n8183), .A3(n8182), .ZN(n8185) );
  OAI21_X1 U9819 ( .B1(n8186), .B2(n8185), .A(n10279), .ZN(n8189) );
  AOI21_X1 U9820 ( .B1(n8202), .B2(n8199), .A(n8187), .ZN(n8188) );
  OAI211_X1 U9821 ( .C1(n8190), .C2(n8204), .A(n8189), .B(n8188), .ZN(n8191)
         );
  AOI21_X1 U9822 ( .B1(n8267), .B2(n8192), .A(n8191), .ZN(n8193) );
  OAI21_X1 U9823 ( .B1(n8194), .B2(n8268), .A(n8193), .ZN(P2_U3198) );
  NOR2_X1 U9824 ( .A1(n8394), .A2(n8197), .ZN(n8220) );
  AOI21_X1 U9825 ( .B1(n8394), .B2(n8197), .A(n8220), .ZN(n8215) );
  OAI21_X1 U9826 ( .B1(n8199), .B2(n8478), .A(n8198), .ZN(n8216) );
  XNOR2_X1 U9827 ( .A(n8216), .B(n8232), .ZN(n8200) );
  NAND2_X1 U9828 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n8200), .ZN(n8218) );
  OAI21_X1 U9829 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8200), .A(n8218), .ZN(
        n8213) );
  INV_X1 U9830 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8205) );
  AOI21_X1 U9831 ( .B1(n8202), .B2(n8232), .A(n8201), .ZN(n8203) );
  OAI21_X1 U9832 ( .B1(n8205), .B2(n8204), .A(n8203), .ZN(n8212) );
  MUX2_X1 U9833 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8255), .Z(n8229) );
  XNOR2_X1 U9834 ( .A(n8229), .B(n8217), .ZN(n8207) );
  AOI21_X1 U9835 ( .B1(n8208), .B2(n8206), .A(n8207), .ZN(n8230) );
  INV_X1 U9836 ( .A(n8230), .ZN(n8210) );
  NAND3_X1 U9837 ( .A1(n8208), .A2(n8207), .A3(n8206), .ZN(n8209) );
  AOI21_X1 U9838 ( .B1(n8210), .B2(n8209), .A(n8264), .ZN(n8211) );
  AOI211_X1 U9839 ( .C1(n8213), .C2(n8267), .A(n8212), .B(n8211), .ZN(n8214)
         );
  OAI21_X1 U9840 ( .B1(n8215), .B2(n8268), .A(n8214), .ZN(P2_U3199) );
  XNOR2_X1 U9841 ( .A(n8253), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8250) );
  NAND2_X1 U9842 ( .A1(n8217), .A2(n8216), .ZN(n8219) );
  NAND2_X1 U9843 ( .A1(n8219), .A2(n8218), .ZN(n8251) );
  XOR2_X1 U9844 ( .A(n8250), .B(n8251), .Z(n8245) );
  INV_X1 U9845 ( .A(n8220), .ZN(n8226) );
  OR2_X1 U9846 ( .A1(n8221), .A2(n8232), .ZN(n8225) );
  NAND2_X1 U9847 ( .A1(n8249), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8247) );
  NAND2_X1 U9848 ( .A1(n8253), .A2(n8222), .ZN(n8223) );
  NAND2_X1 U9849 ( .A1(n8247), .A2(n8223), .ZN(n8224) );
  AND3_X1 U9850 ( .A1(n8226), .A2(n8225), .A3(n8224), .ZN(n8228) );
  INV_X1 U9851 ( .A(n8268), .ZN(n8227) );
  OAI21_X1 U9852 ( .B1(n8248), .B2(n8228), .A(n8227), .ZN(n8244) );
  INV_X1 U9853 ( .A(n8229), .ZN(n8231) );
  AOI21_X1 U9854 ( .B1(n8232), .B2(n8231), .A(n8230), .ZN(n8234) );
  MUX2_X1 U9855 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8255), .Z(n8233) );
  NOR2_X1 U9856 ( .A1(n8234), .A2(n8233), .ZN(n8254) );
  NAND2_X1 U9857 ( .A1(n8234), .A2(n8233), .ZN(n8252) );
  INV_X1 U9858 ( .A(n8252), .ZN(n8235) );
  NOR2_X1 U9859 ( .A1(n8254), .A2(n8235), .ZN(n8238) );
  INV_X1 U9860 ( .A(n8238), .ZN(n8237) );
  OAI21_X1 U9861 ( .B1(n8237), .B2(n8236), .A(n10283), .ZN(n8240) );
  NOR2_X1 U9862 ( .A1(n8238), .A2(n8264), .ZN(n8239) );
  MUX2_X1 U9863 ( .A(n8240), .B(n8239), .S(n8249), .Z(n8241) );
  AOI211_X1 U9864 ( .C1(n10275), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8242), .B(
        n8241), .ZN(n8243) );
  OAI211_X1 U9865 ( .C1(n8246), .C2(n8245), .A(n8244), .B(n8243), .ZN(P2_U3200) );
  XNOR2_X1 U9866 ( .A(n8261), .B(n8382), .ZN(n8257) );
  XNOR2_X1 U9867 ( .A(n8261), .B(n8471), .ZN(n8256) );
  OAI21_X1 U9868 ( .B1(n8254), .B2(n8253), .A(n8252), .ZN(n8259) );
  MUX2_X1 U9869 ( .A(n8257), .B(n8256), .S(n8255), .Z(n8258) );
  XNOR2_X1 U9870 ( .A(n8259), .B(n8258), .ZN(n8265) );
  OAI21_X1 U9871 ( .B1(n10283), .B2(n8261), .A(n8260), .ZN(n8262) );
  AOI21_X1 U9872 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(n10275), .A(n8262), .ZN(
        n8263) );
  OAI21_X1 U9873 ( .B1(n8265), .B2(n8264), .A(n8263), .ZN(n8266) );
  NAND2_X1 U9874 ( .A1(n8270), .A2(n8269), .ZN(n8437) );
  OAI21_X1 U9875 ( .B1(n8437), .B2(n8381), .A(n8271), .ZN(n8274) );
  AOI21_X1 U9876 ( .B1(P2_REG2_REG_31__SCAN_IN), .B2(n8381), .A(n8274), .ZN(
        n8272) );
  OAI21_X1 U9877 ( .B1(n8273), .B2(n8361), .A(n8272), .ZN(P2_U3202) );
  AOI21_X1 U9878 ( .B1(P2_REG2_REG_30__SCAN_IN), .B2(n8381), .A(n8274), .ZN(
        n8275) );
  OAI21_X1 U9879 ( .B1(n8496), .B2(n8361), .A(n8275), .ZN(P2_U3203) );
  XNOR2_X1 U9880 ( .A(n8277), .B(n8276), .ZN(n8279) );
  AOI222_X1 U9881 ( .A1(n10289), .A2(n8279), .B1(n8278), .B2(n10286), .C1(
        n8298), .C2(n10285), .ZN(n8446) );
  XNOR2_X1 U9882 ( .A(n8280), .B(n4920), .ZN(n8444) );
  AOI22_X1 U9883 ( .A1(n8281), .A2(n10294), .B1(n8381), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8282) );
  OAI21_X1 U9884 ( .B1(n8283), .B2(n8361), .A(n8282), .ZN(n8284) );
  AOI21_X1 U9885 ( .B1(n8444), .B2(n10296), .A(n8284), .ZN(n8285) );
  OAI21_X1 U9886 ( .B1(n8446), .B2(n8381), .A(n8285), .ZN(P2_U3206) );
  XNOR2_X1 U9887 ( .A(n8286), .B(n8287), .ZN(n8503) );
  XNOR2_X1 U9888 ( .A(n8288), .B(n8287), .ZN(n8290) );
  AOI222_X1 U9889 ( .A1(n10289), .A2(n8290), .B1(n8312), .B2(n10285), .C1(
        n8289), .C2(n10286), .ZN(n8498) );
  MUX2_X1 U9890 ( .A(n8291), .B(n8498), .S(n10299), .Z(n8294) );
  AOI22_X1 U9891 ( .A1(n8500), .A2(n10292), .B1(n10294), .B2(n8292), .ZN(n8293) );
  OAI211_X1 U9892 ( .C1(n8503), .C2(n8420), .A(n8294), .B(n8293), .ZN(P2_U3207) );
  NOR2_X1 U9893 ( .A1(n8295), .A2(n8308), .ZN(n8301) );
  XNOR2_X1 U9894 ( .A(n8297), .B(n8296), .ZN(n8299) );
  AOI222_X1 U9895 ( .A1(n10289), .A2(n8299), .B1(n8328), .B2(n10285), .C1(
        n8298), .C2(n10286), .ZN(n8504) );
  INV_X1 U9896 ( .A(n8504), .ZN(n8300) );
  AOI211_X1 U9897 ( .C1(n10294), .C2(n8302), .A(n8301), .B(n8300), .ZN(n8307)
         );
  XNOR2_X1 U9898 ( .A(n8303), .B(n8304), .ZN(n8508) );
  INV_X1 U9899 ( .A(n8508), .ZN(n8305) );
  AOI22_X1 U9900 ( .A1(n8305), .A2(n10296), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8381), .ZN(n8306) );
  OAI21_X1 U9901 ( .B1(n8307), .B2(n8381), .A(n8306), .ZN(P2_U3208) );
  INV_X1 U9902 ( .A(n8511), .ZN(n8309) );
  NOR2_X1 U9903 ( .A1(n8309), .A2(n8308), .ZN(n8315) );
  XNOR2_X1 U9904 ( .A(n8311), .B(n8310), .ZN(n8313) );
  AOI222_X1 U9905 ( .A1(n10289), .A2(n8313), .B1(n8337), .B2(n10285), .C1(
        n8312), .C2(n10286), .ZN(n8509) );
  INV_X1 U9906 ( .A(n8509), .ZN(n8314) );
  AOI211_X1 U9907 ( .C1(n10294), .C2(n8316), .A(n8315), .B(n8314), .ZN(n8323)
         );
  NAND2_X1 U9908 ( .A1(n8318), .A2(n8317), .ZN(n8320) );
  XNOR2_X1 U9909 ( .A(n8320), .B(n8319), .ZN(n8514) );
  INV_X1 U9910 ( .A(n8514), .ZN(n8321) );
  AOI22_X1 U9911 ( .A1(n8321), .A2(n10296), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n8381), .ZN(n8322) );
  OAI21_X1 U9912 ( .B1(n8323), .B2(n8381), .A(n8322), .ZN(P2_U3209) );
  XNOR2_X1 U9913 ( .A(n8324), .B(n4758), .ZN(n8520) );
  INV_X1 U9914 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8330) );
  XNOR2_X1 U9915 ( .A(n8326), .B(n8325), .ZN(n8329) );
  AOI222_X1 U9916 ( .A1(n10289), .A2(n8329), .B1(n8328), .B2(n10286), .C1(
        n8327), .C2(n10285), .ZN(n8515) );
  MUX2_X1 U9917 ( .A(n8330), .B(n8515), .S(n10299), .Z(n8333) );
  AOI22_X1 U9918 ( .A1(n8517), .A2(n10292), .B1(n10294), .B2(n8331), .ZN(n8332) );
  OAI211_X1 U9919 ( .C1(n8520), .C2(n8420), .A(n8333), .B(n8332), .ZN(P2_U3210) );
  XNOR2_X1 U9920 ( .A(n8334), .B(n8335), .ZN(n8526) );
  XNOR2_X1 U9921 ( .A(n8336), .B(n8335), .ZN(n8338) );
  AOI222_X1 U9922 ( .A1(n10289), .A2(n8338), .B1(n7576), .B2(n10285), .C1(
        n8337), .C2(n10286), .ZN(n8521) );
  MUX2_X1 U9923 ( .A(n8339), .B(n8521), .S(n10299), .Z(n8342) );
  AOI22_X1 U9924 ( .A1(n8523), .A2(n10292), .B1(n10294), .B2(n8340), .ZN(n8341) );
  OAI211_X1 U9925 ( .C1(n8526), .C2(n8420), .A(n8342), .B(n8341), .ZN(P2_U3211) );
  XOR2_X1 U9926 ( .A(n8343), .B(n8348), .Z(n8344) );
  OAI222_X1 U9927 ( .A1(n8424), .A2(n8346), .B1(n8426), .B2(n8345), .C1(n10301), .C2(n8344), .ZN(n8461) );
  INV_X1 U9928 ( .A(n8461), .ZN(n8353) );
  XOR2_X1 U9929 ( .A(n8347), .B(n8348), .Z(n8462) );
  AOI22_X1 U9930 ( .A1(n8381), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n10294), .B2(
        n8349), .ZN(n8350) );
  OAI21_X1 U9931 ( .B1(n8530), .B2(n8361), .A(n8350), .ZN(n8351) );
  AOI21_X1 U9932 ( .B1(n8462), .B2(n10296), .A(n8351), .ZN(n8352) );
  OAI21_X1 U9933 ( .B1(n8353), .B2(n8381), .A(n8352), .ZN(P2_U3212) );
  OAI21_X1 U9934 ( .B1(n8355), .B2(n8358), .A(n8354), .ZN(n8357) );
  AOI222_X1 U9935 ( .A1(n10289), .A2(n8357), .B1(n7576), .B2(n10286), .C1(
        n8356), .C2(n10285), .ZN(n8465) );
  XOR2_X1 U9936 ( .A(n8359), .B(n8358), .Z(n8467) );
  NOR2_X1 U9937 ( .A1(n7574), .A2(n8361), .ZN(n8365) );
  OAI22_X1 U9938 ( .A1(n8433), .A2(n8363), .B1(n8362), .B2(n8430), .ZN(n8364)
         );
  AOI211_X1 U9939 ( .C1(n8467), .C2(n10296), .A(n8365), .B(n8364), .ZN(n8366)
         );
  OAI21_X1 U9940 ( .B1(n8465), .B2(n8381), .A(n8366), .ZN(P2_U3213) );
  OR2_X1 U9941 ( .A1(n8368), .A2(n8367), .ZN(n8370) );
  NAND2_X1 U9942 ( .A1(n8370), .A2(n8369), .ZN(n8372) );
  XNOR2_X1 U9943 ( .A(n8372), .B(n8371), .ZN(n8540) );
  NOR2_X1 U9944 ( .A1(n8374), .A2(n8373), .ZN(n8376) );
  AOI22_X1 U9945 ( .A1(n8378), .A2(n10286), .B1(n10285), .B2(n8377), .ZN(n8379) );
  MUX2_X1 U9946 ( .A(n8536), .B(n8382), .S(n8381), .Z(n8385) );
  AOI22_X1 U9947 ( .A1(n8537), .A2(n10292), .B1(n10294), .B2(n8383), .ZN(n8384) );
  OAI211_X1 U9948 ( .C1(n8540), .C2(n8420), .A(n8385), .B(n8384), .ZN(P2_U3214) );
  XNOR2_X1 U9949 ( .A(n8387), .B(n8386), .ZN(n8543) );
  XNOR2_X1 U9950 ( .A(n8388), .B(n8389), .ZN(n8390) );
  OAI222_X1 U9951 ( .A1(n8424), .A2(n8392), .B1(n8426), .B2(n8391), .C1(n8390), 
        .C2(n10301), .ZN(n8474) );
  NAND2_X1 U9952 ( .A1(n8474), .A2(n10299), .ZN(n8397) );
  OAI22_X1 U9953 ( .A1(n8433), .A2(n8394), .B1(n8393), .B2(n8430), .ZN(n8395)
         );
  AOI21_X1 U9954 ( .B1(n8475), .B2(n10292), .A(n8395), .ZN(n8396) );
  OAI211_X1 U9955 ( .C1(n8543), .C2(n8420), .A(n8397), .B(n8396), .ZN(P2_U3216) );
  XNOR2_X1 U9956 ( .A(n8398), .B(n8399), .ZN(n8549) );
  XNOR2_X1 U9957 ( .A(n8400), .B(n4886), .ZN(n8403) );
  AOI222_X1 U9958 ( .A1(n10289), .A2(n8403), .B1(n8402), .B2(n10286), .C1(
        n8401), .C2(n10285), .ZN(n8544) );
  MUX2_X1 U9959 ( .A(n8404), .B(n8544), .S(n10299), .Z(n8408) );
  INV_X1 U9960 ( .A(n8405), .ZN(n8406) );
  AOI22_X1 U9961 ( .A1(n8546), .A2(n10292), .B1(n10294), .B2(n8406), .ZN(n8407) );
  OAI211_X1 U9962 ( .C1(n8549), .C2(n8420), .A(n8408), .B(n8407), .ZN(P2_U3217) );
  XOR2_X1 U9963 ( .A(n8409), .B(n8411), .Z(n8556) );
  XNOR2_X1 U9964 ( .A(n8410), .B(n8411), .ZN(n8414) );
  AOI222_X1 U9965 ( .A1(n10289), .A2(n8414), .B1(n8413), .B2(n10285), .C1(
        n8412), .C2(n10286), .ZN(n8550) );
  MUX2_X1 U9966 ( .A(n8415), .B(n8550), .S(n10299), .Z(n8419) );
  INV_X1 U9967 ( .A(n8416), .ZN(n8417) );
  AOI22_X1 U9968 ( .A1(n8552), .A2(n10292), .B1(n10294), .B2(n8417), .ZN(n8418) );
  OAI211_X1 U9969 ( .C1(n8556), .C2(n8420), .A(n8419), .B(n8418), .ZN(P2_U3218) );
  XNOR2_X1 U9970 ( .A(n8421), .B(n8429), .ZN(n8422) );
  OAI222_X1 U9971 ( .A1(n8426), .A2(n8425), .B1(n8424), .B2(n8423), .C1(n8422), 
        .C2(n10301), .ZN(n8485) );
  AOI21_X1 U9972 ( .B1(n8427), .B2(n8558), .A(n8485), .ZN(n8436) );
  XNOR2_X1 U9973 ( .A(n8428), .B(n8429), .ZN(n8561) );
  OAI22_X1 U9974 ( .A1(n8433), .A2(n8432), .B1(n8431), .B2(n8430), .ZN(n8434)
         );
  AOI21_X1 U9975 ( .B1(n8561), .B2(n10296), .A(n8434), .ZN(n8435) );
  OAI21_X1 U9976 ( .B1(n8436), .B2(n8381), .A(n8435), .ZN(P2_U3219) );
  NAND2_X1 U9977 ( .A1(n8490), .A2(n8486), .ZN(n8438) );
  INV_X1 U9978 ( .A(n8437), .ZN(n8491) );
  NAND2_X1 U9979 ( .A1(n8491), .A2(n10386), .ZN(n8440) );
  OAI211_X1 U9980 ( .C1(n10386), .C2(n7676), .A(n8438), .B(n8440), .ZN(
        P2_U3490) );
  INV_X1 U9981 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8442) );
  NAND2_X1 U9982 ( .A1(n8439), .A2(n8486), .ZN(n8441) );
  OAI211_X1 U9983 ( .C1(n10386), .C2(n8442), .A(n8441), .B(n8440), .ZN(
        P2_U3489) );
  AOI22_X1 U9984 ( .A1(n8444), .A2(n10345), .B1(n10366), .B2(n8443), .ZN(n8445) );
  NAND2_X1 U9985 ( .A1(n8446), .A2(n8445), .ZN(n8497) );
  MUX2_X1 U9986 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8497), .S(n10386), .Z(
        P2_U3486) );
  INV_X1 U9987 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8447) );
  MUX2_X1 U9988 ( .A(n8447), .B(n8498), .S(n10386), .Z(n8449) );
  NAND2_X1 U9989 ( .A1(n8500), .A2(n8486), .ZN(n8448) );
  OAI211_X1 U9990 ( .C1(n8503), .C2(n8484), .A(n8449), .B(n8448), .ZN(P2_U3485) );
  INV_X1 U9991 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8450) );
  MUX2_X1 U9992 ( .A(n8450), .B(n8504), .S(n10386), .Z(n8452) );
  NAND2_X1 U9993 ( .A1(n8505), .A2(n8486), .ZN(n8451) );
  OAI211_X1 U9994 ( .C1(n8508), .C2(n8484), .A(n8452), .B(n8451), .ZN(P2_U3484) );
  MUX2_X1 U9995 ( .A(n9690), .B(n8509), .S(n10386), .Z(n8454) );
  NAND2_X1 U9996 ( .A1(n8511), .A2(n8486), .ZN(n8453) );
  OAI211_X1 U9997 ( .C1(n8484), .C2(n8514), .A(n8454), .B(n8453), .ZN(P2_U3483) );
  MUX2_X1 U9998 ( .A(n8455), .B(n8515), .S(n10386), .Z(n8457) );
  NAND2_X1 U9999 ( .A1(n8517), .A2(n8486), .ZN(n8456) );
  OAI211_X1 U10000 ( .C1(n8520), .C2(n8484), .A(n8457), .B(n8456), .ZN(
        P2_U3482) );
  INV_X1 U10001 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8458) );
  MUX2_X1 U10002 ( .A(n8458), .B(n8521), .S(n10386), .Z(n8460) );
  NAND2_X1 U10003 ( .A1(n8523), .A2(n8486), .ZN(n8459) );
  OAI211_X1 U10004 ( .C1(n8526), .C2(n8484), .A(n8460), .B(n8459), .ZN(
        P2_U3481) );
  INV_X1 U10005 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8463) );
  AOI21_X1 U10006 ( .B1(n8462), .B2(n10345), .A(n8461), .ZN(n8527) );
  MUX2_X1 U10007 ( .A(n8463), .B(n8527), .S(n10386), .Z(n8464) );
  OAI21_X1 U10008 ( .B1(n8530), .B2(n8470), .A(n8464), .ZN(P2_U3480) );
  INV_X1 U10009 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8468) );
  INV_X1 U10010 ( .A(n8465), .ZN(n8466) );
  AOI21_X1 U10011 ( .B1(n8467), .B2(n10345), .A(n8466), .ZN(n8531) );
  MUX2_X1 U10012 ( .A(n8468), .B(n8531), .S(n10386), .Z(n8469) );
  OAI21_X1 U10013 ( .B1(n7574), .B2(n8470), .A(n8469), .ZN(P2_U3479) );
  MUX2_X1 U10014 ( .A(n8471), .B(n8536), .S(n10386), .Z(n8473) );
  NAND2_X1 U10015 ( .A1(n8537), .A2(n8486), .ZN(n8472) );
  OAI211_X1 U10016 ( .C1(n8540), .C2(n8484), .A(n8473), .B(n8472), .ZN(
        P2_U3478) );
  AOI21_X1 U10017 ( .B1(n10366), .B2(n8475), .A(n8474), .ZN(n8541) );
  MUX2_X1 U10018 ( .A(n8476), .B(n8541), .S(n10386), .Z(n8477) );
  OAI21_X1 U10019 ( .B1(n8543), .B2(n8484), .A(n8477), .ZN(P2_U3476) );
  MUX2_X1 U10020 ( .A(n8478), .B(n8544), .S(n10386), .Z(n8480) );
  NAND2_X1 U10021 ( .A1(n8546), .A2(n8486), .ZN(n8479) );
  OAI211_X1 U10022 ( .C1(n8549), .C2(n8484), .A(n8480), .B(n8479), .ZN(
        P2_U3475) );
  MUX2_X1 U10023 ( .A(n8481), .B(n8550), .S(n10386), .Z(n8483) );
  NAND2_X1 U10024 ( .A1(n8552), .A2(n8486), .ZN(n8482) );
  OAI211_X1 U10025 ( .C1(n8484), .C2(n8556), .A(n8483), .B(n8482), .ZN(
        P2_U3474) );
  INV_X1 U10026 ( .A(n8485), .ZN(n8557) );
  MUX2_X1 U10027 ( .A(n9471), .B(n8557), .S(n10386), .Z(n8489) );
  AOI22_X1 U10028 ( .A1(n8561), .A2(n8487), .B1(n8486), .B2(n8558), .ZN(n8488)
         );
  NAND2_X1 U10029 ( .A1(n8489), .A2(n8488), .ZN(P2_U3473) );
  INV_X1 U10030 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8493) );
  NAND2_X1 U10031 ( .A1(n8490), .A2(n8559), .ZN(n8492) );
  NAND2_X1 U10032 ( .A1(n8491), .A2(n10367), .ZN(n8494) );
  OAI211_X1 U10033 ( .C1(n8493), .C2(n10367), .A(n8492), .B(n8494), .ZN(
        P2_U3458) );
  NAND2_X1 U10034 ( .A1(n10369), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8495) );
  OAI211_X1 U10035 ( .C1(n8496), .C2(n8534), .A(n8495), .B(n8494), .ZN(
        P2_U3457) );
  MUX2_X1 U10036 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8497), .S(n10367), .Z(
        P2_U3454) );
  INV_X1 U10037 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8499) );
  MUX2_X1 U10038 ( .A(n8499), .B(n8498), .S(n10367), .Z(n8502) );
  NAND2_X1 U10039 ( .A1(n8500), .A2(n8559), .ZN(n8501) );
  OAI211_X1 U10040 ( .C1(n8503), .C2(n8555), .A(n8502), .B(n8501), .ZN(
        P2_U3453) );
  MUX2_X1 U10041 ( .A(n9457), .B(n8504), .S(n10367), .Z(n8507) );
  NAND2_X1 U10042 ( .A1(n8505), .A2(n8559), .ZN(n8506) );
  OAI211_X1 U10043 ( .C1(n8508), .C2(n8555), .A(n8507), .B(n8506), .ZN(
        P2_U3452) );
  INV_X1 U10044 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8510) );
  MUX2_X1 U10045 ( .A(n8510), .B(n8509), .S(n10367), .Z(n8513) );
  NAND2_X1 U10046 ( .A1(n8511), .A2(n8559), .ZN(n8512) );
  OAI211_X1 U10047 ( .C1(n8514), .C2(n8555), .A(n8513), .B(n8512), .ZN(
        P2_U3451) );
  INV_X1 U10048 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8516) );
  MUX2_X1 U10049 ( .A(n8516), .B(n8515), .S(n10367), .Z(n8519) );
  NAND2_X1 U10050 ( .A1(n8517), .A2(n8559), .ZN(n8518) );
  OAI211_X1 U10051 ( .C1(n8520), .C2(n8555), .A(n8519), .B(n8518), .ZN(
        P2_U3450) );
  INV_X1 U10052 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8522) );
  MUX2_X1 U10053 ( .A(n8522), .B(n8521), .S(n10367), .Z(n8525) );
  NAND2_X1 U10054 ( .A1(n8523), .A2(n8559), .ZN(n8524) );
  OAI211_X1 U10055 ( .C1(n8526), .C2(n8555), .A(n8525), .B(n8524), .ZN(
        P2_U3449) );
  INV_X1 U10056 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8528) );
  MUX2_X1 U10057 ( .A(n8528), .B(n8527), .S(n10367), .Z(n8529) );
  OAI21_X1 U10058 ( .B1(n8530), .B2(n8534), .A(n8529), .ZN(P2_U3448) );
  MUX2_X1 U10059 ( .A(n8532), .B(n8531), .S(n10367), .Z(n8533) );
  OAI21_X1 U10060 ( .B1(n7574), .B2(n8534), .A(n8533), .ZN(P2_U3447) );
  INV_X1 U10061 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8535) );
  MUX2_X1 U10062 ( .A(n8536), .B(n8535), .S(n10369), .Z(n8539) );
  NAND2_X1 U10063 ( .A1(n8537), .A2(n8559), .ZN(n8538) );
  OAI211_X1 U10064 ( .C1(n8540), .C2(n8555), .A(n8539), .B(n8538), .ZN(
        P2_U3446) );
  MUX2_X1 U10065 ( .A(n9691), .B(n8541), .S(n10367), .Z(n8542) );
  OAI21_X1 U10066 ( .B1(n8543), .B2(n8555), .A(n8542), .ZN(P2_U3441) );
  INV_X1 U10067 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8545) );
  MUX2_X1 U10068 ( .A(n8545), .B(n8544), .S(n10367), .Z(n8548) );
  NAND2_X1 U10069 ( .A1(n8546), .A2(n8559), .ZN(n8547) );
  OAI211_X1 U10070 ( .C1(n8549), .C2(n8555), .A(n8548), .B(n8547), .ZN(
        P2_U3438) );
  INV_X1 U10071 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8551) );
  MUX2_X1 U10072 ( .A(n8551), .B(n8550), .S(n10367), .Z(n8554) );
  NAND2_X1 U10073 ( .A1(n8552), .A2(n8559), .ZN(n8553) );
  OAI211_X1 U10074 ( .C1(n8556), .C2(n8555), .A(n8554), .B(n8553), .ZN(
        P2_U3435) );
  MUX2_X1 U10075 ( .A(n9623), .B(n8557), .S(n10367), .Z(n8563) );
  AOI22_X1 U10076 ( .A1(n8561), .A2(n8560), .B1(n8559), .B2(n8558), .ZN(n8562)
         );
  NAND2_X1 U10077 ( .A1(n8563), .A2(n8562), .ZN(P2_U3432) );
  NAND2_X1 U10078 ( .A1(n9807), .A2(n8568), .ZN(n8566) );
  OR4_X1 U10079 ( .A1(n8564), .A2(n6279), .A3(P2_U3151), .A4(
        P2_IR_REG_30__SCAN_IN), .ZN(n8565) );
  OAI211_X1 U10080 ( .C1(n8567), .C2(n8578), .A(n8566), .B(n8565), .ZN(
        P2_U3264) );
  NAND2_X1 U10081 ( .A1(n8569), .A2(n8568), .ZN(n8571) );
  OAI211_X1 U10082 ( .C1(n8578), .C2(n9496), .A(n8571), .B(n8570), .ZN(
        P2_U3267) );
  INV_X1 U10083 ( .A(n8572), .ZN(n9816) );
  AOI21_X1 U10084 ( .B1(n8574), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8573), .ZN(
        n8575) );
  OAI21_X1 U10085 ( .B1(n9816), .B2(n8576), .A(n8575), .ZN(P2_U3268) );
  INV_X1 U10086 ( .A(n8577), .ZN(n9819) );
  OAI222_X1 U10087 ( .A1(n8582), .A2(n9819), .B1(P2_U3151), .B2(n8580), .C1(
        n8579), .C2(n8578), .ZN(P2_U3269) );
  MUX2_X1 U10088 ( .A(n8583), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AOI21_X1 U10089 ( .B1(n8586), .B2(n8585), .A(n8584), .ZN(n8587) );
  OAI21_X1 U10090 ( .B1(n8588), .B2(n8587), .A(n8680), .ZN(n8594) );
  INV_X1 U10091 ( .A(n9174), .ZN(n8589) );
  NOR2_X1 U10092 ( .A1(n8589), .A2(n8696), .ZN(n8591) );
  OAI22_X1 U10093 ( .A1(n9123), .A2(n8683), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9616), .ZN(n8590) );
  AOI211_X1 U10094 ( .C1(n8693), .C2(n9180), .A(n8591), .B(n8590), .ZN(n8593)
         );
  NAND2_X1 U10095 ( .A1(n9730), .A2(n8731), .ZN(n8592) );
  NAND3_X1 U10096 ( .A1(n8594), .A2(n8593), .A3(n8592), .ZN(P1_U3214) );
  XNOR2_X1 U10097 ( .A(n8596), .B(n8595), .ZN(n8597) );
  XNOR2_X1 U10098 ( .A(n8598), .B(n8597), .ZN(n8605) );
  NAND2_X1 U10099 ( .A1(n8725), .A2(n8599), .ZN(n8602) );
  NOR2_X1 U10100 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8600), .ZN(n10016) );
  AOI21_X1 U10101 ( .B1(n8726), .B2(n9010), .A(n10016), .ZN(n8601) );
  OAI211_X1 U10102 ( .C1(n10237), .C2(n8729), .A(n8602), .B(n8601), .ZN(n8603)
         );
  AOI21_X1 U10103 ( .B1(n10240), .B2(n8731), .A(n8603), .ZN(n8604) );
  OAI21_X1 U10104 ( .B1(n8605), .B2(n8733), .A(n8604), .ZN(P1_U3215) );
  INV_X1 U10105 ( .A(n8606), .ZN(n8690) );
  INV_X1 U10106 ( .A(n8607), .ZN(n8609) );
  NOR3_X1 U10107 ( .A1(n8690), .A2(n8609), .A3(n8608), .ZN(n8611) );
  INV_X1 U10108 ( .A(n8610), .ZN(n8663) );
  OAI21_X1 U10109 ( .B1(n8611), .B2(n8663), .A(n8680), .ZN(n8616) );
  INV_X1 U10110 ( .A(n9237), .ZN(n8614) );
  AOI22_X1 U10111 ( .A1(n9754), .A2(n8693), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n8612) );
  OAI21_X1 U10112 ( .B1(n9241), .B2(n8683), .A(n8612), .ZN(n8613) );
  AOI21_X1 U10113 ( .B1(n8614), .B2(n8725), .A(n8613), .ZN(n8615) );
  OAI211_X1 U10114 ( .C1(n9757), .C2(n8689), .A(n8616), .B(n8615), .ZN(
        P1_U3216) );
  XNOR2_X1 U10115 ( .A(n8618), .B(n8617), .ZN(n8619) );
  XNOR2_X1 U10116 ( .A(n8620), .B(n8619), .ZN(n8625) );
  NAND2_X1 U10117 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9089) );
  NAND2_X1 U10118 ( .A1(n8693), .A2(n9783), .ZN(n8621) );
  OAI211_X1 U10119 ( .C1(n9889), .C2(n8683), .A(n9089), .B(n8621), .ZN(n8623)
         );
  NOR2_X1 U10120 ( .A1(n9787), .A2(n8689), .ZN(n8622) );
  AOI211_X1 U10121 ( .C1(n9294), .C2(n8725), .A(n8623), .B(n8622), .ZN(n8624)
         );
  OAI21_X1 U10122 ( .B1(n8625), .B2(n8733), .A(n8624), .ZN(P1_U3219) );
  INV_X1 U10123 ( .A(n9272), .ZN(n9770) );
  OAI21_X1 U10124 ( .B1(n8628), .B2(n8627), .A(n8626), .ZN(n8629) );
  NAND2_X1 U10125 ( .A1(n8629), .A2(n8680), .ZN(n8633) );
  AOI22_X1 U10126 ( .A1(n8726), .A2(n9783), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n8630) );
  OAI21_X1 U10127 ( .B1(n9241), .B2(n8729), .A(n8630), .ZN(n8631) );
  AOI21_X1 U10128 ( .B1(n9267), .B2(n8725), .A(n8631), .ZN(n8632) );
  OAI211_X1 U10129 ( .C1(n9770), .C2(n8689), .A(n8633), .B(n8632), .ZN(
        P1_U3223) );
  INV_X1 U10130 ( .A(n9202), .ZN(n9743) );
  OAI21_X1 U10131 ( .B1(n8635), .B2(n8634), .A(n5832), .ZN(n8636) );
  NAND2_X1 U10132 ( .A1(n8636), .A2(n8680), .ZN(n8640) );
  AOI22_X1 U10133 ( .A1(n9741), .A2(n8693), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n8637) );
  OAI21_X1 U10134 ( .B1(n9206), .B2(n8683), .A(n8637), .ZN(n8638) );
  AOI21_X1 U10135 ( .B1(n9203), .B2(n8725), .A(n8638), .ZN(n8639) );
  OAI211_X1 U10136 ( .C1(n9743), .C2(n8689), .A(n8640), .B(n8639), .ZN(
        P1_U3225) );
  XNOR2_X1 U10137 ( .A(n8641), .B(n8642), .ZN(n8724) );
  NOR2_X1 U10138 ( .A1(n8724), .A2(n8723), .ZN(n8722) );
  AOI21_X1 U10139 ( .B1(n8642), .B2(n8641), .A(n8722), .ZN(n8646) );
  XNOR2_X1 U10140 ( .A(n8644), .B(n8643), .ZN(n8645) );
  XNOR2_X1 U10141 ( .A(n8646), .B(n8645), .ZN(n8652) );
  NAND2_X1 U10142 ( .A1(n8693), .A2(n9898), .ZN(n8647) );
  OAI211_X1 U10143 ( .C1(n10237), .C2(n8683), .A(n8648), .B(n8647), .ZN(n8650)
         );
  NOR2_X1 U10144 ( .A1(n4802), .A2(n8689), .ZN(n8649) );
  AOI211_X1 U10145 ( .C1(n9323), .C2(n8725), .A(n8650), .B(n8649), .ZN(n8651)
         );
  OAI21_X1 U10146 ( .B1(n8652), .B2(n8733), .A(n8651), .ZN(P1_U3226) );
  INV_X1 U10147 ( .A(n9892), .ZN(n9313) );
  OAI211_X1 U10148 ( .C1(n8655), .C2(n8654), .A(n8653), .B(n8680), .ZN(n8659)
         );
  NAND2_X1 U10149 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9068) );
  OAI21_X1 U10150 ( .B1(n9908), .B2(n8683), .A(n9068), .ZN(n8657) );
  NOR2_X1 U10151 ( .A1(n8696), .A2(n9307), .ZN(n8656) );
  AOI211_X1 U10152 ( .C1(n8693), .C2(n9784), .A(n8657), .B(n8656), .ZN(n8658)
         );
  OAI211_X1 U10153 ( .C1(n9313), .C2(n8689), .A(n8659), .B(n8658), .ZN(
        P1_U3228) );
  INV_X1 U10154 ( .A(n8660), .ZN(n8662) );
  NOR3_X1 U10155 ( .A1(n8663), .A2(n8662), .A3(n8661), .ZN(n8666) );
  INV_X1 U10156 ( .A(n8664), .ZN(n8665) );
  OAI21_X1 U10157 ( .B1(n8666), .B2(n8665), .A(n8680), .ZN(n8670) );
  AOI22_X1 U10158 ( .A1(n9251), .A2(n8726), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8667) );
  OAI21_X1 U10159 ( .B1(n8837), .B2(n8729), .A(n8667), .ZN(n8668) );
  AOI21_X1 U10160 ( .B1(n9219), .B2(n8725), .A(n8668), .ZN(n8669) );
  OAI211_X1 U10161 ( .C1(n9221), .C2(n8689), .A(n8670), .B(n8669), .ZN(
        P1_U3229) );
  AOI21_X1 U10162 ( .B1(n8672), .B2(n8671), .A(n4589), .ZN(n8677) );
  NAND2_X1 U10163 ( .A1(n8725), .A2(n9280), .ZN(n8674) );
  AOI22_X1 U10164 ( .A1(n8693), .A2(n9775), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n8673) );
  OAI211_X1 U10165 ( .C1(n9283), .C2(n8683), .A(n8674), .B(n8673), .ZN(n8675)
         );
  AOI21_X1 U10166 ( .B1(n9285), .B2(n8731), .A(n8675), .ZN(n8676) );
  OAI21_X1 U10167 ( .B1(n8677), .B2(n8733), .A(n8676), .ZN(P1_U3233) );
  XNOR2_X1 U10168 ( .A(n8679), .B(n8678), .ZN(n8681) );
  NAND2_X1 U10169 ( .A1(n8681), .A2(n8680), .ZN(n8688) );
  OAI22_X1 U10170 ( .A1(n10206), .A2(n8683), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8682), .ZN(n8685) );
  NOR2_X1 U10171 ( .A1(n8729), .A2(n9907), .ZN(n8684) );
  AOI211_X1 U10172 ( .C1(n8686), .C2(n8725), .A(n8685), .B(n8684), .ZN(n8687)
         );
  OAI211_X1 U10173 ( .C1(n10228), .C2(n8689), .A(n8688), .B(n8687), .ZN(
        P1_U3234) );
  AOI21_X1 U10174 ( .B1(n8692), .B2(n8691), .A(n8690), .ZN(n8699) );
  AOI22_X1 U10175 ( .A1(n8726), .A2(n9775), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n8695) );
  NAND2_X1 U10176 ( .A1(n9251), .A2(n8693), .ZN(n8694) );
  OAI211_X1 U10177 ( .C1(n8696), .C2(n9248), .A(n8695), .B(n8694), .ZN(n8697)
         );
  AOI21_X1 U10178 ( .B1(n9763), .B2(n8731), .A(n8697), .ZN(n8698) );
  OAI21_X1 U10179 ( .B1(n8699), .B2(n8733), .A(n8698), .ZN(P1_U3235) );
  AOI21_X1 U10180 ( .B1(n8702), .B2(n8701), .A(n8700), .ZN(n8706) );
  XNOR2_X1 U10181 ( .A(n8704), .B(n8703), .ZN(n8705) );
  XNOR2_X1 U10182 ( .A(n8706), .B(n8705), .ZN(n8712) );
  NAND2_X1 U10183 ( .A1(n8725), .A2(n8707), .ZN(n8709) );
  AOI22_X1 U10184 ( .A1(n8726), .A2(n9012), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n8708) );
  OAI211_X1 U10185 ( .C1(n10206), .C2(n8729), .A(n8709), .B(n8708), .ZN(n8710)
         );
  AOI21_X1 U10186 ( .B1(n10209), .B2(n8731), .A(n8710), .ZN(n8711) );
  OAI21_X1 U10187 ( .B1(n8712), .B2(n8733), .A(n8711), .ZN(P1_U3236) );
  INV_X1 U10188 ( .A(n8713), .ZN(n8714) );
  AOI21_X1 U10189 ( .B1(n8716), .B2(n8715), .A(n8714), .ZN(n8721) );
  NAND2_X1 U10190 ( .A1(n8725), .A2(n9873), .ZN(n8718) );
  AOI22_X1 U10191 ( .A1(n8726), .A2(n9898), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n8717) );
  OAI211_X1 U10192 ( .C1(n9283), .C2(n8729), .A(n8718), .B(n8717), .ZN(n8719)
         );
  AOI21_X1 U10193 ( .B1(n9874), .B2(n8731), .A(n8719), .ZN(n8720) );
  OAI21_X1 U10194 ( .B1(n8721), .B2(n8733), .A(n8720), .ZN(P1_U3238) );
  AOI21_X1 U10195 ( .B1(n8724), .B2(n8723), .A(n8722), .ZN(n8734) );
  NAND2_X1 U10196 ( .A1(n8725), .A2(n9345), .ZN(n8728) );
  AOI22_X1 U10197 ( .A1(n8726), .A2(n9103), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n8727) );
  OAI211_X1 U10198 ( .C1(n9908), .C2(n8729), .A(n8728), .B(n8727), .ZN(n8730)
         );
  AOI21_X1 U10199 ( .B1(n9911), .B2(n8731), .A(n8730), .ZN(n8732) );
  OAI21_X1 U10200 ( .B1(n8734), .B2(n8733), .A(n8732), .ZN(P1_U3241) );
  NAND2_X1 U10201 ( .A1(n9807), .A2(n8738), .ZN(n8736) );
  INV_X1 U10202 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9810) );
  OR2_X1 U10203 ( .A1(n8745), .A2(n9810), .ZN(n8735) );
  AOI211_X1 U10204 ( .C1(n8992), .C2(n8995), .A(n9005), .B(n8737), .ZN(n9002)
         );
  INV_X1 U10205 ( .A(n8855), .ZN(n8860) );
  NAND2_X1 U10206 ( .A1(n9095), .A2(n9094), .ZN(n8864) );
  OR2_X1 U10207 ( .A1(n8745), .A2(n8740), .ZN(n8741) );
  NAND2_X1 U10208 ( .A1(n8744), .A2(n8738), .ZN(n8747) );
  OR2_X1 U10209 ( .A1(n8745), .A2(n9811), .ZN(n8746) );
  NAND4_X1 U10210 ( .A1(n8927), .A2(n9722), .A3(n8855), .A4(n9131), .ZN(n8751)
         );
  NAND2_X1 U10211 ( .A1(n9091), .A2(n9149), .ZN(n8989) );
  NAND2_X1 U10212 ( .A1(n9091), .A2(n9094), .ZN(n8748) );
  NAND2_X1 U10213 ( .A1(n8989), .A2(n8748), .ZN(n8928) );
  NOR3_X1 U10214 ( .A1(n9131), .A2(n9722), .A3(n8855), .ZN(n8749) );
  NAND2_X1 U10215 ( .A1(n8751), .A2(n8750), .ZN(n8752) );
  NAND2_X1 U10216 ( .A1(n9330), .A2(n9908), .ZN(n8907) );
  INV_X1 U10217 ( .A(n8753), .ZN(n8773) );
  NOR2_X1 U10218 ( .A1(n8754), .A2(n8773), .ZN(n8938) );
  NAND2_X1 U10219 ( .A1(n8938), .A2(n8860), .ZN(n8760) );
  INV_X1 U10220 ( .A(n8755), .ZN(n8756) );
  OAI211_X1 U10221 ( .C1(n10087), .C2(n8756), .A(n8943), .B(n8762), .ZN(n8757)
         );
  INV_X1 U10222 ( .A(n8757), .ZN(n8758) );
  AND2_X1 U10223 ( .A1(n8775), .A2(n8761), .ZN(n8948) );
  NAND2_X1 U10224 ( .A1(n8774), .A2(n8948), .ZN(n8767) );
  INV_X1 U10225 ( .A(n8948), .ZN(n8763) );
  OAI21_X1 U10226 ( .B1(n8763), .B2(n8762), .A(n8772), .ZN(n8947) );
  INV_X1 U10227 ( .A(n8777), .ZN(n8764) );
  NOR2_X1 U10228 ( .A1(n8947), .A2(n8764), .ZN(n8766) );
  AOI21_X1 U10229 ( .B1(n8767), .B2(n8766), .A(n8765), .ZN(n8770) );
  OAI21_X1 U10230 ( .B1(n8770), .B2(n8769), .A(n8768), .ZN(n8771) );
  NAND2_X1 U10231 ( .A1(n8771), .A2(n8879), .ZN(n8784) );
  OAI211_X1 U10232 ( .C1(n8774), .C2(n8773), .A(n8944), .B(n8772), .ZN(n8776)
         );
  NAND3_X1 U10233 ( .A1(n8776), .A2(n8775), .A3(n8950), .ZN(n8778) );
  NAND2_X1 U10234 ( .A1(n8778), .A2(n8777), .ZN(n8780) );
  NAND2_X1 U10235 ( .A1(n8780), .A2(n8779), .ZN(n8782) );
  INV_X1 U10236 ( .A(n8956), .ZN(n8785) );
  NAND2_X1 U10237 ( .A1(n8787), .A2(n8953), .ZN(n8788) );
  OAI211_X1 U10238 ( .C1(n8789), .C2(n8788), .A(n8962), .B(n8957), .ZN(n8791)
         );
  AOI21_X1 U10239 ( .B1(n8791), .B2(n8790), .A(n8959), .ZN(n8793) );
  NAND2_X1 U10240 ( .A1(n8887), .A2(n8966), .ZN(n8792) );
  OAI211_X1 U10241 ( .C1(n8793), .C2(n8792), .A(n8855), .B(n8907), .ZN(n8810)
         );
  INV_X1 U10242 ( .A(n8953), .ZN(n8794) );
  AOI21_X1 U10243 ( .B1(n8796), .B2(n8795), .A(n8794), .ZN(n8799) );
  INV_X1 U10244 ( .A(n8797), .ZN(n8798) );
  OAI21_X1 U10245 ( .B1(n8799), .B2(n8798), .A(n8961), .ZN(n8801) );
  INV_X1 U10246 ( .A(n8966), .ZN(n8800) );
  AOI21_X1 U10247 ( .B1(n8801), .B2(n8962), .A(n8800), .ZN(n8805) );
  INV_X1 U10248 ( .A(n8802), .ZN(n8804) );
  OR2_X1 U10249 ( .A1(n9911), .A2(n10237), .ZN(n8812) );
  AND2_X1 U10250 ( .A1(n8967), .A2(n8860), .ZN(n8803) );
  AND2_X1 U10251 ( .A1(n8812), .A2(n8803), .ZN(n8807) );
  OAI211_X1 U10252 ( .C1(n8805), .C2(n8804), .A(n8807), .B(n8973), .ZN(n8809)
         );
  NAND2_X1 U10253 ( .A1(n9911), .A2(n10237), .ZN(n8906) );
  NAND2_X1 U10254 ( .A1(n8906), .A2(n8806), .ZN(n8969) );
  INV_X1 U10255 ( .A(n8807), .ZN(n8808) );
  AOI22_X1 U10256 ( .A1(n8810), .A2(n8809), .B1(n8969), .B2(n8808), .ZN(n8811)
         );
  AOI21_X1 U10257 ( .B1(n4761), .B2(n8860), .A(n8811), .ZN(n8816) );
  INV_X1 U10258 ( .A(n8812), .ZN(n8970) );
  NAND2_X1 U10259 ( .A1(n8907), .A2(n8970), .ZN(n8813) );
  MUX2_X1 U10260 ( .A(n8906), .B(n8813), .S(n8855), .Z(n8814) );
  MUX2_X1 U10261 ( .A(n8860), .B(n8814), .S(n8973), .Z(n8815) );
  INV_X1 U10262 ( .A(n9898), .ZN(n9108) );
  OR2_X1 U10263 ( .A1(n9892), .A2(n9108), .ZN(n9868) );
  NAND2_X1 U10264 ( .A1(n9874), .A2(n9889), .ZN(n8909) );
  INV_X1 U10265 ( .A(n8908), .ZN(n8817) );
  NAND2_X1 U10266 ( .A1(n8909), .A2(n8817), .ZN(n8937) );
  AOI21_X1 U10267 ( .B1(n8822), .B2(n9868), .A(n8937), .ZN(n8818) );
  OR2_X1 U10268 ( .A1(n9298), .A2(n9283), .ZN(n8869) );
  OR2_X1 U10269 ( .A1(n9874), .A2(n9889), .ZN(n8870) );
  NAND2_X1 U10270 ( .A1(n8869), .A2(n8870), .ZN(n8976) );
  NAND2_X1 U10271 ( .A1(n9298), .A2(n9283), .ZN(n8911) );
  INV_X1 U10272 ( .A(n9783), .ZN(n9270) );
  NAND2_X1 U10273 ( .A1(n9285), .A2(n9270), .ZN(n9261) );
  OAI211_X1 U10274 ( .C1(n8818), .C2(n8976), .A(n8911), .B(n9261), .ZN(n8820)
         );
  INV_X1 U10275 ( .A(n9775), .ZN(n8868) );
  OR2_X1 U10276 ( .A1(n9272), .A2(n8868), .ZN(n8913) );
  OR2_X1 U10277 ( .A1(n9285), .A2(n9270), .ZN(n9260) );
  NAND2_X1 U10278 ( .A1(n8913), .A2(n9260), .ZN(n9138) );
  INV_X1 U10279 ( .A(n9138), .ZN(n8819) );
  AND2_X1 U10280 ( .A1(n8870), .A2(n9868), .ZN(n8974) );
  INV_X1 U10281 ( .A(n8974), .ZN(n8821) );
  OAI211_X1 U10282 ( .C1(n8822), .C2(n8821), .A(n8911), .B(n8909), .ZN(n8823)
         );
  NAND3_X1 U10283 ( .A1(n8823), .A2(n8869), .A3(n9260), .ZN(n8825) );
  NAND2_X1 U10284 ( .A1(n9272), .A2(n8868), .ZN(n8826) );
  NAND2_X1 U10285 ( .A1(n8826), .A2(n9261), .ZN(n8914) );
  INV_X1 U10286 ( .A(n8914), .ZN(n8824) );
  MUX2_X1 U10287 ( .A(n8826), .B(n8913), .S(n8855), .Z(n8827) );
  OR2_X1 U10288 ( .A1(n9763), .A2(n9241), .ZN(n8833) );
  NAND2_X1 U10289 ( .A1(n9763), .A2(n9241), .ZN(n8828) );
  NAND2_X1 U10290 ( .A1(n8833), .A2(n8828), .ZN(n9253) );
  INV_X1 U10291 ( .A(n9251), .ZN(n9116) );
  AND2_X1 U10292 ( .A1(n9243), .A2(n9116), .ZN(n8866) );
  INV_X1 U10293 ( .A(n8828), .ZN(n8829) );
  NOR2_X1 U10294 ( .A1(n8866), .A2(n8829), .ZN(n8916) );
  NAND2_X1 U10295 ( .A1(n9750), .A2(n9206), .ZN(n8915) );
  INV_X1 U10296 ( .A(n8915), .ZN(n8830) );
  NOR3_X1 U10297 ( .A1(n8830), .A2(n8866), .A3(n8860), .ZN(n8832) );
  INV_X1 U10298 ( .A(n8900), .ZN(n9141) );
  NOR2_X1 U10299 ( .A1(n9243), .A2(n9116), .ZN(n8867) );
  NOR3_X1 U10300 ( .A1(n9141), .A2(n8867), .A3(n8855), .ZN(n8831) );
  INV_X1 U10301 ( .A(n8833), .ZN(n9139) );
  OR2_X1 U10302 ( .A1(n8867), .A2(n9139), .ZN(n8899) );
  XNOR2_X1 U10303 ( .A(n8915), .B(n8855), .ZN(n8834) );
  INV_X1 U10304 ( .A(n8866), .ZN(n9140) );
  OAI211_X1 U10305 ( .C1(n8899), .C2(n8860), .A(n8834), .B(n9140), .ZN(n8835)
         );
  OAI211_X1 U10306 ( .C1(n8860), .C2(n8900), .A(n8836), .B(n8835), .ZN(n8842)
         );
  NAND2_X1 U10307 ( .A1(n9736), .A2(n9123), .ZN(n8985) );
  INV_X1 U10308 ( .A(n8865), .ZN(n9185) );
  INV_X1 U10309 ( .A(n9143), .ZN(n8839) );
  NOR2_X1 U10310 ( .A1(n9202), .A2(n8837), .ZN(n8912) );
  NAND2_X1 U10311 ( .A1(n9143), .A2(n8912), .ZN(n8838) );
  NOR2_X1 U10312 ( .A1(n9736), .A2(n9123), .ZN(n9142) );
  INV_X1 U10313 ( .A(n9142), .ZN(n8898) );
  AND2_X1 U10314 ( .A1(n8838), .A2(n8898), .ZN(n8840) );
  OAI21_X1 U10315 ( .B1(n8842), .B2(n8839), .A(n8840), .ZN(n8844) );
  INV_X1 U10316 ( .A(n8840), .ZN(n8841) );
  AOI21_X1 U10317 ( .B1(n8842), .B2(n9143), .A(n8841), .ZN(n8843) );
  INV_X1 U10318 ( .A(n8897), .ZN(n8845) );
  NAND2_X1 U10319 ( .A1(n9160), .A2(n9715), .ZN(n9145) );
  NAND2_X1 U10320 ( .A1(n9730), .A2(n9193), .ZN(n9144) );
  AND2_X1 U10321 ( .A1(n9145), .A2(n9144), .ZN(n8848) );
  OAI21_X1 U10322 ( .B1(n8849), .B2(n8845), .A(n8848), .ZN(n8846) );
  NAND2_X1 U10323 ( .A1(n9131), .A2(n9722), .ZN(n8988) );
  AOI211_X1 U10324 ( .C1(n8846), .C2(n8895), .A(n8855), .B(n9146), .ZN(n8847)
         );
  INV_X1 U10325 ( .A(n8848), .ZN(n8923) );
  AOI21_X1 U10326 ( .B1(n8849), .B2(n8897), .A(n8923), .ZN(n8852) );
  NAND3_X1 U10327 ( .A1(n9128), .A2(n8855), .A3(n8895), .ZN(n8850) );
  NAND3_X1 U10328 ( .A1(n8854), .A2(n8853), .A3(n4544), .ZN(n8859) );
  INV_X1 U10329 ( .A(n8928), .ZN(n8856) );
  OAI21_X1 U10330 ( .B1(n8860), .B2(n8864), .A(n8863), .ZN(n9001) );
  INV_X1 U10331 ( .A(n8861), .ZN(n8862) );
  INV_X1 U10332 ( .A(n8864), .ZN(n8930) );
  NOR2_X1 U10333 ( .A1(n8930), .A2(n5126), .ZN(n8994) );
  XNOR2_X1 U10334 ( .A(n9736), .B(n9123), .ZN(n9189) );
  NAND2_X1 U10335 ( .A1(n8895), .A2(n9145), .ZN(n9155) );
  NAND2_X1 U10336 ( .A1(n8897), .A2(n9144), .ZN(n9127) );
  NAND2_X1 U10337 ( .A1(n8900), .A2(n8915), .ZN(n9225) );
  INV_X1 U10338 ( .A(n9225), .ZN(n9214) );
  NOR2_X1 U10339 ( .A1(n8867), .A2(n8866), .ZN(n9234) );
  INV_X1 U10340 ( .A(n9234), .ZN(n9231) );
  XNOR2_X1 U10341 ( .A(n9272), .B(n8868), .ZN(n9264) );
  XNOR2_X1 U10342 ( .A(n9285), .B(n9783), .ZN(n9278) );
  INV_X1 U10343 ( .A(n9868), .ZN(n8871) );
  XNOR2_X1 U10344 ( .A(n9911), .B(n10237), .ZN(n9337) );
  NAND2_X1 U10345 ( .A1(n8973), .A2(n8907), .ZN(n9319) );
  NAND3_X1 U10346 ( .A1(n8872), .A2(n10094), .A3(n8939), .ZN(n8877) );
  NAND2_X1 U10347 ( .A1(n8873), .A2(n10079), .ZN(n8876) );
  NOR4_X1 U10348 ( .A1(n8877), .A2(n8876), .A3(n8875), .A4(n8874), .ZN(n8880)
         );
  NAND4_X1 U10349 ( .A1(n8880), .A2(n8879), .A3(n10068), .A4(n8878), .ZN(n8884) );
  NOR4_X1 U10350 ( .A1(n8884), .A2(n8883), .A3(n8882), .A4(n8881), .ZN(n8888)
         );
  NAND4_X1 U10351 ( .A1(n8888), .A2(n8887), .A3(n8886), .A4(n8885), .ZN(n8889)
         );
  NOR4_X1 U10352 ( .A1(n9304), .A2(n9337), .A3(n9319), .A4(n8889), .ZN(n8890)
         );
  NAND4_X1 U10353 ( .A1(n9278), .A2(n9290), .A3(n9876), .A4(n8890), .ZN(n8891)
         );
  NOR4_X1 U10354 ( .A1(n9231), .A2(n9264), .A3(n9253), .A4(n8891), .ZN(n8892)
         );
  NAND4_X1 U10355 ( .A1(n9179), .A2(n9210), .A3(n9214), .A4(n8892), .ZN(n8893)
         );
  NOR4_X1 U10356 ( .A1(n9146), .A2(n9189), .A3(n9155), .A4(n8893), .ZN(n8894)
         );
  AND4_X1 U10357 ( .A1(n8994), .A2(n8894), .A3(n8933), .A4(n8989), .ZN(n8936)
         );
  NAND2_X1 U10358 ( .A1(n8896), .A2(n8895), .ZN(n8991) );
  NAND2_X1 U10359 ( .A1(n8898), .A2(n8897), .ZN(n8983) );
  INV_X1 U10360 ( .A(n8983), .ZN(n8925) );
  NAND2_X1 U10361 ( .A1(n8899), .A2(n9140), .ZN(n8901) );
  NAND2_X1 U10362 ( .A1(n8901), .A2(n8900), .ZN(n8902) );
  NAND2_X1 U10363 ( .A1(n8902), .A2(n8915), .ZN(n8918) );
  INV_X1 U10364 ( .A(n8918), .ZN(n8904) );
  OR2_X1 U10365 ( .A1(n8912), .A2(n9138), .ZN(n8903) );
  OR2_X1 U10366 ( .A1(n8904), .A2(n8903), .ZN(n8979) );
  NAND2_X1 U10367 ( .A1(n8905), .A2(n8967), .ZN(n9336) );
  OR2_X2 U10368 ( .A1(n9336), .A2(n9337), .ZN(n9334) );
  INV_X1 U10369 ( .A(n9319), .ZN(n9318) );
  NAND2_X1 U10370 ( .A1(n9869), .A2(n8974), .ZN(n8910) );
  NAND2_X1 U10371 ( .A1(n8910), .A2(n8909), .ZN(n9291) );
  INV_X1 U10372 ( .A(n8911), .ZN(n8982) );
  OAI21_X1 U10373 ( .B1(n8979), .B2(n9277), .A(n8985), .ZN(n8924) );
  INV_X1 U10374 ( .A(n8912), .ZN(n8919) );
  NAND2_X1 U10375 ( .A1(n8914), .A2(n8913), .ZN(n9137) );
  NAND3_X1 U10376 ( .A1(n8916), .A2(n8915), .A3(n9137), .ZN(n8917) );
  NAND3_X1 U10377 ( .A1(n8919), .A2(n8918), .A3(n8917), .ZN(n8920) );
  AND2_X1 U10378 ( .A1(n8920), .A2(n9185), .ZN(n8921) );
  NOR2_X1 U10379 ( .A1(n8983), .A2(n8921), .ZN(n8922) );
  OR2_X1 U10380 ( .A1(n8923), .A2(n8922), .ZN(n8987) );
  AOI21_X1 U10381 ( .B1(n8925), .B2(n8924), .A(n8987), .ZN(n8926) );
  OAI21_X1 U10382 ( .B1(n8991), .B2(n8926), .A(n8988), .ZN(n8929) );
  OAI21_X1 U10383 ( .B1(n8929), .B2(n8928), .A(n8927), .ZN(n8932) );
  AOI211_X1 U10384 ( .C1(n8933), .C2(n8932), .A(n8931), .B(n8930), .ZN(n8934)
         );
  OAI21_X1 U10385 ( .B1(n8936), .B2(n8934), .A(n9086), .ZN(n8935) );
  INV_X1 U10386 ( .A(n8937), .ZN(n8978) );
  INV_X1 U10387 ( .A(n8938), .ZN(n8946) );
  AOI21_X1 U10388 ( .B1(n6717), .B2(n10117), .A(n8939), .ZN(n8942) );
  INV_X1 U10389 ( .A(n8940), .ZN(n8941) );
  AND3_X1 U10390 ( .A1(n8943), .A2(n8942), .A3(n8941), .ZN(n8945) );
  OAI21_X1 U10391 ( .B1(n8946), .B2(n8945), .A(n8944), .ZN(n8949) );
  AOI21_X1 U10392 ( .B1(n8949), .B2(n8948), .A(n8947), .ZN(n8955) );
  NAND2_X1 U10393 ( .A1(n8951), .A2(n8950), .ZN(n8954) );
  OAI211_X1 U10394 ( .C1(n8955), .C2(n8954), .A(n8953), .B(n8952), .ZN(n8958)
         );
  NAND4_X1 U10395 ( .A1(n8958), .A2(n8962), .A3(n8957), .A4(n8956), .ZN(n8960)
         );
  OR2_X1 U10396 ( .A1(n8960), .A2(n8959), .ZN(n8968) );
  INV_X1 U10397 ( .A(n8961), .ZN(n8964) );
  NAND3_X1 U10398 ( .A1(n8964), .A2(n8963), .A3(n8962), .ZN(n8965) );
  NAND4_X1 U10399 ( .A1(n8968), .A2(n8967), .A3(n8966), .A4(n8965), .ZN(n8972)
         );
  INV_X1 U10400 ( .A(n8969), .ZN(n8971) );
  AOI21_X1 U10401 ( .B1(n8972), .B2(n8971), .A(n8970), .ZN(n8975) );
  OAI211_X1 U10402 ( .C1(n4761), .C2(n8975), .A(n8974), .B(n8973), .ZN(n8977)
         );
  AOI21_X1 U10403 ( .B1(n8978), .B2(n8977), .A(n8976), .ZN(n8981) );
  INV_X1 U10404 ( .A(n8979), .ZN(n8980) );
  OAI21_X1 U10405 ( .B1(n8982), .B2(n8981), .A(n8980), .ZN(n8984) );
  AOI21_X1 U10406 ( .B1(n8985), .B2(n8984), .A(n8983), .ZN(n8986) );
  NOR2_X1 U10407 ( .A1(n8987), .A2(n8986), .ZN(n8990) );
  OAI211_X1 U10408 ( .C1(n8991), .C2(n8990), .A(n8989), .B(n8988), .ZN(n8993)
         );
  AOI21_X1 U10409 ( .B1(n8994), .B2(n8993), .A(n8992), .ZN(n8996) );
  XNOR2_X1 U10410 ( .A(n8996), .B(n8995), .ZN(n8998) );
  AOI21_X1 U10411 ( .B1(n9002), .B2(n9001), .A(n9000), .ZN(n9008) );
  NAND3_X1 U10412 ( .A1(n9003), .A2(n10194), .A3(n9024), .ZN(n9004) );
  OAI211_X1 U10413 ( .C1(n9005), .C2(n9007), .A(n9004), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9006) );
  OAI21_X1 U10414 ( .B1(n9008), .B2(n9007), .A(n9006), .ZN(P1_U3242) );
  MUX2_X1 U10415 ( .A(n9009), .B(P1_DATAO_REG_29__SCAN_IN), .S(n9030), .Z(
        P1_U3583) );
  MUX2_X1 U10416 ( .A(n9180), .B(P1_DATAO_REG_28__SCAN_IN), .S(n9030), .Z(
        P1_U3582) );
  MUX2_X1 U10417 ( .A(n9735), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9030), .Z(
        P1_U3581) );
  MUX2_X1 U10418 ( .A(n9741), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9030), .Z(
        P1_U3580) );
  MUX2_X1 U10419 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9222), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10420 ( .A(n9754), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9030), .Z(
        P1_U3578) );
  MUX2_X1 U10421 ( .A(n9251), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9030), .Z(
        P1_U3577) );
  MUX2_X1 U10422 ( .A(n9767), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9030), .Z(
        P1_U3576) );
  MUX2_X1 U10423 ( .A(n9775), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9030), .Z(
        P1_U3575) );
  MUX2_X1 U10424 ( .A(n9783), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9030), .Z(
        P1_U3574) );
  MUX2_X1 U10425 ( .A(n9871), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9030), .Z(
        P1_U3573) );
  MUX2_X1 U10426 ( .A(n9784), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9030), .Z(
        P1_U3572) );
  MUX2_X1 U10427 ( .A(n9898), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9030), .Z(
        P1_U3571) );
  MUX2_X1 U10428 ( .A(n9343), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9030), .Z(
        P1_U3570) );
  MUX2_X1 U10429 ( .A(n9897), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9030), .Z(
        P1_U3569) );
  MUX2_X1 U10430 ( .A(n9103), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9030), .Z(
        P1_U3568) );
  MUX2_X1 U10431 ( .A(n9010), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9030), .Z(
        P1_U3567) );
  MUX2_X1 U10432 ( .A(n9011), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9030), .Z(
        P1_U3566) );
  MUX2_X1 U10433 ( .A(n10192), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9030), .Z(
        P1_U3565) );
  MUX2_X1 U10434 ( .A(n9012), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9030), .Z(
        P1_U3564) );
  MUX2_X1 U10435 ( .A(n10193), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9030), .Z(
        P1_U3563) );
  MUX2_X1 U10436 ( .A(n10184), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9030), .Z(
        P1_U3562) );
  MUX2_X1 U10437 ( .A(n10065), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9030), .Z(
        P1_U3561) );
  MUX2_X1 U10438 ( .A(n10166), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9030), .Z(
        P1_U3560) );
  MUX2_X1 U10439 ( .A(n6632), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9030), .Z(
        P1_U3559) );
  MUX2_X1 U10440 ( .A(n5287), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9030), .Z(
        P1_U3558) );
  MUX2_X1 U10441 ( .A(n10089), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9030), .Z(
        P1_U3557) );
  MUX2_X1 U10442 ( .A(n9013), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9030), .Z(
        P1_U3556) );
  MUX2_X1 U10443 ( .A(n6717), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9030), .Z(
        P1_U3555) );
  OAI211_X1 U10444 ( .C1(n9016), .C2(n9015), .A(n9988), .B(n9014), .ZN(n9023)
         );
  AOI22_X1 U10445 ( .A1(n9945), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9022) );
  NAND2_X1 U10446 ( .A1(n10043), .A2(n9017), .ZN(n9021) );
  OAI211_X1 U10447 ( .C1(n9019), .C2(n9025), .A(n9983), .B(n9018), .ZN(n9020)
         );
  NAND4_X1 U10448 ( .A1(n9023), .A2(n9022), .A3(n9021), .A4(n9020), .ZN(
        P1_U3244) );
  MUX2_X1 U10449 ( .A(n9026), .B(n9025), .S(n9024), .Z(n9028) );
  NAND2_X1 U10450 ( .A1(n9028), .A2(n9027), .ZN(n9032) );
  NOR2_X1 U10451 ( .A1(n9924), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9029) );
  OR2_X1 U10452 ( .A1(n9029), .A2(n5872), .ZN(n9925) );
  INV_X1 U10453 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9926) );
  AND2_X1 U10454 ( .A1(n9925), .A2(n9926), .ZN(n9929) );
  NOR2_X1 U10455 ( .A1(n9030), .A2(n9929), .ZN(n9031) );
  NAND2_X1 U10456 ( .A1(n9032), .A2(n9031), .ZN(n9947) );
  INV_X1 U10457 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9034) );
  INV_X1 U10458 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9033) );
  OAI22_X1 U10459 ( .A1(n10046), .A2(n9034), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9033), .ZN(n9035) );
  AOI21_X1 U10460 ( .B1(n9036), .B2(n10043), .A(n9035), .ZN(n9045) );
  OAI211_X1 U10461 ( .C1(n9039), .C2(n9038), .A(n9988), .B(n9037), .ZN(n9044)
         );
  OAI211_X1 U10462 ( .C1(n9042), .C2(n9041), .A(n9983), .B(n9040), .ZN(n9043)
         );
  NAND4_X1 U10463 ( .A1(n9947), .A2(n9045), .A3(n9044), .A4(n9043), .ZN(
        P1_U3245) );
  OAI211_X1 U10464 ( .C1(n9048), .C2(n9047), .A(n9988), .B(n9046), .ZN(n9058)
         );
  INV_X1 U10465 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9050) );
  OAI21_X1 U10466 ( .B1(n10046), .B2(n9050), .A(n9049), .ZN(n9051) );
  AOI21_X1 U10467 ( .B1(n9052), .B2(n10043), .A(n9051), .ZN(n9057) );
  OAI211_X1 U10468 ( .C1(n9055), .C2(n9054), .A(n9983), .B(n9053), .ZN(n9056)
         );
  NAND3_X1 U10469 ( .A1(n9058), .A2(n9057), .A3(n9056), .ZN(P1_U3246) );
  AOI22_X1 U10470 ( .A1(n9080), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9308), .B2(
        n9069), .ZN(n9061) );
  OAI21_X1 U10471 ( .B1(n9061), .B2(n9060), .A(n9075), .ZN(n9062) );
  NAND2_X1 U10472 ( .A1(n9062), .A2(n9983), .ZN(n9074) );
  AOI22_X1 U10473 ( .A1(n9080), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n5608), .B2(
        n9069), .ZN(n9066) );
  OAI21_X1 U10474 ( .B1(n9066), .B2(n9065), .A(n9079), .ZN(n9072) );
  NAND2_X1 U10475 ( .A1(n9945), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9067) );
  OAI211_X1 U10476 ( .C1(n9070), .C2(n9069), .A(n9068), .B(n9067), .ZN(n9071)
         );
  AOI21_X1 U10477 ( .B1(n9072), .B2(n9988), .A(n9071), .ZN(n9073) );
  NAND2_X1 U10478 ( .A1(n9074), .A2(n9073), .ZN(P1_U3260) );
  NAND2_X1 U10479 ( .A1(n10042), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9076) );
  OAI21_X1 U10480 ( .B1(n10042), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9076), .ZN(
        n10038) );
  AOI21_X1 U10481 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n10042), .A(n10037), 
        .ZN(n9077) );
  XNOR2_X1 U10482 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9077), .ZN(n9085) );
  INV_X1 U10483 ( .A(n9085), .ZN(n9083) );
  INV_X1 U10484 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9888) );
  NOR2_X1 U10485 ( .A1(n10042), .A2(n9888), .ZN(n9078) );
  AOI21_X1 U10486 ( .B1(n10042), .B2(n9888), .A(n9078), .ZN(n10034) );
  NOR2_X1 U10487 ( .A1(n10034), .A2(n10035), .ZN(n10033) );
  AOI21_X1 U10488 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n10042), .A(n10033), 
        .ZN(n9081) );
  AOI211_X1 U10489 ( .C1(n9083), .C2(n9983), .A(n10043), .B(n9082), .ZN(n9088)
         );
  AOI22_X1 U10490 ( .A1(n9085), .A2(n9983), .B1(n9988), .B2(n9084), .ZN(n9087)
         );
  MUX2_X1 U10491 ( .A(n9088), .B(n9087), .S(n9086), .Z(n9090) );
  OAI211_X1 U10492 ( .C1(n5168), .C2(n10046), .A(n9090), .B(n9089), .ZN(
        P1_U3262) );
  NAND2_X1 U10493 ( .A1(n9216), .A2(n9221), .ZN(n9217) );
  NAND2_X1 U10494 ( .A1(n9201), .A2(n9195), .ZN(n9194) );
  NOR2_X2 U10495 ( .A1(n9194), .A2(n9730), .ZN(n9173) );
  NAND2_X1 U10496 ( .A1(n9711), .A2(n9130), .ZN(n9098) );
  XOR2_X1 U10497 ( .A(n9095), .B(n9098), .Z(n9092) );
  NAND2_X1 U10498 ( .A1(n9092), .A2(n10097), .ZN(n9354) );
  INV_X1 U10499 ( .A(P1_B_REG_SCAN_IN), .ZN(n9469) );
  OR2_X1 U10500 ( .A1(n9924), .A2(n9469), .ZN(n9093) );
  NAND2_X1 U10501 ( .A1(n10191), .A2(n9093), .ZN(n9148) );
  OR2_X1 U10502 ( .A1(n9094), .A2(n9148), .ZN(n9709) );
  NOR2_X1 U10503 ( .A1(n4495), .A2(n9709), .ZN(n9100) );
  INV_X1 U10504 ( .A(n9095), .ZN(n9355) );
  NOR2_X1 U10505 ( .A1(n9355), .A2(n9341), .ZN(n9096) );
  AOI211_X1 U10506 ( .C1(n4495), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9100), .B(
        n9096), .ZN(n9097) );
  OAI21_X1 U10507 ( .B1(n9354), .B2(n9327), .A(n9097), .ZN(P1_U3263) );
  OAI211_X1 U10508 ( .C1(n9711), .C2(n9130), .A(n10097), .B(n9098), .ZN(n9710)
         );
  NOR2_X1 U10509 ( .A1(n9711), .A2(n9341), .ZN(n9099) );
  AOI211_X1 U10510 ( .C1(n4495), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9100), .B(
        n9099), .ZN(n9101) );
  OAI21_X1 U10511 ( .B1(n9710), .B2(n9327), .A(n9101), .ZN(P1_U3264) );
  NAND2_X1 U10512 ( .A1(n9102), .A2(n9907), .ZN(n9105) );
  NAND2_X1 U10513 ( .A1(n9911), .A2(n9897), .ZN(n9107) );
  INV_X1 U10514 ( .A(n9911), .ZN(n9342) );
  AOI22_X1 U10515 ( .A1(n9338), .A2(n9107), .B1(n9342), .B2(n10237), .ZN(n9320) );
  NAND2_X1 U10516 ( .A1(n9320), .A2(n9319), .ZN(n9321) );
  NOR2_X1 U10517 ( .A1(n9313), .A2(n9108), .ZN(n9109) );
  NOR2_X1 U10518 ( .A1(n9874), .A2(n9784), .ZN(n9110) );
  NOR2_X1 U10519 ( .A1(n9787), .A2(n9283), .ZN(n9111) );
  NAND2_X1 U10520 ( .A1(n9778), .A2(n9270), .ZN(n9113) );
  NOR2_X1 U10521 ( .A1(n9778), .A2(n9270), .ZN(n9112) );
  AOI21_X2 U10522 ( .B1(n9276), .B2(n9113), .A(n9112), .ZN(n9259) );
  NAND2_X1 U10523 ( .A1(n9272), .A2(n9775), .ZN(n9115) );
  NOR2_X1 U10524 ( .A1(n9272), .A2(n9775), .ZN(n9114) );
  NOR2_X1 U10525 ( .A1(n9757), .A2(n9116), .ZN(n9117) );
  NAND2_X1 U10526 ( .A1(n9750), .A2(n9754), .ZN(n9118) );
  NAND2_X1 U10527 ( .A1(n9215), .A2(n9118), .ZN(n9120) );
  NAND2_X1 U10528 ( .A1(n9221), .A2(n9206), .ZN(n9119) );
  NAND2_X1 U10529 ( .A1(n9120), .A2(n9119), .ZN(n9200) );
  NOR2_X1 U10530 ( .A1(n9202), .A2(n9222), .ZN(n9121) );
  NAND2_X1 U10531 ( .A1(n9202), .A2(n9222), .ZN(n9122) );
  NOR2_X1 U10532 ( .A1(n9195), .A2(n9123), .ZN(n9125) );
  NAND2_X1 U10533 ( .A1(n9195), .A2(n9123), .ZN(n9124) );
  NOR2_X1 U10534 ( .A1(n9730), .A2(n9735), .ZN(n9126) );
  NAND2_X1 U10535 ( .A1(n9156), .A2(n9155), .ZN(n9154) );
  NAND2_X1 U10536 ( .A1(n9154), .A2(n5114), .ZN(n9129) );
  XNOR2_X1 U10537 ( .A(n9129), .B(n9128), .ZN(n9714) );
  INV_X1 U10538 ( .A(n9714), .ZN(n9153) );
  AOI211_X1 U10539 ( .C1(n9131), .C2(n9157), .A(n9339), .B(n9130), .ZN(n9718)
         );
  INV_X1 U10540 ( .A(n9131), .ZN(n9716) );
  NOR2_X1 U10541 ( .A1(n9716), .A2(n9341), .ZN(n9136) );
  INV_X1 U10542 ( .A(n9132), .ZN(n9133) );
  AOI22_X1 U10543 ( .A1(n9133), .A2(n10092), .B1(P1_REG2_REG_29__SCAN_IN), 
        .B2(n4495), .ZN(n9134) );
  OAI21_X1 U10544 ( .B1(n9715), .B2(n9348), .A(n9134), .ZN(n9135) );
  AOI211_X1 U10545 ( .C1(n9718), .C2(n10101), .A(n9136), .B(n9135), .ZN(n9152)
         );
  NAND2_X1 U10546 ( .A1(n9233), .A2(n9140), .ZN(n9224) );
  NAND2_X1 U10547 ( .A1(n9177), .A2(n9144), .ZN(n9166) );
  INV_X1 U10548 ( .A(n9155), .ZN(n9167) );
  NAND2_X1 U10549 ( .A1(n9166), .A2(n9167), .ZN(n9165) );
  NAND2_X1 U10550 ( .A1(n9165), .A2(n9145), .ZN(n9147) );
  OAI22_X1 U10551 ( .A1(n9150), .A2(n10222), .B1(n9149), .B2(n9148), .ZN(n9719) );
  NAND2_X1 U10552 ( .A1(n9719), .A2(n9309), .ZN(n9151) );
  OAI211_X1 U10553 ( .C1(n9153), .C2(n9322), .A(n9152), .B(n9151), .ZN(
        P1_U3356) );
  OAI21_X1 U10554 ( .B1(n9156), .B2(n9155), .A(n9154), .ZN(n9728) );
  INV_X1 U10555 ( .A(n9173), .ZN(n9159) );
  INV_X1 U10556 ( .A(n9157), .ZN(n9158) );
  AOI211_X1 U10557 ( .C1(n9160), .C2(n9159), .A(n9339), .B(n9158), .ZN(n9725)
         );
  NAND2_X1 U10558 ( .A1(n9160), .A2(n10090), .ZN(n9164) );
  INV_X1 U10559 ( .A(n9161), .ZN(n9162) );
  AOI22_X1 U10560 ( .A1(n9162), .A2(n10092), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n4495), .ZN(n9163) );
  OAI211_X1 U10561 ( .C1(n9722), .C2(n9192), .A(n9164), .B(n9163), .ZN(n9170)
         );
  OAI21_X1 U10562 ( .B1(n9167), .B2(n9166), .A(n9165), .ZN(n9168) );
  AOI22_X1 U10563 ( .A1(n9168), .A2(n10203), .B1(n10194), .B2(n9735), .ZN(
        n9727) );
  NOR2_X1 U10564 ( .A1(n9727), .A2(n4495), .ZN(n9169) );
  AOI211_X1 U10565 ( .C1(n9725), .C2(n10101), .A(n9170), .B(n9169), .ZN(n9171)
         );
  OAI21_X1 U10566 ( .B1(n9728), .B2(n9322), .A(n9171), .ZN(P1_U3265) );
  XNOR2_X1 U10567 ( .A(n9172), .B(n9179), .ZN(n9733) );
  AOI211_X1 U10568 ( .C1(n9730), .C2(n9194), .A(n9339), .B(n9173), .ZN(n9729)
         );
  AOI22_X1 U10569 ( .A1(n9174), .A2(n10092), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n4495), .ZN(n9175) );
  OAI21_X1 U10570 ( .B1(n9176), .B2(n9341), .A(n9175), .ZN(n9183) );
  OAI21_X1 U10571 ( .B1(n9179), .B2(n9178), .A(n9177), .ZN(n9181) );
  AOI222_X1 U10572 ( .A1(n10203), .A2(n9181), .B1(n9180), .B2(n10191), .C1(
        n9741), .C2(n10194), .ZN(n9732) );
  NOR2_X1 U10573 ( .A1(n9732), .A2(n4495), .ZN(n9182) );
  AOI211_X1 U10574 ( .C1(n10101), .C2(n9729), .A(n9183), .B(n9182), .ZN(n9184)
         );
  OAI21_X1 U10575 ( .B1(n9733), .B2(n9322), .A(n9184), .ZN(P1_U3266) );
  NAND2_X1 U10576 ( .A1(n9209), .A2(n9185), .ZN(n9186) );
  XOR2_X1 U10577 ( .A(n9189), .B(n9186), .Z(n9187) );
  XOR2_X1 U10578 ( .A(n9189), .B(n9188), .Z(n9734) );
  NAND2_X1 U10579 ( .A1(n9734), .A2(n10102), .ZN(n9199) );
  AOI22_X1 U10580 ( .A1(n9190), .A2(n10092), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n4495), .ZN(n9191) );
  OAI21_X1 U10581 ( .B1(n9193), .B2(n9192), .A(n9191), .ZN(n9197) );
  OAI211_X1 U10582 ( .C1(n9201), .C2(n9195), .A(n9194), .B(n10097), .ZN(n9737)
         );
  NOR2_X1 U10583 ( .A1(n9737), .A2(n9327), .ZN(n9196) );
  AOI211_X1 U10584 ( .C1(n10090), .C2(n9736), .A(n9197), .B(n9196), .ZN(n9198)
         );
  OAI211_X1 U10585 ( .C1(n4495), .C2(n9739), .A(n9199), .B(n9198), .ZN(
        P1_U3267) );
  XNOR2_X1 U10586 ( .A(n9200), .B(n9210), .ZN(n9748) );
  AOI211_X1 U10587 ( .C1(n9202), .C2(n9217), .A(n9339), .B(n9201), .ZN(n9745)
         );
  NOR2_X1 U10588 ( .A1(n9743), .A2(n9341), .ZN(n9208) );
  NAND2_X1 U10589 ( .A1(n9344), .A2(n9741), .ZN(n9205) );
  AOI22_X1 U10590 ( .A1(P1_REG2_REG_25__SCAN_IN), .A2(n4495), .B1(n9203), .B2(
        n10092), .ZN(n9204) );
  OAI211_X1 U10591 ( .C1(n9206), .C2(n9348), .A(n9205), .B(n9204), .ZN(n9207)
         );
  AOI211_X1 U10592 ( .C1(n9745), .C2(n10101), .A(n9208), .B(n9207), .ZN(n9213)
         );
  OAI21_X1 U10593 ( .B1(n9211), .B2(n9210), .A(n9209), .ZN(n9746) );
  NAND2_X1 U10594 ( .A1(n9746), .A2(n9301), .ZN(n9212) );
  OAI211_X1 U10595 ( .C1(n9748), .C2(n9322), .A(n9213), .B(n9212), .ZN(
        P1_U3268) );
  XNOR2_X1 U10596 ( .A(n9215), .B(n9214), .ZN(n9753) );
  INV_X1 U10597 ( .A(n9216), .ZN(n9236) );
  INV_X1 U10598 ( .A(n9217), .ZN(n9218) );
  AOI211_X1 U10599 ( .C1(n9750), .C2(n9236), .A(n9339), .B(n9218), .ZN(n9749)
         );
  AOI22_X1 U10600 ( .A1(n4495), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9219), .B2(
        n10092), .ZN(n9220) );
  OAI21_X1 U10601 ( .B1(n9221), .B2(n9341), .A(n9220), .ZN(n9229) );
  AND2_X1 U10602 ( .A1(n9222), .A2(n10191), .ZN(n9227) );
  AOI211_X1 U10603 ( .C1(n9225), .C2(n9224), .A(n10222), .B(n9223), .ZN(n9226)
         );
  AOI211_X1 U10604 ( .C1(n10194), .C2(n9251), .A(n9227), .B(n9226), .ZN(n9752)
         );
  NOR2_X1 U10605 ( .A1(n9752), .A2(n4495), .ZN(n9228) );
  AOI211_X1 U10606 ( .C1(n9749), .C2(n10101), .A(n9229), .B(n9228), .ZN(n9230)
         );
  OAI21_X1 U10607 ( .B1(n9753), .B2(n9322), .A(n9230), .ZN(P1_U3269) );
  XNOR2_X1 U10608 ( .A(n9232), .B(n9231), .ZN(n9761) );
  OAI21_X1 U10609 ( .B1(n9235), .B2(n9234), .A(n9233), .ZN(n9759) );
  OAI211_X1 U10610 ( .C1(n9757), .C2(n4582), .A(n9236), .B(n10097), .ZN(n9756)
         );
  OAI22_X1 U10611 ( .A1(n9309), .A2(n9238), .B1(n9237), .B2(n9306), .ZN(n9239)
         );
  AOI21_X1 U10612 ( .B1(n9344), .B2(n9754), .A(n9239), .ZN(n9240) );
  OAI21_X1 U10613 ( .B1(n9241), .B2(n9348), .A(n9240), .ZN(n9242) );
  AOI21_X1 U10614 ( .B1(n9243), .B2(n10090), .A(n9242), .ZN(n9244) );
  OAI21_X1 U10615 ( .B1(n9756), .B2(n9327), .A(n9244), .ZN(n9245) );
  AOI21_X1 U10616 ( .B1(n9759), .B2(n9301), .A(n9245), .ZN(n9246) );
  OAI21_X1 U10617 ( .B1(n9761), .B2(n9322), .A(n9246), .ZN(P1_U3270) );
  XNOR2_X1 U10618 ( .A(n9247), .B(n9253), .ZN(n9766) );
  AOI211_X1 U10619 ( .C1(n9763), .C2(n9265), .A(n9339), .B(n4582), .ZN(n9762)
         );
  INV_X1 U10620 ( .A(n9248), .ZN(n9249) );
  AOI22_X1 U10621 ( .A1(n4495), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9249), .B2(
        n10092), .ZN(n9250) );
  OAI21_X1 U10622 ( .B1(n4796), .B2(n9341), .A(n9250), .ZN(n9257) );
  AND2_X1 U10623 ( .A1(n9251), .A2(n10191), .ZN(n9255) );
  AOI211_X1 U10624 ( .C1(n9253), .C2(n9252), .A(n10222), .B(n4570), .ZN(n9254)
         );
  AOI211_X1 U10625 ( .C1(n10194), .C2(n9775), .A(n9255), .B(n9254), .ZN(n9765)
         );
  NOR2_X1 U10626 ( .A1(n9765), .A2(n4495), .ZN(n9256) );
  AOI211_X1 U10627 ( .C1(n9762), .C2(n10101), .A(n9257), .B(n9256), .ZN(n9258)
         );
  OAI21_X1 U10628 ( .B1(n9766), .B2(n9322), .A(n9258), .ZN(P1_U3271) );
  XOR2_X1 U10629 ( .A(n9264), .B(n9259), .Z(n9774) );
  INV_X1 U10630 ( .A(n9260), .ZN(n9262) );
  OAI21_X1 U10631 ( .B1(n9277), .B2(n9262), .A(n9261), .ZN(n9263) );
  XOR2_X1 U10632 ( .A(n9264), .B(n9263), .Z(n9772) );
  INV_X1 U10633 ( .A(n9279), .ZN(n9266) );
  OAI211_X1 U10634 ( .C1(n9266), .C2(n9770), .A(n10097), .B(n9265), .ZN(n9769)
         );
  NAND2_X1 U10635 ( .A1(n9344), .A2(n9767), .ZN(n9269) );
  AOI22_X1 U10636 ( .A1(n4495), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9267), .B2(
        n10092), .ZN(n9268) );
  OAI211_X1 U10637 ( .C1(n9270), .C2(n9348), .A(n9269), .B(n9268), .ZN(n9271)
         );
  AOI21_X1 U10638 ( .B1(n9272), .B2(n10090), .A(n9271), .ZN(n9273) );
  OAI21_X1 U10639 ( .B1(n9769), .B2(n9327), .A(n9273), .ZN(n9274) );
  AOI21_X1 U10640 ( .B1(n9772), .B2(n9301), .A(n9274), .ZN(n9275) );
  OAI21_X1 U10641 ( .B1(n9774), .B2(n9322), .A(n9275), .ZN(P1_U3272) );
  XOR2_X1 U10642 ( .A(n9278), .B(n9276), .Z(n9782) );
  XOR2_X1 U10643 ( .A(n9277), .B(n9278), .Z(n9780) );
  OAI211_X1 U10644 ( .C1(n9292), .C2(n9778), .A(n10097), .B(n9279), .ZN(n9777)
         );
  NAND2_X1 U10645 ( .A1(n9344), .A2(n9775), .ZN(n9282) );
  AOI22_X1 U10646 ( .A1(n4495), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9280), .B2(
        n10092), .ZN(n9281) );
  OAI211_X1 U10647 ( .C1(n9283), .C2(n9348), .A(n9282), .B(n9281), .ZN(n9284)
         );
  AOI21_X1 U10648 ( .B1(n9285), .B2(n10090), .A(n9284), .ZN(n9286) );
  OAI21_X1 U10649 ( .B1(n9777), .B2(n9327), .A(n9286), .ZN(n9287) );
  AOI21_X1 U10650 ( .B1(n9780), .B2(n9301), .A(n9287), .ZN(n9288) );
  OAI21_X1 U10651 ( .B1(n9782), .B2(n9322), .A(n9288), .ZN(P1_U3273) );
  XOR2_X1 U10652 ( .A(n9289), .B(n9290), .Z(n9791) );
  XNOR2_X1 U10653 ( .A(n9291), .B(n9290), .ZN(n9789) );
  INV_X1 U10654 ( .A(n9292), .ZN(n9293) );
  OAI211_X1 U10655 ( .C1(n9787), .C2(n9877), .A(n9293), .B(n10097), .ZN(n9786)
         );
  NAND2_X1 U10656 ( .A1(n9344), .A2(n9783), .ZN(n9296) );
  AOI22_X1 U10657 ( .A1(n4495), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9294), .B2(
        n10092), .ZN(n9295) );
  OAI211_X1 U10658 ( .C1(n9889), .C2(n9348), .A(n9296), .B(n9295), .ZN(n9297)
         );
  AOI21_X1 U10659 ( .B1(n9298), .B2(n10090), .A(n9297), .ZN(n9299) );
  OAI21_X1 U10660 ( .B1(n9786), .B2(n9327), .A(n9299), .ZN(n9300) );
  AOI21_X1 U10661 ( .B1(n9789), .B2(n9301), .A(n9300), .ZN(n9302) );
  OAI21_X1 U10662 ( .B1(n9791), .B2(n9322), .A(n9302), .ZN(P1_U3274) );
  XNOR2_X1 U10663 ( .A(n9303), .B(n9304), .ZN(n9894) );
  XOR2_X1 U10664 ( .A(n9305), .B(n9304), .Z(n9896) );
  NAND2_X1 U10665 ( .A1(n9896), .A2(n10102), .ZN(n9316) );
  AOI211_X1 U10666 ( .C1(n9892), .C2(n9326), .A(n9339), .B(n9879), .ZN(n9890)
         );
  NOR2_X1 U10667 ( .A1(n9348), .A2(n9908), .ZN(n9311) );
  OAI22_X1 U10668 ( .A1(n9309), .A2(n9308), .B1(n9307), .B2(n9306), .ZN(n9310)
         );
  AOI211_X1 U10669 ( .C1(n9344), .C2(n9784), .A(n9311), .B(n9310), .ZN(n9312)
         );
  OAI21_X1 U10670 ( .B1(n9313), .B2(n9341), .A(n9312), .ZN(n9314) );
  AOI21_X1 U10671 ( .B1(n9890), .B2(n10101), .A(n9314), .ZN(n9315) );
  OAI211_X1 U10672 ( .C1(n9894), .C2(n9353), .A(n9316), .B(n9315), .ZN(
        P1_U3276) );
  XNOR2_X1 U10673 ( .A(n9317), .B(n9318), .ZN(n9905) );
  INV_X1 U10674 ( .A(n9905), .ZN(n9333) );
  NOR2_X1 U10675 ( .A1(n9320), .A2(n9319), .ZN(n9902) );
  INV_X1 U10676 ( .A(n9321), .ZN(n9901) );
  OR3_X1 U10677 ( .A1(n9902), .A2(n9901), .A3(n9322), .ZN(n9332) );
  NAND2_X1 U10678 ( .A1(n9344), .A2(n9898), .ZN(n9325) );
  AOI22_X1 U10679 ( .A1(n4495), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9323), .B2(
        n10092), .ZN(n9324) );
  OAI211_X1 U10680 ( .C1(n10237), .C2(n9348), .A(n9325), .B(n9324), .ZN(n9329)
         );
  OAI211_X1 U10681 ( .C1(n4581), .C2(n4802), .A(n10097), .B(n9326), .ZN(n9900)
         );
  NOR2_X1 U10682 ( .A1(n9900), .A2(n9327), .ZN(n9328) );
  AOI211_X1 U10683 ( .C1(n10090), .C2(n9330), .A(n9329), .B(n9328), .ZN(n9331)
         );
  OAI211_X1 U10684 ( .C1(n9333), .C2(n9353), .A(n9332), .B(n9331), .ZN(
        P1_U3277) );
  INV_X1 U10685 ( .A(n9334), .ZN(n9335) );
  AOI21_X1 U10686 ( .B1(n9337), .B2(n9336), .A(n9335), .ZN(n9913) );
  XNOR2_X1 U10687 ( .A(n9338), .B(n9337), .ZN(n9915) );
  NAND2_X1 U10688 ( .A1(n9915), .A2(n10102), .ZN(n9352) );
  AOI211_X1 U10689 ( .C1(n9911), .C2(n9340), .A(n9339), .B(n4581), .ZN(n9909)
         );
  NOR2_X1 U10690 ( .A1(n9342), .A2(n9341), .ZN(n9350) );
  NAND2_X1 U10691 ( .A1(n9344), .A2(n9343), .ZN(n9347) );
  AOI22_X1 U10692 ( .A1(n4495), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9345), .B2(
        n10092), .ZN(n9346) );
  OAI211_X1 U10693 ( .C1(n9907), .C2(n9348), .A(n9347), .B(n9346), .ZN(n9349)
         );
  AOI211_X1 U10694 ( .C1(n9909), .C2(n10101), .A(n9350), .B(n9349), .ZN(n9351)
         );
  OAI211_X1 U10695 ( .C1(n9913), .C2(n9353), .A(n9352), .B(n9351), .ZN(
        P1_U3278) );
  OAI211_X1 U10696 ( .C1(n9355), .C2(n10227), .A(n9354), .B(n9709), .ZN(n9792)
         );
  MUX2_X1 U10697 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9792), .S(n10274), .Z(
        P1_U3553) );
  AOI22_X1 U10698 ( .A1(n6878), .A2(keyinput11), .B1(keyinput104), .B2(n9357), 
        .ZN(n9356) );
  OAI221_X1 U10699 ( .B1(n6878), .B2(keyinput11), .C1(n9357), .C2(keyinput104), 
        .A(n9356), .ZN(n9365) );
  INV_X1 U10700 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10111) );
  AOI22_X1 U10701 ( .A1(n8339), .A2(keyinput95), .B1(keyinput33), .B2(n10111), 
        .ZN(n9358) );
  OAI221_X1 U10702 ( .B1(n8339), .B2(keyinput95), .C1(n10111), .C2(keyinput33), 
        .A(n9358), .ZN(n9364) );
  AOI22_X1 U10703 ( .A1(n9683), .A2(keyinput20), .B1(keyinput114), .B2(n9603), 
        .ZN(n9359) );
  OAI221_X1 U10704 ( .B1(n9683), .B2(keyinput20), .C1(n9603), .C2(keyinput114), 
        .A(n9359), .ZN(n9363) );
  INV_X1 U10705 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9361) );
  AOI22_X1 U10706 ( .A1(n9361), .A2(keyinput81), .B1(n9906), .B2(keyinput80), 
        .ZN(n9360) );
  OAI221_X1 U10707 ( .B1(n9361), .B2(keyinput81), .C1(n9906), .C2(keyinput80), 
        .A(n9360), .ZN(n9362) );
  OR4_X1 U10708 ( .A1(n9365), .A2(n9364), .A3(n9363), .A4(n9362), .ZN(n9380)
         );
  AOI22_X1 U10709 ( .A1(n9367), .A2(keyinput28), .B1(keyinput15), .B2(n6110), 
        .ZN(n9366) );
  OAI221_X1 U10710 ( .B1(n9367), .B2(keyinput28), .C1(n6110), .C2(keyinput15), 
        .A(n9366), .ZN(n9379) );
  OAI22_X1 U10711 ( .A1(P1_D_REG_20__SCAN_IN), .A2(keyinput58), .B1(keyinput22), .B2(P1_ADDR_REG_14__SCAN_IN), .ZN(n9368) );
  AOI221_X1 U10712 ( .B1(P1_D_REG_20__SCAN_IN), .B2(keyinput58), .C1(
        P1_ADDR_REG_14__SCAN_IN), .C2(keyinput22), .A(n9368), .ZN(n9375) );
  OAI22_X1 U10713 ( .A1(P2_D_REG_22__SCAN_IN), .A2(keyinput116), .B1(keyinput7), .B2(P1_D_REG_10__SCAN_IN), .ZN(n9369) );
  AOI221_X1 U10714 ( .B1(P2_D_REG_22__SCAN_IN), .B2(keyinput116), .C1(
        P1_D_REG_10__SCAN_IN), .C2(keyinput7), .A(n9369), .ZN(n9374) );
  OAI22_X1 U10715 ( .A1(P1_REG1_REG_25__SCAN_IN), .A2(keyinput62), .B1(
        P2_ADDR_REG_13__SCAN_IN), .B2(keyinput61), .ZN(n9370) );
  AOI221_X1 U10716 ( .B1(P1_REG1_REG_25__SCAN_IN), .B2(keyinput62), .C1(
        keyinput61), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n9370), .ZN(n9373) );
  OAI22_X1 U10717 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput49), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(keyinput40), .ZN(n9371) );
  AOI221_X1 U10718 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput49), .C1(
        keyinput40), .C2(P1_DATAO_REG_29__SCAN_IN), .A(n9371), .ZN(n9372) );
  NAND4_X1 U10719 ( .A1(n9375), .A2(n9374), .A3(n9373), .A4(n9372), .ZN(n9378)
         );
  INV_X1 U10720 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10250) );
  AOI22_X1 U10721 ( .A1(n10250), .A2(keyinput6), .B1(keyinput51), .B2(n9676), 
        .ZN(n9376) );
  OAI221_X1 U10722 ( .B1(n10250), .B2(keyinput6), .C1(n9676), .C2(keyinput51), 
        .A(n9376), .ZN(n9377) );
  NOR4_X1 U10723 ( .A1(n9380), .A2(n9379), .A3(n9378), .A4(n9377), .ZN(n9455)
         );
  OAI22_X1 U10724 ( .A1(n7924), .A2(keyinput66), .B1(n9601), .B2(keyinput70), 
        .ZN(n9381) );
  AOI221_X1 U10725 ( .B1(n7924), .B2(keyinput66), .C1(keyinput70), .C2(n9601), 
        .A(n9381), .ZN(n9454) );
  XOR2_X1 U10726 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput17), .Z(n9391) );
  XNOR2_X1 U10727 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput57), .ZN(n9385) );
  XNOR2_X1 U10728 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput103), .ZN(n9384)
         );
  XNOR2_X1 U10729 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput124), .ZN(n9383) );
  XNOR2_X1 U10730 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(keyinput78), .ZN(n9382) );
  NAND4_X1 U10731 ( .A1(n9385), .A2(n9384), .A3(n9383), .A4(n9382), .ZN(n9390)
         );
  XNOR2_X1 U10732 ( .A(n9386), .B(keyinput90), .ZN(n9389) );
  INV_X1 U10733 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9387) );
  XNOR2_X1 U10734 ( .A(keyinput107), .B(n9387), .ZN(n9388) );
  NOR4_X1 U10735 ( .A1(n9391), .A2(n9390), .A3(n9389), .A4(n9388), .ZN(n9393)
         );
  INV_X1 U10736 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10109) );
  XOR2_X1 U10737 ( .A(keyinput68), .B(n10109), .Z(n9392) );
  NAND2_X1 U10738 ( .A1(n9393), .A2(n9392), .ZN(n9421) );
  OAI22_X1 U10739 ( .A1(P2_REG1_REG_24__SCAN_IN), .A2(keyinput31), .B1(
        P2_ADDR_REG_4__SCAN_IN), .B2(keyinput54), .ZN(n9394) );
  AOI221_X1 U10740 ( .B1(P2_REG1_REG_24__SCAN_IN), .B2(keyinput31), .C1(
        keyinput54), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n9394), .ZN(n9401) );
  OAI22_X1 U10741 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(keyinput63), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(keyinput79), .ZN(n9395) );
  AOI221_X1 U10742 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(keyinput63), .C1(
        keyinput79), .C2(P2_REG3_REG_14__SCAN_IN), .A(n9395), .ZN(n9400) );
  OAI22_X1 U10743 ( .A1(P1_REG1_REG_28__SCAN_IN), .A2(keyinput18), .B1(
        P1_REG0_REG_27__SCAN_IN), .B2(keyinput36), .ZN(n9396) );
  AOI221_X1 U10744 ( .B1(P1_REG1_REG_28__SCAN_IN), .B2(keyinput18), .C1(
        keyinput36), .C2(P1_REG0_REG_27__SCAN_IN), .A(n9396), .ZN(n9399) );
  OAI22_X1 U10745 ( .A1(P2_REG1_REG_23__SCAN_IN), .A2(keyinput74), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(keyinput53), .ZN(n9397) );
  AOI221_X1 U10746 ( .B1(P2_REG1_REG_23__SCAN_IN), .B2(keyinput74), .C1(
        keyinput53), .C2(P1_DATAO_REG_30__SCAN_IN), .A(n9397), .ZN(n9398) );
  NAND4_X1 U10747 ( .A1(n9401), .A2(n9400), .A3(n9399), .A4(n9398), .ZN(n9420)
         );
  OAI22_X1 U10748 ( .A1(P2_REG2_REG_3__SCAN_IN), .A2(keyinput1), .B1(
        keyinput76), .B2(P1_D_REG_2__SCAN_IN), .ZN(n9402) );
  AOI221_X1 U10749 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(keyinput1), .C1(
        P1_D_REG_2__SCAN_IN), .C2(keyinput76), .A(n9402), .ZN(n9409) );
  OAI22_X1 U10750 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput34), .B1(
        keyinput82), .B2(P1_ADDR_REG_18__SCAN_IN), .ZN(n9403) );
  AOI221_X1 U10751 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput34), .C1(
        P1_ADDR_REG_18__SCAN_IN), .C2(keyinput82), .A(n9403), .ZN(n9408) );
  OAI22_X1 U10752 ( .A1(P2_D_REG_30__SCAN_IN), .A2(keyinput60), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(keyinput14), .ZN(n9404) );
  AOI221_X1 U10753 ( .B1(P2_D_REG_30__SCAN_IN), .B2(keyinput60), .C1(
        keyinput14), .C2(P2_DATAO_REG_22__SCAN_IN), .A(n9404), .ZN(n9407) );
  OAI22_X1 U10754 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(keyinput113), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(keyinput71), .ZN(n9405) );
  AOI221_X1 U10755 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(keyinput113), .C1(
        keyinput71), .C2(P1_DATAO_REG_31__SCAN_IN), .A(n9405), .ZN(n9406) );
  NAND4_X1 U10756 ( .A1(n9409), .A2(n9408), .A3(n9407), .A4(n9406), .ZN(n9419)
         );
  OAI22_X1 U10757 ( .A1(P2_REG0_REG_6__SCAN_IN), .A2(keyinput30), .B1(
        keyinput110), .B2(P1_REG1_REG_14__SCAN_IN), .ZN(n9410) );
  AOI221_X1 U10758 ( .B1(P2_REG0_REG_6__SCAN_IN), .B2(keyinput30), .C1(
        P1_REG1_REG_14__SCAN_IN), .C2(keyinput110), .A(n9410), .ZN(n9417) );
  OAI22_X1 U10759 ( .A1(P2_REG0_REG_17__SCAN_IN), .A2(keyinput19), .B1(
        keyinput24), .B2(P2_REG0_REG_14__SCAN_IN), .ZN(n9411) );
  AOI221_X1 U10760 ( .B1(P2_REG0_REG_17__SCAN_IN), .B2(keyinput19), .C1(
        P2_REG0_REG_14__SCAN_IN), .C2(keyinput24), .A(n9411), .ZN(n9416) );
  OAI22_X1 U10761 ( .A1(SI_4_), .A2(keyinput10), .B1(P2_REG1_REG_0__SCAN_IN), 
        .B2(keyinput16), .ZN(n9412) );
  AOI221_X1 U10762 ( .B1(SI_4_), .B2(keyinput10), .C1(keyinput16), .C2(
        P2_REG1_REG_0__SCAN_IN), .A(n9412), .ZN(n9415) );
  OAI22_X1 U10763 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(keyinput84), .B1(
        P1_REG2_REG_13__SCAN_IN), .B2(keyinput56), .ZN(n9413) );
  AOI221_X1 U10764 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(keyinput84), .C1(
        keyinput56), .C2(P1_REG2_REG_13__SCAN_IN), .A(n9413), .ZN(n9414) );
  NAND4_X1 U10765 ( .A1(n9417), .A2(n9416), .A3(n9415), .A4(n9414), .ZN(n9418)
         );
  NOR4_X1 U10766 ( .A1(n9421), .A2(n9420), .A3(n9419), .A4(n9418), .ZN(n9453)
         );
  OAI22_X1 U10767 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(keyinput43), .B1(
        keyinput106), .B2(P1_REG0_REG_10__SCAN_IN), .ZN(n9422) );
  AOI221_X1 U10768 ( .B1(P2_DATAO_REG_14__SCAN_IN), .B2(keyinput43), .C1(
        P1_REG0_REG_10__SCAN_IN), .C2(keyinput106), .A(n9422), .ZN(n9429) );
  OAI22_X1 U10769 ( .A1(P2_REG1_REG_27__SCAN_IN), .A2(keyinput97), .B1(
        P2_REG2_REG_17__SCAN_IN), .B2(keyinput9), .ZN(n9423) );
  AOI221_X1 U10770 ( .B1(P2_REG1_REG_27__SCAN_IN), .B2(keyinput97), .C1(
        keyinput9), .C2(P2_REG2_REG_17__SCAN_IN), .A(n9423), .ZN(n9428) );
  OAI22_X1 U10771 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(keyinput2), .B1(
        P1_REG2_REG_9__SCAN_IN), .B2(keyinput42), .ZN(n9424) );
  AOI221_X1 U10772 ( .B1(P1_REG3_REG_27__SCAN_IN), .B2(keyinput2), .C1(
        keyinput42), .C2(P1_REG2_REG_9__SCAN_IN), .A(n9424), .ZN(n9427) );
  OAI22_X1 U10773 ( .A1(P2_D_REG_25__SCAN_IN), .A2(keyinput65), .B1(keyinput46), .B2(P2_REG1_REG_28__SCAN_IN), .ZN(n9425) );
  AOI221_X1 U10774 ( .B1(P2_D_REG_25__SCAN_IN), .B2(keyinput65), .C1(
        P2_REG1_REG_28__SCAN_IN), .C2(keyinput46), .A(n9425), .ZN(n9426) );
  NAND4_X1 U10775 ( .A1(n9429), .A2(n9428), .A3(n9427), .A4(n9426), .ZN(n9451)
         );
  OAI22_X1 U10776 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput117), .B1(
        keyinput91), .B2(P2_ADDR_REG_17__SCAN_IN), .ZN(n9430) );
  AOI221_X1 U10777 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput117), .C1(
        P2_ADDR_REG_17__SCAN_IN), .C2(keyinput91), .A(n9430), .ZN(n9437) );
  OAI22_X1 U10778 ( .A1(P2_REG2_REG_27__SCAN_IN), .A2(keyinput127), .B1(
        P1_IR_REG_6__SCAN_IN), .B2(keyinput88), .ZN(n9431) );
  AOI221_X1 U10779 ( .B1(P2_REG2_REG_27__SCAN_IN), .B2(keyinput127), .C1(
        keyinput88), .C2(P1_IR_REG_6__SCAN_IN), .A(n9431), .ZN(n9436) );
  OAI22_X1 U10780 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(keyinput12), .B1(
        keyinput120), .B2(P1_ADDR_REG_8__SCAN_IN), .ZN(n9432) );
  AOI221_X1 U10781 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(keyinput12), .C1(
        P1_ADDR_REG_8__SCAN_IN), .C2(keyinput120), .A(n9432), .ZN(n9435) );
  OAI22_X1 U10782 ( .A1(P1_REG0_REG_18__SCAN_IN), .A2(keyinput26), .B1(
        keyinput67), .B2(P1_REG2_REG_14__SCAN_IN), .ZN(n9433) );
  AOI221_X1 U10783 ( .B1(P1_REG0_REG_18__SCAN_IN), .B2(keyinput26), .C1(
        P1_REG2_REG_14__SCAN_IN), .C2(keyinput67), .A(n9433), .ZN(n9434) );
  NAND4_X1 U10784 ( .A1(n9437), .A2(n9436), .A3(n9435), .A4(n9434), .ZN(n9450)
         );
  OAI22_X1 U10785 ( .A1(P2_D_REG_13__SCAN_IN), .A2(keyinput52), .B1(
        P2_REG3_REG_23__SCAN_IN), .B2(keyinput92), .ZN(n9438) );
  AOI221_X1 U10786 ( .B1(P2_D_REG_13__SCAN_IN), .B2(keyinput52), .C1(
        keyinput92), .C2(P2_REG3_REG_23__SCAN_IN), .A(n9438), .ZN(n9445) );
  OAI22_X1 U10787 ( .A1(P2_IR_REG_30__SCAN_IN), .A2(keyinput21), .B1(
        P2_REG0_REG_11__SCAN_IN), .B2(keyinput118), .ZN(n9439) );
  AOI221_X1 U10788 ( .B1(P2_IR_REG_30__SCAN_IN), .B2(keyinput21), .C1(
        keyinput118), .C2(P2_REG0_REG_11__SCAN_IN), .A(n9439), .ZN(n9444) );
  OAI22_X1 U10789 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(keyinput41), .B1(
        keyinput112), .B2(P1_D_REG_12__SCAN_IN), .ZN(n9440) );
  AOI221_X1 U10790 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(keyinput41), .C1(
        P1_D_REG_12__SCAN_IN), .C2(keyinput112), .A(n9440), .ZN(n9443) );
  OAI22_X1 U10791 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput94), .B1(
        keyinput29), .B2(P1_REG0_REG_11__SCAN_IN), .ZN(n9441) );
  AOI221_X1 U10792 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput94), .C1(
        P1_REG0_REG_11__SCAN_IN), .C2(keyinput29), .A(n9441), .ZN(n9442) );
  NAND4_X1 U10793 ( .A1(n9445), .A2(n9444), .A3(n9443), .A4(n9442), .ZN(n9449)
         );
  XOR2_X1 U10794 ( .A(keyinput3), .B(n9679), .Z(n9447) );
  INV_X1 U10795 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10106) );
  XOR2_X1 U10796 ( .A(keyinput35), .B(n10106), .Z(n9446) );
  NAND2_X1 U10797 ( .A1(n9447), .A2(n9446), .ZN(n9448) );
  NOR4_X1 U10798 ( .A1(n9451), .A2(n9450), .A3(n9449), .A4(n9448), .ZN(n9452)
         );
  AND4_X1 U10799 ( .A1(n9455), .A2(n9454), .A3(n9453), .A4(n9452), .ZN(n9492)
         );
  OAI22_X1 U10800 ( .A1(n9457), .A2(keyinput109), .B1(n9640), .B2(keyinput23), 
        .ZN(n9456) );
  AOI221_X1 U10801 ( .B1(n9457), .B2(keyinput109), .C1(keyinput23), .C2(n9640), 
        .A(n9456), .ZN(n9491) );
  OAI22_X1 U10802 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput77), .B1(
        keyinput5), .B2(SI_1_), .ZN(n9458) );
  AOI221_X1 U10803 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput77), .C1(SI_1_), 
        .C2(keyinput5), .A(n9458), .ZN(n9490) );
  INV_X1 U10804 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10105) );
  AOI22_X1 U10805 ( .A1(n10105), .A2(keyinput98), .B1(n5980), .B2(keyinput59), 
        .ZN(n9459) );
  OAI221_X1 U10806 ( .B1(n10105), .B2(keyinput98), .C1(n5980), .C2(keyinput59), 
        .A(n9459), .ZN(n9467) );
  AOI22_X1 U10807 ( .A1(n9462), .A2(keyinput32), .B1(n9461), .B2(keyinput126), 
        .ZN(n9460) );
  OAI221_X1 U10808 ( .B1(n9462), .B2(keyinput32), .C1(n9461), .C2(keyinput126), 
        .A(n9460), .ZN(n9466) );
  XNOR2_X1 U10809 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput48), .ZN(n9464) );
  XNOR2_X1 U10810 ( .A(keyinput96), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9463) );
  NAND2_X1 U10811 ( .A1(n9464), .A2(n9463), .ZN(n9465) );
  NOR3_X1 U10812 ( .A1(n9467), .A2(n9466), .A3(n9465), .ZN(n9488) );
  INV_X1 U10813 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10233) );
  AOI22_X1 U10814 ( .A1(n9469), .A2(keyinput86), .B1(keyinput99), .B2(n10233), 
        .ZN(n9468) );
  OAI221_X1 U10815 ( .B1(n9469), .B2(keyinput86), .C1(n10233), .C2(keyinput99), 
        .A(n9468), .ZN(n9473) );
  AOI22_X1 U10816 ( .A1(n9471), .A2(keyinput119), .B1(n9600), .B2(keyinput93), 
        .ZN(n9470) );
  OAI221_X1 U10817 ( .B1(n9471), .B2(keyinput119), .C1(n9600), .C2(keyinput93), 
        .A(n9470), .ZN(n9472) );
  NOR2_X1 U10818 ( .A1(n9473), .A2(n9472), .ZN(n9487) );
  AOI22_X1 U10819 ( .A1(n9630), .A2(keyinput38), .B1(n6619), .B2(keyinput89), 
        .ZN(n9474) );
  OAI221_X1 U10820 ( .B1(n9630), .B2(keyinput38), .C1(n6619), .C2(keyinput89), 
        .A(n9474), .ZN(n9477) );
  AOI22_X1 U10821 ( .A1(n9836), .A2(keyinput4), .B1(n6411), .B2(keyinput69), 
        .ZN(n9475) );
  OAI221_X1 U10822 ( .B1(n9836), .B2(keyinput4), .C1(n6411), .C2(keyinput69), 
        .A(n9475), .ZN(n9476) );
  NOR2_X1 U10823 ( .A1(n9477), .A2(n9476), .ZN(n9486) );
  AOI22_X1 U10824 ( .A1(n10399), .A2(keyinput75), .B1(n7667), .B2(keyinput8), 
        .ZN(n9478) );
  OAI221_X1 U10825 ( .B1(n10399), .B2(keyinput75), .C1(n7667), .C2(keyinput8), 
        .A(n9478), .ZN(n9484) );
  XNOR2_X1 U10826 ( .A(P2_REG1_REG_1__SCAN_IN), .B(keyinput73), .ZN(n9482) );
  XNOR2_X1 U10827 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput0), .ZN(n9481) );
  XNOR2_X1 U10828 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(keyinput45), .ZN(n9480) );
  XNOR2_X1 U10829 ( .A(keyinput121), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9479) );
  NAND4_X1 U10830 ( .A1(n9482), .A2(n9481), .A3(n9480), .A4(n9479), .ZN(n9483)
         );
  NOR2_X1 U10831 ( .A1(n9484), .A2(n9483), .ZN(n9485) );
  AND4_X1 U10832 ( .A1(n9488), .A2(n9487), .A3(n9486), .A4(n9485), .ZN(n9489)
         );
  AND4_X1 U10833 ( .A1(n9492), .A2(n9491), .A3(n9490), .A4(n9489), .ZN(n9526)
         );
  INV_X1 U10834 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9494) );
  AOI22_X1 U10835 ( .A1(n9665), .A2(keyinput115), .B1(n9494), .B2(keyinput27), 
        .ZN(n9493) );
  OAI221_X1 U10836 ( .B1(n9665), .B2(keyinput115), .C1(n9494), .C2(keyinput27), 
        .A(n9493), .ZN(n9504) );
  AOI22_X1 U10837 ( .A1(n9615), .A2(keyinput55), .B1(n9496), .B2(keyinput100), 
        .ZN(n9495) );
  OAI221_X1 U10838 ( .B1(n9615), .B2(keyinput55), .C1(n9496), .C2(keyinput100), 
        .A(n9495), .ZN(n9503) );
  AOI22_X1 U10839 ( .A1(n9499), .A2(keyinput39), .B1(keyinput47), .B2(n9498), 
        .ZN(n9497) );
  OAI221_X1 U10840 ( .B1(n9499), .B2(keyinput39), .C1(n9498), .C2(keyinput47), 
        .A(n9497), .ZN(n9502) );
  AOI22_X1 U10841 ( .A1(n10258), .A2(keyinput87), .B1(n9654), .B2(keyinput64), 
        .ZN(n9500) );
  OAI221_X1 U10842 ( .B1(n10258), .B2(keyinput87), .C1(n9654), .C2(keyinput64), 
        .A(n9500), .ZN(n9501) );
  NOR4_X1 U10843 ( .A1(n9504), .A2(n9503), .A3(n9502), .A4(n9501), .ZN(n9525)
         );
  INV_X1 U10844 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10108) );
  AOI22_X1 U10845 ( .A1(n9668), .A2(keyinput123), .B1(keyinput72), .B2(n10108), 
        .ZN(n9505) );
  OAI221_X1 U10846 ( .B1(n9668), .B2(keyinput123), .C1(n10108), .C2(keyinput72), .A(n9505), .ZN(n9513) );
  INV_X1 U10847 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9963) );
  AOI22_X1 U10848 ( .A1(n6511), .A2(keyinput101), .B1(keyinput102), .B2(n9963), 
        .ZN(n9506) );
  OAI221_X1 U10849 ( .B1(n6511), .B2(keyinput101), .C1(n9963), .C2(keyinput102), .A(n9506), .ZN(n9512) );
  INV_X1 U10850 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9508) );
  INV_X1 U10851 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10112) );
  AOI22_X1 U10852 ( .A1(n9508), .A2(keyinput122), .B1(n10112), .B2(keyinput105), .ZN(n9507) );
  OAI221_X1 U10853 ( .B1(n9508), .B2(keyinput122), .C1(n10112), .C2(
        keyinput105), .A(n9507), .ZN(n9511) );
  AOI22_X1 U10854 ( .A1(n7112), .A2(keyinput37), .B1(n5988), .B2(keyinput25), 
        .ZN(n9509) );
  OAI221_X1 U10855 ( .B1(n7112), .B2(keyinput37), .C1(n5988), .C2(keyinput25), 
        .A(n9509), .ZN(n9510) );
  NOR4_X1 U10856 ( .A1(n9513), .A2(n9512), .A3(n9511), .A4(n9510), .ZN(n9524)
         );
  AOI22_X1 U10857 ( .A1(n9636), .A2(keyinput111), .B1(keyinput108), .B2(n10371), .ZN(n9514) );
  OAI221_X1 U10858 ( .B1(n9636), .B2(keyinput111), .C1(n10371), .C2(
        keyinput108), .A(n9514), .ZN(n9522) );
  AOI22_X1 U10859 ( .A1(n5146), .A2(keyinput44), .B1(keyinput85), .B2(n10394), 
        .ZN(n9515) );
  OAI221_X1 U10860 ( .B1(n5146), .B2(keyinput44), .C1(n10394), .C2(keyinput85), 
        .A(n9515), .ZN(n9521) );
  AOI22_X1 U10861 ( .A1(n7482), .A2(keyinput50), .B1(n9677), .B2(keyinput125), 
        .ZN(n9516) );
  OAI221_X1 U10862 ( .B1(n7482), .B2(keyinput50), .C1(n9677), .C2(keyinput125), 
        .A(n9516), .ZN(n9520) );
  AOI22_X1 U10863 ( .A1(n9518), .A2(keyinput83), .B1(n10024), .B2(keyinput13), 
        .ZN(n9517) );
  OAI221_X1 U10864 ( .B1(n9518), .B2(keyinput83), .C1(n10024), .C2(keyinput13), 
        .A(n9517), .ZN(n9519) );
  NOR4_X1 U10865 ( .A1(n9522), .A2(n9521), .A3(n9520), .A4(n9519), .ZN(n9523)
         );
  NAND4_X1 U10866 ( .A1(n9526), .A2(n9525), .A3(n9524), .A4(n9523), .ZN(n9708)
         );
  AOI22_X1 U10867 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput218), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(keyinput144), .ZN(n9527) );
  OAI221_X1 U10868 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput218), .C1(
        P2_REG1_REG_0__SCAN_IN), .C2(keyinput144), .A(n9527), .ZN(n9534) );
  AOI22_X1 U10869 ( .A1(P2_REG2_REG_31__SCAN_IN), .A2(keyinput160), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(keyinput169), .ZN(n9528) );
  OAI221_X1 U10870 ( .B1(P2_REG2_REG_31__SCAN_IN), .B2(keyinput160), .C1(
        P2_DATAO_REG_17__SCAN_IN), .C2(keyinput169), .A(n9528), .ZN(n9533) );
  AOI22_X1 U10871 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(keyinput182), .B1(
        P1_REG2_REG_27__SCAN_IN), .B2(keyinput250), .ZN(n9529) );
  OAI221_X1 U10872 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(keyinput182), .C1(
        P1_REG2_REG_27__SCAN_IN), .C2(keyinput250), .A(n9529), .ZN(n9532) );
  AOI22_X1 U10873 ( .A1(P1_REG0_REG_30__SCAN_IN), .A2(keyinput209), .B1(
        P1_IR_REG_30__SCAN_IN), .B2(keyinput172), .ZN(n9530) );
  OAI221_X1 U10874 ( .B1(P1_REG0_REG_30__SCAN_IN), .B2(keyinput209), .C1(
        P1_IR_REG_30__SCAN_IN), .C2(keyinput172), .A(n9530), .ZN(n9531) );
  NOR4_X1 U10875 ( .A1(n9534), .A2(n9533), .A3(n9532), .A4(n9531), .ZN(n9562)
         );
  AOI22_X1 U10876 ( .A1(P2_D_REG_13__SCAN_IN), .A2(keyinput180), .B1(
        P2_IR_REG_23__SCAN_IN), .B2(keyinput153), .ZN(n9535) );
  OAI221_X1 U10877 ( .B1(P2_D_REG_13__SCAN_IN), .B2(keyinput180), .C1(
        P2_IR_REG_23__SCAN_IN), .C2(keyinput153), .A(n9535), .ZN(n9542) );
  AOI22_X1 U10878 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(keyinput187), .B1(
        P2_IR_REG_31__SCAN_IN), .B2(keyinput191), .ZN(n9536) );
  OAI221_X1 U10879 ( .B1(P2_IR_REG_25__SCAN_IN), .B2(keyinput187), .C1(
        P2_IR_REG_31__SCAN_IN), .C2(keyinput191), .A(n9536), .ZN(n9541) );
  AOI22_X1 U10880 ( .A1(SI_6_), .A2(keyinput175), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(keyinput220), .ZN(n9537) );
  OAI221_X1 U10881 ( .B1(SI_6_), .B2(keyinput175), .C1(P2_REG3_REG_23__SCAN_IN), .C2(keyinput220), .A(n9537), .ZN(n9540) );
  AOI22_X1 U10882 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(keyinput181), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(keyinput156), .ZN(n9538) );
  OAI221_X1 U10883 ( .B1(P1_DATAO_REG_30__SCAN_IN), .B2(keyinput181), .C1(
        P1_DATAO_REG_20__SCAN_IN), .C2(keyinput156), .A(n9538), .ZN(n9539) );
  NOR4_X1 U10884 ( .A1(n9542), .A2(n9541), .A3(n9540), .A4(n9539), .ZN(n9561)
         );
  AOI22_X1 U10885 ( .A1(P1_B_REG_SCAN_IN), .A2(keyinput214), .B1(
        P1_IR_REG_1__SCAN_IN), .B2(keyinput249), .ZN(n9543) );
  OAI221_X1 U10886 ( .B1(P1_B_REG_SCAN_IN), .B2(keyinput214), .C1(
        P1_IR_REG_1__SCAN_IN), .C2(keyinput249), .A(n9543), .ZN(n9550) );
  AOI22_X1 U10887 ( .A1(P1_REG1_REG_25__SCAN_IN), .A2(keyinput190), .B1(
        P2_REG3_REG_6__SCAN_IN), .B2(keyinput245), .ZN(n9544) );
  OAI221_X1 U10888 ( .B1(P1_REG1_REG_25__SCAN_IN), .B2(keyinput190), .C1(
        P2_REG3_REG_6__SCAN_IN), .C2(keyinput245), .A(n9544), .ZN(n9549) );
  AOI22_X1 U10889 ( .A1(P1_REG0_REG_11__SCAN_IN), .A2(keyinput157), .B1(
        P2_REG1_REG_27__SCAN_IN), .B2(keyinput225), .ZN(n9545) );
  OAI221_X1 U10890 ( .B1(P1_REG0_REG_11__SCAN_IN), .B2(keyinput157), .C1(
        P2_REG1_REG_27__SCAN_IN), .C2(keyinput225), .A(n9545), .ZN(n9548) );
  AOI22_X1 U10891 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(keyinput235), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(keyinput228), .ZN(n9546) );
  OAI221_X1 U10892 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(keyinput235), .C1(
        P1_DATAO_REG_28__SCAN_IN), .C2(keyinput228), .A(n9546), .ZN(n9547) );
  NOR4_X1 U10893 ( .A1(n9550), .A2(n9549), .A3(n9548), .A4(n9547), .ZN(n9560)
         );
  AOI22_X1 U10894 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput185), .B1(
        P2_REG2_REG_17__SCAN_IN), .B2(keyinput137), .ZN(n9551) );
  OAI221_X1 U10895 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput185), .C1(
        P2_REG2_REG_17__SCAN_IN), .C2(keyinput137), .A(n9551), .ZN(n9558) );
  AOI22_X1 U10896 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(keyinput232), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(keyinput171), .ZN(n9552) );
  OAI221_X1 U10897 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(keyinput232), .C1(
        P2_DATAO_REG_14__SCAN_IN), .C2(keyinput171), .A(n9552), .ZN(n9557) );
  AOI22_X1 U10898 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(keyinput211), .B1(
        P2_REG0_REG_25__SCAN_IN), .B2(keyinput237), .ZN(n9553) );
  OAI221_X1 U10899 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(keyinput211), .C1(
        P2_REG0_REG_25__SCAN_IN), .C2(keyinput237), .A(n9553), .ZN(n9556) );
  AOI22_X1 U10900 ( .A1(P1_REG1_REG_14__SCAN_IN), .A2(keyinput238), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(keyinput162), .ZN(n9554) );
  OAI221_X1 U10901 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(keyinput238), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput162), .A(n9554), .ZN(n9555) );
  NOR4_X1 U10902 ( .A1(n9558), .A2(n9557), .A3(n9556), .A4(n9555), .ZN(n9559)
         );
  NAND4_X1 U10903 ( .A1(n9562), .A2(n9561), .A3(n9560), .A4(n9559), .ZN(n9706)
         );
  AOI22_X1 U10904 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(keyinput216), .B1(
        P2_REG1_REG_7__SCAN_IN), .B2(keyinput139), .ZN(n9563) );
  OAI221_X1 U10905 ( .B1(P1_IR_REG_6__SCAN_IN), .B2(keyinput216), .C1(
        P2_REG1_REG_7__SCAN_IN), .C2(keyinput139), .A(n9563), .ZN(n9570) );
  AOI22_X1 U10906 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(keyinput254), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(keyinput217), .ZN(n9564) );
  OAI221_X1 U10907 ( .B1(P1_REG3_REG_20__SCAN_IN), .B2(keyinput254), .C1(
        P2_REG3_REG_2__SCAN_IN), .C2(keyinput217), .A(n9564), .ZN(n9569) );
  AOI22_X1 U10908 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(keyinput213), .B1(
        P2_REG1_REG_23__SCAN_IN), .B2(keyinput202), .ZN(n9565) );
  OAI221_X1 U10909 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(keyinput213), .C1(
        P2_REG1_REG_23__SCAN_IN), .C2(keyinput202), .A(n9565), .ZN(n9568) );
  AOI22_X1 U10910 ( .A1(P1_REG1_REG_30__SCAN_IN), .A2(keyinput155), .B1(
        P2_REG2_REG_21__SCAN_IN), .B2(keyinput178), .ZN(n9566) );
  OAI221_X1 U10911 ( .B1(P1_REG1_REG_30__SCAN_IN), .B2(keyinput155), .C1(
        P2_REG2_REG_21__SCAN_IN), .C2(keyinput178), .A(n9566), .ZN(n9567) );
  NOR4_X1 U10912 ( .A1(n9570), .A2(n9569), .A3(n9568), .A4(n9567), .ZN(n9598)
         );
  AOI22_X1 U10913 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(keyinput230), .B1(
        P2_REG2_REG_22__SCAN_IN), .B2(keyinput223), .ZN(n9571) );
  OAI221_X1 U10914 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(keyinput230), .C1(
        P2_REG2_REG_22__SCAN_IN), .C2(keyinput223), .A(n9571), .ZN(n9578) );
  AOI22_X1 U10915 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(keyinput210), .B1(
        P2_REG2_REG_27__SCAN_IN), .B2(keyinput255), .ZN(n9572) );
  OAI221_X1 U10916 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(keyinput210), .C1(
        P2_REG2_REG_27__SCAN_IN), .C2(keyinput255), .A(n9572), .ZN(n9577) );
  AOI22_X1 U10917 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(keyinput195), .B1(
        P1_D_REG_12__SCAN_IN), .B2(keyinput240), .ZN(n9573) );
  OAI221_X1 U10918 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(keyinput195), .C1(
        P1_D_REG_12__SCAN_IN), .C2(keyinput240), .A(n9573), .ZN(n9576) );
  AOI22_X1 U10919 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(keyinput199), .B1(SI_4_), .B2(keyinput138), .ZN(n9574) );
  OAI221_X1 U10920 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(keyinput199), .C1(
        SI_4_), .C2(keyinput138), .A(n9574), .ZN(n9575) );
  NOR4_X1 U10921 ( .A1(n9578), .A2(n9577), .A3(n9576), .A4(n9575), .ZN(n9597)
         );
  AOI22_X1 U10922 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(keyinput132), .B1(
        P1_REG2_REG_9__SCAN_IN), .B2(keyinput170), .ZN(n9579) );
  OAI221_X1 U10923 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(keyinput132), .C1(
        P1_REG2_REG_9__SCAN_IN), .C2(keyinput170), .A(n9579), .ZN(n9586) );
  AOI22_X1 U10924 ( .A1(SI_31_), .A2(keyinput136), .B1(P2_REG2_REG_11__SCAN_IN), .B2(keyinput212), .ZN(n9580) );
  OAI221_X1 U10925 ( .B1(SI_31_), .B2(keyinput136), .C1(
        P2_REG2_REG_11__SCAN_IN), .C2(keyinput212), .A(n9580), .ZN(n9585) );
  AOI22_X1 U10926 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(keyinput248), .B1(
        P1_IR_REG_21__SCAN_IN), .B2(keyinput252), .ZN(n9581) );
  OAI221_X1 U10927 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(keyinput248), .C1(
        P1_IR_REG_21__SCAN_IN), .C2(keyinput252), .A(n9581), .ZN(n9584) );
  AOI22_X1 U10928 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(keyinput203), .B1(
        P1_REG0_REG_13__SCAN_IN), .B2(keyinput227), .ZN(n9582) );
  OAI221_X1 U10929 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(keyinput203), .C1(
        P1_REG0_REG_13__SCAN_IN), .C2(keyinput227), .A(n9582), .ZN(n9583) );
  NOR4_X1 U10930 ( .A1(n9586), .A2(n9585), .A3(n9584), .A4(n9583), .ZN(n9596)
         );
  AOI22_X1 U10931 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(keyinput168), .B1(
        P2_D_REG_30__SCAN_IN), .B2(keyinput188), .ZN(n9587) );
  OAI221_X1 U10932 ( .B1(P1_DATAO_REG_29__SCAN_IN), .B2(keyinput168), .C1(
        P2_D_REG_30__SCAN_IN), .C2(keyinput188), .A(n9587), .ZN(n9594) );
  AOI22_X1 U10933 ( .A1(P1_REG0_REG_14__SCAN_IN), .A2(keyinput134), .B1(
        P2_REG0_REG_6__SCAN_IN), .B2(keyinput158), .ZN(n9588) );
  OAI221_X1 U10934 ( .B1(P1_REG0_REG_14__SCAN_IN), .B2(keyinput134), .C1(
        P2_REG0_REG_6__SCAN_IN), .C2(keyinput158), .A(n9588), .ZN(n9593) );
  AOI22_X1 U10935 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(keyinput219), .B1(SI_1_), 
        .B2(keyinput133), .ZN(n9589) );
  OAI221_X1 U10936 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(keyinput219), .C1(SI_1_), .C2(keyinput133), .A(n9589), .ZN(n9592) );
  INV_X1 U10937 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10110) );
  AOI22_X1 U10938 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(keyinput247), .B1(n10110), .B2(keyinput135), .ZN(n9590) );
  OAI221_X1 U10939 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(keyinput247), .C1(
        n10110), .C2(keyinput135), .A(n9590), .ZN(n9591) );
  NOR4_X1 U10940 ( .A1(n9594), .A2(n9593), .A3(n9592), .A4(n9591), .ZN(n9595)
         );
  NAND4_X1 U10941 ( .A1(n9598), .A2(n9597), .A3(n9596), .A4(n9595), .ZN(n9705)
         );
  AOI22_X1 U10942 ( .A1(n9601), .A2(keyinput198), .B1(n9600), .B2(keyinput221), 
        .ZN(n9599) );
  OAI221_X1 U10943 ( .B1(n9601), .B2(keyinput198), .C1(n9600), .C2(keyinput221), .A(n9599), .ZN(n9610) );
  AOI22_X1 U10944 ( .A1(n9604), .A2(keyinput142), .B1(n9603), .B2(keyinput242), 
        .ZN(n9602) );
  OAI221_X1 U10945 ( .B1(n9604), .B2(keyinput142), .C1(n9603), .C2(keyinput242), .A(n9602), .ZN(n9609) );
  AOI22_X1 U10946 ( .A1(n7156), .A2(keyinput246), .B1(keyinput233), .B2(n10112), .ZN(n9605) );
  OAI221_X1 U10947 ( .B1(n7156), .B2(keyinput246), .C1(n10112), .C2(
        keyinput233), .A(n9605), .ZN(n9608) );
  INV_X1 U10948 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10107) );
  AOI22_X1 U10949 ( .A1(n7407), .A2(keyinput140), .B1(n10107), .B2(keyinput186), .ZN(n9606) );
  OAI221_X1 U10950 ( .B1(n7407), .B2(keyinput140), .C1(n10107), .C2(
        keyinput186), .A(n9606), .ZN(n9607) );
  NOR4_X1 U10951 ( .A1(n9610), .A2(n9609), .A3(n9608), .A4(n9607), .ZN(n9650)
         );
  AOI22_X1 U10952 ( .A1(n9612), .A2(keyinput244), .B1(keyinput236), .B2(n10371), .ZN(n9611) );
  OAI221_X1 U10953 ( .B1(n9612), .B2(keyinput244), .C1(n10371), .C2(
        keyinput236), .A(n9611), .ZN(n9621) );
  AOI22_X1 U10954 ( .A1(n10108), .A2(keyinput200), .B1(n6298), .B2(keyinput149), .ZN(n9613) );
  OAI221_X1 U10955 ( .B1(n10108), .B2(keyinput200), .C1(n6298), .C2(
        keyinput149), .A(n9613), .ZN(n9620) );
  AOI22_X1 U10956 ( .A1(n9616), .A2(keyinput130), .B1(n9615), .B2(keyinput183), 
        .ZN(n9614) );
  OAI221_X1 U10957 ( .B1(n9616), .B2(keyinput130), .C1(n9615), .C2(keyinput183), .A(n9614), .ZN(n9619) );
  AOI22_X1 U10958 ( .A1(n10109), .A2(keyinput196), .B1(n10295), .B2(
        keyinput205), .ZN(n9617) );
  OAI221_X1 U10959 ( .B1(n10109), .B2(keyinput196), .C1(n10295), .C2(
        keyinput205), .A(n9617), .ZN(n9618) );
  NOR4_X1 U10960 ( .A1(n9621), .A2(n9620), .A3(n9619), .A4(n9618), .ZN(n9649)
         );
  AOI22_X1 U10961 ( .A1(n9624), .A2(keyinput146), .B1(n9623), .B2(keyinput152), 
        .ZN(n9622) );
  OAI221_X1 U10962 ( .B1(n9624), .B2(keyinput146), .C1(n9623), .C2(keyinput152), .A(n9622), .ZN(n9627) );
  INV_X1 U10963 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10114) );
  XNOR2_X1 U10964 ( .A(n10114), .B(keyinput204), .ZN(n9626) );
  XNOR2_X1 U10965 ( .A(n4670), .B(keyinput173), .ZN(n9625) );
  OR3_X1 U10966 ( .A1(n9627), .A2(n9626), .A3(n9625), .ZN(n9634) );
  AOI22_X1 U10967 ( .A1(n7121), .A2(keyinput184), .B1(n5563), .B2(keyinput224), 
        .ZN(n9628) );
  OAI221_X1 U10968 ( .B1(n7121), .B2(keyinput184), .C1(n5563), .C2(keyinput224), .A(n9628), .ZN(n9633) );
  AOI22_X1 U10969 ( .A1(n9631), .A2(keyinput164), .B1(keyinput166), .B2(n9630), 
        .ZN(n9629) );
  OAI221_X1 U10970 ( .B1(n9631), .B2(keyinput164), .C1(n9630), .C2(keyinput166), .A(n9629), .ZN(n9632) );
  NOR3_X1 U10971 ( .A1(n9634), .A2(n9633), .A3(n9632), .ZN(n9648) );
  INV_X1 U10972 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10204) );
  AOI22_X1 U10973 ( .A1(n10204), .A2(keyinput234), .B1(n9636), .B2(keyinput239), .ZN(n9635) );
  OAI221_X1 U10974 ( .B1(n10204), .B2(keyinput234), .C1(n9636), .C2(
        keyinput239), .A(n9635), .ZN(n9646) );
  AOI22_X1 U10975 ( .A1(n9638), .A2(keyinput174), .B1(keyinput163), .B2(n10106), .ZN(n9637) );
  OAI221_X1 U10976 ( .B1(n9638), .B2(keyinput174), .C1(n10106), .C2(
        keyinput163), .A(n9637), .ZN(n9645) );
  AOI22_X1 U10977 ( .A1(n9641), .A2(keyinput193), .B1(keyinput151), .B2(n9640), 
        .ZN(n9639) );
  OAI221_X1 U10978 ( .B1(n9641), .B2(keyinput193), .C1(n9640), .C2(keyinput151), .A(n9639), .ZN(n9644) );
  AOI22_X1 U10979 ( .A1(n10298), .A2(keyinput129), .B1(n7924), .B2(keyinput194), .ZN(n9642) );
  OAI221_X1 U10980 ( .B1(n10298), .B2(keyinput129), .C1(n7924), .C2(
        keyinput194), .A(n9642), .ZN(n9643) );
  NOR4_X1 U10981 ( .A1(n9646), .A2(n9645), .A3(n9644), .A4(n9643), .ZN(n9647)
         );
  NAND4_X1 U10982 ( .A1(n9650), .A2(n9649), .A3(n9648), .A4(n9647), .ZN(n9704)
         );
  AOI22_X1 U10983 ( .A1(n9652), .A2(keyinput207), .B1(keyinput241), .B2(n6510), 
        .ZN(n9651) );
  OAI221_X1 U10984 ( .B1(n9652), .B2(keyinput207), .C1(n6510), .C2(keyinput241), .A(n9651), .ZN(n9662) );
  AOI22_X1 U10985 ( .A1(n10024), .A2(keyinput141), .B1(n9654), .B2(keyinput192), .ZN(n9653) );
  OAI221_X1 U10986 ( .B1(n10024), .B2(keyinput141), .C1(n9654), .C2(
        keyinput192), .A(n9653), .ZN(n9661) );
  INV_X1 U10987 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9656) );
  AOI22_X1 U10988 ( .A1(n10111), .A2(keyinput161), .B1(n9656), .B2(keyinput177), .ZN(n9655) );
  OAI221_X1 U10989 ( .B1(n10111), .B2(keyinput161), .C1(n9656), .C2(
        keyinput177), .A(n9655), .ZN(n9660) );
  XNOR2_X1 U10990 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(keyinput167), .ZN(n9658)
         );
  XNOR2_X1 U10991 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput231), .ZN(n9657)
         );
  NAND2_X1 U10992 ( .A1(n9658), .A2(n9657), .ZN(n9659) );
  NOR4_X1 U10993 ( .A1(n9662), .A2(n9661), .A3(n9660), .A4(n9659), .ZN(n9702)
         );
  AOI22_X1 U10994 ( .A1(n10019), .A2(keyinput150), .B1(n6110), .B2(keyinput143), .ZN(n9663) );
  OAI221_X1 U10995 ( .B1(n10019), .B2(keyinput150), .C1(n6110), .C2(
        keyinput143), .A(n9663), .ZN(n9674) );
  AOI22_X1 U10996 ( .A1(n9666), .A2(keyinput189), .B1(keyinput243), .B2(n9665), 
        .ZN(n9664) );
  OAI221_X1 U10997 ( .B1(n9666), .B2(keyinput189), .C1(n9665), .C2(keyinput243), .A(n9664), .ZN(n9673) );
  AOI22_X1 U10998 ( .A1(n6511), .A2(keyinput229), .B1(keyinput251), .B2(n9668), 
        .ZN(n9667) );
  OAI221_X1 U10999 ( .B1(n6511), .B2(keyinput229), .C1(n9668), .C2(keyinput251), .A(n9667), .ZN(n9672) );
  INV_X1 U11000 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9916) );
  XOR2_X1 U11001 ( .A(n9916), .B(keyinput154), .Z(n9670) );
  XNOR2_X1 U11002 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput222), .ZN(n9669) );
  NAND2_X1 U11003 ( .A1(n9670), .A2(n9669), .ZN(n9671) );
  NOR4_X1 U11004 ( .A1(n9674), .A2(n9673), .A3(n9672), .A4(n9671), .ZN(n9701)
         );
  AOI22_X1 U11005 ( .A1(n9677), .A2(keyinput253), .B1(keyinput179), .B2(n9676), 
        .ZN(n9675) );
  OAI221_X1 U11006 ( .B1(n9677), .B2(keyinput253), .C1(n9676), .C2(keyinput179), .A(n9675), .ZN(n9687) );
  AOI22_X1 U11007 ( .A1(n9679), .A2(keyinput131), .B1(n10105), .B2(keyinput226), .ZN(n9678) );
  OAI221_X1 U11008 ( .B1(n9679), .B2(keyinput131), .C1(n10105), .C2(
        keyinput226), .A(n9678), .ZN(n9686) );
  XOR2_X1 U11009 ( .A(n6411), .B(keyinput197), .Z(n9682) );
  XNOR2_X1 U11010 ( .A(P2_REG1_REG_1__SCAN_IN), .B(keyinput201), .ZN(n9681) );
  XNOR2_X1 U11011 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput145), .ZN(n9680) );
  NAND3_X1 U11012 ( .A1(n9682), .A2(n9681), .A3(n9680), .ZN(n9685) );
  XNOR2_X1 U11013 ( .A(n9683), .B(keyinput148), .ZN(n9684) );
  NOR4_X1 U11014 ( .A1(n9687), .A2(n9686), .A3(n9685), .A4(n9684), .ZN(n9700)
         );
  AOI22_X1 U11015 ( .A1(n9906), .A2(keyinput208), .B1(keyinput165), .B2(n7112), 
        .ZN(n9688) );
  OAI221_X1 U11016 ( .B1(n9906), .B2(keyinput208), .C1(n7112), .C2(keyinput165), .A(n9688), .ZN(n9698) );
  AOI22_X1 U11017 ( .A1(n9691), .A2(keyinput147), .B1(n9690), .B2(keyinput159), 
        .ZN(n9689) );
  OAI221_X1 U11018 ( .B1(n9691), .B2(keyinput147), .C1(n9690), .C2(keyinput159), .A(n9689), .ZN(n9697) );
  XOR2_X1 U11019 ( .A(n10258), .B(keyinput215), .Z(n9695) );
  XNOR2_X1 U11020 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(keyinput206), .ZN(n9694)
         );
  XNOR2_X1 U11021 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput176), .ZN(n9693)
         );
  XNOR2_X1 U11022 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput128), .ZN(n9692) );
  NAND4_X1 U11023 ( .A1(n9695), .A2(n9694), .A3(n9693), .A4(n9692), .ZN(n9696)
         );
  NOR3_X1 U11024 ( .A1(n9698), .A2(n9697), .A3(n9696), .ZN(n9699) );
  NAND4_X1 U11025 ( .A1(n9702), .A2(n9701), .A3(n9700), .A4(n9699), .ZN(n9703)
         );
  NOR4_X1 U11026 ( .A1(n9706), .A2(n9705), .A3(n9704), .A4(n9703), .ZN(n9707)
         );
  NOR2_X1 U11027 ( .A1(n9708), .A2(n9707), .ZN(n9713) );
  OAI211_X1 U11028 ( .C1(n9711), .C2(n10227), .A(n9710), .B(n9709), .ZN(n9793)
         );
  XOR2_X1 U11029 ( .A(n9713), .B(n9712), .Z(P1_U3552) );
  NAND2_X1 U11030 ( .A1(n9714), .A2(n10231), .ZN(n9721) );
  OAI22_X1 U11031 ( .A1(n9716), .A2(n10227), .B1(n9715), .B2(n10234), .ZN(
        n9717) );
  NAND2_X1 U11032 ( .A1(n9721), .A2(n9720), .ZN(n9794) );
  MUX2_X1 U11033 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9794), .S(n10274), .Z(
        P1_U3551) );
  OAI22_X1 U11034 ( .A1(n9723), .A2(n10227), .B1(n9722), .B2(n10236), .ZN(
        n9724) );
  NOR2_X1 U11035 ( .A1(n9725), .A2(n9724), .ZN(n9726) );
  OAI211_X1 U11036 ( .C1(n9728), .C2(n10198), .A(n9727), .B(n9726), .ZN(n9795)
         );
  MUX2_X1 U11037 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9795), .S(n10274), .Z(
        P1_U3550) );
  AOI21_X1 U11038 ( .B1(n10241), .B2(n9730), .A(n9729), .ZN(n9731) );
  OAI211_X1 U11039 ( .C1(n9733), .C2(n10198), .A(n9732), .B(n9731), .ZN(n9796)
         );
  MUX2_X1 U11040 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9796), .S(n10274), .Z(
        P1_U3549) );
  NAND2_X1 U11041 ( .A1(n9734), .A2(n10231), .ZN(n9740) );
  AOI22_X1 U11042 ( .A1(n9736), .A2(n10241), .B1(n10191), .B2(n9735), .ZN(
        n9738) );
  NAND4_X1 U11043 ( .A1(n9740), .A2(n9739), .A3(n9738), .A4(n9737), .ZN(n9797)
         );
  MUX2_X1 U11044 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9797), .S(n10274), .Z(
        P1_U3548) );
  AOI22_X1 U11045 ( .A1(n9741), .A2(n10191), .B1(n10194), .B2(n9754), .ZN(
        n9742) );
  OAI21_X1 U11046 ( .B1(n9743), .B2(n10227), .A(n9742), .ZN(n9744) );
  AOI211_X1 U11047 ( .C1(n9746), .C2(n10203), .A(n9745), .B(n9744), .ZN(n9747)
         );
  OAI21_X1 U11048 ( .B1(n9748), .B2(n10198), .A(n9747), .ZN(n9798) );
  MUX2_X1 U11049 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9798), .S(n10274), .Z(
        P1_U3547) );
  AOI21_X1 U11050 ( .B1(n10241), .B2(n9750), .A(n9749), .ZN(n9751) );
  OAI211_X1 U11051 ( .C1(n9753), .C2(n10198), .A(n9752), .B(n9751), .ZN(n9799)
         );
  MUX2_X1 U11052 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9799), .S(n10274), .Z(
        P1_U3546) );
  AOI22_X1 U11053 ( .A1(n9754), .A2(n10191), .B1(n10194), .B2(n9767), .ZN(
        n9755) );
  OAI211_X1 U11054 ( .C1(n9757), .C2(n10227), .A(n9756), .B(n9755), .ZN(n9758)
         );
  AOI21_X1 U11055 ( .B1(n9759), .B2(n10203), .A(n9758), .ZN(n9760) );
  OAI21_X1 U11056 ( .B1(n9761), .B2(n10198), .A(n9760), .ZN(n9800) );
  MUX2_X1 U11057 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9800), .S(n10274), .Z(
        P1_U3545) );
  AOI21_X1 U11058 ( .B1(n10241), .B2(n9763), .A(n9762), .ZN(n9764) );
  OAI211_X1 U11059 ( .C1(n9766), .C2(n10198), .A(n9765), .B(n9764), .ZN(n9801)
         );
  MUX2_X1 U11060 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9801), .S(n10274), .Z(
        P1_U3544) );
  AOI22_X1 U11061 ( .A1(n9767), .A2(n10191), .B1(n10194), .B2(n9783), .ZN(
        n9768) );
  OAI211_X1 U11062 ( .C1(n9770), .C2(n10227), .A(n9769), .B(n9768), .ZN(n9771)
         );
  AOI21_X1 U11063 ( .B1(n9772), .B2(n10203), .A(n9771), .ZN(n9773) );
  OAI21_X1 U11064 ( .B1(n9774), .B2(n10198), .A(n9773), .ZN(n9802) );
  MUX2_X1 U11065 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9802), .S(n10274), .Z(
        P1_U3543) );
  AOI22_X1 U11066 ( .A1(n10194), .A2(n9871), .B1(n9775), .B2(n10191), .ZN(
        n9776) );
  OAI211_X1 U11067 ( .C1(n9778), .C2(n10227), .A(n9777), .B(n9776), .ZN(n9779)
         );
  AOI21_X1 U11068 ( .B1(n9780), .B2(n10203), .A(n9779), .ZN(n9781) );
  OAI21_X1 U11069 ( .B1(n9782), .B2(n10198), .A(n9781), .ZN(n9803) );
  MUX2_X1 U11070 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9803), .S(n10274), .Z(
        P1_U3542) );
  AOI22_X1 U11071 ( .A1(n10194), .A2(n9784), .B1(n9783), .B2(n10191), .ZN(
        n9785) );
  OAI211_X1 U11072 ( .C1(n9787), .C2(n10227), .A(n9786), .B(n9785), .ZN(n9788)
         );
  AOI21_X1 U11073 ( .B1(n9789), .B2(n10203), .A(n9788), .ZN(n9790) );
  OAI21_X1 U11074 ( .B1(n9791), .B2(n10198), .A(n9790), .ZN(n9804) );
  MUX2_X1 U11075 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9804), .S(n10274), .Z(
        P1_U3541) );
  MUX2_X1 U11076 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9792), .S(n10251), .Z(
        P1_U3521) );
  MUX2_X1 U11077 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9793), .S(n10251), .Z(
        P1_U3520) );
  MUX2_X1 U11078 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9794), .S(n10251), .Z(
        P1_U3519) );
  MUX2_X1 U11079 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9795), .S(n10251), .Z(
        P1_U3518) );
  MUX2_X1 U11080 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9796), .S(n10251), .Z(
        P1_U3517) );
  MUX2_X1 U11081 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9797), .S(n10251), .Z(
        P1_U3516) );
  MUX2_X1 U11082 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9798), .S(n10251), .Z(
        P1_U3515) );
  MUX2_X1 U11083 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9799), .S(n10251), .Z(
        P1_U3514) );
  MUX2_X1 U11084 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9800), .S(n10251), .Z(
        P1_U3513) );
  MUX2_X1 U11085 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9801), .S(n10251), .Z(
        P1_U3512) );
  MUX2_X1 U11086 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9802), .S(n10251), .Z(
        P1_U3511) );
  MUX2_X1 U11087 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9803), .S(n10251), .Z(
        P1_U3510) );
  MUX2_X1 U11088 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9804), .S(n10251), .Z(
        P1_U3509) );
  MUX2_X1 U11089 ( .A(n9805), .B(P1_D_REG_1__SCAN_IN), .S(n10113), .Z(P1_U3440) );
  NAND2_X1 U11090 ( .A1(n9807), .A2(n9806), .ZN(n9809) );
  NAND4_X1 U11091 ( .A1(n5145), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .A4(n5146), .ZN(n9808) );
  OAI211_X1 U11092 ( .C1(n9810), .C2(n9817), .A(n9809), .B(n9808), .ZN(
        P1_U3324) );
  OAI222_X1 U11093 ( .A1(P1_U3086), .A2(n9813), .B1(n9820), .B2(n9812), .C1(
        n9811), .C2(n9817), .ZN(P1_U3326) );
  OAI222_X1 U11094 ( .A1(n9924), .A2(P1_U3086), .B1(n9820), .B2(n9816), .C1(
        n9815), .C2(n9814), .ZN(P1_U3328) );
  OAI222_X1 U11095 ( .A1(P1_U3086), .A2(n9821), .B1(n9820), .B2(n9819), .C1(
        n9818), .C2(n9817), .ZN(P1_U3329) );
  MUX2_X1 U11096 ( .A(n9823), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI211_X1 U11097 ( .C1(n9826), .C2(n9825), .A(n9824), .B(n10032), .ZN(n9831)
         );
  AOI211_X1 U11098 ( .C1(n9829), .C2(n9828), .A(n9827), .B(n10036), .ZN(n9830)
         );
  AOI211_X1 U11099 ( .C1(n10043), .C2(n9832), .A(n9831), .B(n9830), .ZN(n9835)
         );
  INV_X1 U11100 ( .A(n9833), .ZN(n9834) );
  OAI211_X1 U11101 ( .C1(n9836), .C2(n10046), .A(n9835), .B(n9834), .ZN(
        P1_U3253) );
  INV_X1 U11102 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9851) );
  NAND2_X1 U11103 ( .A1(n10043), .A2(n9837), .ZN(n9848) );
  AOI21_X1 U11104 ( .B1(n9840), .B2(n9839), .A(n9838), .ZN(n9841) );
  NAND2_X1 U11105 ( .A1(n9983), .A2(n9841), .ZN(n9847) );
  AOI21_X1 U11106 ( .B1(n9844), .B2(n9843), .A(n9842), .ZN(n9845) );
  NAND2_X1 U11107 ( .A1(n9988), .A2(n9845), .ZN(n9846) );
  AND3_X1 U11108 ( .A1(n9848), .A2(n9847), .A3(n9846), .ZN(n9850) );
  OAI211_X1 U11109 ( .C1(n10046), .C2(n9851), .A(n9850), .B(n9849), .ZN(
        P1_U3250) );
  AOI21_X1 U11110 ( .B1(n9854), .B2(n9853), .A(n9852), .ZN(n9855) );
  NAND2_X1 U11111 ( .A1(n9983), .A2(n9855), .ZN(n9863) );
  NAND2_X1 U11112 ( .A1(n10043), .A2(n9856), .ZN(n9862) );
  AOI21_X1 U11113 ( .B1(n9859), .B2(n9858), .A(n9857), .ZN(n9860) );
  NAND2_X1 U11114 ( .A1(n9988), .A2(n9860), .ZN(n9861) );
  AND3_X1 U11115 ( .A1(n9863), .A2(n9862), .A3(n9861), .ZN(n9866) );
  INV_X1 U11116 ( .A(n9864), .ZN(n9865) );
  OAI211_X1 U11117 ( .C1(n9867), .C2(n10046), .A(n9866), .B(n9865), .ZN(
        P1_U3251) );
  NAND2_X1 U11118 ( .A1(n9869), .A2(n9868), .ZN(n9870) );
  XOR2_X1 U11119 ( .A(n9876), .B(n9870), .Z(n9872) );
  AOI222_X1 U11120 ( .A1(n10203), .A2(n9872), .B1(n9871), .B2(n10191), .C1(
        n9898), .C2(n10194), .ZN(n9884) );
  AOI222_X1 U11121 ( .A1(n9874), .A2(n10090), .B1(P1_REG2_REG_18__SCAN_IN), 
        .B2(n4495), .C1(n10092), .C2(n9873), .ZN(n9882) );
  XOR2_X1 U11122 ( .A(n9876), .B(n9875), .Z(n9887) );
  INV_X1 U11123 ( .A(n9877), .ZN(n9878) );
  OAI211_X1 U11124 ( .C1(n9885), .C2(n9879), .A(n9878), .B(n10097), .ZN(n9883)
         );
  INV_X1 U11125 ( .A(n9883), .ZN(n9880) );
  AOI22_X1 U11126 ( .A1(n9887), .A2(n10102), .B1(n10101), .B2(n9880), .ZN(
        n9881) );
  OAI211_X1 U11127 ( .C1(n4495), .C2(n9884), .A(n9882), .B(n9881), .ZN(
        P1_U3275) );
  OAI211_X1 U11128 ( .C1(n9885), .C2(n10227), .A(n9884), .B(n9883), .ZN(n9886)
         );
  AOI21_X1 U11129 ( .B1(n9887), .B2(n10231), .A(n9886), .ZN(n9917) );
  AOI22_X1 U11130 ( .A1(n10274), .A2(n9917), .B1(n9888), .B2(n10272), .ZN(
        P1_U3540) );
  OAI22_X1 U11131 ( .A1(n9889), .A2(n10236), .B1(n9908), .B2(n10234), .ZN(
        n9891) );
  AOI211_X1 U11132 ( .C1(n10241), .C2(n9892), .A(n9891), .B(n9890), .ZN(n9893)
         );
  OAI21_X1 U11133 ( .B1(n10222), .B2(n9894), .A(n9893), .ZN(n9895) );
  AOI21_X1 U11134 ( .B1(n9896), .B2(n10231), .A(n9895), .ZN(n9918) );
  AOI22_X1 U11135 ( .A1(n10274), .A2(n9918), .B1(n5608), .B2(n10272), .ZN(
        P1_U3539) );
  AOI22_X1 U11136 ( .A1(n9898), .A2(n10191), .B1(n9897), .B2(n10194), .ZN(
        n9899) );
  OAI211_X1 U11137 ( .C1(n4802), .C2(n10227), .A(n9900), .B(n9899), .ZN(n9904)
         );
  NOR3_X1 U11138 ( .A1(n9902), .A2(n9901), .A3(n10198), .ZN(n9903) );
  AOI211_X1 U11139 ( .C1(n9905), .C2(n10203), .A(n9904), .B(n9903), .ZN(n9920)
         );
  AOI22_X1 U11140 ( .A1(n10274), .A2(n9920), .B1(n9906), .B2(n10272), .ZN(
        P1_U3538) );
  OAI22_X1 U11141 ( .A1(n9908), .A2(n10236), .B1(n9907), .B2(n10234), .ZN(
        n9910) );
  AOI211_X1 U11142 ( .C1(n10241), .C2(n9911), .A(n9910), .B(n9909), .ZN(n9912)
         );
  OAI21_X1 U11143 ( .B1(n10222), .B2(n9913), .A(n9912), .ZN(n9914) );
  AOI21_X1 U11144 ( .B1(n9915), .B2(n10231), .A(n9914), .ZN(n9922) );
  AOI22_X1 U11145 ( .A1(n10274), .A2(n9922), .B1(n10021), .B2(n10272), .ZN(
        P1_U3537) );
  AOI22_X1 U11146 ( .A1(n10251), .A2(n9917), .B1(n9916), .B2(n10249), .ZN(
        P1_U3507) );
  AOI22_X1 U11147 ( .A1(n10251), .A2(n9918), .B1(n5604), .B2(n10249), .ZN(
        P1_U3504) );
  INV_X1 U11148 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9919) );
  AOI22_X1 U11149 ( .A1(n10251), .A2(n9920), .B1(n9919), .B2(n10249), .ZN(
        P1_U3501) );
  INV_X1 U11150 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9921) );
  AOI22_X1 U11151 ( .A1(n10251), .A2(n9922), .B1(n9921), .B2(n10249), .ZN(
        P1_U3498) );
  XNOR2_X1 U11152 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11153 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U11154 ( .A1(n9924), .A2(n9923), .ZN(n9927) );
  NOR2_X1 U11155 ( .A1(n9925), .A2(n9927), .ZN(n9928) );
  MUX2_X1 U11156 ( .A(n9928), .B(n9927), .S(n9926), .Z(n9930) );
  OR2_X1 U11157 ( .A1(n9930), .A2(n9929), .ZN(n9932) );
  AOI22_X1 U11158 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9945), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9931) );
  OAI21_X1 U11159 ( .B1(n9933), .B2(n9932), .A(n9931), .ZN(P1_U3243) );
  OAI211_X1 U11160 ( .C1(n9936), .C2(n9935), .A(n9983), .B(n9934), .ZN(n9943)
         );
  OAI211_X1 U11161 ( .C1(n9939), .C2(n9938), .A(n9988), .B(n9937), .ZN(n9942)
         );
  NAND2_X1 U11162 ( .A1(n10043), .A2(n9940), .ZN(n9941) );
  AND3_X1 U11163 ( .A1(n9943), .A2(n9942), .A3(n9941), .ZN(n9949) );
  AOI21_X1 U11164 ( .B1(n9945), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n9944), .ZN(
        n9946) );
  AND2_X1 U11165 ( .A1(n9947), .A2(n9946), .ZN(n9948) );
  NAND2_X1 U11166 ( .A1(n9949), .A2(n9948), .ZN(P1_U3247) );
  OAI211_X1 U11167 ( .C1(n9952), .C2(n9951), .A(n9988), .B(n9950), .ZN(n9960)
         );
  NAND2_X1 U11168 ( .A1(n10043), .A2(n9953), .ZN(n9959) );
  AOI21_X1 U11169 ( .B1(n9956), .B2(n9955), .A(n9954), .ZN(n9957) );
  NAND2_X1 U11170 ( .A1(n9983), .A2(n9957), .ZN(n9958) );
  AND3_X1 U11171 ( .A1(n9960), .A2(n9959), .A3(n9958), .ZN(n9962) );
  OAI211_X1 U11172 ( .C1(n10046), .C2(n9963), .A(n9962), .B(n9961), .ZN(
        P1_U3248) );
  INV_X1 U11173 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9977) );
  NAND2_X1 U11174 ( .A1(n10043), .A2(n9964), .ZN(n9974) );
  AOI21_X1 U11175 ( .B1(n9966), .B2(n4547), .A(n9965), .ZN(n9967) );
  NAND2_X1 U11176 ( .A1(n9983), .A2(n9967), .ZN(n9973) );
  AOI21_X1 U11177 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(n9971) );
  NAND2_X1 U11178 ( .A1(n9988), .A2(n9971), .ZN(n9972) );
  AND3_X1 U11179 ( .A1(n9974), .A2(n9973), .A3(n9972), .ZN(n9976) );
  OAI211_X1 U11180 ( .C1(n10046), .C2(n9977), .A(n9976), .B(n9975), .ZN(
        P1_U3249) );
  INV_X1 U11181 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9994) );
  NAND2_X1 U11182 ( .A1(n10043), .A2(n9978), .ZN(n9991) );
  AOI21_X1 U11183 ( .B1(n9981), .B2(n9980), .A(n9979), .ZN(n9982) );
  NAND2_X1 U11184 ( .A1(n9983), .A2(n9982), .ZN(n9990) );
  AOI21_X1 U11185 ( .B1(n9986), .B2(n9985), .A(n9984), .ZN(n9987) );
  NAND2_X1 U11186 ( .A1(n9988), .A2(n9987), .ZN(n9989) );
  AND3_X1 U11187 ( .A1(n9991), .A2(n9990), .A3(n9989), .ZN(n9993) );
  NAND2_X1 U11188 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9992) );
  OAI211_X1 U11189 ( .C1(n10046), .C2(n9994), .A(n9993), .B(n9992), .ZN(
        P1_U3254) );
  INV_X1 U11190 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10006) );
  AOI211_X1 U11191 ( .C1(n9997), .C2(n9996), .A(n10032), .B(n9995), .ZN(n10002) );
  AOI211_X1 U11192 ( .C1(n10000), .C2(n9999), .A(n10036), .B(n9998), .ZN(
        n10001) );
  AOI211_X1 U11193 ( .C1(n10043), .C2(n10003), .A(n10002), .B(n10001), .ZN(
        n10005) );
  NAND2_X1 U11194 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n10004)
         );
  OAI211_X1 U11195 ( .C1(n10046), .C2(n10006), .A(n10005), .B(n10004), .ZN(
        P1_U3256) );
  AOI211_X1 U11196 ( .C1(n10009), .C2(n10008), .A(n10007), .B(n10036), .ZN(
        n10014) );
  AOI211_X1 U11197 ( .C1(n10012), .C2(n10011), .A(n10032), .B(n10010), .ZN(
        n10013) );
  AOI211_X1 U11198 ( .C1(n10043), .C2(n10015), .A(n10014), .B(n10013), .ZN(
        n10018) );
  INV_X1 U11199 ( .A(n10016), .ZN(n10017) );
  OAI211_X1 U11200 ( .C1(n10019), .C2(n10046), .A(n10018), .B(n10017), .ZN(
        P1_U3257) );
  INV_X1 U11201 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10031) );
  AOI211_X1 U11202 ( .C1(n10022), .C2(n10021), .A(n10020), .B(n10032), .ZN(
        n10027) );
  AOI211_X1 U11203 ( .C1(n10025), .C2(n10024), .A(n10023), .B(n10036), .ZN(
        n10026) );
  AOI211_X1 U11204 ( .C1(n10043), .C2(n10028), .A(n10027), .B(n10026), .ZN(
        n10030) );
  NAND2_X1 U11205 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n10029)
         );
  OAI211_X1 U11206 ( .C1(n10046), .C2(n10031), .A(n10030), .B(n10029), .ZN(
        P1_U3258) );
  AOI211_X1 U11207 ( .C1(n10035), .C2(n10034), .A(n10033), .B(n10032), .ZN(
        n10041) );
  AOI211_X1 U11208 ( .C1(n10039), .C2(n10038), .A(n10037), .B(n10036), .ZN(
        n10040) );
  AOI211_X1 U11209 ( .C1(n10043), .C2(n10042), .A(n10041), .B(n10040), .ZN(
        n10045) );
  NAND2_X1 U11210 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n10044)
         );
  OAI211_X1 U11211 ( .C1(n10047), .C2(n10046), .A(n10045), .B(n10044), .ZN(
        P1_U3261) );
  OAI211_X1 U11212 ( .C1(n10049), .C2(n10054), .A(n10048), .B(n10203), .ZN(
        n10051) );
  AOI22_X1 U11213 ( .A1(n10194), .A2(n10065), .B1(n10193), .B2(n10191), .ZN(
        n10050) );
  AND2_X1 U11214 ( .A1(n10051), .A2(n10050), .ZN(n10178) );
  AOI222_X1 U11215 ( .A1(n10053), .A2(n10090), .B1(P1_REG2_REG_8__SCAN_IN), 
        .B2(n4495), .C1(n10092), .C2(n10052), .ZN(n10062) );
  XNOR2_X1 U11216 ( .A(n10055), .B(n10054), .ZN(n10181) );
  INV_X1 U11217 ( .A(n10056), .ZN(n10059) );
  INV_X1 U11218 ( .A(n10057), .ZN(n10058) );
  OAI211_X1 U11219 ( .C1(n10179), .C2(n10059), .A(n10058), .B(n10097), .ZN(
        n10177) );
  INV_X1 U11220 ( .A(n10177), .ZN(n10060) );
  AOI22_X1 U11221 ( .A1(n10181), .A2(n10102), .B1(n10101), .B2(n10060), .ZN(
        n10061) );
  OAI211_X1 U11222 ( .C1(n4495), .C2(n10178), .A(n10062), .B(n10061), .ZN(
        P1_U3285) );
  XNOR2_X1 U11223 ( .A(n10063), .B(n10068), .ZN(n10064) );
  AOI222_X1 U11224 ( .A1(n6632), .A2(n10194), .B1(n10065), .B2(n10191), .C1(
        n10203), .C2(n10064), .ZN(n10161) );
  AOI222_X1 U11225 ( .A1(n10067), .A2(n10090), .B1(P1_REG2_REG_6__SCAN_IN), 
        .B2(n4495), .C1(n10066), .C2(n10092), .ZN(n10074) );
  XNOR2_X1 U11226 ( .A(n10069), .B(n10068), .ZN(n10164) );
  OAI211_X1 U11227 ( .C1(n10071), .C2(n10160), .A(n10070), .B(n10097), .ZN(
        n10159) );
  INV_X1 U11228 ( .A(n10159), .ZN(n10072) );
  AOI22_X1 U11229 ( .A1(n10164), .A2(n10102), .B1(n10101), .B2(n10072), .ZN(
        n10073) );
  OAI211_X1 U11230 ( .C1(n4495), .C2(n10161), .A(n10074), .B(n10073), .ZN(
        P1_U3287) );
  XNOR2_X1 U11231 ( .A(n10075), .B(n10079), .ZN(n10076) );
  AOI222_X1 U11232 ( .A1(n10089), .A2(n10194), .B1(n6632), .B2(n10191), .C1(
        n10203), .C2(n10076), .ZN(n10144) );
  AOI222_X1 U11233 ( .A1(n10078), .A2(n10090), .B1(P1_REG2_REG_4__SCAN_IN), 
        .B2(n4495), .C1(n10092), .C2(n10077), .ZN(n10086) );
  XNOR2_X1 U11234 ( .A(n10080), .B(n10079), .ZN(n10147) );
  INV_X1 U11235 ( .A(n10081), .ZN(n10083) );
  OAI211_X1 U11236 ( .C1(n10083), .C2(n10143), .A(n10097), .B(n10082), .ZN(
        n10142) );
  INV_X1 U11237 ( .A(n10142), .ZN(n10084) );
  AOI22_X1 U11238 ( .A1(n10147), .A2(n10102), .B1(n10101), .B2(n10084), .ZN(
        n10085) );
  OAI211_X1 U11239 ( .C1(n4495), .C2(n10144), .A(n10086), .B(n10085), .ZN(
        P1_U3289) );
  XNOR2_X1 U11240 ( .A(n10087), .B(n10094), .ZN(n10088) );
  AOI222_X1 U11241 ( .A1(n6717), .A2(n10194), .B1(n10089), .B2(n10191), .C1(
        n10203), .C2(n10088), .ZN(n10129) );
  AOI222_X1 U11242 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n4495), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10092), .C1(n10091), .C2(n10090), .ZN(
        n10104) );
  XNOR2_X1 U11243 ( .A(n10093), .B(n10094), .ZN(n10132) );
  INV_X1 U11244 ( .A(n10096), .ZN(n10098) );
  OAI211_X1 U11245 ( .C1(n10095), .C2(n10099), .A(n10098), .B(n10097), .ZN(
        n10128) );
  INV_X1 U11246 ( .A(n10128), .ZN(n10100) );
  AOI22_X1 U11247 ( .A1(n10132), .A2(n10102), .B1(n10101), .B2(n10100), .ZN(
        n10103) );
  OAI211_X1 U11248 ( .C1(n4495), .C2(n10129), .A(n10104), .B(n10103), .ZN(
        P1_U3291) );
  AND2_X1 U11249 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10113), .ZN(P1_U3294) );
  NOR2_X1 U11250 ( .A1(n10115), .A2(n10105), .ZN(P1_U3295) );
  AND2_X1 U11251 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10113), .ZN(P1_U3296) );
  AND2_X1 U11252 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10113), .ZN(P1_U3297) );
  AND2_X1 U11253 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10113), .ZN(P1_U3298) );
  AND2_X1 U11254 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10113), .ZN(P1_U3299) );
  AND2_X1 U11255 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10113), .ZN(P1_U3300) );
  AND2_X1 U11256 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10113), .ZN(P1_U3301) );
  NOR2_X1 U11257 ( .A1(n10115), .A2(n10106), .ZN(P1_U3302) );
  AND2_X1 U11258 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10113), .ZN(P1_U3303) );
  AND2_X1 U11259 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10113), .ZN(P1_U3304) );
  NOR2_X1 U11260 ( .A1(n10115), .A2(n10107), .ZN(P1_U3305) );
  AND2_X1 U11261 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10113), .ZN(P1_U3306) );
  NOR2_X1 U11262 ( .A1(n10115), .A2(n10108), .ZN(P1_U3307) );
  NOR2_X1 U11263 ( .A1(n10115), .A2(n10109), .ZN(P1_U3308) );
  AND2_X1 U11264 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10113), .ZN(P1_U3309) );
  AND2_X1 U11265 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10113), .ZN(P1_U3310) );
  AND2_X1 U11266 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10113), .ZN(P1_U3311) );
  AND2_X1 U11267 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10113), .ZN(P1_U3312) );
  AND2_X1 U11268 ( .A1(n10113), .A2(P1_D_REG_12__SCAN_IN), .ZN(P1_U3313) );
  AND2_X1 U11269 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10113), .ZN(P1_U3314) );
  NOR2_X1 U11270 ( .A1(n10115), .A2(n10110), .ZN(P1_U3315) );
  AND2_X1 U11271 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10113), .ZN(P1_U3316) );
  AND2_X1 U11272 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10113), .ZN(P1_U3317) );
  NOR2_X1 U11273 ( .A1(n10115), .A2(n10111), .ZN(P1_U3318) );
  AND2_X1 U11274 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10113), .ZN(P1_U3319) );
  NOR2_X1 U11275 ( .A1(n10115), .A2(n10112), .ZN(P1_U3320) );
  AND2_X1 U11276 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10113), .ZN(P1_U3321) );
  AND2_X1 U11277 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10113), .ZN(P1_U3322) );
  NOR2_X1 U11278 ( .A1(n10115), .A2(n10114), .ZN(P1_U3323) );
  INV_X1 U11279 ( .A(n10116), .ZN(n10248) );
  INV_X1 U11280 ( .A(n10124), .ZN(n10126) );
  OAI22_X1 U11281 ( .A1(n10118), .A2(n10236), .B1(n10117), .B2(n10227), .ZN(
        n10120) );
  AOI211_X1 U11282 ( .C1(n10194), .C2(n10121), .A(n10120), .B(n10119), .ZN(
        n10123) );
  OAI211_X1 U11283 ( .C1(n10124), .C2(n10244), .A(n10123), .B(n10122), .ZN(
        n10125) );
  AOI21_X1 U11284 ( .B1(n10248), .B2(n10126), .A(n10125), .ZN(n10253) );
  INV_X1 U11285 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10127) );
  AOI22_X1 U11286 ( .A1(n10251), .A2(n10253), .B1(n10127), .B2(n10249), .ZN(
        P1_U3456) );
  OAI21_X1 U11287 ( .B1(n10095), .B2(n10227), .A(n10128), .ZN(n10131) );
  INV_X1 U11288 ( .A(n10129), .ZN(n10130) );
  AOI211_X1 U11289 ( .C1(n10231), .C2(n10132), .A(n10131), .B(n10130), .ZN(
        n10255) );
  INV_X1 U11290 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10133) );
  AOI22_X1 U11291 ( .A1(n10251), .A2(n10255), .B1(n10133), .B2(n10249), .ZN(
        P1_U3459) );
  INV_X1 U11292 ( .A(n10134), .ZN(n10140) );
  INV_X1 U11293 ( .A(n10135), .ZN(n10136) );
  OAI211_X1 U11294 ( .C1(n10138), .C2(n10227), .A(n10137), .B(n10136), .ZN(
        n10139) );
  AOI21_X1 U11295 ( .B1(n10231), .B2(n10140), .A(n10139), .ZN(n10257) );
  INV_X1 U11296 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10141) );
  AOI22_X1 U11297 ( .A1(n10251), .A2(n10257), .B1(n10141), .B2(n10249), .ZN(
        P1_U3462) );
  OAI21_X1 U11298 ( .B1(n10143), .B2(n10227), .A(n10142), .ZN(n10146) );
  INV_X1 U11299 ( .A(n10144), .ZN(n10145) );
  AOI211_X1 U11300 ( .C1(n10231), .C2(n10147), .A(n10146), .B(n10145), .ZN(
        n10259) );
  INV_X1 U11301 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10148) );
  AOI22_X1 U11302 ( .A1(n10251), .A2(n10259), .B1(n10148), .B2(n10249), .ZN(
        P1_U3465) );
  OAI22_X1 U11303 ( .A1(n10150), .A2(n10234), .B1(n10149), .B2(n10236), .ZN(
        n10152) );
  AOI211_X1 U11304 ( .C1(n10241), .C2(n10153), .A(n10152), .B(n10151), .ZN(
        n10154) );
  OAI21_X1 U11305 ( .B1(n10155), .B2(n10198), .A(n10154), .ZN(n10156) );
  AOI21_X1 U11306 ( .B1(n10157), .B2(n10203), .A(n10156), .ZN(n10261) );
  INV_X1 U11307 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10158) );
  AOI22_X1 U11308 ( .A1(n10251), .A2(n10261), .B1(n10158), .B2(n10249), .ZN(
        P1_U3468) );
  OAI21_X1 U11309 ( .B1(n10160), .B2(n10227), .A(n10159), .ZN(n10163) );
  INV_X1 U11310 ( .A(n10161), .ZN(n10162) );
  AOI211_X1 U11311 ( .C1(n10231), .C2(n10164), .A(n10163), .B(n10162), .ZN(
        n10262) );
  INV_X1 U11312 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10165) );
  AOI22_X1 U11313 ( .A1(n10251), .A2(n10262), .B1(n10165), .B2(n10249), .ZN(
        P1_U3471) );
  INV_X1 U11314 ( .A(n10173), .ZN(n10175) );
  AOI22_X1 U11315 ( .A1(n10194), .A2(n10166), .B1(n10184), .B2(n10191), .ZN(
        n10167) );
  OAI211_X1 U11316 ( .C1(n10169), .C2(n10227), .A(n10168), .B(n10167), .ZN(
        n10170) );
  NOR2_X1 U11317 ( .A1(n10171), .A2(n10170), .ZN(n10172) );
  OAI21_X1 U11318 ( .B1(n10173), .B2(n10244), .A(n10172), .ZN(n10174) );
  AOI21_X1 U11319 ( .B1(n10248), .B2(n10175), .A(n10174), .ZN(n10263) );
  INV_X1 U11320 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U11321 ( .A1(n10251), .A2(n10263), .B1(n10176), .B2(n10249), .ZN(
        P1_U3474) );
  OAI211_X1 U11322 ( .C1(n10179), .C2(n10227), .A(n10178), .B(n10177), .ZN(
        n10180) );
  AOI21_X1 U11323 ( .B1(n10231), .B2(n10181), .A(n10180), .ZN(n10264) );
  INV_X1 U11324 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10182) );
  AOI22_X1 U11325 ( .A1(n10251), .A2(n10264), .B1(n10182), .B2(n10249), .ZN(
        P1_U3477) );
  AOI22_X1 U11326 ( .A1(n10184), .A2(n10194), .B1(n10241), .B2(n10183), .ZN(
        n10185) );
  OAI211_X1 U11327 ( .C1(n10187), .C2(n10198), .A(n10186), .B(n10185), .ZN(
        n10188) );
  AOI21_X1 U11328 ( .B1(n10203), .B2(n10189), .A(n10188), .ZN(n10266) );
  INV_X1 U11329 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U11330 ( .A1(n10251), .A2(n10266), .B1(n10190), .B2(n10249), .ZN(
        P1_U3480) );
  AOI22_X1 U11331 ( .A1(n10194), .A2(n10193), .B1(n10192), .B2(n10191), .ZN(
        n10195) );
  OAI211_X1 U11332 ( .C1(n10197), .C2(n10227), .A(n10196), .B(n10195), .ZN(
        n10201) );
  NOR2_X1 U11333 ( .A1(n10199), .A2(n10198), .ZN(n10200) );
  AOI211_X1 U11334 ( .C1(n10203), .C2(n10202), .A(n10201), .B(n10200), .ZN(
        n10267) );
  AOI22_X1 U11335 ( .A1(n10251), .A2(n10267), .B1(n10204), .B2(n10249), .ZN(
        P1_U3483) );
  INV_X1 U11336 ( .A(n10212), .ZN(n10214) );
  OAI22_X1 U11337 ( .A1(n10206), .A2(n10236), .B1(n10205), .B2(n10234), .ZN(
        n10208) );
  AOI211_X1 U11338 ( .C1(n10241), .C2(n10209), .A(n10208), .B(n10207), .ZN(
        n10211) );
  OAI211_X1 U11339 ( .C1(n10212), .C2(n10244), .A(n10211), .B(n10210), .ZN(
        n10213) );
  AOI21_X1 U11340 ( .B1(n10248), .B2(n10214), .A(n10213), .ZN(n10268) );
  INV_X1 U11341 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10215) );
  AOI22_X1 U11342 ( .A1(n10251), .A2(n10268), .B1(n10215), .B2(n10249), .ZN(
        P1_U3486) );
  OAI22_X1 U11343 ( .A1(n10235), .A2(n10236), .B1(n10216), .B2(n10234), .ZN(
        n10218) );
  AOI211_X1 U11344 ( .C1(n10241), .C2(n10219), .A(n10218), .B(n10217), .ZN(
        n10220) );
  OAI21_X1 U11345 ( .B1(n10222), .B2(n10221), .A(n10220), .ZN(n10223) );
  AOI21_X1 U11346 ( .B1(n10224), .B2(n10231), .A(n10223), .ZN(n10270) );
  INV_X1 U11347 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10225) );
  AOI22_X1 U11348 ( .A1(n10251), .A2(n10270), .B1(n10225), .B2(n10249), .ZN(
        P1_U3489) );
  OAI21_X1 U11349 ( .B1(n10228), .B2(n10227), .A(n10226), .ZN(n10229) );
  AOI211_X1 U11350 ( .C1(n10232), .C2(n10231), .A(n10230), .B(n10229), .ZN(
        n10271) );
  AOI22_X1 U11351 ( .A1(n10251), .A2(n10271), .B1(n10233), .B2(n10249), .ZN(
        P1_U3492) );
  INV_X1 U11352 ( .A(n10245), .ZN(n10247) );
  OAI22_X1 U11353 ( .A1(n10237), .A2(n10236), .B1(n10235), .B2(n10234), .ZN(
        n10239) );
  AOI211_X1 U11354 ( .C1(n10241), .C2(n10240), .A(n10239), .B(n10238), .ZN(
        n10243) );
  OAI211_X1 U11355 ( .C1(n10245), .C2(n10244), .A(n10243), .B(n10242), .ZN(
        n10246) );
  AOI21_X1 U11356 ( .B1(n10248), .B2(n10247), .A(n10246), .ZN(n10273) );
  AOI22_X1 U11357 ( .A1(n10251), .A2(n10273), .B1(n10250), .B2(n10249), .ZN(
        P1_U3495) );
  AOI22_X1 U11358 ( .A1(n10274), .A2(n10253), .B1(n10252), .B2(n10272), .ZN(
        P1_U3523) );
  AOI22_X1 U11359 ( .A1(n10274), .A2(n10255), .B1(n10254), .B2(n10272), .ZN(
        P1_U3524) );
  AOI22_X1 U11360 ( .A1(n10274), .A2(n10257), .B1(n10256), .B2(n10272), .ZN(
        P1_U3525) );
  AOI22_X1 U11361 ( .A1(n10274), .A2(n10259), .B1(n10258), .B2(n10272), .ZN(
        P1_U3526) );
  AOI22_X1 U11362 ( .A1(n10274), .A2(n10261), .B1(n10260), .B2(n10272), .ZN(
        P1_U3527) );
  AOI22_X1 U11363 ( .A1(n10274), .A2(n10262), .B1(n6109), .B2(n10272), .ZN(
        P1_U3528) );
  AOI22_X1 U11364 ( .A1(n10274), .A2(n10263), .B1(n6110), .B2(n10272), .ZN(
        P1_U3529) );
  AOI22_X1 U11365 ( .A1(n10274), .A2(n10264), .B1(n6111), .B2(n10272), .ZN(
        P1_U3530) );
  AOI22_X1 U11366 ( .A1(n10274), .A2(n10266), .B1(n10265), .B2(n10272), .ZN(
        P1_U3531) );
  AOI22_X1 U11367 ( .A1(n10274), .A2(n10267), .B1(n6363), .B2(n10272), .ZN(
        P1_U3532) );
  AOI22_X1 U11368 ( .A1(n10274), .A2(n10268), .B1(n6366), .B2(n10272), .ZN(
        P1_U3533) );
  AOI22_X1 U11369 ( .A1(n10274), .A2(n10270), .B1(n10269), .B2(n10272), .ZN(
        P1_U3534) );
  AOI22_X1 U11370 ( .A1(n10274), .A2(n10271), .B1(n7112), .B2(n10272), .ZN(
        P1_U3535) );
  AOI22_X1 U11371 ( .A1(n10274), .A2(n10273), .B1(n7113), .B2(n10272), .ZN(
        P1_U3536) );
  AOI22_X1 U11372 ( .A1(n10275), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n10282) );
  NOR2_X1 U11373 ( .A1(n10276), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10277) );
  OAI22_X1 U11374 ( .A1(n10280), .A2(n10279), .B1(n10278), .B2(n10277), .ZN(
        n10281) );
  OAI211_X1 U11375 ( .C1(n10283), .C2(n4966), .A(n10282), .B(n10281), .ZN(
        P2_U3182) );
  XOR2_X1 U11376 ( .A(n10290), .B(n10284), .Z(n10288) );
  AOI222_X1 U11377 ( .A1(n10289), .A2(n10288), .B1(n10287), .B2(n10286), .C1(
        n4512), .C2(n10285), .ZN(n10314) );
  XNOR2_X1 U11378 ( .A(n10291), .B(n10290), .ZN(n10317) );
  AOI222_X1 U11379 ( .A1(n10317), .A2(n10296), .B1(n10295), .B2(n10294), .C1(
        n10293), .C2(n10292), .ZN(n10297) );
  OAI221_X1 U11380 ( .B1(n8381), .B2(n10314), .C1(n10299), .C2(n10298), .A(
        n10297), .ZN(P2_U3230) );
  INV_X1 U11381 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10305) );
  AOI21_X1 U11382 ( .B1(n10301), .B2(n10361), .A(n10300), .ZN(n10302) );
  AOI211_X1 U11383 ( .C1(n10366), .C2(n10304), .A(n10303), .B(n10302), .ZN(
        n10370) );
  AOI22_X1 U11384 ( .A1(n10369), .A2(n10305), .B1(n10370), .B2(n10367), .ZN(
        P2_U3390) );
  INV_X1 U11385 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10307) );
  AOI22_X1 U11386 ( .A1(n10369), .A2(n10307), .B1(n10306), .B2(n10367), .ZN(
        P2_U3393) );
  INV_X1 U11387 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10313) );
  AOI21_X1 U11388 ( .B1(n10351), .B2(n10309), .A(n10308), .ZN(n10311) );
  AOI211_X1 U11389 ( .C1(n10366), .C2(n10312), .A(n10311), .B(n10310), .ZN(
        n10372) );
  AOI22_X1 U11390 ( .A1(n10369), .A2(n10313), .B1(n10372), .B2(n10367), .ZN(
        P2_U3396) );
  INV_X1 U11391 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10318) );
  OAI21_X1 U11392 ( .B1(n10315), .B2(n10356), .A(n10314), .ZN(n10316) );
  AOI21_X1 U11393 ( .B1(n10345), .B2(n10317), .A(n10316), .ZN(n10374) );
  AOI22_X1 U11394 ( .A1(n10369), .A2(n10318), .B1(n10374), .B2(n10367), .ZN(
        P2_U3399) );
  INV_X1 U11395 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10324) );
  INV_X1 U11396 ( .A(n10319), .ZN(n10323) );
  OAI21_X1 U11397 ( .B1(n10321), .B2(n10356), .A(n10320), .ZN(n10322) );
  AOI21_X1 U11398 ( .B1(n10323), .B2(n10345), .A(n10322), .ZN(n10375) );
  AOI22_X1 U11399 ( .A1(n10369), .A2(n10324), .B1(n10375), .B2(n10367), .ZN(
        P2_U3402) );
  INV_X1 U11400 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10329) );
  NOR2_X1 U11401 ( .A1(n10325), .A2(n10356), .ZN(n10327) );
  AOI211_X1 U11402 ( .C1(n10345), .C2(n10328), .A(n10327), .B(n10326), .ZN(
        n10376) );
  AOI22_X1 U11403 ( .A1(n10369), .A2(n10329), .B1(n10376), .B2(n10367), .ZN(
        P2_U3405) );
  NOR2_X1 U11404 ( .A1(n10330), .A2(n10356), .ZN(n10332) );
  AOI211_X1 U11405 ( .C1(n10333), .C2(n10345), .A(n10332), .B(n10331), .ZN(
        n10378) );
  AOI22_X1 U11406 ( .A1(n10369), .A2(n6763), .B1(n10378), .B2(n10367), .ZN(
        P2_U3408) );
  INV_X1 U11407 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10338) );
  OAI22_X1 U11408 ( .A1(n10335), .A2(n10351), .B1(n10334), .B2(n10356), .ZN(
        n10336) );
  NOR2_X1 U11409 ( .A1(n10337), .A2(n10336), .ZN(n10379) );
  AOI22_X1 U11410 ( .A1(n10369), .A2(n10338), .B1(n10379), .B2(n10367), .ZN(
        P2_U3411) );
  INV_X1 U11411 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10343) );
  NOR2_X1 U11412 ( .A1(n10339), .A2(n10356), .ZN(n10341) );
  AOI211_X1 U11413 ( .C1(n10345), .C2(n10342), .A(n10341), .B(n10340), .ZN(
        n10380) );
  AOI22_X1 U11414 ( .A1(n10369), .A2(n10343), .B1(n10380), .B2(n10367), .ZN(
        P2_U3414) );
  INV_X1 U11415 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10349) );
  AND3_X1 U11416 ( .A1(n7145), .A2(n10345), .A3(n10344), .ZN(n10347) );
  AOI211_X1 U11417 ( .C1(n10366), .C2(n10348), .A(n10347), .B(n10346), .ZN(
        n10381) );
  AOI22_X1 U11418 ( .A1(n10369), .A2(n10349), .B1(n10381), .B2(n10367), .ZN(
        P2_U3417) );
  INV_X1 U11419 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10355) );
  OAI22_X1 U11420 ( .A1(n10352), .A2(n10351), .B1(n10350), .B2(n10356), .ZN(
        n10353) );
  NOR2_X1 U11421 ( .A1(n10354), .A2(n10353), .ZN(n10382) );
  AOI22_X1 U11422 ( .A1(n10369), .A2(n10355), .B1(n10382), .B2(n10367), .ZN(
        P2_U3420) );
  OAI22_X1 U11423 ( .A1(n10358), .A2(n10361), .B1(n10357), .B2(n10356), .ZN(
        n10359) );
  NOR2_X1 U11424 ( .A1(n10360), .A2(n10359), .ZN(n10383) );
  AOI22_X1 U11425 ( .A1(n10369), .A2(n7156), .B1(n10383), .B2(n10367), .ZN(
        P2_U3423) );
  INV_X1 U11426 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10368) );
  NOR2_X1 U11427 ( .A1(n10362), .A2(n10361), .ZN(n10364) );
  AOI211_X1 U11428 ( .C1(n10366), .C2(n10365), .A(n10364), .B(n10363), .ZN(
        n10385) );
  AOI22_X1 U11429 ( .A1(n10369), .A2(n10368), .B1(n10385), .B2(n10367), .ZN(
        P2_U3426) );
  AOI22_X1 U11430 ( .A1(n10386), .A2(n10370), .B1(n4931), .B2(n10384), .ZN(
        P2_U3459) );
  AOI22_X1 U11431 ( .A1(n10386), .A2(n10372), .B1(n10371), .B2(n10384), .ZN(
        P2_U3461) );
  INV_X1 U11432 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10373) );
  AOI22_X1 U11433 ( .A1(n10386), .A2(n10374), .B1(n10373), .B2(n10384), .ZN(
        P2_U3462) );
  AOI22_X1 U11434 ( .A1(n10386), .A2(n10375), .B1(n6510), .B2(n10384), .ZN(
        P2_U3463) );
  AOI22_X1 U11435 ( .A1(n10386), .A2(n10376), .B1(n6652), .B2(n10384), .ZN(
        P2_U3464) );
  AOI22_X1 U11436 ( .A1(n10386), .A2(n10378), .B1(n10377), .B2(n10384), .ZN(
        P2_U3465) );
  AOI22_X1 U11437 ( .A1(n10386), .A2(n10379), .B1(n6878), .B2(n10384), .ZN(
        P2_U3466) );
  AOI22_X1 U11438 ( .A1(n10386), .A2(n10380), .B1(n6930), .B2(n10384), .ZN(
        P2_U3467) );
  AOI22_X1 U11439 ( .A1(n10386), .A2(n10381), .B1(n7041), .B2(n10384), .ZN(
        P2_U3468) );
  AOI22_X1 U11440 ( .A1(n10386), .A2(n10382), .B1(n7073), .B2(n10384), .ZN(
        P2_U3469) );
  AOI22_X1 U11441 ( .A1(n10386), .A2(n10383), .B1(n7155), .B2(n10384), .ZN(
        P2_U3470) );
  AOI22_X1 U11442 ( .A1(n10386), .A2(n10385), .B1(n7273), .B2(n10384), .ZN(
        P2_U3471) );
  OAI222_X1 U11443 ( .A1(n10391), .A2(n10390), .B1(n10391), .B2(n10389), .C1(
        n10388), .C2(n10387), .ZN(ADD_1068_U5) );
  AOI21_X1 U11444 ( .B1(n10394), .B2(n10393), .A(n10392), .ZN(ADD_1068_U46) );
  INV_X1 U11445 ( .A(n10397), .ZN(n10396) );
  OAI222_X1 U11446 ( .A1(n10399), .A2(n10398), .B1(n10399), .B2(n10397), .C1(
        n10396), .C2(n10395), .ZN(ADD_1068_U55) );
  OAI21_X1 U11447 ( .B1(n10402), .B2(n10401), .A(n10400), .ZN(ADD_1068_U56) );
  OAI21_X1 U11448 ( .B1(n10405), .B2(n10404), .A(n10403), .ZN(ADD_1068_U57) );
  OAI21_X1 U11449 ( .B1(n10408), .B2(n10407), .A(n10406), .ZN(ADD_1068_U58) );
  OAI21_X1 U11450 ( .B1(n10411), .B2(n10410), .A(n10409), .ZN(ADD_1068_U59) );
  OAI21_X1 U11451 ( .B1(n10414), .B2(n10413), .A(n10412), .ZN(ADD_1068_U60) );
  OAI21_X1 U11452 ( .B1(n10417), .B2(n10416), .A(n10415), .ZN(ADD_1068_U61) );
  OAI21_X1 U11453 ( .B1(n10420), .B2(n10419), .A(n10418), .ZN(ADD_1068_U62) );
  OAI21_X1 U11454 ( .B1(n10423), .B2(n10422), .A(n10421), .ZN(ADD_1068_U63) );
  OAI21_X1 U11455 ( .B1(n10426), .B2(n10425), .A(n10424), .ZN(ADD_1068_U50) );
  OAI21_X1 U11456 ( .B1(n10429), .B2(n10428), .A(n10427), .ZN(ADD_1068_U48) );
  OAI21_X1 U11457 ( .B1(n10432), .B2(n10431), .A(n10430), .ZN(ADD_1068_U51) );
  OAI21_X1 U11458 ( .B1(n10435), .B2(n10434), .A(n10433), .ZN(ADD_1068_U49) );
  OAI21_X1 U11459 ( .B1(n10438), .B2(n10437), .A(n10436), .ZN(ADD_1068_U47) );
  AOI21_X1 U11460 ( .B1(n10441), .B2(n10440), .A(n10439), .ZN(ADD_1068_U54) );
  AOI21_X1 U11461 ( .B1(n10444), .B2(n10443), .A(n10442), .ZN(ADD_1068_U53) );
  OAI21_X1 U11462 ( .B1(n10447), .B2(n10446), .A(n10445), .ZN(ADD_1068_U52) );
  NAND3_X1 U5147 ( .A1(n5081), .A2(n5080), .A3(n5129), .ZN(n5372) );
endmodule

