

module b15_C_AntiSAT_k_128_6 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753;

  INV_X1 U3443 ( .A(n3404), .ZN(n5241) );
  BUF_X1 U3444 ( .A(n3530), .Z(n3612) );
  INV_X1 U34450 ( .A(n3801), .ZN(n4448) );
  CLKBUF_X2 U34460 ( .A(n5196), .Z(n5024) );
  CLKBUF_X2 U34470 ( .A(n3189), .Z(n5195) );
  CLKBUF_X2 U34480 ( .A(n3204), .Z(n2999) );
  CLKBUF_X2 U3449 ( .A(n3203), .Z(n5197) );
  CLKBUF_X2 U3450 ( .A(n3182), .Z(n5198) );
  CLKBUF_X2 U34510 ( .A(n3180), .Z(n5189) );
  CLKBUF_X2 U34520 ( .A(n3205), .Z(n3001) );
  INV_X1 U34530 ( .A(n3973), .ZN(n3636) );
  CLKBUF_X2 U3454 ( .A(n3166), .Z(n5187) );
  AND4_X1 U34550 ( .A1(n3093), .A2(n3092), .A3(n3091), .A4(n3090), .ZN(n3099)
         );
  AND2_X2 U34560 ( .A1(n3898), .A2(n3023), .ZN(n3179) );
  INV_X2 U3457 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3997) );
  NOR2_X1 U3458 ( .A1(n3129), .A2(n3629), .ZN(n3432) );
  AND2_X1 U34590 ( .A1(n5604), .A2(n5601), .ZN(n5592) );
  NOR2_X1 U34600 ( .A1(n5276), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4792) );
  NAND2_X1 U34610 ( .A1(n3674), .A2(n3452), .ZN(n5934) );
  AOI211_X1 U34630 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5331), .A(n5294), .B(
        n5293), .ZN(n5295) );
  INV_X1 U34640 ( .A(n6032), .ZN(n6058) );
  INV_X1 U34650 ( .A(n6079), .ZN(n6101) );
  NAND2_X2 U3466 ( .A1(n5108), .A2(n3921), .ZN(n3765) );
  NOR2_X4 U3467 ( .A1(n4382), .A2(n4381), .ZN(n4509) );
  OR2_X2 U34680 ( .A1(n3302), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6211)
         );
  XNOR2_X2 U34690 ( .A(n3529), .B(n3940), .ZN(n3799) );
  NAND2_X2 U34700 ( .A1(n3525), .A2(n3524), .ZN(n3529) );
  NOR2_X4 U34710 ( .A1(n4506), .A2(n4507), .ZN(n4666) );
  INV_X4 U34720 ( .A(n3950), .ZN(n3624) );
  NAND2_X2 U34730 ( .A1(n3294), .A2(n3293), .ZN(n3309) );
  AND2_X2 U34740 ( .A1(n3242), .A2(n3241), .ZN(n3293) );
  AND2_X2 U3477 ( .A1(n3144), .A2(n3143), .ZN(n3674) );
  INV_X4 U3478 ( .A(n5241), .ZN(n2996) );
  NAND2_X1 U3479 ( .A1(n6111), .A2(n5107), .ZN(n5466) );
  NAND2_X1 U3480 ( .A1(n3236), .A2(n3235), .ZN(n3280) );
  CLKBUF_X2 U3481 ( .A(n3112), .Z(n3979) );
  INV_X1 U3482 ( .A(n3116), .ZN(n3921) );
  CLKBUF_X2 U3483 ( .A(n3179), .Z(n5167) );
  BUF_X2 U3484 ( .A(n3187), .Z(n5185) );
  BUF_X2 U3485 ( .A(n3196), .Z(n2998) );
  CLKBUF_X1 U3486 ( .A(n3425), .Z(n5545) );
  CLKBUF_X1 U3487 ( .A(n5594), .Z(n5612) );
  NOR2_X1 U3488 ( .A1(n4376), .A2(n4375), .ZN(n4377) );
  NAND2_X1 U3489 ( .A1(n3358), .A2(n3357), .ZN(n4157) );
  NAND2_X1 U3490 ( .A1(n3354), .A2(n3353), .ZN(n3356) );
  NAND2_X1 U3491 ( .A1(n3394), .A2(n3393), .ZN(n3404) );
  OR2_X1 U3492 ( .A1(n4050), .A2(n3488), .ZN(n3354) );
  OR2_X1 U3493 ( .A1(n3370), .A2(n3369), .ZN(n3394) );
  NAND2_X2 U3494 ( .A1(n3649), .A2(n3519), .ZN(n6269) );
  NAND2_X1 U3495 ( .A1(n3295), .A2(n3309), .ZN(n4031) );
  NAND2_X1 U3496 ( .A1(n3263), .A2(n3262), .ZN(n3910) );
  NOR2_X2 U3497 ( .A1(n3005), .A2(n4719), .ZN(n4787) );
  OR2_X1 U3498 ( .A1(n3280), .A2(n3279), .ZN(n3241) );
  NAND2_X2 U3499 ( .A1(n3273), .A2(n3272), .ZN(n4398) );
  CLKBUF_X1 U3500 ( .A(n3739), .Z(n5306) );
  NAND2_X1 U3501 ( .A1(n3124), .A2(n3123), .ZN(n3178) );
  CLKBUF_X1 U3502 ( .A(n3154), .Z(n3246) );
  AOI21_X1 U3503 ( .B1(n3016), .B2(n3144), .A(n4452), .ZN(n3126) );
  NAND2_X1 U3504 ( .A1(n3612), .A2(n3538), .ZN(n3941) );
  NAND2_X1 U3505 ( .A1(n3118), .A2(n3117), .ZN(n3144) );
  AND2_X1 U3506 ( .A1(n3113), .A2(n3848), .ZN(n3136) );
  NOR2_X1 U3507 ( .A1(n3846), .A2(n5106), .ZN(n3625) );
  AND2_X1 U3508 ( .A1(n3039), .A2(n3038), .ZN(n3116) );
  AND4_X1 U3509 ( .A1(n3085), .A2(n3084), .A3(n3083), .A4(n3082), .ZN(n3101)
         );
  AND4_X1 U3510 ( .A1(n3037), .A2(n3036), .A3(n3035), .A4(n3034), .ZN(n3038)
         );
  AND4_X1 U3511 ( .A1(n3033), .A2(n3032), .A3(n3031), .A4(n3030), .ZN(n3039)
         );
  BUF_X2 U3512 ( .A(n3181), .Z(n5194) );
  INV_X2 U3513 ( .A(n6238), .ZN(n2997) );
  INV_X2 U3514 ( .A(n6142), .ZN(n6746) );
  BUF_X2 U3515 ( .A(n3165), .Z(n5184) );
  BUF_X2 U3516 ( .A(n3198), .Z(n5186) );
  BUF_X2 U3517 ( .A(n3197), .Z(n3000) );
  AND2_X2 U3518 ( .A1(n3892), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3898)
         );
  NOR2_X2 U3519 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4010) );
  AND2_X2 U3520 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3993) );
  AND2_X2 U3521 ( .A1(n4666), .A2(n4665), .ZN(n4763) );
  AND2_X4 U3522 ( .A1(n3022), .A2(n3893), .ZN(n3166) );
  AND2_X4 U3523 ( .A1(n3893), .A2(n3023), .ZN(n3197) );
  NAND2_X2 U3524 ( .A1(n5413), .A2(n5089), .ZN(n5867) );
  AND2_X2 U3525 ( .A1(n5417), .A2(n5416), .ZN(n5419) );
  NAND2_X4 U3526 ( .A1(n4890), .A2(n4889), .ZN(n5479) );
  NAND2_X2 U3527 ( .A1(n4785), .A2(n4784), .ZN(n4890) );
  AOI211_X2 U3528 ( .C1(n6204), .C2(n5578), .A(n5577), .B(n5576), .ZN(n5579)
         );
  AOI211_X2 U3529 ( .C1(n6204), .C2(n5286), .A(n5282), .B(n5281), .ZN(n5283)
         );
  AND2_X2 U3530 ( .A1(n5371), .A2(n4823), .ZN(n4822) );
  NOR2_X4 U3531 ( .A1(n5369), .A2(n5368), .ZN(n5371) );
  OR2_X2 U3532 ( .A1(n3111), .A2(n3110), .ZN(n3003) );
  NOR2_X4 U3533 ( .A1(n5472), .A2(n3587), .ZN(n5461) );
  OR2_X4 U3534 ( .A1(n5485), .A2(n5387), .ZN(n5472) );
  BUF_X2 U3535 ( .A(n3619), .Z(n5324) );
  OR2_X1 U3536 ( .A1(n3111), .A2(n3110), .ZN(n3004) );
  NOR2_X4 U3537 ( .A1(n5097), .A2(n5096), .ZN(n5417) );
  OR3_X4 U3538 ( .A1(n5429), .A2(n3594), .A3(n3593), .ZN(n5097) );
  NAND2_X1 U3539 ( .A1(n3324), .A2(n3323), .ZN(n3350) );
  NAND3_X1 U3540 ( .A1(n3152), .A2(n3151), .A3(n3150), .ZN(n3222) );
  CLKBUF_X1 U3541 ( .A(n3188), .Z(n5188) );
  OR2_X1 U3542 ( .A1(n3172), .A2(n3171), .ZN(n3264) );
  NAND2_X1 U3543 ( .A1(n4355), .A2(n4354), .ZN(n4376) );
  XNOR2_X1 U3544 ( .A(n3394), .B(n3384), .ZN(n4252) );
  NAND2_X1 U3545 ( .A1(n3394), .A2(n3371), .ZN(n4243) );
  NAND2_X1 U3546 ( .A1(n3370), .A2(n3351), .ZN(n4050) );
  AND2_X1 U3547 ( .A1(n3649), .A2(n3644), .ZN(n3659) );
  NAND2_X1 U3548 ( .A1(n3455), .A2(n3251), .ZN(n3474) );
  NAND2_X1 U3549 ( .A1(n3153), .A2(n3222), .ZN(n3243) );
  OR2_X1 U3550 ( .A1(n4452), .A2(n6540), .ZN(n3251) );
  NOR2_X1 U3551 ( .A1(n4213), .A2(n3645), .ZN(n3871) );
  NOR2_X1 U3552 ( .A1(n4922), .A2(n5575), .ZN(n5040) );
  INV_X1 U3553 ( .A(n4248), .ZN(n4249) );
  NAND2_X1 U3554 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n4249), .ZN(n4349)
         );
  NOR2_X2 U3555 ( .A1(n4256), .A2(n4253), .ZN(n4355) );
  OAI21_X1 U3556 ( .B1(n5587), .B2(n5588), .A(n5239), .ZN(n5582) );
  AND2_X1 U3557 ( .A1(n4812), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3513) );
  INV_X1 U3558 ( .A(n6131), .ZN(n6122) );
  AND2_X1 U3559 ( .A1(n6131), .A2(n3782), .ZN(n5511) );
  CLKBUF_X1 U3560 ( .A(n3188), .Z(n5029) );
  AND2_X2 U3561 ( .A1(n3997), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3024)
         );
  OR2_X1 U3562 ( .A1(n3195), .A2(n3194), .ZN(n3395) );
  INV_X1 U3563 ( .A(n3270), .ZN(n3214) );
  OR2_X1 U3564 ( .A1(n3634), .A2(n3138), .ZN(n3177) );
  OR2_X1 U3565 ( .A1(n4452), .A2(n3452), .ZN(n3675) );
  NAND2_X1 U3566 ( .A1(n4763), .A2(n4762), .ZN(n4771) );
  NAND2_X1 U3567 ( .A1(n4502), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4650)
         );
  NAND2_X1 U3568 ( .A1(n5571), .A2(n5243), .ZN(n5245) );
  NAND2_X1 U3569 ( .A1(n3930), .A2(n3935), .ZN(n3565) );
  OR2_X1 U3570 ( .A1(n3211), .A2(n3210), .ZN(n3285) );
  XNOR2_X1 U3571 ( .A(n3176), .B(n3175), .ZN(n3294) );
  INV_X1 U3572 ( .A(n3281), .ZN(n3282) );
  OAI21_X1 U3573 ( .B1(n6546), .B2(n4028), .A(n6423), .ZN(n3920) );
  XNOR2_X1 U3575 ( .A(n3178), .B(n3177), .ZN(n3739) );
  OR2_X1 U3576 ( .A1(n3808), .A2(n3807), .ZN(n3816) );
  OR2_X1 U3577 ( .A1(n5143), .A2(n5142), .ZN(n5145) );
  AND2_X1 U3578 ( .A1(n5072), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4831)
         );
  NAND2_X1 U3579 ( .A1(n4831), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5139)
         );
  AND2_X1 U3580 ( .A1(n4438), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5059)
         );
  NAND2_X1 U3581 ( .A1(n5040), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5052)
         );
  INV_X1 U3582 ( .A(n4938), .ZN(n4437) );
  NAND2_X1 U3583 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n4436), .ZN(n4938)
         );
  INV_X1 U3584 ( .A(n5018), .ZN(n4436) );
  NOR2_X1 U3585 ( .A1(n4942), .A2(n5972), .ZN(n5019) );
  NAND2_X1 U3586 ( .A1(n5019), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5018)
         );
  AND2_X1 U3587 ( .A1(n5456), .A2(n5455), .ZN(n5467) );
  OR2_X1 U3588 ( .A1(n5480), .A2(n5386), .ZN(n5468) );
  NOR2_X1 U3589 ( .A1(n4650), .A2(n4651), .ZN(n4726) );
  AOI21_X1 U3590 ( .B1(n4252), .B2(n4998), .A(n4251), .ZN(n4253) );
  AOI21_X1 U3591 ( .B1(n4247), .B2(n4998), .A(n4246), .ZN(n4259) );
  OR2_X1 U3592 ( .A1(n4258), .A2(n4259), .ZN(n4256) );
  AOI21_X1 U3593 ( .B1(n4056), .B2(n4998), .A(n4055), .ZN(n4059) );
  INV_X1 U3594 ( .A(n4050), .ZN(n4056) );
  NAND2_X1 U3595 ( .A1(n4058), .A2(n4057), .ZN(n4258) );
  INV_X1 U3596 ( .A(n4059), .ZN(n4057) );
  INV_X1 U3597 ( .A(n4060), .ZN(n4058) );
  NOR2_X1 U3598 ( .A1(n3757), .A2(n3756), .ZN(n3812) );
  INV_X1 U3599 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3756) );
  NAND2_X1 U3600 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3757) );
  NAND2_X1 U3601 ( .A1(n5419), .A2(n5112), .ZN(n5250) );
  AND2_X1 U3602 ( .A1(n5602), .A2(n3417), .ZN(n3418) );
  CLKBUF_X1 U3603 ( .A(n5592), .Z(n5597) );
  AND2_X1 U3604 ( .A1(n2996), .A2(n5610), .ZN(n3414) );
  NAND2_X1 U3605 ( .A1(n5483), .A2(n5482), .ZN(n5485) );
  CLKBUF_X1 U3606 ( .A(n4710), .Z(n4711) );
  CLKBUF_X1 U3607 ( .A(n4514), .Z(n4569) );
  NAND2_X1 U3608 ( .A1(n4158), .A2(n4159), .ZN(n4236) );
  AND2_X1 U3609 ( .A1(n3514), .A2(n6435), .ZN(n3649) );
  NAND2_X1 U3610 ( .A1(n4681), .A2(n6540), .ZN(n3263) );
  CLKBUF_X1 U3611 ( .A(n3911), .Z(n4098) );
  NAND2_X1 U3612 ( .A1(n3245), .A2(n3244), .ZN(n4012) );
  AND2_X1 U3613 ( .A1(n2995), .A2(n4468), .ZN(n4041) );
  INV_X1 U3614 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U3615 ( .A1(n3250), .A2(n3249), .ZN(n4671) );
  AND3_X1 U3616 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6540), .A3(n3920), .ZN(
        n3980) );
  INV_X1 U3617 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n5725) );
  AND2_X1 U3618 ( .A1(n6050), .A2(n4443), .ZN(n6079) );
  NAND2_X1 U3619 ( .A1(n6533), .A2(n4455), .ZN(n6090) );
  AND2_X1 U3620 ( .A1(n5226), .A2(n4449), .ZN(n6088) );
  INV_X1 U3621 ( .A(n6107), .ZN(n6103) );
  INV_X1 U3622 ( .A(n5399), .ZN(n5486) );
  AND2_X1 U3623 ( .A1(n3773), .A2(n3772), .ZN(n3779) );
  INV_X1 U3624 ( .A(n5511), .ZN(n6126) );
  CLKBUF_X1 U3625 ( .A(n6178), .Z(n6164) );
  AND2_X1 U3626 ( .A1(n5448), .A2(n5447), .ZN(n6113) );
  AND2_X1 U3627 ( .A1(n5481), .A2(n5480), .ZN(n5999) );
  INV_X1 U3628 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U3629 ( .A1(n6208), .A2(n5627), .ZN(n6225) );
  AND2_X1 U3630 ( .A1(n5665), .A2(n3661), .ZN(n5660) );
  OR2_X1 U3631 ( .A1(n5682), .A2(n3668), .ZN(n5668) );
  NOR2_X1 U3632 ( .A1(n6226), .A2(n5898), .ZN(n5911) );
  INV_X1 U3633 ( .A(n6288), .ZN(n6303) );
  CLKBUF_X1 U3634 ( .A(n4619), .Z(n5723) );
  INV_X1 U3635 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n4812) );
  NAND2_X1 U3636 ( .A1(n4213), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6423) );
  INV_X1 U3637 ( .A(n5758), .ZN(n5717) );
  INV_X1 U3638 ( .A(n4271), .ZN(n5271) );
  INV_X1 U3639 ( .A(n6350), .ZN(n5272) );
  OR2_X1 U3640 ( .A1(n3952), .A2(n4084), .ZN(n6333) );
  INV_X1 U3641 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6540) );
  INV_X1 U3642 ( .A(n3522), .ZN(n3520) );
  OR2_X2 U3643 ( .A1(n6015), .A2(n6014), .ZN(n3005) );
  NOR2_X4 U3644 ( .A1(n3678), .A2(n4447), .ZN(n6089) );
  INV_X2 U3645 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3882) );
  OR2_X1 U3646 ( .A1(n3663), .A2(n3662), .ZN(n3006) );
  AND4_X1 U3647 ( .A1(n3021), .A2(n3020), .A3(n3019), .A4(n3018), .ZN(n3007)
         );
  NAND2_X1 U3648 ( .A1(n3160), .A2(n3159), .ZN(n3244) );
  NOR2_X1 U3649 ( .A1(n4591), .A2(n3823), .ZN(n3008) );
  OR2_X1 U3650 ( .A1(n5241), .A2(n6567), .ZN(n3009) );
  AND2_X1 U3651 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3010) );
  NOR2_X1 U3652 ( .A1(n4098), .A2(n4097), .ZN(n3011) );
  NOR2_X1 U3653 ( .A1(n5545), .A2(n5546), .ZN(n3012) );
  OR2_X1 U3654 ( .A1(n3941), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3013)
         );
  OR2_X1 U3655 ( .A1(n3147), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3014)
         );
  NOR2_X1 U3656 ( .A1(n3219), .A2(n3285), .ZN(n3015) );
  AND2_X1 U3657 ( .A1(n3141), .A2(n3675), .ZN(n3016) );
  NOR2_X1 U3658 ( .A1(n4582), .A2(n3453), .ZN(n3479) );
  OR2_X1 U3659 ( .A1(n3470), .A2(n3469), .ZN(n3477) );
  AND2_X1 U3660 ( .A1(n6388), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3464)
         );
  OR2_X1 U3661 ( .A1(n3234), .A2(n3233), .ZN(n3284) );
  AND2_X1 U3662 ( .A1(n3765), .A2(n5107), .ZN(n3061) );
  OAI21_X1 U3663 ( .B1(n3119), .B2(n3126), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3121) );
  INV_X1 U3664 ( .A(n5052), .ZN(n4438) );
  AND2_X1 U3665 ( .A1(n3310), .A2(n3910), .ZN(n3324) );
  NAND2_X1 U3666 ( .A1(n3348), .A2(n3347), .ZN(n3370) );
  OR2_X1 U3667 ( .A1(n3515), .A2(n3565), .ZN(n3848) );
  AND2_X1 U3668 ( .A1(n3273), .A2(n3392), .ZN(n3281) );
  AND2_X1 U3669 ( .A1(n3801), .A2(n3565), .ZN(n3598) );
  MUX2_X1 U3670 ( .A(n3615), .B(n3530), .S(EBX_REG_1__SCAN_IN), .Z(n3525) );
  INV_X1 U3671 ( .A(n5439), .ZN(n3621) );
  AND2_X1 U3672 ( .A1(n3536), .A2(n3535), .ZN(n4588) );
  OR2_X1 U3673 ( .A1(n5139), .A2(n5539), .ZN(n5143) );
  AND2_X1 U3674 ( .A1(n6185), .A2(n5882), .ZN(n3407) );
  INV_X1 U3675 ( .A(n5158), .ZN(n5064) );
  OR2_X1 U3676 ( .A1(n3324), .A2(n3323), .ZN(n3325) );
  AND2_X1 U3677 ( .A1(n3930), .A2(n3979), .ZN(n3459) );
  AND2_X1 U3678 ( .A1(n3133), .A2(n5107), .ZN(n3141) );
  AND3_X1 U3679 ( .A1(n3950), .A2(n4452), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3489) );
  AND2_X2 U3680 ( .A1(n3993), .A2(n4007), .ZN(n3205) );
  AOI21_X1 U3681 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n3015), .A(n3214), .ZN(
        n3215) );
  INV_X1 U3682 ( .A(n3598), .ZN(n3608) );
  AND2_X1 U3683 ( .A1(n4801), .A2(n3621), .ZN(n4797) );
  INV_X1 U3684 ( .A(n3615), .ZN(n3618) );
  NAND2_X2 U3685 ( .A1(n3526), .A2(n3520), .ZN(n3615) );
  INV_X1 U3686 ( .A(n3112), .ZN(n5108) );
  INV_X1 U3687 ( .A(n5064), .ZN(n5220) );
  NAND2_X1 U3688 ( .A1(n5059), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5062)
         );
  AND2_X1 U3689 ( .A1(n3406), .A2(n5883), .ZN(n5882) );
  AND2_X1 U3690 ( .A1(n4435), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4502)
         );
  INV_X1 U3691 ( .A(n4243), .ZN(n4247) );
  INV_X1 U3692 ( .A(n3459), .ZN(n3488) );
  AND2_X1 U3693 ( .A1(n3142), .A2(n3141), .ZN(n3143) );
  INV_X1 U3694 ( .A(n3243), .ZN(n3245) );
  AOI22_X1 U3695 ( .A1(n3182), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3196), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3079) );
  AND4_X1 U3696 ( .A1(n3028), .A2(n3027), .A3(n3026), .A4(n3025), .ZN(n3029)
         );
  XNOR2_X1 U3697 ( .A(n3283), .B(n3282), .ZN(n3733) );
  OR2_X1 U3698 ( .A1(n3238), .A2(n3213), .ZN(n3270) );
  OAI21_X1 U3699 ( .B1(n3739), .B2(STATE2_REG_0__SCAN_IN), .A(n3215), .ZN(
        n3218) );
  INV_X1 U3700 ( .A(n4452), .ZN(n3638) );
  NOR2_X1 U3701 ( .A1(n4981), .A2(n5395), .ZN(n4957) );
  NAND2_X1 U3702 ( .A1(n3812), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n4051)
         );
  INV_X1 U3703 ( .A(n6091), .ZN(n6073) );
  OR2_X1 U3704 ( .A1(n6533), .A2(n4434), .ZN(n6050) );
  OR2_X1 U3705 ( .A1(n3619), .A2(n5289), .ZN(n4801) );
  NAND2_X1 U3706 ( .A1(n3116), .A2(n3112), .ZN(n3780) );
  INV_X1 U3707 ( .A(n5145), .ZN(n5181) );
  INV_X1 U3708 ( .A(n5062), .ZN(n5072) );
  NAND2_X1 U3709 ( .A1(n4437), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4922)
         );
  NOR2_X1 U3710 ( .A1(n4764), .A2(n6006), .ZN(n4987) );
  OR2_X1 U3711 ( .A1(n4514), .A2(n3403), .ZN(n6183) );
  NOR2_X1 U3712 ( .A1(n6658), .A2(n4349), .ZN(n4435) );
  OAI21_X1 U3713 ( .B1(n3808), .B2(n3488), .A(n3332), .ZN(n3334) );
  NAND2_X1 U3714 ( .A1(n3423), .A2(n3422), .ZN(n3425) );
  NAND2_X1 U3715 ( .A1(n2996), .A2(n5688), .ZN(n5244) );
  OR2_X1 U3716 ( .A1(n5582), .A2(n5240), .ZN(n5571) );
  NAND2_X1 U3717 ( .A1(n3222), .A2(n3221), .ZN(n3223) );
  INV_X1 U3718 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3892) );
  AND2_X1 U3719 ( .A1(n3881), .A2(n3880), .ZN(n6391) );
  OR2_X1 U3720 ( .A1(n4039), .A2(n4038), .ZN(n4130) );
  NAND2_X1 U3721 ( .A1(n3007), .A2(n3029), .ZN(n3112) );
  OR2_X1 U3722 ( .A1(n4095), .A2(n2995), .ZN(n4103) );
  NAND2_X1 U3723 ( .A1(n3218), .A2(n3269), .ZN(n3273) );
  AND2_X2 U3724 ( .A1(n3452), .A2(n4452), .ZN(n6537) );
  AND2_X1 U3725 ( .A1(n6050), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6091) );
  AND2_X1 U3726 ( .A1(n6050), .A2(n4442), .ZN(n6032) );
  NOR2_X1 U3727 ( .A1(n4051), .A2(n6209), .ZN(n4244) );
  AND2_X1 U3728 ( .A1(n4889), .A2(n4772), .ZN(n4785) );
  AND2_X1 U3729 ( .A1(n6111), .A2(n5489), .ZN(n6107) );
  NAND2_X1 U3730 ( .A1(n5325), .A2(n5280), .ZN(n5312) );
  AND2_X1 U3731 ( .A1(n6131), .A2(n5109), .ZN(n6123) );
  NAND2_X1 U3732 ( .A1(n3816), .A2(n3815), .ZN(n3818) );
  AND2_X1 U3733 ( .A1(n3699), .A2(n3698), .ZN(n6145) );
  AND2_X1 U3734 ( .A1(n5415), .A2(n5414), .ZN(n5864) );
  AOI21_X1 U3735 ( .B1(n5428), .B2(n5427), .A(n5426), .ZN(n5871) );
  AOI21_X1 U3736 ( .B1(n5469), .B2(n5468), .A(n5467), .ZN(n6121) );
  INV_X1 U3737 ( .A(n6225), .ZN(n6204) );
  NAND2_X1 U3738 ( .A1(n3501), .A2(n3500), .ZN(n4213) );
  INV_X1 U3739 ( .A(n6208), .ZN(n6218) );
  BUF_X1 U3740 ( .A(n4790), .Z(n5525) );
  AND2_X1 U3741 ( .A1(n5245), .A2(n5244), .ZN(n5564) );
  INV_X1 U3742 ( .A(n5245), .ZN(n5572) );
  OR2_X1 U3743 ( .A1(n6434), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4216) );
  NAND2_X1 U3744 ( .A1(n3381), .A2(n3380), .ZN(n4230) );
  OR2_X1 U3745 ( .A1(n5916), .A2(n3798), .ZN(n6236) );
  AND2_X1 U3746 ( .A1(n3649), .A2(n3628), .ZN(n6288) );
  NAND2_X1 U3747 ( .A1(n6540), .A2(n3920), .ZN(n4275) );
  INV_X1 U3748 ( .A(n4560), .ZN(n4524) );
  INV_X1 U3749 ( .A(n6331), .ZN(n4557) );
  NOR2_X1 U3750 ( .A1(n4130), .A2(n2995), .ZN(n4136) );
  OAI21_X1 U3751 ( .B1(n5726), .B2(n5725), .A(n5724), .ZN(n5754) );
  OR2_X1 U3752 ( .A1(n4676), .A2(n4675), .ZN(n4703) );
  INV_X1 U3753 ( .A(n4398), .ZN(n4468) );
  INV_X1 U3754 ( .A(n6088), .ZN(n6065) );
  OAI21_X1 U3755 ( .B1(n3822), .B2(n3821), .A(n3820), .ZN(n6111) );
  INV_X1 U3756 ( .A(n5522), .ZN(n5495) );
  OAI21_X1 U3757 ( .B1(n5359), .B2(n5358), .A(n5357), .ZN(n5548) );
  OR2_X1 U3758 ( .A1(n5438), .A2(n5437), .ZN(n5858) );
  NAND2_X1 U3759 ( .A1(n3779), .A2(n3778), .ZN(n6131) );
  OR2_X1 U3760 ( .A1(n6145), .A2(n6746), .ZN(n6750) );
  NAND2_X1 U3761 ( .A1(n6195), .A2(n4217), .ZN(n6208) );
  AND2_X1 U3762 ( .A1(n5932), .A2(n5915), .ZN(n6226) );
  INV_X1 U3763 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U3764 ( .A1(n4136), .A2(n4398), .ZN(n4649) );
  OR2_X1 U3765 ( .A1(n4095), .A2(n4083), .ZN(n6386) );
  OR2_X1 U3766 ( .A1(n4095), .A2(n4084), .ZN(n6352) );
  AND2_X1 U3767 ( .A1(n6422), .A2(n6421), .ZN(n6522) );
  AND2_X2 U3768 ( .A1(n3024), .A2(n4010), .ZN(n3182) );
  AND2_X2 U3769 ( .A1(n3882), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3022)
         );
  AOI22_X1 U3771 ( .A1(n3182), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3196), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3021) );
  AND2_X2 U3772 ( .A1(n3024), .A2(n3898), .ZN(n3187) );
  AND2_X2 U3774 ( .A1(n3023), .A2(n3993), .ZN(n3165) );
  AOI22_X1 U3775 ( .A1(n3187), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3165), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3020) );
  AOI22_X1 U3776 ( .A1(n3179), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3205), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3019) );
  INV_X2 U3777 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3017) );
  AND2_X2 U3778 ( .A1(n3017), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3893)
         );
  AND2_X2 U3779 ( .A1(n3023), .A2(n4010), .ZN(n3198) );
  AOI22_X1 U3780 ( .A1(n3166), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3018) );
  AND2_X2 U3781 ( .A1(n3022), .A2(n3993), .ZN(n3189) );
  AND2_X2 U3782 ( .A1(n3022), .A2(n4010), .ZN(n3180) );
  AOI22_X1 U3783 ( .A1(n3189), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3028) );
  AND2_X2 U3784 ( .A1(n3024), .A2(n3893), .ZN(n3203) );
  AND2_X4 U3785 ( .A1(n3893), .A2(n4007), .ZN(n3181) );
  AOI22_X1 U3786 ( .A1(n3203), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3181), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3027) );
  AND2_X2 U3787 ( .A1(n3898), .A2(n4007), .ZN(n3204) );
  AOI22_X1 U3788 ( .A1(n3204), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3026) );
  AND2_X4 U3789 ( .A1(n3024), .A2(n3993), .ZN(n5196) );
  AND2_X2 U3790 ( .A1(n4010), .A2(n4007), .ZN(n3188) );
  AOI22_X1 U3791 ( .A1(n5196), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3025) );
  AOI22_X1 U3792 ( .A1(n3189), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3033) );
  AOI22_X1 U3793 ( .A1(n3203), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3181), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3032) );
  AOI22_X1 U3794 ( .A1(n3204), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3031) );
  AOI22_X1 U3795 ( .A1(n5196), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3030) );
  AOI22_X1 U3796 ( .A1(n3182), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3196), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3037) );
  AOI22_X1 U3797 ( .A1(n3187), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3165), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3036) );
  AOI22_X1 U3798 ( .A1(n3166), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3035) );
  AOI22_X1 U3799 ( .A1(n3179), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3205), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3034) );
  AOI22_X1 U3800 ( .A1(n3182), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3196), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3043) );
  AOI22_X1 U3801 ( .A1(n3179), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3042) );
  AOI22_X1 U3802 ( .A1(n3204), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3041) );
  AOI22_X1 U3803 ( .A1(n3187), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3165), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3040) );
  NAND4_X1 U3804 ( .A1(n3043), .A2(n3042), .A3(n3041), .A4(n3040), .ZN(n3049)
         );
  AOI22_X1 U3805 ( .A1(n3203), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3181), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3047) );
  AOI22_X1 U3806 ( .A1(n3166), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3046) );
  AOI22_X1 U3807 ( .A1(n5196), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3045) );
  AOI22_X1 U3808 ( .A1(n3180), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3205), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3044) );
  NAND4_X1 U3809 ( .A1(n3047), .A2(n3046), .A3(n3045), .A4(n3044), .ZN(n3048)
         );
  OR2_X2 U3810 ( .A1(n3049), .A2(n3048), .ZN(n5107) );
  AOI22_X1 U3811 ( .A1(n3204), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3053) );
  AOI22_X1 U3812 ( .A1(n3203), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3181), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3052) );
  AOI22_X1 U3813 ( .A1(n3189), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3051) );
  AOI22_X1 U3814 ( .A1(n5196), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3050) );
  NAND4_X1 U3815 ( .A1(n3053), .A2(n3052), .A3(n3051), .A4(n3050), .ZN(n3059)
         );
  AOI22_X1 U3816 ( .A1(n3182), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3196), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3057) );
  AOI22_X1 U3817 ( .A1(n3187), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3165), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3056) );
  AOI22_X1 U3818 ( .A1(n3166), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3055) );
  AOI22_X1 U3819 ( .A1(n3179), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3205), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3054) );
  NAND4_X1 U3820 ( .A1(n3057), .A2(n3056), .A3(n3055), .A4(n3054), .ZN(n3058)
         );
  OR2_X2 U3821 ( .A1(n3059), .A2(n3058), .ZN(n3950) );
  OR2_X1 U3822 ( .A1(n3002), .A2(n3950), .ZN(n3060) );
  NAND2_X1 U3823 ( .A1(n3061), .A2(n3060), .ZN(n3129) );
  AOI22_X1 U3824 ( .A1(n3187), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3166), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3065) );
  AOI22_X1 U3825 ( .A1(n3204), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5196), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3064) );
  AOI22_X1 U3826 ( .A1(n3180), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3181), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3063) );
  AOI22_X1 U3827 ( .A1(n3196), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3062) );
  NAND4_X1 U3828 ( .A1(n3065), .A2(n3064), .A3(n3063), .A4(n3062), .ZN(n3071)
         );
  AOI22_X1 U3829 ( .A1(n3203), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3069) );
  AOI22_X1 U3830 ( .A1(n3182), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3165), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3068) );
  AOI22_X1 U3831 ( .A1(n3197), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3067) );
  AOI22_X1 U3832 ( .A1(n3179), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3205), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3066) );
  NAND4_X1 U3833 ( .A1(n3069), .A2(n3068), .A3(n3067), .A4(n3066), .ZN(n3070)
         );
  OR2_X2 U3834 ( .A1(n3071), .A2(n3070), .ZN(n3973) );
  AOI22_X1 U3835 ( .A1(n3189), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3075) );
  AOI22_X1 U3836 ( .A1(n3203), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3181), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3074) );
  AOI22_X1 U3837 ( .A1(n3204), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3073) );
  AOI22_X1 U3838 ( .A1(n5196), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3072) );
  NAND4_X1 U3839 ( .A1(n3075), .A2(n3074), .A3(n3073), .A4(n3072), .ZN(n3081)
         );
  AOI22_X1 U3840 ( .A1(n3187), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3165), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3078) );
  AOI22_X1 U3841 ( .A1(n3166), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3077) );
  AOI22_X1 U3842 ( .A1(n3179), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3205), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3076) );
  NAND4_X1 U3843 ( .A1(n3079), .A2(n3078), .A3(n3077), .A4(n3076), .ZN(n3080)
         );
  OR2_X2 U3844 ( .A1(n3081), .A2(n3080), .ZN(n3935) );
  NAND2_X1 U3845 ( .A1(n3636), .A2(n3935), .ZN(n3629) );
  NAND3_X1 U3846 ( .A1(n3765), .A2(n3624), .A3(n5107), .ZN(n3434) );
  NAND2_X1 U3847 ( .A1(n3182), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3085) );
  NAND2_X1 U3848 ( .A1(n3196), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3084) );
  NAND2_X1 U3849 ( .A1(n3179), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3083) );
  NAND2_X1 U3850 ( .A1(n3205), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3082)
         );
  NAND2_X1 U3851 ( .A1(n3189), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3089) );
  NAND2_X1 U3852 ( .A1(n3203), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3088)
         );
  NAND2_X1 U3853 ( .A1(n3180), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3087) );
  NAND2_X1 U3854 ( .A1(n3181), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3086)
         );
  AND4_X2 U3855 ( .A1(n3089), .A2(n3088), .A3(n3087), .A4(n3086), .ZN(n3100)
         );
  NAND2_X1 U3856 ( .A1(n3204), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3093)
         );
  NAND2_X1 U3857 ( .A1(n5196), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3092)
         );
  NAND2_X1 U3858 ( .A1(n3197), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3091) );
  NAND2_X1 U3859 ( .A1(n3188), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3090)
         );
  NAND2_X1 U3860 ( .A1(n3187), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3097) );
  NAND2_X1 U3861 ( .A1(n3166), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3096) );
  NAND2_X1 U3862 ( .A1(n3165), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3095) );
  NAND2_X1 U3863 ( .A1(n3198), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3094) );
  AND4_X2 U3864 ( .A1(n3097), .A2(n3096), .A3(n3095), .A4(n3094), .ZN(n3098)
         );
  NAND4_X4 U3865 ( .A1(n3101), .A2(n3100), .A3(n3099), .A4(n3098), .ZN(n3930)
         );
  INV_X2 U3866 ( .A(n3930), .ZN(n3452) );
  AOI22_X1 U3867 ( .A1(n3204), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5196), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3105) );
  AOI22_X1 U3868 ( .A1(n3203), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3197), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3104) );
  AOI22_X1 U3869 ( .A1(n3179), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3165), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3103) );
  AOI22_X1 U3870 ( .A1(n3181), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3205), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3102) );
  NAND4_X1 U3871 ( .A1(n3105), .A2(n3104), .A3(n3103), .A4(n3102), .ZN(n3111)
         );
  AOI22_X1 U3872 ( .A1(n3187), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3166), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3109) );
  AOI22_X1 U3873 ( .A1(n3182), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3180), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3108) );
  AOI22_X1 U3874 ( .A1(n3196), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3198), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3107) );
  AOI22_X1 U3875 ( .A1(n3189), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3188), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3106) );
  NAND4_X1 U3876 ( .A1(n3109), .A2(n3108), .A3(n3107), .A4(n3106), .ZN(n3110)
         );
  OR2_X4 U3877 ( .A1(n3111), .A2(n3110), .ZN(n4452) );
  NAND2_X1 U3878 ( .A1(n3434), .A2(n6537), .ZN(n3113) );
  NAND2_X1 U3879 ( .A1(n3624), .A2(n3979), .ZN(n3515) );
  NAND2_X1 U3880 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6458) );
  OAI21_X1 U3881 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6458), .ZN(n3441) );
  NAND2_X1 U3882 ( .A1(n3452), .A2(n3441), .ZN(n3140) );
  NAND2_X1 U3883 ( .A1(n3140), .A2(n5108), .ZN(n3114) );
  NAND3_X1 U3884 ( .A1(n3432), .A2(n3136), .A3(n3114), .ZN(n3119) );
  NAND2_X1 U3885 ( .A1(n3780), .A2(n3935), .ZN(n3133) );
  OAI21_X1 U3886 ( .B1(n3624), .B2(n3921), .A(n3765), .ZN(n3115) );
  NAND2_X1 U3887 ( .A1(n3115), .A2(n3636), .ZN(n3118) );
  NAND2_X1 U3888 ( .A1(n3116), .A2(n5107), .ZN(n3641) );
  NAND4_X1 U3889 ( .A1(n3641), .A2(n3765), .A3(n3624), .A4(n3973), .ZN(n3117)
         );
  NAND2_X1 U3890 ( .A1(n3002), .A2(n3489), .ZN(n3120) );
  NAND2_X1 U3891 ( .A1(n3121), .A2(n3120), .ZN(n3154) );
  NAND2_X1 U3892 ( .A1(n3154), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3124) );
  INV_X1 U3893 ( .A(n3513), .ZN(n3766) );
  NAND2_X1 U3894 ( .A1(n5725), .A2(n4812), .ZN(n6434) );
  INV_X1 U3895 ( .A(n4216), .ZN(n3158) );
  MUX2_X1 U3896 ( .A(n3766), .B(n3158), .S(n6388), .Z(n3122) );
  INV_X1 U3897 ( .A(n3122), .ZN(n3123) );
  NAND2_X1 U3898 ( .A1(n3459), .A2(n3624), .ZN(n3125) );
  NAND2_X1 U3899 ( .A1(n3126), .A2(n3125), .ZN(n3128) );
  NAND2_X1 U3900 ( .A1(n3973), .A2(n4452), .ZN(n3127) );
  NAND2_X1 U3901 ( .A1(n3128), .A2(n3127), .ZN(n3634) );
  NAND2_X1 U3902 ( .A1(n3002), .A2(n3950), .ZN(n3130) );
  NAND2_X1 U3903 ( .A1(n3130), .A2(n3935), .ZN(n3131) );
  OAI21_X1 U3904 ( .B1(n3129), .B2(n3131), .A(n3930), .ZN(n3137) );
  INV_X1 U3905 ( .A(n3641), .ZN(n3738) );
  INV_X1 U3906 ( .A(n3935), .ZN(n3635) );
  OR2_X1 U3907 ( .A1(n6434), .A2(n6540), .ZN(n3132) );
  AOI21_X1 U3908 ( .B1(n3738), .B2(n3635), .A(n3132), .ZN(n3135) );
  NAND2_X1 U3909 ( .A1(n3133), .A2(n6537), .ZN(n3134) );
  NAND4_X1 U3910 ( .A1(n3137), .A2(n3136), .A3(n3135), .A4(n3134), .ZN(n3138)
         );
  NAND2_X1 U3911 ( .A1(n3178), .A2(n3177), .ZN(n3220) );
  INV_X1 U3912 ( .A(n3629), .ZN(n3286) );
  NAND4_X1 U3913 ( .A1(n3738), .A2(n3286), .A3(n3624), .A4(n3002), .ZN(n3847)
         );
  NOR2_X2 U3914 ( .A1(n3847), .A2(n3638), .ZN(n3879) );
  NOR2_X2 U3915 ( .A1(n3930), .A2(n4452), .ZN(n4582) );
  NOR2_X1 U3916 ( .A1(n3979), .A2(n3935), .ZN(n3139) );
  NAND3_X1 U3917 ( .A1(n4582), .A2(n3636), .A3(n3139), .ZN(n3846) );
  NAND2_X1 U3918 ( .A1(n3921), .A2(n5107), .ZN(n5106) );
  AOI21_X1 U3919 ( .B1(n3879), .B2(n3140), .A(n3625), .ZN(n3145) );
  NOR2_X1 U3920 ( .A1(n3515), .A2(n4452), .ZN(n3142) );
  NAND2_X1 U3921 ( .A1(n3145), .A2(n5934), .ZN(n3149) );
  XNOR2_X1 U3922 ( .A(n6388), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5768)
         );
  AND2_X1 U3923 ( .A1(n3766), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3146)
         );
  AOI21_X1 U3924 ( .B1(n3158), .B2(n5768), .A(n3146), .ZN(n3151) );
  INV_X1 U3925 ( .A(n3151), .ZN(n3147) );
  AND2_X1 U3926 ( .A1(n3014), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3148) );
  NAND2_X1 U3927 ( .A1(n3149), .A2(n3148), .ZN(n3221) );
  NAND2_X1 U3928 ( .A1(n3220), .A2(n3221), .ZN(n3153) );
  NAND2_X1 U3929 ( .A1(n3149), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3152) );
  NAND2_X1 U3930 ( .A1(n3154), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3150) );
  NAND2_X1 U3931 ( .A1(n3246), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3160) );
  AND2_X1 U3932 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3155) );
  INV_X1 U3933 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6400) );
  NAND2_X1 U3934 ( .A1(n3155), .A2(n6400), .ZN(n4072) );
  INV_X1 U3935 ( .A(n3155), .ZN(n3156) );
  NAND2_X1 U3936 ( .A1(n3156), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3157) );
  NAND2_X1 U3937 ( .A1(n4072), .A2(n3157), .ZN(n4174) );
  AOI22_X1 U3938 ( .A1(n3158), .A2(n4174), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3766), .ZN(n3159) );
  XNOR2_X1 U3939 ( .A(n3243), .B(n3244), .ZN(n3911) );
  NAND2_X1 U3940 ( .A1(n3911), .A2(n6540), .ZN(n3174) );
  NAND2_X1 U3941 ( .A1(n3624), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3455) );
  INV_X1 U3942 ( .A(n3455), .ZN(n3770) );
  AOI22_X1 U3943 ( .A1(n5195), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5189), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3164) );
  AOI22_X1 U3944 ( .A1(n5197), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3163) );
  AOI22_X1 U3945 ( .A1(n2999), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3162) );
  AOI22_X1 U3946 ( .A1(n5024), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3161) );
  NAND4_X1 U3947 ( .A1(n3164), .A2(n3163), .A3(n3162), .A4(n3161), .ZN(n3172)
         );
  INV_X1 U3948 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6724) );
  AOI22_X1 U3949 ( .A1(n5198), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3170) );
  AOI22_X1 U3950 ( .A1(n5185), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3169) );
  AOI22_X1 U3951 ( .A1(n5187), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3168) );
  AOI22_X1 U3952 ( .A1(n5167), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3167) );
  NAND4_X1 U3953 ( .A1(n3170), .A2(n3169), .A3(n3168), .A4(n3167), .ZN(n3171)
         );
  NAND2_X1 U3954 ( .A1(n3770), .A2(n3264), .ZN(n3173) );
  NAND2_X1 U3955 ( .A1(n3174), .A2(n3173), .ZN(n3176) );
  INV_X1 U3956 ( .A(n3251), .ZN(n6544) );
  AOI22_X1 U3957 ( .A1(n6544), .A2(n3264), .B1(n3489), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3175) );
  AOI22_X1 U3958 ( .A1(n5167), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5189), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3186) );
  AOI22_X1 U3959 ( .A1(n2999), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n5024), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3185) );
  AOI22_X1 U3960 ( .A1(n5197), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3184) );
  AOI22_X1 U3961 ( .A1(n5198), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3183) );
  NAND4_X1 U3962 ( .A1(n3186), .A2(n3185), .A3(n3184), .A4(n3183), .ZN(n3195)
         );
  AOI22_X1 U3963 ( .A1(n5185), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5187), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3193) );
  AOI22_X1 U3964 ( .A1(n2998), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3192) );
  AOI22_X1 U3965 ( .A1(n3000), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n5188), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3191) );
  AOI22_X1 U3966 ( .A1(n5195), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3190) );
  NAND4_X1 U3967 ( .A1(n3193), .A2(n3192), .A3(n3191), .A4(n3190), .ZN(n3194)
         );
  NAND2_X1 U3968 ( .A1(n3624), .A2(n3395), .ZN(n3219) );
  AOI22_X1 U3969 ( .A1(n5198), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3202) );
  AOI22_X1 U3970 ( .A1(n5167), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n5189), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3201) );
  AOI22_X1 U3971 ( .A1(n5195), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3200) );
  AOI22_X1 U3972 ( .A1(n5186), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3199) );
  NAND4_X1 U3973 ( .A1(n3202), .A2(n3201), .A3(n3200), .A4(n3199), .ZN(n3211)
         );
  AOI22_X1 U3974 ( .A1(n5197), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n2999), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3209) );
  AOI22_X1 U3975 ( .A1(n5185), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5187), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3208) );
  AOI22_X1 U3976 ( .A1(n5194), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3207) );
  AOI22_X1 U3977 ( .A1(n5024), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5188), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3206) );
  NAND4_X1 U3978 ( .A1(n3209), .A2(n3208), .A3(n3207), .A4(n3206), .ZN(n3210)
         );
  INV_X1 U3979 ( .A(n3395), .ZN(n3212) );
  NAND2_X1 U3980 ( .A1(n3770), .A2(n3212), .ZN(n3238) );
  INV_X1 U3981 ( .A(n3285), .ZN(n3213) );
  INV_X1 U3982 ( .A(n3489), .ZN(n3475) );
  INV_X1 U3983 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3217) );
  AOI21_X1 U3984 ( .B1(n3638), .B2(n3285), .A(n6540), .ZN(n3216) );
  OAI211_X1 U3985 ( .C1(n3475), .C2(n3217), .A(n3216), .B(n3219), .ZN(n3269)
         );
  OR2_X1 U3986 ( .A1(n3219), .A2(n6540), .ZN(n3392) );
  INV_X1 U3987 ( .A(n3220), .ZN(n3224) );
  XNOR2_X2 U3988 ( .A(n3224), .B(n3223), .ZN(n4097) );
  NAND2_X1 U3989 ( .A1(n4097), .A2(n6540), .ZN(n3236) );
  AOI22_X1 U3990 ( .A1(n2998), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n5167), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3228) );
  AOI22_X1 U3991 ( .A1(n2999), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5024), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3227) );
  AOI22_X1 U3992 ( .A1(n5185), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5187), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3226) );
  AOI22_X1 U3993 ( .A1(n5197), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3225) );
  NAND4_X1 U3994 ( .A1(n3228), .A2(n3227), .A3(n3226), .A4(n3225), .ZN(n3234)
         );
  AOI22_X1 U3995 ( .A1(n5198), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5189), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3232) );
  AOI22_X1 U3996 ( .A1(n5195), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3231) );
  AOI22_X1 U3997 ( .A1(n5186), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3230) );
  AOI22_X1 U3998 ( .A1(n3000), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3229) );
  NAND4_X1 U3999 ( .A1(n3232), .A2(n3231), .A3(n3230), .A4(n3229), .ZN(n3233)
         );
  NAND2_X1 U4000 ( .A1(n3770), .A2(n3284), .ZN(n3235) );
  INV_X1 U4001 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3239) );
  NAND2_X1 U4002 ( .A1(n6544), .A2(n3284), .ZN(n3237) );
  OAI211_X1 U4003 ( .C1(n3239), .C2(n3475), .A(n3238), .B(n3237), .ZN(n3279)
         );
  NAND2_X1 U4004 ( .A1(n3280), .A2(n3279), .ZN(n3240) );
  NAND2_X1 U4005 ( .A1(n3281), .A2(n3240), .ZN(n3242) );
  NAND2_X1 U4006 ( .A1(n3246), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3250) );
  NAND3_X1 U4007 ( .A1(n5765), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4268) );
  INV_X1 U4008 ( .A(n4268), .ZN(n3913) );
  NAND2_X1 U4009 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3913), .ZN(n6332) );
  NAND2_X1 U4010 ( .A1(n5765), .A2(n6332), .ZN(n3247) );
  NAND3_X1 U4011 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4395) );
  INV_X1 U4012 ( .A(n4395), .ZN(n4401) );
  NAND2_X1 U4013 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4401), .ZN(n4426) );
  NAND2_X1 U4014 ( .A1(n3247), .A2(n4426), .ZN(n4611) );
  OAI22_X1 U4015 ( .A1(n4216), .A2(n4611), .B1(n3513), .B2(n5765), .ZN(n3248)
         );
  INV_X1 U4016 ( .A(n3248), .ZN(n3249) );
  XNOR2_X2 U4017 ( .A(n4012), .B(n4671), .ZN(n4681) );
  AOI22_X1 U4018 ( .A1(n5185), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5198), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3255) );
  AOI22_X1 U4019 ( .A1(n5167), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5195), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3254) );
  AOI22_X1 U4020 ( .A1(n5197), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U4021 ( .A1(n5024), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3252) );
  NAND4_X1 U4022 ( .A1(n3255), .A2(n3254), .A3(n3253), .A4(n3252), .ZN(n3261)
         );
  AOI22_X1 U4023 ( .A1(n5187), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3259) );
  AOI22_X1 U4024 ( .A1(n2998), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3258) );
  AOI22_X1 U4025 ( .A1(n2999), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4026 ( .A1(n5189), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3256) );
  NAND4_X1 U4027 ( .A1(n3259), .A2(n3258), .A3(n3257), .A4(n3256), .ZN(n3260)
         );
  OR2_X1 U4028 ( .A1(n3261), .A2(n3260), .ZN(n3326) );
  AOI22_X1 U4029 ( .A1(n3474), .A2(n3326), .B1(INSTQUEUE_REG_0__3__SCAN_IN), 
        .B2(n3489), .ZN(n3262) );
  XNOR2_X2 U4030 ( .A(n3309), .B(n3910), .ZN(n4039) );
  NAND2_X1 U4031 ( .A1(n4039), .A2(n3459), .ZN(n3268) );
  NAND2_X1 U4032 ( .A1(n3284), .A2(n3285), .ZN(n3296) );
  INV_X1 U4033 ( .A(n3264), .ZN(n3297) );
  NAND2_X1 U4034 ( .A1(n3296), .A2(n3297), .ZN(n3327) );
  INV_X1 U4035 ( .A(n3326), .ZN(n3265) );
  XNOR2_X1 U4036 ( .A(n3327), .B(n3265), .ZN(n3266) );
  NAND2_X1 U4037 ( .A1(n3266), .A2(n6537), .ZN(n3267) );
  NAND2_X1 U4038 ( .A1(n3268), .A2(n3267), .ZN(n3306) );
  XNOR2_X1 U4039 ( .A(n3306), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4211)
         );
  INV_X1 U4040 ( .A(n4211), .ZN(n3305) );
  INV_X1 U4041 ( .A(n3269), .ZN(n3271) );
  NAND2_X1 U4042 ( .A1(n3271), .A2(n3270), .ZN(n3272) );
  INV_X1 U4043 ( .A(n4398), .ZN(n3274) );
  NAND2_X1 U4044 ( .A1(n3274), .A2(n3459), .ZN(n3277) );
  INV_X1 U4045 ( .A(n6537), .ZN(n3436) );
  NAND2_X1 U4046 ( .A1(n3638), .A2(n3935), .ZN(n3298) );
  OAI21_X1 U4047 ( .B1(n3436), .B2(n3285), .A(n3298), .ZN(n3275) );
  INV_X1 U4048 ( .A(n3275), .ZN(n3276) );
  NAND2_X1 U4049 ( .A1(n3277), .A2(n3276), .ZN(n5626) );
  NAND2_X1 U4050 ( .A1(n5626), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6297)
         );
  XNOR2_X1 U4051 ( .A(n6297), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3795)
         );
  INV_X1 U4052 ( .A(n6297), .ZN(n3278) );
  NAND2_X1 U4053 ( .A1(n3278), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3289)
         );
  INV_X1 U4054 ( .A(n3289), .ZN(n3292) );
  XNOR2_X1 U4055 ( .A(n3280), .B(n3279), .ZN(n3283) );
  NAND2_X1 U4056 ( .A1(n4291), .A2(n3459), .ZN(n3793) );
  OAI21_X1 U4057 ( .B1(n3285), .B2(n3284), .A(n3296), .ZN(n3287) );
  OAI211_X1 U4058 ( .C1(n3287), .C2(n3436), .A(n3286), .B(n3979), .ZN(n3288)
         );
  INV_X1 U4059 ( .A(n3288), .ZN(n3792) );
  AND2_X1 U4060 ( .A1(n3792), .A2(n3289), .ZN(n3290) );
  NAND2_X1 U4061 ( .A1(n3793), .A2(n3290), .ZN(n3291) );
  OAI21_X1 U4062 ( .B1(n3795), .B2(n3292), .A(n3291), .ZN(n6213) );
  OR2_X1 U4063 ( .A1(n3294), .A2(n3293), .ZN(n3295) );
  OAI21_X1 U4064 ( .B1(n3297), .B2(n3296), .A(n3327), .ZN(n3300) );
  INV_X1 U4065 ( .A(n3298), .ZN(n3299) );
  AOI21_X1 U4066 ( .B1(n3300), .B2(n6537), .A(n3299), .ZN(n3301) );
  OAI21_X1 U4067 ( .B1(n4031), .B2(n3488), .A(n3301), .ZN(n3302) );
  NAND2_X1 U4068 ( .A1(n3302), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6210)
         );
  NAND2_X1 U4069 ( .A1(n6213), .A2(n6210), .ZN(n3303) );
  NAND2_X1 U4070 ( .A1(n3303), .A2(n6211), .ZN(n4212) );
  INV_X1 U4071 ( .A(n4212), .ZN(n3304) );
  NAND2_X1 U4072 ( .A1(n3305), .A2(n3304), .ZN(n3308) );
  NAND2_X1 U4073 ( .A1(n3306), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3307)
         );
  NAND2_X1 U4074 ( .A1(n3308), .A2(n3307), .ZN(n4224) );
  INV_X1 U4075 ( .A(n3309), .ZN(n3310) );
  AOI22_X1 U4076 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n5195), .B1(n5189), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3314) );
  AOI22_X1 U4077 ( .A1(n5197), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4078 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n2999), .B1(n3000), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3312) );
  AOI22_X1 U4079 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n5024), .B1(n5029), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3311) );
  NAND4_X1 U4080 ( .A1(n3314), .A2(n3313), .A3(n3312), .A4(n3311), .ZN(n3320)
         );
  AOI22_X1 U4081 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5198), .B1(n2998), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4082 ( .A1(n5185), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U4083 ( .A1(n5187), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4084 ( .A1(n5167), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3315) );
  NAND4_X1 U4085 ( .A1(n3318), .A2(n3317), .A3(n3316), .A4(n3315), .ZN(n3319)
         );
  OR2_X1 U4086 ( .A1(n3320), .A2(n3319), .ZN(n3330) );
  NAND2_X1 U4087 ( .A1(n3474), .A2(n3330), .ZN(n3322) );
  NAND2_X1 U4088 ( .A1(n3489), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3321) );
  NAND2_X1 U4089 ( .A1(n3322), .A2(n3321), .ZN(n3323) );
  NAND2_X1 U4090 ( .A1(n3350), .A2(n3325), .ZN(n3808) );
  NAND2_X1 U4091 ( .A1(n3327), .A2(n3326), .ZN(n3329) );
  INV_X1 U4092 ( .A(n3329), .ZN(n3331) );
  INV_X1 U4093 ( .A(n3330), .ZN(n3328) );
  OR2_X1 U4094 ( .A1(n3329), .A2(n3328), .ZN(n3374) );
  OAI211_X1 U4095 ( .C1(n3331), .C2(n3330), .A(n6537), .B(n3374), .ZN(n3332)
         );
  INV_X1 U4096 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3333) );
  XNOR2_X1 U4097 ( .A(n3334), .B(n3333), .ZN(n4223) );
  NAND2_X1 U4098 ( .A1(n4224), .A2(n4223), .ZN(n3336) );
  NAND2_X1 U4099 ( .A1(n3334), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3335)
         );
  NAND2_X1 U4100 ( .A1(n3336), .A2(n3335), .ZN(n6202) );
  INV_X1 U4101 ( .A(n3350), .ZN(n3348) );
  AOI22_X1 U4102 ( .A1(n5195), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5189), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4103 ( .A1(n5197), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3339) );
  AOI22_X1 U4104 ( .A1(n2999), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U4105 ( .A1(n5024), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3337) );
  NAND4_X1 U4106 ( .A1(n3340), .A2(n3339), .A3(n3338), .A4(n3337), .ZN(n3346)
         );
  AOI22_X1 U4107 ( .A1(n5198), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3344) );
  AOI22_X1 U4108 ( .A1(n5185), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3343) );
  AOI22_X1 U4109 ( .A1(n5187), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3342) );
  AOI22_X1 U4110 ( .A1(n5167), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3341) );
  NAND4_X1 U4111 ( .A1(n3344), .A2(n3343), .A3(n3342), .A4(n3341), .ZN(n3345)
         );
  OR2_X1 U4112 ( .A1(n3346), .A2(n3345), .ZN(n3372) );
  AOI22_X1 U4113 ( .A1(n3474), .A2(n3372), .B1(INSTQUEUE_REG_0__5__SCAN_IN), 
        .B2(n3489), .ZN(n3349) );
  INV_X1 U4114 ( .A(n3349), .ZN(n3347) );
  NAND2_X1 U4115 ( .A1(n3350), .A2(n3349), .ZN(n3351) );
  XNOR2_X1 U4116 ( .A(n3374), .B(n3372), .ZN(n3352) );
  NAND2_X1 U4117 ( .A1(n3352), .A2(n6537), .ZN(n3353) );
  INV_X1 U4118 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3355) );
  XNOR2_X1 U4119 ( .A(n3356), .B(n3355), .ZN(n6201) );
  NAND2_X1 U4120 ( .A1(n6202), .A2(n6201), .ZN(n3358) );
  NAND2_X1 U4121 ( .A1(n3356), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3357)
         );
  AOI22_X1 U4122 ( .A1(n5195), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5189), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3362) );
  AOI22_X1 U4123 ( .A1(n5197), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3361) );
  AOI22_X1 U4124 ( .A1(n2999), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4125 ( .A1(n5024), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3359) );
  NAND4_X1 U4126 ( .A1(n3362), .A2(n3361), .A3(n3360), .A4(n3359), .ZN(n3368)
         );
  AOI22_X1 U4127 ( .A1(n5198), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4128 ( .A1(n5185), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3365) );
  AOI22_X1 U4129 ( .A1(n5187), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4130 ( .A1(n5167), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3363) );
  NAND4_X1 U4131 ( .A1(n3366), .A2(n3365), .A3(n3364), .A4(n3363), .ZN(n3367)
         );
  OR2_X1 U4132 ( .A1(n3368), .A2(n3367), .ZN(n3375) );
  AOI22_X1 U4133 ( .A1(n3474), .A2(n3375), .B1(n3489), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3369) );
  NAND2_X1 U4134 ( .A1(n3370), .A2(n3369), .ZN(n3371) );
  INV_X1 U4135 ( .A(n3372), .ZN(n3373) );
  NOR2_X1 U4136 ( .A1(n3374), .A2(n3373), .ZN(n3376) );
  NAND2_X1 U4137 ( .A1(n3376), .A2(n3375), .ZN(n3397) );
  OAI211_X1 U4138 ( .C1(n3376), .C2(n3375), .A(n3397), .B(n6537), .ZN(n3377)
         );
  OAI21_X1 U4139 ( .B1(n4243), .B2(n3488), .A(n3377), .ZN(n3379) );
  INV_X1 U4140 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3378) );
  XNOR2_X1 U4141 ( .A(n3379), .B(n3378), .ZN(n4156) );
  NAND2_X1 U4142 ( .A1(n4157), .A2(n4156), .ZN(n3381) );
  NAND2_X1 U4143 ( .A1(n3379), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3380)
         );
  INV_X1 U4144 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3383) );
  NAND2_X1 U4145 ( .A1(n3474), .A2(n3395), .ZN(n3382) );
  OAI21_X1 U4146 ( .B1(n3383), .B2(n3475), .A(n3382), .ZN(n3384) );
  NAND2_X1 U4147 ( .A1(n4252), .A2(n3459), .ZN(n3387) );
  XNOR2_X1 U4148 ( .A(n3397), .B(n3395), .ZN(n3385) );
  NAND2_X1 U4149 ( .A1(n3385), .A2(n6537), .ZN(n3386) );
  NAND2_X1 U4150 ( .A1(n3387), .A2(n3386), .ZN(n3389) );
  INV_X1 U4151 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3388) );
  XNOR2_X1 U4152 ( .A(n3389), .B(n3388), .ZN(n4229) );
  NAND2_X1 U4153 ( .A1(n4230), .A2(n4229), .ZN(n3391) );
  NAND2_X1 U4154 ( .A1(n3389), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3390)
         );
  NAND2_X1 U4155 ( .A1(n3391), .A2(n3390), .ZN(n4331) );
  NOR2_X1 U4156 ( .A1(n3392), .A2(n3488), .ZN(n3393) );
  NAND2_X1 U4157 ( .A1(n6537), .A2(n3395), .ZN(n3396) );
  OR2_X1 U4158 ( .A1(n3397), .A2(n3396), .ZN(n3398) );
  NAND2_X1 U4159 ( .A1(n3404), .A2(n3398), .ZN(n3399) );
  INV_X1 U4160 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3553) );
  XNOR2_X1 U4161 ( .A(n3399), .B(n3553), .ZN(n4330) );
  NAND2_X1 U4162 ( .A1(n4331), .A2(n4330), .ZN(n3401) );
  NAND2_X1 U4163 ( .A1(n3399), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3400)
         );
  NAND2_X1 U4164 ( .A1(n3401), .A2(n3400), .ZN(n4514) );
  INV_X1 U4165 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6254) );
  NOR2_X1 U4166 ( .A1(n2996), .A2(n6254), .ZN(n4568) );
  NAND2_X1 U4167 ( .A1(n5241), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4572) );
  INV_X1 U4168 ( .A(n4572), .ZN(n3402) );
  OR2_X1 U4169 ( .A1(n4568), .A2(n3402), .ZN(n3403) );
  INV_X1 U4170 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U4171 ( .A1(n2996), .A2(n6234), .ZN(n6184) );
  INV_X1 U4172 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U4173 ( .A1(n2996), .A2(n6246), .ZN(n4573) );
  NAND2_X1 U4174 ( .A1(n2996), .A2(n6254), .ZN(n4570) );
  AND2_X1 U4175 ( .A1(n4573), .A2(n4570), .ZN(n6182) );
  AND2_X1 U4176 ( .A1(n6184), .A2(n6182), .ZN(n3405) );
  NAND2_X1 U4177 ( .A1(n6183), .A2(n3405), .ZN(n4710) );
  NAND2_X1 U4178 ( .A1(n5241), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6185) );
  INV_X1 U4179 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3646) );
  XOR2_X1 U4180 ( .A(n5241), .B(n3646), .Z(n5885) );
  INV_X1 U4181 ( .A(n5885), .ZN(n3406) );
  NAND2_X1 U4182 ( .A1(n5241), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5883) );
  NAND2_X1 U4183 ( .A1(n4710), .A2(n3407), .ZN(n3410) );
  INV_X1 U4184 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6714) );
  NAND2_X1 U4185 ( .A1(n2996), .A2(n6714), .ZN(n5880) );
  NAND2_X1 U4186 ( .A1(n2996), .A2(n3646), .ZN(n3408) );
  AND2_X1 U4187 ( .A1(n5880), .A2(n3408), .ZN(n3409) );
  NAND2_X1 U4188 ( .A1(n3410), .A2(n3409), .ZN(n5618) );
  NAND2_X1 U4189 ( .A1(n5241), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3411) );
  NAND2_X1 U4190 ( .A1(n5618), .A2(n3411), .ZN(n3413) );
  INV_X1 U4191 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5914) );
  NAND2_X1 U4192 ( .A1(n2996), .A2(n5914), .ZN(n3412) );
  NAND2_X1 U4193 ( .A1(n3413), .A2(n3412), .ZN(n5594) );
  NAND2_X1 U4194 ( .A1(n5241), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3415) );
  INV_X1 U4195 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5610) );
  AOI21_X2 U4196 ( .B1(n5594), .B2(n3415), .A(n3414), .ZN(n5604) );
  INV_X1 U4197 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3582) );
  NAND2_X1 U4198 ( .A1(n2996), .A2(n3582), .ZN(n5601) );
  NAND2_X1 U4199 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3667) );
  NAND2_X1 U4200 ( .A1(n2996), .A2(n3667), .ZN(n3416) );
  NAND2_X1 U4201 ( .A1(n5592), .A2(n3416), .ZN(n5555) );
  NAND2_X1 U4202 ( .A1(n5241), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5602) );
  OAI21_X1 U4203 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5241), .ZN(n3417) );
  NAND2_X2 U4204 ( .A1(n5555), .A2(n3418), .ZN(n5587) );
  AND2_X1 U4205 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5694) );
  AND2_X1 U4206 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5676) );
  AND2_X1 U4207 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3660) );
  NAND3_X1 U4208 ( .A1(n5694), .A2(n5676), .A3(n3660), .ZN(n3419) );
  NAND2_X1 U4209 ( .A1(n2996), .A2(n3419), .ZN(n3420) );
  NAND2_X1 U4210 ( .A1(n5587), .A2(n3420), .ZN(n3423) );
  NOR2_X1 U4211 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5693) );
  NOR2_X1 U4212 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5252) );
  NOR2_X1 U4213 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5675) );
  NAND3_X1 U4214 ( .A1(n5693), .A2(n5252), .A3(n5675), .ZN(n3421) );
  NAND2_X1 U4215 ( .A1(n5241), .A2(n3421), .ZN(n3422) );
  INV_X1 U4216 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6649) );
  XNOR2_X1 U4217 ( .A(n2996), .B(n6649), .ZN(n5546) );
  NAND2_X1 U4218 ( .A1(n2996), .A2(n6649), .ZN(n3424) );
  OAI21_X1 U4219 ( .B1(n3425), .B2(n5546), .A(n3424), .ZN(n4790) );
  INV_X1 U4220 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6567) );
  OR2_X2 U4221 ( .A1(n4790), .A2(n3009), .ZN(n5537) );
  NAND2_X1 U4222 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5643) );
  NOR2_X2 U4223 ( .A1(n5537), .A2(n5643), .ZN(n5278) );
  NAND3_X1 U4224 ( .A1(n5278), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3428) );
  NOR2_X1 U4225 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U4226 ( .A1(n5645), .A2(n6567), .ZN(n3426) );
  NOR2_X1 U4227 ( .A1(n2996), .A2(n3426), .ZN(n4791) );
  INV_X1 U4228 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4808) );
  INV_X1 U4229 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5632) );
  NAND4_X1 U4230 ( .A1(n3012), .A2(n4791), .A3(n4808), .A4(n5632), .ZN(n3427)
         );
  NAND2_X1 U4231 ( .A1(n3428), .A2(n3427), .ZN(n3429) );
  XNOR2_X1 U4232 ( .A(n3429), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5268)
         );
  INV_X1 U4233 ( .A(n3674), .ZN(n3686) );
  NAND2_X1 U4234 ( .A1(n3950), .A2(n3979), .ZN(n3430) );
  OR2_X1 U4235 ( .A1(n3641), .A2(n3430), .ZN(n3902) );
  NAND2_X1 U4236 ( .A1(n3902), .A2(n3638), .ZN(n3431) );
  NAND2_X1 U4237 ( .A1(n3432), .A2(n3431), .ZN(n3516) );
  INV_X1 U4238 ( .A(n3002), .ZN(n3433) );
  OR2_X1 U4239 ( .A1(n3434), .A2(n3433), .ZN(n3438) );
  NAND2_X1 U4240 ( .A1(n3002), .A2(n4452), .ZN(n3435) );
  NAND2_X1 U4241 ( .A1(n3436), .A2(n3435), .ZN(n3437) );
  NAND2_X1 U4242 ( .A1(n3438), .A2(n3437), .ZN(n3631) );
  INV_X1 U4243 ( .A(n3631), .ZN(n3439) );
  OR2_X1 U4244 ( .A1(n3516), .A2(n3439), .ZN(n3440) );
  NAND2_X1 U4245 ( .A1(n3686), .A2(n3440), .ZN(n3873) );
  INV_X1 U4246 ( .A(n3847), .ZN(n3626) );
  OR2_X1 U4247 ( .A1(n3441), .A2(STATE_REG_0__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U4248 ( .A1(n3452), .A2(n6539), .ZN(n4454) );
  INV_X1 U4249 ( .A(READY_N), .ZN(n6455) );
  AND2_X1 U4250 ( .A1(n4454), .A2(n6455), .ZN(n3442) );
  NAND2_X1 U4251 ( .A1(n3626), .A2(n3442), .ZN(n3876) );
  NAND3_X1 U4252 ( .A1(n3876), .A2(n4452), .A3(n5106), .ZN(n3502) );
  XNOR2_X1 U4253 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3463) );
  NAND2_X1 U4254 ( .A1(n3464), .A2(n3463), .ZN(n3444) );
  INV_X1 U4255 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6394) );
  NAND2_X1 U4256 ( .A1(n6394), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3443) );
  NAND2_X1 U4257 ( .A1(n3444), .A2(n3443), .ZN(n3473) );
  XNOR2_X1 U4258 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3471) );
  NAND2_X1 U4259 ( .A1(n3473), .A2(n3471), .ZN(n3446) );
  NAND2_X1 U4260 ( .A1(n6400), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3445) );
  NAND2_X1 U4261 ( .A1(n3446), .A2(n3445), .ZN(n3486) );
  XNOR2_X1 U4262 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3484) );
  NAND2_X1 U4263 ( .A1(n3486), .A2(n3484), .ZN(n3448) );
  NAND2_X1 U4264 ( .A1(n5765), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3447) );
  NAND2_X1 U4265 ( .A1(n3448), .A2(n3447), .ZN(n3487) );
  INV_X1 U4266 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6405) );
  AND2_X1 U4267 ( .A1(n6405), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3449)
         );
  OR2_X1 U4268 ( .A1(n3487), .A2(n3449), .ZN(n3451) );
  INV_X1 U4269 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U4270 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n5939), .ZN(n3450) );
  AND2_X1 U4271 ( .A1(n3451), .A2(n3450), .ZN(n3498) );
  NAND2_X1 U4272 ( .A1(n3474), .A2(n3498), .ZN(n3497) );
  AND2_X1 U4273 ( .A1(n3452), .A2(n3979), .ZN(n3453) );
  AND2_X1 U4274 ( .A1(n3017), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3454)
         );
  NOR2_X1 U4275 ( .A1(n3464), .A2(n3454), .ZN(n3458) );
  OAI21_X1 U4276 ( .B1(n3455), .B2(n5108), .A(n3458), .ZN(n3456) );
  NAND2_X1 U4277 ( .A1(n3456), .A2(n4452), .ZN(n3457) );
  NAND2_X1 U4278 ( .A1(n3479), .A2(n3457), .ZN(n3462) );
  NAND2_X1 U4279 ( .A1(n3474), .A2(n3458), .ZN(n3460) );
  NAND2_X1 U4280 ( .A1(n3489), .A2(n3459), .ZN(n3499) );
  NAND2_X1 U4281 ( .A1(n3460), .A2(n3499), .ZN(n3461) );
  NAND2_X1 U4282 ( .A1(n3462), .A2(n3461), .ZN(n3468) );
  AOI21_X1 U4283 ( .B1(n3474), .B2(n3930), .A(n5108), .ZN(n3467) );
  INV_X1 U4284 ( .A(n3463), .ZN(n3465) );
  XNOR2_X1 U4285 ( .A(n3465), .B(n3464), .ZN(n3505) );
  OAI22_X1 U4286 ( .A1(n3468), .A2(n3467), .B1(n3499), .B2(n3505), .ZN(n3470)
         );
  NAND2_X1 U4287 ( .A1(n3505), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3466) );
  AOI21_X1 U4288 ( .B1(n3468), .B2(n3467), .A(n3466), .ZN(n3469) );
  INV_X1 U4289 ( .A(n3471), .ZN(n3472) );
  XNOR2_X1 U4290 ( .A(n3473), .B(n3472), .ZN(n3504) );
  NAND2_X1 U4291 ( .A1(n3474), .A2(n3504), .ZN(n3478) );
  OAI211_X1 U4292 ( .C1(n3504), .C2(n3475), .A(n3479), .B(n3478), .ZN(n3476)
         );
  NAND2_X1 U4293 ( .A1(n3477), .A2(n3476), .ZN(n3483) );
  INV_X1 U4294 ( .A(n3478), .ZN(n3481) );
  INV_X1 U4295 ( .A(n3479), .ZN(n3480) );
  NAND2_X1 U4296 ( .A1(n3481), .A2(n3480), .ZN(n3482) );
  NAND2_X1 U4297 ( .A1(n3483), .A2(n3482), .ZN(n3491) );
  INV_X1 U4298 ( .A(n3491), .ZN(n3494) );
  INV_X1 U4299 ( .A(n3484), .ZN(n3485) );
  XNOR2_X1 U4300 ( .A(n3486), .B(n3485), .ZN(n3506) );
  OR3_X1 U4301 ( .A1(n3487), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(n6405), 
        .ZN(n3503) );
  NAND2_X1 U4302 ( .A1(n3506), .A2(n3503), .ZN(n3493) );
  AOI21_X1 U4303 ( .B1(n3506), .B2(n3503), .A(n3488), .ZN(n3490) );
  OAI21_X1 U4304 ( .B1(n3491), .B2(n3490), .A(n3489), .ZN(n3492) );
  OAI21_X1 U4305 ( .B1(n3494), .B2(n3493), .A(n3492), .ZN(n3495) );
  AOI21_X1 U4306 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6540), .A(n3495), 
        .ZN(n3496) );
  NAND2_X1 U4307 ( .A1(n3497), .A2(n3496), .ZN(n3501) );
  INV_X1 U4308 ( .A(n3498), .ZN(n3508) );
  OR2_X1 U4309 ( .A1(n3499), .A2(n3508), .ZN(n3500) );
  NAND2_X1 U4310 ( .A1(n3502), .A2(n4213), .ZN(n3510) );
  NAND2_X1 U4311 ( .A1(n3930), .A2(n6539), .ZN(n6536) );
  NAND4_X1 U4312 ( .A1(n3506), .A2(n3505), .A3(n3504), .A4(n3503), .ZN(n3507)
         );
  NAND2_X1 U4313 ( .A1(n3508), .A2(n3507), .ZN(n3673) );
  NOR2_X1 U4314 ( .A1(READY_N), .A2(n3673), .ZN(n3774) );
  NAND2_X1 U4315 ( .A1(n6536), .A2(n3774), .ZN(n3509) );
  MUX2_X1 U4316 ( .A(n3510), .B(n3509), .S(n3973), .Z(n3512) );
  INV_X1 U4317 ( .A(n3902), .ZN(n4884) );
  NAND2_X1 U4318 ( .A1(n4884), .A2(n3930), .ZN(n3645) );
  INV_X1 U4319 ( .A(n3871), .ZN(n3511) );
  NAND3_X1 U4320 ( .A1(n3873), .A2(n3512), .A3(n3511), .ZN(n3514) );
  AND2_X1 U4321 ( .A1(n3513), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6435) );
  INV_X1 U4322 ( .A(n4582), .ZN(n3771) );
  NOR2_X1 U4323 ( .A1(n3516), .A2(n3771), .ZN(n3851) );
  INV_X1 U4324 ( .A(n3851), .ZN(n3518) );
  NAND2_X2 U4325 ( .A1(n3003), .A2(n3930), .ZN(n3522) );
  INV_X2 U4326 ( .A(n3522), .ZN(n3801) );
  AOI22_X1 U4327 ( .A1(n3625), .A2(n3950), .B1(n3626), .B2(n3801), .ZN(n3517)
         );
  OR2_X1 U4328 ( .A1(n3516), .A2(n3515), .ZN(n6410) );
  NAND4_X1 U4329 ( .A1(n3518), .A2(n3517), .A3(n5934), .A4(n6410), .ZN(n3519)
         );
  INV_X1 U4330 ( .A(n3565), .ZN(n3526) );
  NAND2_X1 U4331 ( .A1(n3635), .A2(n3004), .ZN(n3530) );
  INV_X1 U4332 ( .A(n3530), .ZN(n3521) );
  NAND2_X1 U4333 ( .A1(n3521), .A2(n3522), .ZN(n3547) );
  NAND3_X1 U4334 ( .A1(n3565), .A2(n3522), .A3(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n3523) );
  AND2_X1 U4335 ( .A1(n3547), .A2(n3523), .ZN(n3524) );
  NAND2_X1 U4336 ( .A1(n3530), .A2(EBX_REG_0__SCAN_IN), .ZN(n3528) );
  INV_X1 U4337 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U4338 ( .A1(n3538), .A2(n5300), .ZN(n3527) );
  NAND2_X1 U4339 ( .A1(n3528), .A2(n3527), .ZN(n3940) );
  NAND2_X1 U4340 ( .A1(n3799), .A2(n3801), .ZN(n3800) );
  NAND2_X2 U4341 ( .A1(n3800), .A2(n3529), .ZN(n4587) );
  MUX2_X1 U4342 ( .A(n3615), .B(n3612), .S(EBX_REG_2__SCAN_IN), .Z(n3533) );
  NAND2_X1 U4343 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n3522), .ZN(n3531)
         );
  AND2_X1 U4344 ( .A1(n3547), .A2(n3531), .ZN(n3532) );
  NAND2_X1 U4345 ( .A1(n3533), .A2(n3532), .ZN(n4589) );
  INV_X1 U4346 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U4347 ( .A1(n3598), .A2(n6112), .ZN(n3536) );
  NAND2_X1 U4348 ( .A1(n3538), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3534)
         );
  OAI211_X1 U4349 ( .C1(n4448), .C2(EBX_REG_3__SCAN_IN), .A(n3612), .B(n3534), 
        .ZN(n3535) );
  NAND2_X1 U4350 ( .A1(n4589), .A2(n4588), .ZN(n3537) );
  NOR2_X4 U4351 ( .A1(n4587), .A2(n3537), .ZN(n3823) );
  INV_X1 U4352 ( .A(n3565), .ZN(n5439) );
  INV_X1 U4353 ( .A(n5439), .ZN(n3538) );
  MUX2_X1 U4354 ( .A(n3608), .B(n3538), .S(EBX_REG_5__SCAN_IN), .Z(n3539) );
  INV_X1 U4355 ( .A(n3539), .ZN(n3541) );
  NOR2_X1 U4356 ( .A1(n3941), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3540)
         );
  NOR2_X1 U4357 ( .A1(n3541), .A2(n3540), .ZN(n4063) );
  MUX2_X1 U4358 ( .A(n3615), .B(n3530), .S(EBX_REG_4__SCAN_IN), .Z(n3544) );
  NAND2_X1 U4359 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n4448), .ZN(n3542)
         );
  AND2_X1 U4360 ( .A1(n3547), .A2(n3542), .ZN(n3543) );
  NAND2_X1 U4361 ( .A1(n3544), .A2(n3543), .ZN(n4064) );
  AND2_X1 U4362 ( .A1(n4063), .A2(n4064), .ZN(n3545) );
  AND2_X2 U4363 ( .A1(n3823), .A2(n3545), .ZN(n4158) );
  MUX2_X1 U4364 ( .A(n3615), .B(n3612), .S(EBX_REG_6__SCAN_IN), .Z(n3549) );
  NAND2_X1 U4365 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4448), .ZN(n3546)
         );
  AND2_X1 U4366 ( .A1(n3547), .A2(n3546), .ZN(n3548) );
  NAND2_X1 U4367 ( .A1(n3549), .A2(n3548), .ZN(n4159) );
  MUX2_X1 U4368 ( .A(n3608), .B(n3621), .S(EBX_REG_7__SCAN_IN), .Z(n3552) );
  INV_X1 U4369 ( .A(n3941), .ZN(n3550) );
  NAND2_X1 U4370 ( .A1(n3550), .A2(n3388), .ZN(n3551) );
  NAND2_X1 U4371 ( .A1(n3552), .A2(n3551), .ZN(n4235) );
  OR2_X2 U4372 ( .A1(n4236), .A2(n4235), .ZN(n4333) );
  INV_X1 U4373 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4358) );
  NAND2_X1 U4374 ( .A1(n3618), .A2(n4358), .ZN(n3557) );
  NAND2_X1 U4375 ( .A1(n3612), .A2(n3553), .ZN(n3555) );
  NAND2_X1 U4376 ( .A1(n3801), .A2(n4358), .ZN(n3554) );
  NAND3_X1 U4377 ( .A1(n3555), .A2(n3621), .A3(n3554), .ZN(n3556) );
  AND2_X1 U4378 ( .A1(n3557), .A2(n3556), .ZN(n4332) );
  OR2_X2 U4379 ( .A1(n4333), .A2(n4332), .ZN(n4382) );
  MUX2_X1 U4380 ( .A(n3608), .B(n3621), .S(EBX_REG_9__SCAN_IN), .Z(n3558) );
  NAND2_X1 U4381 ( .A1(n3013), .A2(n3558), .ZN(n4381) );
  INV_X1 U4382 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4511) );
  NAND2_X1 U4383 ( .A1(n3618), .A2(n4511), .ZN(n3562) );
  NAND2_X1 U4384 ( .A1(n3612), .A2(n6246), .ZN(n3560) );
  NAND2_X1 U4385 ( .A1(n3801), .A2(n4511), .ZN(n3559) );
  NAND3_X1 U4386 ( .A1(n3560), .A2(n3621), .A3(n3559), .ZN(n3561) );
  NAND2_X1 U4387 ( .A1(n3562), .A2(n3561), .ZN(n4508) );
  NAND2_X1 U4388 ( .A1(n4509), .A2(n4508), .ZN(n6015) );
  NAND2_X1 U4389 ( .A1(n3621), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3563) );
  OAI211_X1 U4390 ( .C1(n4448), .C2(EBX_REG_11__SCAN_IN), .A(n3612), .B(n3563), 
        .ZN(n3564) );
  OAI21_X1 U4391 ( .B1(n3608), .B2(EBX_REG_11__SCAN_IN), .A(n3564), .ZN(n6014)
         );
  INV_X1 U4392 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6684) );
  NAND2_X1 U4393 ( .A1(n3618), .A2(n6684), .ZN(n3569) );
  NAND2_X1 U4394 ( .A1(n3612), .A2(n6714), .ZN(n3567) );
  NAND2_X1 U4395 ( .A1(n3801), .A2(n6684), .ZN(n3566) );
  NAND3_X1 U4396 ( .A1(n3567), .A2(n3621), .A3(n3566), .ZN(n3568) );
  AND2_X1 U4397 ( .A1(n3569), .A2(n3568), .ZN(n4719) );
  MUX2_X1 U4398 ( .A(n3608), .B(n3621), .S(EBX_REG_13__SCAN_IN), .Z(n3570) );
  INV_X1 U4399 ( .A(n3570), .ZN(n3572) );
  NOR2_X1 U4400 ( .A1(n3941), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3571)
         );
  NOR2_X1 U4401 ( .A1(n3572), .A2(n3571), .ZN(n4788) );
  AND2_X2 U4402 ( .A1(n4787), .A2(n4788), .ZN(n5483) );
  INV_X1 U4403 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U4404 ( .A1(n3618), .A2(n5996), .ZN(n3576) );
  NAND2_X1 U4405 ( .A1(n3530), .A2(n5914), .ZN(n3574) );
  NAND2_X1 U4406 ( .A1(n3801), .A2(n5996), .ZN(n3573) );
  NAND3_X1 U4407 ( .A1(n3574), .A2(n3621), .A3(n3573), .ZN(n3575) );
  NAND2_X1 U4408 ( .A1(n3576), .A2(n3575), .ZN(n5482) );
  NAND2_X1 U4409 ( .A1(n3621), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3577) );
  OAI211_X1 U4410 ( .C1(n4448), .C2(EBX_REG_15__SCAN_IN), .A(n3612), .B(n3577), 
        .ZN(n3578) );
  OAI21_X1 U4411 ( .B1(n3608), .B2(EBX_REG_15__SCAN_IN), .A(n3578), .ZN(n5387)
         );
  INV_X1 U4412 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U4413 ( .A1(n3598), .A2(n5463), .ZN(n3581) );
  NAND2_X1 U4414 ( .A1(n3621), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3579) );
  OAI211_X1 U4415 ( .C1(n4448), .C2(EBX_REG_17__SCAN_IN), .A(n3612), .B(n3579), 
        .ZN(n3580) );
  AND2_X1 U4416 ( .A1(n3581), .A2(n3580), .ZN(n5459) );
  INV_X1 U4417 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U4418 ( .A1(n3618), .A2(n5986), .ZN(n3586) );
  NAND2_X1 U4419 ( .A1(n3612), .A2(n3582), .ZN(n3584) );
  NAND2_X1 U4420 ( .A1(n3801), .A2(n5986), .ZN(n3583) );
  NAND3_X1 U4421 ( .A1(n3584), .A2(n3621), .A3(n3583), .ZN(n3585) );
  NAND2_X1 U4422 ( .A1(n3586), .A2(n3585), .ZN(n5470) );
  NAND2_X1 U4423 ( .A1(n5459), .A2(n5470), .ZN(n3587) );
  MUX2_X1 U4424 ( .A(n3615), .B(n3612), .S(EBX_REG_19__SCAN_IN), .Z(n3589) );
  NAND2_X1 U4425 ( .A1(n4448), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3588) );
  NAND2_X1 U4426 ( .A1(n3589), .A2(n3588), .ZN(n5443) );
  NAND2_X1 U4427 ( .A1(n5461), .A2(n5443), .ZN(n5429) );
  OR2_X1 U4428 ( .A1(n3941), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3590)
         );
  INV_X1 U4429 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U4430 ( .A1(n3801), .A2(n5453), .ZN(n5440) );
  NAND2_X1 U4431 ( .A1(n3590), .A2(n5440), .ZN(n5441) );
  AND2_X1 U4432 ( .A1(n5441), .A2(n3621), .ZN(n3594) );
  OR2_X1 U4433 ( .A1(n3941), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3592)
         );
  INV_X1 U4434 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U4435 ( .A1(n3801), .A2(n5433), .ZN(n3591) );
  AND2_X1 U4436 ( .A1(n3592), .A2(n3591), .ZN(n5431) );
  OAI22_X1 U4437 ( .A1(n5431), .A2(n5441), .B1(n3621), .B2(n5433), .ZN(n3593)
         );
  MUX2_X1 U4438 ( .A(n3608), .B(n3621), .S(EBX_REG_21__SCAN_IN), .Z(n3595) );
  OAI21_X1 U4439 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n3941), .A(n3595), 
        .ZN(n5096) );
  MUX2_X1 U4440 ( .A(n3615), .B(n3612), .S(EBX_REG_22__SCAN_IN), .Z(n3597) );
  NAND2_X1 U4441 ( .A1(n4448), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3596) );
  NAND2_X1 U4442 ( .A1(n3597), .A2(n3596), .ZN(n5416) );
  INV_X1 U4443 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5115) );
  NAND2_X1 U4444 ( .A1(n3598), .A2(n5115), .ZN(n3601) );
  NAND2_X1 U4445 ( .A1(n3621), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3599) );
  OAI211_X1 U4446 ( .C1(n4448), .C2(EBX_REG_23__SCAN_IN), .A(n3612), .B(n3599), 
        .ZN(n3600) );
  AND2_X1 U4447 ( .A1(n3601), .A2(n3600), .ZN(n5112) );
  MUX2_X1 U4448 ( .A(n3615), .B(n3612), .S(EBX_REG_24__SCAN_IN), .Z(n3603) );
  NAND2_X1 U4449 ( .A1(n4448), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3602) );
  AND2_X1 U4450 ( .A1(n3603), .A2(n3602), .ZN(n5251) );
  OR2_X2 U4451 ( .A1(n5250), .A2(n5251), .ZN(n5369) );
  NAND2_X1 U4452 ( .A1(n3621), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3604) );
  OAI211_X1 U4453 ( .C1(n4448), .C2(EBX_REG_25__SCAN_IN), .A(n3612), .B(n3604), 
        .ZN(n3605) );
  OAI21_X1 U4454 ( .B1(n3608), .B2(EBX_REG_25__SCAN_IN), .A(n3605), .ZN(n5368)
         );
  NAND2_X1 U4455 ( .A1(n3612), .A2(n6567), .ZN(n3606) );
  OAI211_X1 U4456 ( .C1(EBX_REG_26__SCAN_IN), .C2(n4448), .A(n3606), .B(n3621), 
        .ZN(n3607) );
  OAI21_X1 U4457 ( .B1(n3615), .B2(EBX_REG_26__SCAN_IN), .A(n3607), .ZN(n4823)
         );
  MUX2_X1 U4458 ( .A(n3608), .B(n3621), .S(EBX_REG_27__SCAN_IN), .Z(n3609) );
  OAI21_X1 U4459 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n3941), .A(n3609), 
        .ZN(n3610) );
  INV_X1 U4460 ( .A(n3610), .ZN(n5334) );
  AND2_X2 U4461 ( .A1(n4822), .A2(n5334), .ZN(n5336) );
  INV_X1 U4462 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3611) );
  NAND2_X1 U4463 ( .A1(n3612), .A2(n3611), .ZN(n3613) );
  OAI211_X1 U4464 ( .C1(EBX_REG_28__SCAN_IN), .C2(n4448), .A(n3613), .B(n3621), 
        .ZN(n3614) );
  OAI21_X1 U4465 ( .B1(n3615), .B2(EBX_REG_28__SCAN_IN), .A(n3614), .ZN(n5322)
         );
  NAND2_X1 U4466 ( .A1(n5336), .A2(n5322), .ZN(n3619) );
  OR2_X1 U4467 ( .A1(n3941), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3617)
         );
  INV_X1 U4468 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5308) );
  NAND2_X1 U4469 ( .A1(n3801), .A2(n5308), .ZN(n3616) );
  NAND2_X1 U4470 ( .A1(n3617), .A2(n3616), .ZN(n5289) );
  NAND2_X1 U4471 ( .A1(n3618), .A2(n5308), .ZN(n5288) );
  OAI22_X1 U4472 ( .A1(n4801), .A2(n5439), .B1(n5288), .B2(n5324), .ZN(n5292)
         );
  AND2_X1 U4473 ( .A1(n3522), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3620)
         );
  AOI21_X1 U4474 ( .B1(n3941), .B2(EBX_REG_30__SCAN_IN), .A(n3620), .ZN(n4798)
         );
  AOI21_X1 U4475 ( .B1(n5292), .B2(n4798), .A(n4797), .ZN(n3623) );
  AOI22_X1 U4476 ( .A1(n3941), .A2(EBX_REG_31__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n3522), .ZN(n3622) );
  XNOR2_X1 U4477 ( .A(n3623), .B(n3622), .ZN(n5123) );
  NAND2_X1 U4478 ( .A1(n3625), .A2(n3624), .ZN(n3627) );
  NAND2_X1 U4479 ( .A1(n3626), .A2(n6537), .ZN(n6420) );
  NAND2_X1 U4480 ( .A1(n3627), .A2(n6420), .ZN(n3628) );
  AOI22_X1 U4481 ( .A1(n3129), .A2(n5439), .B1(n3973), .B2(n5106), .ZN(n3632)
         );
  NOR2_X1 U4482 ( .A1(n3675), .A2(n3973), .ZN(n3870) );
  OAI21_X1 U4483 ( .B1(n3870), .B2(n3941), .A(n3629), .ZN(n3630) );
  NAND3_X1 U4484 ( .A1(n3632), .A2(n3631), .A3(n3630), .ZN(n3633) );
  OR2_X1 U4485 ( .A1(n3634), .A2(n3633), .ZN(n3822) );
  INV_X1 U4486 ( .A(n3822), .ZN(n3850) );
  AND3_X1 U4487 ( .A1(n3636), .A2(n3635), .A3(n3638), .ZN(n3637) );
  NAND2_X1 U4488 ( .A1(n4884), .A2(n3637), .ZN(n3994) );
  INV_X1 U4489 ( .A(n3848), .ZN(n3639) );
  NAND2_X1 U4490 ( .A1(n3639), .A2(n3638), .ZN(n3640) );
  OAI211_X1 U4491 ( .C1(n3846), .C2(n3641), .A(n3994), .B(n3640), .ZN(n3642)
         );
  INV_X1 U4492 ( .A(n3642), .ZN(n3643) );
  NAND2_X1 U4493 ( .A1(n3850), .A2(n3643), .ZN(n3644) );
  INV_X1 U4494 ( .A(n3659), .ZN(n3648) );
  NOR2_X1 U4495 ( .A1(n3822), .A2(n3645), .ZN(n3852) );
  NAND2_X1 U4496 ( .A1(n3852), .A2(n3649), .ZN(n6283) );
  NAND2_X1 U4497 ( .A1(n3648), .A2(n6283), .ZN(n5916) );
  AND2_X1 U4498 ( .A1(n3674), .A2(n3930), .ZN(n3996) );
  NAND2_X1 U4499 ( .A1(n3649), .A2(n3996), .ZN(n6308) );
  INV_X1 U4500 ( .A(n6308), .ZN(n3798) );
  AND2_X1 U4501 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4825) );
  INV_X1 U4502 ( .A(n6236), .ZN(n5899) );
  NAND2_X1 U4503 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U4504 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6243) );
  NOR2_X1 U4505 ( .A1(n6242), .A2(n6243), .ZN(n3647) );
  INV_X1 U4506 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3896) );
  INV_X1 U4507 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6309) );
  INV_X1 U4508 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6292) );
  OAI21_X1 U4509 ( .B1(n3896), .B2(n6309), .A(n6292), .ZN(n6285) );
  INV_X1 U4510 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6653) );
  NOR4_X1 U4511 ( .A1(n6653), .A2(n3333), .A3(n3355), .A4(n3378), .ZN(n4239)
         );
  AND2_X1 U4512 ( .A1(n6285), .A2(n4239), .ZN(n4234) );
  AND2_X1 U4513 ( .A1(n3647), .A2(n4234), .ZN(n3666) );
  NAND2_X1 U4514 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5924) );
  NOR2_X1 U4515 ( .A1(n3646), .A2(n5924), .ZN(n5918) );
  NAND2_X1 U4516 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5918), .ZN(n5898) );
  NAND2_X1 U4517 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5903) );
  NOR2_X1 U4518 ( .A1(n5898), .A2(n5903), .ZN(n3654) );
  NOR2_X1 U4519 ( .A1(n6292), .A2(n3896), .ZN(n4160) );
  NAND2_X1 U4520 ( .A1(n4160), .A2(n4239), .ZN(n4233) );
  INV_X1 U4521 ( .A(n3647), .ZN(n4715) );
  OR2_X1 U4522 ( .A1(n4233), .A2(n4715), .ZN(n3665) );
  NAND2_X1 U4523 ( .A1(n3648), .A2(n6308), .ZN(n4232) );
  INV_X1 U4524 ( .A(n3654), .ZN(n3652) );
  NAND2_X1 U4525 ( .A1(n3659), .A2(n6309), .ZN(n3651) );
  INV_X1 U4526 ( .A(n3649), .ZN(n3650) );
  OR2_X1 U4527 ( .A1(n4216), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U4528 ( .A1(n3650), .A2(n6238), .ZN(n6307) );
  NAND2_X1 U4529 ( .A1(n3651), .A2(n6307), .ZN(n4231) );
  AOI221_X1 U4530 ( .B1(n3665), .B2(n4232), .C1(n3652), .C2(n4232), .A(n4231), 
        .ZN(n3653) );
  OAI221_X1 U4531 ( .B1(n6283), .B2(n3666), .C1(n6283), .C2(n3654), .A(n3653), 
        .ZN(n5713) );
  INV_X1 U4532 ( .A(n3667), .ZN(n3655) );
  NAND2_X1 U4533 ( .A1(n3655), .A2(n5694), .ZN(n3656) );
  AND2_X1 U4534 ( .A1(n6236), .A2(n3656), .ZN(n3657) );
  NOR2_X1 U4535 ( .A1(n5713), .A2(n3657), .ZN(n5686) );
  INV_X1 U4536 ( .A(n5676), .ZN(n3668) );
  NAND2_X1 U4537 ( .A1(n6236), .A2(n3668), .ZN(n3658) );
  AND2_X1 U4538 ( .A1(n5686), .A2(n3658), .ZN(n5665) );
  NAND2_X1 U4539 ( .A1(n3659), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3664)
         );
  NAND2_X1 U4540 ( .A1(n3664), .A2(n6308), .ZN(n6291) );
  INV_X1 U4541 ( .A(n6283), .ZN(n6264) );
  INV_X1 U4542 ( .A(n3660), .ZN(n3669) );
  OAI21_X1 U4543 ( .B1(n6291), .B2(n6264), .A(n3669), .ZN(n3661) );
  OAI21_X1 U4544 ( .B1(n4825), .B2(n5899), .A(n5660), .ZN(n5654) );
  AOI211_X1 U4545 ( .C1(n5643), .C2(n6236), .A(n5632), .B(n5654), .ZN(n5631)
         );
  INV_X1 U4546 ( .A(n5660), .ZN(n4829) );
  NOR2_X1 U4547 ( .A1(n4829), .A2(n6236), .ZN(n4805) );
  INV_X1 U4548 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n3897) );
  AOI211_X1 U4549 ( .C1(n5631), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n4805), .B(n3897), .ZN(n3663) );
  NAND2_X1 U4550 ( .A1(n2997), .A2(REIP_REG_31__SCAN_IN), .ZN(n5264) );
  INV_X1 U4551 ( .A(n5264), .ZN(n3662) );
  AOI21_X1 U4552 ( .B1(n5123), .B2(n6288), .A(n3006), .ZN(n3671) );
  NOR2_X1 U4553 ( .A1(n6308), .A2(n3665), .ZN(n4717) );
  INV_X1 U4554 ( .A(n4717), .ZN(n5932) );
  OAI21_X1 U4555 ( .B1(n3665), .B2(n3664), .A(n6283), .ZN(n4716) );
  NAND2_X1 U4556 ( .A1(n4716), .A2(n3666), .ZN(n5915) );
  NAND3_X1 U4557 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5911), .ZN(n5891) );
  NOR2_X1 U4558 ( .A1(n5891), .A2(n3667), .ZN(n5705) );
  NAND2_X1 U4559 ( .A1(n5705), .A2(n5694), .ZN(n5682) );
  NOR2_X1 U4560 ( .A1(n5668), .A2(n3669), .ZN(n5662) );
  NAND2_X1 U4561 ( .A1(n5662), .A2(n4825), .ZN(n5651) );
  NOR3_X1 U4562 ( .A1(n5651), .A2(n5643), .A3(n5632), .ZN(n4809) );
  NAND3_X1 U4563 ( .A1(n4809), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n3897), .ZN(n3670) );
  AND2_X1 U4564 ( .A1(n3671), .A2(n3670), .ZN(n3672) );
  OAI21_X1 U4565 ( .B1(n5268), .B2(n6269), .A(n3672), .ZN(U2987) );
  INV_X1 U4566 ( .A(n3673), .ZN(n3687) );
  AND2_X1 U4567 ( .A1(n3674), .A2(n3687), .ZN(n3679) );
  NAND2_X1 U4568 ( .A1(n3679), .A2(n6435), .ZN(n5309) );
  NAND3_X1 U4569 ( .A1(n3879), .A2(n6435), .A3(n4213), .ZN(n5310) );
  NAND2_X1 U4570 ( .A1(n5309), .A2(n5310), .ZN(n6533) );
  INV_X1 U4571 ( .A(n6533), .ZN(n3678) );
  INV_X1 U4572 ( .A(n3675), .ZN(n4581) );
  OR2_X1 U4573 ( .A1(n6537), .A2(n4581), .ZN(n3680) );
  NOR2_X1 U4574 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n4619) );
  NAND2_X1 U4575 ( .A1(n5723), .A2(n4812), .ZN(n5944) );
  INV_X1 U4576 ( .A(n5944), .ZN(n3676) );
  OAI21_X1 U4577 ( .B1(n3676), .B2(READREQUEST_REG_SCAN_IN), .A(n3678), .ZN(
        n3677) );
  OAI21_X1 U4578 ( .B1(n3678), .B2(n3680), .A(n3677), .ZN(U3474) );
  OAI22_X1 U4579 ( .A1(n3679), .A2(n3879), .B1(n4582), .B2(n4213), .ZN(n5942)
         );
  AOI21_X1 U4580 ( .B1(n3680), .B2(n6539), .A(READY_N), .ZN(n3681) );
  NOR2_X1 U4581 ( .A1(n5942), .A2(n3681), .ZN(n6408) );
  INV_X1 U4582 ( .A(n6435), .ZN(n6432) );
  OR2_X1 U4583 ( .A1(n6408), .A2(n6432), .ZN(n3689) );
  INV_X1 U4584 ( .A(n3689), .ZN(n5949) );
  INV_X1 U4585 ( .A(MORE_REG_SCAN_IN), .ZN(n3691) );
  INV_X1 U4586 ( .A(n3879), .ZN(n3682) );
  NAND2_X1 U4587 ( .A1(n6410), .A2(n3682), .ZN(n3684) );
  INV_X1 U4588 ( .A(n4213), .ZN(n3683) );
  OAI21_X1 U4589 ( .B1(n3851), .B2(n3684), .A(n3683), .ZN(n3685) );
  OAI21_X1 U4590 ( .B1(n3687), .B2(n3686), .A(n3685), .ZN(n3688) );
  AOI21_X1 U4591 ( .B1(n3852), .B2(n4213), .A(n3688), .ZN(n6411) );
  OR2_X1 U4592 ( .A1(n3689), .A2(n6411), .ZN(n3690) );
  OAI21_X1 U4593 ( .B1(n5949), .B2(n3691), .A(n3690), .ZN(U3471) );
  NOR2_X1 U4594 ( .A1(n6420), .A2(n6432), .ZN(n3692) );
  NAND2_X1 U4595 ( .A1(n3692), .A2(n4213), .ZN(n6180) );
  INV_X2 U4596 ( .A(n6180), .ZN(n6174) );
  NOR2_X1 U4597 ( .A1(n5310), .A2(READY_N), .ZN(n3693) );
  NOR2_X1 U4598 ( .A1(n6174), .A2(n3693), .ZN(n6178) );
  AOI22_X1 U4599 ( .A1(n6178), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n6174), .ZN(n3695) );
  NAND2_X1 U4600 ( .A1(n3693), .A2(n3930), .ZN(n3773) );
  INV_X1 U4601 ( .A(DATAI_8_), .ZN(n3694) );
  OR2_X1 U4602 ( .A1(n3773), .A2(n3694), .ZN(n3834) );
  NAND2_X1 U4603 ( .A1(n3695), .A2(n3834), .ZN(U2947) );
  AOI22_X1 U4604 ( .A1(n6178), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6174), .ZN(n3696) );
  INV_X1 U4605 ( .A(DATAI_7_), .ZN(n3956) );
  OR2_X1 U4606 ( .A1(n3773), .A2(n3956), .ZN(n3827) );
  NAND2_X1 U4607 ( .A1(n3696), .A2(n3827), .ZN(U2946) );
  AOI22_X1 U4608 ( .A1(n6178), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n6174), .ZN(n3697) );
  INV_X1 U4609 ( .A(n3773), .ZN(n6177) );
  NAND2_X1 U4610 ( .A1(n6177), .A2(DATAI_13_), .ZN(n3730) );
  NAND2_X1 U4611 ( .A1(n3697), .A2(n3730), .ZN(U2952) );
  INV_X1 U4612 ( .A(EAX_REG_17__SCAN_IN), .ZN(n3701) );
  INV_X1 U4613 ( .A(n3996), .ZN(n3906) );
  NAND2_X1 U4614 ( .A1(n3906), .A2(n6420), .ZN(n3699) );
  INV_X1 U4615 ( .A(n6539), .ZN(n4444) );
  AND3_X1 U4616 ( .A1(n4213), .A2(n4444), .A3(n6435), .ZN(n3698) );
  NAND2_X1 U4617 ( .A1(n6145), .A2(n4452), .ZN(n6745) );
  INV_X2 U4618 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6532) );
  NOR2_X1 U4619 ( .A1(n4812), .A2(n6532), .ZN(n4028) );
  NAND2_X1 U4620 ( .A1(n6540), .A2(n4028), .ZN(n6142) );
  INV_X2 U4621 ( .A(n6750), .ZN(n6156) );
  AOI22_X1 U4622 ( .A1(n6746), .A2(UWORD_REG_1__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n3700) );
  OAI21_X1 U4623 ( .B1(n3701), .B2(n6745), .A(n3700), .ZN(U2906) );
  INV_X1 U4624 ( .A(EAX_REG_18__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4625 ( .A1(n6746), .A2(UWORD_REG_2__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n3702) );
  OAI21_X1 U4626 ( .B1(n3703), .B2(n6745), .A(n3702), .ZN(U2905) );
  INV_X1 U4627 ( .A(EAX_REG_23__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4628 ( .A1(n6746), .A2(UWORD_REG_7__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n3704) );
  OAI21_X1 U4629 ( .B1(n3705), .B2(n6745), .A(n3704), .ZN(U2900) );
  INV_X1 U4630 ( .A(EAX_REG_24__SCAN_IN), .ZN(n3707) );
  AOI22_X1 U4631 ( .A1(n6746), .A2(UWORD_REG_8__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n3706) );
  OAI21_X1 U4632 ( .B1(n3707), .B2(n6745), .A(n3706), .ZN(U2899) );
  INV_X1 U4633 ( .A(EAX_REG_19__SCAN_IN), .ZN(n3709) );
  AOI22_X1 U4634 ( .A1(n6746), .A2(UWORD_REG_3__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n3708) );
  OAI21_X1 U4635 ( .B1(n3709), .B2(n6745), .A(n3708), .ZN(U2904) );
  INV_X1 U4636 ( .A(EAX_REG_22__SCAN_IN), .ZN(n3711) );
  AOI22_X1 U4637 ( .A1(n6746), .A2(UWORD_REG_6__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n3710) );
  OAI21_X1 U4638 ( .B1(n3711), .B2(n6745), .A(n3710), .ZN(U2901) );
  INV_X1 U4639 ( .A(EAX_REG_25__SCAN_IN), .ZN(n3713) );
  AOI22_X1 U4640 ( .A1(n6746), .A2(UWORD_REG_9__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n3712) );
  OAI21_X1 U4641 ( .B1(n3713), .B2(n6745), .A(n3712), .ZN(U2898) );
  INV_X1 U4642 ( .A(EAX_REG_16__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4643 ( .A1(n6746), .A2(UWORD_REG_0__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n3714) );
  OAI21_X1 U4644 ( .B1(n3715), .B2(n6745), .A(n3714), .ZN(U2907) );
  INV_X1 U4645 ( .A(EAX_REG_27__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4646 ( .A1(n6746), .A2(UWORD_REG_11__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n3716) );
  OAI21_X1 U4647 ( .B1(n3717), .B2(n6745), .A(n3716), .ZN(U2896) );
  INV_X1 U4648 ( .A(EAX_REG_30__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4649 ( .A1(n6746), .A2(UWORD_REG_14__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n3718) );
  OAI21_X1 U4650 ( .B1(n3719), .B2(n6745), .A(n3718), .ZN(U2893) );
  INV_X1 U4651 ( .A(EAX_REG_28__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4652 ( .A1(n6746), .A2(UWORD_REG_12__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n3720) );
  OAI21_X1 U4653 ( .B1(n3721), .B2(n6745), .A(n3720), .ZN(U2895) );
  INV_X1 U4654 ( .A(EAX_REG_29__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4655 ( .A1(n6746), .A2(UWORD_REG_13__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n3722) );
  OAI21_X1 U4656 ( .B1(n3723), .B2(n6745), .A(n3722), .ZN(U2894) );
  INV_X1 U4657 ( .A(EAX_REG_20__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4658 ( .A1(n6746), .A2(UWORD_REG_4__SCAN_IN), .B1(
        DATAO_REG_20__SCAN_IN), .B2(n6156), .ZN(n3724) );
  OAI21_X1 U4659 ( .B1(n3725), .B2(n6745), .A(n3724), .ZN(U2903) );
  AOI22_X1 U4660 ( .A1(n6164), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6174), .ZN(n3726) );
  NAND2_X1 U4661 ( .A1(n6177), .A2(DATAI_2_), .ZN(n3836) );
  NAND2_X1 U4662 ( .A1(n3726), .A2(n3836), .ZN(U2941) );
  AOI22_X1 U4663 ( .A1(n6164), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6174), .ZN(n3727) );
  INV_X1 U4664 ( .A(DATAI_3_), .ZN(n3934) );
  OR2_X1 U4665 ( .A1(n3773), .A2(n3934), .ZN(n3831) );
  NAND2_X1 U4666 ( .A1(n3727), .A2(n3831), .ZN(U2942) );
  AOI22_X1 U4667 ( .A1(n6164), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6174), .ZN(n3728) );
  NAND2_X1 U4668 ( .A1(n6177), .A2(DATAI_0_), .ZN(n3829) );
  NAND2_X1 U4669 ( .A1(n3728), .A2(n3829), .ZN(U2939) );
  AOI22_X1 U4670 ( .A1(n6164), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6174), .ZN(n3729) );
  INV_X1 U4671 ( .A(DATAI_1_), .ZN(n3929) );
  OR2_X1 U4672 ( .A1(n3773), .A2(n3929), .ZN(n3838) );
  NAND2_X1 U4673 ( .A1(n3729), .A2(n3838), .ZN(U2940) );
  AOI22_X1 U4674 ( .A1(n6164), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n6174), .ZN(n3731) );
  NAND2_X1 U4675 ( .A1(n3731), .A2(n3730), .ZN(U2937) );
  AOI22_X1 U4676 ( .A1(n6164), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6174), .ZN(n3732) );
  INV_X1 U4677 ( .A(DATAI_5_), .ZN(n3977) );
  OR2_X1 U4678 ( .A1(n3773), .A2(n3977), .ZN(n3844) );
  NAND2_X1 U4679 ( .A1(n3732), .A2(n3844), .ZN(U2944) );
  NOR2_X2 U4680 ( .A1(n3921), .A2(n6532), .ZN(n4998) );
  AND2_X1 U4681 ( .A1(n6532), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5219) );
  AOI21_X1 U4682 ( .B1(n4038), .B2(n4998), .A(n5219), .ZN(n3789) );
  NAND2_X1 U4683 ( .A1(n3733), .A2(n4998), .ZN(n3737) );
  NOR2_X1 U4684 ( .A1(n5107), .A2(n6532), .ZN(n5158) );
  AOI22_X1 U4685 ( .A1(n5158), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6532), .ZN(n3735) );
  NOR2_X1 U4686 ( .A1(n5106), .A2(n6532), .ZN(n3755) );
  NAND2_X1 U4687 ( .A1(n3755), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3734) );
  AND2_X1 U4688 ( .A1(n3735), .A2(n3734), .ZN(n3736) );
  NAND2_X1 U4689 ( .A1(n3737), .A2(n3736), .ZN(n3886) );
  NAND2_X1 U4690 ( .A1(n4398), .A2(n3738), .ZN(n3784) );
  INV_X1 U4691 ( .A(n5306), .ZN(n4131) );
  NAND2_X1 U4692 ( .A1(n4131), .A2(n4998), .ZN(n3743) );
  AOI22_X1 U4693 ( .A1(n5158), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6532), .ZN(n3741) );
  NAND2_X1 U4694 ( .A1(n3755), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3740) );
  AND2_X1 U4695 ( .A1(n3741), .A2(n3740), .ZN(n3742) );
  NAND2_X1 U4696 ( .A1(n3743), .A2(n3742), .ZN(n3786) );
  AND2_X1 U4697 ( .A1(n3786), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3744) );
  NAND2_X1 U4698 ( .A1(n3784), .A2(n3744), .ZN(n3785) );
  INV_X1 U4699 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6538) );
  NAND2_X1 U4700 ( .A1(n6532), .A2(n6538), .ZN(n5210) );
  OR2_X1 U4701 ( .A1(n3786), .A2(n5210), .ZN(n3745) );
  NAND2_X1 U4702 ( .A1(n3785), .A2(n3745), .ZN(n3885) );
  NAND2_X1 U4703 ( .A1(n3886), .A2(n3885), .ZN(n3752) );
  NAND2_X1 U4704 ( .A1(n3755), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3750) );
  INV_X1 U4705 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3747) );
  INV_X1 U4706 ( .A(n5219), .ZN(n4768) );
  INV_X2 U4707 ( .A(n5210), .ZN(n5216) );
  OAI21_X1 U4708 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3757), .ZN(n6217) );
  NAND2_X1 U4709 ( .A1(n5216), .A2(n6217), .ZN(n3746) );
  OAI21_X1 U4710 ( .B1(n3747), .B2(n4768), .A(n3746), .ZN(n3748) );
  AOI21_X1 U4711 ( .B1(n5220), .B2(EAX_REG_2__SCAN_IN), .A(n3748), .ZN(n3749)
         );
  AND2_X1 U4712 ( .A1(n3750), .A2(n3749), .ZN(n3788) );
  OR2_X2 U4713 ( .A1(n3752), .A2(n3788), .ZN(n3751) );
  NAND2_X1 U4714 ( .A1(n3789), .A2(n3751), .ZN(n3754) );
  NAND2_X1 U4715 ( .A1(n3752), .A2(n3788), .ZN(n3753) );
  NAND2_X1 U4716 ( .A1(n3754), .A2(n3753), .ZN(n3791) );
  INV_X1 U4717 ( .A(n3755), .ZN(n3811) );
  INV_X1 U4718 ( .A(n3757), .ZN(n3759) );
  INV_X1 U4719 ( .A(n3812), .ZN(n3758) );
  OAI21_X1 U4720 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3759), .A(n3758), 
        .ZN(n4592) );
  AOI22_X1 U4721 ( .A1(n5216), .A2(n4592), .B1(n5219), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3761) );
  NAND2_X1 U4722 ( .A1(n5220), .A2(EAX_REG_3__SCAN_IN), .ZN(n3760) );
  OAI211_X1 U4723 ( .C1(n3811), .C2(n3882), .A(n3761), .B(n3760), .ZN(n3762)
         );
  AOI21_X1 U4724 ( .B1(n4039), .B2(n4998), .A(n3762), .ZN(n3763) );
  NOR2_X2 U4725 ( .A1(n3791), .A2(n3763), .ZN(n3817) );
  AND2_X1 U4726 ( .A1(n3791), .A2(n3763), .ZN(n3764) );
  OR2_X1 U4727 ( .A1(n3817), .A2(n3764), .ZN(n4215) );
  INV_X1 U4728 ( .A(n3765), .ZN(n3769) );
  NOR2_X1 U4729 ( .A1(n5107), .A2(n3766), .ZN(n3768) );
  NOR2_X1 U4730 ( .A1(n3973), .A2(n3935), .ZN(n3767) );
  NAND4_X1 U4731 ( .A1(n3770), .A2(n3769), .A3(n3768), .A4(n3767), .ZN(n3819)
         );
  OR2_X1 U4732 ( .A1(n3819), .A2(n3771), .ZN(n3772) );
  INV_X1 U4733 ( .A(n3774), .ZN(n3775) );
  OR2_X1 U4734 ( .A1(n5934), .A2(n3775), .ZN(n3777) );
  NAND2_X1 U4735 ( .A1(n3851), .A2(n4213), .ZN(n3776) );
  NAND2_X1 U4736 ( .A1(n3777), .A2(n3776), .ZN(n3875) );
  NAND2_X1 U4737 ( .A1(n3875), .A2(n6435), .ZN(n3778) );
  NAND2_X1 U4738 ( .A1(n3002), .A2(n5107), .ZN(n3781) );
  NAND2_X2 U4739 ( .A1(n6131), .A2(n3781), .ZN(n5863) );
  INV_X1 U4740 ( .A(n3781), .ZN(n3782) );
  AOI22_X1 U4741 ( .A1(n5511), .A2(DATAI_3_), .B1(n6122), .B2(
        EAX_REG_3__SCAN_IN), .ZN(n3783) );
  OAI21_X1 U4742 ( .B1(n4215), .B2(n5863), .A(n3783), .ZN(U2888) );
  AND2_X1 U4743 ( .A1(n3784), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3787) );
  OAI21_X1 U4744 ( .B1(n3787), .B2(n3786), .A(n3785), .ZN(n5298) );
  INV_X1 U4745 ( .A(DATAI_0_), .ZN(n3925) );
  INV_X1 U4746 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6159) );
  OAI222_X1 U4747 ( .A1(n5298), .A2(n5863), .B1(n6126), .B2(n3925), .C1(n6131), 
        .C2(n6159), .ZN(U2891) );
  NAND3_X1 U4748 ( .A1(n3789), .A2(n3788), .A3(n3752), .ZN(n3790) );
  AND2_X1 U4749 ( .A1(n3791), .A2(n3790), .ZN(n6214) );
  INV_X1 U4750 ( .A(n6214), .ZN(n3891) );
  INV_X1 U4751 ( .A(DATAI_2_), .ZN(n3972) );
  INV_X1 U4752 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6153) );
  OAI222_X1 U4753 ( .A1(n3891), .A2(n5863), .B1(n6126), .B2(n3972), .C1(n6131), 
        .C2(n6153), .ZN(U2889) );
  INV_X1 U4754 ( .A(n6269), .ZN(n6298) );
  NAND2_X1 U4755 ( .A1(n3793), .A2(n3792), .ZN(n3794) );
  OR2_X1 U4756 ( .A1(n3795), .A2(n3794), .ZN(n3797) );
  NAND2_X1 U4757 ( .A1(n3795), .A2(n3794), .ZN(n3796) );
  AND2_X1 U4758 ( .A1(n3797), .A2(n3796), .ZN(n6222) );
  AOI21_X1 U4759 ( .B1(n5916), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n3798), 
        .ZN(n3803) );
  OAI21_X1 U4760 ( .B1(n3799), .B2(n3801), .A(n3800), .ZN(n3888) );
  AOI22_X1 U4761 ( .A1(n6288), .A2(n3888), .B1(n2997), .B2(REIP_REG_1__SCAN_IN), .ZN(n3802) );
  OAI21_X1 U4762 ( .B1(n3803), .B2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n3802), 
        .ZN(n3805) );
  NAND2_X1 U4763 ( .A1(n5916), .A2(n6309), .ZN(n6301) );
  AOI21_X1 U4764 ( .B1(n6307), .B2(n6301), .A(n3896), .ZN(n3804) );
  AOI211_X1 U4765 ( .C1(n6298), .C2(n6222), .A(n3805), .B(n3804), .ZN(n3806)
         );
  INV_X1 U4766 ( .A(n3806), .ZN(U3017) );
  INV_X1 U4767 ( .A(n4998), .ZN(n3807) );
  NAND2_X1 U4768 ( .A1(n6532), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3810)
         );
  NAND2_X1 U4769 ( .A1(n5220), .A2(EAX_REG_4__SCAN_IN), .ZN(n3809) );
  OAI211_X1 U4770 ( .C1(n3811), .C2(n5939), .A(n3810), .B(n3809), .ZN(n3814)
         );
  OAI21_X1 U4771 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3812), .A(n4051), 
        .ZN(n6078) );
  AND2_X1 U4772 ( .A1(n5216), .A2(n6078), .ZN(n3813) );
  AOI21_X1 U4773 ( .B1(n3814), .B2(n5210), .A(n3813), .ZN(n3815) );
  NAND2_X1 U4774 ( .A1(n3817), .A2(n3818), .ZN(n4060) );
  OAI21_X1 U4775 ( .B1(n3817), .B2(n3818), .A(n4060), .ZN(n4225) );
  NAND2_X1 U4776 ( .A1(n3871), .A2(n6435), .ZN(n3821) );
  OR2_X1 U4777 ( .A1(n3819), .A2(n4448), .ZN(n3820) );
  INV_X1 U4778 ( .A(n4064), .ZN(n3824) );
  XNOR2_X1 U4779 ( .A(n3823), .B(n3824), .ZN(n6266) );
  INV_X1 U4780 ( .A(n5107), .ZN(n5489) );
  INV_X1 U4781 ( .A(n6111), .ZN(n5399) );
  AOI22_X1 U4782 ( .A1(n6266), .A2(n6107), .B1(n5399), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n3825) );
  OAI21_X1 U4783 ( .B1(n4225), .B2(n5466), .A(n3825), .ZN(U2855) );
  AOI22_X1 U4784 ( .A1(n6178), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6174), .ZN(n3826) );
  NAND2_X1 U4785 ( .A1(n6177), .A2(DATAI_4_), .ZN(n3840) );
  NAND2_X1 U4786 ( .A1(n3826), .A2(n3840), .ZN(U2928) );
  AOI22_X1 U4787 ( .A1(n6178), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6174), .ZN(n3828) );
  NAND2_X1 U4788 ( .A1(n3828), .A2(n3827), .ZN(U2931) );
  AOI22_X1 U4789 ( .A1(n6164), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n6174), .ZN(n3830) );
  NAND2_X1 U4790 ( .A1(n3830), .A2(n3829), .ZN(U2924) );
  AOI22_X1 U4791 ( .A1(n6164), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6174), .ZN(n3832) );
  NAND2_X1 U4792 ( .A1(n3832), .A2(n3831), .ZN(U2927) );
  AOI22_X1 U4793 ( .A1(n6164), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6174), .ZN(n3833) );
  NAND2_X1 U4794 ( .A1(n6177), .A2(DATAI_6_), .ZN(n3842) );
  NAND2_X1 U4795 ( .A1(n3833), .A2(n3842), .ZN(U2945) );
  AOI22_X1 U4796 ( .A1(n6164), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n6174), .ZN(n3835) );
  NAND2_X1 U4797 ( .A1(n3835), .A2(n3834), .ZN(U2932) );
  AOI22_X1 U4798 ( .A1(n6164), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6174), .ZN(n3837) );
  NAND2_X1 U4799 ( .A1(n3837), .A2(n3836), .ZN(U2926) );
  AOI22_X1 U4800 ( .A1(n6164), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n6174), .ZN(n3839) );
  NAND2_X1 U4801 ( .A1(n3839), .A2(n3838), .ZN(U2925) );
  AOI22_X1 U4802 ( .A1(n6164), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6174), .ZN(n3841) );
  NAND2_X1 U4803 ( .A1(n3841), .A2(n3840), .ZN(U2943) );
  AOI22_X1 U4804 ( .A1(n6164), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6174), .ZN(n3843) );
  NAND2_X1 U4805 ( .A1(n3843), .A2(n3842), .ZN(U2930) );
  AOI22_X1 U4806 ( .A1(n6164), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6174), .ZN(n3845) );
  NAND2_X1 U4807 ( .A1(n3845), .A2(n3844), .ZN(U2929) );
  AND4_X1 U4808 ( .A1(n5934), .A2(n3848), .A3(n3847), .A4(n3846), .ZN(n3849)
         );
  NAND2_X1 U4809 ( .A1(n3850), .A2(n3849), .ZN(n4001) );
  NAND2_X1 U4810 ( .A1(n4681), .A2(n4001), .ZN(n3867) );
  OR2_X1 U4811 ( .A1(n3852), .A2(n3851), .ZN(n3989) );
  NOR2_X1 U4812 ( .A1(n3993), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3855)
         );
  AND2_X1 U4813 ( .A1(n3989), .A2(n3855), .ZN(n4000) );
  INV_X1 U4814 ( .A(n4000), .ZN(n3854) );
  NAND2_X1 U4815 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3857) );
  NAND2_X1 U4816 ( .A1(n3996), .A2(n3857), .ZN(n3853) );
  NAND2_X1 U4817 ( .A1(n3854), .A2(n3853), .ZN(n3862) );
  INV_X1 U4818 ( .A(n3855), .ZN(n3856) );
  NAND2_X1 U4819 ( .A1(n3989), .A2(n3856), .ZN(n3860) );
  INV_X1 U4820 ( .A(n3857), .ZN(n3858) );
  NAND2_X1 U4821 ( .A1(n3996), .A2(n3858), .ZN(n3859) );
  NAND2_X1 U4822 ( .A1(n3860), .A2(n3859), .ZN(n3861) );
  MUX2_X1 U4823 ( .A(n3862), .B(n3861), .S(n3882), .Z(n3865) );
  AOI21_X1 U4824 ( .B1(n3993), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3882), 
        .ZN(n3863) );
  NOR2_X1 U4825 ( .A1(n5195), .A2(n3863), .ZN(n3868) );
  NOR2_X1 U4826 ( .A1(n3994), .A2(n3868), .ZN(n3864) );
  NOR2_X1 U4827 ( .A1(n3865), .A2(n3864), .ZN(n3866) );
  NAND2_X1 U4828 ( .A1(n3867), .A2(n3866), .ZN(n3988) );
  INV_X1 U4829 ( .A(n6434), .ZN(n5936) );
  NOR2_X1 U4830 ( .A1(n6423), .A2(n3868), .ZN(n3869) );
  AOI21_X1 U4831 ( .B1(n3988), .B2(n5936), .A(n3869), .ZN(n3883) );
  NOR2_X1 U4832 ( .A1(n3871), .A2(n3870), .ZN(n3872) );
  NAND2_X1 U4833 ( .A1(n3873), .A2(n3872), .ZN(n3874) );
  NOR2_X1 U4834 ( .A1(n3875), .A2(n3874), .ZN(n3881) );
  NAND2_X1 U4835 ( .A1(n3996), .A2(n6455), .ZN(n3877) );
  NAND2_X1 U4836 ( .A1(n3877), .A2(n3876), .ZN(n3878) );
  OAI211_X1 U4837 ( .C1(n3879), .C2(n4444), .A(n3878), .B(n4213), .ZN(n3880)
         );
  NAND2_X1 U4838 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4028), .ZN(n6440) );
  INV_X1 U4839 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5948) );
  OAI22_X1 U4840 ( .A1(n6391), .A2(n6432), .B1(n6440), .B2(n5948), .ZN(n5935)
         );
  AOI21_X1 U4841 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6540), .A(n5935), .ZN(
        n4819) );
  MUX2_X1 U4842 ( .A(n3883), .B(n3882), .S(n4819), .Z(n3884) );
  INV_X1 U4843 ( .A(n3884), .ZN(U3456) );
  OR2_X1 U4844 ( .A1(n3886), .A2(n3885), .ZN(n3887) );
  AND2_X1 U4845 ( .A1(n3752), .A2(n3887), .ZN(n6220) );
  INV_X1 U4846 ( .A(n6220), .ZN(n3987) );
  AOI22_X1 U4847 ( .A1(n6107), .A2(n3888), .B1(n5399), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n3889) );
  OAI21_X1 U4848 ( .B1(n3987), .B2(n5466), .A(n3889), .ZN(U2858) );
  XNOR2_X1 U4849 ( .A(n4587), .B(n4589), .ZN(n6287) );
  AOI22_X1 U4850 ( .A1(n6107), .A2(n6287), .B1(n5399), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n3890) );
  OAI21_X1 U4851 ( .B1(n3891), .B2(n5466), .A(n3890), .ZN(U2857) );
  INV_X1 U4852 ( .A(DATAI_4_), .ZN(n3945) );
  INV_X1 U4853 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6149) );
  OAI222_X1 U4854 ( .A1(n4225), .A2(n5863), .B1(n6126), .B2(n3945), .C1(n6149), 
        .C2(n6131), .ZN(U2887) );
  INV_X1 U4855 ( .A(n4097), .ZN(n4609) );
  INV_X1 U4856 ( .A(n4001), .ZN(n3903) );
  AND2_X1 U4857 ( .A1(n3996), .A2(n3892), .ZN(n3991) );
  INV_X1 U4858 ( .A(n3991), .ZN(n3895) );
  OAI21_X1 U4859 ( .B1(n3898), .B2(n3893), .A(n4884), .ZN(n3894) );
  OAI211_X1 U4860 ( .C1(n4609), .C2(n3903), .A(n3895), .B(n3894), .ZN(n6393)
         );
  AOI22_X1 U4861 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n3897), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n3896), .ZN(n4811) );
  NOR2_X1 U4862 ( .A1(n4812), .A2(n6309), .ZN(n3899) );
  INV_X1 U4863 ( .A(n6423), .ZN(n4817) );
  AOI222_X1 U4864 ( .A1(n6393), .A2(n5936), .B1(n4811), .B2(n3899), .C1(n3898), 
        .C2(n4817), .ZN(n3901) );
  INV_X1 U4865 ( .A(n4819), .ZN(n5940) );
  OAI21_X1 U4866 ( .B1(n6423), .B2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(n5940), 
        .ZN(n3904) );
  NAND2_X1 U4867 ( .A1(n3904), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3900) );
  OAI21_X1 U4868 ( .B1(n3901), .B2(n4819), .A(n3900), .ZN(U3460) );
  OAI22_X1 U4869 ( .A1(n5306), .A2(n3903), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n3902), .ZN(n6390) );
  NOR2_X1 U4870 ( .A1(n4812), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3905)
         );
  AOI211_X1 U4871 ( .C1(n6390), .C2(n5936), .A(n3905), .B(n3904), .ZN(n3909)
         );
  NOR2_X1 U4872 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n5940), .ZN(n3908)
         );
  NOR2_X1 U4873 ( .A1(n3906), .A2(n3017), .ZN(n6389) );
  INV_X1 U4874 ( .A(n6389), .ZN(n3907) );
  OAI22_X1 U4875 ( .A1(n3909), .A2(n3908), .B1(n6434), .B2(n3907), .ZN(U3461)
         );
  INV_X1 U4876 ( .A(n3910), .ZN(n4024) );
  NAND2_X1 U4877 ( .A1(n4038), .A2(n4024), .ZN(n3952) );
  NAND2_X1 U4878 ( .A1(n2995), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4068) );
  OR2_X1 U4879 ( .A1(n3952), .A2(n4068), .ZN(n4023) );
  NAND2_X1 U4880 ( .A1(n4023), .A2(n5723), .ZN(n3918) );
  AND2_X1 U4881 ( .A1(n4097), .A2(n4098), .ZN(n4393) );
  INV_X1 U4882 ( .A(n4671), .ZN(n4011) );
  NAND2_X1 U4883 ( .A1(n4393), .A2(n4011), .ZN(n4274) );
  OR2_X1 U4884 ( .A1(n4274), .A2(n5306), .ZN(n3912) );
  NAND2_X1 U4885 ( .A1(n3912), .A2(n6332), .ZN(n3917) );
  INV_X1 U4886 ( .A(n3917), .ZN(n3915) );
  NAND2_X1 U4887 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n3913), .ZN(n3914) );
  OAI21_X1 U4888 ( .B1(n3918), .B2(n3915), .A(n3914), .ZN(n6346) );
  INV_X1 U4889 ( .A(n6346), .ZN(n3939) );
  INV_X1 U4890 ( .A(DATAI_6_), .ZN(n6706) );
  NOR2_X1 U4891 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6546) );
  NOR2_X1 U4892 ( .A1(n6706), .A2(n4275), .ZN(n6373) );
  INV_X1 U4893 ( .A(n6373), .ZN(n5823) );
  AOI21_X1 U4894 ( .B1(n6388), .B2(STATE2_REG_3__SCAN_IN), .A(n4275), .ZN(
        n4462) );
  INV_X1 U4895 ( .A(n4619), .ZN(n5763) );
  NAND2_X1 U4896 ( .A1(n5763), .A2(n4268), .ZN(n3916) );
  OAI211_X1 U4897 ( .C1(n3918), .C2(n3917), .A(n4462), .B(n3916), .ZN(n6347)
         );
  NAND2_X1 U4898 ( .A1(n6347), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3924) );
  NOR2_X1 U4899 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4812), .ZN(n6535) );
  NAND2_X1 U4900 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6535), .ZN(n6443) );
  INV_X1 U4901 ( .A(n6443), .ZN(n3919) );
  NAND2_X1 U4902 ( .A1(n5723), .A2(n3919), .ZN(n6194) );
  INV_X2 U4903 ( .A(n6194), .ZN(n6219) );
  NAND2_X1 U4904 ( .A1(n6219), .A2(DATAI_30_), .ZN(n6376) );
  INV_X1 U4905 ( .A(n6376), .ZN(n5820) );
  NAND2_X1 U4906 ( .A1(n2995), .A2(n4398), .ZN(n4083) );
  OR2_X1 U4907 ( .A1(n3952), .A2(n4083), .ZN(n6350) );
  NAND2_X1 U4908 ( .A1(n3980), .A2(n3921), .ZN(n5818) );
  NAND2_X1 U4909 ( .A1(n6219), .A2(DATAI_22_), .ZN(n5817) );
  INV_X1 U4910 ( .A(n4041), .ZN(n4084) );
  OAI22_X1 U4911 ( .A1(n5818), .A2(n6332), .B1(n5817), .B2(n6333), .ZN(n3922)
         );
  AOI21_X1 U4912 ( .B1(n5820), .B2(n5272), .A(n3922), .ZN(n3923) );
  OAI211_X1 U4913 ( .C1(n3939), .C2(n5823), .A(n3924), .B(n3923), .ZN(U3082)
         );
  NOR2_X1 U4914 ( .A1(n3925), .A2(n4275), .ZN(n6355) );
  INV_X1 U4915 ( .A(n6355), .ZN(n5781) );
  NAND2_X1 U4916 ( .A1(n6347), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3928) );
  NAND2_X1 U4917 ( .A1(n6219), .A2(DATAI_24_), .ZN(n6358) );
  INV_X1 U4918 ( .A(n6358), .ZN(n5778) );
  NAND2_X1 U4919 ( .A1(n3980), .A2(n4452), .ZN(n5776) );
  NAND2_X1 U4920 ( .A1(n6219), .A2(DATAI_16_), .ZN(n5775) );
  OAI22_X1 U4921 ( .A1(n5776), .A2(n6332), .B1(n5775), .B2(n6333), .ZN(n3926)
         );
  AOI21_X1 U4922 ( .B1(n5778), .B2(n5272), .A(n3926), .ZN(n3927) );
  OAI211_X1 U4923 ( .C1(n3939), .C2(n5781), .A(n3928), .B(n3927), .ZN(U3076)
         );
  NOR2_X1 U4924 ( .A1(n3929), .A2(n4275), .ZN(n6313) );
  INV_X1 U4925 ( .A(n6313), .ZN(n5788) );
  NAND2_X1 U4926 ( .A1(n6347), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3933) );
  NAND2_X1 U4927 ( .A1(n6219), .A2(DATAI_25_), .ZN(n6316) );
  INV_X1 U4928 ( .A(n6316), .ZN(n5785) );
  NAND2_X1 U4929 ( .A1(n3980), .A2(n3930), .ZN(n5783) );
  NAND2_X1 U4930 ( .A1(n6219), .A2(DATAI_17_), .ZN(n5782) );
  OAI22_X1 U4931 ( .A1(n5783), .A2(n6332), .B1(n5782), .B2(n6333), .ZN(n3931)
         );
  AOI21_X1 U4932 ( .B1(n5785), .B2(n5272), .A(n3931), .ZN(n3932) );
  OAI211_X1 U4933 ( .C1(n3939), .C2(n5788), .A(n3933), .B(n3932), .ZN(U3077)
         );
  NOR2_X1 U4934 ( .A1(n3934), .A2(n4275), .ZN(n4478) );
  INV_X1 U4935 ( .A(n4478), .ZN(n5802) );
  NAND2_X1 U4936 ( .A1(n6347), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3938) );
  AND2_X1 U4937 ( .A1(n6219), .A2(DATAI_27_), .ZN(n5799) );
  NAND2_X1 U4938 ( .A1(n3980), .A2(n3935), .ZN(n5797) );
  NAND2_X1 U4939 ( .A1(n6219), .A2(DATAI_19_), .ZN(n5796) );
  OAI22_X1 U4940 ( .A1(n5797), .A2(n6332), .B1(n5796), .B2(n6333), .ZN(n3936)
         );
  AOI21_X1 U4941 ( .B1(n5799), .B2(n5272), .A(n3936), .ZN(n3937) );
  OAI211_X1 U4942 ( .C1(n3939), .C2(n5802), .A(n3938), .B(n3937), .ZN(U3079)
         );
  OAI21_X1 U4943 ( .B1(n3941), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n3940), 
        .ZN(n6302) );
  OAI222_X1 U4944 ( .A1(n6302), .A2(n6103), .B1(n5486), .B2(n5300), .C1(n5298), 
        .C2(n5466), .ZN(U2859) );
  NAND2_X1 U4945 ( .A1(n6394), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4465) );
  OR2_X1 U4946 ( .A1(n4465), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5716)
         );
  INV_X1 U4947 ( .A(n5716), .ZN(n3944) );
  NAND2_X1 U4948 ( .A1(n4098), .A2(n4609), .ZN(n4678) );
  NOR2_X1 U4949 ( .A1(n4678), .A2(n4671), .ZN(n5718) );
  NOR2_X1 U4950 ( .A1(n6388), .A2(n5716), .ZN(n3951) );
  AOI21_X1 U4951 ( .B1(n5718), .B2(n4131), .A(n3951), .ZN(n3942) );
  NOR2_X1 U4952 ( .A1(n3942), .A2(n5763), .ZN(n3943) );
  AOI21_X1 U4953 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n3944), .A(n3943), .ZN(
        n3985) );
  NOR2_X1 U4954 ( .A1(n3945), .A2(n4275), .ZN(n6361) );
  INV_X1 U4955 ( .A(n6361), .ZN(n5809) );
  NOR2_X1 U4956 ( .A1(n3952), .A2(n6538), .ZN(n3946) );
  NAND2_X1 U4957 ( .A1(n4619), .A2(n3946), .ZN(n3947) );
  NAND2_X1 U4958 ( .A1(n3947), .A2(n5716), .ZN(n3948) );
  NAND2_X1 U4959 ( .A1(n4462), .A2(n3948), .ZN(n3978) );
  NAND2_X1 U4960 ( .A1(n3978), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3955) );
  NAND2_X1 U4961 ( .A1(n6219), .A2(DATAI_20_), .ZN(n5803) );
  INV_X1 U4962 ( .A(n5803), .ZN(n6359) );
  OR2_X1 U4963 ( .A1(n2995), .A2(n4398), .ZN(n3949) );
  OR2_X1 U4964 ( .A1(n3952), .A2(n3949), .ZN(n4271) );
  NAND2_X1 U4965 ( .A1(n3980), .A2(n3950), .ZN(n5804) );
  INV_X1 U4966 ( .A(n3951), .ZN(n3981) );
  NAND2_X1 U4967 ( .A1(n6219), .A2(DATAI_28_), .ZN(n6364) );
  NOR3_X2 U4968 ( .A1(n3952), .A2(n4468), .A3(n2995), .ZN(n5758) );
  OAI22_X1 U4969 ( .A1(n5804), .A2(n3981), .B1(n6364), .B2(n5717), .ZN(n3953)
         );
  AOI21_X1 U4970 ( .B1(n6359), .B2(n5271), .A(n3953), .ZN(n3954) );
  OAI211_X1 U4971 ( .C1(n3985), .C2(n5809), .A(n3955), .B(n3954), .ZN(U3064)
         );
  NOR2_X1 U4972 ( .A1(n3956), .A2(n4275), .ZN(n6382) );
  INV_X1 U4973 ( .A(n6382), .ZN(n5833) );
  NAND2_X1 U4974 ( .A1(n3978), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3959) );
  NAND2_X1 U4975 ( .A1(n6219), .A2(DATAI_23_), .ZN(n5825) );
  INV_X1 U4976 ( .A(n5825), .ZN(n6378) );
  NAND2_X1 U4977 ( .A1(n3980), .A2(n5107), .ZN(n5827) );
  NAND2_X1 U4978 ( .A1(n6219), .A2(DATAI_31_), .ZN(n6387) );
  OAI22_X1 U4979 ( .A1(n5827), .A2(n3981), .B1(n6387), .B2(n5717), .ZN(n3957)
         );
  AOI21_X1 U4980 ( .B1(n6378), .B2(n5271), .A(n3957), .ZN(n3958) );
  OAI211_X1 U4981 ( .C1(n3985), .C2(n5833), .A(n3959), .B(n3958), .ZN(U3067)
         );
  NAND2_X1 U4982 ( .A1(n3978), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3962) );
  INV_X1 U4983 ( .A(n5817), .ZN(n6371) );
  OAI22_X1 U4984 ( .A1(n5818), .A2(n3981), .B1(n6376), .B2(n5717), .ZN(n3960)
         );
  AOI21_X1 U4985 ( .B1(n6371), .B2(n5271), .A(n3960), .ZN(n3961) );
  OAI211_X1 U4986 ( .C1(n3985), .C2(n5823), .A(n3962), .B(n3961), .ZN(U3066)
         );
  NAND2_X1 U4987 ( .A1(n3978), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3965) );
  OAI22_X1 U4988 ( .A1(n5797), .A2(n3981), .B1(n5796), .B2(n4271), .ZN(n3963)
         );
  AOI21_X1 U4989 ( .B1(n5799), .B2(n5758), .A(n3963), .ZN(n3964) );
  OAI211_X1 U4990 ( .C1(n3985), .C2(n5802), .A(n3965), .B(n3964), .ZN(U3063)
         );
  NAND2_X1 U4991 ( .A1(n3978), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3968) );
  INV_X1 U4992 ( .A(n5775), .ZN(n6353) );
  OAI22_X1 U4993 ( .A1(n5776), .A2(n3981), .B1(n6358), .B2(n5717), .ZN(n3966)
         );
  AOI21_X1 U4994 ( .B1(n6353), .B2(n5271), .A(n3966), .ZN(n3967) );
  OAI211_X1 U4995 ( .C1(n3985), .C2(n5781), .A(n3968), .B(n3967), .ZN(U3060)
         );
  NAND2_X1 U4996 ( .A1(n3978), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3971) );
  INV_X1 U4997 ( .A(n5782), .ZN(n6311) );
  OAI22_X1 U4998 ( .A1(n5783), .A2(n3981), .B1(n6316), .B2(n5717), .ZN(n3969)
         );
  AOI21_X1 U4999 ( .B1(n6311), .B2(n5271), .A(n3969), .ZN(n3970) );
  OAI211_X1 U5000 ( .C1(n3985), .C2(n5788), .A(n3971), .B(n3970), .ZN(U3061)
         );
  NOR2_X1 U5001 ( .A1(n3972), .A2(n4275), .ZN(n6336) );
  INV_X1 U5002 ( .A(n6336), .ZN(n5795) );
  NAND2_X1 U5003 ( .A1(n3978), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3976) );
  NAND2_X1 U5004 ( .A1(n6219), .A2(DATAI_18_), .ZN(n5789) );
  INV_X1 U5005 ( .A(n5789), .ZN(n6334) );
  NAND2_X1 U5006 ( .A1(n3980), .A2(n3973), .ZN(n5790) );
  NAND2_X1 U5007 ( .A1(n6219), .A2(DATAI_26_), .ZN(n6339) );
  OAI22_X1 U5008 ( .A1(n5790), .A2(n3981), .B1(n6339), .B2(n5717), .ZN(n3974)
         );
  AOI21_X1 U5009 ( .B1(n6334), .B2(n5271), .A(n3974), .ZN(n3975) );
  OAI211_X1 U5010 ( .C1(n3985), .C2(n5795), .A(n3976), .B(n3975), .ZN(U3062)
         );
  NOR2_X1 U5011 ( .A1(n3977), .A2(n4275), .ZN(n6367) );
  INV_X1 U5012 ( .A(n6367), .ZN(n5816) );
  NAND2_X1 U5013 ( .A1(n3978), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3984) );
  NAND2_X1 U5014 ( .A1(n6219), .A2(DATAI_21_), .ZN(n5810) );
  INV_X1 U5015 ( .A(n5810), .ZN(n6365) );
  NAND2_X1 U5016 ( .A1(n3980), .A2(n3979), .ZN(n5811) );
  NAND2_X1 U5017 ( .A1(n6219), .A2(DATAI_29_), .ZN(n6370) );
  OAI22_X1 U5018 ( .A1(n5811), .A2(n3981), .B1(n6370), .B2(n5717), .ZN(n3982)
         );
  AOI21_X1 U5019 ( .B1(n6365), .B2(n5271), .A(n3982), .ZN(n3983) );
  OAI211_X1 U5020 ( .C1(n3985), .C2(n5816), .A(n3984), .B(n3983), .ZN(U3065)
         );
  AOI22_X1 U5021 ( .A1(n5511), .A2(DATAI_1_), .B1(n6122), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n3986) );
  OAI21_X1 U5022 ( .B1(n3987), .B2(n5863), .A(n3986), .ZN(U2890) );
  INV_X1 U5023 ( .A(n4068), .ZN(n4124) );
  INV_X1 U5024 ( .A(n4031), .ZN(n4038) );
  XNOR2_X1 U5025 ( .A(n4124), .B(n4038), .ZN(n4022) );
  MUX2_X1 U5026 ( .A(n3988), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6391), 
        .Z(n6401) );
  INV_X1 U5027 ( .A(n3994), .ZN(n3990) );
  MUX2_X1 U5028 ( .A(n3990), .B(n3989), .S(n3993), .Z(n3992) );
  NOR2_X1 U5029 ( .A1(n3992), .A2(n3991), .ZN(n3999) );
  INV_X1 U5030 ( .A(n3993), .ZN(n4816) );
  NOR2_X1 U5031 ( .A1(n3994), .A2(n4816), .ZN(n3995) );
  AOI21_X1 U5032 ( .B1(n3996), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3995), 
        .ZN(n3998) );
  MUX2_X1 U5033 ( .A(n3999), .B(n3998), .S(n3997), .Z(n4003) );
  AOI21_X1 U5034 ( .B1(n4098), .B2(n4001), .A(n4000), .ZN(n4002) );
  NAND2_X1 U5035 ( .A1(n4003), .A2(n4002), .ZN(n4815) );
  NAND2_X1 U5036 ( .A1(n6391), .A2(n3997), .ZN(n4004) );
  OAI21_X1 U5037 ( .B1(n4815), .B2(n6391), .A(n4004), .ZN(n4005) );
  INV_X1 U5038 ( .A(n4005), .ZN(n6399) );
  NAND3_X1 U5039 ( .A1(n6401), .A2(n6399), .A3(n4812), .ZN(n4009) );
  NAND2_X1 U5040 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5948), .ZN(n4014) );
  INV_X1 U5041 ( .A(n4014), .ZN(n4006) );
  NAND2_X1 U5042 ( .A1(n4007), .A2(n4006), .ZN(n4008) );
  NAND2_X1 U5043 ( .A1(n4009), .A2(n4008), .ZN(n6414) );
  INV_X1 U5044 ( .A(n4010), .ZN(n4019) );
  NOR2_X1 U5045 ( .A1(n4012), .A2(n4011), .ZN(n4013) );
  XNOR2_X1 U5046 ( .A(n4013), .B(n5939), .ZN(n6072) );
  NOR2_X1 U5047 ( .A1(n5934), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4017) );
  NAND2_X1 U5048 ( .A1(n6391), .A2(n4812), .ZN(n4015) );
  AOI21_X1 U5049 ( .B1(n4015), .B2(n4014), .A(n5939), .ZN(n4016) );
  AOI21_X1 U5050 ( .B1(n6072), .B2(n4017), .A(n4016), .ZN(n6412) );
  INV_X1 U5051 ( .A(n6412), .ZN(n4018) );
  AOI21_X1 U5052 ( .B1(n6414), .B2(n4019), .A(n4018), .ZN(n6426) );
  NAND2_X1 U5053 ( .A1(n6426), .A2(n5948), .ZN(n4020) );
  INV_X1 U5054 ( .A(n6440), .ZN(n6521) );
  NAND2_X1 U5055 ( .A1(n4020), .A2(n6521), .ZN(n4021) );
  NAND2_X1 U5056 ( .A1(n4275), .A2(n4021), .ZN(n6310) );
  NAND2_X1 U5057 ( .A1(n6310), .A2(n5723), .ZN(n4123) );
  NAND2_X1 U5058 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5725), .ZN(n4027) );
  NAND2_X1 U5059 ( .A1(n6310), .A2(n4027), .ZN(n4129) );
  INV_X1 U5060 ( .A(n4098), .ZN(n6096) );
  OAI222_X1 U5061 ( .A1(n4022), .A2(n4123), .B1(n4129), .B2(n6096), .C1(n6400), 
        .C2(n6310), .ZN(U3463) );
  INV_X1 U5062 ( .A(n4681), .ZN(n5729) );
  INV_X1 U5063 ( .A(n4023), .ZN(n4025) );
  NOR2_X1 U5064 ( .A1(n4031), .A2(n4024), .ZN(n4292) );
  INV_X1 U5065 ( .A(n2995), .ZN(n4125) );
  NAND2_X1 U5066 ( .A1(n4292), .A2(n4125), .ZN(n4469) );
  INV_X1 U5067 ( .A(n4469), .ZN(n4293) );
  NAND2_X1 U5068 ( .A1(n4293), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4463) );
  NAND2_X1 U5069 ( .A1(n4039), .A2(n4031), .ZN(n4095) );
  NAND2_X1 U5070 ( .A1(n4463), .A2(n4095), .ZN(n4033) );
  AOI211_X1 U5071 ( .C1(n4039), .C2(n6538), .A(n4025), .B(n4033), .ZN(n4026)
         );
  OAI222_X1 U5072 ( .A1(n6310), .A2(n5765), .B1(n4129), .B2(n5729), .C1(n4123), 
        .C2(n4026), .ZN(U3462) );
  INV_X1 U5073 ( .A(n6310), .ZN(n4127) );
  AOI222_X1 U5074 ( .A1(n6426), .A2(n4028), .B1(n4131), .B2(n4027), .C1(n4468), 
        .C2(n5723), .ZN(n4030) );
  NAND2_X1 U5075 ( .A1(n4127), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4029) );
  OAI21_X1 U5076 ( .B1(n4127), .B2(n4030), .A(n4029), .ZN(U3465) );
  NAND2_X1 U5077 ( .A1(n4031), .A2(n4124), .ZN(n4032) );
  OAI21_X1 U5078 ( .B1(n4033), .B2(n4032), .A(n5723), .ZN(n4037) );
  OR2_X1 U5079 ( .A1(n4098), .A2(n4609), .ZN(n4070) );
  NOR2_X1 U5080 ( .A1(n4681), .A2(n4070), .ZN(n4531) );
  NOR2_X1 U5081 ( .A1(n4072), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6326)
         );
  AOI21_X1 U5082 ( .B1(n4531), .B2(n4131), .A(n6326), .ZN(n4034) );
  NAND3_X1 U5083 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n5765), .A3(n6400), .ZN(n4522) );
  OAI22_X1 U5084 ( .A1(n4037), .A2(n4034), .B1(n4522), .B2(n6532), .ZN(n6327)
         );
  INV_X1 U5085 ( .A(n6327), .ZN(n4049) );
  INV_X1 U5086 ( .A(n4034), .ZN(n4036) );
  INV_X1 U5087 ( .A(n4462), .ZN(n4079) );
  AOI21_X1 U5088 ( .B1(n4522), .B2(n5763), .A(n4079), .ZN(n4035) );
  OAI21_X1 U5089 ( .B1(n4037), .B2(n4036), .A(n4035), .ZN(n6328) );
  INV_X1 U5090 ( .A(n4130), .ZN(n4042) );
  INV_X1 U5091 ( .A(n4083), .ZN(n4040) );
  NAND2_X1 U5092 ( .A1(n4042), .A2(n4040), .ZN(n6331) );
  INV_X1 U5093 ( .A(n5776), .ZN(n6354) );
  NAND2_X1 U5094 ( .A1(n4042), .A2(n4041), .ZN(n5761) );
  INV_X1 U5095 ( .A(n5761), .ZN(n6325) );
  AOI22_X1 U5096 ( .A1(n6354), .A2(n6326), .B1(n6353), .B2(n6325), .ZN(n4043)
         );
  OAI21_X1 U5097 ( .B1(n6358), .B2(n6331), .A(n4043), .ZN(n4044) );
  AOI21_X1 U5098 ( .B1(n6328), .B2(INSTQUEUE_REG_3__0__SCAN_IN), .A(n4044), 
        .ZN(n4045) );
  OAI21_X1 U5099 ( .B1(n4049), .B2(n5781), .A(n4045), .ZN(U3044) );
  INV_X1 U5100 ( .A(n5799), .ZN(n5744) );
  INV_X1 U5101 ( .A(n5797), .ZN(n4479) );
  INV_X1 U5102 ( .A(n5796), .ZN(n5741) );
  AOI22_X1 U5103 ( .A1(n4479), .A2(n6326), .B1(n5741), .B2(n6325), .ZN(n4046)
         );
  OAI21_X1 U5104 ( .B1(n5744), .B2(n6331), .A(n4046), .ZN(n4047) );
  AOI21_X1 U5105 ( .B1(n6328), .B2(INSTQUEUE_REG_3__3__SCAN_IN), .A(n4047), 
        .ZN(n4048) );
  OAI21_X1 U5106 ( .B1(n4049), .B2(n5802), .A(n4048), .ZN(U3047) );
  INV_X1 U5107 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4062) );
  INV_X1 U5108 ( .A(n4051), .ZN(n4053) );
  INV_X1 U5109 ( .A(n4244), .ZN(n4052) );
  OAI21_X1 U5110 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n4053), .A(n4052), 
        .ZN(n6203) );
  AOI22_X1 U5111 ( .A1(n5216), .A2(n6203), .B1(n5219), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4054) );
  OAI21_X1 U5112 ( .B1(n5064), .B2(n4062), .A(n4054), .ZN(n4055) );
  NAND2_X1 U5113 ( .A1(n4060), .A2(n4059), .ZN(n4061) );
  AND2_X1 U5114 ( .A1(n4258), .A2(n4061), .ZN(n6206) );
  INV_X1 U5115 ( .A(n6206), .ZN(n4067) );
  OAI222_X1 U5116 ( .A1(n4067), .A2(n5863), .B1(n6131), .B2(n4062), .C1(n6126), 
        .C2(n3977), .ZN(U2886) );
  INV_X1 U5117 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4066) );
  AOI21_X1 U5118 ( .B1(n3823), .B2(n4064), .A(n4063), .ZN(n4065) );
  OR2_X1 U5119 ( .A1(n4158), .A2(n4065), .ZN(n6256) );
  OAI222_X1 U5120 ( .A1(n4067), .A2(n5466), .B1(n5486), .B2(n4066), .C1(n6256), 
        .C2(n6103), .ZN(U2854) );
  OR2_X1 U5121 ( .A1(n4095), .A2(n4068), .ZN(n4069) );
  AND2_X1 U5122 ( .A1(n4069), .A2(n5723), .ZN(n4078) );
  INV_X1 U5123 ( .A(n4070), .ZN(n4071) );
  AND2_X1 U5124 ( .A1(n4071), .A2(n4681), .ZN(n5769) );
  NAND2_X1 U5125 ( .A1(n5769), .A2(n4131), .ZN(n4074) );
  INV_X1 U5126 ( .A(n4072), .ZN(n4073) );
  NAND2_X1 U5127 ( .A1(n4073), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6351) );
  NAND2_X1 U5128 ( .A1(n4074), .A2(n6351), .ZN(n4081) );
  NAND2_X1 U5129 ( .A1(n4078), .A2(n4081), .ZN(n4077) );
  NAND3_X1 U5130 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6400), .ZN(n5770) );
  INV_X1 U5131 ( .A(n5770), .ZN(n4075) );
  NAND2_X1 U5132 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4075), .ZN(n4076) );
  NAND2_X1 U5133 ( .A1(n4077), .A2(n4076), .ZN(n6381) );
  INV_X1 U5134 ( .A(n6381), .ZN(n4094) );
  INV_X1 U5135 ( .A(n4078), .ZN(n4082) );
  AOI21_X1 U5136 ( .B1(n5770), .B2(n5763), .A(n4079), .ZN(n4080) );
  OAI21_X1 U5137 ( .B1(n4082), .B2(n4081), .A(n4080), .ZN(n6383) );
  NOR2_X1 U5138 ( .A1(n6386), .A2(n5744), .ZN(n4086) );
  OAI22_X1 U5139 ( .A1(n5797), .A2(n6351), .B1(n5796), .B2(n6352), .ZN(n4085)
         );
  AOI211_X1 U5140 ( .C1(n6383), .C2(INSTQUEUE_REG_11__3__SCAN_IN), .A(n4086), 
        .B(n4085), .ZN(n4087) );
  OAI21_X1 U5141 ( .B1(n4094), .B2(n5802), .A(n4087), .ZN(U3111) );
  NOR2_X1 U5142 ( .A1(n6386), .A2(n6316), .ZN(n4089) );
  OAI22_X1 U5143 ( .A1(n5783), .A2(n6351), .B1(n5782), .B2(n6352), .ZN(n4088)
         );
  AOI211_X1 U5144 ( .C1(n6383), .C2(INSTQUEUE_REG_11__1__SCAN_IN), .A(n4089), 
        .B(n4088), .ZN(n4090) );
  OAI21_X1 U5145 ( .B1(n4094), .B2(n5788), .A(n4090), .ZN(U3109) );
  NOR2_X1 U5146 ( .A1(n6386), .A2(n6339), .ZN(n4092) );
  OAI22_X1 U5147 ( .A1(n5790), .A2(n6351), .B1(n5789), .B2(n6352), .ZN(n4091)
         );
  AOI211_X1 U5148 ( .C1(n6383), .C2(INSTQUEUE_REG_11__2__SCAN_IN), .A(n4092), 
        .B(n4091), .ZN(n4093) );
  OAI21_X1 U5149 ( .B1(n4094), .B2(n5795), .A(n4093), .ZN(U3110) );
  INV_X1 U5150 ( .A(n4103), .ZN(n4096) );
  NAND2_X1 U5151 ( .A1(n4096), .A2(n4398), .ZN(n4173) );
  AOI21_X1 U5152 ( .B1(n4096), .B2(STATEBS16_REG_SCAN_IN), .A(n5763), .ZN(
        n4100) );
  NOR2_X1 U5153 ( .A1(n5729), .A2(n5306), .ZN(n4460) );
  NAND3_X1 U5154 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6400), .A3(n6394), .ZN(n4168) );
  NOR2_X1 U5155 ( .A1(n6388), .A2(n4168), .ZN(n4120) );
  AOI21_X1 U5156 ( .B1(n4460), .B2(n3011), .A(n4120), .ZN(n4102) );
  AOI22_X1 U5157 ( .A1(n4100), .A2(n4102), .B1(n5763), .B2(n4168), .ZN(n4099)
         );
  NAND2_X1 U5158 ( .A1(n4462), .A2(n4099), .ZN(n4119) );
  INV_X1 U5159 ( .A(n4100), .ZN(n4101) );
  OAI22_X1 U5160 ( .A1(n4102), .A2(n4101), .B1(n6532), .B2(n4168), .ZN(n4118)
         );
  AOI22_X1 U5161 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4119), .B1(n6382), 
        .B2(n4118), .ZN(n4105) );
  INV_X1 U5162 ( .A(n5827), .ZN(n6380) );
  NOR2_X2 U5163 ( .A1(n4103), .A2(n4398), .ZN(n5830) );
  AOI22_X1 U5164 ( .A1(n6380), .A2(n4120), .B1(n5830), .B2(n6378), .ZN(n4104)
         );
  OAI211_X1 U5165 ( .C1(n6387), .C2(n4173), .A(n4105), .B(n4104), .ZN(U3099)
         );
  AOI22_X1 U5166 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4119), .B1(n6367), 
        .B2(n4118), .ZN(n4107) );
  INV_X1 U5167 ( .A(n5811), .ZN(n6366) );
  AOI22_X1 U5168 ( .A1(n6366), .A2(n4120), .B1(n5830), .B2(n6365), .ZN(n4106)
         );
  OAI211_X1 U5169 ( .C1(n6370), .C2(n4173), .A(n4107), .B(n4106), .ZN(U3097)
         );
  AOI22_X1 U5170 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4119), .B1(n6361), 
        .B2(n4118), .ZN(n4109) );
  INV_X1 U5171 ( .A(n5804), .ZN(n6360) );
  AOI22_X1 U5172 ( .A1(n6360), .A2(n4120), .B1(n5830), .B2(n6359), .ZN(n4108)
         );
  OAI211_X1 U5173 ( .C1(n6364), .C2(n4173), .A(n4109), .B(n4108), .ZN(U3096)
         );
  AOI22_X1 U5174 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4119), .B1(n4478), 
        .B2(n4118), .ZN(n4111) );
  AOI22_X1 U5175 ( .A1(n4479), .A2(n4120), .B1(n5830), .B2(n5741), .ZN(n4110)
         );
  OAI211_X1 U5176 ( .C1(n5744), .C2(n4173), .A(n4111), .B(n4110), .ZN(U3095)
         );
  AOI22_X1 U5177 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4119), .B1(n6355), 
        .B2(n4118), .ZN(n4113) );
  AOI22_X1 U5178 ( .A1(n6354), .A2(n4120), .B1(n5830), .B2(n6353), .ZN(n4112)
         );
  OAI211_X1 U5179 ( .C1(n6358), .C2(n4173), .A(n4113), .B(n4112), .ZN(U3092)
         );
  AOI22_X1 U5180 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4119), .B1(n6313), 
        .B2(n4118), .ZN(n4115) );
  INV_X1 U5181 ( .A(n5783), .ZN(n6312) );
  AOI22_X1 U5182 ( .A1(n6312), .A2(n4120), .B1(n5830), .B2(n6311), .ZN(n4114)
         );
  OAI211_X1 U5183 ( .C1(n6316), .C2(n4173), .A(n4115), .B(n4114), .ZN(U3093)
         );
  AOI22_X1 U5184 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4119), .B1(n6373), 
        .B2(n4118), .ZN(n4117) );
  INV_X1 U5185 ( .A(n5818), .ZN(n6372) );
  AOI22_X1 U5186 ( .A1(n6372), .A2(n4120), .B1(n5830), .B2(n6371), .ZN(n4116)
         );
  OAI211_X1 U5187 ( .C1(n6376), .C2(n4173), .A(n4117), .B(n4116), .ZN(U3098)
         );
  AOI22_X1 U5188 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4119), .B1(n6336), 
        .B2(n4118), .ZN(n4122) );
  INV_X1 U5189 ( .A(n5790), .ZN(n6335) );
  AOI22_X1 U5190 ( .A1(n6335), .A2(n4120), .B1(n5830), .B2(n6334), .ZN(n4121)
         );
  OAI211_X1 U5191 ( .C1(n6339), .C2(n4173), .A(n4122), .B(n4121), .ZN(U3094)
         );
  AOI211_X1 U5192 ( .C1(n4125), .C2(n6538), .A(n4124), .B(n4123), .ZN(n4126)
         );
  AOI21_X1 U5193 ( .B1(n4127), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n4126), 
        .ZN(n4128) );
  OAI21_X1 U5194 ( .B1(n4609), .B2(n4129), .A(n4128), .ZN(U3464) );
  NAND2_X1 U5195 ( .A1(n5729), .A2(n3011), .ZN(n4615) );
  INV_X1 U5196 ( .A(n4615), .ZN(n4620) );
  NAND3_X1 U5197 ( .A1(n5765), .A2(n6400), .A3(n6394), .ZN(n4610) );
  NOR2_X1 U5198 ( .A1(n6388), .A2(n4610), .ZN(n4153) );
  AOI21_X1 U5199 ( .B1(n4620), .B2(n4131), .A(n4153), .ZN(n4135) );
  AOI21_X1 U5200 ( .B1(n4136), .B2(STATEBS16_REG_SCAN_IN), .A(n5763), .ZN(
        n4133) );
  AOI22_X1 U5201 ( .A1(n4135), .A2(n4133), .B1(n5763), .B2(n4610), .ZN(n4132)
         );
  NAND2_X1 U5202 ( .A1(n4462), .A2(n4132), .ZN(n4152) );
  INV_X1 U5203 ( .A(n4133), .ZN(n4134) );
  OAI22_X1 U5204 ( .A1(n4135), .A2(n4134), .B1(n6532), .B2(n4610), .ZN(n4151)
         );
  AOI22_X1 U5205 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4152), .B1(n6373), 
        .B2(n4151), .ZN(n4138) );
  NAND2_X1 U5206 ( .A1(n4136), .A2(n4468), .ZN(n4560) );
  AOI22_X1 U5207 ( .A1(n6372), .A2(n4153), .B1(n6371), .B2(n4524), .ZN(n4137)
         );
  OAI211_X1 U5208 ( .C1(n6376), .C2(n4649), .A(n4138), .B(n4137), .ZN(U3034)
         );
  AOI22_X1 U5209 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4152), .B1(n6355), 
        .B2(n4151), .ZN(n4140) );
  AOI22_X1 U5210 ( .A1(n6354), .A2(n4153), .B1(n6353), .B2(n4524), .ZN(n4139)
         );
  OAI211_X1 U5211 ( .C1(n6358), .C2(n4649), .A(n4140), .B(n4139), .ZN(U3028)
         );
  AOI22_X1 U5212 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4152), .B1(n6313), 
        .B2(n4151), .ZN(n4142) );
  AOI22_X1 U5213 ( .A1(n6312), .A2(n4153), .B1(n6311), .B2(n4524), .ZN(n4141)
         );
  OAI211_X1 U5214 ( .C1(n6316), .C2(n4649), .A(n4142), .B(n4141), .ZN(U3029)
         );
  AOI22_X1 U5215 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4152), .B1(n4478), 
        .B2(n4151), .ZN(n4144) );
  AOI22_X1 U5216 ( .A1(n4479), .A2(n4153), .B1(n5741), .B2(n4524), .ZN(n4143)
         );
  OAI211_X1 U5217 ( .C1(n5744), .C2(n4649), .A(n4144), .B(n4143), .ZN(U3031)
         );
  AOI22_X1 U5218 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4152), .B1(n6367), 
        .B2(n4151), .ZN(n4146) );
  AOI22_X1 U5219 ( .A1(n6366), .A2(n4153), .B1(n6365), .B2(n4524), .ZN(n4145)
         );
  OAI211_X1 U5220 ( .C1(n6370), .C2(n4649), .A(n4146), .B(n4145), .ZN(U3033)
         );
  AOI22_X1 U5221 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4152), .B1(n6361), 
        .B2(n4151), .ZN(n4148) );
  AOI22_X1 U5222 ( .A1(n6360), .A2(n4153), .B1(n6359), .B2(n4524), .ZN(n4147)
         );
  OAI211_X1 U5223 ( .C1(n6364), .C2(n4649), .A(n4148), .B(n4147), .ZN(U3032)
         );
  AOI22_X1 U5224 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4152), .B1(n6382), 
        .B2(n4151), .ZN(n4150) );
  AOI22_X1 U5225 ( .A1(n6380), .A2(n4153), .B1(n6378), .B2(n4524), .ZN(n4149)
         );
  OAI211_X1 U5226 ( .C1(n6387), .C2(n4649), .A(n4150), .B(n4149), .ZN(U3035)
         );
  AOI22_X1 U5227 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4152), .B1(n6336), 
        .B2(n4151), .ZN(n4155) );
  AOI22_X1 U5228 ( .A1(n6335), .A2(n4153), .B1(n6334), .B2(n4524), .ZN(n4154)
         );
  OAI211_X1 U5229 ( .C1(n6339), .C2(n4649), .A(n4155), .B(n4154), .ZN(U3030)
         );
  XNOR2_X1 U5230 ( .A(n4157), .B(n4156), .ZN(n4266) );
  XOR2_X1 U5231 ( .A(n4159), .B(n4158), .Z(n6062) );
  AND2_X1 U5232 ( .A1(n2997), .A2(REIP_REG_6__SCAN_IN), .ZN(n4261) );
  AOI21_X1 U5233 ( .B1(n4160), .B2(n6291), .A(n6264), .ZN(n4238) );
  NAND4_X1 U5234 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A3(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .A4(n6285), .ZN(n4163) );
  NOR2_X1 U5235 ( .A1(n4238), .A2(n4163), .ZN(n4165) );
  INV_X1 U5236 ( .A(n4160), .ZN(n4161) );
  AOI21_X1 U5237 ( .B1(n4161), .B2(n4232), .A(n4231), .ZN(n4162) );
  INV_X1 U5238 ( .A(n4162), .ZN(n6289) );
  AOI21_X1 U5239 ( .B1(n6236), .B2(n4163), .A(n6289), .ZN(n6262) );
  INV_X1 U5240 ( .A(n6262), .ZN(n4164) );
  MUX2_X1 U5241 ( .A(n4165), .B(n4164), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4166) );
  AOI211_X1 U5242 ( .C1(n6288), .C2(n6062), .A(n4261), .B(n4166), .ZN(n4167)
         );
  OAI21_X1 U5243 ( .B1(n6269), .B2(n4266), .A(n4167), .ZN(U3012) );
  NOR2_X1 U5244 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4168), .ZN(n4204)
         );
  AND2_X1 U5245 ( .A1(n4174), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5728) );
  INV_X1 U5246 ( .A(n5728), .ZN(n4299) );
  OR2_X1 U5247 ( .A1(n5768), .A2(n4611), .ZN(n4679) );
  AOI21_X1 U5248 ( .B1(n4679), .B2(STATE2_REG_2__SCAN_IN), .A(n4275), .ZN(
        n4674) );
  OAI211_X1 U5249 ( .C1(n5725), .C2(n4204), .A(n4299), .B(n4674), .ZN(n4172)
         );
  AOI21_X1 U5250 ( .B1(n4173), .B2(n6333), .A(n6538), .ZN(n4170) );
  NAND2_X1 U5251 ( .A1(n3011), .A2(n4681), .ZN(n4175) );
  INV_X1 U5252 ( .A(n4175), .ZN(n4169) );
  NOR3_X1 U5253 ( .A1(n4170), .A2(n4169), .A3(n5763), .ZN(n4171) );
  NOR2_X1 U5254 ( .A1(n4172), .A2(n4171), .ZN(n4210) );
  INV_X1 U5255 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4179) );
  INV_X1 U5256 ( .A(n4173), .ZN(n4207) );
  NOR2_X1 U5257 ( .A1(n4174), .A2(n6532), .ZN(n5721) );
  INV_X1 U5258 ( .A(n5721), .ZN(n5766) );
  OAI22_X1 U5259 ( .A1(n4175), .A2(n5763), .B1(n5766), .B2(n4679), .ZN(n4203)
         );
  AOI22_X1 U5260 ( .A1(n6312), .A2(n4204), .B1(n6313), .B2(n4203), .ZN(n4176)
         );
  OAI21_X1 U5261 ( .B1(n6316), .B2(n6333), .A(n4176), .ZN(n4177) );
  AOI21_X1 U5262 ( .B1(n6311), .B2(n4207), .A(n4177), .ZN(n4178) );
  OAI21_X1 U5263 ( .B1(n4210), .B2(n4179), .A(n4178), .ZN(U3085) );
  INV_X1 U5264 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4183) );
  AOI22_X1 U5265 ( .A1(n6335), .A2(n4204), .B1(n6336), .B2(n4203), .ZN(n4180)
         );
  OAI21_X1 U5266 ( .B1(n6339), .B2(n6333), .A(n4180), .ZN(n4181) );
  AOI21_X1 U5267 ( .B1(n6334), .B2(n4207), .A(n4181), .ZN(n4182) );
  OAI21_X1 U5268 ( .B1(n4210), .B2(n4183), .A(n4182), .ZN(U3086) );
  INV_X1 U5269 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4187) );
  AOI22_X1 U5270 ( .A1(n6372), .A2(n4204), .B1(n6373), .B2(n4203), .ZN(n4184)
         );
  OAI21_X1 U5271 ( .B1(n6376), .B2(n6333), .A(n4184), .ZN(n4185) );
  AOI21_X1 U5272 ( .B1(n6371), .B2(n4207), .A(n4185), .ZN(n4186) );
  OAI21_X1 U5273 ( .B1(n4210), .B2(n4187), .A(n4186), .ZN(U3090) );
  INV_X1 U5274 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4191) );
  AOI22_X1 U5275 ( .A1(n4479), .A2(n4204), .B1(n4478), .B2(n4203), .ZN(n4188)
         );
  OAI21_X1 U5276 ( .B1(n5744), .B2(n6333), .A(n4188), .ZN(n4189) );
  AOI21_X1 U5277 ( .B1(n5741), .B2(n4207), .A(n4189), .ZN(n4190) );
  OAI21_X1 U5278 ( .B1(n4210), .B2(n4191), .A(n4190), .ZN(U3087) );
  INV_X1 U5279 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4195) );
  AOI22_X1 U5280 ( .A1(n6354), .A2(n4204), .B1(n6355), .B2(n4203), .ZN(n4192)
         );
  OAI21_X1 U5281 ( .B1(n6358), .B2(n6333), .A(n4192), .ZN(n4193) );
  AOI21_X1 U5282 ( .B1(n6353), .B2(n4207), .A(n4193), .ZN(n4194) );
  OAI21_X1 U5283 ( .B1(n4210), .B2(n4195), .A(n4194), .ZN(U3084) );
  INV_X1 U5284 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6722) );
  AOI22_X1 U5285 ( .A1(n6366), .A2(n4204), .B1(n6367), .B2(n4203), .ZN(n4196)
         );
  OAI21_X1 U5286 ( .B1(n6370), .B2(n6333), .A(n4196), .ZN(n4197) );
  AOI21_X1 U5287 ( .B1(n6365), .B2(n4207), .A(n4197), .ZN(n4198) );
  OAI21_X1 U5288 ( .B1(n4210), .B2(n6722), .A(n4198), .ZN(U3089) );
  INV_X1 U5289 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4202) );
  AOI22_X1 U5290 ( .A1(n6360), .A2(n4204), .B1(n6361), .B2(n4203), .ZN(n4199)
         );
  OAI21_X1 U5291 ( .B1(n6364), .B2(n6333), .A(n4199), .ZN(n4200) );
  AOI21_X1 U5292 ( .B1(n6359), .B2(n4207), .A(n4200), .ZN(n4201) );
  OAI21_X1 U5293 ( .B1(n4210), .B2(n4202), .A(n4201), .ZN(U3088) );
  INV_X1 U5294 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4209) );
  AOI22_X1 U5295 ( .A1(n6380), .A2(n4204), .B1(n6382), .B2(n4203), .ZN(n4205)
         );
  OAI21_X1 U5296 ( .B1(n6387), .B2(n6333), .A(n4205), .ZN(n4206) );
  AOI21_X1 U5297 ( .B1(n6378), .B2(n4207), .A(n4206), .ZN(n4208) );
  OAI21_X1 U5298 ( .B1(n4210), .B2(n4209), .A(n4208), .ZN(U3091) );
  XNOR2_X1 U5299 ( .A(n4212), .B(n4211), .ZN(n6276) );
  NOR2_X1 U5300 ( .A1(n6410), .A2(n6432), .ZN(n4214) );
  NAND2_X2 U5301 ( .A1(n4214), .A2(n4213), .ZN(n6195) );
  INV_X1 U5302 ( .A(n4215), .ZN(n6109) );
  NAND2_X1 U5303 ( .A1(n5763), .A2(n4216), .ZN(n6534) );
  NAND2_X1 U5304 ( .A1(n6534), .A2(n6540), .ZN(n4217) );
  NAND2_X1 U5305 ( .A1(n6540), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4219) );
  NAND2_X1 U5306 ( .A1(n6538), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4218) );
  NAND2_X1 U5307 ( .A1(n4219), .A2(n4218), .ZN(n5627) );
  AOI22_X1 U5308 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n2997), 
        .B2(REIP_REG_3__SCAN_IN), .ZN(n4220) );
  OAI21_X1 U5309 ( .B1(n4592), .B2(n6225), .A(n4220), .ZN(n4221) );
  AOI21_X1 U5310 ( .B1(n6109), .B2(n6219), .A(n4221), .ZN(n4222) );
  OAI21_X1 U5311 ( .B1(n6276), .B2(n6195), .A(n4222), .ZN(U2983) );
  XNOR2_X1 U5312 ( .A(n4224), .B(n4223), .ZN(n6270) );
  INV_X1 U5313 ( .A(n4225), .ZN(n6081) );
  AND2_X1 U5314 ( .A1(n2997), .A2(REIP_REG_4__SCAN_IN), .ZN(n6265) );
  AOI21_X1 U5315 ( .B1(n6218), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6265), 
        .ZN(n4226) );
  OAI21_X1 U5316 ( .B1(n6078), .B2(n6225), .A(n4226), .ZN(n4227) );
  AOI21_X1 U5317 ( .B1(n6081), .B2(n6219), .A(n4227), .ZN(n4228) );
  OAI21_X1 U5318 ( .B1(n6195), .B2(n6270), .A(n4228), .ZN(U2982) );
  XNOR2_X1 U5319 ( .A(n4230), .B(n4229), .ZN(n6196) );
  AOI21_X1 U5320 ( .B1(n4233), .B2(n4232), .A(n4231), .ZN(n4713) );
  OAI21_X1 U5321 ( .B1(n4234), .B2(n6283), .A(n4713), .ZN(n6235) );
  NAND2_X1 U5322 ( .A1(n4236), .A2(n4235), .ZN(n4237) );
  NAND2_X1 U5323 ( .A1(n4333), .A2(n4237), .ZN(n6038) );
  NAND2_X1 U5324 ( .A1(n2997), .A2(REIP_REG_7__SCAN_IN), .ZN(n6199) );
  OAI21_X1 U5325 ( .B1(n6038), .B2(n6303), .A(n6199), .ZN(n4241) );
  INV_X1 U5326 ( .A(n6285), .ZN(n6263) );
  NOR2_X1 U5327 ( .A1(n6263), .A2(n4238), .ZN(n6275) );
  NAND2_X1 U5328 ( .A1(n4239), .A2(n6275), .ZN(n6241) );
  NOR2_X1 U5329 ( .A1(n6241), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4240)
         );
  AOI211_X1 U5330 ( .C1(n6235), .C2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n4241), 
        .B(n4240), .ZN(n4242) );
  OAI21_X1 U5331 ( .B1(n6269), .B2(n6196), .A(n4242), .ZN(U3011) );
  NAND2_X1 U5332 ( .A1(n4244), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4248)
         );
  OAI21_X1 U5333 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n4244), .A(n4248), 
        .ZN(n6064) );
  INV_X1 U5334 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4267) );
  INV_X1 U5335 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6054) );
  OAI22_X1 U5336 ( .A1(n5064), .A2(n4267), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6054), .ZN(n4245) );
  MUX2_X1 U5337 ( .A(n6064), .B(n4245), .S(n5210), .Z(n4246) );
  INV_X1 U5338 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4255) );
  OAI21_X1 U5339 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n4249), .A(n4349), 
        .ZN(n6197) );
  AOI22_X1 U5340 ( .A1(n5216), .A2(n6197), .B1(n5219), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4250) );
  OAI21_X1 U5341 ( .B1(n5064), .B2(n4255), .A(n4250), .ZN(n4251) );
  AND2_X1 U5342 ( .A1(n4256), .A2(n4253), .ZN(n4254) );
  OR2_X1 U5343 ( .A1(n4254), .A2(n4355), .ZN(n6193) );
  OAI222_X1 U5344 ( .A1(n6193), .A2(n5863), .B1(n6131), .B2(n4255), .C1(n6126), 
        .C2(n3956), .ZN(U2884) );
  INV_X1 U5345 ( .A(n4256), .ZN(n4257) );
  AOI21_X1 U5346 ( .B1(n4259), .B2(n4258), .A(n4257), .ZN(n4264) );
  INV_X1 U5347 ( .A(n4264), .ZN(n6059) );
  AOI22_X1 U5348 ( .A1(n6062), .A2(n6107), .B1(n5399), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4260) );
  OAI21_X1 U5349 ( .B1(n6059), .B2(n5466), .A(n4260), .ZN(U2853) );
  AOI21_X1 U5350 ( .B1(n6218), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n4261), 
        .ZN(n4262) );
  OAI21_X1 U5351 ( .B1(n6064), .B2(n6225), .A(n4262), .ZN(n4263) );
  AOI21_X1 U5352 ( .B1(n4264), .B2(n6219), .A(n4263), .ZN(n4265) );
  OAI21_X1 U5353 ( .B1(n6195), .B2(n4266), .A(n4265), .ZN(U2980) );
  OAI222_X1 U5354 ( .A1(n6059), .A2(n5863), .B1(n6126), .B2(n6706), .C1(n4267), 
        .C2(n6131), .ZN(U2885) );
  INV_X1 U5355 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6042) );
  OAI222_X1 U5356 ( .A1(n6038), .A2(n6103), .B1(n5486), .B2(n6042), .C1(n5466), 
        .C2(n6193), .ZN(U2852) );
  OR2_X1 U5357 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4268), .ZN(n5275)
         );
  NAND3_X1 U5358 ( .A1(n5729), .A2(n5723), .A3(n4393), .ZN(n4270) );
  NAND3_X1 U5359 ( .A1(n5728), .A2(n5768), .A3(n5765), .ZN(n4269) );
  NAND2_X1 U5360 ( .A1(n4270), .A2(n4269), .ZN(n5270) );
  NAND2_X1 U5361 ( .A1(n5723), .A2(n6538), .ZN(n4523) );
  NAND3_X1 U5362 ( .A1(n5723), .A2(n4271), .A3(n6350), .ZN(n4272) );
  NAND2_X1 U5363 ( .A1(n4523), .A2(n4272), .ZN(n4273) );
  AOI22_X1 U5364 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5275), .B1(n4274), .B2(
        n4273), .ZN(n4276) );
  INV_X1 U5365 ( .A(n4275), .ZN(n4613) );
  OAI21_X1 U5366 ( .B1(n5768), .B2(n6532), .A(n4613), .ZN(n4527) );
  NOR2_X1 U5367 ( .A1(n5721), .A2(n4527), .ZN(n4295) );
  NAND3_X1 U5368 ( .A1(n5765), .A2(n4276), .A3(n4295), .ZN(n5269) );
  AOI22_X1 U5369 ( .A1(n5270), .A2(n6373), .B1(INSTQUEUE_REG_6__6__SCAN_IN), 
        .B2(n5269), .ZN(n4278) );
  AOI22_X1 U5370 ( .A1(n6371), .A2(n5272), .B1(n5271), .B2(n5820), .ZN(n4277)
         );
  OAI211_X1 U5371 ( .C1(n5818), .C2(n5275), .A(n4278), .B(n4277), .ZN(U3074)
         );
  AOI22_X1 U5372 ( .A1(n5270), .A2(n6382), .B1(INSTQUEUE_REG_6__7__SCAN_IN), 
        .B2(n5269), .ZN(n4280) );
  INV_X1 U5373 ( .A(n6387), .ZN(n5829) );
  AOI22_X1 U5374 ( .A1(n6378), .A2(n5272), .B1(n5271), .B2(n5829), .ZN(n4279)
         );
  OAI211_X1 U5375 ( .C1(n5827), .C2(n5275), .A(n4280), .B(n4279), .ZN(U3075)
         );
  AOI22_X1 U5376 ( .A1(n5270), .A2(n4478), .B1(INSTQUEUE_REG_6__3__SCAN_IN), 
        .B2(n5269), .ZN(n4282) );
  AOI22_X1 U5377 ( .A1(n5741), .A2(n5272), .B1(n5271), .B2(n5799), .ZN(n4281)
         );
  OAI211_X1 U5378 ( .C1(n5797), .C2(n5275), .A(n4282), .B(n4281), .ZN(U3071)
         );
  AOI22_X1 U5379 ( .A1(n5270), .A2(n6336), .B1(INSTQUEUE_REG_6__2__SCAN_IN), 
        .B2(n5269), .ZN(n4284) );
  INV_X1 U5380 ( .A(n6339), .ZN(n5792) );
  AOI22_X1 U5381 ( .A1(n6334), .A2(n5272), .B1(n5271), .B2(n5792), .ZN(n4283)
         );
  OAI211_X1 U5382 ( .C1(n5790), .C2(n5275), .A(n4284), .B(n4283), .ZN(U3070)
         );
  AOI22_X1 U5383 ( .A1(n5270), .A2(n6361), .B1(INSTQUEUE_REG_6__4__SCAN_IN), 
        .B2(n5269), .ZN(n4286) );
  INV_X1 U5384 ( .A(n6364), .ZN(n5806) );
  AOI22_X1 U5385 ( .A1(n6359), .A2(n5272), .B1(n5271), .B2(n5806), .ZN(n4285)
         );
  OAI211_X1 U5386 ( .C1(n5804), .C2(n5275), .A(n4286), .B(n4285), .ZN(U3072)
         );
  AOI22_X1 U5387 ( .A1(n5270), .A2(n6313), .B1(INSTQUEUE_REG_6__1__SCAN_IN), 
        .B2(n5269), .ZN(n4288) );
  AOI22_X1 U5388 ( .A1(n6311), .A2(n5272), .B1(n5271), .B2(n5785), .ZN(n4287)
         );
  OAI211_X1 U5389 ( .C1(n5783), .C2(n5275), .A(n4288), .B(n4287), .ZN(U3069)
         );
  AOI22_X1 U5390 ( .A1(n5270), .A2(n6355), .B1(INSTQUEUE_REG_6__0__SCAN_IN), 
        .B2(n5269), .ZN(n4290) );
  AOI22_X1 U5391 ( .A1(n6353), .A2(n5272), .B1(n5271), .B2(n5778), .ZN(n4289)
         );
  OAI211_X1 U5392 ( .C1(n5776), .C2(n5275), .A(n4290), .B(n4289), .ZN(U3068)
         );
  NAND2_X1 U5393 ( .A1(n4292), .A2(n2995), .ZN(n4399) );
  INV_X1 U5394 ( .A(n4399), .ZN(n4394) );
  NAND2_X1 U5395 ( .A1(n4394), .A2(n4398), .ZN(n4430) );
  NAND2_X1 U5396 ( .A1(n4293), .A2(n4468), .ZN(n4491) );
  AOI21_X1 U5397 ( .B1(n4430), .B2(n4491), .A(n6538), .ZN(n4297) );
  NAND2_X1 U5398 ( .A1(n4393), .A2(n4681), .ZN(n4298) );
  NAND2_X1 U5399 ( .A1(n4298), .A2(n5723), .ZN(n4296) );
  OR2_X1 U5400 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4395), .ZN(n4325)
         );
  AOI21_X1 U5401 ( .B1(n4325), .B2(STATE2_REG_3__SCAN_IN), .A(n5765), .ZN(
        n4294) );
  OAI211_X1 U5402 ( .C1(n4297), .C2(n4296), .A(n4295), .B(n4294), .ZN(n4323)
         );
  NAND2_X1 U5403 ( .A1(n4323), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4304)
         );
  INV_X1 U5404 ( .A(n4491), .ZN(n4327) );
  INV_X1 U5405 ( .A(n4298), .ZN(n4301) );
  NOR2_X1 U5406 ( .A1(n4299), .A2(n5765), .ZN(n4300) );
  AOI22_X1 U5407 ( .A1(n4301), .A2(n4619), .B1(n5768), .B2(n4300), .ZN(n4324)
         );
  OAI22_X1 U5408 ( .A1(n5804), .A2(n4325), .B1(n4324), .B2(n5809), .ZN(n4302)
         );
  AOI21_X1 U5409 ( .B1(n5806), .B2(n4327), .A(n4302), .ZN(n4303) );
  OAI211_X1 U5410 ( .C1(n4430), .C2(n5803), .A(n4304), .B(n4303), .ZN(U3136)
         );
  NAND2_X1 U5411 ( .A1(n4323), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4307)
         );
  OAI22_X1 U5412 ( .A1(n5790), .A2(n4325), .B1(n4324), .B2(n5795), .ZN(n4305)
         );
  AOI21_X1 U5413 ( .B1(n5792), .B2(n4327), .A(n4305), .ZN(n4306) );
  OAI211_X1 U5414 ( .C1(n4430), .C2(n5789), .A(n4307), .B(n4306), .ZN(U3134)
         );
  NAND2_X1 U5415 ( .A1(n4323), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4310)
         );
  OAI22_X1 U5416 ( .A1(n5783), .A2(n4325), .B1(n4324), .B2(n5788), .ZN(n4308)
         );
  AOI21_X1 U5417 ( .B1(n5785), .B2(n4327), .A(n4308), .ZN(n4309) );
  OAI211_X1 U5418 ( .C1(n4430), .C2(n5782), .A(n4310), .B(n4309), .ZN(U3133)
         );
  NAND2_X1 U5419 ( .A1(n4323), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4313)
         );
  INV_X1 U5420 ( .A(n6370), .ZN(n5813) );
  OAI22_X1 U5421 ( .A1(n5811), .A2(n4325), .B1(n4324), .B2(n5816), .ZN(n4311)
         );
  AOI21_X1 U5422 ( .B1(n5813), .B2(n4327), .A(n4311), .ZN(n4312) );
  OAI211_X1 U5423 ( .C1(n4430), .C2(n5810), .A(n4313), .B(n4312), .ZN(U3137)
         );
  NAND2_X1 U5424 ( .A1(n4323), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4316)
         );
  OAI22_X1 U5425 ( .A1(n5818), .A2(n4325), .B1(n4324), .B2(n5823), .ZN(n4314)
         );
  AOI21_X1 U5426 ( .B1(n5820), .B2(n4327), .A(n4314), .ZN(n4315) );
  OAI211_X1 U5427 ( .C1(n4430), .C2(n5817), .A(n4316), .B(n4315), .ZN(U3138)
         );
  NAND2_X1 U5428 ( .A1(n4323), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4319)
         );
  OAI22_X1 U5429 ( .A1(n5827), .A2(n4325), .B1(n4324), .B2(n5833), .ZN(n4317)
         );
  AOI21_X1 U5430 ( .B1(n5829), .B2(n4327), .A(n4317), .ZN(n4318) );
  OAI211_X1 U5431 ( .C1(n4430), .C2(n5825), .A(n4319), .B(n4318), .ZN(U3139)
         );
  NAND2_X1 U5432 ( .A1(n4323), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4322)
         );
  OAI22_X1 U5433 ( .A1(n5797), .A2(n4325), .B1(n4324), .B2(n5802), .ZN(n4320)
         );
  AOI21_X1 U5434 ( .B1(n5799), .B2(n4327), .A(n4320), .ZN(n4321) );
  OAI211_X1 U5435 ( .C1(n4430), .C2(n5796), .A(n4322), .B(n4321), .ZN(U3135)
         );
  NAND2_X1 U5436 ( .A1(n4323), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4329)
         );
  OAI22_X1 U5437 ( .A1(n5776), .A2(n4325), .B1(n4324), .B2(n5781), .ZN(n4326)
         );
  AOI21_X1 U5438 ( .B1(n5778), .B2(n4327), .A(n4326), .ZN(n4328) );
  OAI211_X1 U5439 ( .C1(n4430), .C2(n5775), .A(n4329), .B(n4328), .ZN(U3132)
         );
  XNOR2_X1 U5440 ( .A(n4331), .B(n4330), .ZN(n4391) );
  NAND2_X1 U5441 ( .A1(n4333), .A2(n4332), .ZN(n4334) );
  NAND2_X1 U5442 ( .A1(n4382), .A2(n4334), .ZN(n6028) );
  NAND2_X1 U5443 ( .A1(n2997), .A2(REIP_REG_8__SCAN_IN), .ZN(n4388) );
  OAI21_X1 U5444 ( .B1(n6028), .B2(n6303), .A(n4388), .ZN(n4337) );
  OAI21_X1 U5445 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6242), .ZN(n4335) );
  NOR2_X1 U5446 ( .A1(n6241), .A2(n4335), .ZN(n4336) );
  AOI211_X1 U5447 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n6235), .A(n4337), 
        .B(n4336), .ZN(n4338) );
  OAI21_X1 U5448 ( .B1(n6269), .B2(n4391), .A(n4338), .ZN(U3010) );
  INV_X1 U5449 ( .A(EAX_REG_8__SCAN_IN), .ZN(n4385) );
  AOI22_X1 U5450 ( .A1(n5185), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5187), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4342) );
  AOI22_X1 U5451 ( .A1(n5195), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4341) );
  AOI22_X1 U5452 ( .A1(n5197), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4340) );
  AOI22_X1 U5453 ( .A1(n2999), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4339) );
  NAND4_X1 U5454 ( .A1(n4342), .A2(n4341), .A3(n4340), .A4(n4339), .ZN(n4348)
         );
  AOI22_X1 U5455 ( .A1(n5198), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4346) );
  AOI22_X1 U5456 ( .A1(n5024), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5189), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4345) );
  AOI22_X1 U5457 ( .A1(n5186), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4344) );
  AOI22_X1 U5458 ( .A1(n5167), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4343) );
  NAND4_X1 U5459 ( .A1(n4346), .A2(n4345), .A3(n4344), .A4(n4343), .ZN(n4347)
         );
  OAI21_X1 U5460 ( .B1(n4348), .B2(n4347), .A(n4998), .ZN(n4353) );
  INV_X1 U5461 ( .A(n4349), .ZN(n4351) );
  INV_X1 U5462 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6658) );
  INV_X1 U5463 ( .A(n4435), .ZN(n4350) );
  OAI21_X1 U5464 ( .B1(PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n4351), .A(n4350), 
        .ZN(n6030) );
  AOI22_X1 U5465 ( .A1(n5216), .A2(n6030), .B1(n5219), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4352) );
  OAI211_X1 U5466 ( .C1(n5064), .C2(n4385), .A(n4353), .B(n4352), .ZN(n4354)
         );
  INV_X1 U5467 ( .A(n4354), .ZN(n4357) );
  INV_X1 U5468 ( .A(n4355), .ZN(n4356) );
  INV_X1 U5469 ( .A(n4376), .ZN(n4379) );
  AOI21_X1 U5470 ( .B1(n4357), .B2(n4356), .A(n4379), .ZN(n6033) );
  INV_X1 U5471 ( .A(n5466), .ZN(n6108) );
  OAI22_X1 U5472 ( .A1(n6028), .A2(n6103), .B1(n4358), .B2(n5486), .ZN(n4359)
         );
  AOI21_X1 U5473 ( .B1(n6033), .B2(n6108), .A(n4359), .ZN(n4360) );
  INV_X1 U5474 ( .A(n4360), .ZN(U2851) );
  AOI22_X1 U5475 ( .A1(n5197), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4364) );
  AOI22_X1 U5476 ( .A1(n5187), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4363) );
  AOI22_X1 U5477 ( .A1(n5167), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4362) );
  AOI22_X1 U5478 ( .A1(n5024), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4361) );
  NAND4_X1 U5479 ( .A1(n4364), .A2(n4363), .A3(n4362), .A4(n4361), .ZN(n4370)
         );
  AOI22_X1 U5480 ( .A1(n5185), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4368) );
  AOI22_X1 U5481 ( .A1(n5195), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5189), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4367) );
  AOI22_X1 U5482 ( .A1(n2999), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4366) );
  AOI22_X1 U5483 ( .A1(n5198), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4365) );
  NAND4_X1 U5484 ( .A1(n4368), .A2(n4367), .A3(n4366), .A4(n4365), .ZN(n4369)
         );
  OAI21_X1 U5485 ( .B1(n4370), .B2(n4369), .A(n4998), .ZN(n4374) );
  XOR2_X1 U5486 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n4435), .Z(n4517) );
  INV_X1 U5487 ( .A(n4517), .ZN(n4371) );
  AOI22_X1 U5488 ( .A1(n5219), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .B1(n5216), 
        .B2(n4371), .ZN(n4373) );
  NAND2_X1 U5489 ( .A1(n5158), .A2(EAX_REG_9__SCAN_IN), .ZN(n4372) );
  AND3_X1 U5490 ( .A1(n4374), .A2(n4373), .A3(n4372), .ZN(n4375) );
  INV_X1 U5491 ( .A(n4375), .ZN(n4378) );
  INV_X1 U5492 ( .A(n4377), .ZN(n4506) );
  OAI21_X1 U5493 ( .B1(n4379), .B2(n4378), .A(n4506), .ZN(n4520) );
  AOI22_X1 U5494 ( .A1(n5511), .A2(DATAI_9_), .B1(n6122), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4380) );
  OAI21_X1 U5495 ( .B1(n4520), .B2(n5863), .A(n4380), .ZN(U2882) );
  AND2_X1 U5496 ( .A1(n4382), .A2(n4381), .ZN(n4383) );
  NOR2_X1 U5497 ( .A1(n4509), .A2(n4383), .ZN(n6249) );
  AOI22_X1 U5498 ( .A1(n6249), .A2(n6107), .B1(EBX_REG_9__SCAN_IN), .B2(n5399), 
        .ZN(n4384) );
  OAI21_X1 U5499 ( .B1(n4520), .B2(n5466), .A(n4384), .ZN(U2850) );
  INV_X1 U5500 ( .A(n6033), .ZN(n4386) );
  OAI222_X1 U5501 ( .A1(n4386), .A2(n5863), .B1(n6131), .B2(n4385), .C1(n6126), 
        .C2(n3694), .ZN(U2883) );
  NAND2_X1 U5502 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4387)
         );
  OAI211_X1 U5503 ( .C1(n6225), .C2(n6030), .A(n4388), .B(n4387), .ZN(n4389)
         );
  AOI21_X1 U5504 ( .B1(n6033), .B2(n6219), .A(n4389), .ZN(n4390) );
  OAI21_X1 U5505 ( .B1(n6195), .B2(n4391), .A(n4390), .ZN(U2978) );
  INV_X1 U5506 ( .A(n4426), .ZN(n4392) );
  AOI21_X1 U5507 ( .B1(n4460), .B2(n4393), .A(n4392), .ZN(n4400) );
  OAI21_X1 U5508 ( .B1(n4394), .B2(n6194), .A(n4523), .ZN(n4396) );
  AOI22_X1 U5509 ( .A1(n4400), .A2(n4396), .B1(n4395), .B2(n5763), .ZN(n4397)
         );
  NAND2_X1 U5510 ( .A1(n4462), .A2(n4397), .ZN(n4424) );
  NAND2_X1 U5511 ( .A1(n4424), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4405)
         );
  NOR2_X2 U5512 ( .A1(n4399), .A2(n4398), .ZN(n4646) );
  INV_X1 U5513 ( .A(n4400), .ZN(n4402) );
  AOI22_X1 U5514 ( .A1(n4402), .A2(n5723), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4401), .ZN(n4425) );
  OAI22_X1 U5515 ( .A1(n5797), .A2(n4426), .B1(n4425), .B2(n5802), .ZN(n4403)
         );
  AOI21_X1 U5516 ( .B1(n5741), .B2(n4646), .A(n4403), .ZN(n4404) );
  OAI211_X1 U5517 ( .C1(n4430), .C2(n5744), .A(n4405), .B(n4404), .ZN(U3143)
         );
  NAND2_X1 U5518 ( .A1(n4424), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4408)
         );
  OAI22_X1 U5519 ( .A1(n5804), .A2(n4426), .B1(n4425), .B2(n5809), .ZN(n4406)
         );
  AOI21_X1 U5520 ( .B1(n6359), .B2(n4646), .A(n4406), .ZN(n4407) );
  OAI211_X1 U5521 ( .C1(n4430), .C2(n6364), .A(n4408), .B(n4407), .ZN(U3144)
         );
  NAND2_X1 U5522 ( .A1(n4424), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4411)
         );
  OAI22_X1 U5523 ( .A1(n5790), .A2(n4426), .B1(n4425), .B2(n5795), .ZN(n4409)
         );
  AOI21_X1 U5524 ( .B1(n6334), .B2(n4646), .A(n4409), .ZN(n4410) );
  OAI211_X1 U5525 ( .C1(n4430), .C2(n6339), .A(n4411), .B(n4410), .ZN(U3142)
         );
  NAND2_X1 U5526 ( .A1(n4424), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4414)
         );
  OAI22_X1 U5527 ( .A1(n5783), .A2(n4426), .B1(n4425), .B2(n5788), .ZN(n4412)
         );
  AOI21_X1 U5528 ( .B1(n6311), .B2(n4646), .A(n4412), .ZN(n4413) );
  OAI211_X1 U5529 ( .C1(n4430), .C2(n6316), .A(n4414), .B(n4413), .ZN(U3141)
         );
  NAND2_X1 U5530 ( .A1(n4424), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4417)
         );
  OAI22_X1 U5531 ( .A1(n5827), .A2(n4426), .B1(n4425), .B2(n5833), .ZN(n4415)
         );
  AOI21_X1 U5532 ( .B1(n6378), .B2(n4646), .A(n4415), .ZN(n4416) );
  OAI211_X1 U5533 ( .C1(n4430), .C2(n6387), .A(n4417), .B(n4416), .ZN(U3147)
         );
  NAND2_X1 U5534 ( .A1(n4424), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4420)
         );
  OAI22_X1 U5535 ( .A1(n5811), .A2(n4426), .B1(n4425), .B2(n5816), .ZN(n4418)
         );
  AOI21_X1 U5536 ( .B1(n6365), .B2(n4646), .A(n4418), .ZN(n4419) );
  OAI211_X1 U5537 ( .C1(n4430), .C2(n6370), .A(n4420), .B(n4419), .ZN(U3145)
         );
  NAND2_X1 U5538 ( .A1(n4424), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4423)
         );
  OAI22_X1 U5539 ( .A1(n5776), .A2(n4426), .B1(n4425), .B2(n5781), .ZN(n4421)
         );
  AOI21_X1 U5540 ( .B1(n6353), .B2(n4646), .A(n4421), .ZN(n4422) );
  OAI211_X1 U5541 ( .C1(n6358), .C2(n4430), .A(n4423), .B(n4422), .ZN(U3140)
         );
  NAND2_X1 U5542 ( .A1(n4424), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4429)
         );
  OAI22_X1 U5543 ( .A1(n5818), .A2(n4426), .B1(n4425), .B2(n5823), .ZN(n4427)
         );
  AOI21_X1 U5544 ( .B1(n6371), .B2(n4646), .A(n4427), .ZN(n4428) );
  OAI211_X1 U5545 ( .C1(n4430), .C2(n6376), .A(n4429), .B(n4428), .ZN(U3146)
         );
  INV_X1 U5546 ( .A(n6546), .ZN(n6441) );
  NOR3_X1 U5547 ( .A1(n6540), .A2(n5725), .A3(n6441), .ZN(n6425) );
  INV_X1 U5548 ( .A(n6535), .ZN(n4431) );
  OR2_X1 U5549 ( .A1(n5210), .A2(n4431), .ZN(n6438) );
  INV_X1 U5550 ( .A(n6438), .ZN(n4432) );
  OR2_X1 U5551 ( .A1(n2997), .A2(n4432), .ZN(n4433) );
  OR2_X1 U5552 ( .A1(n6425), .A2(n4433), .ZN(n4434) );
  INV_X1 U5553 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4651) );
  NAND2_X1 U5554 ( .A1(n4726), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4764)
         );
  INV_X1 U5555 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U5556 ( .A1(n4987), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4981)
         );
  INV_X1 U5557 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U5558 ( .A1(n4957), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4942)
         );
  INV_X1 U5559 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5972) );
  INV_X1 U5560 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5575) );
  INV_X1 U5561 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5539) );
  INV_X1 U5562 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5142) );
  NAND2_X1 U5563 ( .A1(n5181), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5215)
         );
  INV_X1 U5564 ( .A(n5215), .ZN(n4439) );
  NAND2_X1 U5565 ( .A1(n4439), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4441)
         );
  INV_X1 U5566 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4440) );
  XNOR2_X1 U5567 ( .A(n4441), .B(n4440), .ZN(n5265) );
  NOR2_X1 U5568 ( .A1(n5265), .A2(n4812), .ZN(n4442) );
  AND2_X1 U5569 ( .A1(n5265), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4443) );
  INV_X1 U5570 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4451) );
  NOR2_X1 U5571 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4453) );
  NAND2_X1 U5572 ( .A1(n4444), .A2(n4453), .ZN(n6419) );
  NAND2_X1 U5573 ( .A1(n6537), .A2(n6419), .ZN(n5232) );
  NOR2_X1 U5574 ( .A1(n4453), .A2(EBX_REG_31__SCAN_IN), .ZN(n4445) );
  NAND2_X1 U5575 ( .A1(n4452), .A2(n4445), .ZN(n4446) );
  AND2_X1 U5576 ( .A1(n5232), .A2(n4446), .ZN(n4447) );
  INV_X1 U5577 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5124) );
  NOR2_X1 U5578 ( .A1(n3678), .A2(n5124), .ZN(n5226) );
  NOR2_X1 U5579 ( .A1(n4448), .A2(n4453), .ZN(n4449) );
  AOI22_X1 U5580 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6089), .B1(n6088), .B2(n6249), 
        .ZN(n4450) );
  OAI211_X1 U5581 ( .C1(n6073), .C2(n4451), .A(n4450), .B(n6238), .ZN(n4458)
         );
  INV_X1 U5582 ( .A(n6050), .ZN(n4601) );
  INV_X1 U5583 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6471) );
  INV_X1 U5584 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6652) );
  INV_X1 U5585 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6467) );
  INV_X1 U5586 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6465) );
  NOR3_X1 U5587 ( .A1(n6652), .A2(n6467), .A3(n6465), .ZN(n6082) );
  NAND2_X1 U5588 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6082), .ZN(n6067) );
  NOR2_X1 U5589 ( .A1(n6471), .A2(n6067), .ZN(n6051) );
  NAND4_X1 U5590 ( .A1(n6051), .A2(REIP_REG_8__SCAN_IN), .A3(
        REIP_REG_7__SCAN_IN), .A4(REIP_REG_6__SCAN_IN), .ZN(n4744) );
  AND3_X1 U5591 ( .A1(n4454), .A2(n4453), .A3(n4452), .ZN(n4455) );
  NAND2_X1 U5592 ( .A1(n6090), .A2(n6050), .ZN(n5303) );
  OAI21_X1 U5593 ( .B1(n4601), .B2(n4744), .A(n5303), .ZN(n6036) );
  INV_X1 U5594 ( .A(n6051), .ZN(n4456) );
  NOR2_X1 U5595 ( .A1(n6090), .A2(n4456), .ZN(n6048) );
  NAND4_X1 U5596 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .A4(n6048), .ZN(n6017) );
  INV_X1 U5597 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6477) );
  AOI22_X1 U5598 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6036), .B1(n6017), .B2(n6477), .ZN(n4457) );
  AOI211_X1 U5599 ( .C1(n4517), .C2(n6079), .A(n4458), .B(n4457), .ZN(n4459)
         );
  OAI21_X1 U5600 ( .B1(n6058), .B2(n4520), .A(n4459), .ZN(U2818) );
  NOR2_X1 U5601 ( .A1(n5765), .A2(n4465), .ZN(n4673) );
  INV_X1 U5602 ( .A(n4678), .ZN(n4672) );
  AND2_X1 U5603 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4673), .ZN(n4488)
         );
  AOI21_X1 U5604 ( .B1(n4460), .B2(n4672), .A(n4488), .ZN(n4467) );
  NAND3_X1 U5605 ( .A1(n5723), .A2(n4467), .A3(n4463), .ZN(n4461) );
  OAI211_X1 U5606 ( .C1(n4619), .C2(n4673), .A(n4462), .B(n4461), .ZN(n4487)
         );
  NAND2_X1 U5607 ( .A1(n4619), .A2(n4463), .ZN(n4466) );
  NAND2_X1 U5608 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4464) );
  OAI22_X1 U5609 ( .A1(n4467), .A2(n4466), .B1(n4465), .B2(n4464), .ZN(n4486)
         );
  AOI22_X1 U5610 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4487), .B1(n6373), 
        .B2(n4486), .ZN(n4471) );
  NOR2_X2 U5611 ( .A1(n4469), .A2(n4468), .ZN(n4707) );
  AOI22_X1 U5612 ( .A1(n6372), .A2(n4488), .B1(n5820), .B2(n4707), .ZN(n4470)
         );
  OAI211_X1 U5613 ( .C1(n5817), .C2(n4491), .A(n4471), .B(n4470), .ZN(U3130)
         );
  AOI22_X1 U5614 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4487), .B1(n6361), 
        .B2(n4486), .ZN(n4473) );
  AOI22_X1 U5615 ( .A1(n6360), .A2(n4488), .B1(n5806), .B2(n4707), .ZN(n4472)
         );
  OAI211_X1 U5616 ( .C1(n5803), .C2(n4491), .A(n4473), .B(n4472), .ZN(U3128)
         );
  AOI22_X1 U5617 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4487), .B1(n6382), 
        .B2(n4486), .ZN(n4475) );
  AOI22_X1 U5618 ( .A1(n6380), .A2(n4488), .B1(n5829), .B2(n4707), .ZN(n4474)
         );
  OAI211_X1 U5619 ( .C1(n5825), .C2(n4491), .A(n4475), .B(n4474), .ZN(U3131)
         );
  AOI22_X1 U5620 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4487), .B1(n6367), 
        .B2(n4486), .ZN(n4477) );
  AOI22_X1 U5621 ( .A1(n6366), .A2(n4488), .B1(n5813), .B2(n4707), .ZN(n4476)
         );
  OAI211_X1 U5622 ( .C1(n5810), .C2(n4491), .A(n4477), .B(n4476), .ZN(U3129)
         );
  AOI22_X1 U5623 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4487), .B1(n4478), 
        .B2(n4486), .ZN(n4481) );
  AOI22_X1 U5624 ( .A1(n4479), .A2(n4488), .B1(n5799), .B2(n4707), .ZN(n4480)
         );
  OAI211_X1 U5625 ( .C1(n5796), .C2(n4491), .A(n4481), .B(n4480), .ZN(U3127)
         );
  AOI22_X1 U5626 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4487), .B1(n6336), 
        .B2(n4486), .ZN(n4483) );
  AOI22_X1 U5627 ( .A1(n6335), .A2(n4488), .B1(n5792), .B2(n4707), .ZN(n4482)
         );
  OAI211_X1 U5628 ( .C1(n5789), .C2(n4491), .A(n4483), .B(n4482), .ZN(U3126)
         );
  AOI22_X1 U5629 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4487), .B1(n6313), 
        .B2(n4486), .ZN(n4485) );
  AOI22_X1 U5630 ( .A1(n6312), .A2(n4488), .B1(n5785), .B2(n4707), .ZN(n4484)
         );
  OAI211_X1 U5631 ( .C1(n5782), .C2(n4491), .A(n4485), .B(n4484), .ZN(U3125)
         );
  AOI22_X1 U5632 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4487), .B1(n6355), 
        .B2(n4486), .ZN(n4490) );
  AOI22_X1 U5633 ( .A1(n6354), .A2(n4488), .B1(n5778), .B2(n4707), .ZN(n4489)
         );
  OAI211_X1 U5634 ( .C1(n5775), .C2(n4491), .A(n4490), .B(n4489), .ZN(U3124)
         );
  AOI22_X1 U5635 ( .A1(n5185), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5187), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4495) );
  AOI22_X1 U5636 ( .A1(n2999), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5024), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4494) );
  AOI22_X1 U5637 ( .A1(n5197), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4493) );
  AOI22_X1 U5638 ( .A1(n5195), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4492) );
  NAND4_X1 U5639 ( .A1(n4495), .A2(n4494), .A3(n4493), .A4(n4492), .ZN(n4501)
         );
  AOI22_X1 U5640 ( .A1(n5198), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4499) );
  AOI22_X1 U5641 ( .A1(n5167), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n5189), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4498) );
  AOI22_X1 U5642 ( .A1(n5186), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4497) );
  AOI22_X1 U5643 ( .A1(n5194), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4496) );
  NAND4_X1 U5644 ( .A1(n4499), .A2(n4498), .A3(n4497), .A4(n4496), .ZN(n4500)
         );
  OAI21_X1 U5645 ( .B1(n4501), .B2(n4500), .A(n4998), .ZN(n4505) );
  XNOR2_X1 U5646 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n4502), .ZN(n4577)
         );
  AOI22_X1 U5647 ( .A1(n5216), .A2(n4577), .B1(n5219), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4504) );
  NAND2_X1 U5648 ( .A1(n5158), .A2(EAX_REG_10__SCAN_IN), .ZN(n4503) );
  AND3_X1 U5649 ( .A1(n4505), .A2(n4504), .A3(n4503), .ZN(n4507) );
  AOI21_X1 U5650 ( .B1(n4507), .B2(n4506), .A(n4666), .ZN(n4579) );
  OR2_X1 U5651 ( .A1(n4509), .A2(n4508), .ZN(n4510) );
  NAND2_X1 U5652 ( .A1(n6015), .A2(n4510), .ZN(n6239) );
  OAI22_X1 U5653 ( .A1(n6239), .A2(n6103), .B1(n4511), .B2(n5486), .ZN(n4512)
         );
  AOI21_X1 U5654 ( .B1(n4579), .B2(n6108), .A(n4512), .ZN(n4513) );
  INV_X1 U5655 ( .A(n4513), .ZN(U2849) );
  XNOR2_X1 U5656 ( .A(n2996), .B(n6254), .ZN(n4515) );
  XNOR2_X1 U5657 ( .A(n4569), .B(n4515), .ZN(n6250) );
  INV_X1 U5658 ( .A(n6195), .ZN(n6221) );
  NAND2_X1 U5659 ( .A1(n6250), .A2(n6221), .ZN(n4519) );
  NAND2_X1 U5660 ( .A1(n2997), .A2(REIP_REG_9__SCAN_IN), .ZN(n6247) );
  OAI21_X1 U5661 ( .B1(n6208), .B2(n4451), .A(n6247), .ZN(n4516) );
  AOI21_X1 U5662 ( .B1(n6204), .B2(n4517), .A(n4516), .ZN(n4518) );
  OAI211_X1 U5663 ( .C1(n6194), .C2(n4520), .A(n4519), .B(n4518), .ZN(U2977)
         );
  INV_X1 U5664 ( .A(n4579), .ZN(n4567) );
  AOI22_X1 U5665 ( .A1(n5511), .A2(DATAI_10_), .B1(n6122), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n4521) );
  OAI21_X1 U5666 ( .B1(n4567), .B2(n5863), .A(n4521), .ZN(U2881) );
  NOR2_X1 U5667 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4522), .ZN(n4529)
         );
  OAI21_X1 U5668 ( .B1(n4524), .B2(n4557), .A(n4523), .ZN(n4526) );
  INV_X1 U5669 ( .A(n4531), .ZN(n4525) );
  AOI21_X1 U5670 ( .B1(n4526), .B2(n4525), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4528) );
  NOR2_X1 U5671 ( .A1(n5728), .A2(n4527), .ZN(n5774) );
  OAI21_X1 U5672 ( .B1(n4529), .B2(n4528), .A(n5774), .ZN(n4553) );
  NAND2_X1 U5673 ( .A1(n4553), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4534) );
  INV_X1 U5674 ( .A(n4529), .ZN(n4555) );
  NOR2_X1 U5675 ( .A1(n5766), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4530)
         );
  AOI22_X1 U5676 ( .A1(n4531), .A2(n4619), .B1(n5768), .B2(n4530), .ZN(n4554)
         );
  OAI22_X1 U5677 ( .A1(n5818), .A2(n4555), .B1(n4554), .B2(n5823), .ZN(n4532)
         );
  AOI21_X1 U5678 ( .B1(n6371), .B2(n4557), .A(n4532), .ZN(n4533) );
  OAI211_X1 U5679 ( .C1(n4560), .C2(n6376), .A(n4534), .B(n4533), .ZN(U3042)
         );
  NAND2_X1 U5680 ( .A1(n4553), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4537) );
  OAI22_X1 U5681 ( .A1(n5827), .A2(n4555), .B1(n4554), .B2(n5833), .ZN(n4535)
         );
  AOI21_X1 U5682 ( .B1(n6378), .B2(n4557), .A(n4535), .ZN(n4536) );
  OAI211_X1 U5683 ( .C1(n4560), .C2(n6387), .A(n4537), .B(n4536), .ZN(U3043)
         );
  NAND2_X1 U5684 ( .A1(n4553), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4540) );
  OAI22_X1 U5685 ( .A1(n5811), .A2(n4555), .B1(n4554), .B2(n5816), .ZN(n4538)
         );
  AOI21_X1 U5686 ( .B1(n6365), .B2(n4557), .A(n4538), .ZN(n4539) );
  OAI211_X1 U5687 ( .C1(n4560), .C2(n6370), .A(n4540), .B(n4539), .ZN(U3041)
         );
  NAND2_X1 U5688 ( .A1(n4553), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4543) );
  OAI22_X1 U5689 ( .A1(n5804), .A2(n4555), .B1(n4554), .B2(n5809), .ZN(n4541)
         );
  AOI21_X1 U5690 ( .B1(n6359), .B2(n4557), .A(n4541), .ZN(n4542) );
  OAI211_X1 U5691 ( .C1(n4560), .C2(n6364), .A(n4543), .B(n4542), .ZN(U3040)
         );
  NAND2_X1 U5692 ( .A1(n4553), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4546) );
  OAI22_X1 U5693 ( .A1(n5797), .A2(n4555), .B1(n4554), .B2(n5802), .ZN(n4544)
         );
  AOI21_X1 U5694 ( .B1(n5741), .B2(n4557), .A(n4544), .ZN(n4545) );
  OAI211_X1 U5695 ( .C1(n4560), .C2(n5744), .A(n4546), .B(n4545), .ZN(U3039)
         );
  NAND2_X1 U5696 ( .A1(n4553), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4549) );
  OAI22_X1 U5697 ( .A1(n5783), .A2(n4555), .B1(n4554), .B2(n5788), .ZN(n4547)
         );
  AOI21_X1 U5698 ( .B1(n6311), .B2(n4557), .A(n4547), .ZN(n4548) );
  OAI211_X1 U5699 ( .C1(n4560), .C2(n6316), .A(n4549), .B(n4548), .ZN(U3037)
         );
  NAND2_X1 U5700 ( .A1(n4553), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4552) );
  OAI22_X1 U5701 ( .A1(n5790), .A2(n4555), .B1(n4554), .B2(n5795), .ZN(n4550)
         );
  AOI21_X1 U5702 ( .B1(n6334), .B2(n4557), .A(n4550), .ZN(n4551) );
  OAI211_X1 U5703 ( .C1(n4560), .C2(n6339), .A(n4552), .B(n4551), .ZN(U3038)
         );
  NAND2_X1 U5704 ( .A1(n4553), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4559) );
  OAI22_X1 U5705 ( .A1(n5776), .A2(n4555), .B1(n4554), .B2(n5781), .ZN(n4556)
         );
  AOI21_X1 U5706 ( .B1(n6353), .B2(n4557), .A(n4556), .ZN(n4558) );
  OAI211_X1 U5707 ( .C1(n6358), .C2(n4560), .A(n4559), .B(n4558), .ZN(U3036)
         );
  INV_X1 U5708 ( .A(n4577), .ZN(n4565) );
  AOI22_X1 U5709 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6089), .B1(
        PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n6091), .ZN(n4561) );
  OAI211_X1 U5710 ( .C1(n6065), .C2(n6239), .A(n4561), .B(n6238), .ZN(n4564)
         );
  INV_X1 U5711 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6479) );
  NAND2_X1 U5712 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n6018) );
  OAI21_X1 U5713 ( .B1(REIP_REG_10__SCAN_IN), .B2(REIP_REG_9__SCAN_IN), .A(
        n6018), .ZN(n4562) );
  OAI22_X1 U5714 ( .A1(n6479), .A2(n6036), .B1(n6017), .B2(n4562), .ZN(n4563)
         );
  AOI211_X1 U5715 ( .C1(n6079), .C2(n4565), .A(n4564), .B(n4563), .ZN(n4566)
         );
  OAI21_X1 U5716 ( .B1(n6058), .B2(n4567), .A(n4566), .ZN(U2817) );
  OR2_X1 U5717 ( .A1(n4569), .A2(n4568), .ZN(n4571) );
  NAND2_X1 U5718 ( .A1(n4571), .A2(n4570), .ZN(n4575) );
  NAND2_X1 U5719 ( .A1(n4573), .A2(n4572), .ZN(n4574) );
  XNOR2_X1 U5720 ( .A(n4575), .B(n4574), .ZN(n6237) );
  AOI22_X1 U5721 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n2997), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n4576) );
  OAI21_X1 U5722 ( .B1(n4577), .B2(n6225), .A(n4576), .ZN(n4578) );
  AOI21_X1 U5723 ( .B1(n4579), .B2(n6219), .A(n4578), .ZN(n4580) );
  OAI21_X1 U5724 ( .B1(n6195), .B2(n6237), .A(n4580), .ZN(U2976) );
  NAND2_X1 U5725 ( .A1(n6533), .A2(n4581), .ZN(n6095) );
  NAND2_X1 U5726 ( .A1(n6533), .A2(n4582), .ZN(n4583) );
  NAND2_X1 U5727 ( .A1(n4583), .A2(n6058), .ZN(n6098) );
  NAND2_X1 U5728 ( .A1(n6109), .A2(n6098), .ZN(n4600) );
  OR2_X1 U5729 ( .A1(n6090), .A2(n6082), .ZN(n4584) );
  NAND2_X1 U5730 ( .A1(n4584), .A2(n6050), .ZN(n6077) );
  NAND2_X1 U5731 ( .A1(n6050), .A2(REIP_REG_1__SCAN_IN), .ZN(n4585) );
  NAND2_X1 U5732 ( .A1(n5303), .A2(n4585), .ZN(n4586) );
  NAND2_X1 U5733 ( .A1(n4586), .A2(REIP_REG_2__SCAN_IN), .ZN(n6093) );
  NAND2_X1 U5734 ( .A1(n6093), .A2(n6467), .ZN(n4598) );
  INV_X1 U5735 ( .A(n4587), .ZN(n4590) );
  AOI21_X1 U5736 ( .B1(n4590), .B2(n4589), .A(n4588), .ZN(n4591) );
  NAND2_X1 U5737 ( .A1(n6088), .A2(n3008), .ZN(n4596) );
  INV_X1 U5738 ( .A(n4592), .ZN(n4593) );
  AOI22_X1 U5739 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n6091), .B1(n6079), 
        .B2(n4593), .ZN(n4595) );
  NAND2_X1 U5740 ( .A1(n6089), .A2(EBX_REG_3__SCAN_IN), .ZN(n4594) );
  NAND3_X1 U5741 ( .A1(n4596), .A2(n4595), .A3(n4594), .ZN(n4597) );
  AOI21_X1 U5742 ( .B1(n6077), .B2(n4598), .A(n4597), .ZN(n4599) );
  OAI211_X1 U5743 ( .C1(n5729), .C2(n6095), .A(n4600), .B(n4599), .ZN(U2824)
         );
  NAND2_X1 U5744 ( .A1(n6220), .A2(n6098), .ZN(n4608) );
  NOR2_X1 U5745 ( .A1(n6090), .A2(REIP_REG_1__SCAN_IN), .ZN(n4606) );
  INV_X1 U5746 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4604) );
  AOI22_X1 U5747 ( .A1(EBX_REG_1__SCAN_IN), .A2(n6089), .B1(n4601), .B2(
        REIP_REG_1__SCAN_IN), .ZN(n4603) );
  NAND2_X1 U5748 ( .A1(n6079), .A2(n4604), .ZN(n4602) );
  OAI211_X1 U5749 ( .C1(n6073), .C2(n4604), .A(n4603), .B(n4602), .ZN(n4605)
         );
  AOI211_X1 U5750 ( .C1(n6088), .C2(n3799), .A(n4606), .B(n4605), .ZN(n4607)
         );
  OAI211_X1 U5751 ( .C1(n6095), .C2(n4609), .A(n4608), .B(n4607), .ZN(U2826)
         );
  OR2_X1 U5752 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4610), .ZN(n4644)
         );
  INV_X1 U5753 ( .A(n4611), .ZN(n4612) );
  NOR2_X1 U5754 ( .A1(n5768), .A2(n4612), .ZN(n5727) );
  OAI21_X1 U5755 ( .B1(n5727), .B2(n6532), .A(n4613), .ZN(n5720) );
  AOI211_X1 U5756 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4644), .A(n5728), .B(
        n5720), .ZN(n4618) );
  INV_X1 U5757 ( .A(n4649), .ZN(n4614) );
  OAI21_X1 U5758 ( .B1(n4646), .B2(n4614), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4616) );
  NAND3_X1 U5759 ( .A1(n4616), .A2(n5723), .A3(n4615), .ZN(n4617) );
  NAND2_X1 U5760 ( .A1(n4618), .A2(n4617), .ZN(n4642) );
  NAND2_X1 U5761 ( .A1(n4642), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4623) );
  AOI22_X1 U5762 ( .A1(n4620), .A2(n4619), .B1(n5721), .B2(n5727), .ZN(n4643)
         );
  OAI22_X1 U5763 ( .A1(n5804), .A2(n4644), .B1(n4643), .B2(n5809), .ZN(n4621)
         );
  AOI21_X1 U5764 ( .B1(n5806), .B2(n4646), .A(n4621), .ZN(n4622) );
  OAI211_X1 U5765 ( .C1(n4649), .C2(n5803), .A(n4623), .B(n4622), .ZN(U3024)
         );
  NAND2_X1 U5766 ( .A1(n4642), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4626) );
  OAI22_X1 U5767 ( .A1(n5818), .A2(n4644), .B1(n4643), .B2(n5823), .ZN(n4624)
         );
  AOI21_X1 U5768 ( .B1(n5820), .B2(n4646), .A(n4624), .ZN(n4625) );
  OAI211_X1 U5769 ( .C1(n4649), .C2(n5817), .A(n4626), .B(n4625), .ZN(U3026)
         );
  NAND2_X1 U5770 ( .A1(n4642), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4629) );
  OAI22_X1 U5771 ( .A1(n5811), .A2(n4644), .B1(n4643), .B2(n5816), .ZN(n4627)
         );
  AOI21_X1 U5772 ( .B1(n5813), .B2(n4646), .A(n4627), .ZN(n4628) );
  OAI211_X1 U5773 ( .C1(n4649), .C2(n5810), .A(n4629), .B(n4628), .ZN(U3025)
         );
  NAND2_X1 U5774 ( .A1(n4642), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4632) );
  OAI22_X1 U5775 ( .A1(n5827), .A2(n4644), .B1(n4643), .B2(n5833), .ZN(n4630)
         );
  AOI21_X1 U5776 ( .B1(n5829), .B2(n4646), .A(n4630), .ZN(n4631) );
  OAI211_X1 U5777 ( .C1(n4649), .C2(n5825), .A(n4632), .B(n4631), .ZN(U3027)
         );
  NAND2_X1 U5778 ( .A1(n4642), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4635) );
  OAI22_X1 U5779 ( .A1(n5797), .A2(n4644), .B1(n4643), .B2(n5802), .ZN(n4633)
         );
  AOI21_X1 U5780 ( .B1(n5799), .B2(n4646), .A(n4633), .ZN(n4634) );
  OAI211_X1 U5781 ( .C1(n4649), .C2(n5796), .A(n4635), .B(n4634), .ZN(U3023)
         );
  NAND2_X1 U5782 ( .A1(n4642), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4638) );
  OAI22_X1 U5783 ( .A1(n5776), .A2(n4644), .B1(n4643), .B2(n5781), .ZN(n4636)
         );
  AOI21_X1 U5784 ( .B1(n5778), .B2(n4646), .A(n4636), .ZN(n4637) );
  OAI211_X1 U5785 ( .C1(n4649), .C2(n5775), .A(n4638), .B(n4637), .ZN(U3020)
         );
  NAND2_X1 U5786 ( .A1(n4642), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4641) );
  OAI22_X1 U5787 ( .A1(n5783), .A2(n4644), .B1(n4643), .B2(n5788), .ZN(n4639)
         );
  AOI21_X1 U5788 ( .B1(n5785), .B2(n4646), .A(n4639), .ZN(n4640) );
  OAI211_X1 U5789 ( .C1(n4649), .C2(n5782), .A(n4641), .B(n4640), .ZN(U3021)
         );
  NAND2_X1 U5790 ( .A1(n4642), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4648) );
  OAI22_X1 U5791 ( .A1(n5790), .A2(n4644), .B1(n4643), .B2(n5795), .ZN(n4645)
         );
  AOI21_X1 U5792 ( .B1(n5792), .B2(n4646), .A(n4645), .ZN(n4647) );
  OAI211_X1 U5793 ( .C1(n4649), .C2(n5789), .A(n4648), .B(n4647), .ZN(U3022)
         );
  XOR2_X1 U5794 ( .A(n4651), .B(n4650), .Z(n6023) );
  AOI22_X1 U5795 ( .A1(n5198), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5167), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4655) );
  AOI22_X1 U5796 ( .A1(n5197), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5024), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4654) );
  AOI22_X1 U5797 ( .A1(n5185), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4653) );
  AOI22_X1 U5798 ( .A1(n5187), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4652) );
  NAND4_X1 U5799 ( .A1(n4655), .A2(n4654), .A3(n4653), .A4(n4652), .ZN(n4661)
         );
  AOI22_X1 U5800 ( .A1(n5195), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5189), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4659) );
  AOI22_X1 U5801 ( .A1(n5194), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4658) );
  AOI22_X1 U5802 ( .A1(n2998), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4657) );
  AOI22_X1 U5803 ( .A1(n2999), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4656) );
  NAND4_X1 U5804 ( .A1(n4659), .A2(n4658), .A3(n4657), .A4(n4656), .ZN(n4660)
         );
  OR2_X1 U5805 ( .A1(n4661), .A2(n4660), .ZN(n4662) );
  AOI22_X1 U5806 ( .A1(n4998), .A2(n4662), .B1(n5219), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4664) );
  NAND2_X1 U5807 ( .A1(n5158), .A2(EAX_REG_11__SCAN_IN), .ZN(n4663) );
  OAI211_X1 U5808 ( .C1(n6023), .C2(n5210), .A(n4664), .B(n4663), .ZN(n4665)
         );
  NOR2_X1 U5809 ( .A1(n4666), .A2(n4665), .ZN(n4667) );
  OR2_X1 U5810 ( .A1(n4763), .A2(n4667), .ZN(n6189) );
  AOI22_X1 U5811 ( .A1(n5511), .A2(DATAI_11_), .B1(n6122), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n4668) );
  OAI21_X1 U5812 ( .B1(n6189), .B2(n5863), .A(n4668), .ZN(U2880) );
  INV_X1 U5813 ( .A(n4707), .ZN(n4669) );
  AOI21_X1 U5814 ( .B1(n4669), .B2(n6352), .A(n6538), .ZN(n4670) );
  AOI211_X1 U5815 ( .C1(n4672), .C2(n4671), .A(n5763), .B(n4670), .ZN(n4676)
         );
  AND2_X1 U5816 ( .A1(n6388), .A2(n4673), .ZN(n4677) );
  OAI211_X1 U5817 ( .C1(n5725), .C2(n4677), .A(n5766), .B(n4674), .ZN(n4675)
         );
  NAND2_X1 U5818 ( .A1(n4703), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4684)
         );
  INV_X1 U5819 ( .A(n4677), .ZN(n4705) );
  NOR2_X1 U5820 ( .A1(n4678), .A2(n5763), .ZN(n5730) );
  INV_X1 U5821 ( .A(n4679), .ZN(n4680) );
  AOI22_X1 U5822 ( .A1(n5730), .A2(n4681), .B1(n4680), .B2(n5728), .ZN(n4704)
         );
  OAI22_X1 U5823 ( .A1(n5811), .A2(n4705), .B1(n4704), .B2(n5816), .ZN(n4682)
         );
  AOI21_X1 U5824 ( .B1(n6365), .B2(n4707), .A(n4682), .ZN(n4683) );
  OAI211_X1 U5825 ( .C1(n6352), .C2(n6370), .A(n4684), .B(n4683), .ZN(U3121)
         );
  NAND2_X1 U5826 ( .A1(n4703), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4687)
         );
  OAI22_X1 U5827 ( .A1(n5827), .A2(n4705), .B1(n4704), .B2(n5833), .ZN(n4685)
         );
  AOI21_X1 U5828 ( .B1(n6378), .B2(n4707), .A(n4685), .ZN(n4686) );
  OAI211_X1 U5829 ( .C1(n6352), .C2(n6387), .A(n4687), .B(n4686), .ZN(U3123)
         );
  NAND2_X1 U5830 ( .A1(n4703), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4690)
         );
  OAI22_X1 U5831 ( .A1(n5804), .A2(n4705), .B1(n4704), .B2(n5809), .ZN(n4688)
         );
  AOI21_X1 U5832 ( .B1(n6359), .B2(n4707), .A(n4688), .ZN(n4689) );
  OAI211_X1 U5833 ( .C1(n6352), .C2(n6364), .A(n4690), .B(n4689), .ZN(U3120)
         );
  NAND2_X1 U5834 ( .A1(n4703), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4693)
         );
  OAI22_X1 U5835 ( .A1(n5776), .A2(n4705), .B1(n4704), .B2(n5781), .ZN(n4691)
         );
  AOI21_X1 U5836 ( .B1(n6353), .B2(n4707), .A(n4691), .ZN(n4692) );
  OAI211_X1 U5837 ( .C1(n6352), .C2(n6358), .A(n4693), .B(n4692), .ZN(U3116)
         );
  NAND2_X1 U5838 ( .A1(n4703), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4696)
         );
  OAI22_X1 U5839 ( .A1(n5790), .A2(n4705), .B1(n4704), .B2(n5795), .ZN(n4694)
         );
  AOI21_X1 U5840 ( .B1(n6334), .B2(n4707), .A(n4694), .ZN(n4695) );
  OAI211_X1 U5841 ( .C1(n6352), .C2(n6339), .A(n4696), .B(n4695), .ZN(U3118)
         );
  NAND2_X1 U5842 ( .A1(n4703), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4699)
         );
  OAI22_X1 U5843 ( .A1(n5797), .A2(n4705), .B1(n4704), .B2(n5802), .ZN(n4697)
         );
  AOI21_X1 U5844 ( .B1(n5741), .B2(n4707), .A(n4697), .ZN(n4698) );
  OAI211_X1 U5845 ( .C1(n6352), .C2(n5744), .A(n4699), .B(n4698), .ZN(U3119)
         );
  NAND2_X1 U5846 ( .A1(n4703), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4702)
         );
  OAI22_X1 U5847 ( .A1(n5818), .A2(n4705), .B1(n4704), .B2(n5823), .ZN(n4700)
         );
  AOI21_X1 U5848 ( .B1(n6371), .B2(n4707), .A(n4700), .ZN(n4701) );
  OAI211_X1 U5849 ( .C1(n6352), .C2(n6376), .A(n4702), .B(n4701), .ZN(U3122)
         );
  NAND2_X1 U5850 ( .A1(n4703), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4709)
         );
  OAI22_X1 U5851 ( .A1(n5783), .A2(n4705), .B1(n4704), .B2(n5788), .ZN(n4706)
         );
  AOI21_X1 U5852 ( .B1(n6311), .B2(n4707), .A(n4706), .ZN(n4708) );
  OAI211_X1 U5853 ( .C1(n6352), .C2(n6316), .A(n4709), .B(n4708), .ZN(U3117)
         );
  NAND2_X1 U5854 ( .A1(n4711), .A2(n6185), .ZN(n5881) );
  XNOR2_X1 U5855 ( .A(n2996), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4712)
         );
  XNOR2_X1 U5856 ( .A(n5881), .B(n4712), .ZN(n4761) );
  INV_X1 U5857 ( .A(n4713), .ZN(n4714) );
  OAI22_X1 U5858 ( .A1(n4715), .A2(n6235), .B1(n6236), .B2(n4714), .ZN(n6233)
         );
  OAI21_X1 U5859 ( .B1(n4717), .B2(n4716), .A(n6234), .ZN(n4718) );
  AOI21_X1 U5860 ( .B1(n6233), .B2(n4718), .A(n6714), .ZN(n4724) );
  NAND2_X1 U5861 ( .A1(n2997), .A2(REIP_REG_12__SCAN_IN), .ZN(n4756) );
  INV_X1 U5862 ( .A(n4756), .ZN(n4723) );
  AND2_X1 U5863 ( .A1(n3005), .A2(n4719), .ZN(n4720) );
  OR2_X1 U5864 ( .A1(n4720), .A2(n4787), .ZN(n4745) );
  NOR2_X1 U5865 ( .A1(n4745), .A2(n6303), .ZN(n4722) );
  NOR3_X1 U5866 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6226), .A3(n6234), 
        .ZN(n4721) );
  NOR4_X1 U5867 ( .A1(n4724), .A2(n4723), .A3(n4722), .A4(n4721), .ZN(n4725)
         );
  OAI21_X1 U5868 ( .B1(n4761), .B2(n6269), .A(n4725), .ZN(U3006) );
  AOI22_X1 U5869 ( .A1(n5158), .A2(EAX_REG_12__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6532), .ZN(n4739) );
  XNOR2_X1 U5870 ( .A(n4726), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4757)
         );
  NAND2_X1 U5871 ( .A1(n4757), .A2(n5216), .ZN(n4738) );
  AOI22_X1 U5872 ( .A1(n5185), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4730) );
  AOI22_X1 U5873 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n5167), .B1(n5198), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4729) );
  AOI22_X1 U5874 ( .A1(n5197), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4728) );
  AOI22_X1 U5875 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n3000), .B1(n5029), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4727) );
  NAND4_X1 U5876 ( .A1(n4730), .A2(n4729), .A3(n4728), .A4(n4727), .ZN(n4736)
         );
  AOI22_X1 U5877 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n2999), .B1(n5024), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4734) );
  AOI22_X1 U5878 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5195), .B1(n5189), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4733) );
  AOI22_X1 U5879 ( .A1(n5187), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4732) );
  AOI22_X1 U5880 ( .A1(n5186), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4731) );
  NAND4_X1 U5881 ( .A1(n4734), .A2(n4733), .A3(n4732), .A4(n4731), .ZN(n4735)
         );
  OAI21_X1 U5882 ( .B1(n4736), .B2(n4735), .A(n4998), .ZN(n4737) );
  OAI211_X1 U5883 ( .C1(n5216), .C2(n4739), .A(n4738), .B(n4737), .ZN(n4762)
         );
  XOR2_X1 U5884 ( .A(n4762), .B(n4763), .Z(n4759) );
  INV_X1 U5885 ( .A(n4759), .ZN(n4741) );
  AOI22_X1 U5886 ( .A1(n5511), .A2(DATAI_12_), .B1(n6122), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n4740) );
  OAI21_X1 U5887 ( .B1(n4741), .B2(n5863), .A(n4740), .ZN(U2879) );
  OAI22_X1 U5888 ( .A1(n4745), .A2(n6103), .B1(n6684), .B2(n5486), .ZN(n4742)
         );
  AOI21_X1 U5889 ( .B1(n4759), .B2(n6108), .A(n4742), .ZN(n4743) );
  INV_X1 U5890 ( .A(n4743), .ZN(U2847) );
  NAND3_X1 U5891 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .ZN(n4752) );
  NOR2_X1 U5892 ( .A1(n4744), .A2(n4752), .ZN(n5090) );
  OAI21_X1 U5893 ( .B1(n6090), .B2(n5090), .A(n6050), .ZN(n6019) );
  INV_X1 U5894 ( .A(n6019), .ZN(n4751) );
  INV_X1 U5895 ( .A(REIP_REG_12__SCAN_IN), .ZN(n4750) );
  INV_X1 U5896 ( .A(n4757), .ZN(n4747) );
  NOR2_X1 U5897 ( .A1(n6065), .A2(n4745), .ZN(n4746) );
  AOI211_X1 U5898 ( .C1(n6079), .C2(n4747), .A(n4746), .B(n2997), .ZN(n4749)
         );
  AOI22_X1 U5899 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6089), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6091), .ZN(n4748) );
  OAI211_X1 U5900 ( .C1(n4751), .C2(n4750), .A(n4749), .B(n4748), .ZN(n4753)
         );
  NOR3_X1 U5901 ( .A1(REIP_REG_12__SCAN_IN), .A2(n4752), .A3(n6017), .ZN(n6004) );
  AOI211_X1 U5902 ( .C1(n6032), .C2(n4759), .A(n4753), .B(n6004), .ZN(n4754)
         );
  INV_X1 U5903 ( .A(n4754), .ZN(U2815) );
  NAND2_X1 U5904 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4755)
         );
  OAI211_X1 U5905 ( .C1(n6225), .C2(n4757), .A(n4756), .B(n4755), .ZN(n4758)
         );
  AOI21_X1 U5906 ( .B1(n4759), .B2(n6219), .A(n4758), .ZN(n4760) );
  OAI21_X1 U5907 ( .B1(n4761), .B2(n6195), .A(n4760), .ZN(U2974) );
  INV_X1 U5908 ( .A(n4764), .ZN(n4766) );
  INV_X1 U5909 ( .A(n4987), .ZN(n4765) );
  OAI21_X1 U5910 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n4766), .A(n4765), 
        .ZN(n6009) );
  NAND2_X1 U5911 ( .A1(n5216), .A2(n6009), .ZN(n4767) );
  OAI21_X1 U5912 ( .B1(n4768), .B2(n6006), .A(n4767), .ZN(n4769) );
  AOI21_X1 U5913 ( .B1(n5220), .B2(EAX_REG_13__SCAN_IN), .A(n4769), .ZN(n4770)
         );
  OR2_X2 U5914 ( .A1(n4771), .A2(n4770), .ZN(n4889) );
  NAND2_X1 U5915 ( .A1(n4771), .A2(n4770), .ZN(n4772) );
  AOI22_X1 U5916 ( .A1(n2998), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n5167), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4776) );
  AOI22_X1 U5917 ( .A1(n5189), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4775) );
  AOI22_X1 U5918 ( .A1(n2999), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4774) );
  AOI22_X1 U5919 ( .A1(n5185), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4773) );
  NAND4_X1 U5920 ( .A1(n4776), .A2(n4775), .A3(n4774), .A4(n4773), .ZN(n4782)
         );
  AOI22_X1 U5921 ( .A1(n5197), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5195), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4780) );
  AOI22_X1 U5922 ( .A1(n5187), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4779) );
  AOI22_X1 U5923 ( .A1(n5196), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5188), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4778) );
  AOI22_X1 U5924 ( .A1(n5198), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4777) );
  NAND4_X1 U5925 ( .A1(n4780), .A2(n4779), .A3(n4778), .A4(n4777), .ZN(n4781)
         );
  OR2_X1 U5926 ( .A1(n4782), .A2(n4781), .ZN(n4783) );
  AND2_X1 U5927 ( .A1(n4998), .A2(n4783), .ZN(n4784) );
  OAI21_X1 U5928 ( .B1(n4785), .B2(n4784), .A(n4890), .ZN(n6128) );
  INV_X1 U5929 ( .A(EBX_REG_13__SCAN_IN), .ZN(n4789) );
  INV_X1 U5930 ( .A(n5483), .ZN(n4786) );
  OAI21_X1 U5931 ( .B1(n4788), .B2(n4787), .A(n4786), .ZN(n6013) );
  OAI222_X1 U5932 ( .A1(n6128), .A2(n5466), .B1(n5486), .B2(n4789), .C1(n6103), 
        .C2(n6013), .ZN(U2846) );
  NAND2_X1 U5933 ( .A1(n5525), .A2(n4791), .ZN(n5276) );
  AOI21_X1 U5934 ( .B1(n5278), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n4792), 
        .ZN(n4793) );
  XNOR2_X1 U5935 ( .A(n4793), .B(n4808), .ZN(n5524) );
  INV_X1 U5936 ( .A(n5324), .ZN(n4794) );
  NAND2_X1 U5937 ( .A1(n4801), .A2(n4794), .ZN(n4795) );
  NAND2_X1 U5938 ( .A1(n4795), .A2(n4798), .ZN(n4796) );
  OR2_X1 U5939 ( .A1(n4797), .A2(n4796), .ZN(n4803) );
  INV_X1 U5940 ( .A(n4798), .ZN(n4800) );
  NAND2_X1 U5941 ( .A1(n5324), .A2(n5439), .ZN(n4799) );
  NAND3_X1 U5942 ( .A1(n4801), .A2(n4800), .A3(n4799), .ZN(n4802) );
  NAND2_X1 U5943 ( .A1(n4803), .A2(n4802), .ZN(n5400) );
  INV_X1 U5944 ( .A(n5400), .ZN(n4804) );
  NAND2_X1 U5945 ( .A1(n2997), .A2(REIP_REG_30__SCAN_IN), .ZN(n5518) );
  OAI21_X1 U5946 ( .B1(n4804), .B2(n6303), .A(n5518), .ZN(n4807) );
  NOR3_X1 U5947 ( .A1(n5631), .A2(n4805), .A3(n4808), .ZN(n4806) );
  AOI211_X1 U5948 ( .C1(n4809), .C2(n4808), .A(n4807), .B(n4806), .ZN(n4810)
         );
  OAI21_X1 U5949 ( .B1(n5524), .B2(n6269), .A(n4810), .ZN(U2988) );
  NOR3_X1 U5950 ( .A1(n4812), .A2(n6309), .A3(n4811), .ZN(n4814) );
  NOR3_X1 U5951 ( .A1(n6423), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n4816), 
        .ZN(n4813) );
  AOI211_X1 U5952 ( .C1(n4815), .C2(n5936), .A(n4814), .B(n4813), .ZN(n4820)
         );
  AOI21_X1 U5953 ( .B1(n4817), .B2(n4816), .A(n4819), .ZN(n4818) );
  OAI22_X1 U5954 ( .A1(n4820), .A2(n4819), .B1(n4818), .B2(n3997), .ZN(U3459)
         );
  XNOR2_X1 U5955 ( .A(n2996), .B(n6567), .ZN(n4821) );
  XNOR2_X1 U5956 ( .A(n5525), .B(n4821), .ZN(n5085) );
  NOR2_X1 U5957 ( .A1(n5371), .A2(n4823), .ZN(n4824) );
  OR2_X1 U5958 ( .A1(n4822), .A2(n4824), .ZN(n5405) );
  NAND2_X1 U5959 ( .A1(n2997), .A2(REIP_REG_26__SCAN_IN), .ZN(n5081) );
  OAI21_X1 U5960 ( .B1(n5405), .B2(n6303), .A(n5081), .ZN(n4828) );
  INV_X1 U5961 ( .A(n5662), .ZN(n4826) );
  NOR2_X1 U5962 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5527) );
  NOR3_X1 U5963 ( .A1(n4826), .A2(n4825), .A3(n5527), .ZN(n4827) );
  AOI211_X1 U5964 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n4829), .A(n4828), .B(n4827), .ZN(n4830) );
  OAI21_X1 U5965 ( .B1(n5085), .B2(n6269), .A(n4830), .ZN(U2992) );
  INV_X1 U5966 ( .A(n4831), .ZN(n4832) );
  INV_X1 U5967 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U5968 ( .A1(n4832), .A2(n5349), .ZN(n4833) );
  NAND2_X1 U5969 ( .A1(n5139), .A2(n4833), .ZN(n5348) );
  AOI22_X1 U5970 ( .A1(n5198), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4837) );
  AOI22_X1 U5971 ( .A1(n5185), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4836) );
  AOI22_X1 U5972 ( .A1(n5187), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4835) );
  AOI22_X1 U5973 ( .A1(n5167), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4834) );
  NAND4_X1 U5974 ( .A1(n4837), .A2(n4836), .A3(n4835), .A4(n4834), .ZN(n4843)
         );
  AOI22_X1 U5975 ( .A1(n5195), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5189), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4841) );
  AOI22_X1 U5976 ( .A1(n5197), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4840) );
  AOI22_X1 U5977 ( .A1(n2999), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4839) );
  AOI22_X1 U5978 ( .A1(n5024), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4838) );
  NAND4_X1 U5979 ( .A1(n4841), .A2(n4840), .A3(n4839), .A4(n4838), .ZN(n4842)
         );
  NOR2_X1 U5980 ( .A1(n4843), .A2(n4842), .ZN(n5069) );
  AOI22_X1 U5981 ( .A1(n5198), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5189), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4847) );
  AOI22_X1 U5982 ( .A1(n5194), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4846) );
  AOI22_X1 U5983 ( .A1(n5185), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4845) );
  AOI22_X1 U5984 ( .A1(n2999), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4844) );
  NAND4_X1 U5985 ( .A1(n4847), .A2(n4846), .A3(n4845), .A4(n4844), .ZN(n4853)
         );
  AOI22_X1 U5986 ( .A1(n2998), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5167), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4851) );
  AOI22_X1 U5987 ( .A1(n5197), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5024), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4850) );
  AOI22_X1 U5988 ( .A1(n5187), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4849) );
  AOI22_X1 U5989 ( .A1(n5195), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4848) );
  NAND4_X1 U5990 ( .A1(n4851), .A2(n4850), .A3(n4849), .A4(n4848), .ZN(n4852)
         );
  NOR2_X1 U5991 ( .A1(n4853), .A2(n4852), .ZN(n5047) );
  AOI22_X1 U5992 ( .A1(n5198), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5167), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4857) );
  AOI22_X1 U5993 ( .A1(n5185), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4856) );
  AOI22_X1 U5994 ( .A1(n2999), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4855) );
  AOI22_X1 U5995 ( .A1(n5189), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4854) );
  NAND4_X1 U5996 ( .A1(n4857), .A2(n4856), .A3(n4855), .A4(n4854), .ZN(n4863)
         );
  AOI22_X1 U5997 ( .A1(n2998), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5195), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4861) );
  AOI22_X1 U5998 ( .A1(n5197), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4860) );
  AOI22_X1 U5999 ( .A1(n5024), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4859) );
  AOI22_X1 U6000 ( .A1(n5187), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4858) );
  NAND4_X1 U6001 ( .A1(n4861), .A2(n4860), .A3(n4859), .A4(n4858), .ZN(n4862)
         );
  NOR2_X1 U6002 ( .A1(n4863), .A2(n4862), .ZN(n5046) );
  NOR2_X1 U6003 ( .A1(n5047), .A2(n5046), .ZN(n5058) );
  AOI22_X1 U6004 ( .A1(n5195), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5189), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4867) );
  AOI22_X1 U6005 ( .A1(n5197), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4866) );
  AOI22_X1 U6006 ( .A1(n2999), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4865) );
  AOI22_X1 U6007 ( .A1(n5024), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4864) );
  NAND4_X1 U6008 ( .A1(n4867), .A2(n4866), .A3(n4865), .A4(n4864), .ZN(n4873)
         );
  AOI22_X1 U6009 ( .A1(n5198), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4871) );
  AOI22_X1 U6010 ( .A1(n5185), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4870) );
  AOI22_X1 U6011 ( .A1(n5187), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4869) );
  AOI22_X1 U6012 ( .A1(n5167), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4868) );
  NAND4_X1 U6013 ( .A1(n4871), .A2(n4870), .A3(n4869), .A4(n4868), .ZN(n4872)
         );
  OR2_X1 U6014 ( .A1(n4873), .A2(n4872), .ZN(n5056) );
  NAND2_X1 U6015 ( .A1(n5058), .A2(n5056), .ZN(n5068) );
  NOR2_X1 U6016 ( .A1(n5069), .A2(n5068), .ZN(n5126) );
  AOI22_X1 U6017 ( .A1(n5195), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5189), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4877) );
  AOI22_X1 U6018 ( .A1(n5197), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4876) );
  AOI22_X1 U6019 ( .A1(n2999), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4875) );
  AOI22_X1 U6020 ( .A1(n5024), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5188), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4874) );
  NAND4_X1 U6021 ( .A1(n4877), .A2(n4876), .A3(n4875), .A4(n4874), .ZN(n4883)
         );
  AOI22_X1 U6022 ( .A1(n5198), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4881) );
  AOI22_X1 U6023 ( .A1(n5185), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4880) );
  AOI22_X1 U6024 ( .A1(n5187), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4879) );
  AOI22_X1 U6025 ( .A1(n5167), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4878) );
  NAND4_X1 U6026 ( .A1(n4881), .A2(n4880), .A3(n4879), .A4(n4878), .ZN(n4882)
         );
  OR2_X1 U6027 ( .A1(n4883), .A2(n4882), .ZN(n5125) );
  XNOR2_X1 U6028 ( .A(n5126), .B(n5125), .ZN(n4887) );
  NAND2_X1 U6029 ( .A1(n4884), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5213) );
  AOI21_X1 U6030 ( .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6532), .A(n5216), 
        .ZN(n4886) );
  NAND2_X1 U6031 ( .A1(n5158), .A2(EAX_REG_26__SCAN_IN), .ZN(n4885) );
  OAI211_X1 U6032 ( .C1(n4887), .C2(n5213), .A(n4886), .B(n4885), .ZN(n4888)
         );
  OAI21_X1 U6033 ( .B1(n5210), .B2(n5348), .A(n4888), .ZN(n5080) );
  AOI22_X1 U6034 ( .A1(n5198), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5187), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4894) );
  AOI22_X1 U6035 ( .A1(n5197), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5195), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4893) );
  AOI22_X1 U6036 ( .A1(n5189), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4892) );
  AOI22_X1 U6037 ( .A1(n3000), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4891) );
  NAND4_X1 U6038 ( .A1(n4894), .A2(n4893), .A3(n4892), .A4(n4891), .ZN(n4900)
         );
  AOI22_X1 U6039 ( .A1(n2999), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n5024), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4898) );
  AOI22_X1 U6040 ( .A1(n5167), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4897) );
  AOI22_X1 U6041 ( .A1(n2998), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4896) );
  AOI22_X1 U6042 ( .A1(n5185), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4895) );
  NAND4_X1 U6043 ( .A1(n4898), .A2(n4897), .A3(n4896), .A4(n4895), .ZN(n4899)
         );
  NOR2_X1 U6044 ( .A1(n4900), .A2(n4899), .ZN(n4903) );
  OAI21_X1 U6045 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5575), .A(n5210), .ZN(
        n4901) );
  AOI21_X1 U6046 ( .B1(n5220), .B2(EAX_REG_21__SCAN_IN), .A(n4901), .ZN(n4902)
         );
  OAI21_X1 U6047 ( .B1(n5213), .B2(n4903), .A(n4902), .ZN(n4905) );
  XNOR2_X1 U6048 ( .A(n4922), .B(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5578)
         );
  NAND2_X1 U6049 ( .A1(n5578), .A2(n5216), .ZN(n4904) );
  AND2_X1 U6050 ( .A1(n4905), .A2(n4904), .ZN(n5088) );
  AOI22_X1 U6051 ( .A1(n5198), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4909) );
  AOI22_X1 U6052 ( .A1(n5197), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n5195), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4908) );
  AOI22_X1 U6053 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n5024), .B1(n3000), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4907) );
  AOI22_X1 U6054 ( .A1(n5167), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4906) );
  NAND4_X1 U6055 ( .A1(n4909), .A2(n4908), .A3(n4907), .A4(n4906), .ZN(n4915)
         );
  AOI22_X1 U6056 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5194), .B1(n5189), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4913) );
  AOI22_X1 U6057 ( .A1(n5185), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4912) );
  AOI22_X1 U6058 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5187), .B1(n5186), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4911) );
  AOI22_X1 U6059 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n2999), .B1(n5029), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4910) );
  NAND4_X1 U6060 ( .A1(n4913), .A2(n4912), .A3(n4911), .A4(n4910), .ZN(n4914)
         );
  NOR2_X1 U6061 ( .A1(n4915), .A2(n4914), .ZN(n4919) );
  OAI21_X1 U6062 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6538), .A(n6532), 
        .ZN(n4916) );
  INV_X1 U6063 ( .A(n4916), .ZN(n4917) );
  AOI21_X1 U6064 ( .B1(n5220), .B2(EAX_REG_20__SCAN_IN), .A(n4917), .ZN(n4918)
         );
  OAI21_X1 U6065 ( .B1(n5213), .B2(n4919), .A(n4918), .ZN(n4924) );
  INV_X1 U6066 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4920) );
  NAND2_X1 U6067 ( .A1(n4920), .A2(n4938), .ZN(n4921) );
  AND2_X1 U6068 ( .A1(n4922), .A2(n4921), .ZN(n5849) );
  NAND2_X1 U6069 ( .A1(n5849), .A2(n5216), .ZN(n4923) );
  AND2_X1 U6070 ( .A1(n4924), .A2(n4923), .ZN(n5424) );
  AOI22_X1 U6071 ( .A1(n5195), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5189), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4928) );
  AOI22_X1 U6072 ( .A1(n5197), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4927) );
  AOI22_X1 U6073 ( .A1(n2999), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4926) );
  AOI22_X1 U6074 ( .A1(n5024), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4925) );
  NAND4_X1 U6075 ( .A1(n4928), .A2(n4927), .A3(n4926), .A4(n4925), .ZN(n4934)
         );
  AOI22_X1 U6076 ( .A1(n5198), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4932) );
  AOI22_X1 U6077 ( .A1(n5185), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4931) );
  AOI22_X1 U6078 ( .A1(n5187), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4930) );
  AOI22_X1 U6079 ( .A1(n5167), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4929) );
  NAND4_X1 U6080 ( .A1(n4932), .A2(n4931), .A3(n4930), .A4(n4929), .ZN(n4933)
         );
  NOR2_X1 U6081 ( .A1(n4934), .A2(n4933), .ZN(n4937) );
  INV_X1 U6082 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6553) );
  AOI21_X1 U6083 ( .B1(n6553), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4935) );
  AOI21_X1 U6084 ( .B1(n5220), .B2(EAX_REG_19__SCAN_IN), .A(n4935), .ZN(n4936)
         );
  OAI21_X1 U6085 ( .B1(n5213), .B2(n4937), .A(n4936), .ZN(n4941) );
  NAND2_X1 U6086 ( .A1(n6553), .A2(n5018), .ZN(n4939) );
  AND2_X1 U6087 ( .A1(n4939), .A2(n4938), .ZN(n5860) );
  NAND2_X1 U6088 ( .A1(n5860), .A2(n5216), .ZN(n4940) );
  NAND2_X1 U6089 ( .A1(n4941), .A2(n4940), .ZN(n5436) );
  INV_X1 U6090 ( .A(n5436), .ZN(n5023) );
  XNOR2_X1 U6091 ( .A(n4942), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5977)
         );
  INV_X1 U6092 ( .A(n5213), .ZN(n5178) );
  AOI22_X1 U6093 ( .A1(n5185), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5187), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4946) );
  AOI22_X1 U6094 ( .A1(n5198), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4945) );
  AOI22_X1 U6095 ( .A1(n5195), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5189), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4944) );
  AOI22_X1 U6096 ( .A1(n5024), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4943) );
  NAND4_X1 U6097 ( .A1(n4946), .A2(n4945), .A3(n4944), .A4(n4943), .ZN(n4952)
         );
  AOI22_X1 U6098 ( .A1(n5197), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4950) );
  AOI22_X1 U6099 ( .A1(n5186), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4949) );
  AOI22_X1 U6100 ( .A1(n2999), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4948) );
  AOI22_X1 U6101 ( .A1(n5167), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4947) );
  NAND4_X1 U6102 ( .A1(n4950), .A2(n4949), .A3(n4948), .A4(n4947), .ZN(n4951)
         );
  OR2_X1 U6103 ( .A1(n4952), .A2(n4951), .ZN(n4955) );
  NAND2_X1 U6104 ( .A1(n6532), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4953)
         );
  OAI211_X1 U6105 ( .C1(n5064), .C2(n3701), .A(n5210), .B(n4953), .ZN(n4954)
         );
  AOI21_X1 U6106 ( .B1(n5178), .B2(n4955), .A(n4954), .ZN(n4956) );
  AOI21_X1 U6107 ( .B1(n5977), .B2(n5216), .A(n4956), .ZN(n5458) );
  XOR2_X1 U6108 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n4957), .Z(n5988) );
  INV_X1 U6109 ( .A(n5988), .ZN(n5607) );
  AOI22_X1 U6110 ( .A1(n5198), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4961) );
  AOI22_X1 U6111 ( .A1(n2999), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n5024), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4960) );
  AOI22_X1 U6112 ( .A1(n5185), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5187), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4959) );
  AOI22_X1 U6113 ( .A1(n5167), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4958) );
  NAND4_X1 U6114 ( .A1(n4961), .A2(n4960), .A3(n4959), .A4(n4958), .ZN(n4967)
         );
  AOI22_X1 U6115 ( .A1(n5197), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5195), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4965) );
  AOI22_X1 U6116 ( .A1(n5186), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4964) );
  AOI22_X1 U6117 ( .A1(n3000), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4963) );
  AOI22_X1 U6118 ( .A1(n5189), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4962) );
  NAND4_X1 U6119 ( .A1(n4965), .A2(n4964), .A3(n4963), .A4(n4962), .ZN(n4966)
         );
  NOR2_X1 U6120 ( .A1(n4967), .A2(n4966), .ZN(n4969) );
  AOI22_X1 U6121 ( .A1(n5220), .A2(EAX_REG_16__SCAN_IN), .B1(n5219), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4968) );
  OAI21_X1 U6122 ( .B1(n5213), .B2(n4969), .A(n4968), .ZN(n4970) );
  AOI21_X1 U6123 ( .B1(n5607), .B2(n5216), .A(n4970), .ZN(n5469) );
  AOI22_X1 U6124 ( .A1(n5198), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5195), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4974) );
  AOI22_X1 U6125 ( .A1(n2999), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n5024), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4973) );
  AOI22_X1 U6126 ( .A1(n5197), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4972) );
  AOI22_X1 U6127 ( .A1(n5186), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4971) );
  NAND4_X1 U6128 ( .A1(n4974), .A2(n4973), .A3(n4972), .A4(n4971), .ZN(n4980)
         );
  AOI22_X1 U6129 ( .A1(n2998), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5167), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4978) );
  AOI22_X1 U6130 ( .A1(n5185), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5187), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4977) );
  AOI22_X1 U6131 ( .A1(n5189), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4976) );
  AOI22_X1 U6132 ( .A1(n3000), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4975) );
  NAND4_X1 U6133 ( .A1(n4978), .A2(n4977), .A3(n4976), .A4(n4975), .ZN(n4979)
         );
  OAI21_X1 U6134 ( .B1(n4980), .B2(n4979), .A(n4998), .ZN(n4985) );
  INV_X1 U6135 ( .A(n4981), .ZN(n4982) );
  XNOR2_X1 U6136 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n4982), .ZN(n5614)
         );
  AOI22_X1 U6137 ( .A1(n5216), .A2(n5614), .B1(n5219), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4984) );
  NAND2_X1 U6138 ( .A1(n5220), .A2(EAX_REG_15__SCAN_IN), .ZN(n4983) );
  AND3_X1 U6139 ( .A1(n4985), .A2(n4984), .A3(n4983), .ZN(n5386) );
  NOR2_X1 U6140 ( .A1(n5469), .A2(n5386), .ZN(n5455) );
  AND2_X1 U6141 ( .A1(n5458), .A2(n5455), .ZN(n5003) );
  INV_X1 U6142 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5515) );
  OAI21_X1 U6143 ( .B1(PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n6538), .A(n6532), 
        .ZN(n4986) );
  OAI21_X1 U6144 ( .B1(n5064), .B2(n5515), .A(n4986), .ZN(n4989) );
  XOR2_X1 U6145 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4987), .Z(n5998) );
  NAND2_X1 U6146 ( .A1(n5216), .A2(n5998), .ZN(n4988) );
  NAND2_X1 U6147 ( .A1(n4989), .A2(n4988), .ZN(n5002) );
  AOI22_X1 U6148 ( .A1(n5167), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n5189), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4993) );
  AOI22_X1 U6149 ( .A1(n5197), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4992) );
  AOI22_X1 U6150 ( .A1(n5198), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4991) );
  AOI22_X1 U6151 ( .A1(n5185), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4990) );
  NAND4_X1 U6152 ( .A1(n4993), .A2(n4992), .A3(n4991), .A4(n4990), .ZN(n5000)
         );
  AOI22_X1 U6153 ( .A1(n2998), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5187), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4997) );
  AOI22_X1 U6154 ( .A1(n2999), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4996) );
  AOI22_X1 U6155 ( .A1(n5195), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4995) );
  AOI22_X1 U6156 ( .A1(n5024), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4994) );
  NAND4_X1 U6157 ( .A1(n4997), .A2(n4996), .A3(n4995), .A4(n4994), .ZN(n4999)
         );
  OAI21_X1 U6158 ( .B1(n5000), .B2(n4999), .A(n4998), .ZN(n5001) );
  NAND2_X1 U6159 ( .A1(n5002), .A2(n5001), .ZN(n5478) );
  AND2_X1 U6160 ( .A1(n5003), .A2(n5478), .ZN(n5445) );
  AOI22_X1 U6161 ( .A1(n5198), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5007) );
  AOI22_X1 U6162 ( .A1(n5195), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5006) );
  AOI22_X1 U6163 ( .A1(n5189), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5005) );
  AOI22_X1 U6164 ( .A1(n2999), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5004) );
  NAND4_X1 U6165 ( .A1(n5007), .A2(n5006), .A3(n5005), .A4(n5004), .ZN(n5013)
         );
  AOI22_X1 U6166 ( .A1(n5197), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5024), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5011) );
  AOI22_X1 U6167 ( .A1(n5167), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n5010) );
  AOI22_X1 U6168 ( .A1(n5187), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5009) );
  AOI22_X1 U6169 ( .A1(n5185), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5008) );
  NAND4_X1 U6170 ( .A1(n5011), .A2(n5010), .A3(n5009), .A4(n5008), .ZN(n5012)
         );
  NOR2_X1 U6171 ( .A1(n5013), .A2(n5012), .ZN(n5017) );
  NAND2_X1 U6172 ( .A1(n6532), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5014)
         );
  NAND2_X1 U6173 ( .A1(n5210), .A2(n5014), .ZN(n5015) );
  AOI21_X1 U6174 ( .B1(n5220), .B2(EAX_REG_18__SCAN_IN), .A(n5015), .ZN(n5016)
         );
  OAI21_X1 U6175 ( .B1(n5213), .B2(n5017), .A(n5016), .ZN(n5021) );
  OAI21_X1 U6176 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n5019), .A(n5018), 
        .ZN(n5970) );
  OR2_X1 U6177 ( .A1(n5210), .A2(n5970), .ZN(n5020) );
  NAND2_X1 U6178 ( .A1(n5021), .A2(n5020), .ZN(n5446) );
  INV_X1 U6179 ( .A(n5446), .ZN(n5022) );
  AND2_X1 U6180 ( .A1(n5445), .A2(n5022), .ZN(n5435) );
  AND2_X1 U6181 ( .A1(n5023), .A2(n5435), .ZN(n5425) );
  AND2_X1 U6182 ( .A1(n5424), .A2(n5425), .ZN(n5087) );
  AND2_X1 U6183 ( .A1(n5088), .A2(n5087), .ZN(n5086) );
  AOI22_X1 U6184 ( .A1(n2998), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5187), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n5028) );
  AOI22_X1 U6185 ( .A1(n5198), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5167), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5027) );
  AOI22_X1 U6186 ( .A1(n5024), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5026) );
  AOI22_X1 U6187 ( .A1(n5195), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5025) );
  NAND4_X1 U6188 ( .A1(n5028), .A2(n5027), .A3(n5026), .A4(n5025), .ZN(n5035)
         );
  AOI22_X1 U6189 ( .A1(n5197), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5033) );
  AOI22_X1 U6190 ( .A1(n5185), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5032) );
  AOI22_X1 U6191 ( .A1(n5189), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5031) );
  AOI22_X1 U6192 ( .A1(n2999), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n5029), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5030) );
  NAND4_X1 U6193 ( .A1(n5033), .A2(n5032), .A3(n5031), .A4(n5030), .ZN(n5034)
         );
  NOR2_X1 U6194 ( .A1(n5035), .A2(n5034), .ZN(n5039) );
  NAND2_X1 U6195 ( .A1(n6532), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5036)
         );
  NAND2_X1 U6196 ( .A1(n5210), .A2(n5036), .ZN(n5037) );
  AOI21_X1 U6197 ( .B1(n5220), .B2(EAX_REG_22__SCAN_IN), .A(n5037), .ZN(n5038)
         );
  OAI21_X1 U6198 ( .B1(n5213), .B2(n5039), .A(n5038), .ZN(n5044) );
  INV_X1 U6199 ( .A(n5040), .ZN(n5041) );
  INV_X1 U6200 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U6201 ( .A1(n5041), .A2(n5566), .ZN(n5042) );
  NAND2_X1 U6202 ( .A1(n5052), .A2(n5042), .ZN(n5835) );
  OR2_X1 U6203 ( .A1(n5835), .A2(n5210), .ZN(n5043) );
  NAND2_X1 U6204 ( .A1(n5044), .A2(n5043), .ZN(n5412) );
  INV_X1 U6205 ( .A(n5412), .ZN(n5045) );
  AND2_X1 U6206 ( .A1(n5086), .A2(n5045), .ZN(n5103) );
  XOR2_X1 U6207 ( .A(n5047), .B(n5046), .Z(n5048) );
  NAND2_X1 U6208 ( .A1(n5048), .A2(n5178), .ZN(n5051) );
  INV_X1 U6209 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5557) );
  AOI21_X1 U6210 ( .B1(n5557), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n5049) );
  AOI21_X1 U6211 ( .B1(n5220), .B2(EAX_REG_23__SCAN_IN), .A(n5049), .ZN(n5050)
         );
  NAND2_X1 U6212 ( .A1(n5051), .A2(n5050), .ZN(n5054) );
  XNOR2_X1 U6213 ( .A(n5052), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5561)
         );
  NAND2_X1 U6214 ( .A1(n5561), .A2(n5216), .ZN(n5053) );
  NAND2_X1 U6215 ( .A1(n5054), .A2(n5053), .ZN(n5104) );
  INV_X1 U6216 ( .A(n5104), .ZN(n5055) );
  AND2_X1 U6217 ( .A1(n5103), .A2(n5055), .ZN(n5102) );
  INV_X1 U6218 ( .A(n5056), .ZN(n5057) );
  XNOR2_X1 U6219 ( .A(n5058), .B(n5057), .ZN(n5066) );
  INV_X1 U6220 ( .A(n5059), .ZN(n5060) );
  INV_X1 U6221 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6222 ( .A1(n5060), .A2(n5376), .ZN(n5061) );
  NAND2_X1 U6223 ( .A1(n5062), .A2(n5061), .ZN(n5375) );
  AOI22_X1 U6224 ( .A1(n5375), .A2(n5216), .B1(PHYADDRPOINTER_REG_24__SCAN_IN), 
        .B2(n5219), .ZN(n5063) );
  OAI21_X1 U6225 ( .B1(n5064), .B2(n3707), .A(n5063), .ZN(n5065) );
  AOI21_X1 U6226 ( .B1(n5066), .B2(n5178), .A(n5065), .ZN(n5257) );
  INV_X1 U6227 ( .A(n5257), .ZN(n5067) );
  AND2_X1 U6228 ( .A1(n5102), .A2(n5067), .ZN(n5356) );
  INV_X1 U6229 ( .A(n5356), .ZN(n5076) );
  XOR2_X1 U6230 ( .A(n5069), .B(n5068), .Z(n5070) );
  NAND2_X1 U6231 ( .A1(n5070), .A2(n5178), .ZN(n5074) );
  INV_X1 U6232 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5547) );
  NOR2_X1 U6233 ( .A1(n5547), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5071) );
  AOI211_X1 U6234 ( .C1(n5220), .C2(EAX_REG_25__SCAN_IN), .A(n5216), .B(n5071), 
        .ZN(n5073) );
  XOR2_X1 U6235 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .B(n5072), .Z(n5551) );
  AOI22_X1 U6236 ( .A1(n5074), .A2(n5073), .B1(n5216), .B2(n5551), .ZN(n5358)
         );
  INV_X1 U6237 ( .A(n5358), .ZN(n5075) );
  NOR2_X1 U6238 ( .A1(n5076), .A2(n5075), .ZN(n5078) );
  NAND2_X1 U6239 ( .A1(n5479), .A2(n5078), .ZN(n5357) );
  INV_X1 U6240 ( .A(n5080), .ZN(n5077) );
  AND2_X1 U6241 ( .A1(n5078), .A2(n5077), .ZN(n5079) );
  AND2_X2 U6242 ( .A1(n5479), .A2(n5079), .ZN(n5339) );
  AOI21_X1 U6243 ( .B1(n5080), .B2(n5357), .A(n5339), .ZN(n5404) );
  NOR2_X1 U6244 ( .A1(n6225), .A2(n5348), .ZN(n5083) );
  OAI21_X1 U6245 ( .B1(n6208), .B2(n5349), .A(n5081), .ZN(n5082) );
  AOI211_X1 U6246 ( .C1(n5404), .C2(n6219), .A(n5083), .B(n5082), .ZN(n5084)
         );
  OAI21_X1 U6247 ( .B1(n6195), .B2(n5085), .A(n5084), .ZN(U2960) );
  NAND2_X1 U6248 ( .A1(n5479), .A2(n5086), .ZN(n5413) );
  AND2_X1 U6249 ( .A1(n5479), .A2(n5087), .ZN(n5426) );
  OR2_X1 U6250 ( .A1(n5426), .A2(n5088), .ZN(n5089) );
  INV_X1 U6251 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6487) );
  INV_X1 U6252 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6485) );
  NAND2_X1 U6253 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5090), .ZN(n6003) );
  NOR2_X1 U6254 ( .A1(n6485), .A2(n6003), .ZN(n5993) );
  NAND2_X1 U6255 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5993), .ZN(n5389) );
  NOR2_X1 U6256 ( .A1(n6487), .A2(n5389), .ZN(n5971) );
  NAND3_X1 U6257 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        n5971), .ZN(n5091) );
  NOR2_X1 U6258 ( .A1(n6090), .A2(n5091), .ZN(n5964) );
  NAND4_X1 U6259 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(n5964), .ZN(n5840) );
  NOR2_X1 U6260 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5840), .ZN(n5839) );
  INV_X1 U6261 ( .A(n5091), .ZN(n5092) );
  NAND2_X1 U6262 ( .A1(n6050), .A2(n5092), .ZN(n5093) );
  NAND2_X1 U6263 ( .A1(n5303), .A2(n5093), .ZN(n5973) );
  INV_X1 U6264 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6497) );
  INV_X1 U6265 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6495) );
  INV_X1 U6266 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6492) );
  NOR2_X1 U6267 ( .A1(n6495), .A2(n6492), .ZN(n5846) );
  INV_X1 U6268 ( .A(n5846), .ZN(n5854) );
  OR2_X1 U6269 ( .A1(n6497), .A2(n5854), .ZN(n5094) );
  NAND2_X1 U6270 ( .A1(n5303), .A2(n5094), .ZN(n5095) );
  NAND2_X1 U6271 ( .A1(n5973), .A2(n5095), .ZN(n5838) );
  INV_X1 U6272 ( .A(n5838), .ZN(n5853) );
  INV_X1 U6273 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5841) );
  OAI22_X1 U6274 ( .A1(n5853), .A2(n5841), .B1(n5575), .B2(n6073), .ZN(n5100)
         );
  AOI21_X1 U6275 ( .B1(n5097), .B2(n5096), .A(n5417), .ZN(n5683) );
  INV_X1 U6276 ( .A(n5683), .ZN(n5422) );
  AOI22_X1 U6277 ( .A1(n6089), .A2(EBX_REG_21__SCAN_IN), .B1(n5578), .B2(n6079), .ZN(n5098) );
  OAI21_X1 U6278 ( .B1(n5422), .B2(n6065), .A(n5098), .ZN(n5099) );
  NOR3_X1 U6279 ( .A1(n5839), .A2(n5100), .A3(n5099), .ZN(n5101) );
  OAI21_X1 U6280 ( .B1(n5867), .B2(n6058), .A(n5101), .ZN(U2806) );
  NAND2_X1 U6281 ( .A1(n5479), .A2(n5102), .ZN(n5256) );
  NAND2_X1 U6282 ( .A1(n5479), .A2(n5103), .ZN(n5415) );
  NAND2_X1 U6283 ( .A1(n5415), .A2(n5104), .ZN(n5105) );
  NAND2_X1 U6284 ( .A1(n5256), .A2(n5105), .ZN(n5558) );
  NOR2_X2 U6285 ( .A1(n6122), .A2(n5106), .ZN(n6119) );
  AOI22_X1 U6286 ( .A1(n6119), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6122), .ZN(n5111) );
  AND2_X1 U6287 ( .A1(n5108), .A2(n5107), .ZN(n5109) );
  NAND2_X1 U6288 ( .A1(n6123), .A2(DATAI_7_), .ZN(n5110) );
  OAI211_X1 U6289 ( .C1(n5558), .C2(n5863), .A(n5111), .B(n5110), .ZN(U2868)
         );
  OAI21_X1 U6290 ( .B1(n5419), .B2(n5112), .A(n5250), .ZN(n5667) );
  INV_X1 U6291 ( .A(n5667), .ZN(n5113) );
  AOI22_X1 U6292 ( .A1(n5113), .A2(n6107), .B1(n5399), .B2(EBX_REG_23__SCAN_IN), .ZN(n5114) );
  OAI21_X1 U6293 ( .B1(n5558), .B2(n5466), .A(n5114), .ZN(U2836) );
  INV_X1 U6294 ( .A(n6089), .ZN(n6043) );
  OAI22_X1 U6295 ( .A1(n5115), .A2(n6043), .B1(n5557), .B2(n6073), .ZN(n5117)
         );
  NOR2_X1 U6296 ( .A1(n5667), .A2(n6065), .ZN(n5116) );
  AOI211_X1 U6297 ( .C1(n6079), .C2(n5561), .A(n5117), .B(n5116), .ZN(n5122)
         );
  INV_X1 U6298 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6499) );
  NOR3_X1 U6299 ( .A1(n6499), .A2(n5841), .A3(n5840), .ZN(n5227) );
  NAND2_X1 U6300 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5118) );
  INV_X1 U6301 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6655) );
  OAI21_X1 U6302 ( .B1(n5118), .B2(n6655), .A(n5303), .ZN(n5119) );
  INV_X1 U6303 ( .A(n5119), .ZN(n5120) );
  NOR2_X1 U6304 ( .A1(n5838), .A2(n5120), .ZN(n5377) );
  INV_X1 U6305 ( .A(n5377), .ZN(n5361) );
  OAI21_X1 U6306 ( .B1(n5227), .B2(REIP_REG_23__SCAN_IN), .A(n5361), .ZN(n5121) );
  OAI211_X1 U6307 ( .C1(n5558), .C2(n6058), .A(n5122), .B(n5121), .ZN(U2804)
         );
  INV_X1 U6308 ( .A(n5123), .ZN(n5238) );
  OAI22_X1 U6309 ( .A1(n5238), .A2(n6103), .B1(n5124), .B2(n5486), .ZN(U2828)
         );
  NAND2_X1 U6310 ( .A1(n5126), .A2(n5125), .ZN(n5146) );
  AOI22_X1 U6311 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n2998), .B1(n5167), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5130) );
  AOI22_X1 U6312 ( .A1(n5197), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5129) );
  AOI22_X1 U6313 ( .A1(n5186), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n5128) );
  AOI22_X1 U6314 ( .A1(n5196), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n5188), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5127) );
  NAND4_X1 U6315 ( .A1(n5130), .A2(n5129), .A3(n5128), .A4(n5127), .ZN(n5136)
         );
  AOI22_X1 U6316 ( .A1(n5185), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n5187), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5134) );
  AOI22_X1 U6317 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n5189), .B1(n5195), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n5133) );
  AOI22_X1 U6318 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n2999), .B1(n3000), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5132) );
  AOI22_X1 U6319 ( .A1(n5198), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5131) );
  NAND4_X1 U6320 ( .A1(n5134), .A2(n5133), .A3(n5132), .A4(n5131), .ZN(n5135)
         );
  NOR2_X1 U6321 ( .A1(n5136), .A2(n5135), .ZN(n5147) );
  XOR2_X1 U6322 ( .A(n5146), .B(n5147), .Z(n5137) );
  NAND2_X1 U6323 ( .A1(n5137), .A2(n5178), .ZN(n5141) );
  NOR2_X1 U6324 ( .A1(n5539), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5138) );
  AOI211_X1 U6325 ( .C1(n5220), .C2(EAX_REG_27__SCAN_IN), .A(n5216), .B(n5138), 
        .ZN(n5140) );
  XNOR2_X1 U6326 ( .A(n5139), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5543)
         );
  AOI22_X1 U6327 ( .A1(n5141), .A2(n5140), .B1(n5216), .B2(n5543), .ZN(n5338)
         );
  NAND2_X1 U6328 ( .A1(n5143), .A2(n5142), .ZN(n5144) );
  NAND2_X1 U6329 ( .A1(n5145), .A2(n5144), .ZN(n5532) );
  NOR2_X1 U6330 ( .A1(n5147), .A2(n5146), .ZN(n5166) );
  AOI22_X1 U6331 ( .A1(n5195), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5189), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5151) );
  AOI22_X1 U6332 ( .A1(n5197), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5150) );
  AOI22_X1 U6333 ( .A1(n2999), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5149) );
  AOI22_X1 U6334 ( .A1(n5196), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5188), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5148) );
  NAND4_X1 U6335 ( .A1(n5151), .A2(n5150), .A3(n5149), .A4(n5148), .ZN(n5157)
         );
  AOI22_X1 U6336 ( .A1(n5198), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n2998), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n5155) );
  AOI22_X1 U6337 ( .A1(n5185), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n5154) );
  AOI22_X1 U6338 ( .A1(n5187), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5153) );
  AOI22_X1 U6339 ( .A1(n5167), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5152) );
  NAND4_X1 U6340 ( .A1(n5155), .A2(n5154), .A3(n5153), .A4(n5152), .ZN(n5156)
         );
  OR2_X1 U6341 ( .A1(n5157), .A2(n5156), .ZN(n5165) );
  XNOR2_X1 U6342 ( .A(n5166), .B(n5165), .ZN(n5161) );
  AOI21_X1 U6343 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6532), .A(n5216), 
        .ZN(n5160) );
  NAND2_X1 U6344 ( .A1(n5158), .A2(EAX_REG_28__SCAN_IN), .ZN(n5159) );
  OAI211_X1 U6345 ( .C1(n5161), .C2(n5213), .A(n5160), .B(n5159), .ZN(n5162)
         );
  OAI21_X1 U6346 ( .B1(n5210), .B2(n5532), .A(n5162), .ZN(n5326) );
  INV_X1 U6347 ( .A(n5326), .ZN(n5163) );
  AND2_X1 U6348 ( .A1(n5338), .A2(n5163), .ZN(n5164) );
  AND2_X2 U6349 ( .A1(n5339), .A2(n5164), .ZN(n5325) );
  NAND2_X1 U6350 ( .A1(n5166), .A2(n5165), .ZN(n5205) );
  AOI22_X1 U6351 ( .A1(n2998), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5167), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5171) );
  AOI22_X1 U6352 ( .A1(n5195), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5170) );
  AOI22_X1 U6353 ( .A1(n5185), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5169) );
  AOI22_X1 U6354 ( .A1(n2999), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n5188), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5168) );
  NAND4_X1 U6355 ( .A1(n5171), .A2(n5170), .A3(n5169), .A4(n5168), .ZN(n5177)
         );
  AOI22_X1 U6356 ( .A1(n5197), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5196), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5175) );
  AOI22_X1 U6357 ( .A1(n5189), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5174) );
  AOI22_X1 U6358 ( .A1(n5187), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n5173) );
  AOI22_X1 U6359 ( .A1(n5198), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5172) );
  NAND4_X1 U6360 ( .A1(n5175), .A2(n5174), .A3(n5173), .A4(n5172), .ZN(n5176)
         );
  NOR2_X1 U6361 ( .A1(n5177), .A2(n5176), .ZN(n5206) );
  XOR2_X1 U6362 ( .A(n5205), .B(n5206), .Z(n5179) );
  NAND2_X1 U6363 ( .A1(n5179), .A2(n5178), .ZN(n5183) );
  INV_X1 U6364 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5284) );
  NOR2_X1 U6365 ( .A1(n5284), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5180) );
  AOI211_X1 U6366 ( .C1(n5220), .C2(EAX_REG_29__SCAN_IN), .A(n5216), .B(n5180), 
        .ZN(n5182) );
  XOR2_X1 U6367 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .B(n5181), .Z(n5286) );
  AOI22_X1 U6368 ( .A1(n5183), .A2(n5182), .B1(n5216), .B2(n5286), .ZN(n5280)
         );
  AOI22_X1 U6369 ( .A1(n2998), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5167), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5193) );
  AOI22_X1 U6370 ( .A1(n5185), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5184), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5192) );
  AOI22_X1 U6371 ( .A1(n5187), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5186), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5191) );
  AOI22_X1 U6372 ( .A1(n5189), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5188), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5190) );
  NAND4_X1 U6373 ( .A1(n5193), .A2(n5192), .A3(n5191), .A4(n5190), .ZN(n5204)
         );
  AOI22_X1 U6374 ( .A1(n5195), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5194), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5202) );
  AOI22_X1 U6375 ( .A1(n2999), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n5196), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5201) );
  AOI22_X1 U6376 ( .A1(n5197), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5200) );
  AOI22_X1 U6377 ( .A1(n5198), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3001), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5199) );
  NAND4_X1 U6378 ( .A1(n5202), .A2(n5201), .A3(n5200), .A4(n5199), .ZN(n5203)
         );
  NOR2_X1 U6379 ( .A1(n5204), .A2(n5203), .ZN(n5208) );
  NOR2_X1 U6380 ( .A1(n5206), .A2(n5205), .ZN(n5207) );
  XOR2_X1 U6381 ( .A(n5208), .B(n5207), .Z(n5214) );
  NAND2_X1 U6382 ( .A1(n6532), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5209)
         );
  NAND2_X1 U6383 ( .A1(n5210), .A2(n5209), .ZN(n5211) );
  AOI21_X1 U6384 ( .B1(n5220), .B2(EAX_REG_30__SCAN_IN), .A(n5211), .ZN(n5212)
         );
  OAI21_X1 U6385 ( .B1(n5214), .B2(n5213), .A(n5212), .ZN(n5218) );
  XNOR2_X1 U6386 ( .A(n5215), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5517)
         );
  NAND2_X1 U6387 ( .A1(n5517), .A2(n5216), .ZN(n5217) );
  NAND2_X1 U6388 ( .A1(n5218), .A2(n5217), .ZN(n5313) );
  NOR2_X1 U6389 ( .A1(n5312), .A2(n5313), .ZN(n5222) );
  AOI22_X1 U6390 ( .A1(n5220), .A2(EAX_REG_31__SCAN_IN), .B1(n5219), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5221) );
  XNOR2_X1 U6391 ( .A(n5222), .B(n5221), .ZN(n5490) );
  NAND2_X1 U6392 ( .A1(n5490), .A2(n6032), .ZN(n5237) );
  INV_X1 U6393 ( .A(n6090), .ZN(n6083) );
  INV_X1 U6394 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6512) );
  INV_X1 U6395 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6501) );
  NAND2_X1 U6396 ( .A1(REIP_REG_26__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5229) );
  OAI21_X1 U6397 ( .B1(n6501), .B2(n5229), .A(n5303), .ZN(n5223) );
  NAND2_X1 U6398 ( .A1(n5377), .A2(n5223), .ZN(n5353) );
  NAND2_X1 U6399 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5224) );
  AND2_X1 U6400 ( .A1(n6083), .A2(n5224), .ZN(n5225) );
  OR2_X1 U6401 ( .A1(n5353), .A2(n5225), .ZN(n5331) );
  AOI21_X1 U6402 ( .B1(n6083), .B2(n6512), .A(n5331), .ZN(n5319) );
  OAI21_X1 U6403 ( .B1(REIP_REG_30__SCAN_IN), .B2(n6090), .A(n5319), .ZN(n5235) );
  INV_X1 U6404 ( .A(n5226), .ZN(n5233) );
  NAND2_X1 U6405 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5227), .ZN(n5360) );
  INV_X1 U6406 ( .A(n5360), .ZN(n5228) );
  NAND2_X1 U6407 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5228), .ZN(n5362) );
  NOR2_X1 U6408 ( .A1(n5362), .A2(n5229), .ZN(n5341) );
  NAND3_X1 U6409 ( .A1(n5341), .A2(REIP_REG_28__SCAN_IN), .A3(
        REIP_REG_27__SCAN_IN), .ZN(n5314) );
  INV_X1 U6410 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6516) );
  NOR4_X1 U6411 ( .A1(n5314), .A2(REIP_REG_31__SCAN_IN), .A3(n6516), .A4(n6512), .ZN(n5230) );
  AOI21_X1 U6412 ( .B1(n6091), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5230), 
        .ZN(n5231) );
  OAI21_X1 U6413 ( .B1(n5233), .B2(n5232), .A(n5231), .ZN(n5234) );
  AOI21_X1 U6414 ( .B1(n5235), .B2(REIP_REG_31__SCAN_IN), .A(n5234), .ZN(n5236) );
  OAI211_X1 U6415 ( .C1(n5238), .C2(n6065), .A(n5237), .B(n5236), .ZN(U2796)
         );
  INV_X1 U6416 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5704) );
  XNOR2_X1 U6417 ( .A(n2996), .B(n5704), .ZN(n5588) );
  NAND2_X1 U6418 ( .A1(n2996), .A2(n5704), .ZN(n5239) );
  INV_X1 U6419 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5580) );
  AND2_X1 U6420 ( .A1(n2996), .A2(n5580), .ZN(n5240) );
  INV_X1 U6421 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5688) );
  XNOR2_X1 U6422 ( .A(n2996), .B(n5688), .ZN(n5574) );
  INV_X1 U6423 ( .A(n5574), .ZN(n5242) );
  NAND2_X1 U6424 ( .A1(n5241), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5570) );
  AND2_X1 U6425 ( .A1(n5242), .A2(n5570), .ZN(n5243) );
  NOR2_X1 U6426 ( .A1(n2996), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5563)
         );
  NAND2_X1 U6427 ( .A1(n5572), .A2(n5563), .ZN(n5553) );
  AND2_X1 U6428 ( .A1(n2996), .A2(n3010), .ZN(n5246) );
  NAND2_X1 U6429 ( .A1(n5564), .A2(n5246), .ZN(n5247) );
  OAI21_X1 U6430 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5553), .A(n5247), 
        .ZN(n5248) );
  XNOR2_X1 U6431 ( .A(n5248), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5262)
         );
  INV_X1 U6432 ( .A(n5369), .ZN(n5249) );
  AOI21_X1 U6433 ( .B1(n5251), .B2(n5250), .A(n5249), .ZN(n5410) );
  AND2_X1 U6434 ( .A1(n2997), .A2(REIP_REG_24__SCAN_IN), .ZN(n5258) );
  INV_X1 U6435 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5253) );
  AOI211_X1 U6436 ( .C1(n5253), .C2(n5668), .A(n5252), .B(n5660), .ZN(n5254)
         );
  AOI211_X1 U6437 ( .C1(n6288), .C2(n5410), .A(n5258), .B(n5254), .ZN(n5255)
         );
  OAI21_X1 U6438 ( .B1(n5262), .B2(n6269), .A(n5255), .ZN(U2994) );
  XOR2_X1 U6439 ( .A(n5257), .B(n5256), .Z(n5374) );
  AOI21_X1 U6440 ( .B1(n6218), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5258), 
        .ZN(n5259) );
  OAI21_X1 U6441 ( .B1(n5375), .B2(n6225), .A(n5259), .ZN(n5260) );
  AOI21_X1 U6442 ( .B1(n5374), .B2(n6219), .A(n5260), .ZN(n5261) );
  OAI21_X1 U6443 ( .B1(n5262), .B2(n6195), .A(n5261), .ZN(U2962) );
  NAND2_X1 U6444 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5263)
         );
  OAI211_X1 U6445 ( .C1(n6225), .C2(n5265), .A(n5264), .B(n5263), .ZN(n5266)
         );
  AOI21_X1 U6446 ( .B1(n5490), .B2(n6219), .A(n5266), .ZN(n5267) );
  OAI21_X1 U6447 ( .B1(n5268), .B2(n6195), .A(n5267), .ZN(U2955) );
  AOI22_X1 U6448 ( .A1(n5270), .A2(n6367), .B1(INSTQUEUE_REG_6__5__SCAN_IN), 
        .B2(n5269), .ZN(n5274) );
  AOI22_X1 U6449 ( .A1(n6365), .A2(n5272), .B1(n5271), .B2(n5813), .ZN(n5273)
         );
  OAI211_X1 U6450 ( .C1(n5811), .C2(n5275), .A(n5274), .B(n5273), .ZN(U3073)
         );
  INV_X1 U6451 ( .A(n5276), .ZN(n5277) );
  OR2_X1 U6452 ( .A1(n5278), .A2(n5277), .ZN(n5279) );
  XNOR2_X1 U6453 ( .A(n5279), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5639)
         );
  NAND2_X1 U6454 ( .A1(n2997), .A2(REIP_REG_29__SCAN_IN), .ZN(n5633) );
  OAI21_X1 U6455 ( .B1(n6208), .B2(n5284), .A(n5633), .ZN(n5282) );
  OAI21_X2 U6456 ( .B1(n5325), .B2(n5280), .A(n5312), .ZN(n5307) );
  NOR2_X1 U6457 ( .A1(n5307), .A2(n6194), .ZN(n5281) );
  OAI21_X1 U6458 ( .B1(n5639), .B2(n6195), .A(n5283), .ZN(U2957) );
  OAI22_X1 U6459 ( .A1(n6073), .A2(n5284), .B1(REIP_REG_29__SCAN_IN), .B2(
        n5314), .ZN(n5285) );
  AOI21_X1 U6460 ( .B1(n5286), .B2(n6079), .A(n5285), .ZN(n5287) );
  OAI21_X1 U6461 ( .B1(n6043), .B2(n5308), .A(n5287), .ZN(n5294) );
  OAI211_X1 U6462 ( .C1(n5439), .C2(n5289), .A(n5324), .B(n5288), .ZN(n5290)
         );
  INV_X1 U6463 ( .A(n5290), .ZN(n5291) );
  OR2_X1 U6464 ( .A1(n5292), .A2(n5291), .ZN(n5634) );
  NOR2_X1 U6465 ( .A1(n5634), .A2(n6065), .ZN(n5293) );
  OAI21_X1 U6466 ( .B1(n5307), .B2(n6058), .A(n5295), .ZN(U2798) );
  AOI22_X1 U6467 ( .A1(n6119), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6122), .ZN(n5297) );
  NAND2_X1 U6468 ( .A1(n6123), .A2(DATAI_13_), .ZN(n5296) );
  OAI211_X1 U6469 ( .C1(n5307), .C2(n5863), .A(n5297), .B(n5296), .ZN(U2862)
         );
  INV_X1 U6470 ( .A(n5298), .ZN(n5625) );
  NAND2_X1 U6471 ( .A1(n5625), .A2(n6098), .ZN(n5305) );
  OAI21_X1 U6472 ( .B1(n6091), .B2(n6079), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5299) );
  OAI21_X1 U6473 ( .B1(n6043), .B2(n5300), .A(n5299), .ZN(n5302) );
  NOR2_X1 U6474 ( .A1(n6065), .A2(n6302), .ZN(n5301) );
  AOI211_X1 U6475 ( .C1(REIP_REG_0__SCAN_IN), .C2(n5303), .A(n5302), .B(n5301), 
        .ZN(n5304) );
  OAI211_X1 U6476 ( .C1(n6095), .C2(n5306), .A(n5305), .B(n5304), .ZN(U2827)
         );
  OAI222_X1 U6477 ( .A1(n5308), .A2(n6111), .B1(n6103), .B2(n5634), .C1(n5307), 
        .C2(n5466), .ZN(U2830) );
  NAND2_X1 U6478 ( .A1(n5309), .A2(MEMORYFETCH_REG_SCAN_IN), .ZN(n5311) );
  NAND3_X1 U6479 ( .A1(n5311), .A2(n5310), .A3(n5944), .ZN(U2788) );
  XOR2_X1 U6480 ( .A(n5313), .B(n5312), .Z(n5522) );
  NOR3_X1 U6481 ( .A1(n5314), .A2(REIP_REG_30__SCAN_IN), .A3(n6512), .ZN(n5316) );
  INV_X1 U6482 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5520) );
  NOR2_X1 U6483 ( .A1(n6073), .A2(n5520), .ZN(n5315) );
  AOI211_X1 U6484 ( .C1(n6079), .C2(n5517), .A(n5316), .B(n5315), .ZN(n5318)
         );
  NAND2_X1 U6485 ( .A1(n6089), .A2(EBX_REG_30__SCAN_IN), .ZN(n5317) );
  OAI211_X1 U6486 ( .C1(n5319), .C2(n6516), .A(n5318), .B(n5317), .ZN(n5320)
         );
  AOI21_X1 U6487 ( .B1(n5400), .B2(n6088), .A(n5320), .ZN(n5321) );
  OAI21_X1 U6488 ( .B1(n5495), .B2(n6058), .A(n5321), .ZN(U2797) );
  OR2_X1 U6489 ( .A1(n5336), .A2(n5322), .ZN(n5323) );
  NAND2_X1 U6490 ( .A1(n5324), .A2(n5323), .ZN(n5640) );
  NAND2_X1 U6491 ( .A1(n5339), .A2(n5338), .ZN(n5337) );
  AOI21_X1 U6492 ( .B1(n5326), .B2(n5337), .A(n5325), .ZN(n5534) );
  NAND2_X1 U6493 ( .A1(n5534), .A2(n6032), .ZN(n5333) );
  NAND2_X1 U6494 ( .A1(n6089), .A2(EBX_REG_28__SCAN_IN), .ZN(n5329) );
  INV_X1 U6495 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6556) );
  NOR2_X1 U6496 ( .A1(n6556), .A2(REIP_REG_28__SCAN_IN), .ZN(n5327) );
  AOI22_X1 U6497 ( .A1(n6091), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .B1(n5341), 
        .B2(n5327), .ZN(n5328) );
  OAI211_X1 U6498 ( .C1(n6101), .C2(n5532), .A(n5329), .B(n5328), .ZN(n5330)
         );
  AOI21_X1 U6499 ( .B1(n5331), .B2(REIP_REG_28__SCAN_IN), .A(n5330), .ZN(n5332) );
  OAI211_X1 U6500 ( .C1(n6065), .C2(n5640), .A(n5333), .B(n5332), .ZN(U2799)
         );
  NOR2_X1 U6501 ( .A1(n4822), .A2(n5334), .ZN(n5335) );
  OR2_X1 U6502 ( .A1(n5336), .A2(n5335), .ZN(n5650) );
  OAI21_X1 U6503 ( .B1(n5339), .B2(n5338), .A(n5337), .ZN(n5540) );
  INV_X1 U6504 ( .A(n5540), .ZN(n5340) );
  NAND2_X1 U6505 ( .A1(n5340), .A2(n6032), .ZN(n5347) );
  INV_X1 U6506 ( .A(n5543), .ZN(n5344) );
  NAND2_X1 U6507 ( .A1(n6089), .A2(EBX_REG_27__SCAN_IN), .ZN(n5343) );
  AOI22_X1 U6508 ( .A1(n6091), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .B1(n5341), 
        .B2(n6556), .ZN(n5342) );
  OAI211_X1 U6509 ( .C1(n6101), .C2(n5344), .A(n5343), .B(n5342), .ZN(n5345)
         );
  AOI21_X1 U6510 ( .B1(n5353), .B2(REIP_REG_27__SCAN_IN), .A(n5345), .ZN(n5346) );
  OAI211_X1 U6511 ( .C1(n6065), .C2(n5650), .A(n5347), .B(n5346), .ZN(U2800)
         );
  NAND2_X1 U6512 ( .A1(n5404), .A2(n6032), .ZN(n5355) );
  INV_X1 U6513 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6503) );
  INV_X1 U6514 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6505) );
  OAI21_X1 U6515 ( .B1(n5362), .B2(n6503), .A(n6505), .ZN(n5352) );
  INV_X1 U6516 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5406) );
  NOR2_X1 U6517 ( .A1(n6043), .A2(n5406), .ZN(n5351) );
  OAI22_X1 U6518 ( .A1(n5349), .A2(n6073), .B1(n6101), .B2(n5348), .ZN(n5350)
         );
  AOI211_X1 U6519 ( .C1(n5353), .C2(n5352), .A(n5351), .B(n5350), .ZN(n5354)
         );
  OAI211_X1 U6520 ( .C1(n6065), .C2(n5405), .A(n5355), .B(n5354), .ZN(U2801)
         );
  AND2_X1 U6521 ( .A1(n5479), .A2(n5356), .ZN(n5359) );
  INV_X1 U6522 ( .A(n5551), .ZN(n5366) );
  NOR2_X1 U6523 ( .A1(n5360), .A2(REIP_REG_24__SCAN_IN), .ZN(n5379) );
  OAI21_X1 U6524 ( .B1(n5361), .B2(n5379), .A(REIP_REG_25__SCAN_IN), .ZN(n5365) );
  OAI22_X1 U6525 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5362), .B1(n5547), .B2(
        n6073), .ZN(n5363) );
  INV_X1 U6526 ( .A(n5363), .ZN(n5364) );
  OAI211_X1 U6527 ( .C1(n6101), .C2(n5366), .A(n5365), .B(n5364), .ZN(n5367)
         );
  AOI21_X1 U6528 ( .B1(n6089), .B2(EBX_REG_25__SCAN_IN), .A(n5367), .ZN(n5373)
         );
  AND2_X1 U6529 ( .A1(n5369), .A2(n5368), .ZN(n5370) );
  NOR2_X1 U6530 ( .A1(n5371), .A2(n5370), .ZN(n5657) );
  NAND2_X1 U6531 ( .A1(n5657), .A2(n6088), .ZN(n5372) );
  OAI211_X1 U6532 ( .C1(n5548), .C2(n6058), .A(n5373), .B(n5372), .ZN(U2802)
         );
  INV_X1 U6533 ( .A(n5374), .ZN(n5508) );
  INV_X1 U6534 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5382) );
  INV_X1 U6535 ( .A(n5375), .ZN(n5380) );
  OAI22_X1 U6536 ( .A1(n5377), .A2(n6501), .B1(n5376), .B2(n6073), .ZN(n5378)
         );
  AOI211_X1 U6537 ( .C1(n6079), .C2(n5380), .A(n5379), .B(n5378), .ZN(n5381)
         );
  OAI21_X1 U6538 ( .B1(n6043), .B2(n5382), .A(n5381), .ZN(n5383) );
  AOI21_X1 U6539 ( .B1(n5410), .B2(n6088), .A(n5383), .ZN(n5384) );
  OAI21_X1 U6540 ( .B1(n5508), .B2(n6058), .A(n5384), .ZN(U2803) );
  NAND2_X1 U6541 ( .A1(n5479), .A2(n5478), .ZN(n5480) );
  INV_X1 U6542 ( .A(n5468), .ZN(n5385) );
  AOI21_X1 U6543 ( .B1(n5386), .B2(n5480), .A(n5385), .ZN(n5616) );
  INV_X1 U6544 ( .A(n5616), .ZN(n5513) );
  NAND2_X1 U6545 ( .A1(n5485), .A2(n5387), .ZN(n5388) );
  AND2_X1 U6546 ( .A1(n5472), .A2(n5388), .ZN(n5907) );
  INV_X1 U6547 ( .A(n5389), .ZN(n5392) );
  NAND2_X1 U6548 ( .A1(n5392), .A2(n6487), .ZN(n5390) );
  NOR2_X1 U6549 ( .A1(n6090), .A2(n5390), .ZN(n5982) );
  INV_X1 U6550 ( .A(n5982), .ZN(n5391) );
  OAI21_X1 U6551 ( .B1(n5614), .B2(n6101), .A(n5391), .ZN(n5397) );
  NOR2_X1 U6552 ( .A1(n6090), .A2(n5392), .ZN(n5992) );
  INV_X1 U6553 ( .A(n5992), .ZN(n5393) );
  NAND2_X1 U6554 ( .A1(n6050), .A2(n5393), .ZN(n5994) );
  AOI22_X1 U6555 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6089), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5994), .ZN(n5394) );
  OAI211_X1 U6556 ( .C1(n6073), .C2(n5395), .A(n5394), .B(n6238), .ZN(n5396)
         );
  AOI211_X1 U6557 ( .C1(n5907), .C2(n6088), .A(n5397), .B(n5396), .ZN(n5398)
         );
  OAI21_X1 U6558 ( .B1(n5513), .B2(n6058), .A(n5398), .ZN(U2812) );
  AOI22_X1 U6559 ( .A1(n5400), .A2(n6107), .B1(EBX_REG_30__SCAN_IN), .B2(n5399), .ZN(n5401) );
  OAI21_X1 U6560 ( .B1(n5495), .B2(n5466), .A(n5401), .ZN(U2829) );
  INV_X1 U6561 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5402) );
  INV_X1 U6562 ( .A(n5534), .ZN(n5498) );
  OAI222_X1 U6563 ( .A1(n5402), .A2(n6111), .B1(n6103), .B2(n5640), .C1(n5498), 
        .C2(n5466), .ZN(U2831) );
  INV_X1 U6564 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5403) );
  OAI222_X1 U6565 ( .A1(n5403), .A2(n6111), .B1(n6103), .B2(n5650), .C1(n5540), 
        .C2(n5466), .ZN(U2832) );
  INV_X1 U6566 ( .A(n5404), .ZN(n5503) );
  OAI222_X1 U6567 ( .A1(n5406), .A2(n6111), .B1(n6103), .B2(n5405), .C1(n5503), 
        .C2(n5466), .ZN(U2833) );
  INV_X1 U6568 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5407) );
  NOR2_X1 U6569 ( .A1(n5486), .A2(n5407), .ZN(n5408) );
  AOI21_X1 U6570 ( .B1(n5657), .B2(n6107), .A(n5408), .ZN(n5409) );
  OAI21_X1 U6571 ( .B1(n5548), .B2(n5466), .A(n5409), .ZN(U2834) );
  INV_X1 U6572 ( .A(n5410), .ZN(n5411) );
  OAI222_X1 U6573 ( .A1(n6103), .A2(n5411), .B1(n5466), .B2(n5508), .C1(n5486), 
        .C2(n5382), .ZN(U2835) );
  NAND2_X1 U6574 ( .A1(n5413), .A2(n5412), .ZN(n5414) );
  INV_X1 U6575 ( .A(n5864), .ZN(n5421) );
  INV_X1 U6576 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5420) );
  NOR2_X1 U6577 ( .A1(n5417), .A2(n5416), .ZN(n5418) );
  OR2_X1 U6578 ( .A1(n5419), .A2(n5418), .ZN(n5836) );
  OAI222_X1 U6579 ( .A1(n5466), .A2(n5421), .B1(n5486), .B2(n5420), .C1(n5836), 
        .C2(n6103), .ZN(U2837) );
  INV_X1 U6580 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5423) );
  OAI222_X1 U6581 ( .A1(n5423), .A2(n5486), .B1(n6103), .B2(n5422), .C1(n5867), 
        .C2(n5466), .ZN(U2838) );
  INV_X1 U6582 ( .A(n5424), .ZN(n5428) );
  AND2_X1 U6583 ( .A1(n5479), .A2(n5425), .ZN(n5437) );
  INV_X1 U6584 ( .A(n5437), .ZN(n5427) );
  INV_X1 U6585 ( .A(n5871), .ZN(n5434) );
  INV_X1 U6586 ( .A(n5441), .ZN(n5430) );
  MUX2_X1 U6587 ( .A(n5430), .B(n5439), .S(n5429), .Z(n5432) );
  XNOR2_X1 U6588 ( .A(n5432), .B(n5431), .ZN(n5847) );
  OAI222_X1 U6589 ( .A1(n5466), .A2(n5434), .B1(n5486), .B2(n5433), .C1(n5847), 
        .C2(n6103), .ZN(U2839) );
  NAND2_X1 U6590 ( .A1(n5479), .A2(n5435), .ZN(n5448) );
  AND2_X1 U6591 ( .A1(n5448), .A2(n5436), .ZN(n5438) );
  MUX2_X1 U6592 ( .A(n5441), .B(n5440), .S(n5439), .Z(n5442) );
  INV_X1 U6593 ( .A(n5442), .ZN(n5449) );
  NAND2_X1 U6594 ( .A1(n5461), .A2(n5449), .ZN(n5451) );
  XOR2_X1 U6595 ( .A(n5443), .B(n5451), .Z(n5857) );
  INV_X1 U6596 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5444) );
  OAI222_X1 U6597 ( .A1(n5858), .A2(n5466), .B1(n6103), .B2(n5857), .C1(n5486), 
        .C2(n5444), .ZN(U2840) );
  NAND2_X1 U6598 ( .A1(n5479), .A2(n5445), .ZN(n5457) );
  NAND2_X1 U6599 ( .A1(n5457), .A2(n5446), .ZN(n5447) );
  INV_X1 U6600 ( .A(n6113), .ZN(n5454) );
  OR2_X1 U6601 ( .A1(n5461), .A2(n5449), .ZN(n5450) );
  AND2_X1 U6602 ( .A1(n5451), .A2(n5450), .ZN(n5967) );
  INV_X1 U6603 ( .A(n5967), .ZN(n5452) );
  OAI222_X1 U6604 ( .A1(n5454), .A2(n5466), .B1(n5486), .B2(n5453), .C1(n6103), 
        .C2(n5452), .ZN(U2841) );
  AND2_X1 U6605 ( .A1(n5479), .A2(n5478), .ZN(n5456) );
  OAI21_X1 U6606 ( .B1(n5467), .B2(n5458), .A(n5457), .ZN(n5976) );
  INV_X1 U6607 ( .A(n5472), .ZN(n5460) );
  AOI21_X1 U6608 ( .B1(n5460), .B2(n5470), .A(n5459), .ZN(n5462) );
  OR2_X1 U6609 ( .A1(n5462), .A2(n5461), .ZN(n5980) );
  OAI22_X1 U6610 ( .A1(n5980), .A2(n6103), .B1(n5463), .B2(n5486), .ZN(n5464)
         );
  INV_X1 U6611 ( .A(n5464), .ZN(n5465) );
  OAI21_X1 U6612 ( .B1(n5976), .B2(n5466), .A(n5465), .ZN(U2842) );
  INV_X1 U6613 ( .A(n5470), .ZN(n5471) );
  XNOR2_X1 U6614 ( .A(n5472), .B(n5471), .ZN(n5991) );
  OAI22_X1 U6615 ( .A1(n5991), .A2(n6103), .B1(n5986), .B2(n5486), .ZN(n5473)
         );
  AOI21_X1 U6616 ( .B1(n6121), .B2(n6108), .A(n5473), .ZN(n5474) );
  INV_X1 U6617 ( .A(n5474), .ZN(U2843) );
  INV_X1 U6618 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U6619 ( .A1(n5616), .A2(n6108), .ZN(n5476) );
  NAND2_X1 U6620 ( .A1(n5907), .A2(n6107), .ZN(n5475) );
  OAI211_X1 U6621 ( .C1(n5477), .C2(n5486), .A(n5476), .B(n5475), .ZN(U2844)
         );
  OR2_X1 U6622 ( .A1(n5479), .A2(n5478), .ZN(n5481) );
  OR2_X1 U6623 ( .A1(n5483), .A2(n5482), .ZN(n5484) );
  NAND2_X1 U6624 ( .A1(n5485), .A2(n5484), .ZN(n6002) );
  OAI22_X1 U6625 ( .A1(n6002), .A2(n6103), .B1(n5996), .B2(n5486), .ZN(n5487)
         );
  AOI21_X1 U6626 ( .B1(n5999), .B2(n6108), .A(n5487), .ZN(n5488) );
  INV_X1 U6627 ( .A(n5488), .ZN(U2845) );
  NAND3_X1 U6628 ( .A1(n5490), .A2(n5489), .A3(n6131), .ZN(n5492) );
  AOI22_X1 U6629 ( .A1(n6119), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6122), .ZN(n5491) );
  NAND2_X1 U6630 ( .A1(n5492), .A2(n5491), .ZN(U2860) );
  AOI22_X1 U6631 ( .A1(n6119), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6122), .ZN(n5494) );
  NAND2_X1 U6632 ( .A1(n6123), .A2(DATAI_14_), .ZN(n5493) );
  OAI211_X1 U6633 ( .C1(n5495), .C2(n5863), .A(n5494), .B(n5493), .ZN(U2861)
         );
  AOI22_X1 U6634 ( .A1(n6119), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6122), .ZN(n5497) );
  NAND2_X1 U6635 ( .A1(n6123), .A2(DATAI_12_), .ZN(n5496) );
  OAI211_X1 U6636 ( .C1(n5498), .C2(n5863), .A(n5497), .B(n5496), .ZN(U2863)
         );
  AOI22_X1 U6637 ( .A1(n6119), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6122), .ZN(n5500) );
  NAND2_X1 U6638 ( .A1(n6123), .A2(DATAI_11_), .ZN(n5499) );
  OAI211_X1 U6639 ( .C1(n5540), .C2(n5863), .A(n5500), .B(n5499), .ZN(U2864)
         );
  AOI22_X1 U6640 ( .A1(n6119), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6122), .ZN(n5502) );
  NAND2_X1 U6641 ( .A1(n6123), .A2(DATAI_10_), .ZN(n5501) );
  OAI211_X1 U6642 ( .C1(n5503), .C2(n5863), .A(n5502), .B(n5501), .ZN(U2865)
         );
  AOI22_X1 U6643 ( .A1(n6119), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6122), .ZN(n5505) );
  NAND2_X1 U6644 ( .A1(n6123), .A2(DATAI_9_), .ZN(n5504) );
  OAI211_X1 U6645 ( .C1(n5548), .C2(n5863), .A(n5505), .B(n5504), .ZN(U2866)
         );
  AOI22_X1 U6646 ( .A1(n6119), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6122), .ZN(n5507) );
  NAND2_X1 U6647 ( .A1(n6123), .A2(DATAI_8_), .ZN(n5506) );
  OAI211_X1 U6648 ( .C1(n5508), .C2(n5863), .A(n5507), .B(n5506), .ZN(U2867)
         );
  AOI22_X1 U6649 ( .A1(n6123), .A2(DATAI_3_), .B1(n6122), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U6650 ( .A1(n6119), .A2(DATAI_19_), .ZN(n5509) );
  OAI211_X1 U6651 ( .C1(n5858), .C2(n5863), .A(n5510), .B(n5509), .ZN(U2872)
         );
  AOI22_X1 U6652 ( .A1(n5511), .A2(DATAI_15_), .B1(n6122), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5512) );
  OAI21_X1 U6653 ( .B1(n5513), .B2(n5863), .A(n5512), .ZN(U2876) );
  INV_X1 U6654 ( .A(n5999), .ZN(n5516) );
  INV_X1 U6655 ( .A(DATAI_14_), .ZN(n5514) );
  OAI222_X1 U6656 ( .A1(n5516), .A2(n5863), .B1(n6131), .B2(n5515), .C1(n5514), 
        .C2(n6126), .ZN(U2877) );
  NAND2_X1 U6657 ( .A1(n6204), .A2(n5517), .ZN(n5519) );
  OAI211_X1 U6658 ( .C1(n5520), .C2(n6208), .A(n5519), .B(n5518), .ZN(n5521)
         );
  AOI21_X1 U6659 ( .B1(n5522), .B2(n6219), .A(n5521), .ZN(n5523) );
  OAI21_X1 U6660 ( .B1(n5524), .B2(n6195), .A(n5523), .ZN(U2956) );
  INV_X1 U6661 ( .A(n5525), .ZN(n5526) );
  NAND3_X1 U6662 ( .A1(n5526), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n2996), .ZN(n5529) );
  INV_X1 U6663 ( .A(n5545), .ZN(n5528) );
  NAND3_X1 U6664 ( .A1(n5528), .A2(n5241), .A3(n5527), .ZN(n5536) );
  AOI22_X1 U6665 ( .A1(n5529), .A2(n5536), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n6567), .ZN(n5530) );
  XNOR2_X1 U6666 ( .A(n5530), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5648)
         );
  INV_X1 U6667 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6510) );
  NOR2_X1 U6668 ( .A1(n6238), .A2(n6510), .ZN(n5642) );
  AOI21_X1 U6669 ( .B1(n6218), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5642), 
        .ZN(n5531) );
  OAI21_X1 U6670 ( .B1(n5532), .B2(n6225), .A(n5531), .ZN(n5533) );
  AOI21_X1 U6671 ( .B1(n5534), .B2(n6219), .A(n5533), .ZN(n5535) );
  OAI21_X1 U6672 ( .B1(n6195), .B2(n5648), .A(n5535), .ZN(U2958) );
  NAND2_X1 U6673 ( .A1(n5537), .A2(n5536), .ZN(n5538) );
  XNOR2_X1 U6674 ( .A(n5538), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5656)
         );
  NAND2_X1 U6675 ( .A1(n2997), .A2(REIP_REG_27__SCAN_IN), .ZN(n5649) );
  OAI21_X1 U6676 ( .B1(n6208), .B2(n5539), .A(n5649), .ZN(n5542) );
  NOR2_X1 U6677 ( .A1(n5540), .A2(n6194), .ZN(n5541) );
  AOI211_X1 U6678 ( .C1(n6204), .C2(n5543), .A(n5542), .B(n5541), .ZN(n5544)
         );
  OAI21_X1 U6679 ( .B1(n5656), .B2(n6195), .A(n5544), .ZN(U2959) );
  AOI21_X1 U6680 ( .B1(n5546), .B2(n5545), .A(n3012), .ZN(n5664) );
  NAND2_X1 U6681 ( .A1(n2997), .A2(REIP_REG_25__SCAN_IN), .ZN(n5659) );
  OAI21_X1 U6682 ( .B1(n6208), .B2(n5547), .A(n5659), .ZN(n5550) );
  NOR2_X1 U6683 ( .A1(n5548), .A2(n6194), .ZN(n5549) );
  AOI211_X1 U6684 ( .C1(n6204), .C2(n5551), .A(n5550), .B(n5549), .ZN(n5552)
         );
  OAI21_X1 U6685 ( .B1(n5664), .B2(n6195), .A(n5552), .ZN(U2961) );
  NAND3_X1 U6686 ( .A1(n2996), .A2(n5694), .A3(n5676), .ZN(n5554) );
  OAI21_X1 U6687 ( .B1(n5555), .B2(n5554), .A(n5553), .ZN(n5556) );
  XNOR2_X1 U6688 ( .A(n5556), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5673)
         );
  NAND2_X1 U6689 ( .A1(n2997), .A2(REIP_REG_23__SCAN_IN), .ZN(n5666) );
  OAI21_X1 U6690 ( .B1(n6208), .B2(n5557), .A(n5666), .ZN(n5560) );
  NOR2_X1 U6691 ( .A1(n5558), .A2(n6194), .ZN(n5559) );
  AOI211_X1 U6692 ( .C1(n6204), .C2(n5561), .A(n5560), .B(n5559), .ZN(n5562)
         );
  OAI21_X1 U6693 ( .B1(n5673), .B2(n6195), .A(n5562), .ZN(U2963) );
  AOI21_X1 U6694 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n2996), .A(n5563), 
        .ZN(n5565) );
  XOR2_X1 U6695 ( .A(n5565), .B(n5564), .Z(n5681) );
  NAND2_X1 U6696 ( .A1(n2997), .A2(REIP_REG_22__SCAN_IN), .ZN(n5674) );
  OR2_X1 U6697 ( .A1(n6208), .A2(n5566), .ZN(n5567) );
  OAI211_X1 U6698 ( .C1(n6225), .C2(n5835), .A(n5674), .B(n5567), .ZN(n5568)
         );
  AOI21_X1 U6699 ( .B1(n5864), .B2(n6219), .A(n5568), .ZN(n5569) );
  OAI21_X1 U6700 ( .B1(n5681), .B2(n6195), .A(n5569), .ZN(U2964) );
  NAND2_X1 U6701 ( .A1(n5571), .A2(n5570), .ZN(n5573) );
  AOI21_X1 U6702 ( .B1(n5574), .B2(n5573), .A(n5572), .ZN(n5691) );
  NAND2_X1 U6703 ( .A1(n2997), .A2(REIP_REG_21__SCAN_IN), .ZN(n5685) );
  OAI21_X1 U6704 ( .B1(n6208), .B2(n5575), .A(n5685), .ZN(n5577) );
  NOR2_X1 U6705 ( .A1(n5867), .A2(n6194), .ZN(n5576) );
  OAI21_X1 U6706 ( .B1(n5691), .B2(n6195), .A(n5579), .ZN(U2965) );
  XNOR2_X1 U6707 ( .A(n2996), .B(n5580), .ZN(n5581) );
  XNOR2_X1 U6708 ( .A(n5582), .B(n5581), .ZN(n5699) );
  INV_X1 U6709 ( .A(n5849), .ZN(n5584) );
  NAND2_X1 U6710 ( .A1(n2997), .A2(REIP_REG_20__SCAN_IN), .ZN(n5692) );
  NAND2_X1 U6711 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5583)
         );
  OAI211_X1 U6712 ( .C1(n6225), .C2(n5584), .A(n5692), .B(n5583), .ZN(n5585)
         );
  AOI21_X1 U6713 ( .B1(n5871), .B2(n6219), .A(n5585), .ZN(n5586) );
  OAI21_X1 U6714 ( .B1(n6195), .B2(n5699), .A(n5586), .ZN(U2966) );
  XOR2_X1 U6715 ( .A(n5588), .B(n5587), .Z(n5707) );
  NAND2_X1 U6716 ( .A1(n2997), .A2(REIP_REG_19__SCAN_IN), .ZN(n5701) );
  OAI21_X1 U6717 ( .B1(n6208), .B2(n6553), .A(n5701), .ZN(n5590) );
  NOR2_X1 U6718 ( .A1(n5858), .A2(n6194), .ZN(n5589) );
  AOI211_X1 U6719 ( .C1(n6204), .C2(n5860), .A(n5590), .B(n5589), .ZN(n5591)
         );
  OAI21_X1 U6720 ( .B1(n5707), .B2(n6195), .A(n5591), .ZN(U2967) );
  NAND2_X1 U6721 ( .A1(n2996), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5875) );
  INV_X1 U6722 ( .A(n5597), .ZN(n5876) );
  NAND2_X1 U6723 ( .A1(n5876), .A2(n5602), .ZN(n5593) );
  OAI211_X1 U6724 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n2996), .A(n5593), .B(n5875), .ZN(n5596) );
  NOR4_X1 U6725 ( .A1(n2996), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A4(INSTADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n5595) );
  NAND2_X1 U6726 ( .A1(n5612), .A2(n5595), .ZN(n5874) );
  OAI211_X1 U6727 ( .C1(n5597), .C2(n5875), .A(n5596), .B(n5874), .ZN(n5708)
         );
  NAND2_X1 U6728 ( .A1(n5708), .A2(n6221), .ZN(n5600) );
  NAND2_X1 U6729 ( .A1(n2997), .A2(REIP_REG_17__SCAN_IN), .ZN(n5711) );
  OAI21_X1 U6730 ( .B1(n6208), .B2(n5972), .A(n5711), .ZN(n5598) );
  AOI21_X1 U6731 ( .B1(n5977), .B2(n6204), .A(n5598), .ZN(n5599) );
  OAI211_X1 U6732 ( .C1(n6194), .C2(n5976), .A(n5600), .B(n5599), .ZN(U2969)
         );
  INV_X1 U6733 ( .A(n5602), .ZN(n5605) );
  AND2_X1 U6734 ( .A1(n5602), .A2(n5601), .ZN(n5603) );
  OAI22_X1 U6735 ( .A1(n5876), .A2(n5605), .B1(n5604), .B2(n5603), .ZN(n5901)
         );
  AOI22_X1 U6736 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n2997), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5606) );
  OAI21_X1 U6737 ( .B1(n5607), .B2(n6225), .A(n5606), .ZN(n5608) );
  AOI21_X1 U6738 ( .B1(n6121), .B2(n6219), .A(n5608), .ZN(n5609) );
  OAI21_X1 U6739 ( .B1(n5901), .B2(n6195), .A(n5609), .ZN(U2970) );
  XNOR2_X1 U6740 ( .A(n2996), .B(n5610), .ZN(n5611) );
  XNOR2_X1 U6741 ( .A(n5612), .B(n5611), .ZN(n5906) );
  AOI22_X1 U6742 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n2997), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5613) );
  OAI21_X1 U6743 ( .B1(n5614), .B2(n6225), .A(n5613), .ZN(n5615) );
  AOI21_X1 U6744 ( .B1(n5616), .B2(n6219), .A(n5615), .ZN(n5617) );
  OAI21_X1 U6745 ( .B1(n6195), .B2(n5906), .A(n5617), .ZN(U2971) );
  XNOR2_X1 U6746 ( .A(n2996), .B(n5914), .ZN(n5619) );
  XNOR2_X1 U6747 ( .A(n5618), .B(n5619), .ZN(n5919) );
  INV_X1 U6748 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5621) );
  INV_X1 U6749 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5620) );
  OAI22_X1 U6750 ( .A1(n6208), .A2(n5621), .B1(n6238), .B2(n5620), .ZN(n5622)
         );
  AOI21_X1 U6751 ( .B1(n6204), .B2(n5998), .A(n5622), .ZN(n5624) );
  NAND2_X1 U6752 ( .A1(n5999), .A2(n6219), .ZN(n5623) );
  OAI211_X1 U6753 ( .C1(n5919), .C2(n6195), .A(n5624), .B(n5623), .ZN(U2972)
         );
  NAND2_X1 U6754 ( .A1(n5625), .A2(n6219), .ZN(n5630) );
  OR2_X1 U6755 ( .A1(n5626), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6299)
         );
  NAND3_X1 U6756 ( .A1(n6299), .A2(n6221), .A3(n6297), .ZN(n5629) );
  NAND2_X1 U6757 ( .A1(n2997), .A2(REIP_REG_0__SCAN_IN), .ZN(n6300) );
  OAI21_X1 U6758 ( .B1(n6218), .B2(n5627), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5628) );
  NAND4_X1 U6759 ( .A1(n5630), .A2(n5629), .A3(n6300), .A4(n5628), .ZN(U2986)
         );
  INV_X1 U6760 ( .A(n5631), .ZN(n5637) );
  OAI21_X1 U6761 ( .B1(n5651), .B2(n5643), .A(n5632), .ZN(n5636) );
  OAI21_X1 U6762 ( .B1(n5634), .B2(n6303), .A(n5633), .ZN(n5635) );
  AOI21_X1 U6763 ( .B1(n5637), .B2(n5636), .A(n5635), .ZN(n5638) );
  OAI21_X1 U6764 ( .B1(n5639), .B2(n6269), .A(n5638), .ZN(U2989) );
  NOR2_X1 U6765 ( .A1(n5640), .A2(n6303), .ZN(n5641) );
  AOI211_X1 U6766 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n5654), .A(n5642), .B(n5641), .ZN(n5647) );
  INV_X1 U6767 ( .A(n5643), .ZN(n5644) );
  OR3_X1 U6768 ( .A1(n5651), .A2(n5645), .A3(n5644), .ZN(n5646) );
  OAI211_X1 U6769 ( .C1(n5648), .C2(n6269), .A(n5647), .B(n5646), .ZN(U2990)
         );
  OAI21_X1 U6770 ( .B1(n5650), .B2(n6303), .A(n5649), .ZN(n5653) );
  NOR2_X1 U6771 ( .A1(n5651), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5652)
         );
  AOI211_X1 U6772 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5654), .A(n5653), .B(n5652), .ZN(n5655) );
  OAI21_X1 U6773 ( .B1(n5656), .B2(n6269), .A(n5655), .ZN(U2991) );
  NAND2_X1 U6774 ( .A1(n5657), .A2(n6288), .ZN(n5658) );
  OAI211_X1 U6775 ( .C1(n5660), .C2(n6649), .A(n5659), .B(n5658), .ZN(n5661)
         );
  AOI21_X1 U6776 ( .B1(n5662), .B2(n6649), .A(n5661), .ZN(n5663) );
  OAI21_X1 U6777 ( .B1(n5664), .B2(n6269), .A(n5663), .ZN(U2993) );
  INV_X1 U6778 ( .A(n5665), .ZN(n5671) );
  OAI21_X1 U6779 ( .B1(n5667), .B2(n6303), .A(n5666), .ZN(n5670) );
  NOR2_X1 U6780 ( .A1(n5668), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5669)
         );
  AOI211_X1 U6781 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5671), .A(n5670), .B(n5669), .ZN(n5672) );
  OAI21_X1 U6782 ( .B1(n5673), .B2(n6269), .A(n5672), .ZN(U2995) );
  INV_X1 U6783 ( .A(n5686), .ZN(n5679) );
  OAI21_X1 U6784 ( .B1(n5836), .B2(n6303), .A(n5674), .ZN(n5678) );
  NOR3_X1 U6785 ( .A1(n5682), .A2(n5676), .A3(n5675), .ZN(n5677) );
  AOI211_X1 U6786 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5679), .A(n5678), .B(n5677), .ZN(n5680) );
  OAI21_X1 U6787 ( .B1(n5681), .B2(n6269), .A(n5680), .ZN(U2996) );
  INV_X1 U6788 ( .A(n5682), .ZN(n5689) );
  NAND2_X1 U6789 ( .A1(n5683), .A2(n6288), .ZN(n5684) );
  OAI211_X1 U6790 ( .C1(n5686), .C2(n5688), .A(n5685), .B(n5684), .ZN(n5687)
         );
  AOI21_X1 U6791 ( .B1(n5689), .B2(n5688), .A(n5687), .ZN(n5690) );
  OAI21_X1 U6792 ( .B1(n5691), .B2(n6269), .A(n5690), .ZN(U2997) );
  NOR2_X1 U6793 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5891), .ZN(n5709)
         );
  NOR2_X1 U6794 ( .A1(n5713), .A2(n5709), .ZN(n5897) );
  OAI21_X1 U6795 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5899), .A(n5897), 
        .ZN(n5700) );
  OAI21_X1 U6796 ( .B1(n5847), .B2(n6303), .A(n5692), .ZN(n5697) );
  INV_X1 U6797 ( .A(n5705), .ZN(n5695) );
  NOR3_X1 U6798 ( .A1(n5695), .A2(n5694), .A3(n5693), .ZN(n5696) );
  AOI211_X1 U6799 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n5700), .A(n5697), .B(n5696), .ZN(n5698) );
  OAI21_X1 U6800 ( .B1(n5699), .B2(n6269), .A(n5698), .ZN(U2998) );
  NAND2_X1 U6801 ( .A1(n5700), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5702) );
  OAI211_X1 U6802 ( .C1(n5857), .C2(n6303), .A(n5702), .B(n5701), .ZN(n5703)
         );
  AOI21_X1 U6803 ( .B1(n5705), .B2(n5704), .A(n5703), .ZN(n5706) );
  OAI21_X1 U6804 ( .B1(n5707), .B2(n6269), .A(n5706), .ZN(U2999) );
  INV_X1 U6805 ( .A(n5708), .ZN(n5715) );
  INV_X1 U6806 ( .A(n5709), .ZN(n5710) );
  OAI211_X1 U6807 ( .C1(n5980), .C2(n6303), .A(n5711), .B(n5710), .ZN(n5712)
         );
  AOI21_X1 U6808 ( .B1(n5713), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5712), 
        .ZN(n5714) );
  OAI21_X1 U6809 ( .B1(n5715), .B2(n6269), .A(n5714), .ZN(U3001) );
  NOR2_X1 U6810 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5716), .ZN(n5726)
         );
  AOI21_X1 U6811 ( .B1(n5717), .B2(n5761), .A(n6538), .ZN(n5719) );
  NOR2_X1 U6812 ( .A1(n5719), .A2(n5718), .ZN(n5722) );
  AOI211_X1 U6813 ( .C1(n5723), .C2(n5722), .A(n5721), .B(n5720), .ZN(n5724)
         );
  NAND2_X1 U6814 ( .A1(n5754), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5733) );
  INV_X1 U6815 ( .A(n5726), .ZN(n5756) );
  AOI22_X1 U6816 ( .A1(n5730), .A2(n5729), .B1(n5728), .B2(n5727), .ZN(n5755)
         );
  OAI22_X1 U6817 ( .A1(n5776), .A2(n5756), .B1(n5755), .B2(n5781), .ZN(n5731)
         );
  AOI21_X1 U6818 ( .B1(n6353), .B2(n5758), .A(n5731), .ZN(n5732) );
  OAI211_X1 U6819 ( .C1(n6358), .C2(n5761), .A(n5733), .B(n5732), .ZN(U3052)
         );
  NAND2_X1 U6820 ( .A1(n5754), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5736) );
  OAI22_X1 U6821 ( .A1(n5783), .A2(n5756), .B1(n5755), .B2(n5788), .ZN(n5734)
         );
  AOI21_X1 U6822 ( .B1(n6311), .B2(n5758), .A(n5734), .ZN(n5735) );
  OAI211_X1 U6823 ( .C1(n5761), .C2(n6316), .A(n5736), .B(n5735), .ZN(U3053)
         );
  NAND2_X1 U6824 ( .A1(n5754), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5739) );
  OAI22_X1 U6825 ( .A1(n5790), .A2(n5756), .B1(n5755), .B2(n5795), .ZN(n5737)
         );
  AOI21_X1 U6826 ( .B1(n6334), .B2(n5758), .A(n5737), .ZN(n5738) );
  OAI211_X1 U6827 ( .C1(n5761), .C2(n6339), .A(n5739), .B(n5738), .ZN(U3054)
         );
  NAND2_X1 U6828 ( .A1(n5754), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5743) );
  OAI22_X1 U6829 ( .A1(n5797), .A2(n5756), .B1(n5755), .B2(n5802), .ZN(n5740)
         );
  AOI21_X1 U6830 ( .B1(n5741), .B2(n5758), .A(n5740), .ZN(n5742) );
  OAI211_X1 U6831 ( .C1(n5761), .C2(n5744), .A(n5743), .B(n5742), .ZN(U3055)
         );
  NAND2_X1 U6832 ( .A1(n5754), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5747) );
  OAI22_X1 U6833 ( .A1(n5804), .A2(n5756), .B1(n5755), .B2(n5809), .ZN(n5745)
         );
  AOI21_X1 U6834 ( .B1(n6359), .B2(n5758), .A(n5745), .ZN(n5746) );
  OAI211_X1 U6835 ( .C1(n5761), .C2(n6364), .A(n5747), .B(n5746), .ZN(U3056)
         );
  NAND2_X1 U6836 ( .A1(n5754), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5750) );
  OAI22_X1 U6837 ( .A1(n5811), .A2(n5756), .B1(n5755), .B2(n5816), .ZN(n5748)
         );
  AOI21_X1 U6838 ( .B1(n6365), .B2(n5758), .A(n5748), .ZN(n5749) );
  OAI211_X1 U6839 ( .C1(n5761), .C2(n6370), .A(n5750), .B(n5749), .ZN(U3057)
         );
  NAND2_X1 U6840 ( .A1(n5754), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5753) );
  OAI22_X1 U6841 ( .A1(n5818), .A2(n5756), .B1(n5755), .B2(n5823), .ZN(n5751)
         );
  AOI21_X1 U6842 ( .B1(n6371), .B2(n5758), .A(n5751), .ZN(n5752) );
  OAI211_X1 U6843 ( .C1(n5761), .C2(n6376), .A(n5753), .B(n5752), .ZN(U3058)
         );
  NAND2_X1 U6844 ( .A1(n5754), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5760) );
  OAI22_X1 U6845 ( .A1(n5827), .A2(n5756), .B1(n5755), .B2(n5833), .ZN(n5757)
         );
  AOI21_X1 U6846 ( .B1(n6378), .B2(n5758), .A(n5757), .ZN(n5759) );
  OAI211_X1 U6847 ( .C1(n5761), .C2(n6387), .A(n5760), .B(n5759), .ZN(U3059)
         );
  INV_X1 U6848 ( .A(n5830), .ZN(n5762) );
  NAND2_X1 U6849 ( .A1(n5762), .A2(n6386), .ZN(n5764) );
  AOI21_X1 U6850 ( .B1(n5764), .B2(STATEBS16_REG_SCAN_IN), .A(n5763), .ZN(
        n5772) );
  NOR2_X1 U6851 ( .A1(n5766), .A2(n5765), .ZN(n5767) );
  AOI22_X1 U6852 ( .A1(n5772), .A2(n5769), .B1(n5768), .B2(n5767), .ZN(n5834)
         );
  INV_X1 U6853 ( .A(n5769), .ZN(n5771) );
  OR2_X1 U6854 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5770), .ZN(n5826)
         );
  AOI22_X1 U6855 ( .A1(n5772), .A2(n5771), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5826), .ZN(n5773) );
  OAI211_X1 U6856 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6532), .A(n5774), .B(n5773), .ZN(n5824) );
  NAND2_X1 U6857 ( .A1(n5824), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5780)
         );
  OAI22_X1 U6858 ( .A1(n5776), .A2(n5826), .B1(n6386), .B2(n5775), .ZN(n5777)
         );
  AOI21_X1 U6859 ( .B1(n5830), .B2(n5778), .A(n5777), .ZN(n5779) );
  OAI211_X1 U6860 ( .C1(n5834), .C2(n5781), .A(n5780), .B(n5779), .ZN(U3100)
         );
  NAND2_X1 U6861 ( .A1(n5824), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5787)
         );
  OAI22_X1 U6862 ( .A1(n5783), .A2(n5826), .B1(n6386), .B2(n5782), .ZN(n5784)
         );
  AOI21_X1 U6863 ( .B1(n5830), .B2(n5785), .A(n5784), .ZN(n5786) );
  OAI211_X1 U6864 ( .C1(n5834), .C2(n5788), .A(n5787), .B(n5786), .ZN(U3101)
         );
  NAND2_X1 U6865 ( .A1(n5824), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5794)
         );
  OAI22_X1 U6866 ( .A1(n5790), .A2(n5826), .B1(n6386), .B2(n5789), .ZN(n5791)
         );
  AOI21_X1 U6867 ( .B1(n5830), .B2(n5792), .A(n5791), .ZN(n5793) );
  OAI211_X1 U6868 ( .C1(n5834), .C2(n5795), .A(n5794), .B(n5793), .ZN(U3102)
         );
  NAND2_X1 U6869 ( .A1(n5824), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5801)
         );
  OAI22_X1 U6870 ( .A1(n5797), .A2(n5826), .B1(n6386), .B2(n5796), .ZN(n5798)
         );
  AOI21_X1 U6871 ( .B1(n5830), .B2(n5799), .A(n5798), .ZN(n5800) );
  OAI211_X1 U6872 ( .C1(n5834), .C2(n5802), .A(n5801), .B(n5800), .ZN(U3103)
         );
  NAND2_X1 U6873 ( .A1(n5824), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5808)
         );
  OAI22_X1 U6874 ( .A1(n5804), .A2(n5826), .B1(n6386), .B2(n5803), .ZN(n5805)
         );
  AOI21_X1 U6875 ( .B1(n5830), .B2(n5806), .A(n5805), .ZN(n5807) );
  OAI211_X1 U6876 ( .C1(n5834), .C2(n5809), .A(n5808), .B(n5807), .ZN(U3104)
         );
  NAND2_X1 U6877 ( .A1(n5824), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5815)
         );
  OAI22_X1 U6878 ( .A1(n5811), .A2(n5826), .B1(n6386), .B2(n5810), .ZN(n5812)
         );
  AOI21_X1 U6879 ( .B1(n5830), .B2(n5813), .A(n5812), .ZN(n5814) );
  OAI211_X1 U6880 ( .C1(n5834), .C2(n5816), .A(n5815), .B(n5814), .ZN(U3105)
         );
  NAND2_X1 U6881 ( .A1(n5824), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5822)
         );
  OAI22_X1 U6882 ( .A1(n5818), .A2(n5826), .B1(n6386), .B2(n5817), .ZN(n5819)
         );
  AOI21_X1 U6883 ( .B1(n5830), .B2(n5820), .A(n5819), .ZN(n5821) );
  OAI211_X1 U6884 ( .C1(n5834), .C2(n5823), .A(n5822), .B(n5821), .ZN(U3106)
         );
  NAND2_X1 U6885 ( .A1(n5824), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5832)
         );
  OAI22_X1 U6886 ( .A1(n5827), .A2(n5826), .B1(n6386), .B2(n5825), .ZN(n5828)
         );
  AOI21_X1 U6887 ( .B1(n5830), .B2(n5829), .A(n5828), .ZN(n5831) );
  OAI211_X1 U6888 ( .C1(n5834), .C2(n5833), .A(n5832), .B(n5831), .ZN(U3107)
         );
  AND2_X1 U6889 ( .A1(n6156), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6890 ( .A1(EBX_REG_22__SCAN_IN), .A2(n6089), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6091), .ZN(n5845) );
  OAI22_X1 U6891 ( .A1(n5836), .A2(n6065), .B1(n5835), .B2(n6101), .ZN(n5837)
         );
  AOI21_X1 U6892 ( .B1(n5864), .B2(n6032), .A(n5837), .ZN(n5844) );
  OAI21_X1 U6893 ( .B1(n5839), .B2(n5838), .A(REIP_REG_22__SCAN_IN), .ZN(n5843) );
  OR3_X1 U6894 ( .A1(n5841), .A2(n5840), .A3(REIP_REG_22__SCAN_IN), .ZN(n5842)
         );
  NAND4_X1 U6895 ( .A1(n5845), .A2(n5844), .A3(n5843), .A4(n5842), .ZN(U2805)
         );
  AOI21_X1 U6896 ( .B1(n5846), .B2(n5964), .A(REIP_REG_20__SCAN_IN), .ZN(n5852) );
  AOI22_X1 U6897 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6089), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6091), .ZN(n5851) );
  INV_X1 U6898 ( .A(n5847), .ZN(n5848) );
  AOI222_X1 U6899 ( .A1(n5871), .A2(n6032), .B1(n5849), .B2(n6079), .C1(n6088), 
        .C2(n5848), .ZN(n5850) );
  OAI211_X1 U6900 ( .C1(n5853), .C2(n5852), .A(n5851), .B(n5850), .ZN(U2807)
         );
  OAI211_X1 U6901 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n5964), .B(n5854), .ZN(n5855) );
  OAI211_X1 U6902 ( .C1(n6073), .C2(n6553), .A(n5855), .B(n6238), .ZN(n5856)
         );
  AOI21_X1 U6903 ( .B1(EBX_REG_19__SCAN_IN), .B2(n6089), .A(n5856), .ZN(n5862)
         );
  OAI22_X1 U6904 ( .A1(n5858), .A2(n6058), .B1(n5857), .B2(n6065), .ZN(n5859)
         );
  AOI21_X1 U6905 ( .B1(n5860), .B2(n6079), .A(n5859), .ZN(n5861) );
  OAI211_X1 U6906 ( .C1(n5973), .C2(n6495), .A(n5862), .B(n5861), .ZN(U2808)
         );
  INV_X1 U6907 ( .A(n5863), .ZN(n6120) );
  AOI22_X1 U6908 ( .A1(n5864), .A2(n6120), .B1(n6119), .B2(DATAI_22_), .ZN(
        n5866) );
  AOI22_X1 U6909 ( .A1(n6123), .A2(DATAI_6_), .B1(n6122), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5865) );
  NAND2_X1 U6910 ( .A1(n5866), .A2(n5865), .ZN(U2869) );
  INV_X1 U6911 ( .A(n5867), .ZN(n5868) );
  AOI22_X1 U6912 ( .A1(n5868), .A2(n6120), .B1(n6119), .B2(DATAI_21_), .ZN(
        n5870) );
  AOI22_X1 U6913 ( .A1(n6123), .A2(DATAI_5_), .B1(n6122), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U6914 ( .A1(n5870), .A2(n5869), .ZN(U2870) );
  AOI22_X1 U6915 ( .A1(n5871), .A2(n6120), .B1(n6119), .B2(DATAI_20_), .ZN(
        n5873) );
  AOI22_X1 U6916 ( .A1(n6123), .A2(DATAI_4_), .B1(n6122), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U6917 ( .A1(n5873), .A2(n5872), .ZN(U2871) );
  AOI22_X1 U6918 ( .A1(n2997), .A2(REIP_REG_18__SCAN_IN), .B1(n6218), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5879) );
  OAI21_X1 U6919 ( .B1(n5876), .B2(n5875), .A(n5874), .ZN(n5877) );
  XOR2_X1 U6920 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .B(n5877), .Z(n5893) );
  AOI22_X1 U6921 ( .A1(n5893), .A2(n6221), .B1(n6219), .B2(n6113), .ZN(n5878)
         );
  OAI211_X1 U6922 ( .C1(n6225), .C2(n5970), .A(n5879), .B(n5878), .ZN(U2968)
         );
  NAND2_X1 U6923 ( .A1(n5881), .A2(n5880), .ZN(n5884) );
  NAND2_X1 U6924 ( .A1(n5884), .A2(n5882), .ZN(n5888) );
  NAND2_X1 U6925 ( .A1(n5884), .A2(n5883), .ZN(n5886) );
  NAND2_X1 U6926 ( .A1(n5886), .A2(n5885), .ZN(n5887) );
  NAND2_X1 U6927 ( .A1(n5888), .A2(n5887), .ZN(n5925) );
  OAI22_X1 U6928 ( .A1(n6128), .A2(n6194), .B1(n6009), .B2(n6225), .ZN(n5889)
         );
  AOI21_X1 U6929 ( .B1(n6221), .B2(n5925), .A(n5889), .ZN(n5890) );
  NAND2_X1 U6930 ( .A1(n2997), .A2(REIP_REG_13__SCAN_IN), .ZN(n5930) );
  OAI211_X1 U6931 ( .C1(n6006), .C2(n6208), .A(n5890), .B(n5930), .ZN(U2973)
         );
  INV_X1 U6932 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5896) );
  INV_X1 U6933 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6641) );
  NOR3_X1 U6934 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6641), .A3(n5891), 
        .ZN(n5892) );
  AOI21_X1 U6935 ( .B1(REIP_REG_18__SCAN_IN), .B2(n2997), .A(n5892), .ZN(n5895) );
  AOI22_X1 U6936 ( .A1(n5893), .A2(n6298), .B1(n6288), .B2(n5967), .ZN(n5894)
         );
  OAI211_X1 U6937 ( .C1(n5897), .C2(n5896), .A(n5895), .B(n5894), .ZN(U3000)
         );
  INV_X1 U6938 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6490) );
  INV_X1 U6939 ( .A(n5898), .ZN(n5900) );
  OAI21_X1 U6940 ( .B1(n5900), .B2(n5899), .A(n6233), .ZN(n5910) );
  OAI22_X1 U6941 ( .A1(n5901), .A2(n6269), .B1(n5991), .B2(n6303), .ZN(n5902)
         );
  AOI21_X1 U6942 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n5910), .A(n5902), 
        .ZN(n5905) );
  OAI211_X1 U6943 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5911), .B(n5903), .ZN(n5904) );
  OAI211_X1 U6944 ( .C1(n6490), .C2(n6238), .A(n5905), .B(n5904), .ZN(U3002)
         );
  INV_X1 U6945 ( .A(n5906), .ZN(n5908) );
  AOI22_X1 U6946 ( .A1(n5908), .A2(n6298), .B1(n6288), .B2(n5907), .ZN(n5913)
         );
  NOR2_X1 U6947 ( .A1(n6238), .A2(n6487), .ZN(n5909) );
  AOI221_X1 U6948 ( .B1(n5911), .B2(n5610), .C1(n5910), .C2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5909), .ZN(n5912) );
  NAND2_X1 U6949 ( .A1(n5913), .A2(n5912), .ZN(U3003) );
  NAND2_X1 U6950 ( .A1(n5918), .A2(n5914), .ZN(n5923) );
  NOR3_X1 U6951 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5915), .A3(n5924), 
        .ZN(n5927) );
  AOI21_X1 U6952 ( .B1(n5924), .B2(n5916), .A(n5927), .ZN(n5917) );
  OAI211_X1 U6953 ( .C1(n5918), .C2(n6308), .A(n5917), .B(n6233), .ZN(n5929)
         );
  OAI22_X1 U6954 ( .A1(n5919), .A2(n6269), .B1(n6303), .B2(n6002), .ZN(n5920)
         );
  AOI21_X1 U6955 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n5929), .A(n5920), 
        .ZN(n5922) );
  NAND2_X1 U6956 ( .A1(n2997), .A2(REIP_REG_14__SCAN_IN), .ZN(n5921) );
  OAI211_X1 U6957 ( .C1(n6226), .C2(n5923), .A(n5922), .B(n5921), .ZN(U3004)
         );
  OR2_X1 U6958 ( .A1(n5924), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5933)
         );
  INV_X1 U6959 ( .A(n5925), .ZN(n5926) );
  OAI22_X1 U6960 ( .A1(n5926), .A2(n6269), .B1(n6303), .B2(n6013), .ZN(n5928)
         );
  AOI211_X1 U6961 ( .C1(n5929), .C2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(n5928), .B(n5927), .ZN(n5931) );
  OAI211_X1 U6962 ( .C1(n5933), .C2(n5932), .A(n5931), .B(n5930), .ZN(U3005)
         );
  INV_X1 U6963 ( .A(n5934), .ZN(n5937) );
  NAND4_X1 U6964 ( .A1(n6072), .A2(n5937), .A3(n5936), .A4(n5935), .ZN(n5938)
         );
  OAI21_X1 U6965 ( .B1(n5940), .B2(n5939), .A(n5938), .ZN(U3455) );
  INV_X1 U6966 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6464) );
  INV_X1 U6967 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6450) );
  AOI21_X1 U6968 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6464), .A(n6450), .ZN(n5946) );
  INV_X1 U6969 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5941) );
  NAND2_X1 U6970 ( .A1(n6450), .A2(STATE_REG_1__SCAN_IN), .ZN(n6531) );
  INV_X1 U6971 ( .A(n6531), .ZN(n6504) );
  AOI21_X1 U6972 ( .B1(n5946), .B2(n5941), .A(n6504), .ZN(U2789) );
  OAI21_X1 U6973 ( .B1(n5942), .B2(n6432), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5943) );
  OAI21_X1 U6974 ( .B1(n5944), .B2(n6540), .A(n5943), .ZN(U2790) );
  NOR2_X1 U6975 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5947) );
  INV_X1 U6976 ( .A(n6504), .ZN(n6550) );
  OAI21_X1 U6977 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5947), .A(n6550), .ZN(n5945)
         );
  OAI21_X1 U6978 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6531), .A(n5945), .ZN(
        U2791) );
  NOR2_X1 U6979 ( .A1(n6504), .A2(n5946), .ZN(n6520) );
  OAI21_X1 U6980 ( .B1(n5947), .B2(BS16_N), .A(n6520), .ZN(n6518) );
  OAI21_X1 U6981 ( .B1(n6520), .B2(n6538), .A(n6518), .ZN(U2792) );
  OAI21_X1 U6982 ( .B1(n5949), .B2(n5948), .A(n6195), .ZN(U2793) );
  NOR4_X1 U6983 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n5953) );
  NOR4_X1 U6984 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n5952) );
  NOR4_X1 U6985 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n5951) );
  NOR4_X1 U6986 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_22__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n5950) );
  NAND4_X1 U6987 ( .A1(n5953), .A2(n5952), .A3(n5951), .A4(n5950), .ZN(n5959)
         );
  NOR4_X1 U6988 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(n5957) );
  AOI211_X1 U6989 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_26__SCAN_IN), .B(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n5956) );
  NOR4_X1 U6990 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(n5955)
         );
  NOR4_X1 U6991 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n5954) );
  NAND4_X1 U6992 ( .A1(n5957), .A2(n5956), .A3(n5955), .A4(n5954), .ZN(n5958)
         );
  NOR2_X1 U6993 ( .A1(n5959), .A2(n5958), .ZN(n6529) );
  INV_X1 U6994 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5961) );
  NOR3_X1 U6995 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5962) );
  OAI21_X1 U6996 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5962), .A(n6529), .ZN(n5960)
         );
  OAI21_X1 U6997 ( .B1(n6529), .B2(n5961), .A(n5960), .ZN(U2794) );
  INV_X1 U6998 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6519) );
  AOI21_X1 U6999 ( .B1(n6652), .B2(n6519), .A(n5962), .ZN(n5963) );
  INV_X1 U7000 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6708) );
  INV_X1 U7001 ( .A(n6529), .ZN(n6525) );
  AOI22_X1 U7002 ( .A1(n6529), .A2(n5963), .B1(n6708), .B2(n6525), .ZN(U2795)
         );
  AOI22_X1 U7003 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6089), .B1(n5964), .B2(n6492), .ZN(n5965) );
  OAI21_X1 U7004 ( .B1(n5973), .B2(n6492), .A(n5965), .ZN(n5966) );
  AOI211_X1 U7005 ( .C1(n6091), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n2997), 
        .B(n5966), .ZN(n5969) );
  AOI22_X1 U7006 ( .A1(n6113), .A2(n6032), .B1(n6088), .B2(n5967), .ZN(n5968)
         );
  OAI211_X1 U7007 ( .C1(n5970), .C2(n6101), .A(n5969), .B(n5968), .ZN(U2809)
         );
  AND2_X1 U7008 ( .A1(n6083), .A2(n5971), .ZN(n5981) );
  AOI21_X1 U7009 ( .B1(REIP_REG_16__SCAN_IN), .B2(n5981), .A(
        REIP_REG_17__SCAN_IN), .ZN(n5974) );
  OAI22_X1 U7010 ( .A1(n5974), .A2(n5973), .B1(n5972), .B2(n6073), .ZN(n5975)
         );
  AOI211_X1 U7011 ( .C1(n6089), .C2(EBX_REG_17__SCAN_IN), .A(n2997), .B(n5975), 
        .ZN(n5979) );
  INV_X1 U7012 ( .A(n5976), .ZN(n6116) );
  AOI22_X1 U7013 ( .A1(n6116), .A2(n6032), .B1(n6079), .B2(n5977), .ZN(n5978)
         );
  OAI211_X1 U7014 ( .C1(n6065), .C2(n5980), .A(n5979), .B(n5978), .ZN(U2810)
         );
  INV_X1 U7015 ( .A(n5981), .ZN(n5984) );
  NOR2_X1 U7016 ( .A1(n5982), .A2(n5994), .ZN(n5983) );
  MUX2_X1 U7017 ( .A(n5984), .B(n5983), .S(REIP_REG_16__SCAN_IN), .Z(n5985) );
  OAI21_X1 U7018 ( .B1(n5986), .B2(n6043), .A(n5985), .ZN(n5987) );
  AOI211_X1 U7019 ( .C1(n6091), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n2997), 
        .B(n5987), .ZN(n5990) );
  AOI22_X1 U7020 ( .A1(n6121), .A2(n6032), .B1(n6079), .B2(n5988), .ZN(n5989)
         );
  OAI211_X1 U7021 ( .C1(n6065), .C2(n5991), .A(n5990), .B(n5989), .ZN(U2811)
         );
  AOI22_X1 U7022 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5994), .B1(n5993), .B2(
        n5992), .ZN(n5995) );
  OAI21_X1 U7023 ( .B1(n5996), .B2(n6043), .A(n5995), .ZN(n5997) );
  AOI211_X1 U7024 ( .C1(n6091), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n2997), 
        .B(n5997), .ZN(n6001) );
  AOI22_X1 U7025 ( .A1(n5999), .A2(n6032), .B1(n5998), .B2(n6079), .ZN(n6000)
         );
  OAI211_X1 U7026 ( .C1(n6065), .C2(n6002), .A(n6001), .B(n6000), .ZN(U2813)
         );
  NOR3_X1 U7027 ( .A1(n6090), .A2(REIP_REG_13__SCAN_IN), .A3(n6003), .ZN(n6008) );
  OAI21_X1 U7028 ( .B1(n6004), .B2(n6019), .A(REIP_REG_13__SCAN_IN), .ZN(n6005) );
  OAI211_X1 U7029 ( .C1(n6073), .C2(n6006), .A(n6238), .B(n6005), .ZN(n6007)
         );
  AOI211_X1 U7030 ( .C1(n6089), .C2(EBX_REG_13__SCAN_IN), .A(n6008), .B(n6007), 
        .ZN(n6012) );
  OAI22_X1 U7031 ( .A1(n6128), .A2(n6058), .B1(n6009), .B2(n6101), .ZN(n6010)
         );
  INV_X1 U7032 ( .A(n6010), .ZN(n6011) );
  OAI211_X1 U7033 ( .C1(n6065), .C2(n6013), .A(n6012), .B(n6011), .ZN(U2814)
         );
  NAND2_X1 U7034 ( .A1(n6015), .A2(n6014), .ZN(n6016) );
  AND2_X1 U7035 ( .A1(n3005), .A2(n6016), .ZN(n6102) );
  NOR3_X1 U7036 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6018), .A3(n6017), .ZN(n6022) );
  INV_X1 U7037 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6106) );
  AOI22_X1 U7038 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6091), .B1(
        REIP_REG_11__SCAN_IN), .B2(n6019), .ZN(n6020) );
  OAI211_X1 U7039 ( .C1(n6043), .C2(n6106), .A(n6020), .B(n6238), .ZN(n6021)
         );
  AOI211_X1 U7040 ( .C1(n6102), .C2(n6088), .A(n6022), .B(n6021), .ZN(n6026)
         );
  INV_X1 U7041 ( .A(n6023), .ZN(n6188) );
  OAI22_X1 U7042 ( .A1(n6189), .A2(n6058), .B1(n6101), .B2(n6188), .ZN(n6024)
         );
  INV_X1 U7043 ( .A(n6024), .ZN(n6025) );
  NAND2_X1 U7044 ( .A1(n6026), .A2(n6025), .ZN(U2816) );
  INV_X1 U7045 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6475) );
  INV_X1 U7046 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6473) );
  NOR2_X1 U7047 ( .A1(n6475), .A2(n6473), .ZN(n6027) );
  AOI21_X1 U7048 ( .B1(n6027), .B2(n6048), .A(REIP_REG_8__SCAN_IN), .ZN(n6037)
         );
  OAI22_X1 U7049 ( .A1(n6658), .A2(n6073), .B1(n6065), .B2(n6028), .ZN(n6029)
         );
  AOI211_X1 U7050 ( .C1(n6089), .C2(EBX_REG_8__SCAN_IN), .A(n2997), .B(n6029), 
        .ZN(n6035) );
  INV_X1 U7051 ( .A(n6030), .ZN(n6031) );
  AOI22_X1 U7052 ( .A1(n6033), .A2(n6032), .B1(n6031), .B2(n6079), .ZN(n6034)
         );
  OAI211_X1 U7053 ( .C1(n6037), .C2(n6036), .A(n6035), .B(n6034), .ZN(U2819)
         );
  NAND3_X1 U7054 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6048), .A3(n6475), .ZN(n6046) );
  INV_X1 U7055 ( .A(n6038), .ZN(n6039) );
  NAND2_X1 U7056 ( .A1(n6039), .A2(n6088), .ZN(n6041) );
  AOI21_X1 U7057 ( .B1(n6091), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n2997), 
        .ZN(n6040) );
  OAI211_X1 U7058 ( .C1(n6043), .C2(n6042), .A(n6041), .B(n6040), .ZN(n6044)
         );
  INV_X1 U7059 ( .A(n6044), .ZN(n6045) );
  OAI211_X1 U7060 ( .C1(n6193), .C2(n6058), .A(n6046), .B(n6045), .ZN(n6047)
         );
  INV_X1 U7061 ( .A(n6047), .ZN(n6053) );
  INV_X1 U7062 ( .A(n6048), .ZN(n6049) );
  NOR2_X1 U7063 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6049), .ZN(n6061) );
  OAI21_X1 U7064 ( .B1(n6090), .B2(n6051), .A(n6050), .ZN(n6069) );
  OAI21_X1 U7065 ( .B1(n6061), .B2(n6069), .A(REIP_REG_7__SCAN_IN), .ZN(n6052)
         );
  OAI211_X1 U7066 ( .C1(n6101), .C2(n6197), .A(n6053), .B(n6052), .ZN(U2820)
         );
  NOR2_X1 U7067 ( .A1(n6073), .A2(n6054), .ZN(n6055) );
  AOI211_X1 U7068 ( .C1(n6089), .C2(EBX_REG_6__SCAN_IN), .A(n2997), .B(n6055), 
        .ZN(n6057) );
  NAND2_X1 U7069 ( .A1(n6069), .A2(REIP_REG_6__SCAN_IN), .ZN(n6056) );
  OAI211_X1 U7070 ( .C1(n6059), .C2(n6058), .A(n6057), .B(n6056), .ZN(n6060)
         );
  AOI211_X1 U7071 ( .C1(n6062), .C2(n6088), .A(n6061), .B(n6060), .ZN(n6063)
         );
  OAI21_X1 U7072 ( .B1(n6064), .B2(n6101), .A(n6063), .ZN(U2821) );
  OAI22_X1 U7073 ( .A1(n6209), .A2(n6073), .B1(n6065), .B2(n6256), .ZN(n6066)
         );
  AOI211_X1 U7074 ( .C1(n6089), .C2(EBX_REG_5__SCAN_IN), .A(n2997), .B(n6066), 
        .ZN(n6071) );
  OAI21_X1 U7075 ( .B1(n6090), .B2(n6067), .A(n6471), .ZN(n6068) );
  AOI22_X1 U7076 ( .A1(n6206), .A2(n6098), .B1(n6069), .B2(n6068), .ZN(n6070)
         );
  OAI211_X1 U7077 ( .C1(n6203), .C2(n6101), .A(n6071), .B(n6070), .ZN(U2822)
         );
  AOI22_X1 U7078 ( .A1(EBX_REG_4__SCAN_IN), .A2(n6089), .B1(n6088), .B2(n6266), 
        .ZN(n6087) );
  INV_X1 U7079 ( .A(n6072), .ZN(n6075) );
  INV_X1 U7080 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6074) );
  OAI22_X1 U7081 ( .A1(n6075), .A2(n6095), .B1(n6074), .B2(n6073), .ZN(n6076)
         );
  AOI211_X1 U7082 ( .C1(REIP_REG_4__SCAN_IN), .C2(n6077), .A(n2997), .B(n6076), 
        .ZN(n6086) );
  INV_X1 U7083 ( .A(n6078), .ZN(n6080) );
  AOI22_X1 U7084 ( .A1(n6081), .A2(n6098), .B1(n6080), .B2(n6079), .ZN(n6085)
         );
  INV_X1 U7085 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6469) );
  NAND3_X1 U7086 ( .A1(n6083), .A2(n6469), .A3(n6082), .ZN(n6084) );
  NAND4_X1 U7087 ( .A1(n6087), .A2(n6086), .A3(n6085), .A4(n6084), .ZN(U2823)
         );
  AOI22_X1 U7088 ( .A1(EBX_REG_2__SCAN_IN), .A2(n6089), .B1(n6088), .B2(n6287), 
        .ZN(n6100) );
  OAI21_X1 U7089 ( .B1(n6090), .B2(n6652), .A(n6465), .ZN(n6092) );
  AOI22_X1 U7090 ( .A1(n6093), .A2(n6092), .B1(PHYADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6091), .ZN(n6094) );
  OAI21_X1 U7091 ( .B1(n6096), .B2(n6095), .A(n6094), .ZN(n6097) );
  AOI21_X1 U7092 ( .B1(n6214), .B2(n6098), .A(n6097), .ZN(n6099) );
  OAI211_X1 U7093 ( .C1(n6217), .C2(n6101), .A(n6100), .B(n6099), .ZN(U2825)
         );
  INV_X1 U7094 ( .A(n6102), .ZN(n6227) );
  OAI22_X1 U7095 ( .A1(n6189), .A2(n5466), .B1(n6103), .B2(n6227), .ZN(n6104)
         );
  INV_X1 U7096 ( .A(n6104), .ZN(n6105) );
  OAI21_X1 U7097 ( .B1(n6106), .B2(n6111), .A(n6105), .ZN(U2848) );
  AOI22_X1 U7098 ( .A1(n6109), .A2(n6108), .B1(n6107), .B2(n3008), .ZN(n6110)
         );
  OAI21_X1 U7099 ( .B1(n6112), .B2(n6111), .A(n6110), .ZN(U2856) );
  AOI22_X1 U7100 ( .A1(n6113), .A2(n6120), .B1(n6119), .B2(DATAI_18_), .ZN(
        n6115) );
  AOI22_X1 U7101 ( .A1(n6123), .A2(DATAI_2_), .B1(n6122), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7102 ( .A1(n6115), .A2(n6114), .ZN(U2873) );
  AOI22_X1 U7103 ( .A1(n6116), .A2(n6120), .B1(n6119), .B2(DATAI_17_), .ZN(
        n6118) );
  AOI22_X1 U7104 ( .A1(n6123), .A2(DATAI_1_), .B1(n6122), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U7105 ( .A1(n6118), .A2(n6117), .ZN(U2874) );
  AOI22_X1 U7106 ( .A1(n6121), .A2(n6120), .B1(n6119), .B2(DATAI_16_), .ZN(
        n6125) );
  AOI22_X1 U7107 ( .A1(n6123), .A2(DATAI_0_), .B1(n6122), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U7108 ( .A1(n6125), .A2(n6124), .ZN(U2875) );
  INV_X1 U7109 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6566) );
  INV_X1 U7110 ( .A(DATAI_13_), .ZN(n6127) );
  OAI22_X1 U7111 ( .A1(n6128), .A2(n5863), .B1(n6127), .B2(n6126), .ZN(n6129)
         );
  INV_X1 U7112 ( .A(n6129), .ZN(n6130) );
  OAI21_X1 U7113 ( .B1(n6566), .B2(n6131), .A(n6130), .ZN(U2878) );
  INV_X1 U7114 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n6631) );
  INV_X1 U7115 ( .A(n6745), .ZN(n6132) );
  AOI22_X1 U7116 ( .A1(n6132), .A2(EAX_REG_26__SCAN_IN), .B1(n6746), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6133) );
  OAI21_X1 U7117 ( .B1(n6631), .B2(n6750), .A(n6133), .ZN(U2897) );
  INV_X1 U7118 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6181) );
  INV_X1 U7119 ( .A(n6145), .ZN(n6158) );
  AOI22_X1 U7120 ( .A1(n6746), .A2(LWORD_REG_15__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6134) );
  OAI21_X1 U7121 ( .B1(n6181), .B2(n6158), .A(n6134), .ZN(U2908) );
  INV_X1 U7122 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n6712) );
  AOI22_X1 U7123 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6145), .B1(n6746), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n6135) );
  OAI21_X1 U7124 ( .B1(n6712), .B2(n6750), .A(n6135), .ZN(U2909) );
  AOI22_X1 U7125 ( .A1(n6746), .A2(LWORD_REG_13__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6136) );
  OAI21_X1 U7126 ( .B1(n6566), .B2(n6158), .A(n6136), .ZN(U2910) );
  INV_X1 U7127 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6629) );
  AOI22_X1 U7128 ( .A1(n6746), .A2(LWORD_REG_12__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6137) );
  OAI21_X1 U7129 ( .B1(n6629), .B2(n6158), .A(n6137), .ZN(U2911) );
  INV_X1 U7130 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6139) );
  AOI22_X1 U7131 ( .A1(n6746), .A2(LWORD_REG_11__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6138) );
  OAI21_X1 U7132 ( .B1(n6139), .B2(n6158), .A(n6138), .ZN(U2912) );
  INV_X1 U7133 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n6725) );
  AOI22_X1 U7134 ( .A1(EAX_REG_10__SCAN_IN), .A2(n6145), .B1(n6746), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n6140) );
  OAI21_X1 U7135 ( .B1(n6725), .B2(n6750), .A(n6140), .ZN(U2913) );
  INV_X1 U7136 ( .A(LWORD_REG_9__SCAN_IN), .ZN(n6602) );
  AOI22_X1 U7137 ( .A1(EAX_REG_9__SCAN_IN), .A2(n6145), .B1(
        DATAO_REG_9__SCAN_IN), .B2(n6156), .ZN(n6141) );
  OAI21_X1 U7138 ( .B1(n6142), .B2(n6602), .A(n6141), .ZN(U2914) );
  AOI22_X1 U7139 ( .A1(n6746), .A2(LWORD_REG_8__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6143) );
  OAI21_X1 U7140 ( .B1(n4385), .B2(n6158), .A(n6143), .ZN(U2915) );
  AOI22_X1 U7141 ( .A1(n6746), .A2(LWORD_REG_7__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6144) );
  OAI21_X1 U7142 ( .B1(n4255), .B2(n6158), .A(n6144), .ZN(U2916) );
  AOI222_X1 U7143 ( .A1(n6156), .A2(DATAO_REG_6__SCAN_IN), .B1(n6145), .B2(
        EAX_REG_6__SCAN_IN), .C1(n6746), .C2(LWORD_REG_6__SCAN_IN), .ZN(n6146)
         );
  INV_X1 U7144 ( .A(n6146), .ZN(U2917) );
  AOI22_X1 U7145 ( .A1(n6746), .A2(LWORD_REG_5__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6147) );
  OAI21_X1 U7146 ( .B1(n4062), .B2(n6158), .A(n6147), .ZN(U2918) );
  AOI22_X1 U7147 ( .A1(n6746), .A2(LWORD_REG_4__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6148) );
  OAI21_X1 U7148 ( .B1(n6149), .B2(n6158), .A(n6148), .ZN(U2919) );
  INV_X1 U7149 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6151) );
  AOI22_X1 U7150 ( .A1(n6746), .A2(LWORD_REG_3__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6150) );
  OAI21_X1 U7151 ( .B1(n6151), .B2(n6158), .A(n6150), .ZN(U2920) );
  AOI22_X1 U7152 ( .A1(n6746), .A2(LWORD_REG_2__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6152) );
  OAI21_X1 U7153 ( .B1(n6153), .B2(n6158), .A(n6152), .ZN(U2921) );
  INV_X1 U7154 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6155) );
  AOI22_X1 U7155 ( .A1(n6746), .A2(LWORD_REG_1__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6154) );
  OAI21_X1 U7156 ( .B1(n6155), .B2(n6158), .A(n6154), .ZN(U2922) );
  AOI22_X1 U7157 ( .A1(n6746), .A2(LWORD_REG_0__SCAN_IN), .B1(n6156), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6157) );
  OAI21_X1 U7158 ( .B1(n6159), .B2(n6158), .A(n6157), .ZN(U2923) );
  AOI22_X1 U7159 ( .A1(EAX_REG_25__SCAN_IN), .A2(n6174), .B1(n6164), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U7160 ( .A1(n6177), .A2(DATAI_9_), .ZN(n6166) );
  NAND2_X1 U7161 ( .A1(n6160), .A2(n6166), .ZN(U2933) );
  AOI22_X1 U7162 ( .A1(EAX_REG_26__SCAN_IN), .A2(n6174), .B1(n6164), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7163 ( .A1(n6177), .A2(DATAI_10_), .ZN(n6168) );
  NAND2_X1 U7164 ( .A1(n6161), .A2(n6168), .ZN(U2934) );
  AOI22_X1 U7165 ( .A1(EAX_REG_27__SCAN_IN), .A2(n6174), .B1(n6164), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U7166 ( .A1(n6177), .A2(DATAI_11_), .ZN(n6170) );
  NAND2_X1 U7167 ( .A1(n6162), .A2(n6170), .ZN(U2935) );
  AOI22_X1 U7168 ( .A1(EAX_REG_28__SCAN_IN), .A2(n6174), .B1(n6164), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7169 ( .A1(n6177), .A2(DATAI_12_), .ZN(n6172) );
  NAND2_X1 U7170 ( .A1(n6163), .A2(n6172), .ZN(U2936) );
  AOI22_X1 U7171 ( .A1(EAX_REG_30__SCAN_IN), .A2(n6174), .B1(n6164), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7172 ( .A1(n6177), .A2(DATAI_14_), .ZN(n6175) );
  NAND2_X1 U7173 ( .A1(n6165), .A2(n6175), .ZN(U2938) );
  AOI22_X1 U7174 ( .A1(EAX_REG_9__SCAN_IN), .A2(n6174), .B1(
        LWORD_REG_9__SCAN_IN), .B2(n6178), .ZN(n6167) );
  NAND2_X1 U7175 ( .A1(n6167), .A2(n6166), .ZN(U2948) );
  AOI22_X1 U7176 ( .A1(EAX_REG_10__SCAN_IN), .A2(n6174), .B1(n6178), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U7177 ( .A1(n6169), .A2(n6168), .ZN(U2949) );
  AOI22_X1 U7178 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6174), .B1(n6178), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7179 ( .A1(n6171), .A2(n6170), .ZN(U2950) );
  AOI22_X1 U7180 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6174), .B1(n6178), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7181 ( .A1(n6173), .A2(n6172), .ZN(U2951) );
  AOI22_X1 U7182 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6174), .B1(n6178), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7183 ( .A1(n6176), .A2(n6175), .ZN(U2953) );
  AOI22_X1 U7184 ( .A1(n6178), .A2(LWORD_REG_15__SCAN_IN), .B1(n6177), .B2(
        DATAI_15_), .ZN(n6179) );
  OAI21_X1 U7185 ( .B1(n6181), .B2(n6180), .A(n6179), .ZN(U2954) );
  AND2_X1 U7186 ( .A1(n6183), .A2(n6182), .ZN(n6187) );
  AND2_X1 U7187 ( .A1(n6185), .A2(n6184), .ZN(n6186) );
  XNOR2_X1 U7188 ( .A(n6187), .B(n6186), .ZN(n6228) );
  AOI22_X1 U7189 ( .A1(n2997), .A2(REIP_REG_11__SCAN_IN), .B1(n6218), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6192) );
  OAI22_X1 U7190 ( .A1(n6189), .A2(n6194), .B1(n6225), .B2(n6188), .ZN(n6190)
         );
  INV_X1 U7191 ( .A(n6190), .ZN(n6191) );
  OAI211_X1 U7192 ( .C1(n6228), .C2(n6195), .A(n6192), .B(n6191), .ZN(U2975)
         );
  INV_X1 U7193 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6728) );
  OAI222_X1 U7194 ( .A1(n6225), .A2(n6197), .B1(n6196), .B2(n6195), .C1(n6194), 
        .C2(n6193), .ZN(n6198) );
  INV_X1 U7195 ( .A(n6198), .ZN(n6200) );
  OAI211_X1 U7196 ( .C1(n6728), .C2(n6208), .A(n6200), .B(n6199), .ZN(U2979)
         );
  XOR2_X1 U7197 ( .A(n6202), .B(n6201), .Z(n6258) );
  INV_X1 U7198 ( .A(n6203), .ZN(n6205) );
  AOI222_X1 U7199 ( .A1(n6258), .A2(n6221), .B1(n6219), .B2(n6206), .C1(n6205), 
        .C2(n6204), .ZN(n6207) );
  NAND2_X1 U7200 ( .A1(n2997), .A2(REIP_REG_5__SCAN_IN), .ZN(n6259) );
  OAI211_X1 U7201 ( .C1(n6209), .C2(n6208), .A(n6207), .B(n6259), .ZN(U2981)
         );
  AOI22_X1 U7202 ( .A1(n2997), .A2(REIP_REG_2__SCAN_IN), .B1(n6218), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U7203 ( .A1(n6211), .A2(n6210), .ZN(n6212) );
  XOR2_X1 U7204 ( .A(n6213), .B(n6212), .Z(n6290) );
  AOI22_X1 U7205 ( .A1(n6290), .A2(n6221), .B1(n6219), .B2(n6214), .ZN(n6215)
         );
  OAI211_X1 U7206 ( .C1(n6225), .C2(n6217), .A(n6216), .B(n6215), .ZN(U2984)
         );
  AOI22_X1 U7207 ( .A1(n2997), .A2(REIP_REG_1__SCAN_IN), .B1(n6218), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6224) );
  AOI22_X1 U7208 ( .A1(n6222), .A2(n6221), .B1(n6220), .B2(n6219), .ZN(n6223)
         );
  OAI211_X1 U7209 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6225), .A(n6224), 
        .B(n6223), .ZN(U2985) );
  INV_X1 U7210 ( .A(n6226), .ZN(n6231) );
  INV_X1 U7211 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6482) );
  OAI22_X1 U7212 ( .A1(n6227), .A2(n6303), .B1(n6482), .B2(n6238), .ZN(n6230)
         );
  NOR2_X1 U7213 ( .A1(n6228), .A2(n6269), .ZN(n6229) );
  AOI211_X1 U7214 ( .C1(n6234), .C2(n6231), .A(n6230), .B(n6229), .ZN(n6232)
         );
  OAI21_X1 U7215 ( .B1(n6234), .B2(n6233), .A(n6232), .ZN(U3007) );
  AOI21_X1 U7216 ( .B1(n6242), .B2(n6236), .A(n6235), .ZN(n6255) );
  OAI222_X1 U7217 ( .A1(n6239), .A2(n6303), .B1(n6238), .B2(n6479), .C1(n6269), 
        .C2(n6237), .ZN(n6240) );
  INV_X1 U7218 ( .A(n6240), .ZN(n6245) );
  NOR2_X1 U7219 ( .A1(n6242), .A2(n6241), .ZN(n6251) );
  OAI211_X1 U7220 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6251), .B(n6243), .ZN(n6244) );
  OAI211_X1 U7221 ( .C1(n6255), .C2(n6246), .A(n6245), .B(n6244), .ZN(U3008)
         );
  INV_X1 U7222 ( .A(n6247), .ZN(n6248) );
  AOI21_X1 U7223 ( .B1(n6249), .B2(n6288), .A(n6248), .ZN(n6253) );
  AOI22_X1 U7224 ( .A1(n6251), .A2(n6254), .B1(n6298), .B2(n6250), .ZN(n6252)
         );
  OAI211_X1 U7225 ( .C1(n6255), .C2(n6254), .A(n6253), .B(n6252), .ZN(U3009)
         );
  NOR2_X1 U7226 ( .A1(n6653), .A2(n3333), .ZN(n6274) );
  AOI21_X1 U7227 ( .B1(n6274), .B2(n6275), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6261) );
  INV_X1 U7228 ( .A(n6256), .ZN(n6257) );
  AOI22_X1 U7229 ( .A1(n6258), .A2(n6298), .B1(n6288), .B2(n6257), .ZN(n6260)
         );
  OAI211_X1 U7230 ( .C1(n6262), .C2(n6261), .A(n6260), .B(n6259), .ZN(U3013)
         );
  OAI21_X1 U7231 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6275), .ZN(n6273) );
  AOI21_X1 U7232 ( .B1(n6264), .B2(n6263), .A(n6289), .ZN(n6282) );
  OR2_X1 U7233 ( .A1(n6282), .A2(n3333), .ZN(n6268) );
  AOI21_X1 U7234 ( .B1(n6266), .B2(n6288), .A(n6265), .ZN(n6267) );
  OAI211_X1 U7235 ( .C1(n6270), .C2(n6269), .A(n6268), .B(n6267), .ZN(n6271)
         );
  INV_X1 U7236 ( .A(n6271), .ZN(n6272) );
  OAI21_X1 U7237 ( .B1(n6274), .B2(n6273), .A(n6272), .ZN(U3014) );
  INV_X1 U7238 ( .A(n6275), .ZN(n6279) );
  AOI22_X1 U7239 ( .A1(n3008), .A2(n6288), .B1(n2997), .B2(REIP_REG_3__SCAN_IN), .ZN(n6278) );
  OR2_X1 U7240 ( .A1(n6276), .A2(n6269), .ZN(n6277) );
  OAI211_X1 U7241 ( .C1(n6279), .C2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6278), 
        .B(n6277), .ZN(n6280) );
  INV_X1 U7242 ( .A(n6280), .ZN(n6281) );
  OAI21_X1 U7243 ( .B1(n6282), .B2(n6653), .A(n6281), .ZN(U3015) );
  NAND3_X1 U7244 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A3(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6284) );
  AOI21_X1 U7245 ( .B1(n6285), .B2(n6284), .A(n6283), .ZN(n6286) );
  AOI21_X1 U7246 ( .B1(n6288), .B2(n6287), .A(n6286), .ZN(n6296) );
  AOI22_X1 U7247 ( .A1(n6290), .A2(n6298), .B1(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6289), .ZN(n6295) );
  NAND2_X1 U7248 ( .A1(n2997), .A2(REIP_REG_2__SCAN_IN), .ZN(n6294) );
  NAND3_X1 U7249 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6292), .A3(n6291), 
        .ZN(n6293) );
  NAND4_X1 U7250 ( .A1(n6296), .A2(n6295), .A3(n6294), .A4(n6293), .ZN(U3016)
         );
  AND3_X1 U7251 ( .A1(n6299), .A2(n6298), .A3(n6297), .ZN(n6305) );
  OAI211_X1 U7252 ( .C1(n6303), .C2(n6302), .A(n6301), .B(n6300), .ZN(n6304)
         );
  NOR2_X1 U7253 ( .A1(n6305), .A2(n6304), .ZN(n6306) );
  OAI221_X1 U7254 ( .B1(n6309), .B2(n6308), .C1(n6309), .C2(n6307), .A(n6306), 
        .ZN(U3018) );
  NOR2_X1 U7255 ( .A1(n6405), .A2(n6310), .ZN(U3019) );
  AOI22_X1 U7256 ( .A1(n6312), .A2(n6326), .B1(n6311), .B2(n6325), .ZN(n6315)
         );
  AOI22_X1 U7257 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6328), .B1(n6313), 
        .B2(n6327), .ZN(n6314) );
  OAI211_X1 U7258 ( .C1(n6331), .C2(n6316), .A(n6315), .B(n6314), .ZN(U3045)
         );
  AOI22_X1 U7259 ( .A1(n6335), .A2(n6326), .B1(n6334), .B2(n6325), .ZN(n6318)
         );
  AOI22_X1 U7260 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6328), .B1(n6336), 
        .B2(n6327), .ZN(n6317) );
  OAI211_X1 U7261 ( .C1(n6331), .C2(n6339), .A(n6318), .B(n6317), .ZN(U3046)
         );
  AOI22_X1 U7262 ( .A1(n6360), .A2(n6326), .B1(n6359), .B2(n6325), .ZN(n6320)
         );
  AOI22_X1 U7263 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6328), .B1(n6361), 
        .B2(n6327), .ZN(n6319) );
  OAI211_X1 U7264 ( .C1(n6331), .C2(n6364), .A(n6320), .B(n6319), .ZN(U3048)
         );
  AOI22_X1 U7265 ( .A1(n6366), .A2(n6326), .B1(n6365), .B2(n6325), .ZN(n6322)
         );
  AOI22_X1 U7266 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6328), .B1(n6367), 
        .B2(n6327), .ZN(n6321) );
  OAI211_X1 U7267 ( .C1(n6331), .C2(n6370), .A(n6322), .B(n6321), .ZN(U3049)
         );
  AOI22_X1 U7268 ( .A1(n6372), .A2(n6326), .B1(n6371), .B2(n6325), .ZN(n6324)
         );
  AOI22_X1 U7269 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6328), .B1(n6373), 
        .B2(n6327), .ZN(n6323) );
  OAI211_X1 U7270 ( .C1(n6331), .C2(n6376), .A(n6324), .B(n6323), .ZN(U3050)
         );
  AOI22_X1 U7271 ( .A1(n6380), .A2(n6326), .B1(n6378), .B2(n6325), .ZN(n6330)
         );
  AOI22_X1 U7272 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6328), .B1(n6382), 
        .B2(n6327), .ZN(n6329) );
  OAI211_X1 U7273 ( .C1(n6331), .C2(n6387), .A(n6330), .B(n6329), .ZN(U3051)
         );
  INV_X1 U7274 ( .A(n6332), .ZN(n6345) );
  INV_X1 U7275 ( .A(n6333), .ZN(n6344) );
  AOI22_X1 U7276 ( .A1(n6335), .A2(n6345), .B1(n6334), .B2(n6344), .ZN(n6338)
         );
  AOI22_X1 U7277 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6347), .B1(n6336), 
        .B2(n6346), .ZN(n6337) );
  OAI211_X1 U7278 ( .C1(n6339), .C2(n6350), .A(n6338), .B(n6337), .ZN(U3078)
         );
  AOI22_X1 U7279 ( .A1(n6360), .A2(n6345), .B1(n6359), .B2(n6344), .ZN(n6341)
         );
  AOI22_X1 U7280 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6347), .B1(n6361), 
        .B2(n6346), .ZN(n6340) );
  OAI211_X1 U7281 ( .C1(n6364), .C2(n6350), .A(n6341), .B(n6340), .ZN(U3080)
         );
  AOI22_X1 U7282 ( .A1(n6366), .A2(n6345), .B1(n6365), .B2(n6344), .ZN(n6343)
         );
  AOI22_X1 U7283 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6347), .B1(n6367), 
        .B2(n6346), .ZN(n6342) );
  OAI211_X1 U7284 ( .C1(n6370), .C2(n6350), .A(n6343), .B(n6342), .ZN(U3081)
         );
  AOI22_X1 U7285 ( .A1(n6380), .A2(n6345), .B1(n6378), .B2(n6344), .ZN(n6349)
         );
  AOI22_X1 U7286 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6347), .B1(n6382), 
        .B2(n6346), .ZN(n6348) );
  OAI211_X1 U7287 ( .C1(n6387), .C2(n6350), .A(n6349), .B(n6348), .ZN(U3083)
         );
  INV_X1 U7288 ( .A(n6351), .ZN(n6379) );
  INV_X1 U7289 ( .A(n6352), .ZN(n6377) );
  AOI22_X1 U7290 ( .A1(n6354), .A2(n6379), .B1(n6353), .B2(n6377), .ZN(n6357)
         );
  AOI22_X1 U7291 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6383), .B1(n6355), 
        .B2(n6381), .ZN(n6356) );
  OAI211_X1 U7292 ( .C1(n6358), .C2(n6386), .A(n6357), .B(n6356), .ZN(U3108)
         );
  AOI22_X1 U7293 ( .A1(n6360), .A2(n6379), .B1(n6359), .B2(n6377), .ZN(n6363)
         );
  AOI22_X1 U7294 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6383), .B1(n6361), 
        .B2(n6381), .ZN(n6362) );
  OAI211_X1 U7295 ( .C1(n6364), .C2(n6386), .A(n6363), .B(n6362), .ZN(U3112)
         );
  AOI22_X1 U7296 ( .A1(n6366), .A2(n6379), .B1(n6365), .B2(n6377), .ZN(n6369)
         );
  AOI22_X1 U7297 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6383), .B1(n6367), 
        .B2(n6381), .ZN(n6368) );
  OAI211_X1 U7298 ( .C1(n6370), .C2(n6386), .A(n6369), .B(n6368), .ZN(U3113)
         );
  AOI22_X1 U7299 ( .A1(n6372), .A2(n6379), .B1(n6371), .B2(n6377), .ZN(n6375)
         );
  AOI22_X1 U7300 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6383), .B1(n6373), 
        .B2(n6381), .ZN(n6374) );
  OAI211_X1 U7301 ( .C1(n6376), .C2(n6386), .A(n6375), .B(n6374), .ZN(U3114)
         );
  AOI22_X1 U7302 ( .A1(n6380), .A2(n6379), .B1(n6378), .B2(n6377), .ZN(n6385)
         );
  AOI22_X1 U7303 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6383), .B1(n6382), 
        .B2(n6381), .ZN(n6384) );
  OAI211_X1 U7304 ( .C1(n6387), .C2(n6386), .A(n6385), .B(n6384), .ZN(U3115)
         );
  NOR3_X1 U7305 ( .A1(n6390), .A2(n6389), .A3(n6388), .ZN(n6397) );
  INV_X1 U7306 ( .A(n6397), .ZN(n6395) );
  INV_X1 U7307 ( .A(n6391), .ZN(n6392) );
  OAI211_X1 U7308 ( .C1(n6395), .C2(n6394), .A(n6393), .B(n6392), .ZN(n6396)
         );
  OAI21_X1 U7309 ( .B1(n6397), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6396), 
        .ZN(n6398) );
  AOI222_X1 U7310 ( .A1(n6400), .A2(n6399), .B1(n6400), .B2(n6398), .C1(n6399), 
        .C2(n6398), .ZN(n6404) );
  OR2_X1 U7311 ( .A1(n6404), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6403)
         );
  INV_X1 U7312 ( .A(n6401), .ZN(n6402) );
  NAND2_X1 U7313 ( .A1(n6403), .A2(n6402), .ZN(n6407) );
  NAND2_X1 U7314 ( .A1(n6404), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6406) );
  NAND3_X1 U7315 ( .A1(n6407), .A2(n6406), .A3(n6405), .ZN(n6416) );
  OAI21_X1 U7316 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6408), 
        .ZN(n6409) );
  NAND4_X1 U7317 ( .A1(n6412), .A2(n6411), .A3(n6410), .A4(n6409), .ZN(n6413)
         );
  NOR2_X1 U7318 ( .A1(n6414), .A2(n6413), .ZN(n6415) );
  AND2_X1 U7319 ( .A1(n6416), .A2(n6415), .ZN(n6433) );
  NOR2_X1 U7320 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6455), .ZN(n6445) );
  NAND2_X1 U7321 ( .A1(n6433), .A2(n6435), .ZN(n6418) );
  NAND2_X1 U7322 ( .A1(READY_N), .A2(n6746), .ZN(n6417) );
  NAND2_X1 U7323 ( .A1(n6418), .A2(n6417), .ZN(n6422) );
  OR2_X1 U7324 ( .A1(n6420), .A2(n6419), .ZN(n6421) );
  NOR2_X1 U7325 ( .A1(n6445), .A2(n6522), .ZN(n6429) );
  OAI21_X1 U7326 ( .B1(n6441), .B2(n6423), .A(n6540), .ZN(n6424) );
  OR2_X1 U7327 ( .A1(n6522), .A2(n6424), .ZN(n6428) );
  AOI21_X1 U7328 ( .B1(n6426), .B2(n6521), .A(n6425), .ZN(n6427) );
  OAI211_X1 U7329 ( .C1(n6429), .C2(n6540), .A(n6428), .B(n6427), .ZN(n6430)
         );
  INV_X1 U7330 ( .A(n6430), .ZN(n6431) );
  OAI21_X1 U7331 ( .B1(n6433), .B2(n6432), .A(n6431), .ZN(U3148) );
  NOR2_X1 U7332 ( .A1(n6540), .A2(n6434), .ZN(n6436) );
  AOI21_X1 U7333 ( .B1(n6436), .B2(n6455), .A(n6435), .ZN(n6439) );
  NAND2_X1 U7334 ( .A1(n6540), .A2(n6532), .ZN(n6442) );
  OAI211_X1 U7335 ( .C1(n6522), .C2(n6445), .A(STATE2_REG_1__SCAN_IN), .B(
        n6442), .ZN(n6437) );
  OAI211_X1 U7336 ( .C1(n6522), .C2(n6439), .A(n6438), .B(n6437), .ZN(U3149)
         );
  NAND3_X1 U7337 ( .A1(n6442), .A2(n6441), .A3(n6440), .ZN(n6444) );
  OAI21_X1 U7338 ( .B1(n6445), .B2(n6444), .A(n6443), .ZN(U3150) );
  INV_X1 U7339 ( .A(DATAWIDTH_REG_31__SCAN_IN), .ZN(n6614) );
  NOR2_X1 U7340 ( .A1(n6520), .A2(n6614), .ZN(U3151) );
  INV_X1 U7341 ( .A(n6520), .ZN(n6446) );
  AND2_X1 U7342 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6446), .ZN(U3152) );
  AND2_X1 U7343 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6446), .ZN(U3153) );
  AND2_X1 U7344 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6446), .ZN(U3154) );
  AND2_X1 U7345 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6446), .ZN(U3155) );
  AND2_X1 U7346 ( .A1(n6446), .A2(DATAWIDTH_REG_26__SCAN_IN), .ZN(U3156) );
  AND2_X1 U7347 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6446), .ZN(U3157) );
  AND2_X1 U7348 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6446), .ZN(U3158) );
  INV_X1 U7349 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6628) );
  NOR2_X1 U7350 ( .A1(n6520), .A2(n6628), .ZN(U3159) );
  AND2_X1 U7351 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6446), .ZN(U3160) );
  AND2_X1 U7352 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6446), .ZN(U3161) );
  AND2_X1 U7353 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6446), .ZN(U3162) );
  AND2_X1 U7354 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6446), .ZN(U3163) );
  AND2_X1 U7355 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6446), .ZN(U3164) );
  AND2_X1 U7356 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6446), .ZN(U3165) );
  AND2_X1 U7357 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6446), .ZN(U3166) );
  AND2_X1 U7358 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6446), .ZN(U3167) );
  AND2_X1 U7359 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6446), .ZN(U3168) );
  AND2_X1 U7360 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6446), .ZN(U3169) );
  AND2_X1 U7361 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6446), .ZN(U3170) );
  AND2_X1 U7362 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6446), .ZN(U3171) );
  AND2_X1 U7363 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6446), .ZN(U3172) );
  AND2_X1 U7364 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6446), .ZN(U3173) );
  AND2_X1 U7365 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6446), .ZN(U3174) );
  AND2_X1 U7366 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6446), .ZN(U3175) );
  AND2_X1 U7367 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6446), .ZN(U3176) );
  AND2_X1 U7368 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6446), .ZN(U3177) );
  AND2_X1 U7369 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6446), .ZN(U3178) );
  AND2_X1 U7370 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6446), .ZN(U3179) );
  AND2_X1 U7371 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6446), .ZN(U3180) );
  NAND2_X1 U7372 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6451) );
  NAND2_X1 U7373 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6456) );
  NAND2_X1 U7374 ( .A1(STATE_REG_1__SCAN_IN), .A2(READY_N), .ZN(n6457) );
  NAND2_X1 U7375 ( .A1(n6456), .A2(n6457), .ZN(n6448) );
  INV_X1 U7376 ( .A(NA_N), .ZN(n6447) );
  AOI221_X1 U7377 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6447), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6462) );
  AOI21_X1 U7378 ( .B1(n6458), .B2(n6448), .A(n6462), .ZN(n6449) );
  OAI221_X1 U7379 ( .B1(n6504), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n6504), 
        .C2(n6451), .A(n6449), .ZN(U3181) );
  INV_X1 U7380 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6650) );
  NOR2_X1 U7381 ( .A1(n6450), .A2(n6650), .ZN(n6453) );
  INV_X1 U7382 ( .A(n6451), .ZN(n6452) );
  OAI21_X1 U7383 ( .B1(n6453), .B2(n6452), .A(n6456), .ZN(n6454) );
  NAND3_X1 U7384 ( .A1(n6539), .A2(n6457), .A3(n6454), .ZN(U3182) );
  AOI221_X1 U7385 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6455), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6460) );
  OAI211_X1 U7386 ( .C1(n6458), .C2(n6457), .A(STATE_REG_0__SCAN_IN), .B(n6456), .ZN(n6459) );
  AOI21_X1 U7387 ( .B1(HOLD), .B2(n6460), .A(n6459), .ZN(n6463) );
  NAND4_X1 U7388 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .A3(
        READY_N), .A4(REQUESTPENDING_REG_SCAN_IN), .ZN(n6461) );
  OAI22_X1 U7389 ( .A1(n6463), .A2(n6462), .B1(NA_N), .B2(n6461), .ZN(U3183)
         );
  NOR2_X2 U7390 ( .A1(n6550), .A2(STATE_REG_2__SCAN_IN), .ZN(n6513) );
  INV_X1 U7391 ( .A(n6513), .ZN(n6508) );
  INV_X1 U7392 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6640) );
  NOR2_X1 U7393 ( .A1(n6464), .A2(n6550), .ZN(n6506) );
  INV_X1 U7394 ( .A(n6506), .ZN(n6515) );
  OAI222_X1 U7395 ( .A1(n6508), .A2(n6465), .B1(n6640), .B2(n6504), .C1(n6652), 
        .C2(n6515), .ZN(U3184) );
  INV_X1 U7396 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n6626) );
  OAI222_X1 U7397 ( .A1(n6515), .A2(n6465), .B1(n6626), .B2(n6504), .C1(n6467), 
        .C2(n6508), .ZN(U3185) );
  AOI22_X1 U7398 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6513), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6550), .ZN(n6466) );
  OAI21_X1 U7399 ( .B1(n6467), .B2(n6515), .A(n6466), .ZN(U3186) );
  AOI22_X1 U7400 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6513), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6550), .ZN(n6468) );
  OAI21_X1 U7401 ( .B1(n6469), .B2(n6515), .A(n6468), .ZN(U3187) );
  AOI22_X1 U7402 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6513), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6531), .ZN(n6470) );
  OAI21_X1 U7403 ( .B1(n6471), .B2(n6515), .A(n6470), .ZN(U3188) );
  AOI22_X1 U7404 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6513), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6531), .ZN(n6472) );
  OAI21_X1 U7405 ( .B1(n6473), .B2(n6515), .A(n6472), .ZN(U3189) );
  AOI22_X1 U7406 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6513), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6531), .ZN(n6474) );
  OAI21_X1 U7407 ( .B1(n6475), .B2(n6515), .A(n6474), .ZN(U3190) );
  AOI22_X1 U7408 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6531), .ZN(n6476) );
  OAI21_X1 U7409 ( .B1(n6477), .B2(n6508), .A(n6476), .ZN(U3191) );
  AOI22_X1 U7410 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6531), .ZN(n6478) );
  OAI21_X1 U7411 ( .B1(n6479), .B2(n6508), .A(n6478), .ZN(U3192) );
  AOI22_X1 U7412 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6531), .ZN(n6480) );
  OAI21_X1 U7413 ( .B1(n6482), .B2(n6508), .A(n6480), .ZN(U3193) );
  AOI22_X1 U7414 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6513), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6531), .ZN(n6481) );
  OAI21_X1 U7415 ( .B1(n6482), .B2(n6515), .A(n6481), .ZN(U3194) );
  AOI22_X1 U7416 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6531), .ZN(n6483) );
  OAI21_X1 U7417 ( .B1(n6485), .B2(n6508), .A(n6483), .ZN(U3195) );
  AOI22_X1 U7418 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6513), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6531), .ZN(n6484) );
  OAI21_X1 U7419 ( .B1(n6485), .B2(n6515), .A(n6484), .ZN(U3196) );
  AOI22_X1 U7420 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6531), .ZN(n6486) );
  OAI21_X1 U7421 ( .B1(n6487), .B2(n6508), .A(n6486), .ZN(U3197) );
  AOI22_X1 U7422 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6531), .ZN(n6488) );
  OAI21_X1 U7423 ( .B1(n6490), .B2(n6508), .A(n6488), .ZN(U3198) );
  AOI22_X1 U7424 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6513), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6531), .ZN(n6489) );
  OAI21_X1 U7425 ( .B1(n6490), .B2(n6515), .A(n6489), .ZN(U3199) );
  AOI22_X1 U7426 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6531), .ZN(n6491) );
  OAI21_X1 U7427 ( .B1(n6492), .B2(n6508), .A(n6491), .ZN(U3200) );
  AOI22_X1 U7428 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6531), .ZN(n6493) );
  OAI21_X1 U7429 ( .B1(n6495), .B2(n6508), .A(n6493), .ZN(U3201) );
  AOI22_X1 U7430 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6513), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6531), .ZN(n6494) );
  OAI21_X1 U7431 ( .B1(n6495), .B2(n6515), .A(n6494), .ZN(U3202) );
  AOI22_X1 U7432 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6513), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6531), .ZN(n6496) );
  OAI21_X1 U7433 ( .B1(n6497), .B2(n6515), .A(n6496), .ZN(U3203) );
  AOI22_X1 U7434 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6531), .ZN(n6498) );
  OAI21_X1 U7435 ( .B1(n6499), .B2(n6508), .A(n6498), .ZN(U3204) );
  INV_X1 U7436 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6624) );
  OAI222_X1 U7437 ( .A1(n6515), .A2(n6499), .B1(n6624), .B2(n6504), .C1(n6655), 
        .C2(n6508), .ZN(U3205) );
  AOI22_X1 U7438 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6531), .ZN(n6500) );
  OAI21_X1 U7439 ( .B1(n6501), .B2(n6508), .A(n6500), .ZN(U3206) );
  INV_X1 U7440 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6711) );
  OAI222_X1 U7441 ( .A1(n6508), .A2(n6503), .B1(n6711), .B2(n6504), .C1(n6501), 
        .C2(n6515), .ZN(U3207) );
  AOI22_X1 U7442 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6513), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6550), .ZN(n6502) );
  OAI21_X1 U7443 ( .B1(n6503), .B2(n6515), .A(n6502), .ZN(U3208) );
  INV_X1 U7444 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6721) );
  OAI222_X1 U7445 ( .A1(n6515), .A2(n6505), .B1(n6721), .B2(n6504), .C1(n6556), 
        .C2(n6508), .ZN(U3209) );
  AOI22_X1 U7446 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6506), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6550), .ZN(n6507) );
  OAI21_X1 U7447 ( .B1(n6510), .B2(n6508), .A(n6507), .ZN(U3210) );
  AOI22_X1 U7448 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6513), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6550), .ZN(n6509) );
  OAI21_X1 U7449 ( .B1(n6510), .B2(n6515), .A(n6509), .ZN(U3211) );
  AOI22_X1 U7450 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6513), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6550), .ZN(n6511) );
  OAI21_X1 U7451 ( .B1(n6512), .B2(n6515), .A(n6511), .ZN(U3212) );
  AOI22_X1 U7452 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6513), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6550), .ZN(n6514) );
  OAI21_X1 U7453 ( .B1(n6516), .B2(n6515), .A(n6514), .ZN(U3213) );
  MUX2_X1 U7454 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6550), .Z(U3445) );
  MUX2_X1 U7455 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6550), .Z(U3446) );
  MUX2_X1 U7456 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6550), .Z(U3447) );
  MUX2_X1 U7457 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6550), .Z(U3448) );
  OAI21_X1 U7458 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6520), .A(n6518), .ZN(
        n6517) );
  INV_X1 U7459 ( .A(n6517), .ZN(U3451) );
  OAI21_X1 U7460 ( .B1(n6520), .B2(n6519), .A(n6518), .ZN(U3452) );
  AOI221_X1 U7461 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6540), .C1(
        STATE2_REG_3__SCAN_IN), .C2(n6522), .A(n6521), .ZN(n6523) );
  INV_X1 U7462 ( .A(n6523), .ZN(U3453) );
  AOI21_X1 U7463 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6524) );
  AOI22_X1 U7464 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6524), .B2(n6652), .ZN(n6527) );
  INV_X1 U7465 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6526) );
  AOI22_X1 U7466 ( .A1(n6529), .A2(n6527), .B1(n6526), .B2(n6525), .ZN(U3468)
         );
  INV_X1 U7467 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6730) );
  OAI21_X1 U7468 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6529), .ZN(n6528) );
  OAI21_X1 U7469 ( .B1(n6529), .B2(n6730), .A(n6528), .ZN(U3469) );
  NAND2_X1 U7470 ( .A1(n6531), .A2(W_R_N_REG_SCAN_IN), .ZN(n6530) );
  OAI21_X1 U7471 ( .B1(n6531), .B2(READREQUEST_REG_SCAN_IN), .A(n6530), .ZN(
        U3470) );
  NOR2_X1 U7472 ( .A1(READY_N), .A2(n6532), .ZN(n6541) );
  AOI211_X1 U7473 ( .C1(n6535), .C2(n6541), .A(n6534), .B(n6533), .ZN(n6549)
         );
  INV_X1 U7474 ( .A(n6536), .ZN(n6545) );
  OAI21_X1 U7475 ( .B1(n6539), .B2(n6538), .A(n6537), .ZN(n6542) );
  AOI21_X1 U7476 ( .B1(n6542), .B2(n6541), .A(n6540), .ZN(n6543) );
  AOI21_X1 U7477 ( .B1(n6545), .B2(n6544), .A(n6543), .ZN(n6548) );
  NOR2_X1 U7478 ( .A1(n6549), .A2(n6546), .ZN(n6547) );
  AOI22_X1 U7479 ( .A1(n6650), .A2(n6549), .B1(n6548), .B2(n6547), .ZN(U3472)
         );
  MUX2_X1 U7480 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6550), .Z(U3473) );
  INV_X1 U7481 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6657) );
  OAI22_X1 U7482 ( .A1(n6626), .A2(keyinput61), .B1(n6657), .B2(keyinput52), 
        .ZN(n6551) );
  AOI221_X1 U7483 ( .B1(n6626), .B2(keyinput61), .C1(keyinput52), .C2(n6657), 
        .A(n6551), .ZN(n6562) );
  INV_X1 U7484 ( .A(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n6554) );
  OAI22_X1 U7485 ( .A1(n6554), .A2(keyinput19), .B1(n6553), .B2(keyinput63), 
        .ZN(n6552) );
  AOI221_X1 U7486 ( .B1(n6554), .B2(keyinput19), .C1(keyinput63), .C2(n6553), 
        .A(n6552), .ZN(n6561) );
  OAI22_X1 U7487 ( .A1(n5142), .A2(keyinput48), .B1(n6556), .B2(keyinput28), 
        .ZN(n6555) );
  AOI221_X1 U7488 ( .B1(n5142), .B2(keyinput48), .C1(keyinput28), .C2(n6556), 
        .A(n6555), .ZN(n6560) );
  XNOR2_X1 U7489 ( .A(n3017), .B(keyinput34), .ZN(n6558) );
  XNOR2_X1 U7490 ( .A(keyinput41), .B(n6127), .ZN(n6557) );
  NOR2_X1 U7491 ( .A1(n6558), .A2(n6557), .ZN(n6559) );
  NAND4_X1 U7492 ( .A1(n6562), .A2(n6561), .A3(n6560), .A4(n6559), .ZN(n6743)
         );
  INV_X1 U7493 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n6564) );
  OAI22_X1 U7494 ( .A1(n6564), .A2(keyinput32), .B1(n6684), .B2(keyinput6), 
        .ZN(n6563) );
  AOI221_X1 U7495 ( .B1(n6564), .B2(keyinput32), .C1(keyinput6), .C2(n6684), 
        .A(n6563), .ZN(n6573) );
  OAI22_X1 U7496 ( .A1(n6567), .A2(keyinput23), .B1(n6566), .B2(keyinput3), 
        .ZN(n6565) );
  AOI221_X1 U7497 ( .B1(n6567), .B2(keyinput23), .C1(keyinput3), .C2(n6566), 
        .A(n6565), .ZN(n6572) );
  OAI22_X1 U7498 ( .A1(n4195), .A2(keyinput17), .B1(n6640), .B2(keyinput33), 
        .ZN(n6568) );
  AOI221_X1 U7499 ( .B1(n4195), .B2(keyinput17), .C1(keyinput33), .C2(n6640), 
        .A(n6568), .ZN(n6571) );
  OAI22_X1 U7500 ( .A1(n6624), .A2(keyinput56), .B1(n6614), .B2(keyinput15), 
        .ZN(n6569) );
  AOI221_X1 U7501 ( .B1(n6624), .B2(keyinput56), .C1(keyinput15), .C2(n6614), 
        .A(n6569), .ZN(n6570) );
  NAND4_X1 U7502 ( .A1(n6573), .A2(n6572), .A3(n6571), .A4(n6570), .ZN(n6742)
         );
  AOI22_X1 U7503 ( .A1(EAX_REG_12__SCAN_IN), .A2(keyinput24), .B1(
        PHYADDRPOINTER_REG_8__SCAN_IN), .B2(keyinput42), .ZN(n6574) );
  OAI221_X1 U7504 ( .B1(EAX_REG_12__SCAN_IN), .B2(keyinput24), .C1(
        PHYADDRPOINTER_REG_8__SCAN_IN), .C2(keyinput42), .A(n6574), .ZN(n6581)
         );
  AOI22_X1 U7505 ( .A1(DATAO_REG_6__SCAN_IN), .A2(keyinput53), .B1(DATAI_8_), 
        .B2(keyinput5), .ZN(n6575) );
  OAI221_X1 U7506 ( .B1(DATAO_REG_6__SCAN_IN), .B2(keyinput53), .C1(DATAI_8_), 
        .C2(keyinput5), .A(n6575), .ZN(n6580) );
  AOI22_X1 U7507 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(keyinput54), .B1(
        REIP_REG_8__SCAN_IN), .B2(keyinput51), .ZN(n6576) );
  OAI221_X1 U7508 ( .B1(DATAWIDTH_REG_23__SCAN_IN), .B2(keyinput54), .C1(
        REIP_REG_8__SCAN_IN), .C2(keyinput51), .A(n6576), .ZN(n6579) );
  AOI22_X1 U7509 ( .A1(REIP_REG_23__SCAN_IN), .A2(keyinput58), .B1(
        INSTQUEUE_REG_11__3__SCAN_IN), .B2(keyinput38), .ZN(n6577) );
  OAI221_X1 U7510 ( .B1(REIP_REG_23__SCAN_IN), .B2(keyinput58), .C1(
        INSTQUEUE_REG_11__3__SCAN_IN), .C2(keyinput38), .A(n6577), .ZN(n6578)
         );
  NOR4_X1 U7511 ( .A1(n6581), .A2(n6580), .A3(n6579), .A4(n6578), .ZN(n6610)
         );
  AOI22_X1 U7512 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(keyinput49), .B1(
        INSTADDRPOINTER_REG_16__SCAN_IN), .B2(keyinput50), .ZN(n6582) );
  OAI221_X1 U7513 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(keyinput49), .C1(
        INSTADDRPOINTER_REG_16__SCAN_IN), .C2(keyinput50), .A(n6582), .ZN(
        n6589) );
  AOI22_X1 U7514 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(keyinput7), .B1(
        INSTQUEUE_REG_7__0__SCAN_IN), .B2(keyinput55), .ZN(n6583) );
  OAI221_X1 U7515 ( .B1(INSTQUEUE_REG_7__5__SCAN_IN), .B2(keyinput7), .C1(
        INSTQUEUE_REG_7__0__SCAN_IN), .C2(keyinput55), .A(n6583), .ZN(n6588)
         );
  AOI22_X1 U7516 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(keyinput21), .B1(
        INSTQUEUE_REG_1__0__SCAN_IN), .B2(keyinput44), .ZN(n6584) );
  OAI221_X1 U7517 ( .B1(INSTQUEUE_REG_4__5__SCAN_IN), .B2(keyinput21), .C1(
        INSTQUEUE_REG_1__0__SCAN_IN), .C2(keyinput44), .A(n6584), .ZN(n6587)
         );
  AOI22_X1 U7518 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(keyinput30), .B1(
        INSTQUEUE_REG_11__6__SCAN_IN), .B2(keyinput39), .ZN(n6585) );
  OAI221_X1 U7519 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(keyinput30), 
        .C1(INSTQUEUE_REG_11__6__SCAN_IN), .C2(keyinput39), .A(n6585), .ZN(
        n6586) );
  NOR4_X1 U7520 ( .A1(n6589), .A2(n6588), .A3(n6587), .A4(n6586), .ZN(n6609)
         );
  AOI22_X1 U7521 ( .A1(REIP_REG_14__SCAN_IN), .A2(keyinput10), .B1(
        INSTQUEUE_REG_13__3__SCAN_IN), .B2(keyinput0), .ZN(n6590) );
  OAI221_X1 U7522 ( .B1(REIP_REG_14__SCAN_IN), .B2(keyinput10), .C1(
        INSTQUEUE_REG_13__3__SCAN_IN), .C2(keyinput0), .A(n6590), .ZN(n6597)
         );
  AOI22_X1 U7523 ( .A1(INSTQUEUE_REG_8__3__SCAN_IN), .A2(keyinput22), .B1(
        INSTQUEUE_REG_8__1__SCAN_IN), .B2(keyinput35), .ZN(n6591) );
  OAI221_X1 U7524 ( .B1(INSTQUEUE_REG_8__3__SCAN_IN), .B2(keyinput22), .C1(
        INSTQUEUE_REG_8__1__SCAN_IN), .C2(keyinput35), .A(n6591), .ZN(n6596)
         );
  AOI22_X1 U7525 ( .A1(DATAI_16_), .A2(keyinput43), .B1(
        INSTADDRPOINTER_REG_3__SCAN_IN), .B2(keyinput2), .ZN(n6592) );
  OAI221_X1 U7526 ( .B1(DATAI_16_), .B2(keyinput43), .C1(
        INSTADDRPOINTER_REG_3__SCAN_IN), .C2(keyinput2), .A(n6592), .ZN(n6595)
         );
  AOI22_X1 U7527 ( .A1(UWORD_REG_2__SCAN_IN), .A2(keyinput18), .B1(
        INSTADDRPOINTER_REG_17__SCAN_IN), .B2(keyinput37), .ZN(n6593) );
  OAI221_X1 U7528 ( .B1(UWORD_REG_2__SCAN_IN), .B2(keyinput18), .C1(
        INSTADDRPOINTER_REG_17__SCAN_IN), .C2(keyinput37), .A(n6593), .ZN(
        n6594) );
  NOR4_X1 U7529 ( .A1(n6597), .A2(n6596), .A3(n6595), .A4(n6594), .ZN(n6608)
         );
  AOI22_X1 U7530 ( .A1(REIP_REG_1__SCAN_IN), .A2(keyinput31), .B1(
        REIP_REG_22__SCAN_IN), .B2(keyinput60), .ZN(n6598) );
  OAI221_X1 U7531 ( .B1(REIP_REG_1__SCAN_IN), .B2(keyinput31), .C1(
        REIP_REG_22__SCAN_IN), .C2(keyinput60), .A(n6598), .ZN(n6606) );
  AOI22_X1 U7532 ( .A1(DATAO_REG_20__SCAN_IN), .A2(keyinput59), .B1(
        INSTQUEUE_REG_13__1__SCAN_IN), .B2(keyinput45), .ZN(n6599) );
  OAI221_X1 U7533 ( .B1(DATAO_REG_20__SCAN_IN), .B2(keyinput59), .C1(
        INSTQUEUE_REG_13__1__SCAN_IN), .C2(keyinput45), .A(n6599), .ZN(n6605)
         );
  AOI22_X1 U7534 ( .A1(DATAO_REG_26__SCAN_IN), .A2(keyinput16), .B1(
        DATAWIDTH_REG_26__SCAN_IN), .B2(keyinput1), .ZN(n6600) );
  OAI221_X1 U7535 ( .B1(DATAO_REG_26__SCAN_IN), .B2(keyinput16), .C1(
        DATAWIDTH_REG_26__SCAN_IN), .C2(keyinput1), .A(n6600), .ZN(n6604) );
  AOI22_X1 U7536 ( .A1(DATAO_REG_9__SCAN_IN), .A2(keyinput4), .B1(n6602), .B2(
        keyinput57), .ZN(n6601) );
  OAI221_X1 U7537 ( .B1(DATAO_REG_9__SCAN_IN), .B2(keyinput4), .C1(n6602), 
        .C2(keyinput57), .A(n6601), .ZN(n6603) );
  NOR4_X1 U7538 ( .A1(n6606), .A2(n6605), .A3(n6604), .A4(n6603), .ZN(n6607)
         );
  NAND4_X1 U7539 ( .A1(n6610), .A2(n6609), .A3(n6608), .A4(n6607), .ZN(n6741)
         );
  INV_X1 U7540 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n6612) );
  AOI22_X1 U7541 ( .A1(n6612), .A2(keyinput123), .B1(n6728), .B2(keyinput111), 
        .ZN(n6611) );
  OAI221_X1 U7542 ( .B1(n6612), .B2(keyinput123), .C1(n6728), .C2(keyinput111), 
        .A(n6611), .ZN(n6622) );
  AOI22_X1 U7543 ( .A1(n6725), .A2(keyinput90), .B1(keyinput79), .B2(n6614), 
        .ZN(n6613) );
  OAI221_X1 U7544 ( .B1(n6725), .B2(keyinput90), .C1(n6614), .C2(keyinput79), 
        .A(n6613), .ZN(n6621) );
  INV_X1 U7545 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n6715) );
  AOI22_X1 U7546 ( .A1(n6715), .A2(keyinput84), .B1(keyinput78), .B2(n6711), 
        .ZN(n6615) );
  OAI221_X1 U7547 ( .B1(n6715), .B2(keyinput84), .C1(n6711), .C2(keyinput78), 
        .A(n6615), .ZN(n6620) );
  INV_X1 U7548 ( .A(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n6616) );
  XOR2_X1 U7549 ( .A(n6616), .B(keyinput119), .Z(n6618) );
  XNOR2_X1 U7550 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput98), .ZN(
        n6617) );
  NAND2_X1 U7551 ( .A1(n6618), .A2(n6617), .ZN(n6619) );
  NOR4_X1 U7552 ( .A1(n6622), .A2(n6621), .A3(n6620), .A4(n6619), .ZN(n6666)
         );
  AOI22_X1 U7553 ( .A1(n6624), .A2(keyinput120), .B1(n4179), .B2(keyinput99), 
        .ZN(n6623) );
  OAI221_X1 U7554 ( .B1(n6624), .B2(keyinput120), .C1(n4179), .C2(keyinput99), 
        .A(n6623), .ZN(n6635) );
  AOI22_X1 U7555 ( .A1(n6626), .A2(keyinput125), .B1(keyinput89), .B2(n6721), 
        .ZN(n6625) );
  OAI221_X1 U7556 ( .B1(n6626), .B2(keyinput125), .C1(n6721), .C2(keyinput89), 
        .A(n6625), .ZN(n6634) );
  AOI22_X1 U7557 ( .A1(n6629), .A2(keyinput88), .B1(keyinput118), .B2(n6628), 
        .ZN(n6627) );
  OAI221_X1 U7558 ( .B1(n6629), .B2(keyinput88), .C1(n6628), .C2(keyinput118), 
        .A(n6627), .ZN(n6633) );
  INV_X1 U7559 ( .A(LWORD_REG_2__SCAN_IN), .ZN(n6709) );
  AOI22_X1 U7560 ( .A1(n6709), .A2(keyinput75), .B1(keyinput80), .B2(n6631), 
        .ZN(n6630) );
  OAI221_X1 U7561 ( .B1(n6709), .B2(keyinput75), .C1(n6631), .C2(keyinput80), 
        .A(n6630), .ZN(n6632) );
  NOR4_X1 U7562 ( .A1(n6635), .A2(n6634), .A3(n6633), .A4(n6632), .ZN(n6665)
         );
  AOI22_X1 U7563 ( .A1(n4195), .A2(keyinput81), .B1(keyinput86), .B2(n4191), 
        .ZN(n6636) );
  OAI221_X1 U7564 ( .B1(n4195), .B2(keyinput81), .C1(n4191), .C2(keyinput86), 
        .A(n6636), .ZN(n6647) );
  INV_X1 U7565 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n6638) );
  AOI22_X1 U7566 ( .A1(n6638), .A2(keyinput117), .B1(keyinput104), .B2(n6708), 
        .ZN(n6637) );
  OAI221_X1 U7567 ( .B1(n6638), .B2(keyinput117), .C1(n6708), .C2(keyinput104), 
        .A(n6637), .ZN(n6646) );
  AOI22_X1 U7568 ( .A1(n6641), .A2(keyinput101), .B1(keyinput97), .B2(n6640), 
        .ZN(n6639) );
  OAI221_X1 U7569 ( .B1(n6641), .B2(keyinput101), .C1(n6640), .C2(keyinput97), 
        .A(n6639), .ZN(n6645) );
  INV_X1 U7570 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n6643) );
  AOI22_X1 U7571 ( .A1(n6730), .A2(keyinput93), .B1(n6643), .B2(keyinput108), 
        .ZN(n6642) );
  OAI221_X1 U7572 ( .B1(n6730), .B2(keyinput93), .C1(n6643), .C2(keyinput108), 
        .A(n6642), .ZN(n6644) );
  NOR4_X1 U7573 ( .A1(n6647), .A2(n6646), .A3(n6645), .A4(n6644), .ZN(n6664)
         );
  AOI22_X1 U7574 ( .A1(n6650), .A2(keyinput113), .B1(n6649), .B2(keyinput94), 
        .ZN(n6648) );
  OAI221_X1 U7575 ( .B1(n6650), .B2(keyinput113), .C1(n6649), .C2(keyinput94), 
        .A(n6648), .ZN(n6662) );
  AOI22_X1 U7576 ( .A1(n6653), .A2(keyinput66), .B1(keyinput95), .B2(n6652), 
        .ZN(n6651) );
  OAI221_X1 U7577 ( .B1(n6653), .B2(keyinput66), .C1(n6652), .C2(keyinput95), 
        .A(n6651), .ZN(n6661) );
  AOI22_X1 U7578 ( .A1(n5620), .A2(keyinput74), .B1(n6655), .B2(keyinput122), 
        .ZN(n6654) );
  OAI221_X1 U7579 ( .B1(n5620), .B2(keyinput74), .C1(n6655), .C2(keyinput122), 
        .A(n6654), .ZN(n6660) );
  AOI22_X1 U7580 ( .A1(n6658), .A2(keyinput106), .B1(keyinput116), .B2(n6657), 
        .ZN(n6656) );
  OAI221_X1 U7581 ( .B1(n6658), .B2(keyinput106), .C1(n6657), .C2(keyinput116), 
        .A(n6656), .ZN(n6659) );
  NOR4_X1 U7582 ( .A1(n6662), .A2(n6661), .A3(n6660), .A4(n6659), .ZN(n6663)
         );
  NAND4_X1 U7583 ( .A1(n6666), .A2(n6665), .A3(n6664), .A4(n6663), .ZN(n6739)
         );
  AOI22_X1 U7584 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(keyinput96), .B1(
        INSTQUEUE_REG_4__5__SCAN_IN), .B2(keyinput85), .ZN(n6667) );
  OAI221_X1 U7585 ( .B1(INSTQUEUE_REG_3__3__SCAN_IN), .B2(keyinput96), .C1(
        INSTQUEUE_REG_4__5__SCAN_IN), .C2(keyinput85), .A(n6667), .ZN(n6674)
         );
  AOI22_X1 U7586 ( .A1(UWORD_REG_2__SCAN_IN), .A2(keyinput82), .B1(DATAI_16_), 
        .B2(keyinput107), .ZN(n6668) );
  OAI221_X1 U7587 ( .B1(UWORD_REG_2__SCAN_IN), .B2(keyinput82), .C1(DATAI_16_), 
        .C2(keyinput107), .A(n6668), .ZN(n6673) );
  AOI22_X1 U7588 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(keyinput65), .B1(
        DATAO_REG_14__SCAN_IN), .B2(keyinput100), .ZN(n6669) );
  OAI221_X1 U7589 ( .B1(DATAWIDTH_REG_26__SCAN_IN), .B2(keyinput65), .C1(
        DATAO_REG_14__SCAN_IN), .C2(keyinput100), .A(n6669), .ZN(n6672) );
  AOI22_X1 U7590 ( .A1(REIP_REG_8__SCAN_IN), .A2(keyinput115), .B1(
        INSTQUEUE_REG_11__6__SCAN_IN), .B2(keyinput103), .ZN(n6670) );
  OAI221_X1 U7591 ( .B1(REIP_REG_8__SCAN_IN), .B2(keyinput115), .C1(
        INSTQUEUE_REG_11__6__SCAN_IN), .C2(keyinput103), .A(n6670), .ZN(n6671)
         );
  NOR4_X1 U7592 ( .A1(n6674), .A2(n6673), .A3(n6672), .A4(n6671), .ZN(n6703)
         );
  AOI22_X1 U7593 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(keyinput87), .B1(
        INSTQUEUE_REG_11__3__SCAN_IN), .B2(keyinput102), .ZN(n6675) );
  OAI221_X1 U7594 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(keyinput87), 
        .C1(INSTQUEUE_REG_11__3__SCAN_IN), .C2(keyinput102), .A(n6675), .ZN(
        n6682) );
  AOI22_X1 U7595 ( .A1(EAX_REG_13__SCAN_IN), .A2(keyinput67), .B1(
        INSTQUEUE_REG_9__3__SCAN_IN), .B2(keyinput83), .ZN(n6676) );
  OAI221_X1 U7596 ( .B1(EAX_REG_13__SCAN_IN), .B2(keyinput67), .C1(
        INSTQUEUE_REG_9__3__SCAN_IN), .C2(keyinput83), .A(n6676), .ZN(n6681)
         );
  AOI22_X1 U7597 ( .A1(DATAO_REG_9__SCAN_IN), .A2(keyinput68), .B1(DATAI_30_), 
        .B2(keyinput126), .ZN(n6677) );
  OAI221_X1 U7598 ( .B1(DATAO_REG_9__SCAN_IN), .B2(keyinput68), .C1(DATAI_30_), 
        .C2(keyinput126), .A(n6677), .ZN(n6680) );
  AOI22_X1 U7599 ( .A1(REIP_REG_27__SCAN_IN), .A2(keyinput92), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput127), .ZN(n6678) );
  OAI221_X1 U7600 ( .B1(REIP_REG_27__SCAN_IN), .B2(keyinput92), .C1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .C2(keyinput127), .A(n6678), .ZN(
        n6679) );
  NOR4_X1 U7601 ( .A1(n6682), .A2(n6681), .A3(n6680), .A4(n6679), .ZN(n6702)
         );
  AOI22_X1 U7602 ( .A1(DATAI_8_), .A2(keyinput69), .B1(n6684), .B2(keyinput70), 
        .ZN(n6683) );
  OAI221_X1 U7603 ( .B1(DATAI_8_), .B2(keyinput69), .C1(n6684), .C2(keyinput70), .A(n6683), .ZN(n6691) );
  AOI22_X1 U7604 ( .A1(REIP_REG_22__SCAN_IN), .A2(keyinput124), .B1(
        INSTQUEUE_REG_6__7__SCAN_IN), .B2(keyinput91), .ZN(n6685) );
  OAI221_X1 U7605 ( .B1(REIP_REG_22__SCAN_IN), .B2(keyinput124), .C1(
        INSTQUEUE_REG_6__7__SCAN_IN), .C2(keyinput91), .A(n6685), .ZN(n6690)
         );
  AOI22_X1 U7606 ( .A1(n6724), .A2(keyinput76), .B1(keyinput105), .B2(n6127), 
        .ZN(n6686) );
  OAI221_X1 U7607 ( .B1(n6724), .B2(keyinput76), .C1(n6127), .C2(keyinput105), 
        .A(n6686), .ZN(n6689) );
  AOI22_X1 U7608 ( .A1(n5142), .A2(keyinput112), .B1(n6714), .B2(keyinput110), 
        .ZN(n6687) );
  OAI221_X1 U7609 ( .B1(n5142), .B2(keyinput112), .C1(n6714), .C2(keyinput110), 
        .A(n6687), .ZN(n6688) );
  NOR4_X1 U7610 ( .A1(n6691), .A2(n6690), .A3(n6689), .A4(n6688), .ZN(n6701)
         );
  AOI22_X1 U7611 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(keyinput64), .B1(
        INSTQUEUE_REG_13__1__SCAN_IN), .B2(keyinput109), .ZN(n6692) );
  OAI221_X1 U7612 ( .B1(INSTQUEUE_REG_13__3__SCAN_IN), .B2(keyinput64), .C1(
        INSTQUEUE_REG_13__1__SCAN_IN), .C2(keyinput109), .A(n6692), .ZN(n6699)
         );
  AOI22_X1 U7613 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(keyinput71), .B1(
        INSTQUEUE_REG_8__5__SCAN_IN), .B2(keyinput77), .ZN(n6693) );
  OAI221_X1 U7614 ( .B1(INSTQUEUE_REG_7__5__SCAN_IN), .B2(keyinput71), .C1(
        INSTQUEUE_REG_8__5__SCAN_IN), .C2(keyinput77), .A(n6693), .ZN(n6698)
         );
  AOI22_X1 U7615 ( .A1(LWORD_REG_9__SCAN_IN), .A2(keyinput121), .B1(DATAI_6_), 
        .B2(keyinput73), .ZN(n6694) );
  OAI221_X1 U7616 ( .B1(LWORD_REG_9__SCAN_IN), .B2(keyinput121), .C1(DATAI_6_), 
        .C2(keyinput73), .A(n6694), .ZN(n6697) );
  AOI22_X1 U7617 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(keyinput114), 
        .B1(INSTQUEUE_REG_14__7__SCAN_IN), .B2(keyinput72), .ZN(n6695) );
  OAI221_X1 U7618 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(keyinput114), 
        .C1(INSTQUEUE_REG_14__7__SCAN_IN), .C2(keyinput72), .A(n6695), .ZN(
        n6696) );
  NOR4_X1 U7619 ( .A1(n6699), .A2(n6698), .A3(n6697), .A4(n6696), .ZN(n6700)
         );
  NAND4_X1 U7620 ( .A1(n6703), .A2(n6702), .A3(n6701), .A4(n6700), .ZN(n6738)
         );
  INV_X1 U7621 ( .A(DATAI_30_), .ZN(n6705) );
  AOI22_X1 U7622 ( .A1(n6706), .A2(keyinput9), .B1(n6705), .B2(keyinput62), 
        .ZN(n6704) );
  OAI221_X1 U7623 ( .B1(n6706), .B2(keyinput9), .C1(n6705), .C2(keyinput62), 
        .A(n6704), .ZN(n6719) );
  AOI22_X1 U7624 ( .A1(n6709), .A2(keyinput11), .B1(keyinput40), .B2(n6708), 
        .ZN(n6707) );
  OAI221_X1 U7625 ( .B1(n6709), .B2(keyinput11), .C1(n6708), .C2(keyinput40), 
        .A(n6707), .ZN(n6718) );
  AOI22_X1 U7626 ( .A1(n6712), .A2(keyinput36), .B1(keyinput14), .B2(n6711), 
        .ZN(n6710) );
  OAI221_X1 U7627 ( .B1(n6712), .B2(keyinput36), .C1(n6711), .C2(keyinput14), 
        .A(n6710), .ZN(n6717) );
  AOI22_X1 U7628 ( .A1(n6715), .A2(keyinput20), .B1(keyinput46), .B2(n6714), 
        .ZN(n6713) );
  OAI221_X1 U7629 ( .B1(n6715), .B2(keyinput20), .C1(n6714), .C2(keyinput46), 
        .A(n6713), .ZN(n6716) );
  NOR4_X1 U7630 ( .A1(n6719), .A2(n6718), .A3(n6717), .A4(n6716), .ZN(n6737)
         );
  AOI22_X1 U7631 ( .A1(n6722), .A2(keyinput13), .B1(keyinput25), .B2(n6721), 
        .ZN(n6720) );
  OAI221_X1 U7632 ( .B1(n6722), .B2(keyinput13), .C1(n6721), .C2(keyinput25), 
        .A(n6720), .ZN(n6735) );
  AOI22_X1 U7633 ( .A1(n6725), .A2(keyinput26), .B1(n6724), .B2(keyinput12), 
        .ZN(n6723) );
  OAI221_X1 U7634 ( .B1(n6725), .B2(keyinput26), .C1(n6724), .C2(keyinput12), 
        .A(n6723), .ZN(n6734) );
  INV_X1 U7635 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n6727) );
  AOI22_X1 U7636 ( .A1(n6728), .A2(keyinput47), .B1(n6727), .B2(keyinput27), 
        .ZN(n6726) );
  OAI221_X1 U7637 ( .B1(n6728), .B2(keyinput47), .C1(n6727), .C2(keyinput27), 
        .A(n6726), .ZN(n6733) );
  INV_X1 U7638 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6731) );
  AOI22_X1 U7639 ( .A1(n6731), .A2(keyinput8), .B1(keyinput29), .B2(n6730), 
        .ZN(n6729) );
  OAI221_X1 U7640 ( .B1(n6731), .B2(keyinput8), .C1(n6730), .C2(keyinput29), 
        .A(n6729), .ZN(n6732) );
  NOR4_X1 U7641 ( .A1(n6735), .A2(n6734), .A3(n6733), .A4(n6732), .ZN(n6736)
         );
  OAI211_X1 U7642 ( .C1(n6739), .C2(n6738), .A(n6737), .B(n6736), .ZN(n6740)
         );
  NOR4_X1 U7643 ( .A1(n6743), .A2(n6742), .A3(n6741), .A4(n6740), .ZN(n6753)
         );
  INV_X1 U7644 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n6749) );
  INV_X1 U7645 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6744) );
  OR2_X1 U7646 ( .A1(n6745), .A2(n6744), .ZN(n6748) );
  NAND2_X1 U7647 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n6746), .ZN(n6747) );
  OAI211_X1 U7648 ( .C1(n6750), .C2(n6749), .A(n6748), .B(n6747), .ZN(n6751)
         );
  INV_X1 U7649 ( .A(n6751), .ZN(n6752) );
  XNOR2_X1 U7650 ( .A(n6753), .B(n6752), .ZN(U2902) );
  AND2_X1 U3574 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4007) );
  AND2_X2 U3770 ( .A1(n3022), .A2(n3898), .ZN(n3196) );
  NOR2_X2 U34620 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3023) );
  CLKBUF_X1 U3475 ( .A(n3733), .Z(n4291) );
  CLKBUF_X2 U3476 ( .A(n3780), .Z(n3002) );
  CLKBUF_X1 U3773 ( .A(n4291), .Z(n2995) );
endmodule

