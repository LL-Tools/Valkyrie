

module b14_C_AntiSAT_k_256_4 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2350, n2351, n2352,
         n2353, n2354, n2355, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092;

  INV_X2 U2483 ( .A(n4617), .ZN(n4619) );
  OR2_X1 U2484 ( .A1(n3775), .A2(n3986), .ZN(n2245) );
  AOI211_X1 U2485 ( .C1(n3746), .C2(n3752), .A(n3859), .B(n3854), .ZN(n3755)
         );
  OR2_X1 U2486 ( .A1(n2588), .A2(n2587), .ZN(n2589) );
  OAI21_X1 U2487 ( .B1(n3430), .B2(n3432), .A(n3431), .ZN(n3547) );
  NAND2_X1 U2488 ( .A1(n2330), .A2(n2256), .ZN(n3569) );
  AND2_X1 U2489 ( .A1(n4228), .A2(n4223), .ZN(n2585) );
  NAND2_X1 U2490 ( .A1(n3219), .A2(n2850), .ZN(n3218) );
  INV_X1 U2491 ( .A(n4245), .ZN(n2242) );
  NOR2_X1 U2492 ( .A1(n4266), .A2(n4389), .ZN(n2241) );
  OR2_X1 U2493 ( .A1(n4598), .A2(n3702), .ZN(n3308) );
  INV_X1 U2494 ( .A(n4251), .ZN(n4394) );
  AOI21_X1 U2495 ( .B1(n3185), .B2(n3184), .A(n2260), .ZN(n3696) );
  AND2_X1 U2496 ( .A1(n2828), .A2(n2326), .ZN(n2260) );
  INV_X1 U2497 ( .A(n3069), .ZN(n3065) );
  CLKBUF_X2 U2498 ( .A(n3062), .Z(n2247) );
  OR2_X2 U2499 ( .A1(n2822), .A2(n2813), .ZN(n3071) );
  CLKBUF_X2 U2500 ( .A(n2398), .Z(n2734) );
  CLKBUF_X2 U2502 ( .A(n3741), .Z(n2795) );
  INV_X1 U2503 ( .A(n3118), .ZN(n2822) );
  AND2_X1 U2504 ( .A1(n3883), .A2(n4605), .ZN(n4399) );
  OR2_X1 U2505 ( .A1(n2747), .A2(IR_REG_25__SCAN_IN), .ZN(n2257) );
  OAI21_X1 U2506 ( .B1(n2601), .B2(IR_REG_18__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2680) );
  INV_X2 U2507 ( .A(IR_REG_31__SCAN_IN), .ZN(n2690) );
  NAND2_X1 U2508 ( .A1(n2374), .A2(n3563), .ZN(n2376) );
  BUF_X2 U2509 ( .A(IR_REG_0__SCAN_IN), .Z(n2244) );
  NAND2_X1 U2510 ( .A1(n2276), .A2(n2362), .ZN(n2479) );
  NOR2_X1 U2511 ( .A1(n2242), .A2(n2241), .ZN(n2570) );
  AOI21_X1 U2512 ( .B1(n2591), .B2(n2353), .A(n2243), .ZN(n4183) );
  NOR2_X1 U2513 ( .A1(n4181), .A2(n4186), .ZN(n2243) );
  OAI21_X2 U2514 ( .B1(n3501), .B2(n2283), .A(n2281), .ZN(n3555) );
  AOI21_X2 U2515 ( .B1(n3601), .B2(n3041), .A(n2261), .ZN(n3665) );
  NAND2_X1 U2516 ( .A1(n2864), .A2(n2329), .ZN(n2330) );
  NAND2_X2 U2517 ( .A1(n2964), .A2(n2338), .ZN(n2337) );
  NAND2_X2 U2518 ( .A1(n2267), .A2(n2292), .ZN(n3648) );
  NAND2_X2 U2519 ( .A1(n3061), .A2(n3718), .ZN(n3579) );
  NOR2_X1 U2520 ( .A1(n4206), .A2(n2575), .ZN(n2588) );
  NAND3_X1 U2521 ( .A1(n2262), .A2(n2342), .A3(n2246), .ZN(n2341) );
  INV_X2 U2522 ( .A(n2812), .ZN(n3177) );
  NAND3_X2 U2523 ( .A1(n2391), .A2(n2392), .A3(n2390), .ZN(n2812) );
  OAI21_X2 U2524 ( .B1(n2801), .B2(n4292), .A(n2245), .ZN(n4000) );
  NOR2_X2 U2525 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2347)
         );
  INV_X1 U2526 ( .A(IR_REG_3__SCAN_IN), .ZN(n2410) );
  INV_X1 U2527 ( .A(n4399), .ZN(n4678) );
  AND2_X1 U2528 ( .A1(n2776), .A2(n4080), .ZN(n4075) );
  INV_X1 U2529 ( .A(n3906), .ZN(U4043) );
  AND4_X1 U2530 ( .A1(n2548), .A2(n2365), .A3(n2364), .A4(n2681), .ZN(n2246)
         );
  INV_X8 U2531 ( .A(n3071), .ZN(n2252) );
  AND2_X1 U2532 ( .A1(n2813), .A2(n3118), .ZN(n3062) );
  AND2_X2 U2533 ( .A1(n2249), .A2(n2344), .ZN(n2688) );
  NAND2_X1 U2534 ( .A1(n4243), .A2(n3748), .ZN(n4237) );
  NAND2_X1 U2535 ( .A1(n2714), .A2(n2713), .ZN(n4243) );
  NAND2_X1 U2536 ( .A1(n2698), .A2(n3232), .ZN(n3239) );
  NAND2_X1 U2537 ( .A1(n2278), .A2(n3572), .ZN(n3464) );
  INV_X1 U2538 ( .A(n3907), .ZN(n3243) );
  NAND4_X1 U2539 ( .A1(n2557), .A2(n2556), .A3(n2555), .A4(n2554), .ZN(n4266)
         );
  NAND4_X1 U2540 ( .A1(n2430), .A2(n2429), .A3(n2428), .A4(n2427), .ZN(n3390)
         );
  BUF_X2 U2541 ( .A(n2394), .Z(n3741) );
  INV_X2 U2542 ( .A(n2417), .ZN(n2389) );
  CLKBUF_X3 U2543 ( .A(n2395), .Z(n2248) );
  NAND2_X1 U2544 ( .A1(n2354), .A2(n2731), .ZN(n2793) );
  NAND2_X1 U2545 ( .A1(n2730), .A2(n2729), .ZN(n4021) );
  AND2_X1 U2546 ( .A1(n2288), .A2(n3687), .ZN(n3695) );
  OR2_X1 U2547 ( .A1(n3631), .A2(n3602), .ZN(n3686) );
  AOI21_X1 U2548 ( .B1(n4053), .B2(n2650), .A(n2649), .ZN(n4041) );
  AOI21_X2 U2549 ( .B1(n4073), .B2(n2641), .A(n2640), .ZN(n4053) );
  NAND2_X1 U2550 ( .A1(n2254), .A2(n2264), .ZN(n3998) );
  NAND2_X1 U2551 ( .A1(n2705), .A2(n3845), .ZN(n3475) );
  OR2_X1 U2552 ( .A1(n2576), .A2(n2590), .ZN(n4180) );
  OR2_X1 U2553 ( .A1(n2590), .A2(n2589), .ZN(n4181) );
  AND2_X1 U2554 ( .A1(n2574), .A2(n4225), .ZN(n4206) );
  OR2_X1 U2555 ( .A1(n2573), .A2(n4222), .ZN(n4225) );
  AND2_X2 U2556 ( .A1(n3094), .A2(STATE_REG_SCAN_IN), .ZN(n3736) );
  NAND2_X1 U2557 ( .A1(n2695), .A2(n3818), .ZN(n3797) );
  NAND4_X1 U2558 ( .A1(n2567), .A2(n2566), .A3(n2565), .A4(n2564), .ZN(n4251)
         );
  NAND2_X2 U2559 ( .A1(n2419), .A2(n2418), .ZN(n2842) );
  NAND4_X2 U2560 ( .A1(n2408), .A2(n2407), .A3(n2406), .A4(n2405), .ZN(n3905)
         );
  NAND4_X2 U2561 ( .A1(n2381), .A2(n2380), .A3(n2379), .A4(n2378), .ZN(n2821)
         );
  NAND2_X2 U2562 ( .A1(n2813), .A2(n3101), .ZN(n3069) );
  BUF_X1 U2563 ( .A(n2687), .Z(n3883) );
  INV_X1 U2564 ( .A(n3328), .ZN(n3303) );
  XNOR2_X1 U2565 ( .A(n2680), .B(IR_REG_19__SCAN_IN), .ZN(n4485) );
  INV_X1 U2566 ( .A(n3181), .ZN(n4607) );
  NAND3_X1 U2567 ( .A1(n4481), .A2(n4480), .A3(n2754), .ZN(n3118) );
  NAND2_X1 U2568 ( .A1(n2371), .A2(IR_REG_31__SCAN_IN), .ZN(n2370) );
  MUX2_X1 U2569 ( .A(IR_REG_31__SCAN_IN), .B(n2373), .S(IR_REG_29__SCAN_IN), 
        .Z(n2374) );
  AND2_X1 U2570 ( .A1(n2546), .A2(n2352), .ZN(n2536) );
  NOR2_X1 U2571 ( .A1(n2568), .A2(IR_REG_14__SCAN_IN), .ZN(n2546) );
  NAND2_X1 U2572 ( .A1(n2294), .A2(n2364), .ZN(n2568) );
  INV_X1 U2573 ( .A(n2524), .ZN(n2294) );
  INV_X1 U2574 ( .A(n2479), .ZN(n2274) );
  NOR2_X1 U2575 ( .A1(n2341), .A2(IR_REG_21__SCAN_IN), .ZN(n2275) );
  AND2_X1 U2576 ( .A1(n2363), .A2(n2343), .ZN(n2342) );
  AND2_X1 U2577 ( .A1(n2347), .A2(n2328), .ZN(n2327) );
  NOR3_X1 U2578 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .A3(
        IR_REG_6__SCAN_IN), .ZN(n2361) );
  INV_X1 U2579 ( .A(IR_REG_17__SCAN_IN), .ZN(n2535) );
  INV_X1 U2580 ( .A(IR_REG_16__SCAN_IN), .ZN(n4806) );
  NOR2_X1 U2581 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2363)
         );
  INV_X1 U2582 ( .A(IR_REG_15__SCAN_IN), .ZN(n2548) );
  INV_X1 U2583 ( .A(n2250), .ZN(n2409) );
  AND3_X2 U2584 ( .A1(n2274), .A2(n2275), .A3(n2684), .ZN(n2249) );
  AND2_X2 U2585 ( .A1(n2402), .A2(n2360), .ZN(n2250) );
  OR2_X2 U2586 ( .A1(n4021), .A2(n4020), .ZN(n2354) );
  NOR2_X1 U2587 ( .A1(n4478), .A2(n2376), .ZN(n2395) );
  NOR2_X1 U2588 ( .A1(n4478), .A2(n2376), .ZN(n2251) );
  OR2_X2 U2589 ( .A1(n4034), .A2(n3872), .ZN(n2730) );
  OR2_X1 U2590 ( .A1(n2249), .A2(n2690), .ZN(n2755) );
  AOI21_X2 U2591 ( .B1(n4085), .B2(n2635), .A(n2634), .ZN(n4073) );
  NAND2_X2 U2592 ( .A1(n4235), .A2(n3753), .ZN(n4161) );
  NAND2_X2 U2593 ( .A1(n4237), .A2(n4236), .ZN(n4235) );
  NAND2_X2 U2594 ( .A1(n2700), .A2(n3828), .ZN(n3296) );
  NAND2_X2 U2595 ( .A1(n3177), .A2(n4587), .ZN(n2695) );
  AOI22_X2 U2596 ( .A1(n4041), .A2(n2659), .B1(n3643), .B2(n4048), .ZN(n4019)
         );
  XNOR2_X2 U2597 ( .A(n2792), .B(n2791), .ZN(n3991) );
  AOI21_X2 U2598 ( .B1(n3456), .B2(n3844), .A(n3840), .ZN(n3440) );
  OAI21_X2 U2599 ( .B1(n3401), .B2(n2704), .A(n3839), .ZN(n3456) );
  AOI21_X1 U2600 ( .B1(n2812), .B2(n2840), .A(n2817), .ZN(n2827) );
  AND2_X4 U2601 ( .A1(n3062), .A2(n4678), .ZN(n2840) );
  OAI22_X2 U2602 ( .A1(n3474), .A2(n2492), .B1(n3476), .B2(n3901), .ZN(n3525)
         );
  OAI21_X2 U2603 ( .B1(n3442), .B2(n2483), .A(n2482), .ZN(n3474) );
  INV_X1 U2604 ( .A(IR_REG_9__SCAN_IN), .ZN(n2362) );
  INV_X1 U2605 ( .A(n2477), .ZN(n2276) );
  AOI21_X1 U2606 ( .B1(n2337), .B2(n2334), .A(n2333), .ZN(n3014) );
  NAND2_X1 U2607 ( .A1(n2651), .A2(REG3_REG_26__SCAN_IN), .ZN(n2669) );
  NAND2_X1 U2608 ( .A1(n3144), .A2(n3143), .ZN(n3146) );
  XNOR2_X1 U2609 ( .A(n3349), .B(n4631), .ZN(n4554) );
  AND2_X1 U2610 ( .A1(n4322), .A2(n2648), .ZN(n2649) );
  AND2_X1 U2611 ( .A1(n3890), .A2(n3097), .ZN(n4605) );
  AND2_X1 U2612 ( .A1(n2676), .A2(n2675), .ZN(n4315) );
  NAND2_X1 U2613 ( .A1(n2690), .A2(IR_REG_1__SCAN_IN), .ZN(n2307) );
  XNOR2_X1 U2614 ( .A(n3146), .B(n4493), .ZN(n3208) );
  NAND2_X1 U2615 ( .A1(n4582), .A2(n4583), .ZN(n4580) );
  INV_X1 U2616 ( .A(IR_REG_14__SCAN_IN), .ZN(n2365) );
  INV_X1 U2617 ( .A(IR_REG_19__SCAN_IN), .ZN(n2679) );
  INV_X1 U2618 ( .A(IR_REG_10__SCAN_IN), .ZN(n2343) );
  XNOR2_X1 U2619 ( .A(n2839), .B(n3069), .ZN(n2847) );
  NAND2_X1 U2620 ( .A1(n2838), .A2(n2837), .ZN(n2839) );
  NAND2_X1 U2621 ( .A1(n3622), .A2(n3623), .ZN(n3601) );
  NAND2_X1 U2622 ( .A1(n4313), .A2(n2252), .ZN(n3052) );
  NAND2_X1 U2623 ( .A1(n2252), .A2(n4321), .ZN(n3054) );
  NAND2_X1 U2624 ( .A1(n2252), .A2(n2942), .ZN(n2943) );
  OR2_X1 U2625 ( .A1(n3939), .A2(n4487), .ZN(n2314) );
  NOR2_X1 U2626 ( .A1(n2253), .A2(n2345), .ZN(n2344) );
  NAND2_X1 U2627 ( .A1(n2800), .A2(n2366), .ZN(n2345) );
  NAND2_X1 U2628 ( .A1(n2308), .A2(IR_REG_31__SCAN_IN), .ZN(n2306) );
  NAND2_X1 U2629 ( .A1(n2308), .A2(n2301), .ZN(n2300) );
  NOR2_X1 U2630 ( .A1(n3286), .A2(n2331), .ZN(n2329) );
  NOR2_X1 U2631 ( .A1(n2631), .A2(n3606), .ZN(n2636) );
  NAND2_X1 U2632 ( .A1(n2336), .A2(n2971), .ZN(n2335) );
  INV_X1 U2633 ( .A(n3709), .ZN(n2336) );
  AOI21_X1 U2634 ( .B1(n2821), .B2(n2252), .A(n2820), .ZN(n2824) );
  XNOR2_X1 U2635 ( .A(n2845), .B(n3069), .ZN(n2853) );
  NAND2_X1 U2636 ( .A1(n2844), .A2(n2843), .ZN(n2845) );
  INV_X1 U2637 ( .A(n3062), .ZN(n3068) );
  NAND2_X1 U2638 ( .A1(n3502), .A2(n3503), .ZN(n2284) );
  INV_X1 U2639 ( .A(n3539), .ZN(n2285) );
  AND2_X1 U2640 ( .A1(n2271), .A2(n2963), .ZN(n2338) );
  AND2_X1 U2641 ( .A1(n4483), .A2(n4482), .ZN(n3126) );
  NAND2_X1 U2642 ( .A1(n3555), .A2(n3556), .ZN(n2934) );
  NAND2_X1 U2643 ( .A1(n2303), .A2(n3157), .ZN(n2302) );
  INV_X1 U2644 ( .A(n2307), .ZN(n2303) );
  NAND2_X1 U2645 ( .A1(n3210), .A2(REG1_REG_4__SCAN_IN), .ZN(n3209) );
  OR2_X1 U2646 ( .A1(n3339), .A2(n3338), .ZN(n3340) );
  NAND2_X1 U2647 ( .A1(n4541), .A2(n2309), .ZN(n3374) );
  OR2_X1 U2648 ( .A1(n4549), .A2(n4846), .ZN(n2309) );
  NAND2_X1 U2649 ( .A1(n4544), .A2(n3348), .ZN(n3349) );
  NAND2_X1 U2650 ( .A1(n4554), .A2(REG2_REG_12__SCAN_IN), .ZN(n4553) );
  NAND2_X1 U2651 ( .A1(n4569), .A2(n3376), .ZN(n3420) );
  NAND2_X1 U2652 ( .A1(n2314), .A2(n2313), .ZN(n3940) );
  NAND2_X1 U2653 ( .A1(n3939), .A2(n4487), .ZN(n2313) );
  NOR2_X1 U2654 ( .A1(n3940), .A2(REG1_REG_16__SCAN_IN), .ZN(n3959) );
  NOR2_X1 U2655 ( .A1(n4576), .A2(n4577), .ZN(n4575) );
  AND2_X1 U2656 ( .A1(n4335), .A2(n2775), .ZN(n2634) );
  NAND2_X1 U2657 ( .A1(n4008), .A2(n3992), .ZN(n2277) );
  NAND2_X1 U2658 ( .A1(n4484), .A2(n4605), .ZN(n4288) );
  NAND2_X1 U2659 ( .A1(n2686), .A2(n3981), .ZN(n4594) );
  NAND4_X1 U2660 ( .A1(n3078), .A2(n3235), .A3(n3233), .A4(n3091), .ZN(n2781)
         );
  NAND2_X1 U2661 ( .A1(n2752), .A2(n2754), .ZN(n3122) );
  XNOR2_X1 U2662 ( .A(n2685), .B(n2684), .ZN(n3890) );
  NOR2_X1 U2663 ( .A1(n2479), .A2(IR_REG_10__SCAN_IN), .ZN(n2499) );
  INV_X1 U2664 ( .A(n2942), .ZN(n4274) );
  INV_X1 U2665 ( .A(n5078), .ZN(n2907) );
  XNOR2_X1 U2666 ( .A(n2326), .B(n2827), .ZN(n3185) );
  AND2_X1 U2667 ( .A1(n2652), .A2(n2669), .ZN(n4045) );
  INV_X1 U2668 ( .A(n4485), .ZN(n3981) );
  OAI211_X1 U2669 ( .C1(n4496), .C2(REG2_REG_1__SCAN_IN), .A(n3139), .B(n3196), 
        .ZN(n3918) );
  NAND2_X1 U2670 ( .A1(n3164), .A2(n3165), .ZN(n3362) );
  OAI21_X1 U2671 ( .B1(n3208), .B2(n3145), .A(n3147), .ZN(n3153) );
  XNOR2_X1 U2672 ( .A(n3374), .B(n4631), .ZN(n4559) );
  NAND2_X1 U2673 ( .A1(n4559), .A2(REG1_REG_12__SCAN_IN), .ZN(n4558) );
  OR2_X1 U2674 ( .A1(n3419), .A2(n3418), .ZN(n3945) );
  XNOR2_X1 U2675 ( .A(n3951), .B(n2316), .ZN(n3946) );
  INV_X1 U2676 ( .A(n4487), .ZN(n2316) );
  NAND2_X1 U2677 ( .A1(n3946), .A2(n2541), .ZN(n3952) );
  NAND2_X1 U2678 ( .A1(n3954), .A2(n3955), .ZN(n3974) );
  INV_X1 U2679 ( .A(n4575), .ZN(n2322) );
  AOI21_X1 U2680 ( .B1(n4576), .B2(n4577), .A(n4574), .ZN(n2321) );
  OAI21_X1 U2681 ( .B1(n4585), .B2(n4628), .A(n2325), .ZN(n2324) );
  AOI21_X1 U2682 ( .B1(n4579), .B2(ADDR_REG_18__SCAN_IN), .A(n4578), .ZN(n2325) );
  AND2_X1 U2683 ( .A1(n3152), .A2(n3911), .ZN(n4563) );
  NAND2_X1 U2684 ( .A1(n4580), .A2(n2273), .ZN(n2312) );
  XNOR2_X1 U2685 ( .A(n2787), .B(n2678), .ZN(n4004) );
  NAND2_X1 U2686 ( .A1(n4683), .A2(n3098), .ZN(n4276) );
  AND2_X1 U2687 ( .A1(n3129), .A2(n3097), .ZN(n3098) );
  INV_X1 U2688 ( .A(n4300), .ZN(n4601) );
  NOR2_X1 U2689 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2366)
         );
  NOR2_X1 U2690 ( .A1(n2259), .A2(n3708), .ZN(n2333) );
  NOR2_X1 U2691 ( .A1(n2259), .A2(n2335), .ZN(n2334) );
  NAND2_X1 U2692 ( .A1(n2252), .A2(n4410), .ZN(n2922) );
  AND2_X1 U2693 ( .A1(n2252), .A2(n3702), .ZN(n2832) );
  INV_X1 U2694 ( .A(IR_REG_28__SCAN_IN), .ZN(n2384) );
  NAND2_X1 U2695 ( .A1(n4372), .A2(n2252), .ZN(n2973) );
  NAND2_X1 U2696 ( .A1(n2252), .A2(n4389), .ZN(n2952) );
  OAI21_X1 U2697 ( .B1(n3365), .B2(n3342), .A(n3930), .ZN(n3343) );
  AND2_X1 U2698 ( .A1(n4140), .A2(n2718), .ZN(n3862) );
  INV_X1 U2699 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2470) );
  AND2_X1 U2700 ( .A1(n3315), .A2(n3822), .ZN(n3232) );
  INV_X1 U2701 ( .A(n4098), .ZN(n2775) );
  NAND2_X1 U2702 ( .A1(n2279), .A2(n4234), .ZN(n4209) );
  OAI21_X2 U2703 ( .B1(n2747), .B2(n2253), .A(IR_REG_31__SCAN_IN), .ZN(n2382)
         );
  INV_X1 U2704 ( .A(IR_REG_22__SCAN_IN), .ZN(n2684) );
  XNOR2_X1 U2705 ( .A(n2293), .B(IR_REG_20__SCAN_IN), .ZN(n2687) );
  AOI21_X1 U2706 ( .B1(n2680), .B2(n2679), .A(n2690), .ZN(n2293) );
  NAND2_X1 U2707 ( .A1(n2295), .A2(n2342), .ZN(n2524) );
  INV_X1 U2708 ( .A(n2479), .ZN(n2295) );
  INV_X1 U2709 ( .A(IR_REG_5__SCAN_IN), .ZN(n2328) );
  INV_X1 U2710 ( .A(IR_REG_2__SCAN_IN), .ZN(n2360) );
  INV_X1 U2711 ( .A(REG3_REG_14__SCAN_IN), .ZN(n3354) );
  INV_X1 U2712 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3606) );
  INV_X1 U2713 ( .A(n3476), .ZN(n5086) );
  AND2_X1 U2714 ( .A1(n2252), .A2(n4172), .ZN(n2984) );
  XNOR2_X1 U2715 ( .A(n2816), .B(n3069), .ZN(n2326) );
  NAND2_X1 U2716 ( .A1(n2815), .A2(n2814), .ZN(n2816) );
  XNOR2_X1 U2717 ( .A(n2857), .B(n3069), .ZN(n2862) );
  INV_X1 U2718 ( .A(n3317), .ZN(n3222) );
  AND2_X1 U2719 ( .A1(n2594), .A2(REG3_REG_19__SCAN_IN), .ZN(n2605) );
  XNOR2_X1 U2720 ( .A(n2930), .B(n3065), .ZN(n3556) );
  NAND2_X1 U2721 ( .A1(n2252), .A2(n4412), .ZN(n2929) );
  AND2_X1 U2722 ( .A1(n3019), .A2(n3685), .ZN(n3603) );
  OR2_X1 U2723 ( .A1(n2620), .A2(n3690), .ZN(n2631) );
  NOR2_X1 U2724 ( .A1(n2493), .A2(n4965), .ZN(n2505) );
  AND2_X1 U2725 ( .A1(n2977), .A2(n2978), .ZN(n3709) );
  NOR2_X1 U2726 ( .A1(n2577), .A2(n3712), .ZN(n2594) );
  OR2_X1 U2727 ( .A1(n2540), .A2(n2526), .ZN(n2577) );
  NOR2_X1 U2728 ( .A1(n2561), .A2(n3354), .ZN(n2563) );
  INV_X1 U2729 ( .A(n4625), .ZN(n3103) );
  AND3_X1 U2730 ( .A1(n3745), .A2(n3744), .A3(n3743), .ZN(n3987) );
  OR2_X1 U2731 ( .A1(n2651), .A2(n2643), .ZN(n3641) );
  NAND2_X1 U2732 ( .A1(n3362), .A2(n2296), .ZN(n3364) );
  NAND2_X1 U2733 ( .A1(n4492), .A2(REG1_REG_5__SCAN_IN), .ZN(n2296) );
  NAND2_X1 U2734 ( .A1(n3421), .A2(n3422), .ZN(n3425) );
  INV_X1 U2735 ( .A(n2314), .ZN(n3960) );
  AND2_X1 U2736 ( .A1(n2602), .A2(n3127), .ZN(n3150) );
  OR2_X1 U2737 ( .A1(n2669), .A2(n2668), .ZN(n3997) );
  AND2_X1 U2738 ( .A1(n3691), .A2(n4135), .ZN(n2618) );
  AND2_X1 U2739 ( .A1(n3813), .A2(n3812), .ZN(n4146) );
  INV_X1 U2740 ( .A(n4188), .ZN(n4194) );
  INV_X1 U2741 ( .A(n4246), .ZN(n2713) );
  OR2_X1 U2742 ( .A1(n3784), .A2(n3783), .ZN(n4294) );
  INV_X1 U2743 ( .A(n3394), .ZN(n2278) );
  INV_X1 U2744 ( .A(n2868), .ZN(n3395) );
  INV_X1 U2745 ( .A(n3232), .ZN(n3796) );
  CLKBUF_X1 U2746 ( .A(n3261), .Z(n3262) );
  INV_X1 U2747 ( .A(n4587), .ZN(n4599) );
  AND2_X1 U2748 ( .A1(n2602), .A2(DATAI_30_), .ZN(n4309) );
  AND2_X1 U2749 ( .A1(n3777), .A2(n2732), .ZN(n4292) );
  NAND2_X1 U2750 ( .A1(n2602), .A2(DATAI_29_), .ZN(n3992) );
  NOR2_X1 U2751 ( .A1(n4027), .A2(n2788), .ZN(n2807) );
  OR2_X1 U2752 ( .A1(n4043), .A2(n4312), .ZN(n4027) );
  NAND2_X1 U2753 ( .A1(n4063), .A2(n4048), .ZN(n4043) );
  INV_X1 U2754 ( .A(n4411), .ZN(n4612) );
  NAND2_X1 U2755 ( .A1(n2602), .A2(DATAI_23_), .ZN(n4098) );
  NAND2_X1 U2756 ( .A1(n4129), .A2(n4112), .ZN(n4114) );
  INV_X1 U2757 ( .A(n2774), .ZN(n4174) );
  INV_X1 U2758 ( .A(n2279), .ZN(n4249) );
  INV_X1 U2759 ( .A(n2931), .ZN(n4296) );
  OR2_X1 U2760 ( .A1(n3482), .A2(n2915), .ZN(n3531) );
  NOR2_X2 U2761 ( .A1(n3531), .A2(n4410), .ZN(n4297) );
  INV_X1 U2762 ( .A(n2697), .ZN(n3615) );
  INV_X1 U2763 ( .A(n4288), .ZN(n4588) );
  NAND2_X1 U2764 ( .A1(n4479), .A2(n3126), .ZN(n4393) );
  INV_X1 U2765 ( .A(n3234), .ZN(n3079) );
  OR2_X1 U2766 ( .A1(n2692), .A2(n2369), .ZN(n3189) );
  XNOR2_X1 U2767 ( .A(n2746), .B(n2745), .ZN(n2768) );
  INV_X1 U2768 ( .A(IR_REG_24__SCAN_IN), .ZN(n2745) );
  NAND2_X1 U2769 ( .A1(n2744), .A2(IR_REG_31__SCAN_IN), .ZN(n2746) );
  XNOR2_X1 U2770 ( .A(n2755), .B(n2743), .ZN(n3128) );
  CLKBUF_X1 U2771 ( .A(n2479), .Z(n2480) );
  INV_X1 U2772 ( .A(IR_REG_7__SCAN_IN), .ZN(n4964) );
  AND2_X1 U2773 ( .A1(n3638), .A2(n3056), .ZN(n2339) );
  NAND2_X1 U2774 ( .A1(n2337), .A2(n2332), .ZN(n2280) );
  INV_X1 U2775 ( .A(n2335), .ZN(n2332) );
  INV_X1 U2776 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4790) );
  NAND2_X1 U2777 ( .A1(n3501), .A2(n3503), .ZN(n2286) );
  OAI21_X1 U2778 ( .B1(n3501), .B2(n3503), .A(n3502), .ZN(n2287) );
  XNOR2_X1 U2779 ( .A(n2960), .B(n2961), .ZN(n3652) );
  XNOR2_X1 U2780 ( .A(n3029), .B(n3069), .ZN(n3668) );
  NAND2_X1 U2781 ( .A1(n4058), .A2(n2252), .ZN(n3028) );
  AOI21_X1 U2782 ( .B1(n2285), .B2(n2282), .A(n2272), .ZN(n2281) );
  NAND2_X1 U2783 ( .A1(n2285), .A2(n2284), .ZN(n2283) );
  NOR2_X1 U2784 ( .A1(n3502), .A2(n3503), .ZN(n2282) );
  INV_X1 U2785 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3690) );
  NAND2_X1 U2786 ( .A1(n3688), .A2(n3689), .ZN(n2288) );
  NAND2_X1 U2787 ( .A1(n3686), .A2(n3603), .ZN(n3687) );
  INV_X1 U2788 ( .A(n5077), .ZN(n3699) );
  OR2_X1 U2789 ( .A1(n3586), .A2(n2292), .ZN(n2291) );
  INV_X1 U2790 ( .A(n5080), .ZN(n3732) );
  INV_X1 U2791 ( .A(n5081), .ZN(n3731) );
  INV_X1 U2792 ( .A(n4315), .ZN(n4023) );
  NAND2_X1 U2793 ( .A1(n2665), .A2(n2664), .ZN(n4044) );
  NAND2_X1 U2794 ( .A1(n2658), .A2(n2657), .ZN(n4313) );
  OAI211_X1 U2795 ( .C1(n3742), .C2(n4102), .A(n2633), .B(n2632), .ZN(n4335)
         );
  AND3_X1 U2796 ( .A1(n2416), .A2(n2415), .A3(n2414), .ZN(n2419) );
  OR2_X2 U2797 ( .A1(n3118), .A2(n4625), .ZN(n3906) );
  OR2_X1 U2798 ( .A1(n2417), .A2(n2377), .ZN(n2378) );
  AND2_X1 U2799 ( .A1(n3151), .A2(n3150), .ZN(n3911) );
  NAND2_X1 U2800 ( .A1(n2298), .A2(n2297), .ZN(n3921) );
  NAND2_X1 U2801 ( .A1(n2304), .A2(n2265), .ZN(n2297) );
  AND2_X1 U2802 ( .A1(n2299), .A2(n2302), .ZN(n2298) );
  NAND2_X1 U2803 ( .A1(n3140), .A2(n2315), .ZN(n3199) );
  NAND2_X1 U2804 ( .A1(n3196), .A2(n3918), .ZN(n2315) );
  NAND2_X1 U2805 ( .A1(n3209), .A2(n2266), .ZN(n3164) );
  NOR2_X1 U2806 ( .A1(n3149), .A2(n3148), .ZN(n3339) );
  NAND2_X1 U2807 ( .A1(n4558), .A2(n3375), .ZN(n4570) );
  NAND2_X1 U2808 ( .A1(n4553), .A2(n3350), .ZN(n4565) );
  XNOR2_X1 U2809 ( .A(n3420), .B(n3377), .ZN(n3378) );
  NAND2_X1 U2810 ( .A1(n3378), .A2(REG1_REG_14__SCAN_IN), .ZN(n3421) );
  NOR2_X1 U2811 ( .A1(n3416), .A2(n2319), .ZN(n3415) );
  INV_X1 U2812 ( .A(n3352), .ZN(n2318) );
  AND2_X1 U2813 ( .A1(n2319), .A2(n2317), .ZN(n3419) );
  NAND2_X1 U2814 ( .A1(n3952), .A2(n3953), .ZN(n3954) );
  OAI22_X1 U2815 ( .A1(n3998), .A2(n4300), .B1(n3997), .B2(n4276), .ZN(n3999)
         );
  INV_X1 U2816 ( .A(n4312), .ZN(n4028) );
  NAND2_X1 U2817 ( .A1(n2602), .A2(DATAI_26_), .ZN(n4048) );
  NAND2_X1 U2818 ( .A1(n2602), .A2(DATAI_21_), .ZN(n4135) );
  NAND2_X1 U2819 ( .A1(n4617), .A2(n3238), .ZN(n4241) );
  AND2_X1 U2820 ( .A1(n4617), .A2(n3260), .ZN(n4615) );
  INV_X1 U2821 ( .A(n4276), .ZN(n4614) );
  OR2_X1 U2822 ( .A1(n4404), .A2(n4403), .ZN(n4468) );
  NAND2_X1 U2823 ( .A1(n3122), .A2(n3129), .ZN(n4622) );
  INV_X1 U2824 ( .A(n3189), .ZN(n4479) );
  NAND2_X1 U2825 ( .A1(n2257), .A2(IR_REG_31__SCAN_IN), .ZN(n2751) );
  INV_X1 U2826 ( .A(n2753), .ZN(n4480) );
  INV_X1 U2827 ( .A(n2768), .ZN(n4481) );
  NAND2_X1 U2828 ( .A1(n3128), .A2(STATE_REG_SCAN_IN), .ZN(n4625) );
  INV_X1 U2829 ( .A(n3097), .ZN(n4483) );
  INV_X1 U2830 ( .A(n3359), .ZN(n4630) );
  AND2_X1 U2831 ( .A1(n2502), .A2(n2511), .ZN(n4490) );
  AND2_X1 U2832 ( .A1(n2420), .A2(n2412), .ZN(n4494) );
  NAND2_X1 U2833 ( .A1(n2304), .A2(n2307), .ZN(n4496) );
  INV_X2 U2834 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U2835 ( .A(n2324), .ZN(n2323) );
  NAND2_X1 U2836 ( .A1(n2322), .A2(n2321), .ZN(n2320) );
  OAI21_X1 U2837 ( .B1(n2310), .B2(n4500), .A(n3984), .ZN(U3259) );
  XNOR2_X1 U2838 ( .A(n2312), .B(n2311), .ZN(n2310) );
  INV_X1 U2839 ( .A(n3973), .ZN(n2311) );
  AOI22_X1 U2840 ( .A1(n4497), .A2(n4601), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4619), .ZN(n4498) );
  OR2_X1 U2841 ( .A1(n4005), .A2(n4408), .ZN(n2784) );
  NOR2_X1 U2842 ( .A1(n4685), .A2(n3113), .ZN(n3114) );
  OR2_X1 U2843 ( .A1(n4005), .A2(n4472), .ZN(n2779) );
  INV_X2 U2844 ( .A(n2647), .ZN(n2398) );
  OR2_X1 U2845 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2253)
         );
  OR2_X2 U2846 ( .A1(n4027), .A2(n2277), .ZN(n2254) );
  AND2_X1 U2847 ( .A1(n2305), .A2(n3157), .ZN(n2255) );
  INV_X1 U2848 ( .A(IR_REG_1__SCAN_IN), .ZN(n2308) );
  AND2_X1 U2849 ( .A1(n2879), .A2(n3285), .ZN(n2256) );
  NAND2_X1 U2850 ( .A1(n3299), .A2(n3395), .ZN(n3394) );
  AND2_X1 U2851 ( .A1(n2250), .A2(n2327), .ZN(n2433) );
  NAND2_X1 U2852 ( .A1(n2274), .A2(n2275), .ZN(n2258) );
  NAND2_X1 U2853 ( .A1(n2687), .A2(n4483), .ZN(n2813) );
  NAND2_X1 U2854 ( .A1(n3623), .A2(n3006), .ZN(n2259) );
  NOR2_X1 U2855 ( .A1(n3040), .A2(n3039), .ZN(n2261) );
  NAND2_X1 U2856 ( .A1(n2280), .A2(n3708), .ZN(n3622) );
  NAND2_X1 U2857 ( .A1(n2337), .A2(n2971), .ZN(n3707) );
  AND4_X1 U2858 ( .A1(n2679), .A2(n4805), .A3(n2535), .A4(n4806), .ZN(n2262)
         );
  OR2_X1 U2859 ( .A1(n2480), .A2(n2341), .ZN(n2263) );
  NAND2_X1 U2860 ( .A1(n3120), .A2(n4478), .ZN(n2647) );
  NAND2_X1 U2861 ( .A1(n2250), .A2(n2347), .ZN(n2431) );
  OR2_X1 U2862 ( .A1(n2807), .A2(n3992), .ZN(n2264) );
  AND2_X1 U2863 ( .A1(REG1_REG_1__SCAN_IN), .A2(n2307), .ZN(n2265) );
  OR2_X1 U2864 ( .A1(n3163), .A2(n3213), .ZN(n2266) );
  AND2_X1 U2865 ( .A1(n2290), .A2(n3586), .ZN(n2267) );
  OR2_X1 U2866 ( .A1(n2382), .A2(n2800), .ZN(n2269) );
  AND2_X1 U2867 ( .A1(n2907), .A2(n2901), .ZN(n2270) );
  AND2_X1 U2868 ( .A1(n2289), .A2(n2291), .ZN(n3650) );
  INV_X1 U2869 ( .A(n2958), .ZN(n2292) );
  NAND2_X1 U2870 ( .A1(n2287), .A2(n2286), .ZN(n3538) );
  AND2_X1 U2871 ( .A1(n2938), .A2(n2937), .ZN(n3585) );
  INV_X1 U2872 ( .A(IR_REG_20__SCAN_IN), .ZN(n2681) );
  NAND2_X1 U2873 ( .A1(n2902), .A2(n2901), .ZN(n5076) );
  INV_X1 U2874 ( .A(n2776), .ZN(n4097) );
  NOR2_X1 U2875 ( .A1(n4114), .A2(n2775), .ZN(n2776) );
  NAND2_X1 U2876 ( .A1(n3659), .A2(n3658), .ZN(n2271) );
  AND2_X1 U2877 ( .A1(n2435), .A2(n2434), .ZN(n4492) );
  NAND2_X1 U2878 ( .A1(n4210), .A2(n4194), .ZN(n4171) );
  NAND2_X1 U2879 ( .A1(n5089), .A2(n2912), .ZN(n3501) );
  AND2_X1 U2880 ( .A1(n4297), .A2(n4296), .ZN(n4273) );
  INV_X1 U2881 ( .A(IR_REG_27__SCAN_IN), .ZN(n2800) );
  AND2_X1 U2882 ( .A1(n4668), .A2(n3549), .ZN(n3443) );
  AND2_X1 U2883 ( .A1(n3303), .A2(n3298), .ZN(n3299) );
  INV_X1 U2884 ( .A(n2840), .ZN(n2858) );
  NAND2_X1 U2885 ( .A1(n3569), .A2(n2884), .ZN(n3430) );
  AND2_X1 U2886 ( .A1(n2927), .A2(n2926), .ZN(n2272) );
  NAND2_X1 U2887 ( .A1(n2330), .A2(n3285), .ZN(n3567) );
  AND2_X1 U2888 ( .A1(n2835), .A2(n2836), .ZN(n3697) );
  INV_X1 U2889 ( .A(n3680), .ZN(n4151) );
  INV_X1 U2890 ( .A(IR_REG_23__SCAN_IN), .ZN(n2743) );
  OR2_X1 U2891 ( .A1(n4628), .A2(n3972), .ZN(n2273) );
  AND2_X1 U2892 ( .A1(n2602), .A2(DATAI_28_), .ZN(n2788) );
  INV_X1 U2893 ( .A(n2788), .ZN(n4008) );
  BUF_X1 U2894 ( .A(n2371), .Z(n3563) );
  INV_X1 U2895 ( .A(n2376), .ZN(n3120) );
  INV_X1 U2896 ( .A(n2244), .ZN(n2301) );
  NAND2_X1 U2897 ( .A1(n2383), .A2(n2269), .ZN(n2386) );
  NOR2_X2 U2898 ( .A1(n3308), .A2(n2773), .ZN(n3298) );
  NOR2_X2 U2899 ( .A1(n4209), .A2(n4371), .ZN(n4210) );
  NOR2_X2 U2900 ( .A1(n4248), .A2(n4389), .ZN(n2279) );
  AND2_X2 U2901 ( .A1(n4128), .A2(n4135), .ZN(n4129) );
  AND2_X2 U2902 ( .A1(n2774), .A2(n3680), .ZN(n4128) );
  AND2_X2 U2903 ( .A1(n4075), .A2(n4065), .ZN(n4063) );
  NAND4_X1 U2904 ( .A1(n2938), .A2(n2937), .A3(n2958), .A4(n3587), .ZN(n2289)
         );
  NAND3_X1 U2905 ( .A1(n2938), .A2(n2937), .A3(n3587), .ZN(n2290) );
  NAND2_X1 U2906 ( .A1(n3921), .A2(n3920), .ZN(n3919) );
  NAND2_X1 U2907 ( .A1(n2300), .A2(n2305), .ZN(n2304) );
  NAND2_X1 U2908 ( .A1(n2255), .A2(n2300), .ZN(n2299) );
  NAND2_X1 U2909 ( .A1(n2306), .A2(n2244), .ZN(n2305) );
  INV_X1 U2910 ( .A(n3416), .ZN(n2317) );
  OR2_X1 U2911 ( .A1(n3416), .A2(n2318), .ZN(n3353) );
  NAND2_X1 U2912 ( .A1(n3352), .A2(REG2_REG_14__SCAN_IN), .ZN(n2319) );
  NAND3_X1 U2913 ( .A1(n4584), .A2(n2323), .A3(n2320), .ZN(U3258) );
  NAND3_X1 U2914 ( .A1(n2327), .A2(n2250), .A3(n2361), .ZN(n2477) );
  NAND2_X1 U2915 ( .A1(n2864), .A2(n2863), .ZN(n3284) );
  INV_X1 U2916 ( .A(n2863), .ZN(n2331) );
  NAND2_X1 U2917 ( .A1(n2964), .A2(n2963), .ZN(n3657) );
  NAND2_X1 U2918 ( .A1(n2902), .A2(n2270), .ZN(n5089) );
  NAND2_X1 U2919 ( .A1(n3639), .A2(n3637), .ZN(n2340) );
  NAND2_X1 U2920 ( .A1(n2340), .A2(n3638), .ZN(n3717) );
  NAND2_X1 U2921 ( .A1(n2340), .A2(n2339), .ZN(n3061) );
  NAND2_X1 U2922 ( .A1(n2249), .A2(n2366), .ZN(n2747) );
  NAND2_X1 U2923 ( .A1(n3243), .A2(n3702), .ZN(n3820) );
  CLKBUF_X1 U2924 ( .A(n3797), .Z(n4593) );
  NAND2_X1 U2926 ( .A1(n2389), .A2(REG2_REG_2__SCAN_IN), .ZN(n2399) );
  OR2_X1 U2927 ( .A1(n2834), .A2(n2833), .ZN(n2835) );
  AND2_X1 U2928 ( .A1(n2631), .A2(n3606), .ZN(n2346) );
  OR4_X1 U2929 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n2348) );
  NOR2_X1 U2930 ( .A1(n2552), .A2(n2551), .ZN(n2350) );
  AND2_X1 U2931 ( .A1(n3085), .A2(n3084), .ZN(n2351) );
  AND2_X1 U2932 ( .A1(n2548), .A2(n4806), .ZN(n2352) );
  NOR2_X1 U2933 ( .A1(n4180), .A2(n4186), .ZN(n2353) );
  OR2_X1 U2934 ( .A1(n4325), .A2(n4028), .ZN(n2355) );
  NAND2_X1 U2935 ( .A1(n4702), .A2(n4399), .ZN(n4408) );
  INV_X1 U2936 ( .A(n2786), .ZN(n2678) );
  INV_X1 U2937 ( .A(D_REG_0__SCAN_IN), .ZN(n2766) );
  NOR2_X1 U2938 ( .A1(n3602), .A2(n3020), .ZN(n2357) );
  NOR2_X1 U2939 ( .A1(n2605), .A2(n2595), .ZN(n2358) );
  NAND2_X1 U2940 ( .A1(n2602), .A2(DATAI_24_), .ZN(n4080) );
  INV_X1 U2941 ( .A(n4080), .ZN(n4334) );
  AND2_X1 U2942 ( .A1(n3109), .A2(n3108), .ZN(n2359) );
  NAND2_X1 U2943 ( .A1(n2602), .A2(DATAI_22_), .ZN(n4112) );
  INV_X1 U2944 ( .A(IR_REG_13__SCAN_IN), .ZN(n2364) );
  INV_X1 U2945 ( .A(IR_REG_18__SCAN_IN), .ZN(n4805) );
  NAND2_X1 U2946 ( .A1(n2842), .A2(n2252), .ZN(n2844) );
  INV_X1 U2947 ( .A(n4112), .ZN(n2627) );
  INV_X1 U2948 ( .A(n3568), .ZN(n2879) );
  INV_X1 U2949 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2484) );
  NAND2_X1 U2950 ( .A1(n4352), .A2(n2627), .ZN(n2628) );
  AND2_X1 U2951 ( .A1(n3088), .A2(n3699), .ZN(n3084) );
  INV_X1 U2952 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2526) );
  OR2_X1 U2953 ( .A1(n2471), .A2(n2470), .ZN(n2485) );
  INV_X1 U2954 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2515) );
  AND2_X1 U2955 ( .A1(n2563), .A2(REG3_REG_15__SCAN_IN), .ZN(n2552) );
  OR2_X1 U2956 ( .A1(n4485), .A2(n3890), .ZN(n3101) );
  OR2_X1 U2957 ( .A1(n2485), .A2(n2484), .ZN(n2493) );
  NOR2_X1 U2958 ( .A1(n3363), .A2(n3337), .ZN(n3338) );
  AND2_X1 U2959 ( .A1(n3975), .A2(REG2_REG_18__SCAN_IN), .ZN(n3976) );
  AND2_X1 U2960 ( .A1(n2670), .A2(n3997), .ZN(n4006) );
  NOR2_X1 U2961 ( .A1(n4058), .A2(n4334), .ZN(n2640) );
  AOI21_X1 U2962 ( .B1(n4126), .B2(n2619), .A(n2618), .ZN(n4118) );
  OR2_X1 U2963 ( .A1(n4179), .A2(n4204), .ZN(n4221) );
  NAND2_X1 U2964 ( .A1(n4023), .A2(n2788), .ZN(n2789) );
  INV_X1 U2965 ( .A(n4215), .ZN(n4371) );
  INV_X1 U2966 ( .A(n4393), .ZN(n4589) );
  AND2_X1 U2967 ( .A1(n3189), .A2(n3126), .ZN(n4411) );
  OR2_X1 U2968 ( .A1(n2611), .A2(n4790), .ZN(n2620) );
  AND3_X1 U2969 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2439) );
  OR2_X1 U2970 ( .A1(n2516), .A2(n2515), .ZN(n2561) );
  INV_X1 U2971 ( .A(n2915), .ZN(n3532) );
  NAND2_X1 U2972 ( .A1(n3105), .A2(n4479), .ZN(n5081) );
  AND2_X1 U2973 ( .A1(n2642), .A2(REG3_REG_25__SCAN_IN), .ZN(n2651) );
  AND2_X1 U2974 ( .A1(n2636), .A2(REG3_REG_24__SCAN_IN), .ZN(n2642) );
  INV_X1 U2975 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4939) );
  INV_X1 U2976 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4965) );
  INV_X1 U2977 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3712) );
  INV_X1 U2978 ( .A(n4044), .ZN(n4325) );
  INV_X1 U2979 ( .A(n3995), .ZN(n4256) );
  AND2_X1 U2980 ( .A1(n2602), .A2(DATAI_27_), .ZN(n4312) );
  AND2_X1 U2981 ( .A1(n3092), .A2(n3129), .ZN(n3235) );
  OR2_X1 U2982 ( .A1(n3129), .A2(n3891), .ZN(n3151) );
  NOR2_X1 U2983 ( .A1(n3104), .A2(n3893), .ZN(n3105) );
  AND3_X1 U2984 ( .A1(n2799), .A2(n2798), .A3(n2797), .ZN(n3775) );
  AND2_X1 U2985 ( .A1(n3911), .A2(n3908), .ZN(n4581) );
  INV_X1 U2986 ( .A(n3814), .ZN(n4186) );
  INV_X1 U2987 ( .A(n4241), .ZN(n4302) );
  INV_X1 U2988 ( .A(n4292), .ZN(n4609) );
  INV_X1 U2989 ( .A(n4408), .ZN(n2808) );
  NAND2_X1 U2990 ( .A1(n2771), .A2(n2770), .ZN(n3234) );
  NAND2_X1 U2991 ( .A1(n2602), .A2(DATAI_25_), .ZN(n4065) );
  NAND2_X1 U2992 ( .A1(n4594), .A2(n4643), .ZN(n4665) );
  AND2_X1 U2993 ( .A1(n3308), .A2(n3272), .ZN(n4689) );
  AND2_X1 U2994 ( .A1(n3118), .A2(n3103), .ZN(n3129) );
  XNOR2_X1 U2995 ( .A(n2751), .B(IR_REG_26__SCAN_IN), .ZN(n2754) );
  AND2_X1 U2996 ( .A1(n2525), .A2(n2568), .ZN(n3359) );
  AND2_X1 U2997 ( .A1(n3130), .A2(n3151), .ZN(n4579) );
  NAND2_X1 U2998 ( .A1(n3105), .A2(n3189), .ZN(n5080) );
  OR2_X1 U2999 ( .A1(n3104), .A2(n3083), .ZN(n5077) );
  NAND4_X1 U3000 ( .A1(n2600), .A2(n2599), .A3(n2598), .A4(n2597), .ZN(n4189)
         );
  INV_X1 U3001 ( .A(n4563), .ZN(n4574) );
  NAND2_X1 U3002 ( .A1(n3911), .A2(n3189), .ZN(n4585) );
  OR2_X1 U3003 ( .A1(n4197), .A2(n4678), .ZN(n4300) );
  NAND2_X2 U3004 ( .A1(n3237), .A2(n4276), .ZN(n4617) );
  INV_X1 U3005 ( .A(n4702), .ZN(n4700) );
  OR2_X1 U3006 ( .A1(n2781), .A2(n3079), .ZN(n4684) );
  INV_X1 U3007 ( .A(n4622), .ZN(n4624) );
  INV_X1 U3008 ( .A(n3890), .ZN(n4482) );
  AND2_X1 U3009 ( .A1(n2560), .A2(n2559), .ZN(n4488) );
  AND2_X1 U3010 ( .A1(n2466), .A2(n2457), .ZN(n4491) );
  INV_X1 U3011 ( .A(REG0_REG_28__SCAN_IN), .ZN(n2772) );
  NOR2_X2 U3012 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2402)
         );
  INV_X1 U3013 ( .A(IR_REG_26__SCAN_IN), .ZN(n2367) );
  NAND2_X1 U3014 ( .A1(n2688), .A2(n2384), .ZN(n2372) );
  INV_X1 U3015 ( .A(n2372), .ZN(n2369) );
  INV_X1 U3016 ( .A(IR_REG_29__SCAN_IN), .ZN(n2368) );
  NAND2_X1 U3017 ( .A1(n2369), .A2(n2368), .ZN(n2371) );
  XNOR2_X2 U3018 ( .A(n2370), .B(IR_REG_30__SCAN_IN), .ZN(n4478) );
  NAND2_X1 U3019 ( .A1(n2372), .A2(IR_REG_31__SCAN_IN), .ZN(n2373) );
  NAND2_X1 U3020 ( .A1(n2248), .A2(REG1_REG_0__SCAN_IN), .ZN(n2381) );
  NAND2_X1 U3021 ( .A1(n2398), .A2(REG3_REG_0__SCAN_IN), .ZN(n2380) );
  NOR2_X2 U3023 ( .A1(n3120), .A2(n4478), .ZN(n2394) );
  NAND2_X1 U3024 ( .A1(n3741), .A2(REG0_REG_0__SCAN_IN), .ZN(n2379) );
  NAND2_X1 U3025 ( .A1(n4478), .A2(n2376), .ZN(n2417) );
  INV_X1 U3026 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2377) );
  NAND2_X1 U3027 ( .A1(n2382), .A2(n2384), .ZN(n2383) );
  NAND2_X1 U3028 ( .A1(n2384), .A2(IR_REG_27__SCAN_IN), .ZN(n2385) );
  NAND2_X2 U3029 ( .A1(n2386), .A2(n2385), .ZN(n2436) );
  MUX2_X1 U3030 ( .A(n2244), .B(DATAI_0_), .S(n2436), .Z(n3181) );
  AND2_X1 U3031 ( .A1(n2821), .A2(n3181), .ZN(n4592) );
  NAND2_X1 U3032 ( .A1(n2394), .A2(REG0_REG_1__SCAN_IN), .ZN(n2388) );
  NAND2_X1 U3033 ( .A1(n2251), .A2(REG1_REG_1__SCAN_IN), .ZN(n2387) );
  AND2_X1 U3034 ( .A1(n2388), .A2(n2387), .ZN(n2392) );
  NAND2_X1 U3035 ( .A1(n2398), .A2(REG3_REG_1__SCAN_IN), .ZN(n2391) );
  NAND2_X1 U3036 ( .A1(n2389), .A2(REG2_REG_1__SCAN_IN), .ZN(n2390) );
  MUX2_X1 U3037 ( .A(n4496), .B(DATAI_1_), .S(n2436), .Z(n4587) );
  NAND2_X1 U3038 ( .A1(n2812), .A2(n4599), .ZN(n3818) );
  NAND2_X1 U3039 ( .A1(n4592), .A2(n3797), .ZN(n4591) );
  NAND2_X1 U3040 ( .A1(n2812), .A2(n4587), .ZN(n2393) );
  NAND2_X1 U3041 ( .A1(n4591), .A2(n2393), .ZN(n3257) );
  INV_X1 U3042 ( .A(n3257), .ZN(n2404) );
  NAND2_X1 U3043 ( .A1(n2394), .A2(REG0_REG_2__SCAN_IN), .ZN(n2397) );
  NAND2_X1 U3044 ( .A1(n2251), .A2(REG1_REG_2__SCAN_IN), .ZN(n2396) );
  AND2_X1 U3045 ( .A1(n2397), .A2(n2396), .ZN(n2401) );
  NAND2_X1 U3046 ( .A1(n2398), .A2(REG3_REG_2__SCAN_IN), .ZN(n2400) );
  NAND3_X2 U3047 ( .A1(n2401), .A2(n2400), .A3(n2399), .ZN(n3907) );
  OR2_X1 U3048 ( .A1(n2402), .A2(n2690), .ZN(n2403) );
  MUX2_X1 U3050 ( .A(n4495), .B(DATAI_2_), .S(n2436), .Z(n3702) );
  INV_X1 U3051 ( .A(n3702), .ZN(n3266) );
  NAND2_X1 U3052 ( .A1(n3907), .A2(n3266), .ZN(n3823) );
  NAND2_X1 U3053 ( .A1(n3820), .A2(n3823), .ZN(n3799) );
  NAND2_X1 U3054 ( .A1(n2404), .A2(n3799), .ZN(n3229) );
  INV_X1 U3055 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3618) );
  NAND2_X1 U3056 ( .A1(n2398), .A2(n3618), .ZN(n2408) );
  NAND2_X1 U3057 ( .A1(n3741), .A2(REG0_REG_3__SCAN_IN), .ZN(n2407) );
  NAND2_X1 U3058 ( .A1(n3740), .A2(REG1_REG_3__SCAN_IN), .ZN(n2406) );
  INV_X1 U3059 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3242) );
  OR2_X1 U3060 ( .A1(n2417), .A2(n3242), .ZN(n2405) );
  NAND2_X1 U3061 ( .A1(n2409), .A2(IR_REG_31__SCAN_IN), .ZN(n2411) );
  NAND2_X1 U3062 ( .A1(n2411), .A2(n2410), .ZN(n2420) );
  OR2_X1 U3063 ( .A1(n2411), .A2(n2410), .ZN(n2412) );
  MUX2_X1 U3064 ( .A(n4494), .B(DATAI_3_), .S(n2436), .Z(n2697) );
  NAND2_X1 U3065 ( .A1(n3905), .A2(n2697), .ZN(n3311) );
  INV_X1 U3066 ( .A(n3311), .ZN(n2423) );
  NOR2_X1 U3067 ( .A1(n3907), .A2(n3702), .ZN(n3230) );
  NOR2_X1 U3068 ( .A1(n3905), .A2(n2697), .ZN(n3312) );
  AOI21_X1 U3069 ( .B1(n3230), .B2(n3311), .A(n3312), .ZN(n2422) );
  NAND2_X1 U3070 ( .A1(n3741), .A2(REG0_REG_4__SCAN_IN), .ZN(n2416) );
  INV_X1 U3071 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2413) );
  XNOR2_X1 U3072 ( .A(n2413), .B(REG3_REG_3__SCAN_IN), .ZN(n3324) );
  NAND2_X1 U3073 ( .A1(n2398), .A2(n3324), .ZN(n2415) );
  NAND2_X1 U3074 ( .A1(n2248), .A2(REG1_REG_4__SCAN_IN), .ZN(n2414) );
  INV_X1 U3075 ( .A(REG2_REG_4__SCAN_IN), .ZN(n3145) );
  OR2_X1 U3076 ( .A1(n2417), .A2(n3145), .ZN(n2418) );
  INV_X1 U3077 ( .A(n2842), .ZN(n3330) );
  NAND2_X1 U3078 ( .A1(n2420), .A2(IR_REG_31__SCAN_IN), .ZN(n2421) );
  XNOR2_X1 U3079 ( .A(n2421), .B(IR_REG_4__SCAN_IN), .ZN(n4493) );
  MUX2_X1 U3080 ( .A(n4493), .B(DATAI_4_), .S(n2436), .Z(n3317) );
  NAND2_X1 U3081 ( .A1(n3330), .A2(n3317), .ZN(n2699) );
  NAND2_X1 U3082 ( .A1(n2842), .A2(n3222), .ZN(n3828) );
  NAND2_X1 U3083 ( .A1(n2699), .A2(n3828), .ZN(n3793) );
  OAI211_X1 U3084 ( .C1(n3229), .C2(n2423), .A(n2422), .B(n3793), .ZN(n2425)
         );
  NAND2_X1 U3085 ( .A1(n2842), .A2(n3317), .ZN(n2424) );
  NAND2_X1 U3086 ( .A1(n2425), .A2(n2424), .ZN(n3295) );
  NAND2_X1 U3088 ( .A1(n3740), .A2(REG1_REG_5__SCAN_IN), .ZN(n2430) );
  AOI21_X1 U3089 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        REG3_REG_5__SCAN_IN), .ZN(n2426) );
  NOR2_X1 U3090 ( .A1(n2426), .A2(n2439), .ZN(n3300) );
  NAND2_X1 U3091 ( .A1(n2734), .A2(n3300), .ZN(n2429) );
  NAND2_X1 U3092 ( .A1(n2795), .A2(REG0_REG_5__SCAN_IN), .ZN(n2428) );
  INV_X1 U3093 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3337) );
  OR2_X1 U3094 ( .A1(n3742), .A2(n3337), .ZN(n2427) );
  NAND2_X1 U3095 ( .A1(n2431), .A2(IR_REG_31__SCAN_IN), .ZN(n2432) );
  MUX2_X1 U3096 ( .A(IR_REG_31__SCAN_IN), .B(n2432), .S(IR_REG_5__SCAN_IN), 
        .Z(n2435) );
  INV_X1 U3097 ( .A(n2433), .ZN(n2434) );
  CLKBUF_X3 U3098 ( .A(n2436), .Z(n2602) );
  MUX2_X1 U3099 ( .A(n4492), .B(DATAI_5_), .S(n2602), .Z(n3328) );
  AND2_X1 U3100 ( .A1(n3390), .A2(n3328), .ZN(n2438) );
  INV_X1 U3101 ( .A(n3390), .ZN(n2701) );
  NAND2_X1 U3102 ( .A1(n2701), .A2(n3303), .ZN(n2437) );
  OAI21_X1 U3103 ( .B1(n3295), .B2(n2438), .A(n2437), .ZN(n3388) );
  NAND2_X1 U3104 ( .A1(n3740), .A2(REG1_REG_6__SCAN_IN), .ZN(n2445) );
  NAND2_X1 U3105 ( .A1(n2795), .A2(REG0_REG_6__SCAN_IN), .ZN(n2444) );
  NAND2_X1 U3106 ( .A1(n2439), .A2(REG3_REG_6__SCAN_IN), .ZN(n2448) );
  OAI21_X1 U3107 ( .B1(n2439), .B2(REG3_REG_6__SCAN_IN), .A(n2448), .ZN(n2440)
         );
  INV_X1 U3108 ( .A(n2440), .ZN(n3396) );
  NAND2_X1 U3109 ( .A1(n2734), .A2(n3396), .ZN(n2443) );
  INV_X1 U3110 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2441) );
  OR2_X1 U3111 ( .A1(n3742), .A2(n2441), .ZN(n2442) );
  NAND4_X1 U3112 ( .A1(n2445), .A2(n2444), .A3(n2443), .A4(n2442), .ZN(n3571)
         );
  OR2_X1 U3113 ( .A1(n2433), .A2(n2690), .ZN(n2446) );
  XNOR2_X1 U3114 ( .A(n2446), .B(IR_REG_6__SCAN_IN), .ZN(n4635) );
  MUX2_X1 U3115 ( .A(n4635), .B(DATAI_6_), .S(n2602), .Z(n2868) );
  NOR2_X1 U3116 ( .A1(n3571), .A2(n2868), .ZN(n2447) );
  INV_X1 U3117 ( .A(n3571), .ZN(n3405) );
  OAI22_X2 U3118 ( .A1(n3388), .A2(n2447), .B1(n3405), .B2(n3395), .ZN(n3411)
         );
  NAND2_X1 U3119 ( .A1(n3740), .A2(REG1_REG_7__SCAN_IN), .ZN(n2453) );
  NAND2_X1 U3120 ( .A1(n2795), .A2(REG0_REG_7__SCAN_IN), .ZN(n2452) );
  NOR2_X1 U3121 ( .A1(n2448), .A2(n4939), .ZN(n2460) );
  AND2_X1 U3122 ( .A1(n2448), .A2(n4939), .ZN(n2449) );
  NOR2_X1 U3123 ( .A1(n2460), .A2(n2449), .ZN(n3574) );
  NAND2_X1 U3124 ( .A1(n2734), .A2(n3574), .ZN(n2451) );
  INV_X1 U3125 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3342) );
  OR2_X1 U3126 ( .A1(n3742), .A2(n3342), .ZN(n2450) );
  NAND4_X1 U3127 ( .A1(n2453), .A2(n2452), .A3(n2451), .A4(n2450), .ZN(n3904)
         );
  INV_X1 U3128 ( .A(n3904), .ZN(n3459) );
  INV_X1 U3129 ( .A(IR_REG_6__SCAN_IN), .ZN(n2454) );
  NAND2_X1 U3130 ( .A1(n2433), .A2(n2454), .ZN(n2455) );
  NAND2_X1 U3131 ( .A1(n2455), .A2(IR_REG_31__SCAN_IN), .ZN(n2456) );
  NAND2_X1 U3132 ( .A1(n2456), .A2(n4964), .ZN(n2466) );
  OR2_X1 U3133 ( .A1(n2456), .A2(n4964), .ZN(n2457) );
  MUX2_X1 U3134 ( .A(n4491), .B(DATAI_7_), .S(n2602), .Z(n3406) );
  NAND2_X1 U3135 ( .A1(n3459), .A2(n3406), .ZN(n2703) );
  INV_X1 U3136 ( .A(n3406), .ZN(n3572) );
  NAND2_X1 U3137 ( .A1(n3904), .A2(n3572), .ZN(n3839) );
  NAND2_X1 U3138 ( .A1(n2703), .A2(n3839), .ZN(n3794) );
  NAND2_X1 U3139 ( .A1(n3411), .A2(n3794), .ZN(n2459) );
  NAND2_X1 U3140 ( .A1(n3904), .A2(n3406), .ZN(n2458) );
  NAND2_X1 U3141 ( .A1(n2459), .A2(n2458), .ZN(n3454) );
  NAND2_X1 U3142 ( .A1(n3740), .A2(REG1_REG_8__SCAN_IN), .ZN(n2465) );
  NAND2_X1 U3143 ( .A1(n2460), .A2(REG3_REG_8__SCAN_IN), .ZN(n2471) );
  OR2_X1 U3144 ( .A1(n2460), .A2(REG3_REG_8__SCAN_IN), .ZN(n2461) );
  AND2_X1 U3145 ( .A1(n2471), .A2(n2461), .ZN(n3467) );
  NAND2_X1 U3146 ( .A1(n2734), .A2(n3467), .ZN(n2464) );
  NAND2_X1 U3147 ( .A1(n2795), .A2(REG0_REG_8__SCAN_IN), .ZN(n2463) );
  INV_X1 U31480 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3469) );
  OR2_X1 U31490 ( .A1(n3742), .A2(n3469), .ZN(n2462) );
  NAND4_X1 U3150 ( .A1(n2465), .A2(n2464), .A3(n2463), .A4(n2462), .ZN(n3903)
         );
  NAND2_X1 U3151 ( .A1(n2466), .A2(IR_REG_31__SCAN_IN), .ZN(n2467) );
  XNOR2_X1 U3152 ( .A(n2467), .B(IR_REG_8__SCAN_IN), .ZN(n3367) );
  MUX2_X1 U3153 ( .A(n3367), .B(DATAI_8_), .S(n2602), .Z(n3457) );
  AND2_X1 U3154 ( .A1(n3903), .A2(n3457), .ZN(n2469) );
  INV_X1 U3155 ( .A(n3903), .ZN(n3447) );
  INV_X1 U3156 ( .A(n3457), .ZN(n3465) );
  NAND2_X1 U3157 ( .A1(n3447), .A2(n3465), .ZN(n2468) );
  OAI21_X1 U3158 ( .B1(n3454), .B2(n2469), .A(n2468), .ZN(n3442) );
  NAND2_X1 U3159 ( .A1(n2471), .A2(n2470), .ZN(n2472) );
  NAND2_X1 U3160 ( .A1(n2485), .A2(n2472), .ZN(n3445) );
  INV_X1 U3161 ( .A(n3445), .ZN(n3551) );
  NAND2_X1 U3162 ( .A1(n2734), .A2(n3551), .ZN(n2476) );
  NAND2_X1 U3163 ( .A1(n2795), .A2(REG0_REG_9__SCAN_IN), .ZN(n2475) );
  NAND2_X1 U3164 ( .A1(n3740), .A2(REG1_REG_9__SCAN_IN), .ZN(n2474) );
  INV_X1 U3165 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3336) );
  OR2_X1 U3166 ( .A1(n3742), .A2(n3336), .ZN(n2473) );
  NAND4_X1 U3167 ( .A1(n2476), .A2(n2475), .A3(n2474), .A4(n2473), .ZN(n3902)
         );
  NAND2_X1 U3168 ( .A1(n2477), .A2(IR_REG_31__SCAN_IN), .ZN(n2478) );
  MUX2_X1 U3169 ( .A(IR_REG_31__SCAN_IN), .B(n2478), .S(IR_REG_9__SCAN_IN), 
        .Z(n2481) );
  AND2_X1 U3170 ( .A1(n2481), .A2(n2480), .ZN(n4519) );
  MUX2_X1 U3171 ( .A(n4519), .B(DATAI_9_), .S(n2602), .Z(n3490) );
  NOR2_X1 U3172 ( .A1(n3902), .A2(n3490), .ZN(n2483) );
  NAND2_X1 U3173 ( .A1(n3902), .A2(n3490), .ZN(n2482) );
  NAND2_X1 U3174 ( .A1(n2248), .A2(REG1_REG_10__SCAN_IN), .ZN(n2490) );
  NAND2_X1 U3175 ( .A1(n2485), .A2(n2484), .ZN(n2486) );
  AND2_X1 U3176 ( .A1(n2493), .A2(n2486), .ZN(n5083) );
  NAND2_X1 U3177 ( .A1(n2734), .A2(n5083), .ZN(n2489) );
  NAND2_X1 U3178 ( .A1(n2795), .A2(REG0_REG_10__SCAN_IN), .ZN(n2488) );
  INV_X1 U3179 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3484) );
  OR2_X1 U3180 ( .A1(n3742), .A2(n3484), .ZN(n2487) );
  NAND4_X1 U3181 ( .A1(n2490), .A2(n2489), .A3(n2488), .A4(n2487), .ZN(n3901)
         );
  NAND2_X1 U3182 ( .A1(n2480), .A2(IR_REG_31__SCAN_IN), .ZN(n2491) );
  XNOR2_X1 U3183 ( .A(n2491), .B(IR_REG_10__SCAN_IN), .ZN(n4632) );
  MUX2_X1 U3184 ( .A(n4632), .B(DATAI_10_), .S(n2602), .Z(n3476) );
  AND2_X1 U3185 ( .A1(n3901), .A2(n3476), .ZN(n2492) );
  NAND2_X1 U3186 ( .A1(n2248), .A2(REG1_REG_11__SCAN_IN), .ZN(n2498) );
  AND2_X1 U3187 ( .A1(n2493), .A2(n4965), .ZN(n2494) );
  NOR2_X1 U3188 ( .A1(n2505), .A2(n2494), .ZN(n3533) );
  NAND2_X1 U3189 ( .A1(n2734), .A2(n3533), .ZN(n2497) );
  NAND2_X1 U3190 ( .A1(n2795), .A2(REG0_REG_11__SCAN_IN), .ZN(n2496) );
  INV_X1 U3191 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3335) );
  OR2_X1 U3192 ( .A1(n3742), .A2(n3335), .ZN(n2495) );
  NAND4_X1 U3193 ( .A1(n2498), .A2(n2497), .A3(n2496), .A4(n2495), .ZN(n4413)
         );
  INV_X1 U3194 ( .A(n4413), .ZN(n5079) );
  OR2_X1 U3195 ( .A1(n2499), .A2(n2690), .ZN(n2501) );
  INV_X1 U3196 ( .A(IR_REG_11__SCAN_IN), .ZN(n2500) );
  OR2_X1 U3197 ( .A1(n2501), .A2(n2500), .ZN(n2502) );
  NAND2_X1 U3198 ( .A1(n2501), .A2(n2500), .ZN(n2511) );
  MUX2_X1 U3199 ( .A(n4490), .B(DATAI_11_), .S(n2602), .Z(n2915) );
  NAND2_X1 U3200 ( .A1(n5079), .A2(n2915), .ZN(n3510) );
  NAND2_X1 U3201 ( .A1(n4413), .A2(n3532), .ZN(n3512) );
  NAND2_X1 U3202 ( .A1(n3510), .A2(n3512), .ZN(n3795) );
  NAND2_X1 U3203 ( .A1(n3525), .A2(n3795), .ZN(n2504) );
  NAND2_X1 U3204 ( .A1(n5079), .A2(n3532), .ZN(n2503) );
  NAND2_X1 U3205 ( .A1(n2504), .A2(n2503), .ZN(n3515) );
  NAND2_X1 U3206 ( .A1(n2248), .A2(REG1_REG_12__SCAN_IN), .ZN(n2510) );
  NAND2_X1 U3207 ( .A1(n2795), .A2(REG0_REG_12__SCAN_IN), .ZN(n2509) );
  OR2_X1 U3208 ( .A1(n2505), .A2(REG3_REG_12__SCAN_IN), .ZN(n2506) );
  NAND2_X1 U3209 ( .A1(n2505), .A2(REG3_REG_12__SCAN_IN), .ZN(n2516) );
  AND2_X1 U32100 ( .A1(n2506), .A2(n2516), .ZN(n3544) );
  NAND2_X1 U32110 ( .A1(n2734), .A2(n3544), .ZN(n2508) );
  INV_X1 U32120 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3518) );
  OR2_X1 U32130 ( .A1(n3742), .A2(n3518), .ZN(n2507) );
  NAND4_X1 U32140 ( .A1(n2510), .A2(n2509), .A3(n2508), .A4(n2507), .ZN(n4290)
         );
  NAND2_X1 U32150 ( .A1(n2511), .A2(IR_REG_31__SCAN_IN), .ZN(n2512) );
  XNOR2_X1 U32160 ( .A(n2512), .B(IR_REG_12__SCAN_IN), .ZN(n3373) );
  MUX2_X1 U32170 ( .A(n3373), .B(DATAI_12_), .S(n2602), .Z(n4410) );
  NOR2_X1 U32180 ( .A1(n4290), .A2(n4410), .ZN(n2514) );
  NAND2_X1 U32190 ( .A1(n4290), .A2(n4410), .ZN(n2513) );
  OAI21_X2 U32200 ( .B1(n3515), .B2(n2514), .A(n2513), .ZN(n4179) );
  INV_X1 U32210 ( .A(n4179), .ZN(n2591) );
  NAND2_X1 U32220 ( .A1(n3740), .A2(REG1_REG_13__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U32230 ( .A1(n2516), .A2(n2515), .ZN(n2517) );
  AND2_X1 U32240 ( .A1(n2561), .A2(n2517), .ZN(n4298) );
  NAND2_X1 U32250 ( .A1(n2734), .A2(n4298), .ZN(n2521) );
  NAND2_X1 U32260 ( .A1(n2795), .A2(REG0_REG_13__SCAN_IN), .ZN(n2520) );
  INV_X1 U32270 ( .A(REG2_REG_13__SCAN_IN), .ZN(n2518) );
  OR2_X1 U32280 ( .A1(n3742), .A2(n2518), .ZN(n2519) );
  NAND4_X1 U32290 ( .A1(n2522), .A2(n2521), .A3(n2520), .A4(n2519), .ZN(n4412)
         );
  NAND2_X1 U32300 ( .A1(n2524), .A2(IR_REG_31__SCAN_IN), .ZN(n2523) );
  MUX2_X1 U32310 ( .A(IR_REG_31__SCAN_IN), .B(n2523), .S(IR_REG_13__SCAN_IN), 
        .Z(n2525) );
  MUX2_X1 U32320 ( .A(n3359), .B(DATAI_13_), .S(n2602), .Z(n2931) );
  AND2_X1 U32330 ( .A1(n4412), .A2(n2931), .ZN(n4204) );
  NAND2_X1 U32340 ( .A1(n3740), .A2(REG1_REG_17__SCAN_IN), .ZN(n2532) );
  NAND2_X1 U32350 ( .A1(n2795), .A2(REG0_REG_17__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U32360 ( .A1(n2552), .A2(REG3_REG_16__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U32370 ( .A1(n2540), .A2(n2526), .ZN(n2527) );
  AND2_X1 U32380 ( .A1(n2577), .A2(n2527), .ZN(n4212) );
  NAND2_X1 U32390 ( .A1(n2734), .A2(n4212), .ZN(n2530) );
  INV_X1 U32400 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2528) );
  OR2_X1 U32410 ( .A1(n3742), .A2(n2528), .ZN(n2529) );
  NAND4_X1 U32420 ( .A1(n2532), .A2(n2531), .A3(n2530), .A4(n2529), .ZN(n4380)
         );
  INV_X1 U32430 ( .A(n4380), .ZN(n4191) );
  NOR2_X1 U32440 ( .A1(n2536), .A2(n2690), .ZN(n2533) );
  MUX2_X1 U32450 ( .A(n2690), .B(n2533), .S(IR_REG_17__SCAN_IN), .Z(n2534) );
  INV_X1 U32460 ( .A(n2534), .ZN(n2537) );
  NAND2_X1 U32470 ( .A1(n2536), .A2(n2535), .ZN(n2601) );
  NAND2_X1 U32480 ( .A1(n2537), .A2(n2601), .ZN(n3968) );
  INV_X1 U32490 ( .A(DATAI_17_), .ZN(n2538) );
  MUX2_X1 U32500 ( .A(n3968), .B(n2538), .S(n2602), .Z(n4215) );
  NAND2_X1 U32510 ( .A1(n4191), .A2(n4215), .ZN(n2586) );
  INV_X1 U32520 ( .A(n2586), .ZN(n2575) );
  NAND2_X1 U32530 ( .A1(n3740), .A2(REG1_REG_16__SCAN_IN), .ZN(n2545) );
  OR2_X1 U32540 ( .A1(n2552), .A2(REG3_REG_16__SCAN_IN), .ZN(n2539) );
  AND2_X1 U32550 ( .A1(n2540), .A2(n2539), .ZN(n4231) );
  NAND2_X1 U32560 ( .A1(n2734), .A2(n4231), .ZN(n2544) );
  NAND2_X1 U32570 ( .A1(n2795), .A2(REG0_REG_16__SCAN_IN), .ZN(n2543) );
  INV_X1 U32580 ( .A(REG2_REG_16__SCAN_IN), .ZN(n2541) );
  OR2_X1 U32590 ( .A1(n3742), .A2(n2541), .ZN(n2542) );
  NAND4_X1 U32600 ( .A1(n2545), .A2(n2544), .A3(n2543), .A4(n2542), .ZN(n4390)
         );
  INV_X1 U32610 ( .A(n2546), .ZN(n2547) );
  AND2_X1 U32620 ( .A1(n2547), .A2(IR_REG_31__SCAN_IN), .ZN(n2558) );
  INV_X1 U32630 ( .A(n2558), .ZN(n2549) );
  NAND2_X1 U32640 ( .A1(n2549), .A2(n2548), .ZN(n2559) );
  NAND2_X1 U32650 ( .A1(n2559), .A2(IR_REG_31__SCAN_IN), .ZN(n2550) );
  XNOR2_X1 U32660 ( .A(n2550), .B(IR_REG_16__SCAN_IN), .ZN(n4487) );
  MUX2_X1 U32670 ( .A(n4487), .B(DATAI_16_), .S(n2602), .Z(n4379) );
  NAND2_X1 U32680 ( .A1(n4390), .A2(n4379), .ZN(n2574) );
  INV_X1 U32690 ( .A(n4390), .ZN(n4375) );
  NAND2_X1 U32700 ( .A1(n4375), .A2(n4379), .ZN(n3749) );
  INV_X1 U32710 ( .A(n4379), .ZN(n4234) );
  NAND2_X1 U32720 ( .A1(n4390), .A2(n4234), .ZN(n4201) );
  NAND2_X1 U32730 ( .A1(n3749), .A2(n4201), .ZN(n4228) );
  NAND2_X1 U32740 ( .A1(n3740), .A2(REG1_REG_15__SCAN_IN), .ZN(n2557) );
  NAND2_X1 U32750 ( .A1(n2795), .A2(REG0_REG_15__SCAN_IN), .ZN(n2556) );
  NOR2_X1 U32760 ( .A1(n2563), .A2(REG3_REG_15__SCAN_IN), .ZN(n2551) );
  NAND2_X1 U32770 ( .A1(n2734), .A2(n2350), .ZN(n2555) );
  INV_X1 U32780 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2553) );
  OR2_X1 U32790 ( .A1(n3742), .A2(n2553), .ZN(n2554) );
  NAND2_X1 U32800 ( .A1(n2558), .A2(IR_REG_15__SCAN_IN), .ZN(n2560) );
  MUX2_X1 U32810 ( .A(n4488), .B(DATAI_15_), .S(n2602), .Z(n4389) );
  NAND2_X1 U32820 ( .A1(n4266), .A2(n4389), .ZN(n2572) );
  INV_X1 U32830 ( .A(n2572), .ZN(n2571) );
  NAND2_X1 U32840 ( .A1(n3740), .A2(REG1_REG_14__SCAN_IN), .ZN(n2567) );
  AND2_X1 U32850 ( .A1(n2561), .A2(n3354), .ZN(n2562) );
  NOR2_X1 U32860 ( .A1(n2563), .A2(n2562), .ZN(n4275) );
  NAND2_X1 U32870 ( .A1(n2734), .A2(n4275), .ZN(n2566) );
  NAND2_X1 U32880 ( .A1(n2795), .A2(REG0_REG_14__SCAN_IN), .ZN(n2565) );
  INV_X1 U32890 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4278) );
  OR2_X1 U32900 ( .A1(n3742), .A2(n4278), .ZN(n2564) );
  NAND2_X1 U32910 ( .A1(n2568), .A2(IR_REG_31__SCAN_IN), .ZN(n2569) );
  XNOR2_X1 U32920 ( .A(n2569), .B(IR_REG_14__SCAN_IN), .ZN(n4489) );
  MUX2_X1 U32930 ( .A(n4489), .B(DATAI_14_), .S(n2602), .Z(n2942) );
  NAND2_X1 U32940 ( .A1(n4394), .A2(n4274), .ZN(n4245) );
  OR2_X1 U32950 ( .A1(n2571), .A2(n2570), .ZN(n4223) );
  INV_X1 U32960 ( .A(n2585), .ZN(n2573) );
  NAND2_X1 U32970 ( .A1(n4394), .A2(n2942), .ZN(n3751) );
  NAND2_X1 U32980 ( .A1(n4251), .A2(n4274), .ZN(n3747) );
  NAND2_X1 U32990 ( .A1(n3751), .A2(n3747), .ZN(n4263) );
  AND2_X1 U33000 ( .A1(n4263), .A2(n2572), .ZN(n4222) );
  OR2_X1 U33010 ( .A1(n4204), .A2(n2588), .ZN(n2576) );
  AND2_X1 U33020 ( .A1(n4380), .A2(n4371), .ZN(n2590) );
  NAND2_X1 U33030 ( .A1(n2248), .A2(REG1_REG_18__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U33040 ( .A1(n2795), .A2(REG0_REG_18__SCAN_IN), .ZN(n2582) );
  AND2_X1 U33050 ( .A1(n2577), .A2(n3712), .ZN(n2578) );
  NOR2_X1 U33060 ( .A1(n2594), .A2(n2578), .ZN(n4195) );
  NAND2_X1 U33070 ( .A1(n2734), .A2(n4195), .ZN(n2581) );
  INV_X1 U33080 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2579) );
  OR2_X1 U33090 ( .A1(n3742), .A2(n2579), .ZN(n2580) );
  NAND4_X1 U33100 ( .A1(n2583), .A2(n2582), .A3(n2581), .A4(n2580), .ZN(n4372)
         );
  INV_X1 U33110 ( .A(n4372), .ZN(n2592) );
  NAND2_X1 U33120 ( .A1(n2601), .A2(IR_REG_31__SCAN_IN), .ZN(n2584) );
  XNOR2_X1 U33130 ( .A(n2584), .B(IR_REG_18__SCAN_IN), .ZN(n3975) );
  MUX2_X1 U33140 ( .A(n3975), .B(DATAI_18_), .S(n2602), .Z(n4188) );
  NAND2_X1 U33150 ( .A1(n2592), .A2(n4188), .ZN(n4162) );
  NAND2_X1 U33160 ( .A1(n4372), .A2(n4194), .ZN(n4163) );
  NAND2_X1 U33170 ( .A1(n4162), .A2(n4163), .ZN(n3814) );
  INV_X1 U33180 ( .A(n4412), .ZN(n3591) );
  NAND2_X1 U33190 ( .A1(n3591), .A2(n4296), .ZN(n4220) );
  AND2_X1 U33200 ( .A1(n4220), .A2(n2585), .ZN(n4205) );
  AND2_X1 U33210 ( .A1(n4205), .A2(n2586), .ZN(n2587) );
  NAND2_X1 U33220 ( .A1(n2592), .A2(n4194), .ZN(n2593) );
  NAND2_X1 U33230 ( .A1(n4183), .A2(n2593), .ZN(n4159) );
  NAND2_X1 U33240 ( .A1(n2248), .A2(REG1_REG_19__SCAN_IN), .ZN(n2600) );
  NOR2_X1 U33250 ( .A1(n2594), .A2(REG3_REG_19__SCAN_IN), .ZN(n2595) );
  NAND2_X1 U33260 ( .A1(n2734), .A2(n2358), .ZN(n2599) );
  NAND2_X1 U33270 ( .A1(n2795), .A2(REG0_REG_19__SCAN_IN), .ZN(n2598) );
  INV_X1 U33280 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2596) );
  OR2_X1 U33290 ( .A1(n3742), .A2(n2596), .ZN(n2597) );
  MUX2_X1 U33300 ( .A(n4485), .B(DATAI_19_), .S(n2602), .Z(n4172) );
  NAND2_X1 U33310 ( .A1(n4189), .A2(n4172), .ZN(n2604) );
  NOR2_X1 U33320 ( .A1(n4189), .A2(n4172), .ZN(n2603) );
  AOI21_X1 U33330 ( .B1(n4159), .B2(n2604), .A(n2603), .ZN(n4147) );
  NAND2_X1 U33340 ( .A1(n2248), .A2(REG1_REG_20__SCAN_IN), .ZN(n2610) );
  NAND2_X1 U33350 ( .A1(n2605), .A2(REG3_REG_20__SCAN_IN), .ZN(n2611) );
  OR2_X1 U33360 ( .A1(n2605), .A2(REG3_REG_20__SCAN_IN), .ZN(n2606) );
  AND2_X1 U33370 ( .A1(n2611), .A2(n2606), .ZN(n4152) );
  NAND2_X1 U33380 ( .A1(n2734), .A2(n4152), .ZN(n2609) );
  NAND2_X1 U33390 ( .A1(n2795), .A2(REG0_REG_20__SCAN_IN), .ZN(n2608) );
  INV_X1 U33400 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4154) );
  OR2_X1 U33410 ( .A1(n3742), .A2(n4154), .ZN(n2607) );
  NAND4_X1 U33420 ( .A1(n2610), .A2(n2609), .A3(n2608), .A4(n2607), .ZN(n4131)
         );
  NAND2_X1 U33430 ( .A1(n2602), .A2(DATAI_20_), .ZN(n3680) );
  AND2_X1 U33440 ( .A1(n4131), .A2(n4151), .ZN(n3811) );
  INV_X1 U33450 ( .A(n4131), .ZN(n4355) );
  NAND2_X1 U33460 ( .A1(n4355), .A2(n3680), .ZN(n3812) );
  OAI21_X1 U33470 ( .B1(n4147), .B2(n3811), .A(n3812), .ZN(n4126) );
  NAND2_X1 U33480 ( .A1(n2248), .A2(REG1_REG_21__SCAN_IN), .ZN(n2617) );
  NAND2_X1 U33490 ( .A1(n2611), .A2(n4790), .ZN(n2612) );
  AND2_X1 U33500 ( .A1(n2620), .A2(n2612), .ZN(n4132) );
  NAND2_X1 U33510 ( .A1(n2734), .A2(n4132), .ZN(n2616) );
  NAND2_X1 U33520 ( .A1(n2795), .A2(REG0_REG_21__SCAN_IN), .ZN(n2615) );
  INV_X1 U3353 ( .A(REG2_REG_21__SCAN_IN), .ZN(n2613) );
  OR2_X1 U33540 ( .A1(n3742), .A2(n2613), .ZN(n2614) );
  NAND4_X1 U3355 ( .A1(n2617), .A2(n2616), .A3(n2615), .A4(n2614), .ZN(n4143)
         );
  INV_X1 U3356 ( .A(n4135), .ZN(n4351) );
  NAND2_X1 U3357 ( .A1(n4143), .A2(n4351), .ZN(n2619) );
  INV_X1 U3358 ( .A(n4143), .ZN(n3691) );
  NAND2_X1 U3359 ( .A1(n2248), .A2(REG1_REG_22__SCAN_IN), .ZN(n2626) );
  NAND2_X1 U3360 ( .A1(n2795), .A2(REG0_REG_22__SCAN_IN), .ZN(n2625) );
  NAND2_X1 U3361 ( .A1(n2620), .A2(n3690), .ZN(n2621) );
  AND2_X1 U3362 ( .A1(n2631), .A2(n2621), .ZN(n4115) );
  NAND2_X1 U3363 ( .A1(n2734), .A2(n4115), .ZN(n2624) );
  INV_X1 U3364 ( .A(REG2_REG_22__SCAN_IN), .ZN(n2622) );
  OR2_X1 U3365 ( .A1(n3742), .A2(n2622), .ZN(n2623) );
  NAND4_X1 U3366 ( .A1(n2626), .A2(n2625), .A3(n2624), .A4(n2623), .ZN(n4352)
         );
  INV_X1 U3367 ( .A(n4352), .ZN(n3632) );
  NAND2_X1 U3368 ( .A1(n3632), .A2(n2627), .ZN(n4088) );
  NAND2_X1 U3369 ( .A1(n4352), .A2(n4112), .ZN(n2722) );
  NAND2_X1 U3370 ( .A1(n4088), .A2(n2722), .ZN(n4117) );
  NAND2_X1 U3371 ( .A1(n4118), .A2(n4117), .ZN(n4119) );
  NAND2_X1 U3372 ( .A1(n4119), .A2(n2628), .ZN(n4085) );
  INV_X1 U3373 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4102) );
  NAND2_X1 U3374 ( .A1(n2248), .A2(REG1_REG_23__SCAN_IN), .ZN(n2630) );
  NAND2_X1 U3375 ( .A1(n2795), .A2(REG0_REG_23__SCAN_IN), .ZN(n2629) );
  AND2_X1 U3376 ( .A1(n2630), .A2(n2629), .ZN(n2633) );
  NOR2_X1 U3377 ( .A1(n2636), .A2(n2346), .ZN(n4100) );
  NAND2_X1 U3378 ( .A1(n4100), .A2(n2734), .ZN(n2632) );
  INV_X1 U3379 ( .A(n4335), .ZN(n4108) );
  NAND2_X1 U3380 ( .A1(n4108), .A2(n4098), .ZN(n2635) );
  NOR2_X1 U3381 ( .A1(n2636), .A2(REG3_REG_24__SCAN_IN), .ZN(n2637) );
  OR2_X1 U3382 ( .A1(n2642), .A2(n2637), .ZN(n3669) );
  AOI22_X1 U3383 ( .A1(n2389), .A2(REG2_REG_24__SCAN_IN), .B1(n2248), .B2(
        REG1_REG_24__SCAN_IN), .ZN(n2639) );
  NAND2_X1 U3384 ( .A1(n2795), .A2(REG0_REG_24__SCAN_IN), .ZN(n2638) );
  OAI211_X1 U3385 ( .C1(n3669), .C2(n2647), .A(n2639), .B(n2638), .ZN(n4058)
         );
  NAND2_X1 U3386 ( .A1(n4058), .A2(n4334), .ZN(n2641) );
  INV_X1 U3387 ( .A(n4058), .ZN(n4093) );
  NOR2_X1 U3388 ( .A1(n2642), .A2(REG3_REG_25__SCAN_IN), .ZN(n2643) );
  AOI22_X1 U3389 ( .A1(n2248), .A2(REG1_REG_25__SCAN_IN), .B1(n2795), .B2(
        REG0_REG_25__SCAN_IN), .ZN(n2646) );
  INV_X1 U3390 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2644) );
  OR2_X1 U3391 ( .A1(n3742), .A2(n2644), .ZN(n2645) );
  OAI211_X1 U3392 ( .C1(n2647), .C2(n3641), .A(n2646), .B(n2645), .ZN(n4322)
         );
  INV_X1 U3393 ( .A(n4322), .ZN(n4338) );
  NAND2_X1 U3394 ( .A1(n4338), .A2(n4065), .ZN(n2650) );
  INV_X1 U3395 ( .A(n4065), .ZN(n2648) );
  OR2_X1 U3396 ( .A1(n2651), .A2(REG3_REG_26__SCAN_IN), .ZN(n2652) );
  NAND2_X1 U3397 ( .A1(n4045), .A2(n2734), .ZN(n2658) );
  INV_X1 U3398 ( .A(REG2_REG_26__SCAN_IN), .ZN(n2655) );
  NAND2_X1 U3399 ( .A1(n2248), .A2(REG1_REG_26__SCAN_IN), .ZN(n2654) );
  NAND2_X1 U3400 ( .A1(n2795), .A2(REG0_REG_26__SCAN_IN), .ZN(n2653) );
  OAI211_X1 U3401 ( .C1(n2655), .C2(n3742), .A(n2654), .B(n2653), .ZN(n2656)
         );
  INV_X1 U3402 ( .A(n2656), .ZN(n2657) );
  INV_X1 U3403 ( .A(n4048), .ZN(n4321) );
  NAND2_X1 U3404 ( .A1(n4313), .A2(n4321), .ZN(n2659) );
  INV_X1 U3405 ( .A(n4313), .ZN(n3643) );
  XNOR2_X1 U3406 ( .A(n2669), .B(REG3_REG_27__SCAN_IN), .ZN(n4024) );
  NAND2_X1 U3407 ( .A1(n4024), .A2(n2734), .ZN(n2665) );
  INV_X1 U3408 ( .A(REG2_REG_27__SCAN_IN), .ZN(n2662) );
  NAND2_X1 U3409 ( .A1(n2248), .A2(REG1_REG_27__SCAN_IN), .ZN(n2661) );
  NAND2_X1 U3410 ( .A1(n2795), .A2(REG0_REG_27__SCAN_IN), .ZN(n2660) );
  OAI211_X1 U3411 ( .C1(n2662), .C2(n3742), .A(n2661), .B(n2660), .ZN(n2663)
         );
  INV_X1 U3412 ( .A(n2663), .ZN(n2664) );
  OR2_X1 U3413 ( .A1(n4044), .A2(n4312), .ZN(n2666) );
  NAND2_X1 U3414 ( .A1(n4019), .A2(n2666), .ZN(n2667) );
  NAND2_X1 U3415 ( .A1(n2667), .A2(n2355), .ZN(n2787) );
  INV_X1 U3416 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3580) );
  INV_X1 U3417 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3100) );
  OAI21_X1 U3418 ( .B1(n2669), .B2(n3580), .A(n3100), .ZN(n2670) );
  NAND2_X1 U3419 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_28__SCAN_IN), .ZN(
        n2668) );
  NAND2_X1 U3420 ( .A1(n4006), .A2(n2734), .ZN(n2676) );
  INV_X1 U3421 ( .A(REG2_REG_28__SCAN_IN), .ZN(n2673) );
  NAND2_X1 U3422 ( .A1(n3741), .A2(REG0_REG_28__SCAN_IN), .ZN(n2672) );
  NAND2_X1 U3423 ( .A1(n2248), .A2(REG1_REG_28__SCAN_IN), .ZN(n2671) );
  OAI211_X1 U3424 ( .C1(n3742), .C2(n2673), .A(n2672), .B(n2671), .ZN(n2674)
         );
  INV_X1 U3425 ( .A(n2674), .ZN(n2675) );
  AND2_X1 U3426 ( .A1(n4315), .A2(n2788), .ZN(n3762) );
  INV_X1 U3427 ( .A(n3762), .ZN(n2677) );
  NAND2_X1 U3428 ( .A1(n4023), .A2(n4008), .ZN(n3767) );
  NAND2_X1 U3429 ( .A1(n2677), .A2(n3767), .ZN(n2786) );
  NAND2_X1 U3430 ( .A1(n2263), .A2(IR_REG_31__SCAN_IN), .ZN(n2682) );
  MUX2_X1 U3431 ( .A(IR_REG_31__SCAN_IN), .B(n2682), .S(IR_REG_21__SCAN_IN), 
        .Z(n2683) );
  NAND2_X1 U3432 ( .A1(n2683), .A2(n2258), .ZN(n3097) );
  NAND2_X1 U3433 ( .A1(n2258), .A2(IR_REG_31__SCAN_IN), .ZN(n2685) );
  XNOR2_X1 U3434 ( .A(n2813), .B(n4482), .ZN(n2686) );
  AND2_X1 U3435 ( .A1(n3883), .A2(n4485), .ZN(n4608) );
  AND2_X1 U3436 ( .A1(n4608), .A2(n3890), .ZN(n4683) );
  INV_X1 U3437 ( .A(n4683), .ZN(n4643) );
  NOR2_X1 U3438 ( .A1(n2688), .A2(n2690), .ZN(n2689) );
  MUX2_X1 U3439 ( .A(n2690), .B(n2689), .S(IR_REG_28__SCAN_IN), .Z(n2692) );
  INV_X1 U3440 ( .A(n2821), .ZN(n2693) );
  NAND2_X1 U3441 ( .A1(n2693), .A2(n3181), .ZN(n3798) );
  INV_X1 U3442 ( .A(n3798), .ZN(n4586) );
  INV_X1 U3443 ( .A(n3797), .ZN(n2694) );
  NAND2_X1 U3444 ( .A1(n4586), .A2(n2694), .ZN(n3261) );
  NAND2_X1 U3445 ( .A1(n3261), .A2(n2695), .ZN(n2696) );
  INV_X1 U3446 ( .A(n3799), .ZN(n3256) );
  NAND2_X1 U3447 ( .A1(n2696), .A2(n3256), .ZN(n3240) );
  NAND2_X1 U3448 ( .A1(n3240), .A2(n3820), .ZN(n2698) );
  INV_X1 U3449 ( .A(n3905), .ZN(n3319) );
  NAND2_X1 U3450 ( .A1(n3319), .A2(n2697), .ZN(n3315) );
  NAND2_X1 U3451 ( .A1(n3905), .A2(n3615), .ZN(n3822) );
  AND2_X1 U3452 ( .A1(n3315), .A2(n2699), .ZN(n3825) );
  NAND2_X1 U3453 ( .A1(n3239), .A2(n3825), .ZN(n2700) );
  AND2_X1 U3454 ( .A1(n3390), .A2(n3303), .ZN(n3294) );
  NAND2_X1 U3455 ( .A1(n2701), .A2(n3328), .ZN(n3834) );
  OAI21_X2 U3456 ( .B1(n3296), .B2(n3294), .A(n3834), .ZN(n3387) );
  NAND2_X1 U3457 ( .A1(n3571), .A2(n3395), .ZN(n3833) );
  NAND2_X1 U34580 ( .A1(n3387), .A2(n3833), .ZN(n2702) );
  NAND2_X1 U34590 ( .A1(n3405), .A2(n2868), .ZN(n3830) );
  NAND2_X1 U3460 ( .A1(n2702), .A2(n3830), .ZN(n3401) );
  INV_X1 U3461 ( .A(n2703), .ZN(n2704) );
  NAND2_X1 U3462 ( .A1(n3447), .A2(n3457), .ZN(n3844) );
  AND2_X1 U3463 ( .A1(n3903), .A2(n3465), .ZN(n3840) );
  INV_X1 U3464 ( .A(n3490), .ZN(n3549) );
  NAND2_X1 U3465 ( .A1(n3902), .A2(n3549), .ZN(n3846) );
  NAND2_X1 U3466 ( .A1(n3440), .A2(n3846), .ZN(n2705) );
  INV_X1 U34670 ( .A(n3902), .ZN(n5082) );
  NAND2_X1 U3468 ( .A1(n5082), .A2(n3490), .ZN(n3845) );
  NAND2_X1 U34690 ( .A1(n3901), .A2(n5086), .ZN(n3851) );
  NAND2_X1 U3470 ( .A1(n3475), .A2(n3851), .ZN(n2706) );
  INV_X1 U34710 ( .A(n3901), .ZN(n3446) );
  NAND2_X1 U3472 ( .A1(n3446), .A2(n3476), .ZN(n3850) );
  NAND2_X1 U34730 ( .A1(n2706), .A2(n3850), .ZN(n3509) );
  INV_X1 U3474 ( .A(n4410), .ZN(n3541) );
  NAND2_X1 U34750 ( .A1(n4290), .A2(n3541), .ZN(n4283) );
  NAND2_X1 U3476 ( .A1(n4412), .A2(n4296), .ZN(n3782) );
  NAND2_X1 U34770 ( .A1(n4283), .A2(n3782), .ZN(n2708) );
  INV_X1 U3478 ( .A(n3512), .ZN(n2707) );
  NOR2_X1 U34790 ( .A1(n2708), .A2(n2707), .ZN(n3852) );
  NAND2_X1 U3480 ( .A1(n3509), .A2(n3852), .ZN(n2711) );
  INV_X1 U34810 ( .A(n4290), .ZN(n3526) );
  NAND2_X1 U3482 ( .A1(n3526), .A2(n4410), .ZN(n4285) );
  NAND2_X1 U34830 ( .A1(n3510), .A2(n4285), .ZN(n2710) );
  INV_X1 U3484 ( .A(n2708), .ZN(n2709) );
  NOR2_X1 U34850 ( .A1(n4412), .A2(n4296), .ZN(n3783) );
  AOI21_X1 U3486 ( .B1(n2710), .B2(n2709), .A(n3783), .ZN(n3858) );
  NAND2_X1 U34870 ( .A1(n2711), .A2(n3858), .ZN(n3746) );
  INV_X1 U3488 ( .A(n4263), .ZN(n4265) );
  NAND2_X1 U34890 ( .A1(n3746), .A2(n4265), .ZN(n2712) );
  NAND2_X1 U3490 ( .A1(n2712), .A2(n3751), .ZN(n4242) );
  INV_X1 U34910 ( .A(n4242), .ZN(n2714) );
  INV_X1 U3492 ( .A(n4266), .ZN(n4382) );
  NAND2_X1 U34930 ( .A1(n4382), .A2(n4389), .ZN(n3750) );
  INV_X1 U3494 ( .A(n4389), .ZN(n4257) );
  NAND2_X1 U34950 ( .A1(n4266), .A2(n4257), .ZN(n3748) );
  NAND2_X1 U3496 ( .A1(n3750), .A2(n3748), .ZN(n4246) );
  INV_X1 U34970 ( .A(n4228), .ZN(n4236) );
  NAND2_X1 U3498 ( .A1(n4380), .A2(n4215), .ZN(n3861) );
  AND2_X1 U34990 ( .A1(n4201), .A2(n3861), .ZN(n3753) );
  NAND2_X1 U3500 ( .A1(n4191), .A2(n4371), .ZN(n4160) );
  NAND2_X1 U35010 ( .A1(n4162), .A2(n4160), .ZN(n2717) );
  INV_X1 U3502 ( .A(n4172), .ZN(n4167) );
  NAND2_X1 U35030 ( .A1(n4189), .A2(n4167), .ZN(n2715) );
  AND2_X1 U3504 ( .A1(n4163), .A2(n2715), .ZN(n2719) );
  NOR2_X1 U35050 ( .A1(n4189), .A2(n4167), .ZN(n2716) );
  AOI21_X1 U35060 ( .B1(n2717), .B2(n2719), .A(n2716), .ZN(n4140) );
  NAND2_X1 U35070 ( .A1(n4355), .A2(n4151), .ZN(n2718) );
  NAND2_X1 U35080 ( .A1(n4161), .A2(n3862), .ZN(n2721) );
  INV_X1 U35090 ( .A(n2719), .ZN(n4141) );
  AND2_X1 U35100 ( .A1(n4131), .A2(n3680), .ZN(n2720) );
  AOI21_X1 U35110 ( .B1(n3862), .B2(n4141), .A(n2720), .ZN(n3866) );
  NAND2_X1 U35120 ( .A1(n2721), .A2(n3866), .ZN(n4124) );
  NAND2_X1 U35130 ( .A1(n3691), .A2(n4351), .ZN(n4086) );
  AND2_X1 U35140 ( .A1(n4088), .A2(n4086), .ZN(n3869) );
  NAND2_X1 U35150 ( .A1(n4124), .A2(n3869), .ZN(n2725) );
  NAND2_X1 U35160 ( .A1(n4335), .A2(n4098), .ZN(n3809) );
  AND2_X1 U35170 ( .A1(n3809), .A2(n2722), .ZN(n3874) );
  AND2_X1 U35180 ( .A1(n4143), .A2(n4135), .ZN(n4087) );
  NAND2_X1 U35190 ( .A1(n4088), .A2(n4087), .ZN(n2723) );
  NAND2_X1 U35200 ( .A1(n3874), .A2(n2723), .ZN(n3760) );
  INV_X1 U35210 ( .A(n3760), .ZN(n2724) );
  NAND2_X1 U35220 ( .A1(n2725), .A2(n2724), .ZN(n2726) );
  OR2_X1 U35230 ( .A1(n4335), .A2(n4098), .ZN(n3810) );
  NAND2_X1 U35240 ( .A1(n2726), .A2(n3810), .ZN(n4071) );
  INV_X1 U35250 ( .A(n4071), .ZN(n2727) );
  OR2_X1 U35260 ( .A1(n4058), .A2(n4080), .ZN(n3808) );
  INV_X1 U35270 ( .A(n3808), .ZN(n3758) );
  NAND2_X1 U35280 ( .A1(n2727), .A2(n3808), .ZN(n4034) );
  OR2_X1 U35290 ( .A1(n4322), .A2(n4065), .ZN(n4036) );
  OAI21_X1 U35300 ( .B1(n4313), .B2(n4048), .A(n4036), .ZN(n3872) );
  NAND2_X1 U35310 ( .A1(n4322), .A2(n4065), .ZN(n3780) );
  NAND2_X1 U35320 ( .A1(n4058), .A2(n4080), .ZN(n4054) );
  AND2_X1 U35330 ( .A1(n3780), .A2(n4054), .ZN(n4035) );
  OR2_X1 U35340 ( .A1(n3872), .A2(n4035), .ZN(n2728) );
  NAND2_X1 U35350 ( .A1(n4313), .A2(n4048), .ZN(n3768) );
  NAND2_X1 U35360 ( .A1(n2728), .A2(n3768), .ZN(n3877) );
  INV_X1 U35370 ( .A(n3877), .ZN(n2729) );
  XNOR2_X1 U35380 ( .A(n4044), .B(n4312), .ZN(n4018) );
  INV_X1 U35390 ( .A(n4018), .ZN(n4020) );
  NOR2_X1 U35400 ( .A1(n4044), .A2(n4028), .ZN(n3761) );
  INV_X1 U35410 ( .A(n3761), .ZN(n2731) );
  XNOR2_X1 U35420 ( .A(n2793), .B(n2678), .ZN(n2733) );
  INV_X1 U35430 ( .A(n3883), .ZN(n4484) );
  NAND2_X1 U35440 ( .A1(n4484), .A2(n4483), .ZN(n3777) );
  NAND2_X1 U35450 ( .A1(n4485), .A2(n4482), .ZN(n2732) );
  NAND2_X1 U35460 ( .A1(n2733), .A2(n4609), .ZN(n4017) );
  INV_X1 U35470 ( .A(n3997), .ZN(n2735) );
  NAND2_X1 U35480 ( .A1(n2735), .A2(n2734), .ZN(n2740) );
  INV_X1 U35490 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3993) );
  NAND2_X1 U35500 ( .A1(n3741), .A2(REG0_REG_29__SCAN_IN), .ZN(n2737) );
  NAND2_X1 U35510 ( .A1(n2248), .A2(REG1_REG_29__SCAN_IN), .ZN(n2736) );
  OAI211_X1 U35520 ( .C1(n3742), .C2(n3993), .A(n2737), .B(n2736), .ZN(n2738)
         );
  INV_X1 U35530 ( .A(n2738), .ZN(n2739) );
  NAND2_X1 U35540 ( .A1(n2740), .A2(n2739), .ZN(n3900) );
  AOI22_X1 U35550 ( .A1(n3900), .A2(n4411), .B1(n4588), .B2(n2788), .ZN(n2741)
         );
  OAI211_X1 U35560 ( .C1(n4325), .C2(n4393), .A(n4017), .B(n2741), .ZN(n2742)
         );
  AOI21_X1 U35570 ( .B1(n4004), .B2(n4665), .A(n2742), .ZN(n2782) );
  NAND2_X1 U35580 ( .A1(n2755), .A2(n2743), .ZN(n2744) );
  NAND2_X1 U35590 ( .A1(n2747), .A2(IR_REG_31__SCAN_IN), .ZN(n2748) );
  MUX2_X1 U35600 ( .A(IR_REG_31__SCAN_IN), .B(n2748), .S(IR_REG_25__SCAN_IN), 
        .Z(n2749) );
  NAND2_X1 U35610 ( .A1(n2749), .A2(n2257), .ZN(n2753) );
  NAND2_X1 U35620 ( .A1(n2768), .A2(n2753), .ZN(n2750) );
  MUX2_X1 U35630 ( .A(n2768), .B(n2750), .S(B_REG_SCAN_IN), .Z(n2752) );
  OAI22_X1 U35640 ( .A1(n3122), .A2(D_REG_1__SCAN_IN), .B1(n4480), .B2(n2754), 
        .ZN(n3078) );
  NAND2_X1 U35650 ( .A1(n3883), .A2(n3981), .ZN(n3080) );
  NAND2_X1 U35660 ( .A1(n3080), .A2(n3126), .ZN(n3092) );
  INV_X1 U35670 ( .A(n3122), .ZN(n2767) );
  NOR4_X1 U35680 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2764) );
  NOR4_X1 U35690 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2763) );
  INV_X1 U35700 ( .A(D_REG_13__SCAN_IN), .ZN(n4620) );
  INV_X1 U35710 ( .A(D_REG_7__SCAN_IN), .ZN(n4621) );
  INV_X1 U35720 ( .A(D_REG_2__SCAN_IN), .ZN(n4623) );
  INV_X1 U35730 ( .A(D_REG_12__SCAN_IN), .ZN(n4822) );
  NAND4_X1 U35740 ( .A1(n4620), .A2(n4621), .A3(n4623), .A4(n4822), .ZN(n2761)
         );
  NOR4_X1 U35750 ( .A1(D_REG_3__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2759) );
  NOR4_X1 U35760 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2758) );
  NOR4_X1 U35770 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2757) );
  NOR4_X1 U35780 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2756) );
  NAND4_X1 U35790 ( .A1(n2759), .A2(n2758), .A3(n2757), .A4(n2756), .ZN(n2760)
         );
  NOR4_X1 U35800 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(n2761), 
        .A4(n2760), .ZN(n2762) );
  NAND3_X1 U35810 ( .A1(n2764), .A2(n2763), .A3(n2762), .ZN(n2765) );
  NAND2_X1 U3582 ( .A1(n2767), .A2(n2765), .ZN(n3233) );
  NAND3_X1 U3583 ( .A1(n4288), .A2(n4605), .A3(n4485), .ZN(n3091) );
  NAND2_X1 U3584 ( .A1(n2767), .A2(n2766), .ZN(n2771) );
  INV_X1 U3585 ( .A(n2754), .ZN(n2769) );
  NAND2_X1 U3586 ( .A1(n2769), .A2(n2768), .ZN(n2770) );
  MUX2_X1 U3587 ( .A(n2772), .B(n2782), .S(n4685), .Z(n2780) );
  NAND2_X1 U3588 ( .A1(n4607), .A2(n4599), .ZN(n4598) );
  NAND2_X1 U3589 ( .A1(n3222), .A2(n3615), .ZN(n2773) );
  NOR2_X4 U3590 ( .A1(n3464), .A2(n3457), .ZN(n4668) );
  NAND2_X1 U3591 ( .A1(n3443), .A2(n5086), .ZN(n3482) );
  NAND2_X1 U3592 ( .A1(n4273), .A2(n4274), .ZN(n4248) );
  NOR2_X2 U3593 ( .A1(n4171), .A2(n4172), .ZN(n2774) );
  INV_X1 U3594 ( .A(n4027), .ZN(n2778) );
  INV_X1 U3595 ( .A(n2807), .ZN(n2777) );
  OAI21_X1 U3596 ( .B1(n2778), .B2(n4008), .A(n2777), .ZN(n4005) );
  NAND2_X1 U3597 ( .A1(n4685), .A2(n4399), .ZN(n4472) );
  NAND2_X1 U3598 ( .A1(n2780), .A2(n2779), .ZN(U3514) );
  INV_X1 U3599 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2783) );
  NOR2_X4 U3600 ( .A1(n2781), .A2(n3234), .ZN(n4702) );
  MUX2_X1 U3601 ( .A(n2783), .B(n2782), .S(n4702), .Z(n2785) );
  NAND2_X1 U3602 ( .A1(n2785), .A2(n2784), .ZN(U3546) );
  NAND2_X1 U3603 ( .A1(n2787), .A2(n2786), .ZN(n2790) );
  NAND2_X1 U3604 ( .A1(n2790), .A2(n2789), .ZN(n2792) );
  XNOR2_X1 U3605 ( .A(n3900), .B(n3992), .ZN(n3806) );
  INV_X1 U3606 ( .A(n3806), .ZN(n2791) );
  NAND2_X1 U3607 ( .A1(n3991), .A2(n4665), .ZN(n2803) );
  AOI21_X1 U3608 ( .B1(n2793), .B2(n3767), .A(n3762), .ZN(n2794) );
  XOR2_X1 U3609 ( .A(n3806), .B(n2794), .Z(n2801) );
  NAND2_X1 U3610 ( .A1(n2248), .A2(REG1_REG_30__SCAN_IN), .ZN(n2799) );
  NAND2_X1 U3611 ( .A1(n2795), .A2(REG0_REG_30__SCAN_IN), .ZN(n2798) );
  INV_X1 U3612 ( .A(REG2_REG_30__SCAN_IN), .ZN(n2796) );
  OR2_X1 U3613 ( .A1(n3742), .A2(n2796), .ZN(n2797) );
  XNOR2_X1 U3614 ( .A(n2382), .B(n2800), .ZN(n3908) );
  INV_X1 U3615 ( .A(B_REG_SCAN_IN), .ZN(n3889) );
  OAI21_X1 U3616 ( .B1(n3908), .B2(n3889), .A(n4411), .ZN(n3986) );
  OAI22_X1 U3617 ( .A1(n4315), .A2(n4393), .B1(n3992), .B2(n4288), .ZN(n3112)
         );
  NOR3_X1 U3618 ( .A1(n4000), .A2(n3112), .A3(n4700), .ZN(n2802) );
  NAND2_X1 U3619 ( .A1(n2803), .A2(n2802), .ZN(n2806) );
  INV_X1 U3620 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2804) );
  NAND2_X1 U3621 ( .A1(n4700), .A2(n2804), .ZN(n2805) );
  NAND2_X1 U3622 ( .A1(n2806), .A2(n2805), .ZN(n2811) );
  INV_X1 U3623 ( .A(n3998), .ZN(n2809) );
  NAND2_X1 U3624 ( .A1(n2809), .A2(n2808), .ZN(n2810) );
  NAND2_X1 U3625 ( .A1(n2811), .A2(n2810), .ZN(U3547) );
  NAND2_X1 U3626 ( .A1(n2812), .A2(n2252), .ZN(n2815) );
  NAND2_X1 U3627 ( .A1(n4587), .A2(n3062), .ZN(n2814) );
  AND2_X1 U3628 ( .A1(n4587), .A2(n2252), .ZN(n2817) );
  NAND2_X1 U3629 ( .A1(n2821), .A2(n2840), .ZN(n2819) );
  AOI22_X1 U3630 ( .A1(n3181), .A2(n2252), .B1(n2822), .B2(n2244), .ZN(n2818)
         );
  NAND2_X1 U3631 ( .A1(n2819), .A2(n2818), .ZN(n3178) );
  AND2_X1 U3632 ( .A1(n3181), .A2(n2247), .ZN(n2820) );
  NAND2_X1 U3633 ( .A1(n2822), .A2(REG1_REG_0__SCAN_IN), .ZN(n2823) );
  NAND2_X1 U3634 ( .A1(n2824), .A2(n2823), .ZN(n3179) );
  NAND2_X1 U3635 ( .A1(n3178), .A2(n3179), .ZN(n2826) );
  NAND2_X1 U3636 ( .A1(n2824), .A2(n3065), .ZN(n2825) );
  NAND2_X1 U3637 ( .A1(n2826), .A2(n2825), .ZN(n3184) );
  INV_X1 U3638 ( .A(n2827), .ZN(n2828) );
  NAND2_X1 U3639 ( .A1(n3907), .A2(n2252), .ZN(n2830) );
  NAND2_X1 U3640 ( .A1(n3702), .A2(n2247), .ZN(n2829) );
  NAND2_X1 U3641 ( .A1(n2830), .A2(n2829), .ZN(n2831) );
  XNOR2_X1 U3642 ( .A(n2831), .B(n3065), .ZN(n2834) );
  AOI21_X1 U3643 ( .B1(n3907), .B2(n2840), .A(n2832), .ZN(n2833) );
  NAND2_X1 U3644 ( .A1(n2834), .A2(n2833), .ZN(n2836) );
  NAND2_X1 U3645 ( .A1(n3696), .A2(n3697), .ZN(n3698) );
  NAND2_X1 U3646 ( .A1(n3698), .A2(n2836), .ZN(n3612) );
  NAND2_X1 U3647 ( .A1(n3905), .A2(n2252), .ZN(n2838) );
  NAND2_X1 U3648 ( .A1(n2697), .A2(n2247), .ZN(n2837) );
  AND2_X1 U3649 ( .A1(n2697), .A2(n2252), .ZN(n2841) );
  AOI21_X1 U3650 ( .B1(n3905), .B2(n2840), .A(n2841), .ZN(n2848) );
  XNOR2_X1 U3651 ( .A(n2847), .B(n2848), .ZN(n3613) );
  NAND2_X1 U3652 ( .A1(n3612), .A2(n3613), .ZN(n3219) );
  NAND2_X1 U3653 ( .A1(n3317), .A2(n2247), .ZN(n2843) );
  AND2_X1 U3654 ( .A1(n3317), .A2(n2252), .ZN(n2846) );
  AOI21_X1 U3655 ( .B1(n2842), .B2(n2840), .A(n2846), .ZN(n2851) );
  XNOR2_X1 U3656 ( .A(n2853), .B(n2851), .ZN(n3220) );
  INV_X1 U3657 ( .A(n2847), .ZN(n2849) );
  NAND2_X1 U3658 ( .A1(n2849), .A2(n2848), .ZN(n3221) );
  AND2_X1 U3659 ( .A1(n3220), .A2(n3221), .ZN(n2850) );
  INV_X1 U3660 ( .A(n2851), .ZN(n2852) );
  NAND2_X1 U3661 ( .A1(n2853), .A2(n2852), .ZN(n2854) );
  NAND2_X1 U3662 ( .A1(n3218), .A2(n2854), .ZN(n3277) );
  NAND2_X1 U3663 ( .A1(n3390), .A2(n2252), .ZN(n2856) );
  NAND2_X1 U3664 ( .A1(n3328), .A2(n2247), .ZN(n2855) );
  NAND2_X1 U3665 ( .A1(n2856), .A2(n2855), .ZN(n2857) );
  AND2_X1 U3666 ( .A1(n3328), .A2(n2252), .ZN(n2859) );
  AOI21_X1 U3667 ( .B1(n3390), .B2(n2840), .A(n2859), .ZN(n2860) );
  XNOR2_X1 U3668 ( .A(n2862), .B(n2860), .ZN(n3278) );
  NAND2_X1 U3669 ( .A1(n3277), .A2(n3278), .ZN(n2864) );
  INV_X1 U3670 ( .A(n2860), .ZN(n2861) );
  NAND2_X1 U3671 ( .A1(n2862), .A2(n2861), .ZN(n2863) );
  NAND2_X1 U3672 ( .A1(n3571), .A2(n2252), .ZN(n2866) );
  NAND2_X1 U3673 ( .A1(n2868), .A2(n3062), .ZN(n2865) );
  NAND2_X1 U3674 ( .A1(n2866), .A2(n2865), .ZN(n2867) );
  XNOR2_X1 U3675 ( .A(n2867), .B(n3069), .ZN(n2871) );
  NAND2_X1 U3676 ( .A1(n3571), .A2(n2840), .ZN(n2870) );
  NAND2_X1 U3677 ( .A1(n2868), .A2(n2252), .ZN(n2869) );
  NAND2_X1 U3678 ( .A1(n2870), .A2(n2869), .ZN(n2872) );
  AND2_X1 U3679 ( .A1(n2871), .A2(n2872), .ZN(n3286) );
  INV_X1 U3680 ( .A(n2871), .ZN(n2874) );
  INV_X1 U3681 ( .A(n2872), .ZN(n2873) );
  NAND2_X1 U3682 ( .A1(n2874), .A2(n2873), .ZN(n3285) );
  NAND2_X1 U3683 ( .A1(n3904), .A2(n2252), .ZN(n2876) );
  NAND2_X1 U3684 ( .A1(n3406), .A2(n3062), .ZN(n2875) );
  NAND2_X1 U3685 ( .A1(n2876), .A2(n2875), .ZN(n2877) );
  XNOR2_X1 U3686 ( .A(n2877), .B(n3065), .ZN(n2880) );
  AND2_X1 U3687 ( .A1(n3406), .A2(n2252), .ZN(n2878) );
  AOI21_X1 U3688 ( .B1(n3904), .B2(n2840), .A(n2878), .ZN(n2881) );
  XNOR2_X1 U3689 ( .A(n2880), .B(n2881), .ZN(n3568) );
  INV_X1 U3690 ( .A(n2880), .ZN(n2883) );
  INV_X1 U3691 ( .A(n2881), .ZN(n2882) );
  NAND2_X1 U3692 ( .A1(n2883), .A2(n2882), .ZN(n2884) );
  NAND2_X1 U3693 ( .A1(n3903), .A2(n2252), .ZN(n2886) );
  NAND2_X1 U3694 ( .A1(n3457), .A2(n2247), .ZN(n2885) );
  NAND2_X1 U3695 ( .A1(n2886), .A2(n2885), .ZN(n2887) );
  XNOR2_X1 U3696 ( .A(n2887), .B(n3069), .ZN(n2890) );
  NAND2_X1 U3697 ( .A1(n3903), .A2(n2840), .ZN(n2889) );
  NAND2_X1 U3698 ( .A1(n3457), .A2(n2252), .ZN(n2888) );
  NAND2_X1 U3699 ( .A1(n2889), .A2(n2888), .ZN(n2891) );
  AND2_X1 U3700 ( .A1(n2890), .A2(n2891), .ZN(n3432) );
  INV_X1 U3701 ( .A(n2890), .ZN(n2893) );
  INV_X1 U3702 ( .A(n2891), .ZN(n2892) );
  NAND2_X1 U3703 ( .A1(n2893), .A2(n2892), .ZN(n3431) );
  NAND2_X1 U3704 ( .A1(n3902), .A2(n2252), .ZN(n2895) );
  NAND2_X1 U3705 ( .A1(n3490), .A2(n2247), .ZN(n2894) );
  NAND2_X1 U3706 ( .A1(n2895), .A2(n2894), .ZN(n2896) );
  XNOR2_X1 U3707 ( .A(n2896), .B(n3069), .ZN(n2898) );
  AND2_X1 U3708 ( .A1(n3490), .A2(n2252), .ZN(n2897) );
  AOI21_X1 U3709 ( .B1(n3902), .B2(n2840), .A(n2897), .ZN(n2899) );
  XNOR2_X1 U3710 ( .A(n2898), .B(n2899), .ZN(n3548) );
  NAND2_X1 U3711 ( .A1(n3547), .A2(n3548), .ZN(n2902) );
  INV_X1 U3712 ( .A(n2898), .ZN(n2900) );
  NAND2_X1 U3713 ( .A1(n2900), .A2(n2899), .ZN(n2901) );
  NAND2_X1 U3714 ( .A1(n3901), .A2(n2252), .ZN(n2904) );
  NAND2_X1 U3715 ( .A1(n3476), .A2(n3062), .ZN(n2903) );
  NAND2_X1 U3716 ( .A1(n2904), .A2(n2903), .ZN(n2905) );
  XNOR2_X1 U3717 ( .A(n2905), .B(n3065), .ZN(n2908) );
  AND2_X1 U3718 ( .A1(n3476), .A2(n2252), .ZN(n2906) );
  AOI21_X1 U3719 ( .B1(n3901), .B2(n2840), .A(n2906), .ZN(n2909) );
  XNOR2_X1 U3720 ( .A(n2908), .B(n2909), .ZN(n5078) );
  INV_X1 U3721 ( .A(n2908), .ZN(n2911) );
  INV_X1 U3722 ( .A(n2909), .ZN(n2910) );
  NAND2_X1 U3723 ( .A1(n2911), .A2(n2910), .ZN(n2912) );
  NAND2_X1 U3724 ( .A1(n4413), .A2(n2840), .ZN(n2914) );
  NAND2_X1 U3725 ( .A1(n2915), .A2(n2252), .ZN(n2913) );
  NAND2_X1 U3726 ( .A1(n2914), .A2(n2913), .ZN(n3503) );
  NAND2_X1 U3727 ( .A1(n4413), .A2(n2252), .ZN(n2917) );
  NAND2_X1 U3728 ( .A1(n2915), .A2(n3062), .ZN(n2916) );
  NAND2_X1 U3729 ( .A1(n2917), .A2(n2916), .ZN(n2918) );
  XNOR2_X1 U3730 ( .A(n2918), .B(n3069), .ZN(n3502) );
  NAND2_X1 U3731 ( .A1(n4290), .A2(n2252), .ZN(n2920) );
  NAND2_X1 U3732 ( .A1(n4410), .A2(n2247), .ZN(n2919) );
  NAND2_X1 U3733 ( .A1(n2920), .A2(n2919), .ZN(n2921) );
  XNOR2_X1 U3734 ( .A(n2921), .B(n3069), .ZN(n2924) );
  NAND2_X1 U3735 ( .A1(n4290), .A2(n2840), .ZN(n2923) );
  NAND2_X1 U3736 ( .A1(n2923), .A2(n2922), .ZN(n2925) );
  AND2_X1 U3737 ( .A1(n2924), .A2(n2925), .ZN(n3539) );
  INV_X1 U3738 ( .A(n2924), .ZN(n2927) );
  INV_X1 U3739 ( .A(n2925), .ZN(n2926) );
  NAND2_X1 U3740 ( .A1(n2931), .A2(n2247), .ZN(n2928) );
  NAND2_X1 U3741 ( .A1(n2929), .A2(n2928), .ZN(n2930) );
  NAND2_X1 U3742 ( .A1(n4412), .A2(n2840), .ZN(n2933) );
  NAND2_X1 U3743 ( .A1(n2931), .A2(n2252), .ZN(n2932) );
  NAND2_X1 U3744 ( .A1(n2933), .A2(n2932), .ZN(n3557) );
  NAND2_X1 U3745 ( .A1(n2934), .A2(n3557), .ZN(n2938) );
  INV_X1 U3746 ( .A(n3555), .ZN(n2936) );
  INV_X1 U3747 ( .A(n3556), .ZN(n2935) );
  NAND2_X1 U3748 ( .A1(n2936), .A2(n2935), .ZN(n2937) );
  NAND2_X1 U3749 ( .A1(n4251), .A2(n2252), .ZN(n2940) );
  NAND2_X1 U3750 ( .A1(n2942), .A2(n3062), .ZN(n2939) );
  NAND2_X1 U3751 ( .A1(n2940), .A2(n2939), .ZN(n2941) );
  XNOR2_X1 U3752 ( .A(n2941), .B(n3069), .ZN(n2945) );
  NAND2_X1 U3753 ( .A1(n4251), .A2(n2840), .ZN(n2944) );
  NAND2_X1 U3754 ( .A1(n2944), .A2(n2943), .ZN(n2946) );
  NAND2_X1 U3755 ( .A1(n2945), .A2(n2946), .ZN(n3587) );
  INV_X1 U3756 ( .A(n2945), .ZN(n2948) );
  INV_X1 U3757 ( .A(n2946), .ZN(n2947) );
  NAND2_X1 U3758 ( .A1(n2948), .A2(n2947), .ZN(n3586) );
  NAND2_X1 U3759 ( .A1(n4266), .A2(n2252), .ZN(n2950) );
  NAND2_X1 U3760 ( .A1(n4389), .A2(n2247), .ZN(n2949) );
  NAND2_X1 U3761 ( .A1(n2950), .A2(n2949), .ZN(n2951) );
  XNOR2_X1 U3762 ( .A(n2951), .B(n3065), .ZN(n2958) );
  NAND2_X1 U3763 ( .A1(n4266), .A2(n2840), .ZN(n2953) );
  NAND2_X1 U3764 ( .A1(n2953), .A2(n2952), .ZN(n3649) );
  NAND2_X1 U3765 ( .A1(n3650), .A2(n3649), .ZN(n2959) );
  NAND2_X1 U3766 ( .A1(n4390), .A2(n2252), .ZN(n2955) );
  NAND2_X1 U3767 ( .A1(n4379), .A2(n3062), .ZN(n2954) );
  NAND2_X1 U3768 ( .A1(n2955), .A2(n2954), .ZN(n2956) );
  XNOR2_X1 U3769 ( .A(n2956), .B(n3069), .ZN(n2960) );
  AND2_X1 U3770 ( .A1(n4379), .A2(n2252), .ZN(n2957) );
  AOI21_X1 U3771 ( .B1(n4390), .B2(n2840), .A(n2957), .ZN(n2961) );
  NAND3_X1 U3772 ( .A1(n2959), .A2(n3652), .A3(n3648), .ZN(n2964) );
  INV_X1 U3773 ( .A(n2960), .ZN(n2962) );
  NAND2_X1 U3774 ( .A1(n2962), .A2(n2961), .ZN(n2963) );
  NAND2_X1 U3775 ( .A1(n4380), .A2(n2252), .ZN(n2966) );
  OR2_X1 U3776 ( .A1(n4215), .A2(n3068), .ZN(n2965) );
  NAND2_X1 U3777 ( .A1(n2966), .A2(n2965), .ZN(n2967) );
  XNOR2_X1 U3778 ( .A(n2967), .B(n3065), .ZN(n3659) );
  NOR2_X1 U3779 ( .A1(n4215), .A2(n3071), .ZN(n2968) );
  AOI21_X1 U3780 ( .B1(n4380), .B2(n2840), .A(n2968), .ZN(n3658) );
  INV_X1 U3781 ( .A(n3659), .ZN(n2970) );
  INV_X1 U3782 ( .A(n3658), .ZN(n2969) );
  NAND2_X1 U3783 ( .A1(n2970), .A2(n2969), .ZN(n2971) );
  NAND2_X1 U3784 ( .A1(n4188), .A2(n3062), .ZN(n2972) );
  NAND2_X1 U3785 ( .A1(n2973), .A2(n2972), .ZN(n2974) );
  XNOR2_X1 U3786 ( .A(n2974), .B(n3069), .ZN(n2977) );
  NAND2_X1 U3787 ( .A1(n4372), .A2(n2840), .ZN(n2976) );
  NAND2_X1 U3788 ( .A1(n4188), .A2(n2252), .ZN(n2975) );
  NAND2_X1 U3789 ( .A1(n2976), .A2(n2975), .ZN(n2978) );
  INV_X1 U3790 ( .A(n2977), .ZN(n2980) );
  INV_X1 U3791 ( .A(n2978), .ZN(n2979) );
  NAND2_X1 U3792 ( .A1(n2980), .A2(n2979), .ZN(n3708) );
  NAND2_X1 U3793 ( .A1(n4189), .A2(n2252), .ZN(n2982) );
  NAND2_X1 U3794 ( .A1(n4172), .A2(n2247), .ZN(n2981) );
  NAND2_X1 U3795 ( .A1(n2982), .A2(n2981), .ZN(n2983) );
  XNOR2_X1 U3796 ( .A(n2983), .B(n3069), .ZN(n3007) );
  AOI21_X1 U3797 ( .B1(n4189), .B2(n2840), .A(n2984), .ZN(n3008) );
  XNOR2_X1 U3798 ( .A(n3007), .B(n3008), .ZN(n3623) );
  NAND2_X1 U3799 ( .A1(n4131), .A2(n2252), .ZN(n2986) );
  OR2_X1 U3800 ( .A1(n3680), .A2(n3068), .ZN(n2985) );
  NAND2_X1 U3801 ( .A1(n2986), .A2(n2985), .ZN(n2987) );
  XNOR2_X1 U3802 ( .A(n2987), .B(n3069), .ZN(n3005) );
  INV_X1 U3803 ( .A(n3005), .ZN(n2991) );
  NAND2_X1 U3804 ( .A1(n4131), .A2(n2840), .ZN(n2989) );
  NAND2_X1 U3805 ( .A1(n4151), .A2(n2252), .ZN(n2988) );
  NAND2_X1 U3806 ( .A1(n2989), .A2(n2988), .ZN(n3004) );
  INV_X1 U3807 ( .A(n3004), .ZN(n2990) );
  NAND2_X1 U3808 ( .A1(n2991), .A2(n2990), .ZN(n3678) );
  NAND2_X1 U3809 ( .A1(n4143), .A2(n2252), .ZN(n2993) );
  OR2_X1 U3810 ( .A1(n4135), .A2(n3068), .ZN(n2992) );
  NAND2_X1 U3811 ( .A1(n2993), .A2(n2992), .ZN(n2994) );
  XNOR2_X1 U3812 ( .A(n2994), .B(n3065), .ZN(n3629) );
  NOR2_X1 U3813 ( .A1(n4135), .A2(n3071), .ZN(n2995) );
  AOI21_X1 U3814 ( .B1(n4143), .B2(n2840), .A(n2995), .ZN(n3628) );
  AND2_X1 U3815 ( .A1(n3629), .A2(n3628), .ZN(n3602) );
  NAND2_X1 U3816 ( .A1(n4335), .A2(n2252), .ZN(n2997) );
  OR2_X1 U3817 ( .A1(n4098), .A2(n3068), .ZN(n2996) );
  NAND2_X1 U3818 ( .A1(n2997), .A2(n2996), .ZN(n2998) );
  XNOR2_X1 U3819 ( .A(n2998), .B(n3069), .ZN(n3023) );
  NOR2_X1 U3820 ( .A1(n4098), .A2(n3071), .ZN(n2999) );
  AOI21_X1 U3821 ( .B1(n4335), .B2(n2840), .A(n2999), .ZN(n3021) );
  XNOR2_X1 U3822 ( .A(n3023), .B(n3021), .ZN(n3604) );
  NAND2_X1 U3823 ( .A1(n4352), .A2(n2252), .ZN(n3001) );
  OR2_X1 U3824 ( .A1(n4112), .A2(n3068), .ZN(n3000) );
  NAND2_X1 U3825 ( .A1(n3001), .A2(n3000), .ZN(n3002) );
  XNOR2_X1 U3826 ( .A(n3002), .B(n3065), .ZN(n3016) );
  NOR2_X1 U3827 ( .A1(n4112), .A2(n3071), .ZN(n3003) );
  AOI21_X1 U3828 ( .B1(n4352), .B2(n2840), .A(n3003), .ZN(n3015) );
  NAND2_X1 U3829 ( .A1(n3016), .A2(n3015), .ZN(n3605) );
  NAND2_X1 U3830 ( .A1(n3604), .A2(n3605), .ZN(n3020) );
  AND2_X1 U3831 ( .A1(n3678), .A2(n2357), .ZN(n3010) );
  INV_X1 U3832 ( .A(n3010), .ZN(n3034) );
  NAND2_X1 U3833 ( .A1(n3005), .A2(n3004), .ZN(n3676) );
  OR2_X1 U3834 ( .A1(n3034), .A2(n3676), .ZN(n3006) );
  INV_X1 U3835 ( .A(n3006), .ZN(n3012) );
  INV_X1 U3836 ( .A(n3007), .ZN(n3009) );
  NAND2_X1 U3837 ( .A1(n3009), .A2(n3008), .ZN(n3600) );
  AND2_X1 U3838 ( .A1(n3600), .A2(n3010), .ZN(n3011) );
  OR2_X1 U3839 ( .A1(n3012), .A2(n3011), .ZN(n3013) );
  NAND2_X1 U3840 ( .A1(n3014), .A2(n3013), .ZN(n3596) );
  XNOR2_X1 U3841 ( .A(n3016), .B(n3015), .ZN(n3689) );
  INV_X1 U3842 ( .A(n3689), .ZN(n3019) );
  INV_X1 U3843 ( .A(n3629), .ZN(n3018) );
  INV_X1 U3844 ( .A(n3628), .ZN(n3017) );
  NAND2_X1 U3845 ( .A1(n3018), .A2(n3017), .ZN(n3685) );
  NOR2_X1 U3846 ( .A1(n3020), .A2(n3603), .ZN(n3597) );
  INV_X1 U3847 ( .A(n3021), .ZN(n3022) );
  NAND2_X1 U3848 ( .A1(n3023), .A2(n3022), .ZN(n3030) );
  NOR2_X1 U3849 ( .A1(n4080), .A2(n3071), .ZN(n3024) );
  AOI21_X1 U3850 ( .B1(n4058), .B2(n2840), .A(n3024), .ZN(n3033) );
  NAND2_X1 U3851 ( .A1(n3030), .A2(n3033), .ZN(n3025) );
  NOR2_X1 U3852 ( .A1(n3597), .A2(n3025), .ZN(n3026) );
  NAND2_X1 U3853 ( .A1(n3596), .A2(n3026), .ZN(n3666) );
  OR2_X1 U3854 ( .A1(n4080), .A2(n3068), .ZN(n3027) );
  NAND2_X1 U3855 ( .A1(n3028), .A2(n3027), .ZN(n3029) );
  NAND2_X1 U3856 ( .A1(n3666), .A2(n3668), .ZN(n3042) );
  INV_X1 U3857 ( .A(n3030), .ZN(n3031) );
  NOR2_X1 U3858 ( .A1(n3597), .A2(n3031), .ZN(n3032) );
  OR2_X1 U3859 ( .A1(n3033), .A2(n3032), .ZN(n3038) );
  INV_X1 U3860 ( .A(n3038), .ZN(n3036) );
  NOR2_X1 U3861 ( .A1(n3034), .A2(n3033), .ZN(n3035) );
  OR2_X1 U3862 ( .A1(n3036), .A2(n3035), .ZN(n3037) );
  AND2_X1 U3863 ( .A1(n3600), .A2(n3037), .ZN(n3041) );
  INV_X1 U3864 ( .A(n3037), .ZN(n3040) );
  AND2_X1 U3865 ( .A1(n3676), .A2(n3038), .ZN(n3039) );
  NAND2_X1 U3866 ( .A1(n3042), .A2(n3665), .ZN(n3639) );
  NAND2_X1 U3867 ( .A1(n4322), .A2(n2252), .ZN(n3044) );
  OR2_X1 U3868 ( .A1(n4065), .A2(n3068), .ZN(n3043) );
  NAND2_X1 U3869 ( .A1(n3044), .A2(n3043), .ZN(n3045) );
  XNOR2_X1 U3870 ( .A(n3045), .B(n3065), .ZN(n3047) );
  NOR2_X1 U3871 ( .A1(n4065), .A2(n3071), .ZN(n3046) );
  AOI21_X1 U3872 ( .B1(n4322), .B2(n2840), .A(n3046), .ZN(n3048) );
  NAND2_X1 U3873 ( .A1(n3047), .A2(n3048), .ZN(n3637) );
  INV_X1 U3874 ( .A(n3047), .ZN(n3050) );
  INV_X1 U3875 ( .A(n3048), .ZN(n3049) );
  NAND2_X1 U3876 ( .A1(n3050), .A2(n3049), .ZN(n3638) );
  OR2_X1 U3877 ( .A1(n4048), .A2(n3068), .ZN(n3051) );
  NAND2_X1 U3878 ( .A1(n3052), .A2(n3051), .ZN(n3053) );
  XNOR2_X1 U3879 ( .A(n3053), .B(n3069), .ZN(n3057) );
  NAND2_X1 U3880 ( .A1(n4313), .A2(n2840), .ZN(n3055) );
  NAND2_X1 U3881 ( .A1(n3055), .A2(n3054), .ZN(n3058) );
  AND2_X1 U3882 ( .A1(n3057), .A2(n3058), .ZN(n3719) );
  INV_X1 U3883 ( .A(n3719), .ZN(n3056) );
  INV_X1 U3884 ( .A(n3057), .ZN(n3060) );
  INV_X1 U3885 ( .A(n3058), .ZN(n3059) );
  NAND2_X1 U3886 ( .A1(n3060), .A2(n3059), .ZN(n3718) );
  NAND2_X1 U3887 ( .A1(n4044), .A2(n2252), .ZN(n3064) );
  NAND2_X1 U3888 ( .A1(n4312), .A2(n2247), .ZN(n3063) );
  NAND2_X1 U3889 ( .A1(n3064), .A2(n3063), .ZN(n3066) );
  XNOR2_X1 U3890 ( .A(n3066), .B(n3065), .ZN(n3074) );
  AND2_X1 U3891 ( .A1(n4312), .A2(n2252), .ZN(n3067) );
  AOI21_X1 U3892 ( .B1(n4044), .B2(n2840), .A(n3067), .ZN(n3075) );
  XNOR2_X1 U3893 ( .A(n3074), .B(n3075), .ZN(n3578) );
  NOR2_X1 U3894 ( .A1(n3579), .A2(n3578), .ZN(n3087) );
  INV_X1 U3895 ( .A(n3087), .ZN(n3086) );
  OAI22_X1 U3896 ( .A1(n4315), .A2(n3071), .B1(n3068), .B2(n4008), .ZN(n3070)
         );
  XNOR2_X1 U3897 ( .A(n3070), .B(n3069), .ZN(n3073) );
  OAI22_X1 U3898 ( .A1(n4315), .A2(n2858), .B1(n3071), .B2(n4008), .ZN(n3072)
         );
  XNOR2_X1 U3899 ( .A(n3073), .B(n3072), .ZN(n3090) );
  INV_X1 U3900 ( .A(n3090), .ZN(n3085) );
  INV_X1 U3901 ( .A(n3074), .ZN(n3077) );
  INV_X1 U3902 ( .A(n3075), .ZN(n3076) );
  NAND2_X1 U3903 ( .A1(n3077), .A2(n3076), .ZN(n3088) );
  INV_X1 U3904 ( .A(n3078), .ZN(n3236) );
  NAND3_X1 U3905 ( .A1(n3236), .A2(n3079), .A3(n3233), .ZN(n3104) );
  NAND2_X1 U3906 ( .A1(n3080), .A2(n4605), .ZN(n3082) );
  INV_X1 U3907 ( .A(n3126), .ZN(n3081) );
  NAND3_X1 U3908 ( .A1(n3082), .A2(n3129), .A3(n3081), .ZN(n3083) );
  NAND2_X1 U3909 ( .A1(n3086), .A2(n2351), .ZN(n3111) );
  NAND3_X1 U3910 ( .A1(n3087), .A2(n3699), .A3(n3090), .ZN(n3110) );
  INV_X1 U3911 ( .A(n3088), .ZN(n3089) );
  NAND3_X1 U3912 ( .A1(n3090), .A2(n3699), .A3(n3089), .ZN(n3109) );
  NAND2_X1 U3913 ( .A1(n3104), .A2(n3091), .ZN(n3180) );
  AND3_X1 U3914 ( .A1(n3092), .A2(n3128), .A3(n3118), .ZN(n3093) );
  NAND2_X1 U3915 ( .A1(n3180), .A2(n3093), .ZN(n3094) );
  INV_X1 U3916 ( .A(n3104), .ZN(n3096) );
  AND2_X1 U3917 ( .A1(n4588), .A2(n3129), .ZN(n3095) );
  NAND2_X1 U3918 ( .A1(n3096), .A2(n3095), .ZN(n3099) );
  AND2_X2 U3919 ( .A1(n3099), .A2(n4276), .ZN(n3733) );
  OAI22_X1 U3920 ( .A1(n3733), .A2(n4008), .B1(STATE_REG_SCAN_IN), .B2(n3100), 
        .ZN(n3107) );
  INV_X1 U3921 ( .A(n3101), .ZN(n3102) );
  NAND3_X1 U3922 ( .A1(n2252), .A2(n3103), .A3(n3102), .ZN(n3893) );
  INV_X1 U3923 ( .A(n3900), .ZN(n4010) );
  OAI22_X1 U3924 ( .A1(n4325), .A2(n5081), .B1(n4010), .B2(n5080), .ZN(n3106)
         );
  AOI211_X1 U3925 ( .C1(n4006), .C2(n3736), .A(n3107), .B(n3106), .ZN(n3108)
         );
  NAND3_X1 U3926 ( .A1(n3111), .A2(n3110), .A3(n2359), .ZN(U3217) );
  AOI211_X1 U3927 ( .C1(n3991), .C2(n4665), .A(n4000), .B(n3112), .ZN(n3117)
         );
  NOR2_X1 U3928 ( .A1(n3998), .A2(n4472), .ZN(n3115) );
  INV_X1 U3929 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3113) );
  NOR2_X1 U3930 ( .A1(n3115), .A2(n3114), .ZN(n3116) );
  OAI21_X1 U3931 ( .B1(n3117), .B2(n4684), .A(n3116), .ZN(U3515) );
  INV_X1 U3932 ( .A(DATAI_27_), .ZN(n4784) );
  INV_X1 U3933 ( .A(n3908), .ZN(n3190) );
  NAND2_X1 U3934 ( .A1(n3190), .A2(STATE_REG_SCAN_IN), .ZN(n3119) );
  OAI21_X1 U3935 ( .B1(STATE_REG_SCAN_IN), .B2(n4784), .A(n3119), .ZN(U3325)
         );
  INV_X1 U3936 ( .A(DATAI_29_), .ZN(n4953) );
  NAND2_X1 U3937 ( .A1(n3120), .A2(STATE_REG_SCAN_IN), .ZN(n3121) );
  OAI21_X1 U3938 ( .B1(STATE_REG_SCAN_IN), .B2(n4953), .A(n3121), .ZN(U3323)
         );
  INV_X1 U3939 ( .A(D_REG_1__SCAN_IN), .ZN(n3124) );
  NOR3_X1 U3940 ( .A1(n2754), .A2(n4480), .A3(n4625), .ZN(n3123) );
  AOI21_X1 U3941 ( .B1(n4622), .B2(n3124), .A(n3123), .ZN(U3459) );
  NOR3_X1 U3942 ( .A1(n4481), .A2(n2754), .A3(n4625), .ZN(n3125) );
  AOI21_X1 U3943 ( .B1(n4622), .B2(n2766), .A(n3125), .ZN(U3458) );
  NAND2_X1 U3944 ( .A1(n3128), .A2(n3126), .ZN(n3127) );
  INV_X1 U3945 ( .A(n3150), .ZN(n3130) );
  NOR2_X1 U3946 ( .A1(n3128), .A2(U3149), .ZN(n3891) );
  NOR2_X1 U3947 ( .A1(n4579), .A2(U4043), .ZN(U3148) );
  INV_X1 U3948 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n4937) );
  NAND2_X1 U3949 ( .A1(n2821), .A2(U4043), .ZN(n3131) );
  OAI21_X1 U3950 ( .B1(U4043), .B2(n4937), .A(n3131), .ZN(U3550) );
  INV_X1 U3951 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n4857) );
  NAND2_X1 U3952 ( .A1(n2812), .A2(U4043), .ZN(n3132) );
  OAI21_X1 U3953 ( .B1(U4043), .B2(n4857), .A(n3132), .ZN(U3551) );
  INV_X1 U3954 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4923) );
  NAND2_X1 U3955 ( .A1(n4131), .A2(U4043), .ZN(n3133) );
  OAI21_X1 U3956 ( .B1(U4043), .B2(n4923), .A(n3133), .ZN(U3570) );
  INV_X1 U3957 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4856) );
  NAND2_X1 U3958 ( .A1(n4380), .A2(U4043), .ZN(n3134) );
  OAI21_X1 U3959 ( .B1(U4043), .B2(n4856), .A(n3134), .ZN(U3567) );
  INV_X1 U3960 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n4972) );
  NAND2_X1 U3961 ( .A1(n3571), .A2(U4043), .ZN(n3135) );
  OAI21_X1 U3962 ( .B1(U4043), .B2(n4972), .A(n3135), .ZN(U3556) );
  INV_X1 U3963 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n4951) );
  NAND2_X1 U3964 ( .A1(n3390), .A2(U4043), .ZN(n3136) );
  OAI21_X1 U3965 ( .B1(U4043), .B2(n4951), .A(n3136), .ZN(U3555) );
  INV_X1 U3966 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n4948) );
  NAND2_X1 U3967 ( .A1(n4390), .A2(U4043), .ZN(n3137) );
  OAI21_X1 U3968 ( .B1(U4043), .B2(n4948), .A(n3137), .ZN(U3566) );
  INV_X1 U3969 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3138) );
  AND2_X1 U3970 ( .A1(REG2_REG_0__SCAN_IN), .A2(n2244), .ZN(n3139) );
  NAND2_X1 U3971 ( .A1(n4496), .A2(REG2_REG_1__SCAN_IN), .ZN(n3196) );
  INV_X1 U3972 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3271) );
  MUX2_X1 U3973 ( .A(REG2_REG_2__SCAN_IN), .B(n3271), .S(n4495), .Z(n3140) );
  NAND2_X1 U3974 ( .A1(n4495), .A2(REG2_REG_2__SCAN_IN), .ZN(n3141) );
  NAND2_X1 U3975 ( .A1(n3199), .A2(n3141), .ZN(n3142) );
  INV_X1 U3976 ( .A(n4494), .ZN(n3170) );
  XNOR2_X1 U3977 ( .A(n3142), .B(n3170), .ZN(n3169) );
  NAND2_X1 U3978 ( .A1(n3169), .A2(REG2_REG_3__SCAN_IN), .ZN(n3144) );
  NAND2_X1 U3979 ( .A1(n3142), .A2(n4494), .ZN(n3143) );
  NAND2_X1 U3980 ( .A1(n3146), .A2(n4493), .ZN(n3147) );
  INV_X1 U3981 ( .A(n3153), .ZN(n3149) );
  MUX2_X1 U3982 ( .A(n3337), .B(REG2_REG_5__SCAN_IN), .S(n4492), .Z(n3148) );
  MUX2_X1 U3983 ( .A(REG2_REG_5__SCAN_IN), .B(n3337), .S(n4492), .Z(n3154) );
  NAND2_X1 U3984 ( .A1(n4479), .A2(n3190), .ZN(n3894) );
  INV_X1 U3985 ( .A(n3894), .ZN(n3152) );
  OAI21_X1 U3986 ( .B1(n3154), .B2(n3153), .A(n4563), .ZN(n3168) );
  AND2_X1 U3987 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3280) );
  INV_X1 U3988 ( .A(n4492), .ZN(n3363) );
  NOR2_X1 U3989 ( .A1(n4585), .A2(n3363), .ZN(n3155) );
  AOI211_X1 U3990 ( .C1(n4579), .C2(ADDR_REG_5__SCAN_IN), .A(n3280), .B(n3155), 
        .ZN(n3167) );
  XOR2_X1 U3991 ( .A(REG1_REG_5__SCAN_IN), .B(n4492), .Z(n3165) );
  INV_X1 U3992 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3156) );
  MUX2_X1 U3993 ( .A(REG1_REG_2__SCAN_IN), .B(n3156), .S(n4495), .Z(n3202) );
  INV_X1 U3994 ( .A(REG1_REG_1__SCAN_IN), .ZN(n3157) );
  AND2_X1 U3995 ( .A1(n2244), .A2(REG1_REG_0__SCAN_IN), .ZN(n3920) );
  NAND2_X1 U3996 ( .A1(n4496), .A2(REG1_REG_1__SCAN_IN), .ZN(n3158) );
  NAND2_X1 U3997 ( .A1(n3919), .A2(n3158), .ZN(n3201) );
  NAND2_X1 U3998 ( .A1(n3202), .A2(n3201), .ZN(n3200) );
  NAND2_X1 U3999 ( .A1(n4495), .A2(REG1_REG_2__SCAN_IN), .ZN(n3159) );
  NAND2_X1 U4000 ( .A1(n3200), .A2(n3159), .ZN(n3160) );
  XNOR2_X1 U4001 ( .A(n3160), .B(n3170), .ZN(n3173) );
  NAND2_X1 U4002 ( .A1(n3173), .A2(REG1_REG_3__SCAN_IN), .ZN(n3172) );
  NAND2_X1 U4003 ( .A1(n3160), .A2(n4494), .ZN(n3161) );
  NAND2_X1 U4004 ( .A1(n3172), .A2(n3161), .ZN(n3162) );
  INV_X1 U4005 ( .A(n3162), .ZN(n3163) );
  INV_X1 U4006 ( .A(n4493), .ZN(n3213) );
  XNOR2_X1 U4007 ( .A(n3162), .B(n3213), .ZN(n3210) );
  OAI211_X1 U4008 ( .C1(n3165), .C2(n3164), .A(n4581), .B(n3362), .ZN(n3166)
         );
  OAI211_X1 U4009 ( .C1(n3339), .C2(n3168), .A(n3167), .B(n3166), .ZN(U3245)
         );
  XNOR2_X1 U4010 ( .A(n3169), .B(REG2_REG_3__SCAN_IN), .ZN(n3176) );
  NOR2_X1 U4011 ( .A1(STATE_REG_SCAN_IN), .A2(n3618), .ZN(n3617) );
  NOR2_X1 U4012 ( .A1(n4585), .A2(n3170), .ZN(n3171) );
  AOI211_X1 U4013 ( .C1(n4579), .C2(ADDR_REG_3__SCAN_IN), .A(n3617), .B(n3171), 
        .ZN(n3175) );
  OAI211_X1 U4014 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3173), .A(n4581), .B(n3172), 
        .ZN(n3174) );
  OAI211_X1 U4015 ( .C1(n3176), .C2(n4574), .A(n3175), .B(n3174), .ZN(U3243)
         );
  XOR2_X1 U4016 ( .A(n3178), .B(n3179), .Z(n3191) );
  NAND2_X1 U4017 ( .A1(n3191), .A2(n3699), .ZN(n3183) );
  INV_X1 U4018 ( .A(n3733), .ZN(n3703) );
  NAND2_X1 U4019 ( .A1(n3180), .A2(n3235), .ZN(n3701) );
  AOI22_X1 U4020 ( .A1(n3703), .A2(n3181), .B1(REG3_REG_0__SCAN_IN), .B2(n3701), .ZN(n3182) );
  OAI211_X1 U4021 ( .C1(n3177), .C2(n5080), .A(n3183), .B(n3182), .ZN(U3229)
         );
  XNOR2_X1 U4022 ( .A(n3185), .B(n3184), .ZN(n3188) );
  AOI22_X1 U4023 ( .A1(n3703), .A2(n4587), .B1(REG3_REG_1__SCAN_IN), .B2(n3701), .ZN(n3187) );
  AOI22_X1 U4024 ( .A1(n3731), .A2(n2821), .B1(n3732), .B2(n3907), .ZN(n3186)
         );
  OAI211_X1 U4025 ( .C1(n3188), .C2(n5077), .A(n3187), .B(n3186), .ZN(U3219)
         );
  NOR3_X1 U4026 ( .A1(n3191), .A2(n3190), .A3(n3189), .ZN(n3195) );
  OR2_X1 U4027 ( .A1(n3908), .A2(REG2_REG_0__SCAN_IN), .ZN(n3192) );
  NAND2_X1 U4028 ( .A1(n4479), .A2(n3192), .ZN(n3909) );
  NOR2_X1 U4029 ( .A1(n3894), .A2(n2377), .ZN(n3193) );
  MUX2_X1 U4030 ( .A(n3909), .B(n3193), .S(n2244), .Z(n3194) );
  NOR3_X1 U4031 ( .A1(n3195), .A2(n3194), .A3(n3906), .ZN(n3214) );
  MUX2_X1 U4032 ( .A(n3271), .B(REG2_REG_2__SCAN_IN), .S(n4495), .Z(n3197) );
  NAND3_X1 U4033 ( .A1(n3197), .A2(n3918), .A3(n3196), .ZN(n3198) );
  NAND3_X1 U4034 ( .A1(n4563), .A2(n3199), .A3(n3198), .ZN(n3206) );
  AOI22_X1 U4035 ( .A1(n4579), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3205) );
  INV_X1 U4036 ( .A(n4585), .ZN(n3949) );
  NAND2_X1 U4037 ( .A1(n3949), .A2(n4495), .ZN(n3204) );
  OAI211_X1 U4038 ( .C1(n3202), .C2(n3201), .A(n4581), .B(n3200), .ZN(n3203)
         );
  NAND4_X1 U4039 ( .A1(n3206), .A2(n3205), .A3(n3204), .A4(n3203), .ZN(n3207)
         );
  OR2_X1 U4040 ( .A1(n3214), .A2(n3207), .ZN(U3242) );
  XNOR2_X1 U4041 ( .A(n3208), .B(REG2_REG_4__SCAN_IN), .ZN(n3216) );
  OAI211_X1 U4042 ( .C1(n3210), .C2(REG1_REG_4__SCAN_IN), .A(n4581), .B(n3209), 
        .ZN(n3212) );
  AND2_X1 U40430 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3224) );
  AOI21_X1 U4044 ( .B1(n4579), .B2(ADDR_REG_4__SCAN_IN), .A(n3224), .ZN(n3211)
         );
  OAI211_X1 U4045 ( .C1(n4585), .C2(n3213), .A(n3212), .B(n3211), .ZN(n3215)
         );
  AOI211_X1 U4046 ( .C1(n4563), .C2(n3216), .A(n3215), .B(n3214), .ZN(n3217)
         );
  INV_X1 U4047 ( .A(n3217), .ZN(U3244) );
  NAND2_X1 U4048 ( .A1(n3218), .A2(n3699), .ZN(n3228) );
  AOI21_X1 U4049 ( .B1(n3219), .B2(n3221), .A(n3220), .ZN(n3227) );
  AOI22_X1 U4050 ( .A1(n3732), .A2(n3390), .B1(n3731), .B2(n3905), .ZN(n3226)
         );
  NOR2_X1 U4051 ( .A1(n3733), .A2(n3222), .ZN(n3223) );
  AOI211_X1 U4052 ( .C1(n3736), .C2(n3324), .A(n3224), .B(n3223), .ZN(n3225)
         );
  OAI211_X1 U4053 ( .C1(n3228), .C2(n3227), .A(n3226), .B(n3225), .ZN(U3227)
         );
  INV_X1 U4054 ( .A(n3230), .ZN(n3231) );
  NAND2_X1 U4055 ( .A1(n3229), .A2(n3231), .ZN(n3313) );
  XNOR2_X1 U4056 ( .A(n3313), .B(n3796), .ZN(n3254) );
  INV_X1 U4057 ( .A(n3254), .ZN(n3250) );
  NAND4_X1 U4058 ( .A1(n3236), .A2(n3235), .A3(n3234), .A4(n3233), .ZN(n3237)
         );
  OR2_X1 U4059 ( .A1(n2813), .A2(n3981), .ZN(n3259) );
  NAND2_X1 U4060 ( .A1(n4594), .A2(n3259), .ZN(n3238) );
  NAND3_X1 U4061 ( .A1(n3240), .A2(n3820), .A3(n3796), .ZN(n3241) );
  AOI21_X1 U4062 ( .B1(n3239), .B2(n3241), .A(n4292), .ZN(n3252) );
  XNOR2_X1 U4063 ( .A(n3308), .B(n3615), .ZN(n3381) );
  INV_X1 U4064 ( .A(n3381), .ZN(n3247) );
  NAND2_X1 U4065 ( .A1(n4617), .A2(n3981), .ZN(n4197) );
  AND2_X1 U4066 ( .A1(n4617), .A2(n4588), .ZN(n3995) );
  OAI22_X1 U4067 ( .A1(n4617), .A2(n3242), .B1(n4276), .B2(REG3_REG_3__SCAN_IN), .ZN(n3245) );
  NAND2_X1 U4068 ( .A1(n4617), .A2(n4589), .ZN(n4011) );
  NAND2_X1 U4069 ( .A1(n4617), .A2(n4411), .ZN(n4009) );
  OAI22_X1 U4070 ( .A1(n3243), .A2(n4011), .B1(n3330), .B2(n4009), .ZN(n3244)
         );
  AOI211_X1 U4071 ( .C1(n2697), .C2(n3995), .A(n3245), .B(n3244), .ZN(n3246)
         );
  OAI21_X1 U4072 ( .B1(n3247), .B2(n4300), .A(n3246), .ZN(n3248) );
  AOI21_X1 U4073 ( .B1(n3252), .B2(n4617), .A(n3248), .ZN(n3249) );
  OAI21_X1 U4074 ( .B1(n3250), .B2(n4241), .A(n3249), .ZN(U3287) );
  AOI22_X1 U4075 ( .A1(n2842), .A2(n4411), .B1(n4588), .B2(n2697), .ZN(n3251)
         );
  OAI21_X1 U4076 ( .B1(n3243), .B2(n4393), .A(n3251), .ZN(n3253) );
  AOI211_X1 U4077 ( .C1(n4665), .C2(n3254), .A(n3253), .B(n3252), .ZN(n3383)
         );
  INV_X1 U4078 ( .A(n4472), .ZN(n4651) );
  AOI22_X1 U4079 ( .A1(n4651), .A2(n3381), .B1(REG0_REG_3__SCAN_IN), .B2(n4684), .ZN(n3255) );
  OAI21_X1 U4080 ( .B1(n3383), .B2(n4684), .A(n3255), .ZN(U3473) );
  NAND2_X1 U4081 ( .A1(n3257), .A2(n3256), .ZN(n3258) );
  NAND2_X1 U4082 ( .A1(n3229), .A2(n3258), .ZN(n4650) );
  INV_X1 U4083 ( .A(n4650), .ZN(n3276) );
  INV_X1 U4084 ( .A(n3259), .ZN(n3260) );
  INV_X1 U4085 ( .A(n4615), .ZN(n3275) );
  NAND3_X1 U4086 ( .A1(n3799), .A2(n2695), .A3(n3262), .ZN(n3263) );
  NAND2_X1 U4087 ( .A1(n3240), .A2(n3263), .ZN(n3268) );
  NAND2_X1 U4088 ( .A1(n2812), .A2(n4589), .ZN(n3265) );
  NAND2_X1 U4089 ( .A1(n3905), .A2(n4411), .ZN(n3264) );
  OAI211_X1 U4090 ( .C1(n4288), .C2(n3266), .A(n3265), .B(n3264), .ZN(n3267)
         );
  AOI21_X1 U4091 ( .B1(n3268), .B2(n4609), .A(n3267), .ZN(n3270) );
  INV_X1 U4092 ( .A(n4594), .ZN(n4610) );
  NAND2_X1 U4093 ( .A1(n4650), .A2(n4610), .ZN(n3269) );
  AND2_X1 U4094 ( .A1(n3270), .A2(n3269), .ZN(n4648) );
  MUX2_X1 U4095 ( .A(n4648), .B(n3271), .S(n4619), .Z(n3274) );
  NAND2_X1 U4096 ( .A1(n4598), .A2(n3702), .ZN(n3272) );
  AOI22_X1 U4097 ( .A1(n4601), .A2(n4689), .B1(REG3_REG_2__SCAN_IN), .B2(n4614), .ZN(n3273) );
  OAI211_X1 U4098 ( .C1(n3276), .C2(n3275), .A(n3274), .B(n3273), .ZN(U3288)
         );
  XNOR2_X1 U4099 ( .A(n3278), .B(n3277), .ZN(n3283) );
  AOI22_X1 U4100 ( .A1(n3731), .A2(n2842), .B1(n3732), .B2(n3571), .ZN(n3282)
         );
  NOR2_X1 U4101 ( .A1(n3733), .A2(n3303), .ZN(n3279) );
  AOI211_X1 U4102 ( .C1(n3736), .C2(n3300), .A(n3280), .B(n3279), .ZN(n3281)
         );
  OAI211_X1 U4103 ( .C1(n3283), .C2(n5077), .A(n3282), .B(n3281), .ZN(U3224)
         );
  INV_X1 U4104 ( .A(n3285), .ZN(n3287) );
  NOR2_X1 U4105 ( .A1(n3287), .A2(n3286), .ZN(n3288) );
  XNOR2_X1 U4106 ( .A(n3284), .B(n3288), .ZN(n3293) );
  AOI22_X1 U4107 ( .A1(n3731), .A2(n3390), .B1(n3732), .B2(n3904), .ZN(n3292)
         );
  INV_X1 U4108 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3289) );
  NOR2_X1 U4109 ( .A1(STATE_REG_SCAN_IN), .A2(n3289), .ZN(n4504) );
  NOR2_X1 U4110 ( .A1(n3733), .A2(n3395), .ZN(n3290) );
  AOI211_X1 U4111 ( .C1(n3736), .C2(n3396), .A(n4504), .B(n3290), .ZN(n3291)
         );
  OAI211_X1 U4112 ( .C1(n3293), .C2(n5077), .A(n3292), .B(n3291), .ZN(U3236)
         );
  INV_X1 U4113 ( .A(n3294), .ZN(n3827) );
  NAND2_X1 U4114 ( .A1(n3827), .A2(n3834), .ZN(n3791) );
  XOR2_X1 U4115 ( .A(n3791), .B(n3295), .Z(n3333) );
  INV_X1 U4116 ( .A(n3333), .ZN(n3307) );
  XOR2_X1 U4117 ( .A(n3791), .B(n3296), .Z(n3297) );
  NOR2_X1 U4118 ( .A1(n3297), .A2(n4292), .ZN(n3331) );
  NAND2_X1 U4119 ( .A1(n3331), .A2(n4617), .ZN(n3306) );
  INV_X1 U4120 ( .A(n3298), .ZN(n3310) );
  AOI21_X1 U4121 ( .B1(n3328), .B2(n3310), .A(n3299), .ZN(n3384) );
  INV_X1 U4122 ( .A(n4011), .ZN(n4252) );
  INV_X1 U4123 ( .A(n4009), .ZN(n4253) );
  AOI22_X1 U4124 ( .A1(n4252), .A2(n2842), .B1(n4253), .B2(n3571), .ZN(n3302)
         );
  AOI22_X1 U4125 ( .A1(n4619), .A2(REG2_REG_5__SCAN_IN), .B1(n3300), .B2(n4614), .ZN(n3301) );
  OAI211_X1 U4126 ( .C1(n3303), .C2(n4256), .A(n3302), .B(n3301), .ZN(n3304)
         );
  AOI21_X1 U4127 ( .B1(n3384), .B2(n4601), .A(n3304), .ZN(n3305) );
  OAI211_X1 U4128 ( .C1(n3307), .C2(n4241), .A(n3306), .B(n3305), .ZN(U3285)
         );
  OAI21_X1 U4129 ( .B1(n3308), .B2(n2697), .A(n3317), .ZN(n3309) );
  NAND3_X1 U4130 ( .A1(n3310), .A2(n4399), .A3(n3309), .ZN(n4653) );
  NOR2_X1 U4131 ( .A1(n4653), .A2(n4485), .ZN(n3323) );
  OAI21_X1 U4132 ( .B1(n3313), .B2(n3312), .A(n3311), .ZN(n3314) );
  XNOR2_X1 U4133 ( .A(n3793), .B(n3314), .ZN(n3325) );
  NAND2_X1 U4134 ( .A1(n3239), .A2(n3315), .ZN(n3316) );
  XOR2_X1 U4135 ( .A(n3793), .B(n3316), .Z(n3321) );
  AOI22_X1 U4136 ( .A1(n3390), .A2(n4411), .B1(n3317), .B2(n4588), .ZN(n3318)
         );
  OAI21_X1 U4137 ( .B1(n3319), .B2(n4393), .A(n3318), .ZN(n3320) );
  AOI21_X1 U4138 ( .B1(n3321), .B2(n4609), .A(n3320), .ZN(n3322) );
  OAI21_X1 U4139 ( .B1(n4594), .B2(n3325), .A(n3322), .ZN(n4654) );
  AOI211_X1 U4140 ( .C1(n4614), .C2(n3324), .A(n3323), .B(n4654), .ZN(n3327)
         );
  INV_X1 U4141 ( .A(n3325), .ZN(n4656) );
  AOI22_X1 U4142 ( .A1(n4656), .A2(n4615), .B1(REG2_REG_4__SCAN_IN), .B2(n4619), .ZN(n3326) );
  OAI21_X1 U4143 ( .B1(n3327), .B2(n4619), .A(n3326), .ZN(U3286) );
  AOI22_X1 U4144 ( .A1(n3571), .A2(n4411), .B1(n4588), .B2(n3328), .ZN(n3329)
         );
  OAI21_X1 U4145 ( .B1(n3330), .B2(n4393), .A(n3329), .ZN(n3332) );
  AOI211_X1 U4146 ( .C1(n3333), .C2(n4665), .A(n3332), .B(n3331), .ZN(n3386)
         );
  AOI22_X1 U4147 ( .A1(n3384), .A2(n4651), .B1(REG0_REG_5__SCAN_IN), .B2(n4684), .ZN(n3334) );
  OAI21_X1 U4148 ( .B1(n3386), .B2(n4684), .A(n3334), .ZN(U3477) );
  NAND2_X1 U4149 ( .A1(n4490), .A2(REG2_REG_11__SCAN_IN), .ZN(n3348) );
  MUX2_X1 U4150 ( .A(REG2_REG_11__SCAN_IN), .B(n3335), .S(n4490), .Z(n4545) );
  NAND2_X1 U4151 ( .A1(n4519), .A2(REG2_REG_9__SCAN_IN), .ZN(n3345) );
  MUX2_X1 U4152 ( .A(REG2_REG_9__SCAN_IN), .B(n3336), .S(n4519), .Z(n4524) );
  INV_X1 U4153 ( .A(n4491), .ZN(n3365) );
  NAND2_X1 U4154 ( .A1(n4635), .A2(n3340), .ZN(n3341) );
  INV_X1 U4155 ( .A(n4635), .ZN(n4509) );
  XNOR2_X1 U4156 ( .A(n3340), .B(n4509), .ZN(n4506) );
  NAND2_X1 U4157 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4506), .ZN(n4505) );
  NAND2_X1 U4158 ( .A1(n3341), .A2(n4505), .ZN(n3932) );
  MUX2_X1 U4159 ( .A(REG2_REG_7__SCAN_IN), .B(n3342), .S(n4491), .Z(n3931) );
  NAND2_X1 U4160 ( .A1(n3932), .A2(n3931), .ZN(n3930) );
  NAND2_X1 U4161 ( .A1(n3367), .A2(n3343), .ZN(n3344) );
  INV_X1 U4162 ( .A(n3367), .ZN(n4634) );
  XNOR2_X1 U4163 ( .A(n3343), .B(n4634), .ZN(n4511) );
  NAND2_X1 U4164 ( .A1(REG2_REG_8__SCAN_IN), .A2(n4511), .ZN(n4510) );
  NAND2_X1 U4165 ( .A1(n3344), .A2(n4510), .ZN(n4525) );
  NAND2_X1 U4166 ( .A1(n4524), .A2(n4525), .ZN(n4523) );
  NAND2_X1 U4167 ( .A1(n3345), .A2(n4523), .ZN(n3346) );
  NAND2_X1 U4168 ( .A1(n4632), .A2(n3346), .ZN(n3347) );
  INV_X1 U4169 ( .A(n4632), .ZN(n4540) );
  XNOR2_X1 U4170 ( .A(n3346), .B(n4540), .ZN(n4533) );
  NAND2_X1 U4171 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4533), .ZN(n4532) );
  NAND2_X1 U4172 ( .A1(n3347), .A2(n4532), .ZN(n4546) );
  NAND2_X1 U4173 ( .A1(n4545), .A2(n4546), .ZN(n4544) );
  NAND2_X1 U4174 ( .A1(n3373), .A2(n3349), .ZN(n3350) );
  INV_X1 U4175 ( .A(n3373), .ZN(n4631) );
  NOR2_X1 U4176 ( .A1(n2518), .A2(n4630), .ZN(n4562) );
  OAI22_X1 U4177 ( .A1(n4565), .A2(n4562), .B1(REG2_REG_13__SCAN_IN), .B2(
        n3359), .ZN(n3351) );
  INV_X1 U4178 ( .A(n4489), .ZN(n3377) );
  NOR2_X1 U4179 ( .A1(n3351), .A2(n3377), .ZN(n3416) );
  NAND2_X1 U4180 ( .A1(n3351), .A2(n3377), .ZN(n3352) );
  AOI211_X1 U4181 ( .C1(n4278), .C2(n3353), .A(n3415), .B(n4574), .ZN(n3357)
         );
  NOR2_X1 U4182 ( .A1(n3354), .A2(STATE_REG_SCAN_IN), .ZN(n3589) );
  AOI21_X1 U4183 ( .B1(n4579), .B2(ADDR_REG_14__SCAN_IN), .A(n3589), .ZN(n3355) );
  OAI21_X1 U4184 ( .B1(n3377), .B2(n4585), .A(n3355), .ZN(n3356) );
  NOR2_X1 U4185 ( .A1(n3357), .A2(n3356), .ZN(n3380) );
  NAND2_X1 U4186 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3359), .ZN(n3376) );
  INV_X1 U4187 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4188 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3359), .B1(n4630), .B2(
        n3358), .ZN(n4571) );
  INV_X1 U4189 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4846) );
  INV_X1 U4190 ( .A(n4490), .ZN(n4549) );
  NAND2_X1 U4191 ( .A1(n4519), .A2(REG1_REG_9__SCAN_IN), .ZN(n3370) );
  INV_X1 U4192 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3360) );
  MUX2_X1 U4193 ( .A(n3360), .B(REG1_REG_9__SCAN_IN), .S(n4519), .Z(n3361) );
  INV_X1 U4194 ( .A(n3361), .ZN(n4521) );
  INV_X1 U4195 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4877) );
  XNOR2_X1 U4196 ( .A(n3364), .B(n4635), .ZN(n4502) );
  NOR2_X1 U4197 ( .A1(n4877), .A2(n4502), .ZN(n4501) );
  AOI21_X1 U4198 ( .B1(n4635), .B2(n3364), .A(n4501), .ZN(n3927) );
  NOR2_X1 U4199 ( .A1(n4491), .A2(REG1_REG_7__SCAN_IN), .ZN(n3366) );
  INV_X1 U4200 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4695) );
  OAI22_X1 U4201 ( .A1(n3927), .A2(n3366), .B1(n4695), .B2(n3365), .ZN(n3368)
         );
  NAND2_X1 U4202 ( .A1(n3368), .A2(n3367), .ZN(n3369) );
  XNOR2_X1 U4203 ( .A(n3368), .B(n4634), .ZN(n4516) );
  NAND2_X1 U4204 ( .A1(REG1_REG_8__SCAN_IN), .A2(n4516), .ZN(n4515) );
  NAND2_X1 U4205 ( .A1(n3369), .A2(n4515), .ZN(n4522) );
  NAND2_X1 U4206 ( .A1(n4521), .A2(n4522), .ZN(n4520) );
  NAND2_X1 U4207 ( .A1(n3370), .A2(n4520), .ZN(n3371) );
  NAND2_X1 U4208 ( .A1(n4632), .A2(n3371), .ZN(n3372) );
  XNOR2_X1 U4209 ( .A(n3371), .B(n4540), .ZN(n4537) );
  NAND2_X1 U4210 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4537), .ZN(n4536) );
  NAND2_X1 U4211 ( .A1(n3372), .A2(n4536), .ZN(n4543) );
  MUX2_X1 U4212 ( .A(REG1_REG_11__SCAN_IN), .B(n4846), .S(n4490), .Z(n4542) );
  NAND2_X1 U4213 ( .A1(n4543), .A2(n4542), .ZN(n4541) );
  NAND2_X1 U4214 ( .A1(n3373), .A2(n3374), .ZN(n3375) );
  NAND2_X1 U4215 ( .A1(n4571), .A2(n4570), .ZN(n4569) );
  OAI211_X1 U4216 ( .C1(n3378), .C2(REG1_REG_14__SCAN_IN), .A(n4581), .B(n3421), .ZN(n3379) );
  NAND2_X1 U4217 ( .A1(n3380), .A2(n3379), .ZN(U3254) );
  AOI22_X1 U4218 ( .A1(n2808), .A2(n3381), .B1(REG1_REG_3__SCAN_IN), .B2(n4700), .ZN(n3382) );
  OAI21_X1 U4219 ( .B1(n3383), .B2(n4700), .A(n3382), .ZN(U3521) );
  AOI22_X1 U4220 ( .A1(n3384), .A2(n2808), .B1(REG1_REG_5__SCAN_IN), .B2(n4700), .ZN(n3385) );
  OAI21_X1 U4221 ( .B1(n3386), .B2(n4700), .A(n3385), .ZN(U3523) );
  NAND2_X1 U4222 ( .A1(n3830), .A2(n3833), .ZN(n3800) );
  XNOR2_X1 U4223 ( .A(n3387), .B(n3800), .ZN(n3393) );
  XNOR2_X1 U4224 ( .A(n3388), .B(n3800), .ZN(n4661) );
  NAND2_X1 U4225 ( .A1(n4661), .A2(n4610), .ZN(n3392) );
  OAI22_X1 U4226 ( .A1(n3459), .A2(n4612), .B1(n4288), .B2(n3395), .ZN(n3389)
         );
  AOI21_X1 U4227 ( .B1(n4589), .B2(n3390), .A(n3389), .ZN(n3391) );
  OAI211_X1 U4228 ( .C1(n3393), .C2(n4292), .A(n3392), .B(n3391), .ZN(n4659)
         );
  INV_X1 U4229 ( .A(n4659), .ZN(n3400) );
  OAI21_X1 U4230 ( .B1(n3299), .B2(n3395), .A(n3394), .ZN(n4658) );
  AOI22_X1 U4231 ( .A1(n4619), .A2(REG2_REG_6__SCAN_IN), .B1(n3396), .B2(n4614), .ZN(n3397) );
  OAI21_X1 U4232 ( .B1(n4658), .B2(n4300), .A(n3397), .ZN(n3398) );
  AOI21_X1 U4233 ( .B1(n4661), .B2(n4615), .A(n3398), .ZN(n3399) );
  OAI21_X1 U4234 ( .B1(n3400), .B2(n4619), .A(n3399), .ZN(U3284) );
  INV_X1 U4235 ( .A(n3794), .ZN(n3831) );
  XNOR2_X1 U4236 ( .A(n3401), .B(n3831), .ZN(n3402) );
  NAND2_X1 U4237 ( .A1(n3402), .A2(n4609), .ZN(n3404) );
  AOI22_X1 U4238 ( .A1(n3903), .A2(n4411), .B1(n4588), .B2(n3406), .ZN(n3403)
         );
  OAI211_X1 U4239 ( .C1(n3405), .C2(n4393), .A(n3404), .B(n3403), .ZN(n4663)
         );
  INV_X1 U4240 ( .A(n4663), .ZN(n3414) );
  AOI21_X1 U4241 ( .B1(n3394), .B2(n3406), .A(n4678), .ZN(n3407) );
  AND2_X1 U4242 ( .A1(n3407), .A2(n3464), .ZN(n4664) );
  INV_X1 U4243 ( .A(n4197), .ZN(n3410) );
  INV_X1 U4244 ( .A(n3574), .ZN(n3408) );
  OAI22_X1 U4245 ( .A1(n4617), .A2(n3342), .B1(n3408), .B2(n4276), .ZN(n3409)
         );
  AOI21_X1 U4246 ( .B1(n4664), .B2(n3410), .A(n3409), .ZN(n3413) );
  XOR2_X1 U4247 ( .A(n3411), .B(n3794), .Z(n4666) );
  NAND2_X1 U4248 ( .A1(n4666), .A2(n4302), .ZN(n3412) );
  OAI211_X1 U4249 ( .C1(n3414), .C2(n4619), .A(n3413), .B(n3412), .ZN(U3283)
         );
  NAND2_X1 U4250 ( .A1(n4488), .A2(REG2_REG_15__SCAN_IN), .ZN(n3944) );
  OAI21_X1 U4251 ( .B1(n4488), .B2(REG2_REG_15__SCAN_IN), .A(n3944), .ZN(n3418) );
  INV_X1 U4252 ( .A(n3945), .ZN(n3417) );
  AOI211_X1 U4253 ( .C1(n3419), .C2(n3418), .A(n3417), .B(n4574), .ZN(n3429)
         );
  INV_X1 U4254 ( .A(n4488), .ZN(n3938) );
  NAND2_X1 U4255 ( .A1(n4489), .A2(n3420), .ZN(n3422) );
  INV_X1 U4256 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4891) );
  NOR2_X1 U4257 ( .A1(n3938), .A2(n4891), .ZN(n3423) );
  AOI21_X1 U4258 ( .B1(n4891), .B2(n3938), .A(n3423), .ZN(n3424) );
  NAND2_X1 U4259 ( .A1(n3424), .A2(n3425), .ZN(n3937) );
  OAI211_X1 U4260 ( .C1(n3425), .C2(n3424), .A(n4581), .B(n3937), .ZN(n3427)
         );
  AND2_X1 U4261 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n3735) );
  AOI21_X1 U4262 ( .B1(n4579), .B2(ADDR_REG_15__SCAN_IN), .A(n3735), .ZN(n3426) );
  OAI211_X1 U4263 ( .C1(n4585), .C2(n3938), .A(n3427), .B(n3426), .ZN(n3428)
         );
  OR2_X1 U4264 ( .A1(n3429), .A2(n3428), .ZN(U3255) );
  INV_X1 U4265 ( .A(n3431), .ZN(n3433) );
  NOR2_X1 U4266 ( .A1(n3433), .A2(n3432), .ZN(n3434) );
  XNOR2_X1 U4267 ( .A(n3430), .B(n3434), .ZN(n3438) );
  NAND2_X1 U4268 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4512) );
  OAI21_X1 U4269 ( .B1(n3733), .B2(n3465), .A(n4512), .ZN(n3436) );
  OAI22_X1 U4270 ( .A1(n5082), .A2(n5080), .B1(n5081), .B2(n3459), .ZN(n3435)
         );
  AOI211_X1 U4271 ( .C1(n3467), .C2(n3736), .A(n3436), .B(n3435), .ZN(n3437)
         );
  OAI21_X1 U4272 ( .B1(n3438), .B2(n5077), .A(n3437), .ZN(U3218) );
  NAND2_X1 U4273 ( .A1(n3845), .A2(n3846), .ZN(n3790) );
  INV_X1 U4274 ( .A(n3790), .ZN(n3439) );
  XNOR2_X1 U4275 ( .A(n3440), .B(n3439), .ZN(n3441) );
  NAND2_X1 U4276 ( .A1(n3441), .A2(n4609), .ZN(n3494) );
  XNOR2_X1 U4277 ( .A(n3442), .B(n3790), .ZN(n3489) );
  INV_X1 U4278 ( .A(n4668), .ZN(n3444) );
  AOI21_X1 U4279 ( .B1(n3490), .B2(n3444), .A(n3443), .ZN(n3499) );
  INV_X1 U4280 ( .A(n3499), .ZN(n3451) );
  OAI22_X1 U4281 ( .A1(n3445), .A2(n4276), .B1(n3336), .B2(n4617), .ZN(n3449)
         );
  OAI22_X1 U4282 ( .A1(n3447), .A2(n4011), .B1(n3446), .B2(n4009), .ZN(n3448)
         );
  AOI211_X1 U4283 ( .C1(n3995), .C2(n3490), .A(n3449), .B(n3448), .ZN(n3450)
         );
  OAI21_X1 U4284 ( .B1(n3451), .B2(n4300), .A(n3450), .ZN(n3452) );
  AOI21_X1 U4285 ( .B1(n3489), .B2(n4302), .A(n3452), .ZN(n3453) );
  OAI21_X1 U4286 ( .B1(n3494), .B2(n4619), .A(n3453), .ZN(U3281) );
  INV_X1 U4287 ( .A(n3840), .ZN(n3455) );
  NAND2_X1 U4288 ( .A1(n3455), .A2(n3844), .ZN(n3792) );
  XNOR2_X1 U4289 ( .A(n3454), .B(n3792), .ZN(n3463) );
  XNOR2_X1 U4290 ( .A(n3456), .B(n3792), .ZN(n3461) );
  AOI22_X1 U4291 ( .A1(n3902), .A2(n4411), .B1(n3457), .B2(n4588), .ZN(n3458)
         );
  OAI21_X1 U4292 ( .B1(n3459), .B2(n4393), .A(n3458), .ZN(n3460) );
  AOI21_X1 U4293 ( .B1(n3461), .B2(n4609), .A(n3460), .ZN(n3462) );
  OAI21_X1 U4294 ( .B1(n3463), .B2(n4594), .A(n3462), .ZN(n4670) );
  INV_X1 U4295 ( .A(n4670), .ZN(n3473) );
  INV_X1 U4296 ( .A(n3463), .ZN(n4672) );
  INV_X1 U4297 ( .A(n3464), .ZN(n3466) );
  NOR2_X1 U4298 ( .A1(n3466), .A2(n3465), .ZN(n4669) );
  NOR3_X1 U4299 ( .A1(n4669), .A2(n4668), .A3(n4300), .ZN(n3471) );
  INV_X1 U4300 ( .A(n3467), .ZN(n3468) );
  OAI22_X1 U4301 ( .A1(n4617), .A2(n3469), .B1(n3468), .B2(n4276), .ZN(n3470)
         );
  AOI211_X1 U4302 ( .C1(n4672), .C2(n4615), .A(n3471), .B(n3470), .ZN(n3472)
         );
  OAI21_X1 U4303 ( .B1(n3473), .B2(n4619), .A(n3472), .ZN(U3282) );
  NAND2_X1 U4304 ( .A1(n3850), .A2(n3851), .ZN(n3786) );
  XNOR2_X1 U4305 ( .A(n3474), .B(n3786), .ZN(n3481) );
  XOR2_X1 U4306 ( .A(n3786), .B(n3475), .Z(n3479) );
  AOI22_X1 U4307 ( .A1(n4413), .A2(n4411), .B1(n4588), .B2(n3476), .ZN(n3477)
         );
  OAI21_X1 U4308 ( .B1(n5082), .B2(n4393), .A(n3477), .ZN(n3478) );
  AOI21_X1 U4309 ( .B1(n3479), .B2(n4609), .A(n3478), .ZN(n3480) );
  OAI21_X1 U4310 ( .B1(n4594), .B2(n3481), .A(n3480), .ZN(n4675) );
  INV_X1 U4311 ( .A(n4675), .ZN(n3488) );
  INV_X1 U4312 ( .A(n3481), .ZN(n4677) );
  NOR2_X1 U4313 ( .A1(n3443), .A2(n5086), .ZN(n4674) );
  INV_X1 U4314 ( .A(n3482), .ZN(n4673) );
  NOR3_X1 U4315 ( .A1(n4674), .A2(n4673), .A3(n4300), .ZN(n3486) );
  INV_X1 U4316 ( .A(n5083), .ZN(n3483) );
  OAI22_X1 U4317 ( .A1(n4617), .A2(n3484), .B1(n3483), .B2(n4276), .ZN(n3485)
         );
  AOI211_X1 U4318 ( .C1(n4677), .C2(n4615), .A(n3486), .B(n3485), .ZN(n3487)
         );
  OAI21_X1 U4319 ( .B1(n3488), .B2(n4619), .A(n3487), .ZN(U3280) );
  NAND2_X1 U4320 ( .A1(n3489), .A2(n4665), .ZN(n3493) );
  AOI22_X1 U4321 ( .A1(n3901), .A2(n4411), .B1(n4588), .B2(n3490), .ZN(n3492)
         );
  NAND2_X1 U4322 ( .A1(n3903), .A2(n4589), .ZN(n3491) );
  NAND4_X1 U4323 ( .A1(n3494), .A2(n3493), .A3(n3492), .A4(n3491), .ZN(n3497)
         );
  INV_X2 U4324 ( .A(n4684), .ZN(n4685) );
  MUX2_X1 U4325 ( .A(REG0_REG_9__SCAN_IN), .B(n3497), .S(n4685), .Z(n3495) );
  AOI21_X1 U4326 ( .B1(n3499), .B2(n4651), .A(n3495), .ZN(n3496) );
  INV_X1 U4327 ( .A(n3496), .ZN(U3485) );
  MUX2_X1 U4328 ( .A(REG1_REG_9__SCAN_IN), .B(n3497), .S(n4702), .Z(n3498) );
  AOI21_X1 U4329 ( .B1(n2808), .B2(n3499), .A(n3498), .ZN(n3500) );
  INV_X1 U4330 ( .A(n3500), .ZN(U3527) );
  XOR2_X1 U4331 ( .A(n3503), .B(n3502), .Z(n3504) );
  XNOR2_X1 U4332 ( .A(n3501), .B(n3504), .ZN(n3508) );
  AOI22_X1 U4333 ( .A1(n3731), .A2(n3901), .B1(n3732), .B2(n4290), .ZN(n3507)
         );
  NOR2_X1 U4334 ( .A1(STATE_REG_SCAN_IN), .A2(n4965), .ZN(n4551) );
  NOR2_X1 U4335 ( .A1(n3733), .A2(n3532), .ZN(n3505) );
  AOI211_X1 U4336 ( .C1(n3736), .C2(n3533), .A(n4551), .B(n3505), .ZN(n3506)
         );
  OAI211_X1 U4337 ( .C1(n3508), .C2(n5077), .A(n3507), .B(n3506), .ZN(U3233)
         );
  INV_X1 U4338 ( .A(n3510), .ZN(n3511) );
  OR2_X1 U4339 ( .A1(n3509), .A2(n3511), .ZN(n3513) );
  NAND2_X1 U4340 ( .A1(n3513), .A2(n3512), .ZN(n4286) );
  NAND2_X1 U4341 ( .A1(n4285), .A2(n4283), .ZN(n3787) );
  XNOR2_X1 U4342 ( .A(n4286), .B(n3787), .ZN(n3514) );
  NAND2_X1 U4343 ( .A1(n3514), .A2(n4609), .ZN(n4415) );
  XNOR2_X1 U4344 ( .A(n3515), .B(n3787), .ZN(n4409) );
  AND2_X1 U4345 ( .A1(n3531), .A2(n4410), .ZN(n3516) );
  NOR2_X1 U4346 ( .A1(n4297), .A2(n3516), .ZN(n4476) );
  NAND2_X1 U4347 ( .A1(n4476), .A2(n4601), .ZN(n3522) );
  INV_X1 U4348 ( .A(n3544), .ZN(n3517) );
  OAI22_X1 U4349 ( .A1(n4617), .A2(n3518), .B1(n3517), .B2(n4276), .ZN(n3519)
         );
  AOI21_X1 U4350 ( .B1(n4410), .B2(n3995), .A(n3519), .ZN(n3521) );
  AOI22_X1 U4351 ( .A1(n4252), .A2(n4413), .B1(n4253), .B2(n4412), .ZN(n3520)
         );
  NAND3_X1 U4352 ( .A1(n3522), .A2(n3521), .A3(n3520), .ZN(n3523) );
  AOI21_X1 U4353 ( .B1(n4409), .B2(n4302), .A(n3523), .ZN(n3524) );
  OAI21_X1 U4354 ( .B1(n4619), .B2(n4415), .A(n3524), .ZN(U3278) );
  XNOR2_X1 U4355 ( .A(n3509), .B(n3795), .ZN(n3530) );
  XNOR2_X1 U4356 ( .A(n3525), .B(n3795), .ZN(n4682) );
  NAND2_X1 U4357 ( .A1(n4682), .A2(n4610), .ZN(n3529) );
  OAI22_X1 U4358 ( .A1(n3526), .A2(n4612), .B1(n4288), .B2(n3532), .ZN(n3527)
         );
  AOI21_X1 U4359 ( .B1(n4589), .B2(n3901), .A(n3527), .ZN(n3528) );
  OAI211_X1 U4360 ( .C1(n4292), .C2(n3530), .A(n3529), .B(n3528), .ZN(n4680)
         );
  INV_X1 U4361 ( .A(n4680), .ZN(n3537) );
  OAI21_X1 U4362 ( .B1(n4673), .B2(n3532), .A(n3531), .ZN(n4679) );
  AOI22_X1 U4363 ( .A1(n4619), .A2(REG2_REG_11__SCAN_IN), .B1(n3533), .B2(
        n4614), .ZN(n3534) );
  OAI21_X1 U4364 ( .B1(n4679), .B2(n4300), .A(n3534), .ZN(n3535) );
  AOI21_X1 U4365 ( .B1(n4682), .B2(n4615), .A(n3535), .ZN(n3536) );
  OAI21_X1 U4366 ( .B1(n3537), .B2(n4619), .A(n3536), .ZN(U3279) );
  NOR2_X1 U4367 ( .A1(n2272), .A2(n3539), .ZN(n3540) );
  XNOR2_X1 U4368 ( .A(n3538), .B(n3540), .ZN(n3546) );
  NAND2_X1 U4369 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4555) );
  OAI21_X1 U4370 ( .B1(n3733), .B2(n3541), .A(n4555), .ZN(n3543) );
  OAI22_X1 U4371 ( .A1(n5079), .A2(n5081), .B1(n5080), .B2(n3591), .ZN(n3542)
         );
  AOI211_X1 U4372 ( .C1(n3544), .C2(n3736), .A(n3543), .B(n3542), .ZN(n3545)
         );
  OAI21_X1 U4373 ( .B1(n3546), .B2(n5077), .A(n3545), .ZN(U3221) );
  XOR2_X1 U4374 ( .A(n3547), .B(n3548), .Z(n3554) );
  AOI22_X1 U4375 ( .A1(n3731), .A2(n3903), .B1(n3732), .B2(n3901), .ZN(n3553)
         );
  AND2_X1 U4376 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4530) );
  NOR2_X1 U4377 ( .A1(n3733), .A2(n3549), .ZN(n3550) );
  AOI211_X1 U4378 ( .C1(n3736), .C2(n3551), .A(n4530), .B(n3550), .ZN(n3552)
         );
  OAI211_X1 U4379 ( .C1(n3554), .C2(n5077), .A(n3553), .B(n3552), .ZN(U3228)
         );
  XOR2_X1 U4380 ( .A(n3557), .B(n3556), .Z(n3558) );
  XNOR2_X1 U4381 ( .A(n3555), .B(n3558), .ZN(n3562) );
  AOI22_X1 U4382 ( .A1(n3731), .A2(n4290), .B1(n3732), .B2(n4251), .ZN(n3561)
         );
  AND2_X1 U4383 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n4568) );
  NOR2_X1 U4384 ( .A1(n3733), .A2(n4296), .ZN(n3559) );
  AOI211_X1 U4385 ( .C1(n3736), .C2(n4298), .A(n4568), .B(n3559), .ZN(n3560)
         );
  OAI211_X1 U4386 ( .C1(n3562), .C2(n5077), .A(n3561), .B(n3560), .ZN(U3231)
         );
  INV_X1 U4387 ( .A(IR_REG_30__SCAN_IN), .ZN(n3564) );
  NAND3_X1 U4388 ( .A1(n3564), .A2(STATE_REG_SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n3566) );
  INV_X1 U4389 ( .A(DATAI_31_), .ZN(n3565) );
  OAI22_X1 U4390 ( .A1(n3563), .A2(n3566), .B1(STATE_REG_SCAN_IN), .B2(n3565), 
        .ZN(U3321) );
  AOI21_X1 U4391 ( .B1(n3567), .B2(n3568), .A(n5077), .ZN(n3570) );
  NAND2_X1 U4392 ( .A1(n3570), .A2(n3569), .ZN(n3577) );
  AOI22_X1 U4393 ( .A1(n3731), .A2(n3571), .B1(n3732), .B2(n3903), .ZN(n3576)
         );
  NOR2_X1 U4394 ( .A1(STATE_REG_SCAN_IN), .A2(n4939), .ZN(n3929) );
  NOR2_X1 U4395 ( .A1(n3733), .A2(n3572), .ZN(n3573) );
  AOI211_X1 U4396 ( .C1(n3736), .C2(n3574), .A(n3929), .B(n3573), .ZN(n3575)
         );
  NAND3_X1 U4397 ( .A1(n3577), .A2(n3576), .A3(n3575), .ZN(U3210) );
  XNOR2_X1 U4398 ( .A(n3579), .B(n3578), .ZN(n3584) );
  OAI22_X1 U4399 ( .A1(n3733), .A2(n4028), .B1(STATE_REG_SCAN_IN), .B2(n3580), 
        .ZN(n3582) );
  OAI22_X1 U4400 ( .A1(n4315), .A2(n5080), .B1(n3643), .B2(n5081), .ZN(n3581)
         );
  AOI211_X1 U4401 ( .C1(n4024), .C2(n3736), .A(n3582), .B(n3581), .ZN(n3583)
         );
  OAI21_X1 U4402 ( .B1(n3584), .B2(n5077), .A(n3583), .ZN(U3211) );
  NAND2_X1 U4403 ( .A1(n3587), .A2(n3586), .ZN(n3588) );
  XNOR2_X1 U4404 ( .A(n3585), .B(n3588), .ZN(n3595) );
  INV_X1 U4405 ( .A(n3589), .ZN(n3590) );
  OAI21_X1 U4406 ( .B1(n3733), .B2(n4274), .A(n3590), .ZN(n3593) );
  OAI22_X1 U4407 ( .A1(n3591), .A2(n5081), .B1(n5080), .B2(n4382), .ZN(n3592)
         );
  AOI211_X1 U4408 ( .C1(n4275), .C2(n3736), .A(n3593), .B(n3592), .ZN(n3594)
         );
  OAI21_X1 U4409 ( .B1(n3595), .B2(n5077), .A(n3594), .ZN(U3212) );
  INV_X1 U4410 ( .A(n3596), .ZN(n3598) );
  NOR2_X1 U4411 ( .A1(n3598), .A2(n3597), .ZN(n3599) );
  NAND2_X1 U4412 ( .A1(n3599), .A2(n3699), .ZN(n3611) );
  NAND2_X1 U4413 ( .A1(n3601), .A2(n3600), .ZN(n3675) );
  NAND2_X1 U4414 ( .A1(n3675), .A2(n3676), .ZN(n3674) );
  NAND2_X1 U4415 ( .A1(n3674), .A2(n3678), .ZN(n3631) );
  AOI21_X1 U4416 ( .B1(n3687), .B2(n3605), .A(n3604), .ZN(n3610) );
  OAI22_X1 U4417 ( .A1(n3733), .A2(n4098), .B1(STATE_REG_SCAN_IN), .B2(n3606), 
        .ZN(n3608) );
  OAI22_X1 U4418 ( .A1(n4093), .A2(n5080), .B1(n3632), .B2(n5081), .ZN(n3607)
         );
  AOI211_X1 U4419 ( .C1(n4100), .C2(n3736), .A(n3608), .B(n3607), .ZN(n3609)
         );
  OAI21_X1 U4420 ( .B1(n3611), .B2(n3610), .A(n3609), .ZN(U3213) );
  OAI21_X1 U4421 ( .B1(n3613), .B2(n3612), .A(n3219), .ZN(n3614) );
  NAND2_X1 U4422 ( .A1(n3614), .A2(n3699), .ZN(n3621) );
  AOI22_X1 U4423 ( .A1(n3731), .A2(n3907), .B1(n3732), .B2(n2842), .ZN(n3620)
         );
  NOR2_X1 U4424 ( .A1(n3733), .A2(n3615), .ZN(n3616) );
  AOI211_X1 U4425 ( .C1(n3736), .C2(n3618), .A(n3617), .B(n3616), .ZN(n3619)
         );
  NAND3_X1 U4426 ( .A1(n3621), .A2(n3620), .A3(n3619), .ZN(U3215) );
  XOR2_X1 U4427 ( .A(n3623), .B(n3622), .Z(n3627) );
  AOI22_X1 U4428 ( .A1(n3731), .A2(n4372), .B1(n3732), .B2(n4131), .ZN(n3626)
         );
  INV_X1 U4429 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4905) );
  NOR2_X1 U4430 ( .A1(n4905), .A2(STATE_REG_SCAN_IN), .ZN(n3979) );
  NOR2_X1 U4431 ( .A1(n3733), .A2(n4167), .ZN(n3624) );
  AOI211_X1 U4432 ( .C1(n3736), .C2(n2358), .A(n3979), .B(n3624), .ZN(n3625)
         );
  OAI211_X1 U4433 ( .C1(n3627), .C2(n5077), .A(n3626), .B(n3625), .ZN(U3216)
         );
  XNOR2_X1 U4434 ( .A(n3629), .B(n3628), .ZN(n3630) );
  XNOR2_X1 U4435 ( .A(n3631), .B(n3630), .ZN(n3636) );
  OAI22_X1 U4436 ( .A1(n3733), .A2(n4135), .B1(STATE_REG_SCAN_IN), .B2(n4790), 
        .ZN(n3634) );
  OAI22_X1 U4437 ( .A1(n4355), .A2(n5081), .B1(n5080), .B2(n3632), .ZN(n3633)
         );
  AOI211_X1 U4438 ( .C1(n4132), .C2(n3736), .A(n3634), .B(n3633), .ZN(n3635)
         );
  OAI21_X1 U4439 ( .B1(n3636), .B2(n5077), .A(n3635), .ZN(U3220) );
  NAND2_X1 U4440 ( .A1(n3638), .A2(n3637), .ZN(n3640) );
  XOR2_X1 U4441 ( .A(n3640), .B(n3639), .Z(n3647) );
  INV_X1 U4442 ( .A(n3641), .ZN(n4066) );
  INV_X1 U4443 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3642) );
  OAI22_X1 U4444 ( .A1(n3733), .A2(n4065), .B1(STATE_REG_SCAN_IN), .B2(n3642), 
        .ZN(n3645) );
  OAI22_X1 U4445 ( .A1(n3643), .A2(n5080), .B1(n4093), .B2(n5081), .ZN(n3644)
         );
  AOI211_X1 U4446 ( .C1(n4066), .C2(n3736), .A(n3645), .B(n3644), .ZN(n3646)
         );
  OAI21_X1 U4447 ( .B1(n3647), .B2(n5077), .A(n3646), .ZN(U3222) );
  INV_X1 U4448 ( .A(n3649), .ZN(n3728) );
  NAND2_X1 U4449 ( .A1(n3648), .A2(n3728), .ZN(n3727) );
  NAND2_X1 U4450 ( .A1(n3727), .A2(n3650), .ZN(n3651) );
  XOR2_X1 U4451 ( .A(n3652), .B(n3651), .Z(n3656) );
  AOI22_X1 U4452 ( .A1(n3731), .A2(n4266), .B1(n3732), .B2(n4380), .ZN(n3655)
         );
  INV_X1 U4453 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4984) );
  NOR2_X1 U4454 ( .A1(STATE_REG_SCAN_IN), .A2(n4984), .ZN(n3941) );
  NOR2_X1 U4455 ( .A1(n3733), .A2(n4234), .ZN(n3653) );
  AOI211_X1 U4456 ( .C1(n3736), .C2(n4231), .A(n3941), .B(n3653), .ZN(n3654)
         );
  OAI211_X1 U4457 ( .C1(n3656), .C2(n5077), .A(n3655), .B(n3654), .ZN(U3223)
         );
  XNOR2_X1 U4458 ( .A(n3659), .B(n3658), .ZN(n3660) );
  XNOR2_X1 U4459 ( .A(n3657), .B(n3660), .ZN(n3664) );
  AOI22_X1 U4460 ( .A1(n3731), .A2(n4390), .B1(n3732), .B2(n4372), .ZN(n3663)
         );
  AND2_X1 U4461 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n3965) );
  NOR2_X1 U4462 ( .A1(n3733), .A2(n4215), .ZN(n3661) );
  AOI211_X1 U4463 ( .C1(n3736), .C2(n4212), .A(n3965), .B(n3661), .ZN(n3662)
         );
  OAI211_X1 U4464 ( .C1(n3664), .C2(n5077), .A(n3663), .B(n3662), .ZN(U3225)
         );
  NAND2_X1 U4465 ( .A1(n3665), .A2(n3666), .ZN(n3667) );
  XOR2_X1 U4466 ( .A(n3668), .B(n3667), .Z(n3673) );
  INV_X1 U4467 ( .A(n3669), .ZN(n4077) );
  INV_X1 U4468 ( .A(REG3_REG_24__SCAN_IN), .ZN(n5047) );
  OAI22_X1 U4469 ( .A1(n3733), .A2(n4080), .B1(STATE_REG_SCAN_IN), .B2(n5047), 
        .ZN(n3671) );
  OAI22_X1 U4470 ( .A1(n4338), .A2(n5080), .B1(n4108), .B2(n5081), .ZN(n3670)
         );
  AOI211_X1 U4471 ( .C1(n4077), .C2(n3736), .A(n3671), .B(n3670), .ZN(n3672)
         );
  OAI21_X1 U4472 ( .B1(n3673), .B2(n5077), .A(n3672), .ZN(U3226) );
  INV_X1 U4473 ( .A(n3674), .ZN(n3679) );
  AOI21_X1 U4474 ( .B1(n3678), .B2(n3676), .A(n3675), .ZN(n3677) );
  AOI21_X1 U4475 ( .B1(n3679), .B2(n3678), .A(n3677), .ZN(n3684) );
  AOI22_X1 U4476 ( .A1(n3731), .A2(n4189), .B1(n3732), .B2(n4143), .ZN(n3683)
         );
  INV_X1 U4477 ( .A(REG3_REG_20__SCAN_IN), .ZN(n5045) );
  OAI22_X1 U4478 ( .A1(n3733), .A2(n3680), .B1(STATE_REG_SCAN_IN), .B2(n5045), 
        .ZN(n3681) );
  AOI21_X1 U4479 ( .B1(n4152), .B2(n3736), .A(n3681), .ZN(n3682) );
  OAI211_X1 U4480 ( .C1(n3684), .C2(n5077), .A(n3683), .B(n3682), .ZN(U3230)
         );
  NAND2_X1 U4481 ( .A1(n3686), .A2(n3685), .ZN(n3688) );
  OAI22_X1 U4482 ( .A1(n3733), .A2(n4112), .B1(STATE_REG_SCAN_IN), .B2(n3690), 
        .ZN(n3693) );
  OAI22_X1 U4483 ( .A1(n4108), .A2(n5080), .B1(n5081), .B2(n3691), .ZN(n3692)
         );
  AOI211_X1 U4484 ( .C1(n4115), .C2(n3736), .A(n3693), .B(n3692), .ZN(n3694)
         );
  OAI21_X1 U4485 ( .B1(n3695), .B2(n5077), .A(n3694), .ZN(U3232) );
  OAI21_X1 U4486 ( .B1(n3696), .B2(n3697), .A(n3698), .ZN(n3700) );
  NAND2_X1 U4487 ( .A1(n3700), .A2(n3699), .ZN(n3706) );
  AOI22_X1 U4488 ( .A1(n3703), .A2(n3702), .B1(REG3_REG_2__SCAN_IN), .B2(n3701), .ZN(n3705) );
  AOI22_X1 U4489 ( .A1(n3732), .A2(n3905), .B1(n3731), .B2(n2812), .ZN(n3704)
         );
  NAND3_X1 U4490 ( .A1(n3706), .A2(n3705), .A3(n3704), .ZN(U3234) );
  INV_X1 U4491 ( .A(n3708), .ZN(n3710) );
  NOR2_X1 U4492 ( .A1(n3710), .A2(n3709), .ZN(n3711) );
  XNOR2_X1 U4493 ( .A(n3707), .B(n3711), .ZN(n3716) );
  AOI22_X1 U4494 ( .A1(n3732), .A2(n4189), .B1(n3731), .B2(n4380), .ZN(n3715)
         );
  NOR2_X1 U4495 ( .A1(n3712), .A2(STATE_REG_SCAN_IN), .ZN(n4578) );
  NOR2_X1 U4496 ( .A1(n3733), .A2(n4194), .ZN(n3713) );
  AOI211_X1 U4497 ( .C1(n3736), .C2(n4195), .A(n4578), .B(n3713), .ZN(n3714)
         );
  OAI211_X1 U4498 ( .C1(n3716), .C2(n5077), .A(n3715), .B(n3714), .ZN(U3235)
         );
  INV_X1 U4499 ( .A(n3718), .ZN(n3720) );
  NOR2_X1 U4500 ( .A1(n3720), .A2(n3719), .ZN(n3721) );
  XNOR2_X1 U4501 ( .A(n3717), .B(n3721), .ZN(n3726) );
  INV_X1 U4502 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3722) );
  OAI22_X1 U4503 ( .A1(n3733), .A2(n4048), .B1(STATE_REG_SCAN_IN), .B2(n3722), 
        .ZN(n3724) );
  OAI22_X1 U4504 ( .A1(n4325), .A2(n5080), .B1(n4338), .B2(n5081), .ZN(n3723)
         );
  AOI211_X1 U4505 ( .C1(n4045), .C2(n3736), .A(n3724), .B(n3723), .ZN(n3725)
         );
  OAI21_X1 U4506 ( .B1(n3726), .B2(n5077), .A(n3725), .ZN(U3237) );
  INV_X1 U4507 ( .A(n3727), .ZN(n3730) );
  AOI21_X1 U4508 ( .B1(n3648), .B2(n3650), .A(n3728), .ZN(n3729) );
  AOI21_X1 U4509 ( .B1(n3730), .B2(n3650), .A(n3729), .ZN(n3739) );
  AOI22_X1 U4510 ( .A1(n3732), .A2(n4390), .B1(n3731), .B2(n4251), .ZN(n3738)
         );
  NOR2_X1 U4511 ( .A1(n3733), .A2(n4257), .ZN(n3734) );
  AOI211_X1 U4512 ( .C1(n3736), .C2(n2350), .A(n3735), .B(n3734), .ZN(n3737)
         );
  OAI211_X1 U4513 ( .C1(n3739), .C2(n5077), .A(n3738), .B(n3737), .ZN(U3238)
         );
  NAND2_X1 U4514 ( .A1(n2248), .A2(REG1_REG_31__SCAN_IN), .ZN(n3745) );
  NAND2_X1 U4515 ( .A1(n3741), .A2(REG0_REG_31__SCAN_IN), .ZN(n3744) );
  INV_X1 U4516 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3989) );
  OR2_X1 U4517 ( .A1(n3742), .A2(n3989), .ZN(n3743) );
  NAND2_X1 U4518 ( .A1(n3748), .A2(n3747), .ZN(n3843) );
  AND2_X1 U4519 ( .A1(n3843), .A2(n3750), .ZN(n3857) );
  INV_X1 U4520 ( .A(n3857), .ZN(n3752) );
  INV_X1 U4521 ( .A(n3749), .ZN(n3859) );
  AOI21_X1 U4522 ( .B1(n3751), .B2(n3750), .A(n3857), .ZN(n3854) );
  INV_X1 U4523 ( .A(n3753), .ZN(n3754) );
  OAI21_X1 U4524 ( .B1(n3755), .B2(n3754), .A(n3862), .ZN(n3756) );
  NAND2_X1 U4525 ( .A1(n3756), .A2(n3866), .ZN(n3759) );
  INV_X1 U4526 ( .A(n3810), .ZN(n3757) );
  NOR2_X1 U4527 ( .A1(n3758), .A2(n3757), .ZN(n3870) );
  OAI221_X1 U4528 ( .B1(n3760), .B2(n3869), .C1(n3760), .C2(n3759), .A(n3870), 
        .ZN(n3765) );
  OR2_X1 U4529 ( .A1(n3762), .A2(n3761), .ZN(n3770) );
  NAND2_X1 U4530 ( .A1(n3775), .A2(n4309), .ZN(n3763) );
  INV_X1 U4531 ( .A(n3987), .ZN(n3898) );
  NAND2_X1 U4532 ( .A1(n2602), .A2(DATAI_31_), .ZN(n3985) );
  NAND2_X1 U4533 ( .A1(n3898), .A2(n3985), .ZN(n3880) );
  NAND2_X1 U4534 ( .A1(n3763), .A2(n3880), .ZN(n3785) );
  INV_X1 U4535 ( .A(n3785), .ZN(n3764) );
  OAI21_X1 U4536 ( .B1(n3900), .B2(n3992), .A(n3764), .ZN(n3769) );
  AOI211_X1 U4537 ( .C1(n4035), .C2(n3765), .A(n3770), .B(n3769), .ZN(n3773)
         );
  INV_X1 U4538 ( .A(n3872), .ZN(n3772) );
  NAND2_X1 U4539 ( .A1(n3900), .A2(n3992), .ZN(n3766) );
  AND2_X1 U4540 ( .A1(n3767), .A2(n3766), .ZN(n3875) );
  NAND3_X1 U4541 ( .A1(n4018), .A2(n3875), .A3(n3768), .ZN(n3771) );
  AOI21_X1 U4542 ( .B1(n3875), .B2(n3770), .A(n3769), .ZN(n3882) );
  AOI22_X1 U4543 ( .A1(n3773), .A2(n3772), .B1(n3771), .B2(n3882), .ZN(n3774)
         );
  AOI21_X1 U4544 ( .B1(n3987), .B2(n4309), .A(n3774), .ZN(n3779) );
  INV_X1 U4545 ( .A(n3775), .ZN(n3899) );
  INV_X1 U4546 ( .A(n4309), .ZN(n3776) );
  NAND2_X1 U4547 ( .A1(n3899), .A2(n3776), .ZN(n3781) );
  AOI21_X1 U4548 ( .B1(n3781), .B2(n3898), .A(n3985), .ZN(n3778) );
  NOR3_X1 U4549 ( .A1(n3779), .A2(n3778), .A3(n3777), .ZN(n3887) );
  NAND2_X1 U4550 ( .A1(n4036), .A2(n3780), .ZN(n4055) );
  OAI21_X1 U4551 ( .B1(n3985), .B2(n3898), .A(n3781), .ZN(n3881) );
  NOR3_X1 U4552 ( .A1(n4055), .A2(n4483), .A3(n3881), .ZN(n3789) );
  INV_X1 U4553 ( .A(n3782), .ZN(n3784) );
  NOR4_X1 U4554 ( .A1(n4294), .A2(n3787), .A3(n3786), .A4(n3785), .ZN(n3788)
         );
  NAND3_X1 U4555 ( .A1(n2678), .A2(n3789), .A3(n3788), .ZN(n3807) );
  XNOR2_X1 U4556 ( .A(n4313), .B(n4048), .ZN(n4042) );
  NOR4_X1 U4557 ( .A1(n3792), .A2(n3791), .A3(n4263), .A4(n3790), .ZN(n3804)
         );
  NOR4_X1 U4558 ( .A1(n3796), .A2(n3795), .A3(n3794), .A4(n3793), .ZN(n3803)
         );
  NAND2_X1 U4559 ( .A1(n2821), .A2(n4607), .ZN(n3819) );
  NAND2_X1 U4560 ( .A1(n3798), .A2(n3819), .ZN(n4639) );
  NOR4_X1 U4561 ( .A1(n3799), .A2(n4593), .A3(n4639), .A4(n4228), .ZN(n3802)
         );
  INV_X1 U4562 ( .A(n4087), .ZN(n3865) );
  NAND2_X1 U4563 ( .A1(n3865), .A2(n4086), .ZN(n4127) );
  NOR4_X1 U4564 ( .A1(n4117), .A2(n4127), .A3(n4246), .A4(n3800), .ZN(n3801)
         );
  NAND4_X1 U4565 ( .A1(n3804), .A2(n3803), .A3(n3802), .A4(n3801), .ZN(n3805)
         );
  OR4_X1 U4566 ( .A1(n3807), .A2(n3806), .A3(n4042), .A4(n3805), .ZN(n3817) );
  AND2_X1 U4567 ( .A1(n3808), .A2(n4054), .ZN(n4074) );
  AND2_X1 U4568 ( .A1(n3810), .A2(n3809), .ZN(n4091) );
  INV_X1 U4569 ( .A(n3811), .ZN(n3813) );
  XNOR2_X1 U4570 ( .A(n4189), .B(n4167), .ZN(n4166) );
  NAND2_X1 U4571 ( .A1(n4160), .A2(n3861), .ZN(n4208) );
  NOR4_X1 U4572 ( .A1(n4146), .A2(n3814), .A3(n4166), .A4(n4208), .ZN(n3815)
         );
  NAND3_X1 U4573 ( .A1(n4074), .A2(n4091), .A3(n3815), .ZN(n3816) );
  NOR3_X1 U4574 ( .A1(n3817), .A2(n3816), .A3(n4020), .ZN(n3885) );
  NOR2_X1 U4575 ( .A1(n4325), .A2(n4312), .ZN(n3879) );
  OAI211_X1 U4576 ( .C1(n4586), .C2(n4483), .A(n3819), .B(n3818), .ZN(n3821)
         );
  NAND3_X1 U4577 ( .A1(n3821), .A2(n3820), .A3(n2695), .ZN(n3824) );
  NAND3_X1 U4578 ( .A1(n3824), .A2(n3823), .A3(n3822), .ZN(n3826) );
  NAND2_X1 U4579 ( .A1(n3826), .A2(n3825), .ZN(n3829) );
  NAND4_X1 U4580 ( .A1(n3829), .A2(n3828), .A3(n3827), .A4(n3833), .ZN(n3832)
         );
  NAND3_X1 U4581 ( .A1(n3832), .A2(n3831), .A3(n3830), .ZN(n3838) );
  INV_X1 U4582 ( .A(n3843), .ZN(n3837) );
  INV_X1 U4583 ( .A(n3833), .ZN(n3835) );
  NOR3_X1 U4584 ( .A1(n3857), .A2(n3835), .A3(n3834), .ZN(n3836) );
  AOI21_X1 U4585 ( .B1(n3838), .B2(n3837), .A(n3836), .ZN(n3842) );
  INV_X1 U4586 ( .A(n3839), .ZN(n3841) );
  NOR3_X1 U4587 ( .A1(n3842), .A2(n3841), .A3(n3840), .ZN(n3848) );
  AOI21_X1 U4588 ( .B1(n3845), .B2(n3844), .A(n3843), .ZN(n3847) );
  OAI21_X1 U4589 ( .B1(n3848), .B2(n3847), .A(n3846), .ZN(n3849) );
  OAI21_X1 U4590 ( .B1(n3857), .B2(n3850), .A(n3849), .ZN(n3853) );
  NAND3_X1 U4591 ( .A1(n3853), .A2(n3852), .A3(n3851), .ZN(n3856) );
  INV_X1 U4592 ( .A(n3854), .ZN(n3855) );
  OAI211_X1 U4593 ( .C1(n3858), .C2(n3857), .A(n3856), .B(n3855), .ZN(n3860)
         );
  AOI21_X1 U4594 ( .B1(n3860), .B2(n4201), .A(n3859), .ZN(n3864) );
  INV_X1 U4595 ( .A(n3861), .ZN(n3863) );
  OAI21_X1 U4596 ( .B1(n3864), .B2(n3863), .A(n3862), .ZN(n3867) );
  NAND3_X1 U4597 ( .A1(n3867), .A2(n3866), .A3(n3865), .ZN(n3868) );
  NAND2_X1 U4598 ( .A1(n3869), .A2(n3868), .ZN(n3873) );
  INV_X1 U4599 ( .A(n3870), .ZN(n3871) );
  AOI211_X1 U4600 ( .C1(n3874), .C2(n3873), .A(n3872), .B(n3871), .ZN(n3878)
         );
  INV_X1 U4601 ( .A(n3875), .ZN(n3876) );
  AOI22_X1 U4602 ( .A1(n2348), .A2(n3882), .B1(n3881), .B2(n3880), .ZN(n3884)
         );
  MUX2_X1 U4603 ( .A(n3885), .B(n3884), .S(n3883), .Z(n3886) );
  NOR2_X1 U4604 ( .A1(n3887), .A2(n3886), .ZN(n3888) );
  XNOR2_X1 U4605 ( .A(n3888), .B(n3981), .ZN(n3897) );
  INV_X1 U4606 ( .A(n3891), .ZN(n3896) );
  AOI21_X1 U4607 ( .B1(n3891), .B2(n3890), .A(n3889), .ZN(n3892) );
  OAI21_X1 U4608 ( .B1(n3894), .B2(n3893), .A(n3892), .ZN(n3895) );
  OAI21_X1 U4609 ( .B1(n3897), .B2(n3896), .A(n3895), .ZN(U3239) );
  MUX2_X1 U4610 ( .A(DATAO_REG_31__SCAN_IN), .B(n3898), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4611 ( .A(DATAO_REG_30__SCAN_IN), .B(n3899), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4612 ( .A(DATAO_REG_29__SCAN_IN), .B(n3900), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4613 ( .A(n4023), .B(DATAO_REG_28__SCAN_IN), .S(n3906), .Z(U3578)
         );
  MUX2_X1 U4614 ( .A(n4044), .B(DATAO_REG_27__SCAN_IN), .S(n3906), .Z(U3577)
         );
  MUX2_X1 U4615 ( .A(n4313), .B(DATAO_REG_26__SCAN_IN), .S(n3906), .Z(U3576)
         );
  MUX2_X1 U4616 ( .A(n4322), .B(DATAO_REG_25__SCAN_IN), .S(n3906), .Z(U3575)
         );
  MUX2_X1 U4617 ( .A(n4058), .B(DATAO_REG_24__SCAN_IN), .S(n3906), .Z(U3574)
         );
  MUX2_X1 U4618 ( .A(n4335), .B(DATAO_REG_23__SCAN_IN), .S(n3906), .Z(U3573)
         );
  MUX2_X1 U4619 ( .A(n4352), .B(DATAO_REG_22__SCAN_IN), .S(n3906), .Z(U3572)
         );
  MUX2_X1 U4620 ( .A(n4143), .B(DATAO_REG_21__SCAN_IN), .S(n3906), .Z(U3571)
         );
  MUX2_X1 U4621 ( .A(n4189), .B(DATAO_REG_19__SCAN_IN), .S(n3906), .Z(U3569)
         );
  MUX2_X1 U4622 ( .A(n4372), .B(DATAO_REG_18__SCAN_IN), .S(n3906), .Z(U3568)
         );
  MUX2_X1 U4623 ( .A(n4266), .B(DATAO_REG_15__SCAN_IN), .S(n3906), .Z(U3565)
         );
  MUX2_X1 U4624 ( .A(n4251), .B(DATAO_REG_14__SCAN_IN), .S(n3906), .Z(U3564)
         );
  MUX2_X1 U4625 ( .A(n4412), .B(DATAO_REG_13__SCAN_IN), .S(n3906), .Z(U3563)
         );
  MUX2_X1 U4626 ( .A(n4290), .B(DATAO_REG_12__SCAN_IN), .S(n3906), .Z(U3562)
         );
  MUX2_X1 U4627 ( .A(n4413), .B(DATAO_REG_11__SCAN_IN), .S(n3906), .Z(U3561)
         );
  MUX2_X1 U4628 ( .A(n3901), .B(DATAO_REG_10__SCAN_IN), .S(n3906), .Z(U3560)
         );
  MUX2_X1 U4629 ( .A(n3902), .B(DATAO_REG_9__SCAN_IN), .S(n3906), .Z(U3559) );
  MUX2_X1 U4630 ( .A(n3903), .B(DATAO_REG_8__SCAN_IN), .S(n3906), .Z(U3558) );
  MUX2_X1 U4631 ( .A(n3904), .B(DATAO_REG_7__SCAN_IN), .S(n3906), .Z(U3557) );
  MUX2_X1 U4632 ( .A(n2842), .B(DATAO_REG_4__SCAN_IN), .S(n3906), .Z(U3554) );
  MUX2_X1 U4633 ( .A(n3905), .B(DATAO_REG_3__SCAN_IN), .S(n3906), .Z(U3553) );
  MUX2_X1 U4634 ( .A(n3907), .B(DATAO_REG_2__SCAN_IN), .S(n3906), .Z(U3552) );
  INV_X1 U4635 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4686) );
  AOI21_X1 U4636 ( .B1(n4686), .B2(n3908), .A(n3909), .ZN(n3910) );
  MUX2_X1 U4637 ( .A(n3910), .B(n3909), .S(n2244), .Z(n3912) );
  NAND2_X1 U4638 ( .A1(n3912), .A2(n3911), .ZN(n3915) );
  AOI22_X1 U4639 ( .A1(n4579), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n3914) );
  NAND3_X1 U4640 ( .A1(n4581), .A2(n2244), .A3(n4686), .ZN(n3913) );
  NAND3_X1 U4641 ( .A1(n3915), .A2(n3914), .A3(n3913), .ZN(U3240) );
  MUX2_X1 U4642 ( .A(n3138), .B(REG2_REG_1__SCAN_IN), .S(n4496), .Z(n3916) );
  OAI21_X1 U4643 ( .B1(n2377), .B2(n2301), .A(n3916), .ZN(n3917) );
  NAND3_X1 U4644 ( .A1(n4563), .A2(n3918), .A3(n3917), .ZN(n3925) );
  AOI22_X1 U4645 ( .A1(n4579), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3924) );
  NAND2_X1 U4646 ( .A1(n3949), .A2(n4496), .ZN(n3923) );
  OAI211_X1 U4647 ( .C1(n3921), .C2(n3920), .A(n4581), .B(n3919), .ZN(n3922)
         );
  NAND4_X1 U4648 ( .A1(n3925), .A2(n3924), .A3(n3923), .A4(n3922), .ZN(U3241)
         );
  MUX2_X1 U4649 ( .A(REG1_REG_7__SCAN_IN), .B(n4695), .S(n4491), .Z(n3926) );
  XNOR2_X1 U4650 ( .A(n3927), .B(n3926), .ZN(n3928) );
  NAND2_X1 U4651 ( .A1(n3928), .A2(n4581), .ZN(n3936) );
  AOI21_X1 U4652 ( .B1(n4579), .B2(ADDR_REG_7__SCAN_IN), .A(n3929), .ZN(n3935)
         );
  OAI211_X1 U4653 ( .C1(n3932), .C2(n3931), .A(n4563), .B(n3930), .ZN(n3934)
         );
  NAND2_X1 U4654 ( .A1(n3949), .A2(n4491), .ZN(n3933) );
  NAND4_X1 U4655 ( .A1(n3936), .A2(n3935), .A3(n3934), .A4(n3933), .ZN(U3247)
         );
  INV_X1 U4656 ( .A(n4581), .ZN(n4500) );
  OAI21_X1 U4657 ( .B1(n3938), .B2(n4891), .A(n3937), .ZN(n3939) );
  AOI21_X1 U4658 ( .B1(n3940), .B2(REG1_REG_16__SCAN_IN), .A(n3959), .ZN(n3943) );
  AOI21_X1 U4659 ( .B1(n4579), .B2(ADDR_REG_16__SCAN_IN), .A(n3941), .ZN(n3942) );
  OAI21_X1 U4660 ( .B1(n4500), .B2(n3943), .A(n3942), .ZN(n3948) );
  NAND2_X1 U4661 ( .A1(n3945), .A2(n3944), .ZN(n3951) );
  AOI221_X1 U4662 ( .B1(n3946), .B2(n3952), .C1(n2541), .C2(n3952), .A(n4574), 
        .ZN(n3947) );
  AOI211_X1 U4663 ( .C1(n3949), .C2(n4487), .A(n3948), .B(n3947), .ZN(n3950)
         );
  INV_X1 U4664 ( .A(n3950), .ZN(U3256) );
  XNOR2_X1 U4665 ( .A(n3968), .B(REG2_REG_17__SCAN_IN), .ZN(n3955) );
  OR2_X1 U4666 ( .A1(n3951), .A2(n4487), .ZN(n3953) );
  AOI221_X1 U4667 ( .B1(n3955), .B2(n3974), .C1(n3954), .C2(n3974), .A(n4574), 
        .ZN(n3956) );
  INV_X1 U4668 ( .A(n3956), .ZN(n3967) );
  INV_X1 U4669 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3958) );
  INV_X1 U4670 ( .A(n3968), .ZN(n4486) );
  NOR2_X1 U4671 ( .A1(n4486), .A2(REG1_REG_17__SCAN_IN), .ZN(n3971) );
  INV_X1 U4672 ( .A(n3971), .ZN(n3957) );
  OAI21_X1 U4673 ( .B1(n3958), .B2(n3968), .A(n3957), .ZN(n3962) );
  NOR2_X1 U4674 ( .A1(n3960), .A2(n3959), .ZN(n3961) );
  NOR2_X1 U4675 ( .A1(n3961), .A2(n3962), .ZN(n3970) );
  AOI21_X1 U4676 ( .B1(n3962), .B2(n3961), .A(n3970), .ZN(n3963) );
  NOR2_X1 U4677 ( .A1(n4500), .A2(n3963), .ZN(n3964) );
  AOI211_X1 U4678 ( .C1(n4579), .C2(ADDR_REG_17__SCAN_IN), .A(n3965), .B(n3964), .ZN(n3966) );
  OAI211_X1 U4679 ( .C1(n4585), .C2(n3968), .A(n3967), .B(n3966), .ZN(U3257)
         );
  INV_X1 U4680 ( .A(REG1_REG_19__SCAN_IN), .ZN(n3969) );
  MUX2_X1 U4681 ( .A(n3969), .B(REG1_REG_19__SCAN_IN), .S(n4485), .Z(n3973) );
  INV_X1 U4682 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3972) );
  INV_X1 U4683 ( .A(n3975), .ZN(n4628) );
  AOI22_X1 U4684 ( .A1(REG1_REG_18__SCAN_IN), .A2(n3975), .B1(n4628), .B2(
        n3972), .ZN(n4583) );
  NOR2_X1 U4685 ( .A1(n3971), .A2(n3970), .ZN(n4582) );
  AOI22_X1 U4686 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4628), .B1(n3975), .B2(
        n2579), .ZN(n4577) );
  OAI21_X1 U4687 ( .B1(n4486), .B2(REG2_REG_17__SCAN_IN), .A(n3974), .ZN(n4576) );
  NOR2_X1 U4688 ( .A1(n4575), .A2(n3976), .ZN(n3978) );
  MUX2_X1 U4689 ( .A(REG2_REG_19__SCAN_IN), .B(n2596), .S(n4485), .Z(n3977) );
  XNOR2_X1 U4690 ( .A(n3978), .B(n3977), .ZN(n3983) );
  AOI21_X1 U4691 ( .B1(n4579), .B2(ADDR_REG_19__SCAN_IN), .A(n3979), .ZN(n3980) );
  OAI21_X1 U4692 ( .B1(n3981), .B2(n4585), .A(n3980), .ZN(n3982) );
  AOI21_X1 U4693 ( .B1(n3983), .B2(n4563), .A(n3982), .ZN(n3984) );
  NOR2_X2 U4694 ( .A1(n2254), .A2(n4309), .ZN(n4307) );
  XNOR2_X1 U4695 ( .A(n4307), .B(n3985), .ZN(n4423) );
  INV_X1 U4696 ( .A(n3985), .ZN(n3988) );
  NOR2_X1 U4697 ( .A1(n3987), .A2(n3986), .ZN(n4308) );
  AOI21_X1 U4698 ( .B1(n3988), .B2(n4588), .A(n4308), .ZN(n4420) );
  MUX2_X1 U4699 ( .A(n3989), .B(n4420), .S(n4617), .Z(n3990) );
  OAI21_X1 U4700 ( .B1(n4423), .B2(n4300), .A(n3990), .ZN(U3260) );
  INV_X1 U4701 ( .A(n3991), .ZN(n4003) );
  INV_X1 U4702 ( .A(n3992), .ZN(n3996) );
  OAI22_X1 U4703 ( .A1(n4315), .A2(n4011), .B1(n4617), .B2(n3993), .ZN(n3994)
         );
  AOI21_X1 U4704 ( .B1(n3996), .B2(n3995), .A(n3994), .ZN(n4002) );
  OAI21_X1 U4705 ( .B1(n4000), .B2(n3999), .A(n4617), .ZN(n4001) );
  OAI211_X1 U4706 ( .C1(n4003), .C2(n4241), .A(n4002), .B(n4001), .ZN(U3354)
         );
  NAND2_X1 U4707 ( .A1(n4004), .A2(n4302), .ZN(n4016) );
  INV_X1 U4708 ( .A(n4005), .ZN(n4014) );
  AOI22_X1 U4709 ( .A1(n4006), .A2(n4614), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4619), .ZN(n4007) );
  OAI21_X1 U4710 ( .B1(n4008), .B2(n4256), .A(n4007), .ZN(n4013) );
  OAI22_X1 U4711 ( .A1(n4325), .A2(n4011), .B1(n4010), .B2(n4009), .ZN(n4012)
         );
  AOI211_X1 U4712 ( .C1(n4014), .C2(n4601), .A(n4013), .B(n4012), .ZN(n4015)
         );
  OAI211_X1 U4713 ( .C1(n4619), .C2(n4017), .A(n4016), .B(n4015), .ZN(U3262)
         );
  XNOR2_X1 U4714 ( .A(n4019), .B(n4018), .ZN(n4318) );
  INV_X1 U4715 ( .A(n4318), .ZN(n4033) );
  NAND2_X1 U4716 ( .A1(n4021), .A2(n4020), .ZN(n4022) );
  AOI21_X1 U4717 ( .B1(n2354), .B2(n4022), .A(n4292), .ZN(n4317) );
  AOI22_X1 U4718 ( .A1(n4023), .A2(n4253), .B1(n4252), .B2(n4313), .ZN(n4026)
         );
  AOI22_X1 U4719 ( .A1(n4024), .A2(n4614), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4619), .ZN(n4025) );
  OAI211_X1 U4720 ( .C1(n4028), .C2(n4256), .A(n4026), .B(n4025), .ZN(n4031)
         );
  INV_X1 U4721 ( .A(n4043), .ZN(n4029) );
  OAI21_X1 U4722 ( .B1(n4029), .B2(n4028), .A(n4027), .ZN(n4429) );
  NOR2_X1 U4723 ( .A1(n4429), .A2(n4300), .ZN(n4030) );
  AOI211_X1 U4724 ( .C1(n4317), .C2(n4617), .A(n4031), .B(n4030), .ZN(n4032)
         );
  OAI21_X1 U4725 ( .B1(n4033), .B2(n4241), .A(n4032), .ZN(U3263) );
  NAND2_X1 U4726 ( .A1(n4034), .A2(n4035), .ZN(n4037) );
  NAND2_X1 U4727 ( .A1(n4037), .A2(n4036), .ZN(n4039) );
  INV_X1 U4728 ( .A(n4042), .ZN(n4038) );
  XNOR2_X1 U4729 ( .A(n4039), .B(n4038), .ZN(n4040) );
  NAND2_X1 U4730 ( .A1(n4040), .A2(n4609), .ZN(n4324) );
  XNOR2_X1 U4731 ( .A(n4041), .B(n4042), .ZN(n4327) );
  NAND2_X1 U4732 ( .A1(n4327), .A2(n4302), .ZN(n4052) );
  OAI21_X1 U4733 ( .B1(n4063), .B2(n4048), .A(n4043), .ZN(n4433) );
  INV_X1 U4734 ( .A(n4433), .ZN(n4050) );
  AOI22_X1 U4735 ( .A1(n4044), .A2(n4253), .B1(n4252), .B2(n4322), .ZN(n4047)
         );
  AOI22_X1 U4736 ( .A1(n4045), .A2(n4614), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4619), .ZN(n4046) );
  OAI211_X1 U4737 ( .C1(n4048), .C2(n4256), .A(n4047), .B(n4046), .ZN(n4049)
         );
  AOI21_X1 U4738 ( .B1(n4050), .B2(n4601), .A(n4049), .ZN(n4051) );
  OAI211_X1 U4739 ( .C1(n4619), .C2(n4324), .A(n4052), .B(n4051), .ZN(U3264)
         );
  XOR2_X1 U4740 ( .A(n4053), .B(n4055), .Z(n4331) );
  INV_X1 U4741 ( .A(n4331), .ZN(n4070) );
  NAND2_X1 U4742 ( .A1(n4034), .A2(n4054), .ZN(n4056) );
  XNOR2_X1 U4743 ( .A(n4056), .B(n4055), .ZN(n4057) );
  NAND2_X1 U4744 ( .A1(n4057), .A2(n4609), .ZN(n4062) );
  NAND2_X1 U4745 ( .A1(n4058), .A2(n4589), .ZN(n4059) );
  OAI21_X1 U4746 ( .B1(n4288), .B2(n4065), .A(n4059), .ZN(n4060) );
  AOI21_X1 U4747 ( .B1(n4411), .B2(n4313), .A(n4060), .ZN(n4061) );
  NAND2_X1 U4748 ( .A1(n4062), .A2(n4061), .ZN(n4330) );
  INV_X1 U4749 ( .A(n4063), .ZN(n4064) );
  OAI21_X1 U4750 ( .B1(n4075), .B2(n4065), .A(n4064), .ZN(n4437) );
  AOI22_X1 U4751 ( .A1(n4066), .A2(n4614), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4619), .ZN(n4067) );
  OAI21_X1 U4752 ( .B1(n4437), .B2(n4300), .A(n4067), .ZN(n4068) );
  AOI21_X1 U4753 ( .B1(n4330), .B2(n4617), .A(n4068), .ZN(n4069) );
  OAI21_X1 U4754 ( .B1(n4070), .B2(n4241), .A(n4069), .ZN(U3265) );
  XNOR2_X1 U4755 ( .A(n4071), .B(n4074), .ZN(n4072) );
  NAND2_X1 U4756 ( .A1(n4072), .A2(n4609), .ZN(n4337) );
  XOR2_X1 U4757 ( .A(n4074), .B(n4073), .Z(n4340) );
  NAND2_X1 U4758 ( .A1(n4340), .A2(n4302), .ZN(n4084) );
  INV_X1 U4759 ( .A(n4075), .ZN(n4076) );
  OAI21_X1 U4760 ( .B1(n2776), .B2(n4080), .A(n4076), .ZN(n4440) );
  INV_X1 U4761 ( .A(n4440), .ZN(n4082) );
  AOI22_X1 U4762 ( .A1(n4322), .A2(n4253), .B1(n4252), .B2(n4335), .ZN(n4079)
         );
  AOI22_X1 U4763 ( .A1(REG2_REG_24__SCAN_IN), .A2(n4619), .B1(n4077), .B2(
        n4614), .ZN(n4078) );
  OAI211_X1 U4764 ( .C1(n4080), .C2(n4256), .A(n4079), .B(n4078), .ZN(n4081)
         );
  AOI21_X1 U4765 ( .B1(n4082), .B2(n4601), .A(n4081), .ZN(n4083) );
  OAI211_X1 U4766 ( .C1(n4619), .C2(n4337), .A(n4084), .B(n4083), .ZN(U3266)
         );
  XNOR2_X1 U4767 ( .A(n4085), .B(n4091), .ZN(n4343) );
  INV_X1 U4768 ( .A(n4343), .ZN(n4106) );
  OAI21_X1 U4769 ( .B1(n4124), .B2(n4087), .A(n4086), .ZN(n4107) );
  INV_X1 U4770 ( .A(n4117), .ZN(n4090) );
  INV_X1 U4771 ( .A(n4088), .ZN(n4089) );
  AOI21_X1 U4772 ( .B1(n4107), .B2(n4090), .A(n4089), .ZN(n4092) );
  XNOR2_X1 U4773 ( .A(n4092), .B(n4091), .ZN(n4096) );
  OAI22_X1 U4774 ( .A1(n4093), .A2(n4612), .B1(n4098), .B2(n4288), .ZN(n4094)
         );
  AOI21_X1 U4775 ( .B1(n4589), .B2(n4352), .A(n4094), .ZN(n4095) );
  OAI21_X1 U4776 ( .B1(n4096), .B2(n4292), .A(n4095), .ZN(n4342) );
  INV_X1 U4777 ( .A(n4114), .ZN(n4099) );
  OAI21_X1 U4778 ( .B1(n4099), .B2(n4098), .A(n4097), .ZN(n4444) );
  NOR2_X1 U4779 ( .A1(n4444), .A2(n4300), .ZN(n4104) );
  NAND2_X1 U4780 ( .A1(n4100), .A2(n4614), .ZN(n4101) );
  OAI21_X1 U4781 ( .B1(n4617), .B2(n4102), .A(n4101), .ZN(n4103) );
  AOI211_X1 U4782 ( .C1(n4342), .C2(n4617), .A(n4104), .B(n4103), .ZN(n4105)
         );
  OAI21_X1 U4783 ( .B1(n4106), .B2(n4241), .A(n4105), .ZN(U3267) );
  XNOR2_X1 U4784 ( .A(n4107), .B(n4117), .ZN(n4111) );
  OAI22_X1 U4785 ( .A1(n4108), .A2(n4612), .B1(n4112), .B2(n4288), .ZN(n4109)
         );
  AOI21_X1 U4786 ( .B1(n4589), .B2(n4143), .A(n4109), .ZN(n4110) );
  OAI21_X1 U4787 ( .B1(n4111), .B2(n4292), .A(n4110), .ZN(n4347) );
  OR2_X1 U4788 ( .A1(n4129), .A2(n4112), .ZN(n4113) );
  NAND2_X1 U4789 ( .A1(n4114), .A2(n4113), .ZN(n4448) );
  AOI22_X1 U4790 ( .A1(n4619), .A2(REG2_REG_22__SCAN_IN), .B1(n4115), .B2(
        n4614), .ZN(n4116) );
  OAI21_X1 U4791 ( .B1(n4448), .B2(n4300), .A(n4116), .ZN(n4122) );
  NOR2_X1 U4792 ( .A1(n4118), .A2(n4117), .ZN(n4346) );
  INV_X1 U4793 ( .A(n4119), .ZN(n4120) );
  NOR3_X1 U4794 ( .A1(n4346), .A2(n4120), .A3(n4241), .ZN(n4121) );
  AOI211_X1 U4795 ( .C1(n4617), .C2(n4347), .A(n4122), .B(n4121), .ZN(n4123)
         );
  INV_X1 U4796 ( .A(n4123), .ZN(U3268) );
  XNOR2_X1 U4797 ( .A(n4124), .B(n4127), .ZN(n4125) );
  NAND2_X1 U4798 ( .A1(n4125), .A2(n4609), .ZN(n4354) );
  XNOR2_X1 U4799 ( .A(n4126), .B(n4127), .ZN(n4357) );
  NAND2_X1 U4800 ( .A1(n4357), .A2(n4302), .ZN(n4139) );
  INV_X1 U4801 ( .A(n4129), .ZN(n4130) );
  OAI21_X1 U4802 ( .B1(n4128), .B2(n4135), .A(n4130), .ZN(n4452) );
  INV_X1 U4803 ( .A(n4452), .ZN(n4137) );
  AOI22_X1 U4804 ( .A1(n4252), .A2(n4131), .B1(n4253), .B2(n4352), .ZN(n4134)
         );
  AOI22_X1 U4805 ( .A1(n4619), .A2(REG2_REG_21__SCAN_IN), .B1(n4132), .B2(
        n4614), .ZN(n4133) );
  OAI211_X1 U4806 ( .C1(n4135), .C2(n4256), .A(n4134), .B(n4133), .ZN(n4136)
         );
  AOI21_X1 U4807 ( .B1(n4137), .B2(n4601), .A(n4136), .ZN(n4138) );
  OAI211_X1 U4808 ( .C1(n4619), .C2(n4354), .A(n4139), .B(n4138), .ZN(U3269)
         );
  OAI21_X1 U4809 ( .B1(n4161), .B2(n4141), .A(n4140), .ZN(n4142) );
  XOR2_X1 U4810 ( .A(n4146), .B(n4142), .Z(n4150) );
  INV_X1 U4811 ( .A(n4189), .ZN(n4145) );
  AOI22_X1 U4812 ( .A1(n4143), .A2(n4411), .B1(n4588), .B2(n4151), .ZN(n4144)
         );
  OAI21_X1 U4813 ( .B1(n4145), .B2(n4393), .A(n4144), .ZN(n4149) );
  XNOR2_X1 U4814 ( .A(n4147), .B(n4146), .ZN(n4364) );
  NOR2_X1 U4815 ( .A1(n4364), .A2(n4594), .ZN(n4148) );
  AOI211_X1 U4816 ( .C1(n4609), .C2(n4150), .A(n4149), .B(n4148), .ZN(n4363)
         );
  INV_X1 U4817 ( .A(n4364), .ZN(n4157) );
  INV_X1 U4818 ( .A(n4128), .ZN(n4361) );
  NAND2_X1 U4819 ( .A1(n4174), .A2(n4151), .ZN(n4360) );
  AND3_X1 U4820 ( .A1(n4361), .A2(n4601), .A3(n4360), .ZN(n4156) );
  INV_X1 U4821 ( .A(n4152), .ZN(n4153) );
  OAI22_X1 U4822 ( .A1(n4617), .A2(n4154), .B1(n4153), .B2(n4276), .ZN(n4155)
         );
  AOI211_X1 U4823 ( .C1(n4157), .C2(n4615), .A(n4156), .B(n4155), .ZN(n4158)
         );
  OAI21_X1 U4824 ( .B1(n4363), .B2(n4619), .A(n4158), .ZN(U3270) );
  XNOR2_X1 U4825 ( .A(n4159), .B(n4166), .ZN(n4366) );
  INV_X1 U4826 ( .A(n4366), .ZN(n4178) );
  NAND2_X1 U4827 ( .A1(n4161), .A2(n4160), .ZN(n4187) );
  INV_X1 U4828 ( .A(n4162), .ZN(n4164) );
  OAI21_X1 U4829 ( .B1(n4187), .B2(n4164), .A(n4163), .ZN(n4165) );
  XOR2_X1 U4830 ( .A(n4166), .B(n4165), .Z(n4170) );
  OAI22_X1 U4831 ( .A1(n4355), .A2(n4612), .B1(n4288), .B2(n4167), .ZN(n4168)
         );
  AOI21_X1 U4832 ( .B1(n4589), .B2(n4372), .A(n4168), .ZN(n4169) );
  OAI21_X1 U4833 ( .B1(n4170), .B2(n4292), .A(n4169), .ZN(n4365) );
  NAND2_X1 U4834 ( .A1(n4171), .A2(n4172), .ZN(n4173) );
  NAND2_X1 U4835 ( .A1(n4174), .A2(n4173), .ZN(n4457) );
  AOI22_X1 U4836 ( .A1(n4619), .A2(REG2_REG_19__SCAN_IN), .B1(n2358), .B2(
        n4614), .ZN(n4175) );
  OAI21_X1 U4837 ( .B1(n4457), .B2(n4300), .A(n4175), .ZN(n4176) );
  AOI21_X1 U4838 ( .B1(n4365), .B2(n4617), .A(n4176), .ZN(n4177) );
  OAI21_X1 U4839 ( .B1(n4178), .B2(n4241), .A(n4177), .ZN(U3271) );
  OR2_X1 U4840 ( .A1(n4179), .A2(n4180), .ZN(n4182) );
  AND2_X1 U4841 ( .A1(n4182), .A2(n4181), .ZN(n4185) );
  INV_X1 U4842 ( .A(n4183), .ZN(n4184) );
  AOI21_X1 U4843 ( .B1(n4186), .B2(n4185), .A(n4184), .ZN(n4370) );
  XNOR2_X1 U4844 ( .A(n4187), .B(n4186), .ZN(n4193) );
  AOI22_X1 U4845 ( .A1(n4189), .A2(n4411), .B1(n4188), .B2(n4588), .ZN(n4190)
         );
  OAI21_X1 U4846 ( .B1(n4191), .B2(n4393), .A(n4190), .ZN(n4192) );
  AOI21_X1 U4847 ( .B1(n4193), .B2(n4609), .A(n4192), .ZN(n4369) );
  INV_X1 U4848 ( .A(n4369), .ZN(n4199) );
  OAI211_X1 U4849 ( .C1(n4210), .C2(n4194), .A(n4171), .B(n4399), .ZN(n4368)
         );
  AOI22_X1 U4850 ( .A1(n4619), .A2(REG2_REG_18__SCAN_IN), .B1(n4195), .B2(
        n4614), .ZN(n4196) );
  OAI21_X1 U4851 ( .B1(n4368), .B2(n4197), .A(n4196), .ZN(n4198) );
  AOI21_X1 U4852 ( .B1(n4199), .B2(n4617), .A(n4198), .ZN(n4200) );
  OAI21_X1 U4853 ( .B1(n4370), .B2(n4241), .A(n4200), .ZN(U3272) );
  NAND2_X1 U4854 ( .A1(n4235), .A2(n4201), .ZN(n4202) );
  XNOR2_X1 U4855 ( .A(n4202), .B(n4208), .ZN(n4203) );
  NAND2_X1 U4856 ( .A1(n4203), .A2(n4609), .ZN(n4374) );
  NAND2_X1 U4857 ( .A1(n4221), .A2(n4205), .ZN(n4226) );
  NAND2_X1 U4858 ( .A1(n4226), .A2(n4206), .ZN(n4207) );
  XOR2_X1 U4859 ( .A(n4208), .B(n4207), .Z(n4377) );
  NAND2_X1 U4860 ( .A1(n4377), .A2(n4302), .ZN(n4219) );
  INV_X1 U4861 ( .A(n4209), .ZN(n4230) );
  INV_X1 U4862 ( .A(n4210), .ZN(n4211) );
  OAI21_X1 U4863 ( .B1(n4230), .B2(n4215), .A(n4211), .ZN(n4462) );
  INV_X1 U4864 ( .A(n4462), .ZN(n4217) );
  AOI22_X1 U4865 ( .A1(n4252), .A2(n4390), .B1(n4253), .B2(n4372), .ZN(n4214)
         );
  AOI22_X1 U4866 ( .A1(n4619), .A2(REG2_REG_17__SCAN_IN), .B1(n4212), .B2(
        n4614), .ZN(n4213) );
  OAI211_X1 U4867 ( .C1(n4215), .C2(n4256), .A(n4214), .B(n4213), .ZN(n4216)
         );
  AOI21_X1 U4868 ( .B1(n4217), .B2(n4601), .A(n4216), .ZN(n4218) );
  OAI211_X1 U4869 ( .C1(n4619), .C2(n4374), .A(n4219), .B(n4218), .ZN(U3273)
         );
  NAND2_X1 U4870 ( .A1(n4221), .A2(n4220), .ZN(n4264) );
  NAND2_X1 U4871 ( .A1(n4264), .A2(n4222), .ZN(n4224) );
  AND2_X1 U4872 ( .A1(n4224), .A2(n4223), .ZN(n4229) );
  AND2_X1 U4873 ( .A1(n4226), .A2(n4225), .ZN(n4227) );
  OAI21_X1 U4874 ( .B1(n4229), .B2(n4228), .A(n4227), .ZN(n4388) );
  AOI21_X1 U4875 ( .B1(n4379), .B2(n4249), .A(n4230), .ZN(n4384) );
  AOI22_X1 U4876 ( .A1(n4252), .A2(n4266), .B1(n4253), .B2(n4380), .ZN(n4233)
         );
  AOI22_X1 U4877 ( .A1(n4619), .A2(REG2_REG_16__SCAN_IN), .B1(n4231), .B2(
        n4614), .ZN(n4232) );
  OAI211_X1 U4878 ( .C1(n4234), .C2(n4256), .A(n4233), .B(n4232), .ZN(n4239)
         );
  OAI211_X1 U4879 ( .C1(n4237), .C2(n4236), .A(n4235), .B(n4609), .ZN(n4385)
         );
  NOR2_X1 U4880 ( .A1(n4385), .A2(n4619), .ZN(n4238) );
  AOI211_X1 U4881 ( .C1(n4384), .C2(n4601), .A(n4239), .B(n4238), .ZN(n4240)
         );
  OAI21_X1 U4882 ( .B1(n4241), .B2(n4388), .A(n4240), .ZN(U3274) );
  AOI21_X1 U4883 ( .B1(n4242), .B2(n4246), .A(n4292), .ZN(n4244) );
  NAND2_X1 U4884 ( .A1(n4244), .A2(n4243), .ZN(n4392) );
  NAND2_X1 U4885 ( .A1(n4264), .A2(n4263), .ZN(n4262) );
  NAND2_X1 U4886 ( .A1(n4262), .A2(n4245), .ZN(n4247) );
  XNOR2_X1 U4887 ( .A(n4247), .B(n4246), .ZN(n4396) );
  NAND2_X1 U4888 ( .A1(n4396), .A2(n4302), .ZN(n4261) );
  INV_X1 U4889 ( .A(n4248), .ZN(n4250) );
  OAI21_X1 U4890 ( .B1(n4250), .B2(n4257), .A(n4249), .ZN(n4467) );
  INV_X1 U4891 ( .A(n4467), .ZN(n4259) );
  AOI22_X1 U4892 ( .A1(n4253), .A2(n4390), .B1(n4252), .B2(n4251), .ZN(n4255)
         );
  AOI22_X1 U4893 ( .A1(n4619), .A2(REG2_REG_15__SCAN_IN), .B1(n2350), .B2(
        n4614), .ZN(n4254) );
  OAI211_X1 U4894 ( .C1(n4257), .C2(n4256), .A(n4255), .B(n4254), .ZN(n4258)
         );
  AOI21_X1 U4895 ( .B1(n4259), .B2(n4601), .A(n4258), .ZN(n4260) );
  OAI211_X1 U4896 ( .C1(n4619), .C2(n4392), .A(n4261), .B(n4260), .ZN(U3275)
         );
  OAI21_X1 U4897 ( .B1(n4264), .B2(n4263), .A(n4262), .ZN(n4398) );
  NAND2_X1 U4898 ( .A1(n4398), .A2(n4610), .ZN(n4272) );
  XNOR2_X1 U4899 ( .A(n3746), .B(n4265), .ZN(n4270) );
  NAND2_X1 U4900 ( .A1(n4412), .A2(n4589), .ZN(n4268) );
  NAND2_X1 U4901 ( .A1(n4266), .A2(n4411), .ZN(n4267) );
  OAI211_X1 U4902 ( .C1(n4288), .C2(n4274), .A(n4268), .B(n4267), .ZN(n4269)
         );
  AOI21_X1 U4903 ( .B1(n4270), .B2(n4609), .A(n4269), .ZN(n4271) );
  NAND2_X1 U4904 ( .A1(n4272), .A2(n4271), .ZN(n4404) );
  INV_X1 U4905 ( .A(n4404), .ZN(n4282) );
  OR2_X1 U4906 ( .A1(n4273), .A2(n4274), .ZN(n4400) );
  AND3_X1 U4907 ( .A1(n4400), .A2(n4248), .A3(n4601), .ZN(n4280) );
  INV_X1 U4908 ( .A(n4275), .ZN(n4277) );
  OAI22_X1 U4909 ( .A1(n4617), .A2(n4278), .B1(n4277), .B2(n4276), .ZN(n4279)
         );
  AOI211_X1 U4910 ( .C1(n4398), .C2(n4615), .A(n4280), .B(n4279), .ZN(n4281)
         );
  OAI21_X1 U4911 ( .B1(n4282), .B2(n4619), .A(n4281), .ZN(U3276) );
  INV_X1 U4912 ( .A(n4283), .ZN(n4284) );
  AOI21_X1 U4913 ( .B1(n4286), .B2(n4285), .A(n4284), .ZN(n4287) );
  XNOR2_X1 U4914 ( .A(n4287), .B(n4294), .ZN(n4293) );
  OAI22_X1 U4915 ( .A1(n4394), .A2(n4612), .B1(n4288), .B2(n4296), .ZN(n4289)
         );
  AOI21_X1 U4916 ( .B1(n4589), .B2(n4290), .A(n4289), .ZN(n4291) );
  OAI21_X1 U4917 ( .B1(n4293), .B2(n4292), .A(n4291), .ZN(n4405) );
  INV_X1 U4918 ( .A(n4405), .ZN(n4304) );
  XOR2_X1 U4919 ( .A(n4294), .B(n4179), .Z(n4406) );
  INV_X1 U4920 ( .A(n4273), .ZN(n4295) );
  OAI21_X1 U4921 ( .B1(n4297), .B2(n4296), .A(n4295), .ZN(n4473) );
  AOI22_X1 U4922 ( .A1(n4619), .A2(REG2_REG_13__SCAN_IN), .B1(n4298), .B2(
        n4614), .ZN(n4299) );
  OAI21_X1 U4923 ( .B1(n4473), .B2(n4300), .A(n4299), .ZN(n4301) );
  AOI21_X1 U4924 ( .B1(n4406), .B2(n4302), .A(n4301), .ZN(n4303) );
  OAI21_X1 U4925 ( .B1(n4619), .B2(n4304), .A(n4303), .ZN(U3277) );
  NOR2_X1 U4926 ( .A1(n4420), .A2(n4700), .ZN(n4305) );
  AOI21_X1 U4927 ( .B1(REG1_REG_31__SCAN_IN), .B2(n4700), .A(n4305), .ZN(n4306) );
  OAI21_X1 U4928 ( .B1(n4423), .B2(n4408), .A(n4306), .ZN(U3549) );
  AOI21_X1 U4929 ( .B1(n4309), .B2(n2254), .A(n4307), .ZN(n4497) );
  INV_X1 U4930 ( .A(n4497), .ZN(n4425) );
  INV_X1 U4931 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4310) );
  AOI21_X1 U4932 ( .B1(n4309), .B2(n4588), .A(n4308), .ZN(n4499) );
  MUX2_X1 U4933 ( .A(n4310), .B(n4499), .S(n4702), .Z(n4311) );
  OAI21_X1 U4934 ( .B1(n4425), .B2(n4408), .A(n4311), .ZN(U3548) );
  INV_X1 U4935 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4319) );
  AOI22_X1 U4936 ( .A1(n4313), .A2(n4589), .B1(n4312), .B2(n4588), .ZN(n4314)
         );
  OAI21_X1 U4937 ( .B1(n4315), .B2(n4612), .A(n4314), .ZN(n4316) );
  AOI211_X1 U4938 ( .C1(n4318), .C2(n4665), .A(n4317), .B(n4316), .ZN(n4426)
         );
  MUX2_X1 U4939 ( .A(n4319), .B(n4426), .S(n4702), .Z(n4320) );
  OAI21_X1 U4940 ( .B1(n4408), .B2(n4429), .A(n4320), .ZN(U3545) );
  INV_X1 U4941 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4328) );
  AOI22_X1 U4942 ( .A1(n4322), .A2(n4589), .B1(n4321), .B2(n4588), .ZN(n4323)
         );
  OAI211_X1 U4943 ( .C1(n4325), .C2(n4612), .A(n4324), .B(n4323), .ZN(n4326)
         );
  AOI21_X1 U4944 ( .B1(n4327), .B2(n4665), .A(n4326), .ZN(n4430) );
  MUX2_X1 U4945 ( .A(n4328), .B(n4430), .S(n4702), .Z(n4329) );
  OAI21_X1 U4946 ( .B1(n4408), .B2(n4433), .A(n4329), .ZN(U3544) );
  INV_X1 U4947 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4332) );
  AOI21_X1 U4948 ( .B1(n4331), .B2(n4665), .A(n4330), .ZN(n4434) );
  MUX2_X1 U4949 ( .A(n4332), .B(n4434), .S(n4702), .Z(n4333) );
  OAI21_X1 U4950 ( .B1(n4408), .B2(n4437), .A(n4333), .ZN(U3543) );
  INV_X1 U4951 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4918) );
  AOI22_X1 U4952 ( .A1(n4335), .A2(n4589), .B1(n4588), .B2(n4334), .ZN(n4336)
         );
  OAI211_X1 U4953 ( .C1(n4338), .C2(n4612), .A(n4337), .B(n4336), .ZN(n4339)
         );
  AOI21_X1 U4954 ( .B1(n4340), .B2(n4665), .A(n4339), .ZN(n4438) );
  MUX2_X1 U4955 ( .A(n4918), .B(n4438), .S(n4702), .Z(n4341) );
  OAI21_X1 U4956 ( .B1(n4408), .B2(n4440), .A(n4341), .ZN(U3542) );
  INV_X1 U4957 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4344) );
  AOI21_X1 U4958 ( .B1(n4343), .B2(n4665), .A(n4342), .ZN(n4441) );
  MUX2_X1 U4959 ( .A(n4344), .B(n4441), .S(n4702), .Z(n4345) );
  OAI21_X1 U4960 ( .B1(n4408), .B2(n4444), .A(n4345), .ZN(U3541) );
  INV_X1 U4961 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4349) );
  INV_X1 U4962 ( .A(n4665), .ZN(n4387) );
  NOR2_X1 U4963 ( .A1(n4346), .A2(n4387), .ZN(n4348) );
  AOI21_X1 U4964 ( .B1(n4348), .B2(n4119), .A(n4347), .ZN(n4445) );
  MUX2_X1 U4965 ( .A(n4349), .B(n4445), .S(n4702), .Z(n4350) );
  OAI21_X1 U4966 ( .B1(n4408), .B2(n4448), .A(n4350), .ZN(U3540) );
  INV_X1 U4967 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4358) );
  AOI22_X1 U4968 ( .A1(n4352), .A2(n4411), .B1(n4588), .B2(n4351), .ZN(n4353)
         );
  OAI211_X1 U4969 ( .C1(n4355), .C2(n4393), .A(n4354), .B(n4353), .ZN(n4356)
         );
  AOI21_X1 U4970 ( .B1(n4357), .B2(n4665), .A(n4356), .ZN(n4449) );
  MUX2_X1 U4971 ( .A(n4358), .B(n4449), .S(n4702), .Z(n4359) );
  OAI21_X1 U4972 ( .B1(n4408), .B2(n4452), .A(n4359), .ZN(U3539) );
  NAND3_X1 U4973 ( .A1(n4361), .A2(n4360), .A3(n4399), .ZN(n4362) );
  OAI211_X1 U4974 ( .C1(n4364), .C2(n4643), .A(n4363), .B(n4362), .ZN(n4453)
         );
  MUX2_X1 U4975 ( .A(REG1_REG_20__SCAN_IN), .B(n4453), .S(n4702), .Z(U3538) );
  AOI21_X1 U4976 ( .B1(n4366), .B2(n4665), .A(n4365), .ZN(n4455) );
  MUX2_X1 U4977 ( .A(n4455), .B(n3969), .S(n4700), .Z(n4367) );
  OAI21_X1 U4978 ( .B1(n4408), .B2(n4457), .A(n4367), .ZN(U3537) );
  OAI211_X1 U4979 ( .C1(n4370), .C2(n4387), .A(n4369), .B(n4368), .ZN(n4458)
         );
  MUX2_X1 U4980 ( .A(REG1_REG_18__SCAN_IN), .B(n4458), .S(n4702), .Z(U3536) );
  AOI22_X1 U4981 ( .A1(n4372), .A2(n4411), .B1(n4588), .B2(n4371), .ZN(n4373)
         );
  OAI211_X1 U4982 ( .C1(n4375), .C2(n4393), .A(n4374), .B(n4373), .ZN(n4376)
         );
  AOI21_X1 U4983 ( .B1(n4377), .B2(n4665), .A(n4376), .ZN(n4460) );
  MUX2_X1 U4984 ( .A(n4460), .B(n3958), .S(n4700), .Z(n4378) );
  OAI21_X1 U4985 ( .B1(n4408), .B2(n4462), .A(n4378), .ZN(U3535) );
  AOI22_X1 U4986 ( .A1(n4380), .A2(n4411), .B1(n4588), .B2(n4379), .ZN(n4381)
         );
  OAI21_X1 U4987 ( .B1(n4382), .B2(n4393), .A(n4381), .ZN(n4383) );
  AOI21_X1 U4988 ( .B1(n4384), .B2(n4399), .A(n4383), .ZN(n4386) );
  OAI211_X1 U4989 ( .C1(n4388), .C2(n4387), .A(n4386), .B(n4385), .ZN(n4463)
         );
  MUX2_X1 U4990 ( .A(REG1_REG_16__SCAN_IN), .B(n4463), .S(n4702), .Z(U3534) );
  AOI22_X1 U4991 ( .A1(n4390), .A2(n4411), .B1(n4389), .B2(n4588), .ZN(n4391)
         );
  OAI211_X1 U4992 ( .C1(n4394), .C2(n4393), .A(n4392), .B(n4391), .ZN(n4395)
         );
  AOI21_X1 U4993 ( .B1(n4396), .B2(n4665), .A(n4395), .ZN(n4464) );
  MUX2_X1 U4994 ( .A(n4891), .B(n4464), .S(n4702), .Z(n4397) );
  OAI21_X1 U4995 ( .B1(n4408), .B2(n4467), .A(n4397), .ZN(U3533) );
  NAND2_X1 U4996 ( .A1(n4398), .A2(n4683), .ZN(n4402) );
  NAND3_X1 U4997 ( .A1(n4400), .A2(n4248), .A3(n4399), .ZN(n4401) );
  NAND2_X1 U4998 ( .A1(n4402), .A2(n4401), .ZN(n4403) );
  MUX2_X1 U4999 ( .A(REG1_REG_14__SCAN_IN), .B(n4468), .S(n4702), .Z(U3532) );
  AOI21_X1 U5000 ( .B1(n4406), .B2(n4665), .A(n4405), .ZN(n4469) );
  MUX2_X1 U5001 ( .A(n3358), .B(n4469), .S(n4702), .Z(n4407) );
  OAI21_X1 U5002 ( .B1(n4408), .B2(n4473), .A(n4407), .ZN(U3531) );
  NAND2_X1 U5003 ( .A1(n4409), .A2(n4665), .ZN(n4417) );
  AOI22_X1 U5004 ( .A1(n4412), .A2(n4411), .B1(n4588), .B2(n4410), .ZN(n4416)
         );
  NAND2_X1 U5005 ( .A1(n4413), .A2(n4589), .ZN(n4414) );
  NAND4_X1 U5006 ( .A1(n4417), .A2(n4416), .A3(n4415), .A4(n4414), .ZN(n4474)
         );
  MUX2_X1 U5007 ( .A(REG1_REG_12__SCAN_IN), .B(n4474), .S(n4702), .Z(n4418) );
  AOI21_X1 U5008 ( .B1(n4476), .B2(n2808), .A(n4418), .ZN(n4419) );
  INV_X1 U5009 ( .A(n4419), .ZN(U3530) );
  NOR2_X1 U5010 ( .A1(n4420), .A2(n4684), .ZN(n4421) );
  AOI21_X1 U5011 ( .B1(REG0_REG_31__SCAN_IN), .B2(n4684), .A(n4421), .ZN(n4422) );
  OAI21_X1 U5012 ( .B1(n4423), .B2(n4472), .A(n4422), .ZN(U3517) );
  INV_X1 U5013 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4920) );
  MUX2_X1 U5014 ( .A(n4920), .B(n4499), .S(n4685), .Z(n4424) );
  OAI21_X1 U5015 ( .B1(n4425), .B2(n4472), .A(n4424), .ZN(U3516) );
  INV_X1 U5016 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4427) );
  MUX2_X1 U5017 ( .A(n4427), .B(n4426), .S(n4685), .Z(n4428) );
  OAI21_X1 U5018 ( .B1(n4429), .B2(n4472), .A(n4428), .ZN(U3513) );
  INV_X1 U5019 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4431) );
  MUX2_X1 U5020 ( .A(n4431), .B(n4430), .S(n4685), .Z(n4432) );
  OAI21_X1 U5021 ( .B1(n4433), .B2(n4472), .A(n4432), .ZN(U3512) );
  INV_X1 U5022 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4435) );
  MUX2_X1 U5023 ( .A(n4435), .B(n4434), .S(n4685), .Z(n4436) );
  OAI21_X1 U5024 ( .B1(n4437), .B2(n4472), .A(n4436), .ZN(U3511) );
  INV_X1 U5025 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4917) );
  MUX2_X1 U5026 ( .A(n4917), .B(n4438), .S(n4685), .Z(n4439) );
  OAI21_X1 U5027 ( .B1(n4440), .B2(n4472), .A(n4439), .ZN(U3510) );
  INV_X1 U5028 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4442) );
  MUX2_X1 U5029 ( .A(n4442), .B(n4441), .S(n4685), .Z(n4443) );
  OAI21_X1 U5030 ( .B1(n4444), .B2(n4472), .A(n4443), .ZN(U3509) );
  INV_X1 U5031 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4446) );
  MUX2_X1 U5032 ( .A(n4446), .B(n4445), .S(n4685), .Z(n4447) );
  OAI21_X1 U5033 ( .B1(n4448), .B2(n4472), .A(n4447), .ZN(U3508) );
  INV_X1 U5034 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4450) );
  MUX2_X1 U5035 ( .A(n4450), .B(n4449), .S(n4685), .Z(n4451) );
  OAI21_X1 U5036 ( .B1(n4452), .B2(n4472), .A(n4451), .ZN(U3507) );
  MUX2_X1 U5037 ( .A(REG0_REG_20__SCAN_IN), .B(n4453), .S(n4685), .Z(U3506) );
  INV_X1 U5038 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4454) );
  MUX2_X1 U5039 ( .A(n4455), .B(n4454), .S(n4684), .Z(n4456) );
  OAI21_X1 U5040 ( .B1(n4457), .B2(n4472), .A(n4456), .ZN(U3505) );
  MUX2_X1 U5041 ( .A(REG0_REG_18__SCAN_IN), .B(n4458), .S(n4685), .Z(U3503) );
  INV_X1 U5042 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4459) );
  MUX2_X1 U5043 ( .A(n4460), .B(n4459), .S(n4684), .Z(n4461) );
  OAI21_X1 U5044 ( .B1(n4462), .B2(n4472), .A(n4461), .ZN(U3501) );
  MUX2_X1 U5045 ( .A(REG0_REG_16__SCAN_IN), .B(n4463), .S(n4685), .Z(U3499) );
  INV_X1 U5046 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4465) );
  MUX2_X1 U5047 ( .A(n4465), .B(n4464), .S(n4685), .Z(n4466) );
  OAI21_X1 U5048 ( .B1(n4467), .B2(n4472), .A(n4466), .ZN(U3497) );
  MUX2_X1 U5049 ( .A(n4468), .B(REG0_REG_14__SCAN_IN), .S(n4684), .Z(U3495) );
  INV_X1 U5050 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4470) );
  MUX2_X1 U5051 ( .A(n4470), .B(n4469), .S(n4685), .Z(n4471) );
  OAI21_X1 U5052 ( .B1(n4473), .B2(n4472), .A(n4471), .ZN(U3493) );
  MUX2_X1 U5053 ( .A(REG0_REG_12__SCAN_IN), .B(n4474), .S(n4685), .Z(n4475) );
  AOI21_X1 U5054 ( .B1(n4476), .B2(n4651), .A(n4475), .ZN(n4477) );
  INV_X1 U5055 ( .A(n4477), .ZN(U3491) );
  MUX2_X1 U5056 ( .A(DATAI_30_), .B(n4478), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U5057 ( .A(n4479), .B(DATAI_28_), .S(U3149), .Z(U3324) );
  MUX2_X1 U5058 ( .A(n2754), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5059 ( .A(n4480), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U5060 ( .A(DATAI_24_), .B(n4481), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U5061 ( .A(DATAI_22_), .B(n4482), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U5062 ( .A(n4483), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5063 ( .A(DATAI_20_), .B(n4484), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5064 ( .A(n4485), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5065 ( .A(n4486), .B(DATAI_17_), .S(U3149), .Z(U3335) );
  MUX2_X1 U5066 ( .A(n4487), .B(DATAI_16_), .S(U3149), .Z(U3336) );
  MUX2_X1 U5067 ( .A(n4488), .B(DATAI_15_), .S(U3149), .Z(U3337) );
  MUX2_X1 U5068 ( .A(n4489), .B(DATAI_14_), .S(U3149), .Z(U3338) );
  MUX2_X1 U5069 ( .A(n4490), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U5070 ( .A(n4519), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5071 ( .A(n4491), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5072 ( .A(n4492), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5073 ( .A(DATAI_4_), .B(n4493), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5074 ( .A(n4494), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5075 ( .A(n4495), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5076 ( .A(n4496), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U5077 ( .A(DATAI_0_), .B(n2244), .S(STATE_REG_SCAN_IN), .Z(U3352) );
  OAI21_X1 U5078 ( .B1(n4619), .B2(n4499), .A(n4498), .ZN(U3261) );
  AOI211_X1 U5079 ( .C1(n4877), .C2(n4502), .A(n4501), .B(n4500), .ZN(n4503)
         );
  AOI211_X1 U5080 ( .C1(ADDR_REG_6__SCAN_IN), .C2(n4579), .A(n4504), .B(n4503), 
        .ZN(n4508) );
  OAI211_X1 U5081 ( .C1(REG2_REG_6__SCAN_IN), .C2(n4506), .A(n4563), .B(n4505), 
        .ZN(n4507) );
  OAI211_X1 U5082 ( .C1(n4585), .C2(n4509), .A(n4508), .B(n4507), .ZN(U3246)
         );
  OAI211_X1 U5083 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4511), .A(n4563), .B(n4510), 
        .ZN(n4513) );
  NAND2_X1 U5084 ( .A1(n4513), .A2(n4512), .ZN(n4514) );
  AOI21_X1 U5085 ( .B1(n4579), .B2(ADDR_REG_8__SCAN_IN), .A(n4514), .ZN(n4518)
         );
  OAI211_X1 U5086 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4516), .A(n4581), .B(n4515), 
        .ZN(n4517) );
  OAI211_X1 U5087 ( .C1(n4585), .C2(n4634), .A(n4518), .B(n4517), .ZN(U3248)
         );
  INV_X1 U5088 ( .A(n4519), .ZN(n4528) );
  OAI211_X1 U5089 ( .C1(n4522), .C2(n4521), .A(n4581), .B(n4520), .ZN(n4527)
         );
  OAI211_X1 U5090 ( .C1(n4525), .C2(n4524), .A(n4563), .B(n4523), .ZN(n4526)
         );
  OAI211_X1 U5091 ( .C1(n4585), .C2(n4528), .A(n4527), .B(n4526), .ZN(n4529)
         );
  AOI211_X1 U5092 ( .C1(n4579), .C2(ADDR_REG_9__SCAN_IN), .A(n4530), .B(n4529), 
        .ZN(n4531) );
  INV_X1 U5093 ( .A(n4531), .ZN(U3249) );
  NAND2_X1 U5094 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n5084) );
  OAI211_X1 U5095 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4533), .A(n4563), .B(n4532), .ZN(n4534) );
  NAND2_X1 U5096 ( .A1(n5084), .A2(n4534), .ZN(n4535) );
  AOI21_X1 U5097 ( .B1(ADDR_REG_10__SCAN_IN), .B2(n4579), .A(n4535), .ZN(n4539) );
  OAI211_X1 U5098 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4537), .A(n4581), .B(n4536), .ZN(n4538) );
  OAI211_X1 U5099 ( .C1(n4585), .C2(n4540), .A(n4539), .B(n4538), .ZN(U3250)
         );
  OAI211_X1 U5100 ( .C1(n4543), .C2(n4542), .A(n4541), .B(n4581), .ZN(n4548)
         );
  OAI211_X1 U5101 ( .C1(n4546), .C2(n4545), .A(n4563), .B(n4544), .ZN(n4547)
         );
  OAI211_X1 U5102 ( .C1(n4585), .C2(n4549), .A(n4548), .B(n4547), .ZN(n4550)
         );
  AOI211_X1 U5103 ( .C1(n4579), .C2(ADDR_REG_11__SCAN_IN), .A(n4551), .B(n4550), .ZN(n4552) );
  INV_X1 U5104 ( .A(n4552), .ZN(U3251) );
  OAI211_X1 U5105 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4554), .A(n4563), .B(n4553), .ZN(n4556) );
  NAND2_X1 U5106 ( .A1(n4556), .A2(n4555), .ZN(n4557) );
  AOI21_X1 U5107 ( .B1(n4579), .B2(ADDR_REG_12__SCAN_IN), .A(n4557), .ZN(n4561) );
  OAI211_X1 U5108 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4559), .A(n4581), .B(n4558), .ZN(n4560) );
  OAI211_X1 U5109 ( .C1(n4585), .C2(n4631), .A(n4561), .B(n4560), .ZN(U3252)
         );
  AOI21_X1 U5110 ( .B1(n2518), .B2(n4630), .A(n4562), .ZN(n4566) );
  OAI21_X1 U5111 ( .B1(n4566), .B2(n4565), .A(n4563), .ZN(n4564) );
  AOI21_X1 U5112 ( .B1(n4566), .B2(n4565), .A(n4564), .ZN(n4567) );
  AOI211_X1 U5113 ( .C1(n4579), .C2(ADDR_REG_13__SCAN_IN), .A(n4568), .B(n4567), .ZN(n4573) );
  OAI211_X1 U5114 ( .C1(n4571), .C2(n4570), .A(n4581), .B(n4569), .ZN(n4572)
         );
  OAI211_X1 U5115 ( .C1(n4585), .C2(n4630), .A(n4573), .B(n4572), .ZN(U3253)
         );
  OAI211_X1 U5116 ( .C1(n4583), .C2(n4582), .A(n4581), .B(n4580), .ZN(n4584)
         );
  OAI21_X1 U5117 ( .B1(n2694), .B2(n4586), .A(n3262), .ZN(n4597) );
  AOI22_X1 U5118 ( .A1(n2821), .A2(n4589), .B1(n4588), .B2(n4587), .ZN(n4590)
         );
  OAI21_X1 U5119 ( .B1(n3243), .B2(n4612), .A(n4590), .ZN(n4596) );
  OAI21_X1 U5120 ( .B1(n4593), .B2(n4592), .A(n4591), .ZN(n4644) );
  NOR2_X1 U5121 ( .A1(n4644), .A2(n4594), .ZN(n4595) );
  AOI211_X1 U5122 ( .C1(n4609), .C2(n4597), .A(n4596), .B(n4595), .ZN(n4641)
         );
  AOI22_X1 U5123 ( .A1(REG2_REG_1__SCAN_IN), .A2(n4619), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4614), .ZN(n4604) );
  INV_X1 U5124 ( .A(n4644), .ZN(n4602) );
  OAI21_X1 U5125 ( .B1(n4599), .B2(n4607), .A(n4598), .ZN(n4642) );
  INV_X1 U5126 ( .A(n4642), .ZN(n4600) );
  AOI22_X1 U5127 ( .A1(n4602), .A2(n4615), .B1(n4601), .B2(n4600), .ZN(n4603)
         );
  OAI211_X1 U5128 ( .C1(n4619), .C2(n4641), .A(n4604), .B(n4603), .ZN(U3289)
         );
  INV_X1 U5129 ( .A(n4605), .ZN(n4606) );
  NOR2_X1 U5130 ( .A1(n4607), .A2(n4606), .ZN(n4638) );
  INV_X1 U5131 ( .A(n4608), .ZN(n4613) );
  OAI21_X1 U5132 ( .B1(n4610), .B2(n4609), .A(n4639), .ZN(n4611) );
  OAI21_X1 U5133 ( .B1(n3177), .B2(n4612), .A(n4611), .ZN(n4637) );
  AOI21_X1 U5134 ( .B1(n4638), .B2(n4613), .A(n4637), .ZN(n4618) );
  AOI22_X1 U5135 ( .A1(n4639), .A2(n4615), .B1(REG3_REG_0__SCAN_IN), .B2(n4614), .ZN(n4616) );
  OAI221_X1 U5136 ( .B1(n4619), .B2(n4618), .C1(n4617), .C2(n2377), .A(n4616), 
        .ZN(U3290) );
  INV_X1 U5137 ( .A(D_REG_31__SCAN_IN), .ZN(n4983) );
  NOR2_X1 U5138 ( .A1(n4624), .A2(n4983), .ZN(U3291) );
  AND2_X1 U5139 ( .A1(D_REG_30__SCAN_IN), .A2(n4622), .ZN(U3292) );
  INV_X1 U5140 ( .A(D_REG_29__SCAN_IN), .ZN(n4952) );
  NOR2_X1 U5141 ( .A1(n4624), .A2(n4952), .ZN(U3293) );
  AND2_X1 U5142 ( .A1(D_REG_28__SCAN_IN), .A2(n4622), .ZN(U3294) );
  INV_X1 U5143 ( .A(D_REG_27__SCAN_IN), .ZN(n4824) );
  NOR2_X1 U5144 ( .A1(n4624), .A2(n4824), .ZN(U3295) );
  AND2_X1 U5145 ( .A1(D_REG_26__SCAN_IN), .A2(n4622), .ZN(U3296) );
  INV_X1 U5146 ( .A(D_REG_25__SCAN_IN), .ZN(n4978) );
  NOR2_X1 U5147 ( .A1(n4624), .A2(n4978), .ZN(U3297) );
  AND2_X1 U5148 ( .A1(D_REG_24__SCAN_IN), .A2(n4622), .ZN(U3298) );
  AND2_X1 U5149 ( .A1(D_REG_23__SCAN_IN), .A2(n4622), .ZN(U3299) );
  AND2_X1 U5150 ( .A1(D_REG_22__SCAN_IN), .A2(n4622), .ZN(U3300) );
  AND2_X1 U5151 ( .A1(D_REG_21__SCAN_IN), .A2(n4622), .ZN(U3301) );
  AND2_X1 U5152 ( .A1(D_REG_20__SCAN_IN), .A2(n4622), .ZN(U3302) );
  INV_X1 U5153 ( .A(D_REG_19__SCAN_IN), .ZN(n4957) );
  NOR2_X1 U5154 ( .A1(n4624), .A2(n4957), .ZN(U3303) );
  AND2_X1 U5155 ( .A1(D_REG_18__SCAN_IN), .A2(n4622), .ZN(U3304) );
  AND2_X1 U5156 ( .A1(D_REG_17__SCAN_IN), .A2(n4622), .ZN(U3305) );
  INV_X1 U5157 ( .A(D_REG_16__SCAN_IN), .ZN(n4936) );
  NOR2_X1 U5158 ( .A1(n4624), .A2(n4936), .ZN(U3306) );
  AND2_X1 U5159 ( .A1(D_REG_15__SCAN_IN), .A2(n4622), .ZN(U3307) );
  INV_X1 U5160 ( .A(D_REG_14__SCAN_IN), .ZN(n4986) );
  NOR2_X1 U5161 ( .A1(n4624), .A2(n4986), .ZN(U3308) );
  NOR2_X1 U5162 ( .A1(n4624), .A2(n4620), .ZN(U3309) );
  NOR2_X1 U5163 ( .A1(n4624), .A2(n4822), .ZN(U3310) );
  INV_X1 U5164 ( .A(D_REG_11__SCAN_IN), .ZN(n4977) );
  NOR2_X1 U5165 ( .A1(n4624), .A2(n4977), .ZN(U3311) );
  INV_X1 U5166 ( .A(D_REG_10__SCAN_IN), .ZN(n4940) );
  NOR2_X1 U5167 ( .A1(n4624), .A2(n4940), .ZN(U3312) );
  AND2_X1 U5168 ( .A1(D_REG_9__SCAN_IN), .A2(n4622), .ZN(U3313) );
  AND2_X1 U5169 ( .A1(D_REG_8__SCAN_IN), .A2(n4622), .ZN(U3314) );
  NOR2_X1 U5170 ( .A1(n4624), .A2(n4621), .ZN(U3315) );
  INV_X1 U5171 ( .A(D_REG_6__SCAN_IN), .ZN(n4933) );
  NOR2_X1 U5172 ( .A1(n4624), .A2(n4933), .ZN(U3316) );
  AND2_X1 U5173 ( .A1(D_REG_5__SCAN_IN), .A2(n4622), .ZN(U3317) );
  INV_X1 U5174 ( .A(D_REG_4__SCAN_IN), .ZN(n4934) );
  NOR2_X1 U5175 ( .A1(n4624), .A2(n4934), .ZN(U3318) );
  AND2_X1 U5176 ( .A1(D_REG_3__SCAN_IN), .A2(n4622), .ZN(U3319) );
  NOR2_X1 U5177 ( .A1(n4624), .A2(n4623), .ZN(U3320) );
  OAI21_X1 U5178 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4625), .ZN(
        n4626) );
  INV_X1 U5179 ( .A(n4626), .ZN(U3329) );
  INV_X1 U5180 ( .A(DATAI_18_), .ZN(n4627) );
  AOI22_X1 U5181 ( .A1(STATE_REG_SCAN_IN), .A2(n4628), .B1(n4627), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5182 ( .A(DATAI_13_), .ZN(n4629) );
  AOI22_X1 U5183 ( .A1(STATE_REG_SCAN_IN), .A2(n4630), .B1(n4629), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5184 ( .A(DATAI_12_), .ZN(n4906) );
  AOI22_X1 U5185 ( .A1(STATE_REG_SCAN_IN), .A2(n4631), .B1(n4906), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5186 ( .A1(U3149), .A2(n4632), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4633) );
  INV_X1 U5187 ( .A(n4633), .ZN(U3342) );
  INV_X1 U5188 ( .A(DATAI_8_), .ZN(n4788) );
  AOI22_X1 U5189 ( .A1(STATE_REG_SCAN_IN), .A2(n4634), .B1(n4788), .B2(U3149), 
        .ZN(U3344) );
  OAI22_X1 U5190 ( .A1(U3149), .A2(n4635), .B1(DATAI_6_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4636) );
  INV_X1 U5191 ( .A(n4636), .ZN(U3346) );
  AOI211_X1 U5192 ( .C1(n4683), .C2(n4639), .A(n4638), .B(n4637), .ZN(n4687)
         );
  INV_X1 U5193 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4640) );
  AOI22_X1 U5194 ( .A1(n4685), .A2(n4687), .B1(n4640), .B2(n4684), .ZN(U3467)
         );
  INV_X1 U5195 ( .A(n4641), .ZN(n4646) );
  OAI22_X1 U5196 ( .A1(n4644), .A2(n4643), .B1(n4678), .B2(n4642), .ZN(n4645)
         );
  NOR2_X1 U5197 ( .A1(n4646), .A2(n4645), .ZN(n4688) );
  INV_X1 U5198 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4647) );
  AOI22_X1 U5199 ( .A1(n4685), .A2(n4688), .B1(n4647), .B2(n4684), .ZN(U3469)
         );
  INV_X1 U5200 ( .A(n4648), .ZN(n4649) );
  AOI21_X1 U5201 ( .B1(n4683), .B2(n4650), .A(n4649), .ZN(n4691) );
  AOI22_X1 U5202 ( .A1(n4651), .A2(n4689), .B1(REG0_REG_2__SCAN_IN), .B2(n4684), .ZN(n4652) );
  OAI21_X1 U5203 ( .B1(n4691), .B2(n4684), .A(n4652), .ZN(U3471) );
  INV_X1 U5204 ( .A(n4653), .ZN(n4655) );
  AOI211_X1 U5205 ( .C1(n4656), .C2(n4683), .A(n4655), .B(n4654), .ZN(n4693)
         );
  INV_X1 U5206 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4657) );
  AOI22_X1 U5207 ( .A1(n4685), .A2(n4693), .B1(n4657), .B2(n4684), .ZN(U3475)
         );
  NOR2_X1 U5208 ( .A1(n4658), .A2(n4678), .ZN(n4660) );
  AOI211_X1 U5209 ( .C1(n4683), .C2(n4661), .A(n4660), .B(n4659), .ZN(n4694)
         );
  INV_X1 U5210 ( .A(REG0_REG_6__SCAN_IN), .ZN(n4662) );
  AOI22_X1 U5211 ( .A1(n4685), .A2(n4694), .B1(n4662), .B2(n4684), .ZN(U3479)
         );
  AOI211_X1 U5212 ( .C1(n4666), .C2(n4665), .A(n4664), .B(n4663), .ZN(n4696)
         );
  INV_X1 U5213 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4667) );
  AOI22_X1 U5214 ( .A1(n4685), .A2(n4696), .B1(n4667), .B2(n4684), .ZN(U3481)
         );
  NOR3_X1 U5215 ( .A1(n4669), .A2(n4668), .A3(n4678), .ZN(n4671) );
  AOI211_X1 U5216 ( .C1(n4672), .C2(n4683), .A(n4671), .B(n4670), .ZN(n4697)
         );
  INV_X1 U5217 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4826) );
  AOI22_X1 U5218 ( .A1(n4685), .A2(n4697), .B1(n4826), .B2(n4684), .ZN(U3483)
         );
  NOR3_X1 U5219 ( .A1(n4674), .A2(n4673), .A3(n4678), .ZN(n4676) );
  AOI211_X1 U5220 ( .C1(n4677), .C2(n4683), .A(n4676), .B(n4675), .ZN(n4699)
         );
  INV_X1 U5221 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4829) );
  AOI22_X1 U5222 ( .A1(n4685), .A2(n4699), .B1(n4829), .B2(n4684), .ZN(U3487)
         );
  NOR2_X1 U5223 ( .A1(n4679), .A2(n4678), .ZN(n4681) );
  AOI211_X1 U5224 ( .C1(n4683), .C2(n4682), .A(n4681), .B(n4680), .ZN(n4701)
         );
  INV_X1 U5225 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4963) );
  AOI22_X1 U5226 ( .A1(n4685), .A2(n4701), .B1(n4963), .B2(n4684), .ZN(U3489)
         );
  AOI22_X1 U5227 ( .A1(n4702), .A2(n4687), .B1(n4686), .B2(n4700), .ZN(U3518)
         );
  AOI22_X1 U5228 ( .A1(n4702), .A2(n4688), .B1(n3157), .B2(n4700), .ZN(U3519)
         );
  AOI22_X1 U5229 ( .A1(n2808), .A2(n4689), .B1(REG1_REG_2__SCAN_IN), .B2(n4700), .ZN(n4690) );
  OAI21_X1 U5230 ( .B1(n4691), .B2(n4700), .A(n4690), .ZN(U3520) );
  INV_X1 U5231 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4692) );
  AOI22_X1 U5232 ( .A1(n4702), .A2(n4693), .B1(n4692), .B2(n4700), .ZN(U3522)
         );
  AOI22_X1 U5233 ( .A1(n4702), .A2(n4694), .B1(n4877), .B2(n4700), .ZN(U3524)
         );
  AOI22_X1 U5234 ( .A1(n4702), .A2(n4696), .B1(n4695), .B2(n4700), .ZN(U3525)
         );
  INV_X1 U5235 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4839) );
  AOI22_X1 U5236 ( .A1(n4702), .A2(n4697), .B1(n4839), .B2(n4700), .ZN(U3526)
         );
  INV_X1 U5237 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4698) );
  AOI22_X1 U5238 ( .A1(n4702), .A2(n4699), .B1(n4698), .B2(n4700), .ZN(U3528)
         );
  AOI22_X1 U5239 ( .A1(n4702), .A2(n4701), .B1(n4846), .B2(n4700), .ZN(U3529)
         );
  AOI22_X1 U5240 ( .A1(DATAI_19_), .A2(keyinput237), .B1(DATAI_29_), .B2(
        keyinput192), .ZN(n4703) );
  OAI221_X1 U5241 ( .B1(DATAI_19_), .B2(keyinput237), .C1(DATAI_29_), .C2(
        keyinput192), .A(n4703), .ZN(n4710) );
  AOI22_X1 U5242 ( .A1(DATAI_15_), .A2(keyinput226), .B1(DATAI_14_), .B2(
        keyinput230), .ZN(n4704) );
  OAI221_X1 U5243 ( .B1(DATAI_15_), .B2(keyinput226), .C1(DATAI_14_), .C2(
        keyinput230), .A(n4704), .ZN(n4709) );
  AOI22_X1 U5244 ( .A1(DATAI_4_), .A2(keyinput201), .B1(DATAI_10_), .B2(
        keyinput150), .ZN(n4705) );
  OAI221_X1 U5245 ( .B1(DATAI_4_), .B2(keyinput201), .C1(DATAI_10_), .C2(
        keyinput150), .A(n4705), .ZN(n4708) );
  AOI22_X1 U5246 ( .A1(DATAI_2_), .A2(keyinput136), .B1(REG3_REG_14__SCAN_IN), 
        .B2(keyinput247), .ZN(n4706) );
  OAI221_X1 U5247 ( .B1(DATAI_2_), .B2(keyinput136), .C1(REG3_REG_14__SCAN_IN), 
        .C2(keyinput247), .A(n4706), .ZN(n4707) );
  NOR4_X1 U5248 ( .A1(n4710), .A2(n4709), .A3(n4708), .A4(n4707), .ZN(n4738)
         );
  AOI22_X1 U5249 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput161), .B1(
        REG3_REG_7__SCAN_IN), .B2(keyinput152), .ZN(n4711) );
  OAI221_X1 U5250 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput161), .C1(
        REG3_REG_7__SCAN_IN), .C2(keyinput152), .A(n4711), .ZN(n4718) );
  AOI22_X1 U5251 ( .A1(n2244), .A2(keyinput148), .B1(IR_REG_5__SCAN_IN), .B2(
        keyinput179), .ZN(n4712) );
  OAI221_X1 U5252 ( .B1(n2244), .B2(keyinput148), .C1(IR_REG_5__SCAN_IN), .C2(
        keyinput179), .A(n4712), .ZN(n4717) );
  AOI22_X1 U5253 ( .A1(IR_REG_9__SCAN_IN), .A2(keyinput204), .B1(
        IR_REG_10__SCAN_IN), .B2(keyinput196), .ZN(n4713) );
  OAI221_X1 U5254 ( .B1(IR_REG_9__SCAN_IN), .B2(keyinput204), .C1(
        IR_REG_10__SCAN_IN), .C2(keyinput196), .A(n4713), .ZN(n4716) );
  AOI22_X1 U5255 ( .A1(IR_REG_12__SCAN_IN), .A2(keyinput178), .B1(
        IR_REG_15__SCAN_IN), .B2(keyinput234), .ZN(n4714) );
  OAI221_X1 U5256 ( .B1(IR_REG_12__SCAN_IN), .B2(keyinput178), .C1(
        IR_REG_15__SCAN_IN), .C2(keyinput234), .A(n4714), .ZN(n4715) );
  NOR4_X1 U5257 ( .A1(n4718), .A2(n4717), .A3(n4716), .A4(n4715), .ZN(n4737)
         );
  AOI22_X1 U5258 ( .A1(IR_REG_19__SCAN_IN), .A2(keyinput155), .B1(
        IR_REG_22__SCAN_IN), .B2(keyinput252), .ZN(n4719) );
  OAI221_X1 U5259 ( .B1(IR_REG_19__SCAN_IN), .B2(keyinput155), .C1(
        IR_REG_22__SCAN_IN), .C2(keyinput252), .A(n4719), .ZN(n4726) );
  AOI22_X1 U5260 ( .A1(IR_REG_27__SCAN_IN), .A2(keyinput177), .B1(
        IR_REG_26__SCAN_IN), .B2(keyinput173), .ZN(n4720) );
  OAI221_X1 U5261 ( .B1(IR_REG_27__SCAN_IN), .B2(keyinput177), .C1(
        IR_REG_26__SCAN_IN), .C2(keyinput173), .A(n4720), .ZN(n4725) );
  AOI22_X1 U5262 ( .A1(IR_REG_28__SCAN_IN), .A2(keyinput232), .B1(
        D_REG_0__SCAN_IN), .B2(keyinput141), .ZN(n4721) );
  OAI221_X1 U5263 ( .B1(IR_REG_28__SCAN_IN), .B2(keyinput232), .C1(
        D_REG_0__SCAN_IN), .C2(keyinput141), .A(n4721), .ZN(n4724) );
  AOI22_X1 U5264 ( .A1(D_REG_2__SCAN_IN), .A2(keyinput215), .B1(
        D_REG_7__SCAN_IN), .B2(keyinput235), .ZN(n4722) );
  OAI221_X1 U5265 ( .B1(D_REG_2__SCAN_IN), .B2(keyinput215), .C1(
        D_REG_7__SCAN_IN), .C2(keyinput235), .A(n4722), .ZN(n4723) );
  NOR4_X1 U5266 ( .A1(n4726), .A2(n4725), .A3(n4724), .A4(n4723), .ZN(n4736)
         );
  AOI22_X1 U5267 ( .A1(D_REG_11__SCAN_IN), .A2(keyinput229), .B1(
        D_REG_6__SCAN_IN), .B2(keyinput160), .ZN(n4727) );
  OAI221_X1 U5268 ( .B1(D_REG_11__SCAN_IN), .B2(keyinput229), .C1(
        D_REG_6__SCAN_IN), .C2(keyinput160), .A(n4727), .ZN(n4734) );
  AOI22_X1 U5269 ( .A1(D_REG_14__SCAN_IN), .A2(keyinput153), .B1(
        D_REG_13__SCAN_IN), .B2(keyinput248), .ZN(n4728) );
  OAI221_X1 U5270 ( .B1(D_REG_14__SCAN_IN), .B2(keyinput153), .C1(
        D_REG_13__SCAN_IN), .C2(keyinput248), .A(n4728), .ZN(n4733) );
  AOI22_X1 U5271 ( .A1(D_REG_25__SCAN_IN), .A2(keyinput149), .B1(
        D_REG_19__SCAN_IN), .B2(keyinput244), .ZN(n4729) );
  OAI221_X1 U5272 ( .B1(D_REG_25__SCAN_IN), .B2(keyinput149), .C1(
        D_REG_19__SCAN_IN), .C2(keyinput244), .A(n4729), .ZN(n4732) );
  AOI22_X1 U5273 ( .A1(D_REG_31__SCAN_IN), .A2(keyinput225), .B1(
        D_REG_29__SCAN_IN), .B2(keyinput158), .ZN(n4730) );
  OAI221_X1 U5274 ( .B1(D_REG_31__SCAN_IN), .B2(keyinput225), .C1(
        D_REG_29__SCAN_IN), .C2(keyinput158), .A(n4730), .ZN(n4731) );
  NOR4_X1 U5275 ( .A1(n4734), .A2(n4733), .A3(n4732), .A4(n4731), .ZN(n4735)
         );
  NAND4_X1 U5276 ( .A1(n4738), .A2(n4737), .A3(n4736), .A4(n4735), .ZN(n4875)
         );
  AOI22_X1 U5277 ( .A1(REG0_REG_3__SCAN_IN), .A2(keyinput133), .B1(
        REG0_REG_17__SCAN_IN), .B2(keyinput190), .ZN(n4739) );
  OAI221_X1 U5278 ( .B1(REG0_REG_3__SCAN_IN), .B2(keyinput133), .C1(
        REG0_REG_17__SCAN_IN), .C2(keyinput190), .A(n4739), .ZN(n4746) );
  AOI22_X1 U5279 ( .A1(REG0_REG_21__SCAN_IN), .A2(keyinput236), .B1(
        REG0_REG_25__SCAN_IN), .B2(keyinput200), .ZN(n4740) );
  OAI221_X1 U5280 ( .B1(REG0_REG_21__SCAN_IN), .B2(keyinput236), .C1(
        REG0_REG_25__SCAN_IN), .C2(keyinput200), .A(n4740), .ZN(n4745) );
  AOI22_X1 U5281 ( .A1(REG1_REG_6__SCAN_IN), .A2(keyinput254), .B1(
        REG1_REG_10__SCAN_IN), .B2(keyinput221), .ZN(n4741) );
  OAI221_X1 U5282 ( .B1(REG1_REG_6__SCAN_IN), .B2(keyinput254), .C1(
        REG1_REG_10__SCAN_IN), .C2(keyinput221), .A(n4741), .ZN(n4744) );
  AOI22_X1 U5283 ( .A1(REG1_REG_15__SCAN_IN), .A2(keyinput245), .B1(
        REG1_REG_12__SCAN_IN), .B2(keyinput175), .ZN(n4742) );
  OAI221_X1 U5284 ( .B1(REG1_REG_15__SCAN_IN), .B2(keyinput245), .C1(
        REG1_REG_12__SCAN_IN), .C2(keyinput175), .A(n4742), .ZN(n4743) );
  NOR4_X1 U5285 ( .A1(n4746), .A2(n4745), .A3(n4744), .A4(n4743), .ZN(n4774)
         );
  AOI22_X1 U5286 ( .A1(REG1_REG_18__SCAN_IN), .A2(keyinput191), .B1(
        REG1_REG_20__SCAN_IN), .B2(keyinput241), .ZN(n4747) );
  OAI221_X1 U5287 ( .B1(REG1_REG_18__SCAN_IN), .B2(keyinput191), .C1(
        REG1_REG_20__SCAN_IN), .C2(keyinput241), .A(n4747), .ZN(n4754) );
  AOI22_X1 U5288 ( .A1(REG1_REG_24__SCAN_IN), .A2(keyinput217), .B1(
        REG1_REG_23__SCAN_IN), .B2(keyinput139), .ZN(n4748) );
  OAI221_X1 U5289 ( .B1(REG1_REG_24__SCAN_IN), .B2(keyinput217), .C1(
        REG1_REG_23__SCAN_IN), .C2(keyinput139), .A(n4748), .ZN(n4753) );
  AOI22_X1 U5290 ( .A1(REG1_REG_30__SCAN_IN), .A2(keyinput172), .B1(
        REG2_REG_9__SCAN_IN), .B2(keyinput216), .ZN(n4749) );
  OAI221_X1 U5291 ( .B1(REG1_REG_30__SCAN_IN), .B2(keyinput172), .C1(
        REG2_REG_9__SCAN_IN), .C2(keyinput216), .A(n4749), .ZN(n4752) );
  AOI22_X1 U5292 ( .A1(REG2_REG_11__SCAN_IN), .A2(keyinput176), .B1(
        REG2_REG_10__SCAN_IN), .B2(keyinput210), .ZN(n4750) );
  OAI221_X1 U5293 ( .B1(REG2_REG_11__SCAN_IN), .B2(keyinput176), .C1(
        REG2_REG_10__SCAN_IN), .C2(keyinput210), .A(n4750), .ZN(n4751) );
  NOR4_X1 U5294 ( .A1(n4754), .A2(n4753), .A3(n4752), .A4(n4751), .ZN(n4773)
         );
  AOI22_X1 U5295 ( .A1(REG2_REG_18__SCAN_IN), .A2(keyinput197), .B1(
        REG2_REG_14__SCAN_IN), .B2(keyinput128), .ZN(n4755) );
  OAI221_X1 U5296 ( .B1(REG2_REG_18__SCAN_IN), .B2(keyinput197), .C1(
        REG2_REG_14__SCAN_IN), .C2(keyinput128), .A(n4755), .ZN(n4762) );
  AOI22_X1 U5297 ( .A1(REG2_REG_20__SCAN_IN), .A2(keyinput212), .B1(
        REG2_REG_27__SCAN_IN), .B2(keyinput255), .ZN(n4756) );
  OAI221_X1 U5298 ( .B1(REG2_REG_20__SCAN_IN), .B2(keyinput212), .C1(
        REG2_REG_27__SCAN_IN), .C2(keyinput255), .A(n4756), .ZN(n4761) );
  AOI22_X1 U5299 ( .A1(ADDR_REG_17__SCAN_IN), .A2(keyinput165), .B1(
        REG2_REG_29__SCAN_IN), .B2(keyinput180), .ZN(n4757) );
  OAI221_X1 U5300 ( .B1(ADDR_REG_17__SCAN_IN), .B2(keyinput165), .C1(
        REG2_REG_29__SCAN_IN), .C2(keyinput180), .A(n4757), .ZN(n4760) );
  AOI22_X1 U5301 ( .A1(ADDR_REG_15__SCAN_IN), .A2(keyinput220), .B1(
        ADDR_REG_13__SCAN_IN), .B2(keyinput227), .ZN(n4758) );
  OAI221_X1 U5302 ( .B1(ADDR_REG_15__SCAN_IN), .B2(keyinput220), .C1(
        ADDR_REG_13__SCAN_IN), .C2(keyinput227), .A(n4758), .ZN(n4759) );
  NOR4_X1 U5303 ( .A1(n4762), .A2(n4761), .A3(n4760), .A4(n4759), .ZN(n4772)
         );
  AOI22_X1 U5304 ( .A1(ADDR_REG_6__SCAN_IN), .A2(keyinput187), .B1(
        ADDR_REG_4__SCAN_IN), .B2(keyinput130), .ZN(n4763) );
  OAI221_X1 U5305 ( .B1(ADDR_REG_6__SCAN_IN), .B2(keyinput187), .C1(
        ADDR_REG_4__SCAN_IN), .C2(keyinput130), .A(n4763), .ZN(n4770) );
  AOI22_X1 U5306 ( .A1(DATAO_REG_2__SCAN_IN), .A2(keyinput181), .B1(
        DATAO_REG_0__SCAN_IN), .B2(keyinput222), .ZN(n4764) );
  OAI221_X1 U5307 ( .B1(DATAO_REG_2__SCAN_IN), .B2(keyinput181), .C1(
        DATAO_REG_0__SCAN_IN), .C2(keyinput222), .A(n4764), .ZN(n4769) );
  AOI22_X1 U5308 ( .A1(DATAO_REG_6__SCAN_IN), .A2(keyinput182), .B1(
        DATAO_REG_5__SCAN_IN), .B2(keyinput167), .ZN(n4765) );
  OAI221_X1 U5309 ( .B1(DATAO_REG_6__SCAN_IN), .B2(keyinput182), .C1(
        DATAO_REG_5__SCAN_IN), .C2(keyinput167), .A(n4765), .ZN(n4768) );
  AOI22_X1 U5310 ( .A1(DATAO_REG_13__SCAN_IN), .A2(keyinput202), .B1(
        DATAO_REG_8__SCAN_IN), .B2(keyinput219), .ZN(n4766) );
  OAI221_X1 U5311 ( .B1(DATAO_REG_13__SCAN_IN), .B2(keyinput202), .C1(
        DATAO_REG_8__SCAN_IN), .C2(keyinput219), .A(n4766), .ZN(n4767) );
  NOR4_X1 U5312 ( .A1(n4770), .A2(n4769), .A3(n4768), .A4(n4767), .ZN(n4771)
         );
  NAND4_X1 U5313 ( .A1(n4774), .A2(n4773), .A3(n4772), .A4(n4771), .ZN(n4874)
         );
  AOI22_X1 U5314 ( .A1(DATAO_REG_18__SCAN_IN), .A2(keyinput143), .B1(
        DATAO_REG_16__SCAN_IN), .B2(keyinput135), .ZN(n4775) );
  OAI221_X1 U5315 ( .B1(DATAO_REG_18__SCAN_IN), .B2(keyinput143), .C1(
        DATAO_REG_16__SCAN_IN), .C2(keyinput135), .A(n4775), .ZN(n4782) );
  AOI22_X1 U5316 ( .A1(DATAO_REG_27__SCAN_IN), .A2(keyinput147), .B1(
        DATAO_REG_20__SCAN_IN), .B2(keyinput250), .ZN(n4776) );
  OAI221_X1 U5317 ( .B1(DATAO_REG_27__SCAN_IN), .B2(keyinput147), .C1(
        DATAO_REG_20__SCAN_IN), .C2(keyinput250), .A(n4776), .ZN(n4781) );
  AOI22_X1 U5318 ( .A1(REG3_REG_11__SCAN_IN), .A2(keyinput183), .B1(
        REG3_REG_22__SCAN_IN), .B2(keyinput169), .ZN(n4777) );
  OAI221_X1 U5319 ( .B1(REG3_REG_11__SCAN_IN), .B2(keyinput183), .C1(
        REG3_REG_22__SCAN_IN), .C2(keyinput169), .A(n4777), .ZN(n4780) );
  AOI22_X1 U5320 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput195), .B1(
        IR_REG_2__SCAN_IN), .B2(keyinput137), .ZN(n4778) );
  OAI221_X1 U5321 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput195), .C1(
        IR_REG_2__SCAN_IN), .C2(keyinput137), .A(n4778), .ZN(n4779) );
  NOR4_X1 U5322 ( .A1(n4782), .A2(n4781), .A3(n4780), .A4(n4779), .ZN(n4820)
         );
  AOI22_X1 U5323 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput134), .B1(n4784), 
        .B2(keyinput199), .ZN(n4783) );
  OAI221_X1 U5324 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput134), .C1(n4784), 
        .C2(keyinput199), .A(n4783), .ZN(n4794) );
  INV_X1 U5325 ( .A(DATAI_9_), .ZN(n4922) );
  AOI22_X1 U5326 ( .A1(n4906), .A2(keyinput168), .B1(keyinput251), .B2(n4922), 
        .ZN(n4785) );
  OAI221_X1 U5327 ( .B1(n4906), .B2(keyinput168), .C1(n4922), .C2(keyinput251), 
        .A(n4785), .ZN(n4793) );
  INV_X1 U5328 ( .A(DATAI_7_), .ZN(n4787) );
  AOI22_X1 U5329 ( .A1(n4788), .A2(keyinput253), .B1(keyinput185), .B2(n4787), 
        .ZN(n4786) );
  OAI221_X1 U5330 ( .B1(n4788), .B2(keyinput253), .C1(n4787), .C2(keyinput185), 
        .A(n4786), .ZN(n4792) );
  AOI22_X1 U5331 ( .A1(n4790), .A2(keyinput166), .B1(keyinput206), .B2(n3618), 
        .ZN(n4789) );
  OAI221_X1 U5332 ( .B1(n4790), .B2(keyinput166), .C1(n3618), .C2(keyinput206), 
        .A(n4789), .ZN(n4791) );
  NOR4_X1 U5333 ( .A1(n4794), .A2(n4793), .A3(n4792), .A4(n4791), .ZN(n4819)
         );
  AOI22_X1 U5334 ( .A1(n5047), .A2(keyinput238), .B1(keyinput231), .B2(n5045), 
        .ZN(n4795) );
  OAI221_X1 U5335 ( .B1(n5047), .B2(keyinput238), .C1(n5045), .C2(keyinput231), 
        .A(n4795), .ZN(n4804) );
  INV_X1 U5336 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4797) );
  AOI22_X1 U5337 ( .A1(n4797), .A2(keyinput164), .B1(n4984), .B2(keyinput140), 
        .ZN(n4796) );
  OAI221_X1 U5338 ( .B1(n4797), .B2(keyinput164), .C1(n4984), .C2(keyinput140), 
        .A(n4796), .ZN(n4803) );
  XNOR2_X1 U5339 ( .A(IR_REG_1__SCAN_IN), .B(keyinput157), .ZN(n4801) );
  XNOR2_X1 U5340 ( .A(IR_REG_3__SCAN_IN), .B(keyinput151), .ZN(n4800) );
  XNOR2_X1 U5341 ( .A(IR_REG_11__SCAN_IN), .B(keyinput208), .ZN(n4799) );
  XNOR2_X1 U5342 ( .A(IR_REG_7__SCAN_IN), .B(keyinput203), .ZN(n4798) );
  NAND4_X1 U5343 ( .A1(n4801), .A2(n4800), .A3(n4799), .A4(n4798), .ZN(n4802)
         );
  NOR3_X1 U5344 ( .A1(n4804), .A2(n4803), .A3(n4802), .ZN(n4818) );
  XOR2_X1 U5345 ( .A(IR_REG_25__SCAN_IN), .B(keyinput228), .Z(n4810) );
  XOR2_X1 U5346 ( .A(IR_REG_21__SCAN_IN), .B(keyinput240), .Z(n4809) );
  XNOR2_X1 U5347 ( .A(n4805), .B(keyinput132), .ZN(n4808) );
  XNOR2_X1 U5348 ( .A(n4806), .B(keyinput242), .ZN(n4807) );
  NOR4_X1 U5349 ( .A1(n4810), .A2(n4809), .A3(n4808), .A4(n4807), .ZN(n4814)
         );
  XOR2_X1 U5350 ( .A(n2743), .B(keyinput211), .Z(n4813) );
  XNOR2_X1 U5351 ( .A(IR_REG_14__SCAN_IN), .B(keyinput207), .ZN(n4812) );
  XNOR2_X1 U5352 ( .A(IR_REG_17__SCAN_IN), .B(keyinput209), .ZN(n4811) );
  NAND4_X1 U5353 ( .A1(n4814), .A2(n4813), .A3(n4812), .A4(n4811), .ZN(n4816)
         );
  XNOR2_X1 U5354 ( .A(n4934), .B(keyinput184), .ZN(n4815) );
  NOR2_X1 U5355 ( .A1(n4816), .A2(n4815), .ZN(n4817) );
  NAND4_X1 U5356 ( .A1(n4820), .A2(n4819), .A3(n4818), .A4(n4817), .ZN(n4873)
         );
  AOI22_X1 U5357 ( .A1(n4940), .A2(keyinput156), .B1(n4822), .B2(keyinput129), 
        .ZN(n4821) );
  OAI221_X1 U5358 ( .B1(n4940), .B2(keyinput156), .C1(n4822), .C2(keyinput129), 
        .A(n4821), .ZN(n4833) );
  AOI22_X1 U5359 ( .A1(n4936), .A2(keyinput214), .B1(n4824), .B2(keyinput171), 
        .ZN(n4823) );
  OAI221_X1 U5360 ( .B1(n4936), .B2(keyinput214), .C1(n4824), .C2(keyinput171), 
        .A(n4823), .ZN(n4832) );
  INV_X1 U5361 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4827) );
  AOI22_X1 U5362 ( .A1(n4827), .A2(keyinput223), .B1(n4826), .B2(keyinput142), 
        .ZN(n4825) );
  OAI221_X1 U5363 ( .B1(n4827), .B2(keyinput223), .C1(n4826), .C2(keyinput142), 
        .A(n4825), .ZN(n4831) );
  AOI22_X1 U5364 ( .A1(n4829), .A2(keyinput213), .B1(keyinput198), .B2(n4963), 
        .ZN(n4828) );
  OAI221_X1 U5365 ( .B1(n4829), .B2(keyinput213), .C1(n4963), .C2(keyinput198), 
        .A(n4828), .ZN(n4830) );
  NOR4_X1 U5366 ( .A1(n4833), .A2(n4832), .A3(n4831), .A4(n4830), .ZN(n4871)
         );
  INV_X1 U5367 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4902) );
  AOI22_X1 U5368 ( .A1(n4902), .A2(keyinput154), .B1(n4470), .B2(keyinput159), 
        .ZN(n4834) );
  OAI221_X1 U5369 ( .B1(n4902), .B2(keyinput154), .C1(n4470), .C2(keyinput159), 
        .A(n4834), .ZN(n4843) );
  INV_X1 U5370 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4836) );
  AOI22_X1 U5371 ( .A1(n4836), .A2(keyinput144), .B1(keyinput205), .B2(n4917), 
        .ZN(n4835) );
  OAI221_X1 U5372 ( .B1(n4836), .B2(keyinput144), .C1(n4917), .C2(keyinput205), 
        .A(n4835), .ZN(n4842) );
  INV_X1 U5373 ( .A(REG1_REG_3__SCAN_IN), .ZN(n5043) );
  AOI22_X1 U5374 ( .A1(n4427), .A2(keyinput138), .B1(keyinput233), .B2(n5043), 
        .ZN(n4837) );
  OAI221_X1 U5375 ( .B1(n4427), .B2(keyinput138), .C1(n5043), .C2(keyinput233), 
        .A(n4837), .ZN(n4841) );
  AOI22_X1 U5376 ( .A1(n4920), .A2(keyinput186), .B1(n4839), .B2(keyinput170), 
        .ZN(n4838) );
  OAI221_X1 U5377 ( .B1(n4920), .B2(keyinput186), .C1(n4839), .C2(keyinput170), 
        .A(n4838), .ZN(n4840) );
  NOR4_X1 U5378 ( .A1(n4843), .A2(n4842), .A3(n4841), .A4(n4840), .ZN(n4870)
         );
  INV_X1 U5379 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4845) );
  AOI22_X1 U5380 ( .A1(n4846), .A2(keyinput218), .B1(n4845), .B2(keyinput224), 
        .ZN(n4844) );
  OAI221_X1 U5381 ( .B1(n4846), .B2(keyinput218), .C1(n4845), .C2(keyinput224), 
        .A(n4844), .ZN(n4854) );
  INV_X1 U5382 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4848) );
  AOI22_X1 U5383 ( .A1(n4848), .A2(keyinput239), .B1(keyinput194), .B2(n3271), 
        .ZN(n4847) );
  OAI221_X1 U5384 ( .B1(n4848), .B2(keyinput239), .C1(n3271), .C2(keyinput194), 
        .A(n4847), .ZN(n4853) );
  AOI22_X1 U5385 ( .A1(n3342), .A2(keyinput189), .B1(n2528), .B2(keyinput131), 
        .ZN(n4849) );
  OAI221_X1 U5386 ( .B1(n3342), .B2(keyinput189), .C1(n2528), .C2(keyinput131), 
        .A(n4849), .ZN(n4852) );
  AOI22_X1 U5387 ( .A1(n4102), .A2(keyinput174), .B1(keyinput146), .B2(n2622), 
        .ZN(n4850) );
  OAI221_X1 U5388 ( .B1(n4102), .B2(keyinput174), .C1(n2622), .C2(keyinput146), 
        .A(n4850), .ZN(n4851) );
  NOR4_X1 U5389 ( .A1(n4854), .A2(n4853), .A3(n4852), .A4(n4851), .ZN(n4869)
         );
  AOI22_X1 U5390 ( .A1(n4857), .A2(keyinput188), .B1(keyinput243), .B2(n4856), 
        .ZN(n4855) );
  OAI221_X1 U5391 ( .B1(n4857), .B2(keyinput188), .C1(n4856), .C2(keyinput243), 
        .A(n4855), .ZN(n4867) );
  INV_X1 U5392 ( .A(ADDR_REG_18__SCAN_IN), .ZN(n4949) );
  INV_X1 U5393 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n4880) );
  AOI22_X1 U5394 ( .A1(n4949), .A2(keyinput162), .B1(keyinput249), .B2(n4880), 
        .ZN(n4858) );
  OAI221_X1 U5395 ( .B1(n4949), .B2(keyinput162), .C1(n4880), .C2(keyinput249), 
        .A(n4858), .ZN(n4866) );
  INV_X1 U5396 ( .A(ADDR_REG_10__SCAN_IN), .ZN(n4861) );
  INV_X1 U5397 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n4860) );
  AOI22_X1 U5398 ( .A1(n4861), .A2(keyinput163), .B1(keyinput193), .B2(n4860), 
        .ZN(n4859) );
  OAI221_X1 U5399 ( .B1(n4861), .B2(keyinput163), .C1(n4860), .C2(keyinput193), 
        .A(n4859), .ZN(n4865) );
  XNOR2_X1 U5400 ( .A(REG3_REG_18__SCAN_IN), .B(keyinput246), .ZN(n4863) );
  XNOR2_X1 U5401 ( .A(IR_REG_30__SCAN_IN), .B(keyinput145), .ZN(n4862) );
  NAND2_X1 U5402 ( .A1(n4863), .A2(n4862), .ZN(n4864) );
  NOR4_X1 U5403 ( .A1(n4867), .A2(n4866), .A3(n4865), .A4(n4864), .ZN(n4868)
         );
  NAND4_X1 U5404 ( .A1(n4871), .A2(n4870), .A3(n4869), .A4(n4868), .ZN(n4872)
         );
  NOR4_X1 U5405 ( .A1(n4875), .A2(n4874), .A3(n4873), .A4(n4872), .ZN(n5075)
         );
  INV_X1 U5406 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4878) );
  AOI22_X1 U5407 ( .A1(n4878), .A2(keyinput2), .B1(n4877), .B2(keyinput126), 
        .ZN(n4876) );
  OAI221_X1 U5408 ( .B1(n4878), .B2(keyinput2), .C1(n4877), .C2(keyinput126), 
        .A(n4876), .ZN(n4889) );
  INV_X1 U5409 ( .A(ADDR_REG_6__SCAN_IN), .ZN(n4881) );
  AOI22_X1 U5410 ( .A1(n4881), .A2(keyinput59), .B1(keyinput121), .B2(n4880), 
        .ZN(n4879) );
  OAI221_X1 U5411 ( .B1(n4881), .B2(keyinput59), .C1(n4880), .C2(keyinput121), 
        .A(n4879), .ZN(n4888) );
  INV_X1 U5412 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4884) );
  INV_X1 U5413 ( .A(ADDR_REG_17__SCAN_IN), .ZN(n4883) );
  AOI22_X1 U5414 ( .A1(n4884), .A2(keyinput99), .B1(n4883), .B2(keyinput37), 
        .ZN(n4882) );
  OAI221_X1 U5415 ( .B1(n4884), .B2(keyinput99), .C1(n4883), .C2(keyinput37), 
        .A(n4882), .ZN(n4887) );
  AOI22_X1 U5416 ( .A1(n3271), .A2(keyinput66), .B1(n3342), .B2(keyinput61), 
        .ZN(n4885) );
  OAI221_X1 U5417 ( .B1(n3271), .B2(keyinput66), .C1(n3342), .C2(keyinput61), 
        .A(n4885), .ZN(n4886) );
  NOR4_X1 U5418 ( .A1(n4889), .A2(n4888), .A3(n4887), .A4(n4886), .ZN(n4931)
         );
  AOI22_X1 U5419 ( .A1(n3335), .A2(keyinput48), .B1(keyinput117), .B2(n4891), 
        .ZN(n4890) );
  OAI221_X1 U5420 ( .B1(n3335), .B2(keyinput48), .C1(n4891), .C2(keyinput117), 
        .A(n4890), .ZN(n4900) );
  INV_X1 U5421 ( .A(DATAI_15_), .ZN(n4893) );
  AOI22_X1 U5422 ( .A1(n4893), .A2(keyinput98), .B1(n4278), .B2(keyinput0), 
        .ZN(n4892) );
  OAI221_X1 U5423 ( .B1(n4893), .B2(keyinput98), .C1(n4278), .C2(keyinput0), 
        .A(n4892), .ZN(n4899) );
  XNOR2_X1 U5424 ( .A(IR_REG_17__SCAN_IN), .B(keyinput81), .ZN(n4897) );
  XNOR2_X1 U5425 ( .A(IR_REG_18__SCAN_IN), .B(keyinput4), .ZN(n4896) );
  XNOR2_X1 U5426 ( .A(IR_REG_16__SCAN_IN), .B(keyinput114), .ZN(n4895) );
  XNOR2_X1 U5427 ( .A(IR_REG_15__SCAN_IN), .B(keyinput106), .ZN(n4894) );
  NAND4_X1 U5428 ( .A1(n4897), .A2(n4896), .A3(n4895), .A4(n4894), .ZN(n4898)
         );
  NOR3_X1 U5429 ( .A1(n4900), .A2(n4899), .A3(n4898), .ZN(n4930) );
  INV_X1 U5430 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4903) );
  AOI22_X1 U5431 ( .A1(n4903), .A2(keyinput47), .B1(n4902), .B2(keyinput26), 
        .ZN(n4901) );
  OAI221_X1 U5432 ( .B1(n4903), .B2(keyinput47), .C1(n4902), .C2(keyinput26), 
        .A(n4901), .ZN(n4913) );
  AOI22_X1 U5433 ( .A1(n4470), .A2(keyinput31), .B1(n4905), .B2(keyinput6), 
        .ZN(n4904) );
  OAI221_X1 U5434 ( .B1(n4470), .B2(keyinput31), .C1(n4905), .C2(keyinput6), 
        .A(n4904), .ZN(n4912) );
  XOR2_X1 U5435 ( .A(n4906), .B(keyinput40), .Z(n4910) );
  XNOR2_X1 U5436 ( .A(IR_REG_14__SCAN_IN), .B(keyinput79), .ZN(n4909) );
  XNOR2_X1 U5437 ( .A(REG1_REG_14__SCAN_IN), .B(keyinput96), .ZN(n4908) );
  XNOR2_X1 U5438 ( .A(IR_REG_11__SCAN_IN), .B(keyinput80), .ZN(n4907) );
  NAND4_X1 U5439 ( .A1(n4910), .A2(n4909), .A3(n4908), .A4(n4907), .ZN(n4911)
         );
  NOR3_X1 U5440 ( .A1(n4913), .A2(n4912), .A3(n4911), .ZN(n4929) );
  INV_X1 U5441 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4915) );
  AOI22_X1 U5442 ( .A1(n4915), .A2(keyinput113), .B1(n4344), .B2(keyinput11), 
        .ZN(n4914) );
  OAI221_X1 U5443 ( .B1(n4915), .B2(keyinput113), .C1(n4344), .C2(keyinput11), 
        .A(n4914), .ZN(n4927) );
  AOI22_X1 U5444 ( .A1(n4918), .A2(keyinput89), .B1(n4917), .B2(keyinput77), 
        .ZN(n4916) );
  OAI221_X1 U5445 ( .B1(n4918), .B2(keyinput89), .C1(n4917), .C2(keyinput77), 
        .A(n4916), .ZN(n4926) );
  AOI22_X1 U5446 ( .A1(n4435), .A2(keyinput72), .B1(keyinput58), .B2(n4920), 
        .ZN(n4919) );
  OAI221_X1 U5447 ( .B1(n4435), .B2(keyinput72), .C1(n4920), .C2(keyinput58), 
        .A(n4919), .ZN(n4925) );
  AOI22_X1 U5448 ( .A1(n4923), .A2(keyinput122), .B1(n4922), .B2(keyinput123), 
        .ZN(n4921) );
  OAI221_X1 U5449 ( .B1(n4923), .B2(keyinput122), .C1(n4922), .C2(keyinput123), 
        .A(n4921), .ZN(n4924) );
  NOR4_X1 U5450 ( .A1(n4927), .A2(n4926), .A3(n4925), .A4(n4924), .ZN(n4928)
         );
  NAND4_X1 U5451 ( .A1(n4931), .A2(n4930), .A3(n4929), .A4(n4928), .ZN(n5074)
         );
  AOI22_X1 U5452 ( .A1(n4934), .A2(keyinput56), .B1(keyinput32), .B2(n4933), 
        .ZN(n4932) );
  OAI221_X1 U5453 ( .B1(n4934), .B2(keyinput56), .C1(n4933), .C2(keyinput32), 
        .A(n4932), .ZN(n4946) );
  AOI22_X1 U5454 ( .A1(n4937), .A2(keyinput94), .B1(n4936), .B2(keyinput86), 
        .ZN(n4935) );
  OAI221_X1 U5455 ( .B1(n4937), .B2(keyinput94), .C1(n4936), .C2(keyinput86), 
        .A(n4935), .ZN(n4945) );
  AOI22_X1 U5456 ( .A1(n4940), .A2(keyinput28), .B1(keyinput24), .B2(n4939), 
        .ZN(n4938) );
  OAI221_X1 U5457 ( .B1(n4940), .B2(keyinput28), .C1(n4939), .C2(keyinput24), 
        .A(n4938), .ZN(n4944) );
  XNOR2_X1 U5458 ( .A(IR_REG_22__SCAN_IN), .B(keyinput124), .ZN(n4942) );
  XNOR2_X1 U5459 ( .A(IR_REG_21__SCAN_IN), .B(keyinput112), .ZN(n4941) );
  NAND2_X1 U5460 ( .A1(n4942), .A2(n4941), .ZN(n4943) );
  NOR4_X1 U5461 ( .A1(n4946), .A2(n4945), .A3(n4944), .A4(n4943), .ZN(n4993)
         );
  AOI22_X1 U5462 ( .A1(n4949), .A2(keyinput34), .B1(keyinput7), .B2(n4948), 
        .ZN(n4947) );
  OAI221_X1 U5463 ( .B1(n4949), .B2(keyinput34), .C1(n4948), .C2(keyinput7), 
        .A(n4947), .ZN(n4961) );
  AOI22_X1 U5464 ( .A1(n4952), .A2(keyinput30), .B1(keyinput39), .B2(n4951), 
        .ZN(n4950) );
  OAI221_X1 U5465 ( .B1(n4952), .B2(keyinput30), .C1(n4951), .C2(keyinput39), 
        .A(n4950), .ZN(n4960) );
  XOR2_X1 U5466 ( .A(n4953), .B(keyinput64), .Z(n4956) );
  XNOR2_X1 U5467 ( .A(IR_REG_25__SCAN_IN), .B(keyinput100), .ZN(n4955) );
  XNOR2_X1 U5468 ( .A(IR_REG_28__SCAN_IN), .B(keyinput104), .ZN(n4954) );
  NAND3_X1 U5469 ( .A1(n4956), .A2(n4955), .A3(n4954), .ZN(n4959) );
  XNOR2_X1 U5470 ( .A(n4957), .B(keyinput116), .ZN(n4958) );
  NOR4_X1 U5471 ( .A1(n4961), .A2(n4960), .A3(n4959), .A4(n4958), .ZN(n4992)
         );
  AOI22_X1 U5472 ( .A1(n4964), .A2(keyinput75), .B1(keyinput70), .B2(n4963), 
        .ZN(n4962) );
  OAI221_X1 U5473 ( .B1(n4964), .B2(keyinput75), .C1(n4963), .C2(keyinput70), 
        .A(n4962), .ZN(n4975) );
  XOR2_X1 U5474 ( .A(DATAI_2_), .B(keyinput8), .Z(n4967) );
  XNOR2_X1 U5475 ( .A(n4965), .B(keyinput55), .ZN(n4966) );
  NOR2_X1 U5476 ( .A1(n4967), .A2(n4966), .ZN(n4971) );
  XNOR2_X1 U5477 ( .A(keyinput14), .B(REG0_REG_8__SCAN_IN), .ZN(n4970) );
  XNOR2_X1 U5478 ( .A(IR_REG_5__SCAN_IN), .B(keyinput51), .ZN(n4969) );
  XNOR2_X1 U5479 ( .A(IR_REG_3__SCAN_IN), .B(keyinput23), .ZN(n4968) );
  NAND4_X1 U5480 ( .A1(n4971), .A2(n4970), .A3(n4969), .A4(n4968), .ZN(n4974)
         );
  XNOR2_X1 U5481 ( .A(n4972), .B(keyinput54), .ZN(n4973) );
  NOR3_X1 U5482 ( .A1(n4975), .A2(n4974), .A3(n4973), .ZN(n4991) );
  AOI22_X1 U5483 ( .A1(n4977), .A2(keyinput101), .B1(n2367), .B2(keyinput45), 
        .ZN(n4976) );
  OAI221_X1 U5484 ( .B1(n4977), .B2(keyinput101), .C1(n2367), .C2(keyinput45), 
        .A(n4976), .ZN(n4981) );
  XNOR2_X1 U5485 ( .A(n4978), .B(keyinput21), .ZN(n4980) );
  XOR2_X1 U5486 ( .A(IR_REG_1__SCAN_IN), .B(keyinput29), .Z(n4979) );
  OR3_X1 U5487 ( .A1(n4981), .A2(n4980), .A3(n4979), .ZN(n4989) );
  AOI22_X1 U5488 ( .A1(n4984), .A2(keyinput12), .B1(n4983), .B2(keyinput97), 
        .ZN(n4982) );
  OAI221_X1 U5489 ( .B1(n4984), .B2(keyinput12), .C1(n4983), .C2(keyinput97), 
        .A(n4982), .ZN(n4988) );
  AOI22_X1 U5490 ( .A1(n4986), .A2(keyinput25), .B1(n2766), .B2(keyinput13), 
        .ZN(n4985) );
  OAI221_X1 U5491 ( .B1(n4986), .B2(keyinput25), .C1(n2766), .C2(keyinput13), 
        .A(n4985), .ZN(n4987) );
  NOR3_X1 U5492 ( .A1(n4989), .A2(n4988), .A3(n4987), .ZN(n4990) );
  NAND4_X1 U5493 ( .A1(n4993), .A2(n4992), .A3(n4991), .A4(n4990), .ZN(n5073)
         );
  AOI22_X1 U5494 ( .A1(REG3_REG_21__SCAN_IN), .A2(keyinput38), .B1(
        REG3_REG_22__SCAN_IN), .B2(keyinput41), .ZN(n4994) );
  OAI221_X1 U5495 ( .B1(REG3_REG_21__SCAN_IN), .B2(keyinput38), .C1(
        REG3_REG_22__SCAN_IN), .C2(keyinput41), .A(n4994), .ZN(n5001) );
  AOI22_X1 U5496 ( .A1(DATAO_REG_13__SCAN_IN), .A2(keyinput74), .B1(
        REG3_REG_27__SCAN_IN), .B2(keyinput67), .ZN(n4995) );
  OAI221_X1 U5497 ( .B1(DATAO_REG_13__SCAN_IN), .B2(keyinput74), .C1(
        REG3_REG_27__SCAN_IN), .C2(keyinput67), .A(n4995), .ZN(n5000) );
  AOI22_X1 U5498 ( .A1(REG1_REG_30__SCAN_IN), .A2(keyinput44), .B1(
        REG2_REG_20__SCAN_IN), .B2(keyinput84), .ZN(n4996) );
  OAI221_X1 U5499 ( .B1(REG1_REG_30__SCAN_IN), .B2(keyinput44), .C1(
        REG2_REG_20__SCAN_IN), .C2(keyinput84), .A(n4996), .ZN(n4999) );
  AOI22_X1 U5500 ( .A1(REG2_REG_23__SCAN_IN), .A2(keyinput46), .B1(
        REG3_REG_18__SCAN_IN), .B2(keyinput118), .ZN(n4997) );
  OAI221_X1 U5501 ( .B1(REG2_REG_23__SCAN_IN), .B2(keyinput46), .C1(
        REG3_REG_18__SCAN_IN), .C2(keyinput118), .A(n4997), .ZN(n4998) );
  NOR4_X1 U5502 ( .A1(n5001), .A2(n5000), .A3(n4999), .A4(n4998), .ZN(n5071)
         );
  AOI22_X1 U5503 ( .A1(REG2_REG_17__SCAN_IN), .A2(keyinput3), .B1(
        REG2_REG_27__SCAN_IN), .B2(keyinput127), .ZN(n5002) );
  OAI221_X1 U5504 ( .B1(REG2_REG_17__SCAN_IN), .B2(keyinput3), .C1(
        REG2_REG_27__SCAN_IN), .C2(keyinput127), .A(n5002), .ZN(n5009) );
  AOI22_X1 U5505 ( .A1(REG1_REG_18__SCAN_IN), .A2(keyinput63), .B1(DATAI_4_), 
        .B2(keyinput73), .ZN(n5003) );
  OAI221_X1 U5506 ( .B1(REG1_REG_18__SCAN_IN), .B2(keyinput63), .C1(DATAI_4_), 
        .C2(keyinput73), .A(n5003), .ZN(n5008) );
  AOI22_X1 U5507 ( .A1(DATAO_REG_8__SCAN_IN), .A2(keyinput91), .B1(
        DATAO_REG_2__SCAN_IN), .B2(keyinput53), .ZN(n5004) );
  OAI221_X1 U5508 ( .B1(DATAO_REG_8__SCAN_IN), .B2(keyinput91), .C1(
        DATAO_REG_2__SCAN_IN), .C2(keyinput53), .A(n5004), .ZN(n5007) );
  AOI22_X1 U5509 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput33), .B1(DATAI_19_), 
        .B2(keyinput109), .ZN(n5005) );
  OAI221_X1 U5510 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput33), .C1(DATAI_19_), 
        .C2(keyinput109), .A(n5005), .ZN(n5006) );
  NOR4_X1 U5511 ( .A1(n5009), .A2(n5008), .A3(n5007), .A4(n5006), .ZN(n5070)
         );
  OAI22_X1 U5512 ( .A1(D_REG_13__SCAN_IN), .A2(keyinput120), .B1(keyinput90), 
        .B2(REG1_REG_11__SCAN_IN), .ZN(n5010) );
  AOI221_X1 U5513 ( .B1(D_REG_13__SCAN_IN), .B2(keyinput120), .C1(
        REG1_REG_11__SCAN_IN), .C2(keyinput90), .A(n5010), .ZN(n5017) );
  OAI22_X1 U5514 ( .A1(IR_REG_27__SCAN_IN), .A2(keyinput49), .B1(keyinput88), 
        .B2(REG2_REG_9__SCAN_IN), .ZN(n5011) );
  AOI221_X1 U5515 ( .B1(IR_REG_27__SCAN_IN), .B2(keyinput49), .C1(
        REG2_REG_9__SCAN_IN), .C2(keyinput88), .A(n5011), .ZN(n5016) );
  OAI22_X1 U5516 ( .A1(DATAI_14_), .A2(keyinput102), .B1(DATAI_10_), .B2(
        keyinput22), .ZN(n5012) );
  AOI221_X1 U5517 ( .B1(DATAI_14_), .B2(keyinput102), .C1(keyinput22), .C2(
        DATAI_10_), .A(n5012), .ZN(n5015) );
  OAI22_X1 U5518 ( .A1(D_REG_7__SCAN_IN), .A2(keyinput107), .B1(
        D_REG_2__SCAN_IN), .B2(keyinput87), .ZN(n5013) );
  AOI221_X1 U5519 ( .B1(D_REG_7__SCAN_IN), .B2(keyinput107), .C1(keyinput87), 
        .C2(D_REG_2__SCAN_IN), .A(n5013), .ZN(n5014) );
  NAND4_X1 U5520 ( .A1(n5017), .A2(n5016), .A3(n5015), .A4(n5014), .ZN(n5068)
         );
  OAI22_X1 U5521 ( .A1(REG3_REG_3__SCAN_IN), .A2(keyinput78), .B1(keyinput62), 
        .B2(REG0_REG_17__SCAN_IN), .ZN(n5018) );
  AOI221_X1 U5522 ( .B1(REG3_REG_3__SCAN_IN), .B2(keyinput78), .C1(
        REG0_REG_17__SCAN_IN), .C2(keyinput62), .A(n5018), .ZN(n5025) );
  OAI22_X1 U5523 ( .A1(DATAI_27_), .A2(keyinput71), .B1(REG0_REG_21__SCAN_IN), 
        .B2(keyinput108), .ZN(n5019) );
  AOI221_X1 U5524 ( .B1(DATAI_27_), .B2(keyinput71), .C1(keyinput108), .C2(
        REG0_REG_21__SCAN_IN), .A(n5019), .ZN(n5024) );
  OAI22_X1 U5525 ( .A1(ADDR_REG_15__SCAN_IN), .A2(keyinput92), .B1(keyinput35), 
        .B2(ADDR_REG_10__SCAN_IN), .ZN(n5020) );
  AOI221_X1 U5526 ( .B1(ADDR_REG_15__SCAN_IN), .B2(keyinput92), .C1(
        ADDR_REG_10__SCAN_IN), .C2(keyinput35), .A(n5020), .ZN(n5023) );
  OAI22_X1 U5527 ( .A1(REG3_REG_12__SCAN_IN), .A2(keyinput36), .B1(
        REG2_REG_10__SCAN_IN), .B2(keyinput82), .ZN(n5021) );
  AOI221_X1 U5528 ( .B1(REG3_REG_12__SCAN_IN), .B2(keyinput36), .C1(keyinput82), .C2(REG2_REG_10__SCAN_IN), .A(n5021), .ZN(n5022) );
  NAND4_X1 U5529 ( .A1(n5025), .A2(n5024), .A3(n5023), .A4(n5022), .ZN(n5067)
         );
  AOI22_X1 U5530 ( .A1(ADDR_REG_3__SCAN_IN), .A2(keyinput65), .B1(
        IR_REG_30__SCAN_IN), .B2(keyinput17), .ZN(n5026) );
  OAI221_X1 U5531 ( .B1(ADDR_REG_3__SCAN_IN), .B2(keyinput65), .C1(
        IR_REG_30__SCAN_IN), .C2(keyinput17), .A(n5026), .ZN(n5033) );
  AOI22_X1 U5532 ( .A1(DATAI_7_), .A2(keyinput57), .B1(REG0_REG_10__SCAN_IN), 
        .B2(keyinput85), .ZN(n5027) );
  OAI221_X1 U5533 ( .B1(DATAI_7_), .B2(keyinput57), .C1(REG0_REG_10__SCAN_IN), 
        .C2(keyinput85), .A(n5027), .ZN(n5032) );
  AOI22_X1 U5534 ( .A1(DATAO_REG_17__SCAN_IN), .A2(keyinput115), .B1(
        REG0_REG_2__SCAN_IN), .B2(keyinput95), .ZN(n5028) );
  OAI221_X1 U5535 ( .B1(DATAO_REG_17__SCAN_IN), .B2(keyinput115), .C1(
        REG0_REG_2__SCAN_IN), .C2(keyinput95), .A(n5028), .ZN(n5031) );
  AOI22_X1 U5536 ( .A1(D_REG_12__SCAN_IN), .A2(keyinput1), .B1(
        IR_REG_2__SCAN_IN), .B2(keyinput9), .ZN(n5029) );
  OAI221_X1 U5537 ( .B1(D_REG_12__SCAN_IN), .B2(keyinput1), .C1(
        IR_REG_2__SCAN_IN), .C2(keyinput9), .A(n5029), .ZN(n5030) );
  NOR4_X1 U5538 ( .A1(n5033), .A2(n5032), .A3(n5031), .A4(n5030), .ZN(n5065)
         );
  AOI22_X1 U5539 ( .A1(REG0_REG_14__SCAN_IN), .A2(keyinput16), .B1(
        REG1_REG_16__SCAN_IN), .B2(keyinput111), .ZN(n5034) );
  OAI221_X1 U5540 ( .B1(REG0_REG_14__SCAN_IN), .B2(keyinput16), .C1(
        REG1_REG_16__SCAN_IN), .C2(keyinput111), .A(n5034), .ZN(n5041) );
  AOI22_X1 U5541 ( .A1(REG0_REG_3__SCAN_IN), .A2(keyinput5), .B1(
        REG1_REG_10__SCAN_IN), .B2(keyinput93), .ZN(n5035) );
  OAI221_X1 U5542 ( .B1(REG0_REG_3__SCAN_IN), .B2(keyinput5), .C1(
        REG1_REG_10__SCAN_IN), .C2(keyinput93), .A(n5035), .ZN(n5040) );
  AOI22_X1 U5543 ( .A1(DATAI_8_), .A2(keyinput125), .B1(REG0_REG_27__SCAN_IN), 
        .B2(keyinput10), .ZN(n5036) );
  OAI221_X1 U5544 ( .B1(DATAI_8_), .B2(keyinput125), .C1(REG0_REG_27__SCAN_IN), 
        .C2(keyinput10), .A(n5036), .ZN(n5039) );
  AOI22_X1 U5545 ( .A1(DATAO_REG_27__SCAN_IN), .A2(keyinput19), .B1(
        DATAO_REG_18__SCAN_IN), .B2(keyinput15), .ZN(n5037) );
  OAI221_X1 U5546 ( .B1(DATAO_REG_27__SCAN_IN), .B2(keyinput19), .C1(
        DATAO_REG_18__SCAN_IN), .C2(keyinput15), .A(n5037), .ZN(n5038) );
  NOR4_X1 U5547 ( .A1(n5041), .A2(n5040), .A3(n5039), .A4(n5038), .ZN(n5064)
         );
  AOI22_X1 U5548 ( .A1(n2579), .A2(keyinput69), .B1(n5043), .B2(keyinput105), 
        .ZN(n5042) );
  OAI221_X1 U5549 ( .B1(n2579), .B2(keyinput69), .C1(n5043), .C2(keyinput105), 
        .A(n5042), .ZN(n5053) );
  AOI22_X1 U5550 ( .A1(n5045), .A2(keyinput103), .B1(keyinput18), .B2(n2622), 
        .ZN(n5044) );
  OAI221_X1 U5551 ( .B1(n5045), .B2(keyinput103), .C1(n2622), .C2(keyinput18), 
        .A(n5044), .ZN(n5052) );
  AOI22_X1 U5552 ( .A1(n3993), .A2(keyinput52), .B1(keyinput110), .B2(n5047), 
        .ZN(n5046) );
  OAI221_X1 U5553 ( .B1(n3993), .B2(keyinput52), .C1(n5047), .C2(keyinput110), 
        .A(n5046), .ZN(n5051) );
  XNOR2_X1 U5554 ( .A(n2244), .B(keyinput20), .ZN(n5049) );
  XNOR2_X1 U5555 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput119), .ZN(n5048) );
  NAND2_X1 U5556 ( .A1(n5049), .A2(n5048), .ZN(n5050) );
  NOR4_X1 U5557 ( .A1(n5053), .A2(n5052), .A3(n5051), .A4(n5050), .ZN(n5063)
         );
  AOI22_X1 U5558 ( .A1(DATAO_REG_1__SCAN_IN), .A2(keyinput60), .B1(
        REG1_REG_8__SCAN_IN), .B2(keyinput42), .ZN(n5054) );
  OAI221_X1 U5559 ( .B1(DATAO_REG_1__SCAN_IN), .B2(keyinput60), .C1(
        REG1_REG_8__SCAN_IN), .C2(keyinput42), .A(n5054), .ZN(n5061) );
  AOI22_X1 U5560 ( .A1(IR_REG_9__SCAN_IN), .A2(keyinput76), .B1(
        IR_REG_10__SCAN_IN), .B2(keyinput68), .ZN(n5055) );
  OAI221_X1 U5561 ( .B1(IR_REG_9__SCAN_IN), .B2(keyinput76), .C1(
        IR_REG_10__SCAN_IN), .C2(keyinput68), .A(n5055), .ZN(n5060) );
  AOI22_X1 U5562 ( .A1(D_REG_27__SCAN_IN), .A2(keyinput43), .B1(
        IR_REG_23__SCAN_IN), .B2(keyinput83), .ZN(n5056) );
  OAI221_X1 U5563 ( .B1(D_REG_27__SCAN_IN), .B2(keyinput43), .C1(
        IR_REG_23__SCAN_IN), .C2(keyinput83), .A(n5056), .ZN(n5059) );
  AOI22_X1 U5564 ( .A1(IR_REG_12__SCAN_IN), .A2(keyinput50), .B1(
        IR_REG_19__SCAN_IN), .B2(keyinput27), .ZN(n5057) );
  OAI221_X1 U5565 ( .B1(IR_REG_12__SCAN_IN), .B2(keyinput50), .C1(
        IR_REG_19__SCAN_IN), .C2(keyinput27), .A(n5057), .ZN(n5058) );
  NOR4_X1 U5566 ( .A1(n5061), .A2(n5060), .A3(n5059), .A4(n5058), .ZN(n5062)
         );
  NAND4_X1 U5567 ( .A1(n5065), .A2(n5064), .A3(n5063), .A4(n5062), .ZN(n5066)
         );
  NOR3_X1 U5568 ( .A1(n5068), .A2(n5067), .A3(n5066), .ZN(n5069) );
  NAND3_X1 U5569 ( .A1(n5071), .A2(n5070), .A3(n5069), .ZN(n5072) );
  NOR4_X1 U5570 ( .A1(n5075), .A2(n5074), .A3(n5073), .A4(n5072), .ZN(n5092)
         );
  AOI21_X1 U5571 ( .B1(n5076), .B2(n5078), .A(n5077), .ZN(n5090) );
  OAI22_X1 U5572 ( .A1(n5082), .A2(n5081), .B1(n5080), .B2(n5079), .ZN(n5088)
         );
  NAND2_X1 U5573 ( .A1(n3736), .A2(n5083), .ZN(n5085) );
  OAI211_X1 U5574 ( .C1(n3733), .C2(n5086), .A(n5085), .B(n5084), .ZN(n5087)
         );
  AOI211_X1 U5575 ( .C1(n5090), .C2(n5089), .A(n5088), .B(n5087), .ZN(n5091)
         );
  XNOR2_X1 U5576 ( .A(n5092), .B(n5091), .ZN(U3214) );
  CLKBUF_X2 U2501 ( .A(n2248), .Z(n3740) );
  CLKBUF_X1 U2925 ( .A(n2417), .Z(n3742) );
  XNOR2_X1 U3022 ( .A(n2403), .B(IR_REG_2__SCAN_IN), .ZN(n4495) );
endmodule

