

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD, 
        READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN, 
        M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN, 
        STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN, 
        W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N,
         BS16_N, READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN,
         CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN,
         REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN,
         FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191;

  AND2_X1 U34550 ( .A1(n5857), .A2(n4291), .ZN(n3504) );
  NAND2_X1 U34560 ( .A1(n3483), .A2(n3481), .ZN(n5854) );
  NAND2_X2 U3457 ( .A1(n4500), .A2(n4521), .ZN(n4540) );
  OR2_X1 U3458 ( .A1(n6493), .A2(n6492), .ZN(n6495) );
  CLKBUF_X1 U34590 ( .A(n4366), .Z(n4444) );
  CLKBUF_X2 U34600 ( .A(n4459), .Z(n4890) );
  INV_X1 U34610 ( .A(n4359), .ZN(n4850) );
  CLKBUF_X2 U34620 ( .A(n3582), .Z(n4666) );
  CLKBUF_X1 U34630 ( .A(n3577), .Z(n3773) );
  CLKBUF_X2 U34640 ( .A(n3617), .Z(n3448) );
  CLKBUF_X2 U34650 ( .A(n3778), .Z(n3425) );
  INV_X1 U3466 ( .A(n3676), .ZN(n4908) );
  AND2_X1 U3467 ( .A1(n4968), .A2(n3520), .ZN(n3778) );
  AND2_X1 U34680 ( .A1(n4968), .A2(n4964), .ZN(n3583) );
  AND2_X1 U34690 ( .A1(n6181), .A2(n4964), .ZN(n3699) );
  AND2_X2 U34700 ( .A1(n3519), .A2(n4968), .ZN(n3617) );
  AND2_X2 U34710 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4941) );
  CLKBUF_X1 U34720 ( .A(n5345), .Z(n3421) );
  NOR2_X1 U34730 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), 
        .ZN(n5345) );
  CLKBUF_X1 U34740 ( .A(n6960), .Z(n3422) );
  OAI211_X1 U3475 ( .C1(n4880), .C2(n4879), .A(n4878), .B(n4877), .ZN(n6960)
         );
  NOR2_X2 U3476 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3520) );
  AND2_X1 U3478 ( .A1(n4941), .A2(n4964), .ZN(n3714) );
  AND2_X1 U3479 ( .A1(n6181), .A2(n3520), .ZN(n3811) );
  NOR2_X1 U3480 ( .A1(n3698), .A2(n6923), .ZN(n4329) );
  NAND4_X1 U3481 ( .A1(n3611), .A2(n3610), .A3(n3609), .A4(n3608), .ZN(n3658)
         );
  BUF_X1 U3482 ( .A(n3681), .Z(n3446) );
  INV_X1 U3483 ( .A(n3757), .ZN(n4691) );
  INV_X2 U3484 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4950) );
  INV_X1 U3485 ( .A(n3658), .ZN(n3480) );
  INV_X1 U3486 ( .A(n4540), .ZN(n6019) );
  AND2_X1 U3487 ( .A1(n5445), .A2(n5444), .ZN(n5497) );
  NOR2_X2 U3488 ( .A1(n5674), .A2(n5708), .ZN(n5686) );
  INV_X1 U3489 ( .A(n6865), .ZN(n6827) );
  INV_X1 U3490 ( .A(n6861), .ZN(n6833) );
  OR2_X2 U3491 ( .A1(n3732), .A2(n3731), .ZN(n3733) );
  NAND2_X2 U3492 ( .A1(n3671), .A2(n3670), .ZN(n3732) );
  AND4_X2 U3493 ( .A1(n3534), .A2(n3533), .A3(n3532), .A4(n3531), .ZN(n3545)
         );
  AOI21_X2 U3494 ( .B1(n3691), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3665), 
        .ZN(n3667) );
  XNOR2_X2 U3495 ( .A(n4627), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5988)
         );
  CLKBUF_X1 U3496 ( .A(n3811), .Z(n3423) );
  CLKBUF_X1 U3497 ( .A(n3811), .Z(n3424) );
  BUF_X2 U3498 ( .A(n4540), .Z(n3449) );
  NAND2_X1 U3499 ( .A1(n3820), .A2(n3821), .ZN(n3854) );
  OR2_X1 U3500 ( .A1(n5532), .A2(n5533), .ZN(n5645) );
  NAND2_X2 U3501 ( .A1(n3436), .A2(n3733), .ZN(n3792) );
  NAND2_X1 U3502 ( .A1(n4345), .A2(n4344), .ZN(n5817) );
  NOR2_X2 U3503 ( .A1(n4845), .A2(n4844), .ZN(n6504) );
  OR2_X1 U3504 ( .A1(n4834), .A2(n4827), .ZN(n4845) );
  CLKBUF_X2 U3505 ( .A(n3679), .Z(n6581) );
  CLKBUF_X2 U3506 ( .A(n3480), .Z(n4886) );
  INV_X1 U3507 ( .A(n3659), .ZN(n4913) );
  NAND2_X4 U3508 ( .A1(n3447), .A2(n3659), .ZN(n4359) );
  BUF_X2 U3509 ( .A(n3712), .Z(n4231) );
  BUF_X2 U3510 ( .A(n3612), .Z(n4267) );
  CLKBUF_X2 U3511 ( .A(n3576), .Z(n4650) );
  AND2_X2 U3512 ( .A1(n6180), .A2(n3520), .ZN(n3762) );
  NAND2_X1 U3514 ( .A1(n6009), .A2(n4543), .ZN(n5996) );
  NAND2_X1 U3515 ( .A1(n3438), .A2(n6010), .ZN(n6009) );
  INV_X1 U3516 ( .A(n5929), .ZN(n3483) );
  AOI21_X1 U3517 ( .B1(n5940), .B2(n3498), .A(n3453), .ZN(n6973) );
  AND2_X1 U3518 ( .A1(n5946), .A2(n5947), .ZN(n5938) );
  NAND2_X1 U3519 ( .A1(n5632), .A2(n4004), .ZN(n5652) );
  AND2_X1 U3520 ( .A1(n3427), .A2(n3428), .ZN(n5674) );
  OR2_X1 U3521 ( .A1(n3429), .A2(n4004), .ZN(n3428) );
  NAND2_X1 U3522 ( .A1(n3909), .A2(n3908), .ZN(n5084) );
  NAND2_X1 U3523 ( .A1(n5869), .A2(n3464), .ZN(n5793) );
  NOR2_X2 U3524 ( .A1(n5883), .A2(n4439), .ZN(n5869) );
  NOR2_X1 U3525 ( .A1(n4529), .A2(n3458), .ZN(n3470) );
  OAI21_X1 U3526 ( .B1(n4516), .B2(n4519), .A(n4515), .ZN(n4517) );
  AOI21_X1 U3527 ( .B1(n4492), .B2(n4028), .A(n3876), .ZN(n5043) );
  NAND2_X1 U3528 ( .A1(n3907), .A2(n3906), .ZN(n5085) );
  NAND2_X1 U3529 ( .A1(n4540), .A2(n6096), .ZN(n4544) );
  NOR2_X1 U3530 ( .A1(n3867), .A2(n3479), .ZN(n4492) );
  XNOR2_X1 U3531 ( .A(n4500), .B(n3892), .ZN(n4510) );
  XNOR2_X1 U3532 ( .A(n3854), .B(n3843), .ZN(n4486) );
  NAND2_X1 U3533 ( .A1(n3741), .A2(n3740), .ZN(n4988) );
  NAND2_X1 U3534 ( .A1(n3819), .A2(n3818), .ZN(n3821) );
  CLKBUF_X1 U3535 ( .A(n4891), .Z(n5548) );
  AND2_X1 U3536 ( .A1(n4811), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4810)
         );
  NAND2_X1 U3537 ( .A1(n3729), .A2(n3728), .ZN(n3754) );
  OAI21_X2 U3538 ( .B1(n3792), .B2(STATE2_REG_0__SCAN_IN), .A(n3791), .ZN(
        n5746) );
  NAND2_X1 U3539 ( .A1(n5817), .A2(n5829), .ZN(n4880) );
  AOI21_X1 U3540 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6923), .A(n4333), 
        .ZN(n4342) );
  CLKBUF_X1 U3541 ( .A(n4746), .Z(n3432) );
  NOR2_X1 U3542 ( .A1(n4346), .A2(n3657), .ZN(n3663) );
  NAND2_X1 U3543 ( .A1(n4561), .A2(n3641), .ZN(n3672) );
  AND2_X1 U3544 ( .A1(n3661), .A2(n4355), .ZN(n3688) );
  NAND2_X1 U3545 ( .A1(n3640), .A2(n6183), .ZN(n4561) );
  INV_X1 U3546 ( .A(n3653), .ZN(n4351) );
  NAND2_X2 U3547 ( .A1(n3480), .A2(n4913), .ZN(n3673) );
  NAND2_X1 U3548 ( .A1(n3635), .A2(n3636), .ZN(n3660) );
  AND2_X1 U3549 ( .A1(n3698), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4340) );
  CLKBUF_X1 U3550 ( .A(n3636), .Z(n4455) );
  OR2_X1 U3551 ( .A1(n3725), .A2(n3724), .ZN(n4454) );
  NAND2_X2 U3552 ( .A1(n3506), .A2(n3507), .ZN(n3746) );
  OR2_X1 U3553 ( .A1(n3785), .A2(n3784), .ZN(n4523) );
  AND4_X1 U3554 ( .A1(n3629), .A2(n3628), .A3(n3627), .A4(n3626), .ZN(n3630)
         );
  AND4_X1 U3555 ( .A1(n3625), .A2(n3624), .A3(n3623), .A4(n3622), .ZN(n3631)
         );
  AND4_X1 U3556 ( .A1(n3607), .A2(n3606), .A3(n3605), .A4(n3604), .ZN(n3608)
         );
  AND4_X1 U3557 ( .A1(n3602), .A2(n3601), .A3(n3600), .A4(n3599), .ZN(n3609)
         );
  AND4_X1 U3558 ( .A1(n3598), .A2(n3597), .A3(n3596), .A4(n3595), .ZN(n3610)
         );
  AND4_X1 U3559 ( .A1(n3594), .A2(n3593), .A3(n3592), .A4(n3591), .ZN(n3611)
         );
  AND4_X1 U3560 ( .A1(n3587), .A2(n3586), .A3(n3585), .A4(n3584), .ZN(n3455)
         );
  AND4_X1 U3561 ( .A1(n3570), .A2(n3569), .A3(n3568), .A4(n3567), .ZN(n3506)
         );
  AND4_X1 U3562 ( .A1(n3524), .A2(n3523), .A3(n3522), .A4(n3521), .ZN(n3525)
         );
  AND4_X1 U3563 ( .A1(n3517), .A2(n3516), .A3(n3515), .A4(n3514), .ZN(n3526)
         );
  AND4_X1 U3564 ( .A1(n3542), .A2(n3541), .A3(n3540), .A4(n3539), .ZN(n3543)
         );
  AND4_X1 U3565 ( .A1(n3530), .A2(n3529), .A3(n3528), .A4(n3527), .ZN(n3546)
         );
  AND4_X1 U3566 ( .A1(n3555), .A2(n3554), .A3(n3553), .A4(n3552), .ZN(n3556)
         );
  AND4_X1 U3567 ( .A1(n3550), .A2(n3549), .A3(n3548), .A4(n3547), .ZN(n3557)
         );
  AND4_X1 U3568 ( .A1(n3616), .A2(n3615), .A3(n3614), .A4(n3613), .ZN(n3633)
         );
  AND4_X1 U3569 ( .A1(n3538), .A2(n3537), .A3(n3536), .A4(n3535), .ZN(n3544)
         );
  AND4_X1 U3570 ( .A1(n3621), .A2(n3620), .A3(n3619), .A4(n3618), .ZN(n3632)
         );
  BUF_X2 U3571 ( .A(n3762), .Z(n3441) );
  BUF_X2 U3572 ( .A(n3699), .Z(n4673) );
  CLKBUF_X2 U3573 ( .A(n3762), .Z(n3440) );
  BUF_X2 U3574 ( .A(n3583), .Z(n4667) );
  BUF_X2 U3575 ( .A(n3714), .Z(n3779) );
  AND2_X2 U3576 ( .A1(n3518), .A2(n4941), .ZN(n3443) );
  AND2_X2 U3577 ( .A1(n3518), .A2(n4941), .ZN(n3719) );
  AND2_X2 U3578 ( .A1(n6181), .A2(n3518), .ZN(n3445) );
  AND2_X2 U3579 ( .A1(n3518), .A2(n4968), .ZN(n3713) );
  AND2_X2 U3580 ( .A1(n6181), .A2(n3519), .ZN(n3582) );
  AND2_X2 U3581 ( .A1(n6181), .A2(n3518), .ZN(n4072) );
  OR2_X2 U3582 ( .A1(n6571), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6821) );
  AND2_X2 U3583 ( .A1(n3512), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3518)
         );
  AND2_X2 U3584 ( .A1(n3511), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n6181)
         );
  AND2_X1 U3585 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4964) );
  CLKBUF_X1 U3586 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n5774) );
  AND2_X1 U3587 ( .A1(n3497), .A2(n5947), .ZN(n3426) );
  NAND2_X1 U3588 ( .A1(n5628), .A2(n3430), .ZN(n3427) );
  INV_X1 U3589 ( .A(n3499), .ZN(n3429) );
  AND2_X1 U3590 ( .A1(n5629), .A2(n3499), .ZN(n3430) );
  NAND2_X1 U3591 ( .A1(n3694), .A2(n3693), .ZN(n3431) );
  NAND2_X1 U3592 ( .A1(n3694), .A2(n3693), .ZN(n4970) );
  NAND2_X1 U3593 ( .A1(n3642), .A2(n4596), .ZN(n4746) );
  NAND2_X2 U3594 ( .A1(n3668), .A2(n3690), .ZN(n3711) );
  NAND2_X1 U3595 ( .A1(n6008), .A2(n6010), .ZN(n3433) );
  AND2_X2 U3596 ( .A1(n3433), .A2(n3434), .ZN(n4640) );
  AND2_X1 U3597 ( .A1(n4544), .A2(n4543), .ZN(n3434) );
  CLKBUF_X1 U3598 ( .A(n5333), .Z(n3435) );
  NAND2_X1 U3599 ( .A1(n3732), .A2(n3731), .ZN(n3436) );
  CLKBUF_X1 U3600 ( .A(n6538), .Z(n3437) );
  NOR2_X1 U3601 ( .A1(n4542), .A2(n3457), .ZN(n3438) );
  NOR2_X1 U3602 ( .A1(n4542), .A2(n3457), .ZN(n6008) );
  NAND2_X1 U3603 ( .A1(n3739), .A2(n3738), .ZN(n3755) );
  NAND2_X1 U3604 ( .A1(n4713), .A2(n4746), .ZN(n4584) );
  OAI21_X1 U3605 ( .B1(n4706), .B2(n6942), .A(n4583), .ZN(n3647) );
  AND2_X1 U3606 ( .A1(n3518), .A2(n6180), .ZN(n3439) );
  NAND2_X2 U3607 ( .A1(n3526), .A2(n3525), .ZN(n3634) );
  AND2_X1 U3608 ( .A1(n3518), .A2(n4941), .ZN(n3442) );
  AND2_X1 U3609 ( .A1(n6181), .A2(n3518), .ZN(n3444) );
  NAND2_X2 U3610 ( .A1(n6527), .A2(n6525), .ZN(n6526) );
  NAND2_X1 U3611 ( .A1(n6518), .A2(n4491), .ZN(n6527) );
  AND3_X2 U3612 ( .A1(n6029), .A2(n6155), .A3(n4620), .ZN(n3457) );
  NAND2_X1 U3613 ( .A1(n4468), .A2(n4467), .ZN(n6511) );
  NOR2_X2 U3614 ( .A1(n5723), .A2(n5724), .ZN(n5946) );
  INV_X2 U3615 ( .A(n3636), .ZN(n5155) );
  OAI222_X1 U3616 ( .A1(n5741), .A2(n4892), .B1(n5150), .B2(n6883), .C1(n5745), 
        .C2(n4983), .ZN(U3463) );
  AOI21_X1 U3617 ( .B1(n3691), .B2(n5774), .A(n3692), .ZN(n3695) );
  AND2_X2 U3618 ( .A1(n3664), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3691) );
  XNOR2_X1 U3619 ( .A(n4490), .B(n6627), .ZN(n6519) );
  NAND2_X1 U3620 ( .A1(n4489), .A2(n4488), .ZN(n4490) );
  AOI21_X2 U3621 ( .B1(n4459), .B2(n4574), .A(n4458), .ZN(n5523) );
  XNOR2_X2 U3622 ( .A(n3756), .B(n3755), .ZN(n4459) );
  AND2_X2 U3623 ( .A1(n4988), .A2(n3822), .ZN(n4888) );
  NAND4_X1 U3624 ( .A1(n3611), .A2(n3610), .A3(n3609), .A4(n3608), .ZN(n3447)
         );
  NAND2_X2 U3625 ( .A1(n3500), .A2(n3636), .ZN(n3653) );
  INV_X2 U3626 ( .A(n3634), .ZN(n3500) );
  NOR2_X4 U3627 ( .A1(n4292), .A2(n3504), .ZN(n5986) );
  NAND4_X4 U3628 ( .A1(n3546), .A2(n3545), .A3(n3544), .A4(n3543), .ZN(n3636)
         );
  OAI21_X2 U3629 ( .B1(n5538), .B2(n3469), .A(n3468), .ZN(n6552) );
  NAND2_X2 U3630 ( .A1(n5590), .A2(n4528), .ZN(n5538) );
  OAI21_X2 U3631 ( .B1(n5699), .B2(n5695), .A(n5696), .ZN(n6072) );
  OAI21_X2 U3632 ( .B1(n5637), .B2(n4535), .A(n4534), .ZN(n5699) );
  NOR2_X2 U3633 ( .A1(n5084), .A2(n3493), .ZN(n5459) );
  AND2_X2 U3634 ( .A1(n4289), .A2(n3490), .ZN(n3451) );
  NOR2_X4 U3635 ( .A1(n5854), .A2(n5855), .ZN(n4289) );
  INV_X2 U3636 ( .A(n3654), .ZN(n5160) );
  NAND2_X4 U3637 ( .A1(n3588), .A2(n3455), .ZN(n3654) );
  NAND2_X2 U3638 ( .A1(n4970), .A2(n3697), .ZN(n4892) );
  XNOR2_X2 U3639 ( .A(n3711), .B(n3730), .ZN(n4893) );
  AND2_X4 U3640 ( .A1(n6180), .A2(n4964), .ZN(n3577) );
  INV_X1 U3641 ( .A(n3421), .ZN(n4685) );
  AND2_X1 U3642 ( .A1(n3842), .A2(n3841), .ZN(n3853) );
  NAND2_X1 U3643 ( .A1(n6071), .A2(n3459), .ZN(n3476) );
  INV_X1 U3644 ( .A(n5930), .ZN(n4186) );
  NAND2_X1 U3645 ( .A1(n3995), .A2(n3502), .ZN(n4004) );
  NAND2_X1 U3646 ( .A1(n3496), .A2(n5443), .ZN(n3495) );
  INV_X1 U3647 ( .A(n5250), .ZN(n3496) );
  AND2_X1 U3648 ( .A1(n3659), .A2(n4455), .ZN(n4574) );
  NAND2_X1 U3649 ( .A1(n3634), .A2(n3746), .ZN(n4357) );
  AND2_X1 U3650 ( .A1(n3755), .A2(n3754), .ZN(n3743) );
  AND2_X1 U3651 ( .A1(n4329), .A2(n4574), .ZN(n4343) );
  OR2_X1 U3652 ( .A1(n5817), .A2(n5824), .ZN(n4757) );
  AND2_X1 U3653 ( .A1(n3421), .A2(n6007), .ZN(n4222) );
  AND2_X1 U3654 ( .A1(n5881), .A2(n3485), .ZN(n3484) );
  INV_X1 U3655 ( .A(n6026), .ZN(n3485) );
  NAND2_X1 U3656 ( .A1(n5459), .A2(n5494), .ZN(n3998) );
  OR2_X1 U3657 ( .A1(n3840), .A2(n3839), .ZN(n4493) );
  NAND2_X1 U3658 ( .A1(n4460), .A2(n3659), .ZN(n4383) );
  NAND2_X1 U3659 ( .A1(n3653), .A2(n3654), .ZN(n3683) );
  OR2_X1 U3660 ( .A1(n3660), .A2(n4383), .ZN(n4355) );
  INV_X1 U3661 ( .A(n5043), .ZN(n3877) );
  AND2_X1 U3662 ( .A1(n3745), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3793) );
  INV_X1 U3663 ( .A(n3475), .ZN(n3474) );
  OAI21_X1 U3664 ( .B1(n4536), .B2(n3476), .A(n4538), .ZN(n3475) );
  AND2_X1 U3665 ( .A1(n4557), .A2(n4913), .ZN(n3641) );
  OR2_X1 U3666 ( .A1(n3817), .A2(n3816), .ZN(n4480) );
  OAI22_X1 U3667 ( .A1(n4332), .A2(n4331), .B1(n4330), .B2(n4569), .ZN(n4333)
         );
  NOR2_X1 U3668 ( .A1(n3480), .A2(n3659), .ZN(n3679) );
  OR2_X1 U3669 ( .A1(n6910), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4694) );
  AND2_X1 U3670 ( .A1(n5869), .A2(n3463), .ZN(n4590) );
  AND2_X1 U3671 ( .A1(n4121), .A2(n4120), .ZN(n5947) );
  AND2_X1 U3672 ( .A1(n4381), .A2(n4380), .ZN(n6503) );
  OAI211_X1 U3673 ( .C1(n4359), .C2(EBX_REG_5__SCAN_IN), .A(n4444), .B(n4379), 
        .ZN(n4380) );
  NAND2_X1 U3674 ( .A1(n4444), .A2(n4374), .ZN(n5790) );
  NOR2_X1 U3675 ( .A1(n3489), .A2(n3492), .ZN(n3488) );
  INV_X1 U3676 ( .A(n3490), .ZN(n3489) );
  NOR2_X1 U3677 ( .A1(n3482), .A2(n5867), .ZN(n3481) );
  INV_X1 U3678 ( .A(n3484), .ZN(n3482) );
  NAND2_X1 U3679 ( .A1(n4188), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4221)
         );
  AND2_X1 U3680 ( .A1(n4083), .A2(n5687), .ZN(n4084) );
  NAND2_X1 U3681 ( .A1(n5460), .A2(n3494), .ZN(n3493) );
  INV_X1 U3682 ( .A(n3495), .ZN(n3494) );
  NAND2_X1 U3683 ( .A1(n5793), .A2(n4595), .ZN(n5791) );
  AND2_X1 U3684 ( .A1(n5978), .A2(n4547), .ZN(n5747) );
  AND2_X1 U3685 ( .A1(n5869), .A2(n4628), .ZN(n4630) );
  NAND2_X1 U3686 ( .A1(n6552), .A2(n6553), .ZN(n4533) );
  NAND2_X1 U3687 ( .A1(n6526), .A2(n4499), .ZN(n6533) );
  NAND2_X1 U3688 ( .A1(n6533), .A2(n6532), .ZN(n6531) );
  OR2_X1 U3689 ( .A1(n5152), .A2(n4889), .ZN(n4923) );
  INV_X1 U3690 ( .A(n6080), .ZN(n4451) );
  OR2_X1 U3691 ( .A1(n4362), .A2(n4361), .ZN(n6510) );
  AND2_X1 U3692 ( .A1(n4606), .A2(n4594), .ZN(n6721) );
  INV_X1 U3693 ( .A(n4890), .ZN(n5152) );
  AOI21_X1 U3694 ( .B1(n4328), .B2(n4327), .A(n4326), .ZN(n4335) );
  AND2_X1 U3695 ( .A1(n3673), .A2(n4307), .ZN(n4321) );
  NOR2_X1 U3696 ( .A1(n4317), .A2(n4564), .ZN(n4319) );
  AND2_X1 U3697 ( .A1(n3575), .A2(n3746), .ZN(n3650) );
  INV_X1 U3698 ( .A(n4346), .ZN(n4556) );
  OAI21_X1 U3699 ( .B1(n3659), .B2(n3655), .A(n5155), .ZN(n3656) );
  NAND2_X1 U3700 ( .A1(n3441), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U3701 ( .A1(n3445), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3762), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3564) );
  AND2_X1 U3702 ( .A1(n3713), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3551) );
  NAND2_X1 U3703 ( .A1(n3441), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3529) );
  AOI22_X1 U3704 ( .A1(n3444), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3762), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3517) );
  NAND2_X1 U3705 ( .A1(n3650), .A2(n5160), .ZN(n4350) );
  AOI22_X1 U3706 ( .A1(n3576), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3568) );
  NAND2_X1 U3707 ( .A1(n3778), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3605) );
  NAND2_X1 U3708 ( .A1(n3583), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3604)
         );
  AND2_X1 U3709 ( .A1(n3491), .A2(n4290), .ZN(n3490) );
  INV_X1 U3710 ( .A(n5760), .ZN(n3491) );
  NOR2_X1 U3711 ( .A1(n4283), .A2(n5989), .ZN(n4284) );
  NAND2_X1 U3712 ( .A1(n3898), .A2(n3900), .ZN(n4501) );
  INV_X1 U3713 ( .A(n6073), .ZN(n4536) );
  AND2_X1 U3714 ( .A1(n3868), .A2(n3899), .ZN(n3501) );
  OR2_X1 U3715 ( .A1(n3709), .A2(n3708), .ZN(n4476) );
  AOI22_X1 U3716 ( .A1(n4072), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3441), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U3717 ( .A1(n3617), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3585) );
  AND2_X1 U3718 ( .A1(n4603), .A2(n4356), .ZN(n4749) );
  AND2_X2 U3719 ( .A1(n4950), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3519)
         );
  NAND2_X1 U3720 ( .A1(n3727), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3728) );
  NAND2_X1 U3721 ( .A1(n3737), .A2(n3736), .ZN(n3739) );
  AOI21_X1 U3722 ( .B1(n6925), .B2(n6914), .A(n5778), .ZN(n4887) );
  INV_X1 U3723 ( .A(n4946), .ZN(n5824) );
  CLKBUF_X1 U3724 ( .A(n4706), .Z(n5818) );
  OR2_X1 U3725 ( .A1(n4850), .A2(n4363), .ZN(n4364) );
  NAND2_X1 U3726 ( .A1(n4366), .A2(EBX_REG_0__SCAN_IN), .ZN(n4368) );
  AND2_X1 U3727 ( .A1(n4857), .A2(n5827), .ZN(n6406) );
  INV_X1 U3728 ( .A(n4877), .ZN(n4795) );
  OR2_X1 U3729 ( .A1(n4354), .A2(n4359), .ZN(n4713) );
  OR2_X1 U3730 ( .A1(n4687), .A2(n5839), .ZN(n4698) );
  AND2_X1 U3731 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n4243), .ZN(n4244)
         );
  INV_X1 U3732 ( .A(n4242), .ZN(n4243) );
  NAND2_X1 U3733 ( .A1(n4244), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4283)
         );
  OR2_X1 U3734 ( .A1(n4221), .A2(n6024), .ZN(n4242) );
  AND2_X1 U3735 ( .A1(n4205), .A2(n4204), .ZN(n6026) );
  OR2_X1 U3736 ( .A1(n6862), .A2(n4685), .ZN(n4205) );
  NOR2_X1 U3737 ( .A1(n5894), .A2(n3498), .ZN(n3497) );
  NOR2_X1 U3738 ( .A1(n4102), .A2(n4101), .ZN(n4103) );
  AND2_X1 U3739 ( .A1(n4103), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4138)
         );
  NAND2_X1 U3740 ( .A1(n4051), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4102)
         );
  NAND2_X1 U3741 ( .A1(n4050), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4067)
         );
  AND2_X1 U3742 ( .A1(n4036), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4050)
         );
  NOR2_X1 U3743 ( .A1(n4019), .A2(n5660), .ZN(n4036) );
  AND2_X1 U3744 ( .A1(n4035), .A2(n5651), .ZN(n3499) );
  INV_X1 U3745 ( .A(n5676), .ZN(n4035) );
  NOR2_X1 U3746 ( .A1(n4000), .A2(n3968), .ZN(n4001) );
  NAND2_X1 U3747 ( .A1(n4001), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4019)
         );
  AND2_X1 U3748 ( .A1(n4004), .A2(n3999), .ZN(n5628) );
  NAND2_X1 U3749 ( .A1(n3967), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4000)
         );
  NAND2_X1 U3750 ( .A1(n3949), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3953)
         );
  NOR2_X1 U3751 ( .A1(n3925), .A2(n3920), .ZN(n3949) );
  AND4_X1 U3752 ( .A1(n3924), .A2(n3923), .A3(n3922), .A4(n3921), .ZN(n5250)
         );
  OR2_X1 U3753 ( .A1(n3903), .A2(n6771), .ZN(n3925) );
  AND2_X1 U3754 ( .A1(n5086), .A2(n5085), .ZN(n3908) );
  NAND2_X1 U3755 ( .A1(n3901), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3903)
         );
  INV_X1 U3756 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3871) );
  NOR2_X1 U3757 ( .A1(n3872), .A2(n3871), .ZN(n3901) );
  CLKBUF_X1 U3758 ( .A(n5041), .Z(n5042) );
  AND3_X1 U3759 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A3(PHYADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n3848) );
  AOI21_X1 U3760 ( .B1(n4978), .B2(n4028), .A(n3830), .ZN(n4832) );
  NOR2_X2 U3761 ( .A1(n4831), .A2(n4832), .ZN(n4843) );
  OAI211_X1 U3762 ( .C1(n4359), .C2(EBX_REG_27__SCAN_IN), .A(n4441), .B(n4444), 
        .ZN(n4442) );
  NAND2_X1 U3763 ( .A1(n3467), .A2(n3465), .ZN(n5883) );
  NOR2_X1 U3764 ( .A1(n4541), .A2(n3449), .ZN(n4542) );
  INV_X1 U3765 ( .A(n3467), .ZN(n6112) );
  NAND2_X1 U3766 ( .A1(n5943), .A2(n5896), .ZN(n5933) );
  OR2_X1 U3767 ( .A1(n5950), .A2(n5949), .ZN(n5952) );
  OAI211_X1 U3768 ( .C1(n4359), .C2(EBX_REG_19__SCAN_IN), .A(n4418), .B(n4444), 
        .ZN(n4419) );
  NAND2_X1 U3769 ( .A1(n5725), .A2(n5726), .ZN(n5950) );
  OR2_X1 U3770 ( .A1(n3449), .A2(n6707), .ZN(n6071) );
  OR2_X1 U3771 ( .A1(n4540), .A2(n5635), .ZN(n4534) );
  NOR2_X1 U3772 ( .A1(n3449), .A2(n6700), .ZN(n5695) );
  OAI211_X1 U3773 ( .C1(n4359), .C2(EBX_REG_15__SCAN_IN), .A(n4408), .B(n4444), 
        .ZN(n4409) );
  AOI21_X1 U3774 ( .B1(n3470), .B2(n3452), .A(n3461), .ZN(n3468) );
  INV_X1 U3775 ( .A(n3470), .ZN(n3469) );
  XNOR2_X1 U3776 ( .A(n3449), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6553)
         );
  AND2_X1 U3777 ( .A1(n4402), .A2(n4401), .ZN(n5533) );
  NAND2_X1 U3778 ( .A1(n5497), .A2(n4399), .ZN(n5532) );
  AND2_X1 U3779 ( .A1(n4390), .A2(n4389), .ZN(n5264) );
  NOR2_X2 U3780 ( .A1(n6495), .A2(n5264), .ZN(n5445) );
  NAND2_X1 U3781 ( .A1(n6504), .A2(n3460), .ZN(n6493) );
  AND2_X1 U3782 ( .A1(n6504), .A2(n6503), .ZN(n6506) );
  OR2_X1 U3783 ( .A1(n5790), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4375)
         );
  OAI21_X1 U3784 ( .B1(n4482), .B2(n4519), .A(n4481), .ZN(n4823) );
  OR3_X1 U3785 ( .A1(n4880), .A2(n4580), .A3(n3676), .ZN(n4581) );
  INV_X1 U3786 ( .A(n4329), .ZN(n4297) );
  INV_X1 U3787 ( .A(n3669), .ZN(n3670) );
  AND4_X1 U3788 ( .A1(n3688), .A2(n3687), .A3(n3686), .A4(n3685), .ZN(n3689)
         );
  INV_X1 U3789 ( .A(n3695), .ZN(n3693) );
  AND2_X2 U3790 ( .A1(n3513), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6180)
         );
  INV_X1 U3791 ( .A(n5256), .ZN(n5212) );
  NOR2_X1 U3792 ( .A1(n4989), .A2(n4978), .ZN(n7040) );
  NOR2_X1 U3793 ( .A1(n5451), .A2(n7052), .ZN(n5127) );
  OR2_X1 U3794 ( .A1(n5548), .A2(n7052), .ZN(n5553) );
  AND2_X1 U3795 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7041) );
  INV_X1 U3796 ( .A(n7162), .ZN(n5162) );
  AND2_X1 U3797 ( .A1(n4977), .A2(n5152), .ZN(n5221) );
  INV_X1 U3798 ( .A(n5746), .ZN(n6990) );
  OR3_X1 U3799 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4887), .A3(n6916), .ZN(n5161) );
  NAND2_X1 U3800 ( .A1(n4342), .A2(n4341), .ZN(n4345) );
  AND2_X1 U3801 ( .A1(n5348), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4358) );
  AND2_X1 U3802 ( .A1(n6756), .A2(n5354), .ZN(n6861) );
  NAND2_X1 U3803 ( .A1(n5352), .A2(n5351), .ZN(n6847) );
  AND2_X1 U3804 ( .A1(n6583), .A2(n5360), .ZN(n6855) );
  NAND2_X1 U3805 ( .A1(n5791), .A2(n3466), .ZN(n5794) );
  OR2_X1 U3806 ( .A1(n5793), .A2(n5792), .ZN(n3466) );
  INV_X1 U3807 ( .A(n6510), .ZN(n6200) );
  INV_X1 U3808 ( .A(n3746), .ZN(n5812) );
  AND2_X1 U3809 ( .A1(n3422), .A2(n3745), .ZN(n7077) );
  INV_X1 U3810 ( .A(n7078), .ZN(n5976) );
  CLKBUF_X1 U3811 ( .A(n4764), .Z(n4806) );
  OR2_X1 U3812 ( .A1(n4880), .A2(n6904), .ZN(n4856) );
  INV_X1 U3813 ( .A(n4764), .ZN(n4743) );
  OR2_X1 U3814 ( .A1(n3488), .A2(n4692), .ZN(n3487) );
  NAND2_X1 U3815 ( .A1(n3483), .A2(n3484), .ZN(n5866) );
  INV_X1 U3816 ( .A(n6828), .ZN(n6970) );
  INV_X1 U3817 ( .A(n6869), .ZN(n6562) );
  OR2_X1 U3818 ( .A1(n4880), .A2(n6891), .ZN(n6869) );
  INV_X2 U3819 ( .A(n6069), .ZN(n6561) );
  XNOR2_X1 U3820 ( .A(n4592), .B(n5792), .ZN(n5920) );
  XNOR2_X1 U3821 ( .A(n5750), .B(n5749), .ZN(n5765) );
  AOI22_X1 U3822 ( .A1(n5979), .A2(n5747), .B1(n6082), .B2(n3449), .ZN(n5750)
         );
  NAND2_X1 U3823 ( .A1(n6531), .A2(n4509), .ZN(n6540) );
  NAND2_X1 U3824 ( .A1(n4606), .A2(n4946), .ZN(n6651) );
  OR2_X1 U3825 ( .A1(n6725), .A2(n6727), .ZN(n6694) );
  INV_X1 U3826 ( .A(n4893), .ZN(n5357) );
  INV_X1 U3827 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5348) );
  INV_X1 U3828 ( .A(n6924), .ZN(n5778) );
  INV_X1 U3829 ( .A(n7035), .ZN(n7177) );
  INV_X1 U3830 ( .A(n7036), .ZN(n7175) );
  NOR2_X1 U3831 ( .A1(n4923), .A2(n4899), .ZN(n5312) );
  INV_X1 U3832 ( .A(n6997), .ZN(n7168) );
  AND2_X1 U3833 ( .A1(n5221), .A2(n6990), .ZN(n7154) );
  INV_X1 U3834 ( .A(n7059), .ZN(n5578) );
  INV_X1 U3835 ( .A(n7076), .ZN(n5570) );
  INV_X1 U3836 ( .A(n7111), .ZN(n5574) );
  INV_X1 U3837 ( .A(n7125), .ZN(n5558) );
  INV_X1 U3838 ( .A(n7153), .ZN(n5566) );
  INV_X1 U3839 ( .A(n5255), .ZN(n5274) );
  INV_X1 U3840 ( .A(n5005), .ZN(n5283) );
  NAND2_X1 U3841 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5817), .ZN(n6924) );
  INV_X1 U3842 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6916) );
  XNOR2_X1 U3843 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n6942) );
  NAND2_X1 U3844 ( .A1(n5986), .A2(n6508), .ZN(n4453) );
  INV_X1 U3845 ( .A(n4633), .ZN(n4634) );
  OAI21_X1 U3846 ( .B1(n5926), .B2(n6709), .A(n4632), .ZN(n4633) );
  AND2_X2 U3847 ( .A1(n4941), .A2(n3520), .ZN(n3603) );
  NOR2_X1 U3848 ( .A1(n4460), .A2(n3676), .ZN(n3681) );
  NAND2_X1 U3849 ( .A1(n3477), .A2(n4536), .ZN(n6070) );
  NOR2_X1 U3850 ( .A1(n6019), .A2(n4530), .ZN(n3452) );
  NOR2_X1 U3851 ( .A1(n5084), .A2(n5250), .ZN(n5249) );
  AND2_X1 U3852 ( .A1(n5938), .A2(n5939), .ZN(n3453) );
  NOR2_X1 U3853 ( .A1(n5929), .A2(n6026), .ZN(n5880) );
  NAND2_X1 U3854 ( .A1(n6070), .A2(n6071), .ZN(n6058) );
  AND2_X2 U3855 ( .A1(n3519), .A2(n6180), .ZN(n3576) );
  AND4_X1 U3856 ( .A1(n3565), .A2(n3564), .A3(n3563), .A4(n3562), .ZN(n3454)
         );
  OR2_X1 U3857 ( .A1(n4473), .A2(n4472), .ZN(n3456) );
  NAND2_X1 U3858 ( .A1(n4289), .A2(n4290), .ZN(n4663) );
  AND2_X1 U3859 ( .A1(n3500), .A2(n3746), .ZN(n3680) );
  OAI21_X1 U3860 ( .B1(n3478), .B2(n3867), .A(n4497), .ZN(n4498) );
  AND2_X1 U3861 ( .A1(n6019), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3458)
         );
  OR2_X1 U3862 ( .A1(n4540), .A2(n4537), .ZN(n3459) );
  AND2_X1 U3863 ( .A1(n6503), .A2(n5048), .ZN(n3460) );
  AND2_X1 U3864 ( .A1(n4540), .A2(n5618), .ZN(n3461) );
  INV_X1 U3865 ( .A(n4509), .ZN(n3473) );
  CLKBUF_X3 U3866 ( .A(n4383), .Z(n4374) );
  NOR2_X1 U3867 ( .A1(n5084), .A2(n3495), .ZN(n5441) );
  NAND2_X1 U3868 ( .A1(n5652), .A2(n5651), .ZN(n5650) );
  OR2_X1 U3869 ( .A1(n5711), .A2(n5710), .ZN(n3462) );
  OAI21_X1 U3870 ( .B1(n5538), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6019), 
        .ZN(n5605) );
  NAND2_X1 U3871 ( .A1(n3653), .A2(n4460), .ZN(n4557) );
  INV_X1 U3872 ( .A(n4357), .ZN(n3745) );
  AND2_X1 U3873 ( .A1(n5908), .A2(n5907), .ZN(n5725) );
  INV_X1 U3874 ( .A(n5939), .ZN(n3498) );
  INV_X1 U3875 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6923) );
  INV_X1 U3876 ( .A(n3821), .ZN(n4976) );
  OR2_X1 U3877 ( .A1(n4874), .A2(n4357), .ZN(n4583) );
  AND2_X1 U3878 ( .A1(n4628), .A2(n4447), .ZN(n3463) );
  AND2_X1 U3879 ( .A1(n3463), .A2(n5754), .ZN(n3464) );
  AND2_X1 U3880 ( .A1(n5884), .A2(n6111), .ZN(n3465) );
  MUX2_X1 U3881 ( .A(n4374), .B(n4444), .S(EBX_REG_16__SCAN_IN), .Z(n4412) );
  MUX2_X1 U3882 ( .A(n4374), .B(n4366), .S(EBX_REG_2__SCAN_IN), .Z(n4373) );
  MUX2_X1 U3883 ( .A(n4374), .B(n4444), .S(EBX_REG_8__SCAN_IN), .Z(n4390) );
  MUX2_X1 U3884 ( .A(n4374), .B(n4444), .S(EBX_REG_10__SCAN_IN), .Z(n4397) );
  MUX2_X1 U3885 ( .A(n4374), .B(n4444), .S(EBX_REG_22__SCAN_IN), .Z(n4428) );
  MUX2_X1 U3886 ( .A(n4374), .B(n4444), .S(EBX_REG_26__SCAN_IN), .Z(n4438) );
  NOR3_X2 U3887 ( .A1(n5711), .A2(n5688), .A3(n5710), .ZN(n5908) );
  NOR2_X2 U3888 ( .A1(n5933), .A2(n5932), .ZN(n3467) );
  NOR2_X2 U3889 ( .A1(n5952), .A2(n5941), .ZN(n5943) );
  NAND2_X2 U3890 ( .A1(n3557), .A2(n3556), .ZN(n4460) );
  NAND3_X1 U3891 ( .A1(n3472), .A2(n6539), .A3(n3471), .ZN(n6538) );
  OR2_X1 U3892 ( .A1(n3473), .A2(n6532), .ZN(n3471) );
  NAND3_X1 U3893 ( .A1(n4509), .A2(n6526), .A3(n4499), .ZN(n3472) );
  OAI21_X2 U3894 ( .B1(n3477), .B2(n3476), .A(n3474), .ZN(n6014) );
  INV_X1 U3895 ( .A(n6072), .ZN(n3477) );
  NAND2_X1 U3896 ( .A1(n3898), .A2(n4574), .ZN(n3478) );
  INV_X1 U3897 ( .A(n3898), .ZN(n3479) );
  NAND2_X1 U3898 ( .A1(n3869), .A2(n3868), .ZN(n3898) );
  OAI211_X1 U3899 ( .C1(n4289), .C2(n4692), .A(n3487), .B(n3486), .ZN(n5813)
         );
  NAND3_X1 U3900 ( .A1(n4289), .A2(n4692), .A3(n3488), .ZN(n3486) );
  INV_X1 U3901 ( .A(n5766), .ZN(n3492) );
  NAND2_X1 U3902 ( .A1(n3426), .A2(n5946), .ZN(n5895) );
  INV_X1 U3903 ( .A(n5895), .ZN(n4187) );
  NAND2_X1 U3904 ( .A1(n3869), .A2(n3501), .ZN(n4500) );
  INV_X1 U3905 ( .A(n5960), .ZN(n5922) );
  NAND2_X1 U3906 ( .A1(n4485), .A2(n4821), .ZN(n6520) );
  OAI21_X1 U3907 ( .B1(n6019), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n4640), 
        .ZN(n5979) );
  AOI21_X1 U3908 ( .B1(n4639), .B2(n4638), .A(n4637), .ZN(n4642) );
  OAI21_X1 U3909 ( .B1(n6511), .B2(n6661), .A(n6512), .ZN(n4475) );
  XNOR2_X1 U3910 ( .A(n3492), .B(n3451), .ZN(n5960) );
  AND2_X1 U3911 ( .A1(n6014), .A2(n3505), .ZN(n4541) );
  AOI21_X1 U3912 ( .B1(n4888), .B2(n4028), .A(n3744), .ZN(n3799) );
  NAND2_X2 U3913 ( .A1(n4533), .A2(n4532), .ZN(n5637) );
  AND2_X1 U3914 ( .A1(n5531), .A2(n3994), .ZN(n3502) );
  AND2_X1 U3915 ( .A1(n4908), .A2(n4460), .ZN(n3503) );
  AND3_X1 U3916 ( .A1(n6132), .A2(n6156), .A3(n4539), .ZN(n3505) );
  INV_X1 U3917 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4638) );
  NOR2_X2 U3918 ( .A1(n3634), .A2(n6906), .ZN(n4028) );
  AND4_X1 U3919 ( .A1(n3574), .A2(n3573), .A3(n3572), .A4(n3571), .ZN(n3507)
         );
  AND4_X1 U3920 ( .A1(n3561), .A2(n3560), .A3(n3559), .A4(n3558), .ZN(n3508)
         );
  INV_X1 U3921 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7025) );
  INV_X1 U3922 ( .A(n5894), .ZN(n4156) );
  NOR2_X1 U3923 ( .A1(n3746), .A2(n6906), .ZN(n3870) );
  INV_X1 U3924 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5172) );
  AND2_X2 U3925 ( .A1(n6869), .A2(n4695), .ZN(n6560) );
  INV_X1 U3926 ( .A(n6507), .ZN(n5956) );
  AND2_X1 U3927 ( .A1(n6510), .A2(n5812), .ZN(n6507) );
  OR2_X1 U3928 ( .A1(n3665), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3509)
         );
  AND2_X1 U3929 ( .A1(n4625), .A2(n4624), .ZN(n3510) );
  OR2_X1 U3930 ( .A1(n4297), .A2(n5262), .ZN(n3842) );
  OR2_X1 U3931 ( .A1(n3864), .A2(n3863), .ZN(n4503) );
  INV_X1 U3932 ( .A(n4303), .ZN(n4298) );
  OR2_X1 U3933 ( .A1(n4297), .A2(n5254), .ZN(n3866) );
  NAND2_X1 U3934 ( .A1(n3735), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3736) );
  OR2_X1 U3935 ( .A1(n3888), .A2(n3887), .ZN(n4512) );
  AOI21_X1 U3936 ( .B1(n3582), .B2(INSTQUEUE_REG_6__3__SCAN_IN), .A(n3551), 
        .ZN(n3555) );
  AOI22_X1 U3937 ( .A1(n3712), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3582), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3573) );
  OR2_X1 U3938 ( .A1(n4218), .A2(n4217), .ZN(n4225) );
  OR2_X1 U3939 ( .A1(n6834), .A2(n4685), .ZN(n4121) );
  INV_X1 U3940 ( .A(n4201), .ZN(n3744) );
  NAND2_X1 U3941 ( .A1(n3654), .A2(n3658), .ZN(n3698) );
  OR2_X1 U3942 ( .A1(n4334), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4569)
         );
  INV_X1 U3943 ( .A(n3673), .ZN(n3645) );
  AND2_X1 U3944 ( .A1(n5831), .A2(n3421), .ZN(n4688) );
  INV_X1 U3945 ( .A(n4178), .ZN(n4682) );
  INV_X1 U3946 ( .A(n3870), .ZN(n3757) );
  OAI21_X1 U3947 ( .B1(n3998), .B2(n3997), .A(n3996), .ZN(n3999) );
  INV_X1 U3948 ( .A(n4886), .ZN(n3643) );
  NAND2_X1 U3949 ( .A1(n4138), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4139)
         );
  INV_X1 U3950 ( .A(n6756), .ZN(n5658) );
  AND2_X1 U3951 ( .A1(n4378), .A2(n4377), .ZN(n4844) );
  AND2_X1 U3952 ( .A1(n3982), .A2(n3981), .ZN(n3997) );
  NAND2_X1 U3953 ( .A1(n4501), .A2(n4028), .ZN(n3907) );
  NAND2_X1 U3954 ( .A1(n4850), .A2(n4374), .ZN(n4440) );
  AND2_X1 U3955 ( .A1(n4410), .A2(n4409), .ZN(n5677) );
  OAI21_X1 U3956 ( .B1(n3806), .B2(n4950), .A(n3805), .ZN(n4971) );
  AND2_X1 U3957 ( .A1(n4892), .A2(n5357), .ZN(n5170) );
  AND2_X1 U3958 ( .A1(n5821), .A2(n5816), .ZN(n4710) );
  AND2_X1 U3959 ( .A1(n4749), .A2(n4580), .ZN(n4946) );
  NOR2_X1 U3960 ( .A1(n4139), .A2(n4151), .ZN(n4188) );
  OR2_X1 U3961 ( .A1(n6802), .A2(n5681), .ZN(n5730) );
  INV_X1 U3962 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5463) );
  OR2_X1 U3963 ( .A1(n6583), .A2(n5347), .ZN(n6756) );
  NAND2_X1 U3964 ( .A1(n6583), .A2(n5364), .ZN(n6802) );
  AND2_X1 U3965 ( .A1(n4393), .A2(n4392), .ZN(n5444) );
  OR2_X1 U3966 ( .A1(n4248), .A2(n4247), .ZN(n5867) );
  NOR2_X1 U3967 ( .A1(n4067), .A2(n6064), .ZN(n4051) );
  AND2_X1 U3968 ( .A1(n4540), .A2(n6707), .ZN(n6073) );
  NOR2_X1 U3969 ( .A1(n3953), .A2(n5463), .ZN(n3967) );
  AOI21_X1 U3970 ( .B1(n5979), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5748), 
        .ZN(n4641) );
  INV_X1 U3971 ( .A(n6694), .ZN(n6674) );
  INV_X1 U3972 ( .A(n4888), .ZN(n4889) );
  AND2_X1 U3973 ( .A1(n5055), .A2(n5152), .ZN(n5183) );
  INV_X1 U3974 ( .A(n5546), .ZN(n7043) );
  INV_X1 U3975 ( .A(n5312), .ZN(n5317) );
  INV_X1 U3976 ( .A(n5372), .ZN(n5424) );
  INV_X1 U3977 ( .A(n7156), .ZN(n5325) );
  INV_X1 U3978 ( .A(n5553), .ZN(n5374) );
  INV_X1 U3979 ( .A(n6928), .ZN(n5829) );
  AND2_X1 U3980 ( .A1(n6756), .A2(n5349), .ZN(n6865) );
  AND2_X1 U3981 ( .A1(n6756), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6856) );
  INV_X1 U3982 ( .A(n6847), .ZN(n6864) );
  NOR2_X1 U3983 ( .A1(n6510), .A2(n4449), .ZN(n4450) );
  INV_X1 U3984 ( .A(n5958), .ZN(n6508) );
  NOR2_X1 U3985 ( .A1(n4757), .A2(n6928), .ZN(n4362) );
  INV_X1 U3986 ( .A(n3422), .ZN(n7080) );
  INV_X1 U3987 ( .A(n6963), .ZN(n7081) );
  AND2_X1 U3988 ( .A1(n3422), .A2(n4881), .ZN(n7078) );
  NAND2_X1 U3989 ( .A1(n5331), .A2(n4527), .ZN(n5592) );
  NAND2_X1 U3990 ( .A1(n3848), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3872)
         );
  INV_X1 U3991 ( .A(n6566), .ZN(n6548) );
  INV_X1 U3992 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4643) );
  NOR2_X1 U3993 ( .A1(n6651), .A2(n4616), .ZN(n6595) );
  NAND2_X1 U3994 ( .A1(n6538), .A2(n4518), .ZN(n5333) );
  NAND2_X1 U3995 ( .A1(n4582), .A2(n4581), .ZN(n4606) );
  INV_X1 U3996 ( .A(n6651), .ZN(n6612) );
  INV_X1 U3997 ( .A(n6702), .ZN(n6723) );
  AND2_X1 U3998 ( .A1(n5221), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6980) );
  AND2_X1 U3999 ( .A1(n5183), .A2(n6990), .ZN(n5582) );
  AND2_X1 U4000 ( .A1(n7040), .A2(n5746), .ZN(n7184) );
  INV_X1 U4001 ( .A(n4995), .ZN(n7185) );
  INV_X1 U4002 ( .A(n4994), .ZN(n7176) );
  NOR2_X1 U4003 ( .A1(n4923), .A2(n4900), .ZN(n5372) );
  INV_X1 U4004 ( .A(n7013), .ZN(n7169) );
  AND3_X1 U4005 ( .A1(n4978), .A2(n4890), .A3(n5096), .ZN(n7162) );
  NOR2_X1 U4006 ( .A1(n5222), .A2(n6990), .ZN(n7156) );
  NOR2_X2 U4007 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4887), .ZN(n5175) );
  INV_X1 U4008 ( .A(n7097), .ZN(n5554) );
  INV_X1 U4009 ( .A(n7139), .ZN(n5562) );
  INV_X1 U4010 ( .A(n7190), .ZN(n5584) );
  OR2_X1 U4011 ( .A1(n4880), .A2(n5818), .ZN(n5343) );
  NAND2_X1 U4012 ( .A1(n5343), .A2(n5342), .ZN(n6583) );
  INV_X1 U4013 ( .A(n6955), .ZN(n6938) );
  OR2_X1 U4014 ( .A1(n4590), .A2(n4448), .ZN(n6080) );
  INV_X1 U4015 ( .A(n6856), .ZN(n6854) );
  INV_X1 U4016 ( .A(n6855), .ZN(n6796) );
  AOI21_X1 U4017 ( .B1(n4451), .B2(n6507), .A(n4450), .ZN(n4452) );
  NAND2_X1 U4018 ( .A1(n6510), .A2(n3746), .ZN(n5958) );
  AND2_X1 U4019 ( .A1(n4883), .A2(n6963), .ZN(n5975) );
  INV_X1 U4020 ( .A(n6406), .ZN(n6427) );
  OR3_X1 U4021 ( .A1(n4880), .A2(READY_N), .A3(n4713), .ZN(n4877) );
  OR2_X1 U4022 ( .A1(n6560), .A2(n4813), .ZN(n6566) );
  INV_X1 U4023 ( .A(n6721), .ZN(n6709) );
  NAND2_X1 U4024 ( .A1(n4606), .A2(n4587), .ZN(n6702) );
  INV_X1 U4025 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6883) );
  INV_X1 U4026 ( .A(n5774), .ZN(n5780) );
  NOR2_X1 U4027 ( .A1(n5177), .A2(n5176), .ZN(n5219) );
  INV_X1 U4028 ( .A(n6952), .ZN(n6955) );
  NAND2_X1 U4029 ( .A1(n4453), .A2(n4452), .ZN(U2831) );
  INV_X1 U4030 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3511) );
  INV_X1 U4031 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3512) );
  INV_X1 U4032 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4033 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(n3713), .B1(n3576), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3516) );
  AND2_X4 U4034 ( .A1(n3519), .A2(n4941), .ZN(n3612) );
  AOI22_X1 U4035 ( .A1(n3699), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3612), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4036 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n3442), .B1(n3577), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3514) );
  AND2_X2 U4037 ( .A1(n3518), .A2(n6180), .ZN(n3712) );
  AOI22_X1 U4038 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n3439), .B1(n3582), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3524) );
  AOI22_X1 U4039 ( .A1(n3811), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3523) );
  AOI22_X1 U4040 ( .A1(n3617), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U4041 ( .A1(n3778), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3583), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3521) );
  NAND2_X1 U4042 ( .A1(n4072), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3530)
         );
  NAND2_X1 U4043 ( .A1(n3576), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3528) );
  NAND2_X1 U4044 ( .A1(n3612), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3527) );
  NAND2_X1 U4045 ( .A1(n3713), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3534) );
  NAND2_X1 U4046 ( .A1(n3699), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3533)
         );
  NAND2_X1 U4047 ( .A1(n3443), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3532)
         );
  NAND2_X1 U4048 ( .A1(n3603), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3531) );
  NAND2_X1 U4049 ( .A1(n3712), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3538) );
  NAND2_X1 U4050 ( .A1(n3582), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3537) );
  NAND2_X1 U4051 ( .A1(n3617), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3536) );
  NAND2_X1 U4052 ( .A1(n3778), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3535) );
  NAND2_X1 U4053 ( .A1(n3811), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3542) );
  NAND2_X1 U4054 ( .A1(n3577), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3541)
         );
  NAND2_X1 U4055 ( .A1(n3583), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3540)
         );
  NAND2_X1 U4056 ( .A1(n3714), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3539)
         );
  AOI22_X1 U4057 ( .A1(n3699), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3612), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4058 ( .A1(n3443), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3576), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4059 ( .A1(n3445), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3548) );
  AOI22_X1 U4060 ( .A1(n3811), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3547) );
  AOI22_X1 U4061 ( .A1(n3617), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3583), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4062 ( .A1(n3577), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3778), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4063 ( .A1(n3439), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3552) );
  AOI22_X1 U4064 ( .A1(n3583), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3778), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4065 ( .A1(n3617), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4066 ( .A1(n3712), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3582), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U4067 ( .A1(n3811), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3558) );
  AOI22_X1 U4068 ( .A1(n3699), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3612), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4069 ( .A1(n3713), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3576), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4070 ( .A1(n3719), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3577), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3562) );
  NAND2_X2 U4071 ( .A1(n3508), .A2(n3454), .ZN(n3676) );
  NAND2_X1 U4072 ( .A1(n3500), .A2(n4908), .ZN(n3566) );
  NOR2_X1 U4073 ( .A1(n4557), .A2(n3566), .ZN(n3590) );
  NAND2_X1 U4074 ( .A1(n5155), .A2(n3634), .ZN(n3575) );
  AOI22_X1 U4075 ( .A1(n3699), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3612), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4076 ( .A1(n3719), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3617), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4077 ( .A1(n3811), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3778), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3567) );
  AOI22_X1 U4078 ( .A1(n4072), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3713), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3574) );
  AOI22_X1 U4079 ( .A1(n3577), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3572) );
  AOI22_X1 U4080 ( .A1(n3583), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3571) );
  AOI22_X1 U4081 ( .A1(n3713), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3576), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4082 ( .A1(n3699), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3612), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3579) );
  AOI22_X1 U4083 ( .A1(n3719), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3577), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3578) );
  AND4_X2 U4084 ( .A1(n3581), .A2(n3580), .A3(n3579), .A4(n3578), .ZN(n3588)
         );
  AOI22_X1 U4085 ( .A1(n3712), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3582), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4086 ( .A1(n3778), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3583), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4087 ( .A1(n3811), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3714), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3584) );
  INV_X1 U4088 ( .A(n4350), .ZN(n3589) );
  NAND2_X1 U4089 ( .A1(n3590), .A2(n3589), .ZN(n4354) );
  NAND2_X1 U4090 ( .A1(n3699), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3594)
         );
  NAND2_X1 U4091 ( .A1(n3445), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3593)
         );
  NAND2_X1 U4092 ( .A1(n3612), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3592) );
  NAND2_X1 U4093 ( .A1(n3441), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3591) );
  NAND2_X1 U4094 ( .A1(n3811), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3598) );
  NAND2_X1 U4095 ( .A1(n3712), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3597) );
  NAND2_X1 U4096 ( .A1(n3582), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3596) );
  NAND2_X1 U4097 ( .A1(n3714), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3595)
         );
  NAND2_X1 U4098 ( .A1(n3713), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3602) );
  NAND2_X1 U4099 ( .A1(n3719), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3601)
         );
  NAND2_X1 U4100 ( .A1(n3576), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3600) );
  NAND2_X1 U4101 ( .A1(n3577), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3599)
         );
  NAND2_X1 U4102 ( .A1(n3617), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3607) );
  NAND2_X1 U4103 ( .A1(n3603), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3606) );
  NAND2_X1 U4104 ( .A1(n3699), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3616)
         );
  NAND2_X1 U4105 ( .A1(n4072), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3615)
         );
  NAND2_X1 U4106 ( .A1(n3612), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3614) );
  NAND2_X1 U4107 ( .A1(n3576), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3613) );
  NAND2_X1 U4108 ( .A1(n3719), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3621)
         );
  NAND2_X1 U4109 ( .A1(n3582), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3620) );
  NAND2_X1 U4110 ( .A1(n3617), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3619) );
  NAND2_X1 U4111 ( .A1(n3583), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3618)
         );
  NAND2_X1 U4112 ( .A1(n3713), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3625) );
  NAND2_X1 U4113 ( .A1(n3577), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3623)
         );
  NAND2_X1 U4114 ( .A1(n3603), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3622) );
  NAND2_X1 U4115 ( .A1(n3712), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3629) );
  NAND2_X1 U4116 ( .A1(n3811), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3628) );
  NAND2_X1 U4117 ( .A1(n3714), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3627)
         );
  NAND2_X1 U4118 ( .A1(n3778), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3626) );
  NAND4_X4 U4119 ( .A1(n3633), .A2(n3632), .A3(n3631), .A4(n3630), .ZN(n3659)
         );
  INV_X1 U4120 ( .A(n3654), .ZN(n3635) );
  NAND2_X1 U4121 ( .A1(n3660), .A2(n3676), .ZN(n3638) );
  NAND2_X1 U4122 ( .A1(n3636), .A2(n4908), .ZN(n3637) );
  NAND3_X1 U4123 ( .A1(n3745), .A2(n3638), .A3(n3637), .ZN(n3640) );
  NOR2_X2 U4124 ( .A1(n3676), .A2(n5160), .ZN(n3639) );
  NAND2_X2 U4125 ( .A1(n3680), .A2(n3639), .ZN(n6183) );
  INV_X1 U4126 ( .A(n3672), .ZN(n3642) );
  OR2_X1 U4127 ( .A1(n3660), .A2(n3447), .ZN(n4558) );
  INV_X1 U4128 ( .A(n4558), .ZN(n4596) );
  INV_X1 U4129 ( .A(n4354), .ZN(n3644) );
  NAND2_X1 U4130 ( .A1(n3644), .A2(n3658), .ZN(n4706) );
  NAND2_X1 U4131 ( .A1(n3446), .A2(n5155), .ZN(n4360) );
  INV_X1 U4132 ( .A(n4360), .ZN(n3646) );
  NAND2_X1 U4133 ( .A1(n3646), .A2(n3645), .ZN(n4874) );
  OAI21_X2 U4134 ( .B1(n4584), .B2(n3647), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3666) );
  INV_X1 U4135 ( .A(n3666), .ZN(n3649) );
  INV_X1 U4136 ( .A(n7041), .ZN(n3648) );
  NAND2_X1 U4137 ( .A1(n5172), .A2(n7025), .ZN(n5052) );
  NAND2_X1 U4138 ( .A1(n3648), .A2(n5052), .ZN(n5227) );
  NAND2_X1 U4139 ( .A1(n5348), .A2(n6916), .ZN(n6910) );
  OAI22_X1 U4140 ( .A1(n5227), .A2(n4694), .B1(n4358), .B2(n5172), .ZN(n3665)
         );
  NAND2_X1 U4141 ( .A1(n3649), .A2(n3509), .ZN(n3668) );
  NAND2_X1 U4142 ( .A1(n4351), .A2(n5160), .ZN(n3651) );
  NAND2_X1 U4143 ( .A1(n3651), .A2(n3650), .ZN(n3682) );
  INV_X1 U4144 ( .A(n3682), .ZN(n3652) );
  NAND2_X1 U4145 ( .A1(n3652), .A2(n3503), .ZN(n4346) );
  INV_X1 U4146 ( .A(n6942), .ZN(n3655) );
  NAND2_X1 U4147 ( .A1(n3683), .A2(n3656), .ZN(n3657) );
  NAND2_X1 U4148 ( .A1(n3672), .A2(n4886), .ZN(n3662) );
  NAND2_X1 U4149 ( .A1(n4350), .A2(n3679), .ZN(n3661) );
  NAND3_X1 U4150 ( .A1(n3663), .A2(n3662), .A3(n3688), .ZN(n3664) );
  NAND2_X1 U4151 ( .A1(n3667), .A2(n3666), .ZN(n3690) );
  NAND2_X1 U4152 ( .A1(n3691), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3671) );
  INV_X1 U4153 ( .A(n4358), .ZN(n3803) );
  INV_X1 U4154 ( .A(n4694), .ZN(n3804) );
  MUX2_X1 U4155 ( .A(n3803), .B(n3804), .S(n7025), .Z(n3669) );
  NAND2_X1 U4156 ( .A1(n3660), .A2(n4886), .ZN(n3674) );
  NAND2_X1 U4157 ( .A1(n3674), .A2(n3673), .ZN(n3675) );
  NAND2_X1 U4158 ( .A1(n3672), .A2(n3675), .ZN(n4747) );
  INV_X1 U4159 ( .A(n4460), .ZN(n4905) );
  NAND2_X1 U4160 ( .A1(n3676), .A2(n3658), .ZN(n3677) );
  INV_X1 U4161 ( .A(n6910), .ZN(n5775) );
  NAND3_X1 U4162 ( .A1(n3677), .A2(n5775), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3678) );
  AOI21_X1 U4163 ( .B1(n4905), .B2(n3673), .A(n3678), .ZN(n3687) );
  AOI22_X1 U4164 ( .A1(n4351), .A2(n6581), .B1(n3680), .B2(n3446), .ZN(n3686)
         );
  INV_X1 U4165 ( .A(n3683), .ZN(n3684) );
  OAI21_X1 U4166 ( .B1(n3682), .B2(n3684), .A(n3659), .ZN(n3685) );
  NAND2_X1 U4167 ( .A1(n4747), .A2(n3689), .ZN(n3731) );
  AND2_X2 U4168 ( .A1(n3732), .A2(n3731), .ZN(n3730) );
  OAI21_X2 U4169 ( .B1(n3711), .B2(n3730), .A(n3690), .ZN(n3696) );
  INV_X1 U4170 ( .A(n3696), .ZN(n3694) );
  NAND2_X1 U4171 ( .A1(n7041), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4918) );
  OAI21_X1 U4172 ( .B1(n7041), .B2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(n4918), 
        .ZN(n4993) );
  OAI22_X1 U4173 ( .A1(n4993), .A2(n4694), .B1(n4358), .B2(n6883), .ZN(n3692)
         );
  NAND2_X1 U4174 ( .A1(n3696), .A2(n3695), .ZN(n3697) );
  AOI22_X1 U4175 ( .A1(n4673), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4645), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4176 ( .A1(n3712), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4666), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4177 ( .A1(n3443), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4178 ( .A1(n3423), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3700) );
  NAND4_X1 U4179 ( .A1(n3703), .A2(n3702), .A3(n3701), .A4(n3700), .ZN(n3709)
         );
  AOI22_X1 U4180 ( .A1(n3445), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3707) );
  AOI22_X1 U4181 ( .A1(n4267), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4182 ( .A1(n3448), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4183 ( .A1(n3773), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3704) );
  NAND4_X1 U4184 ( .A1(n3707), .A2(n3706), .A3(n3705), .A4(n3704), .ZN(n3708)
         );
  AOI22_X1 U4185 ( .A1(n4329), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4340), 
        .B2(n4476), .ZN(n3710) );
  OAI21_X2 U4186 ( .B1(n4892), .B2(STATE2_REG_0__SCAN_IN), .A(n3710), .ZN(
        n3742) );
  INV_X1 U4187 ( .A(n3742), .ZN(n3741) );
  NAND2_X1 U4188 ( .A1(n4893), .A2(n6923), .ZN(n3729) );
  AOI22_X1 U4189 ( .A1(n3439), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4666), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4190 ( .A1(n4673), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3717) );
  BUF_X1 U4191 ( .A(n3713), .Z(n4645) );
  AOI22_X1 U4192 ( .A1(n4645), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4193 ( .A1(n3424), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3715) );
  NAND4_X1 U4194 ( .A1(n3718), .A2(n3717), .A3(n3716), .A4(n3715), .ZN(n3725)
         );
  AOI22_X1 U4195 ( .A1(n4072), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3719), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4197 ( .A1(n4267), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4198 ( .A1(n3773), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4199 ( .A1(n3448), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3720) );
  NAND4_X1 U4200 ( .A1(n3723), .A2(n3722), .A3(n3721), .A4(n3720), .ZN(n3724)
         );
  INV_X1 U4201 ( .A(n4454), .ZN(n3726) );
  NOR2_X1 U4202 ( .A1(n3726), .A2(n3654), .ZN(n3727) );
  NAND2_X1 U4203 ( .A1(n3792), .A2(n6923), .ZN(n3737) );
  NAND2_X1 U4204 ( .A1(n4886), .A2(n4454), .ZN(n3734) );
  AND2_X1 U4205 ( .A1(n3734), .A2(n3654), .ZN(n3735) );
  NAND2_X1 U4206 ( .A1(n4329), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3738) );
  NAND2_X1 U4207 ( .A1(n3754), .A2(n3755), .ZN(n3740) );
  NAND2_X1 U4208 ( .A1(n3743), .A2(n3742), .ZN(n3822) );
  INV_X2 U4209 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6906) );
  INV_X1 U4210 ( .A(n4028), .ZN(n4018) );
  NAND2_X1 U4211 ( .A1(n6906), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4201) );
  INV_X1 U4212 ( .A(n3799), .ZN(n3753) );
  NAND2_X1 U4213 ( .A1(n3793), .A2(n5774), .ZN(n3751) );
  INV_X1 U4214 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3748) );
  NAND2_X1 U4215 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3824) );
  OAI21_X1 U4216 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3824), .ZN(n6517) );
  NAND2_X1 U4217 ( .A1(n3421), .A2(n6517), .ZN(n3747) );
  OAI21_X1 U4218 ( .B1(n3748), .B2(n4201), .A(n3747), .ZN(n3749) );
  AOI21_X1 U4219 ( .B1(n4691), .B2(EAX_REG_2__SCAN_IN), .A(n3749), .ZN(n3750)
         );
  AND2_X1 U4220 ( .A1(n3751), .A2(n3750), .ZN(n3798) );
  INV_X1 U4221 ( .A(n3798), .ZN(n3752) );
  NAND2_X1 U4222 ( .A1(n3753), .A2(n3752), .ZN(n3797) );
  INV_X1 U4223 ( .A(n3754), .ZN(n3756) );
  NAND2_X1 U4224 ( .A1(n4890), .A2(n4028), .ZN(n3761) );
  AOI22_X1 U4225 ( .A1(n4691), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6906), .ZN(n3759) );
  NAND2_X1 U4226 ( .A1(n3793), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3758) );
  AND2_X1 U4227 ( .A1(n3759), .A2(n3758), .ZN(n3760) );
  NAND2_X1 U4228 ( .A1(n3761), .A2(n3760), .ZN(n4853) );
  INV_X1 U4229 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5067) );
  AOI22_X1 U4230 ( .A1(n3576), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4231 ( .A1(n3712), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3582), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4232 ( .A1(n4645), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4233 ( .A1(n3603), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3763) );
  NAND4_X1 U4234 ( .A1(n3766), .A2(n3765), .A3(n3764), .A4(n3763), .ZN(n3772)
         );
  AOI22_X1 U4235 ( .A1(n3445), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3719), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4236 ( .A1(n4673), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3612), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4237 ( .A1(n3448), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3768) );
  AOI22_X1 U4238 ( .A1(n3424), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3767) );
  NAND4_X1 U4239 ( .A1(n3770), .A2(n3769), .A3(n3768), .A4(n3767), .ZN(n3771)
         );
  OR2_X1 U4240 ( .A1(n3772), .A2(n3771), .ZN(n4462) );
  AOI21_X1 U4241 ( .B1(n4886), .B2(n4462), .A(n6923), .ZN(n3786) );
  AOI22_X1 U4242 ( .A1(n4072), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4645), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4243 ( .A1(n3423), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3582), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4244 ( .A1(n3612), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4245 ( .A1(n3773), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3774) );
  NAND4_X1 U4246 ( .A1(n3777), .A2(n3776), .A3(n3775), .A4(n3774), .ZN(n3785)
         );
  AOI22_X1 U4247 ( .A1(n4673), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4248 ( .A1(n3448), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4249 ( .A1(n3443), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4250 ( .A1(n3439), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3780) );
  NAND4_X1 U4251 ( .A1(n3783), .A2(n3782), .A3(n3781), .A4(n3780), .ZN(n3784)
         );
  NAND2_X1 U4252 ( .A1(n5160), .A2(n4523), .ZN(n4520) );
  OAI211_X1 U4253 ( .C1(n4297), .C2(n5067), .A(n3786), .B(n4520), .ZN(n3790)
         );
  INV_X1 U4254 ( .A(n4523), .ZN(n3787) );
  XNOR2_X1 U4255 ( .A(n3787), .B(n4462), .ZN(n3788) );
  NAND3_X1 U4256 ( .A1(n3788), .A2(STATE2_REG_0__SCAN_IN), .A3(n5160), .ZN(
        n3789) );
  XNOR2_X1 U4257 ( .A(n3790), .B(n3789), .ZN(n3791) );
  AOI21_X1 U4258 ( .B1(n5746), .B2(n3680), .A(n6906), .ZN(n4815) );
  INV_X1 U4259 ( .A(n3792), .ZN(n5093) );
  INV_X1 U4260 ( .A(n3793), .ZN(n3847) );
  NAND2_X1 U4261 ( .A1(n6906), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3795)
         );
  NAND2_X1 U4262 ( .A1(n3870), .A2(EAX_REG_0__SCAN_IN), .ZN(n3794) );
  OAI211_X1 U4263 ( .C1(n3847), .C2(n3511), .A(n3795), .B(n3794), .ZN(n3796)
         );
  AOI21_X1 U4264 ( .B1(n5093), .B2(n4028), .A(n3796), .ZN(n4816) );
  MUX2_X1 U4265 ( .A(n4815), .B(n3421), .S(n4816), .Z(n4852) );
  NAND2_X1 U4266 ( .A1(n4853), .A2(n4852), .ZN(n4851) );
  NAND2_X1 U4267 ( .A1(n3797), .A2(n4851), .ZN(n3800) );
  NAND2_X1 U4268 ( .A1(n3799), .A2(n3798), .ZN(n4837) );
  NAND2_X1 U4269 ( .A1(n3800), .A2(n4837), .ZN(n4831) );
  INV_X1 U4270 ( .A(n3822), .ZN(n3820) );
  INV_X1 U4271 ( .A(n3691), .ZN(n3806) );
  NAND2_X1 U4272 ( .A1(n4918), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3802) );
  INV_X1 U4273 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6889) );
  NAND2_X1 U4274 ( .A1(n6889), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n7024) );
  INV_X1 U4275 ( .A(n7024), .ZN(n3801) );
  NAND2_X1 U4276 ( .A1(n7041), .A2(n3801), .ZN(n5315) );
  NAND2_X1 U4277 ( .A1(n3802), .A2(n5315), .ZN(n5228) );
  AOI22_X1 U4278 ( .A1(n5228), .A2(n3804), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3803), .ZN(n3805) );
  XNOR2_X1 U4279 ( .A(n3431), .B(n4971), .ZN(n4891) );
  NAND2_X1 U4280 ( .A1(n4891), .A2(n6923), .ZN(n3819) );
  AOI22_X1 U4281 ( .A1(n4673), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4267), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4282 ( .A1(n4072), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4283 ( .A1(n4645), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4284 ( .A1(n3443), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3807) );
  NAND4_X1 U4285 ( .A1(n3810), .A2(n3809), .A3(n3808), .A4(n3807), .ZN(n3817)
         );
  AOI22_X1 U4286 ( .A1(n3439), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4666), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4287 ( .A1(n3448), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4288 ( .A1(n3425), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4289 ( .A1(n3424), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3812) );
  NAND4_X1 U4290 ( .A1(n3815), .A2(n3814), .A3(n3813), .A4(n3812), .ZN(n3816)
         );
  AOI22_X1 U4291 ( .A1(n4329), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4340), 
        .B2(n4480), .ZN(n3818) );
  NAND2_X1 U4292 ( .A1(n4976), .A2(n3822), .ZN(n3823) );
  NAND2_X1 U4293 ( .A1(n3854), .A2(n3823), .ZN(n4482) );
  INV_X2 U4294 ( .A(n4482), .ZN(n4978) );
  INV_X1 U4295 ( .A(n3848), .ZN(n3827) );
  INV_X1 U4296 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3825) );
  NAND2_X1 U4297 ( .A1(n3825), .A2(n3824), .ZN(n3826) );
  NAND2_X1 U4298 ( .A1(n3827), .A2(n3826), .ZN(n5483) );
  AOI22_X1 U4299 ( .A1(n5483), .A2(n3421), .B1(n3744), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3829) );
  NAND2_X1 U4300 ( .A1(n3870), .A2(EAX_REG_3__SCAN_IN), .ZN(n3828) );
  OAI211_X1 U4301 ( .C1(n3847), .C2(n4950), .A(n3829), .B(n3828), .ZN(n3830)
         );
  INV_X1 U4302 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5262) );
  AOI22_X1 U4303 ( .A1(n4673), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4267), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4304 ( .A1(n3445), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4305 ( .A1(n4645), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4306 ( .A1(n3719), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3831) );
  NAND4_X1 U4307 ( .A1(n3834), .A2(n3833), .A3(n3832), .A4(n3831), .ZN(n3840)
         );
  AOI22_X1 U4308 ( .A1(n3712), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4666), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4309 ( .A1(n3448), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4310 ( .A1(n3425), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4311 ( .A1(n3423), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3835) );
  NAND4_X1 U4312 ( .A1(n3838), .A2(n3837), .A3(n3836), .A4(n3835), .ZN(n3839)
         );
  NAND2_X1 U4313 ( .A1(n4340), .A2(n4493), .ZN(n3841) );
  INV_X1 U4314 ( .A(n3853), .ZN(n3843) );
  NAND2_X1 U4315 ( .A1(n4486), .A2(n4028), .ZN(n3852) );
  INV_X1 U4316 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3846) );
  NAND2_X1 U4317 ( .A1(n6906), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3845)
         );
  NAND2_X1 U4318 ( .A1(n3870), .A2(EAX_REG_4__SCAN_IN), .ZN(n3844) );
  OAI211_X1 U4319 ( .C1(n3847), .C2(n3846), .A(n3845), .B(n3844), .ZN(n3850)
         );
  OAI21_X1 U4320 ( .B1(n3848), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3872), 
        .ZN(n6745) );
  AND2_X1 U4321 ( .A1(n6745), .A2(n3421), .ZN(n3849) );
  AOI21_X1 U4322 ( .B1(n3850), .B2(n4685), .A(n3849), .ZN(n3851) );
  NAND2_X1 U4323 ( .A1(n3852), .A2(n3851), .ZN(n4841) );
  NAND2_X1 U4324 ( .A1(n4843), .A2(n4841), .ZN(n5044) );
  INV_X1 U4325 ( .A(n5044), .ZN(n3878) );
  NOR2_X2 U4326 ( .A1(n3854), .A2(n3853), .ZN(n3869) );
  INV_X1 U4327 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5254) );
  AOI22_X1 U4328 ( .A1(n4231), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4329 ( .A1(n4645), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3719), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4330 ( .A1(n4267), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4331 ( .A1(n4650), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3855) );
  NAND4_X1 U4332 ( .A1(n3858), .A2(n3857), .A3(n3856), .A4(n3855), .ZN(n3864)
         );
  AOI22_X1 U4333 ( .A1(n4673), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3424), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4334 ( .A1(n3425), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4335 ( .A1(n4072), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4336 ( .A1(n4666), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3859) );
  NAND4_X1 U4337 ( .A1(n3862), .A2(n3861), .A3(n3860), .A4(n3859), .ZN(n3863)
         );
  NAND2_X1 U4338 ( .A1(n4340), .A2(n4503), .ZN(n3865) );
  NAND2_X1 U4339 ( .A1(n3866), .A2(n3865), .ZN(n3868) );
  NOR2_X1 U4340 ( .A1(n3869), .A2(n3868), .ZN(n3867) );
  INV_X1 U4341 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3875) );
  AND2_X1 U4342 ( .A1(n3872), .A2(n3871), .ZN(n3873) );
  OR2_X1 U4343 ( .A1(n3873), .A2(n3901), .ZN(n6760) );
  AOI22_X1 U4344 ( .A1(n6760), .A2(n3421), .B1(n3744), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3874) );
  OAI21_X1 U4345 ( .B1(n3757), .B2(n3875), .A(n3874), .ZN(n3876) );
  NAND2_X1 U4346 ( .A1(n3878), .A2(n3877), .ZN(n5041) );
  INV_X1 U4347 ( .A(n5041), .ZN(n3909) );
  INV_X1 U4348 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5075) );
  OR2_X1 U4349 ( .A1(n4297), .A2(n5075), .ZN(n3890) );
  AOI22_X1 U4350 ( .A1(n4673), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4267), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4351 ( .A1(n3445), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4352 ( .A1(n4645), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4353 ( .A1(n3719), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3879) );
  NAND4_X1 U4354 ( .A1(n3882), .A2(n3881), .A3(n3880), .A4(n3879), .ZN(n3888)
         );
  AOI22_X1 U4355 ( .A1(n3439), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4666), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4356 ( .A1(n3448), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4357 ( .A1(n3425), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4358 ( .A1(n3423), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3883) );
  NAND4_X1 U4359 ( .A1(n3886), .A2(n3885), .A3(n3884), .A4(n3883), .ZN(n3887)
         );
  NAND2_X1 U4360 ( .A1(n4340), .A2(n4512), .ZN(n3889) );
  NAND2_X1 U4361 ( .A1(n3890), .A2(n3889), .ZN(n3899) );
  INV_X1 U4362 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5071) );
  NAND2_X1 U4363 ( .A1(n4340), .A2(n4523), .ZN(n3891) );
  OAI21_X1 U4364 ( .B1(n4297), .B2(n5071), .A(n3891), .ZN(n3892) );
  NAND2_X1 U4365 ( .A1(n4510), .A2(n4028), .ZN(n3897) );
  NAND2_X1 U4366 ( .A1(n3903), .A2(n6771), .ZN(n3893) );
  NAND2_X1 U4367 ( .A1(n3925), .A2(n3893), .ZN(n6784) );
  NAND2_X1 U4368 ( .A1(n6784), .A2(n3421), .ZN(n3894) );
  OAI21_X1 U4369 ( .B1(n6771), .B2(n4201), .A(n3894), .ZN(n3895) );
  AOI21_X1 U4370 ( .B1(n3870), .B2(EAX_REG_7__SCAN_IN), .A(n3895), .ZN(n3896)
         );
  NAND2_X1 U4371 ( .A1(n3897), .A2(n3896), .ZN(n5086) );
  INV_X1 U4372 ( .A(n3899), .ZN(n3900) );
  OR2_X1 U4373 ( .A1(n3901), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3902) );
  NAND2_X1 U4374 ( .A1(n3903), .A2(n3902), .ZN(n6765) );
  INV_X1 U4375 ( .A(n6765), .ZN(n3905) );
  AOI22_X1 U4376 ( .A1(n4691), .A2(EAX_REG_6__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6906), .ZN(n3904) );
  MUX2_X1 U4377 ( .A(n3905), .B(n3904), .S(n4685), .Z(n3906) );
  AOI22_X1 U4378 ( .A1(n4673), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4267), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4379 ( .A1(n3443), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4380 ( .A1(n3448), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4381 ( .A1(n4666), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3910) );
  NAND4_X1 U4382 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3919)
         );
  AOI22_X1 U4383 ( .A1(n4645), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4384 ( .A1(n3424), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4231), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4385 ( .A1(n4072), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4386 ( .A1(n3425), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3914) );
  NAND4_X1 U4387 ( .A1(n3917), .A2(n3916), .A3(n3915), .A4(n3914), .ZN(n3918)
         );
  OAI21_X1 U4388 ( .B1(n3919), .B2(n3918), .A(n4028), .ZN(n3924) );
  NAND2_X1 U4389 ( .A1(n3870), .A2(EAX_REG_8__SCAN_IN), .ZN(n3923) );
  INV_X1 U4390 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3920) );
  XNOR2_X1 U4391 ( .A(n3925), .B(n3920), .ZN(n5511) );
  NAND2_X1 U4392 ( .A1(n5511), .A2(n3421), .ZN(n3922) );
  NAND2_X1 U4393 ( .A1(n3744), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3921)
         );
  XOR2_X1 U4394 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3949), .Z(n6793) );
  AOI22_X1 U4395 ( .A1(n4673), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4267), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4396 ( .A1(n3423), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4231), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4397 ( .A1(n4650), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4398 ( .A1(n3448), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3926) );
  NAND4_X1 U4399 ( .A1(n3929), .A2(n3928), .A3(n3927), .A4(n3926), .ZN(n3935)
         );
  AOI22_X1 U4400 ( .A1(n4072), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4645), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4401 ( .A1(n3719), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4402 ( .A1(n3425), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4403 ( .A1(n4666), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3930) );
  NAND4_X1 U4404 ( .A1(n3933), .A2(n3932), .A3(n3931), .A4(n3930), .ZN(n3934)
         );
  OR2_X1 U4405 ( .A1(n3935), .A2(n3934), .ZN(n3936) );
  AOI22_X1 U4406 ( .A1(n4028), .A2(n3936), .B1(n3744), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3938) );
  NAND2_X1 U4407 ( .A1(n3870), .A2(EAX_REG_9__SCAN_IN), .ZN(n3937) );
  OAI211_X1 U4408 ( .C1(n6793), .C2(n4685), .A(n3938), .B(n3937), .ZN(n5443)
         );
  AOI22_X1 U4409 ( .A1(n4673), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4410 ( .A1(n4231), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4666), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4411 ( .A1(n3443), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4412 ( .A1(n3424), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3939) );
  NAND4_X1 U4413 ( .A1(n3942), .A2(n3941), .A3(n3940), .A4(n3939), .ZN(n3948)
         );
  AOI22_X1 U4414 ( .A1(n3445), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4267), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4415 ( .A1(n4645), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4416 ( .A1(n3448), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4417 ( .A1(n3425), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3943) );
  NAND4_X1 U4418 ( .A1(n3946), .A2(n3945), .A3(n3944), .A4(n3943), .ZN(n3947)
         );
  NOR2_X1 U4419 ( .A1(n3948), .A2(n3947), .ZN(n3952) );
  XNOR2_X1 U4420 ( .A(n3953), .B(n5463), .ZN(n5541) );
  NAND2_X1 U4421 ( .A1(n5541), .A2(n3421), .ZN(n3951) );
  AOI22_X1 U4422 ( .A1(n4691), .A2(EAX_REG_10__SCAN_IN), .B1(n3744), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3950) );
  OAI211_X1 U4423 ( .C1(n3952), .C2(n4018), .A(n3951), .B(n3950), .ZN(n5460)
         );
  XOR2_X1 U4424 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3967), .Z(n6547) );
  AOI22_X1 U4425 ( .A1(n4267), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4426 ( .A1(n3423), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4666), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4427 ( .A1(n3448), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4428 ( .A1(n4667), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3954) );
  NAND4_X1 U4429 ( .A1(n3957), .A2(n3956), .A3(n3955), .A4(n3954), .ZN(n3963)
         );
  AOI22_X1 U4430 ( .A1(n4072), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4673), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4431 ( .A1(n4645), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4432 ( .A1(n3719), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4433 ( .A1(n4231), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3958) );
  NAND4_X1 U4434 ( .A1(n3961), .A2(n3960), .A3(n3959), .A4(n3958), .ZN(n3962)
         );
  OR2_X1 U4435 ( .A1(n3963), .A2(n3962), .ZN(n3964) );
  AOI22_X1 U4436 ( .A1(n4028), .A2(n3964), .B1(n3744), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3966) );
  NAND2_X1 U4437 ( .A1(n3870), .A2(EAX_REG_11__SCAN_IN), .ZN(n3965) );
  OAI211_X1 U4438 ( .C1(n6547), .C2(n4685), .A(n3966), .B(n3965), .ZN(n5494)
         );
  INV_X1 U4439 ( .A(n3998), .ZN(n3995) );
  INV_X1 U4440 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3968) );
  XNOR2_X1 U4441 ( .A(n4000), .B(n3968), .ZN(n5614) );
  AOI21_X1 U4442 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n3968), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3970) );
  AND2_X1 U4443 ( .A1(n3870), .A2(EAX_REG_12__SCAN_IN), .ZN(n3969) );
  OAI22_X1 U4444 ( .A1(n5614), .A2(n4685), .B1(n3970), .B2(n3969), .ZN(n3982)
         );
  AOI22_X1 U4445 ( .A1(n4650), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U4446 ( .A1(n4231), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4666), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4447 ( .A1(n3444), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4448 ( .A1(n3425), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3971) );
  NAND4_X1 U4449 ( .A1(n3974), .A2(n3973), .A3(n3972), .A4(n3971), .ZN(n3980)
         );
  AOI22_X1 U4450 ( .A1(n4645), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3719), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4451 ( .A1(n4673), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4267), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4452 ( .A1(n3773), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4453 ( .A1(n3424), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3975) );
  NAND4_X1 U4454 ( .A1(n3978), .A2(n3977), .A3(n3976), .A4(n3975), .ZN(n3979)
         );
  OAI21_X1 U4455 ( .B1(n3980), .B2(n3979), .A(n4028), .ZN(n3981) );
  INV_X1 U4456 ( .A(n3997), .ZN(n5531) );
  AOI22_X1 U4457 ( .A1(n4673), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U4458 ( .A1(n4072), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4459 ( .A1(n4645), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4460 ( .A1(n4231), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3983) );
  NAND4_X1 U4461 ( .A1(n3986), .A2(n3985), .A3(n3984), .A4(n3983), .ZN(n3992)
         );
  AOI22_X1 U4462 ( .A1(n3423), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4666), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U4463 ( .A1(n3443), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4267), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U4464 ( .A1(n3448), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U4465 ( .A1(n3425), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3987) );
  NAND4_X1 U4466 ( .A1(n3990), .A2(n3989), .A3(n3988), .A4(n3987), .ZN(n3991)
         );
  OR2_X1 U4467 ( .A1(n3992), .A2(n3991), .ZN(n3993) );
  NAND2_X1 U4468 ( .A1(n4028), .A2(n3993), .ZN(n3996) );
  INV_X1 U4469 ( .A(n3996), .ZN(n3994) );
  NAND2_X1 U4470 ( .A1(n4691), .A2(EAX_REG_13__SCAN_IN), .ZN(n4003) );
  OAI21_X1 U4471 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n4001), .A(n4019), 
        .ZN(n6813) );
  AOI22_X1 U4472 ( .A1(n3421), .A2(n6813), .B1(n3744), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4002) );
  NAND2_X1 U4473 ( .A1(n4003), .A2(n4002), .ZN(n5629) );
  NAND2_X1 U4474 ( .A1(n5628), .A2(n5629), .ZN(n5632) );
  AOI22_X1 U4475 ( .A1(n3444), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4673), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4476 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(n4666), .B1(n3423), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4007) );
  AOI22_X1 U4477 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n3773), .B1(n4667), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4478 ( .A1(n3425), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4005) );
  NAND4_X1 U4479 ( .A1(n4008), .A2(n4007), .A3(n4006), .A4(n4005), .ZN(n4014)
         );
  AOI22_X1 U4480 ( .A1(n4645), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4481 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n4231), .B1(n3448), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4482 ( .A1(n4267), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U4483 ( .A1(n3443), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4009) );
  NAND4_X1 U4484 ( .A1(n4012), .A2(n4011), .A3(n4010), .A4(n4009), .ZN(n4013)
         );
  NOR2_X1 U4485 ( .A1(n4014), .A2(n4013), .ZN(n4017) );
  XNOR2_X1 U4486 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4019), .ZN(n5668)
         );
  INV_X1 U4487 ( .A(n5668), .ZN(n5656) );
  AOI22_X1 U4488 ( .A1(n3744), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n3421), 
        .B2(n5656), .ZN(n4016) );
  NAND2_X1 U4489 ( .A1(n4691), .A2(EAX_REG_14__SCAN_IN), .ZN(n4015) );
  OAI211_X1 U4490 ( .C1(n4018), .C2(n4017), .A(n4016), .B(n4015), .ZN(n5651)
         );
  INV_X1 U4491 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5660) );
  XNOR2_X1 U4492 ( .A(n4036), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5701)
         );
  AOI22_X1 U4493 ( .A1(n3443), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U4494 ( .A1(n4231), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4666), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U4495 ( .A1(n4673), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U4496 ( .A1(n3425), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4020) );
  NAND4_X1 U4497 ( .A1(n4023), .A2(n4022), .A3(n4021), .A4(n4020), .ZN(n4030)
         );
  AOI22_X1 U4498 ( .A1(n3445), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4267), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U4499 ( .A1(n3713), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U4500 ( .A1(n3448), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U4501 ( .A1(n3423), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4024) );
  NAND4_X1 U4502 ( .A1(n4027), .A2(n4026), .A3(n4025), .A4(n4024), .ZN(n4029)
         );
  OAI21_X1 U4503 ( .B1(n4030), .B2(n4029), .A(n4028), .ZN(n4033) );
  NAND2_X1 U4504 ( .A1(n4691), .A2(EAX_REG_15__SCAN_IN), .ZN(n4032) );
  NAND2_X1 U4505 ( .A1(n3744), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4031)
         );
  NAND3_X1 U4506 ( .A1(n4033), .A2(n4032), .A3(n4031), .ZN(n4034) );
  AOI21_X1 U4507 ( .B1(n5701), .B2(n3421), .A(n4034), .ZN(n5676) );
  XNOR2_X1 U4508 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n4050), .ZN(n6077)
         );
  INV_X1 U4509 ( .A(n6183), .ZN(n4575) );
  NAND2_X1 U4510 ( .A1(n4575), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4178) );
  AOI22_X1 U4511 ( .A1(n3445), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4267), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U4512 ( .A1(n3713), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U4513 ( .A1(n3719), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U4514 ( .A1(n3423), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4037) );
  NAND4_X1 U4515 ( .A1(n4040), .A2(n4039), .A3(n4038), .A4(n4037), .ZN(n4046)
         );
  AOI22_X1 U4516 ( .A1(n4231), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3582), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U4517 ( .A1(n4673), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U4518 ( .A1(n3773), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U4519 ( .A1(n3448), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4041) );
  NAND4_X1 U4520 ( .A1(n4044), .A2(n4043), .A3(n4042), .A4(n4041), .ZN(n4045)
         );
  NOR2_X1 U4521 ( .A1(n4046), .A2(n4045), .ZN(n4048) );
  AOI22_X1 U4522 ( .A1(n4691), .A2(EAX_REG_16__SCAN_IN), .B1(n3744), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4047) );
  OAI21_X1 U4523 ( .B1(n4178), .B2(n4048), .A(n4047), .ZN(n4049) );
  AOI21_X1 U4524 ( .B1(n6077), .B2(n3421), .A(n4049), .ZN(n5708) );
  OR2_X1 U4525 ( .A1(n4051), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4052)
         );
  NAND2_X1 U4526 ( .A1(n4052), .A2(n4102), .ZN(n6559) );
  AOI22_X1 U4527 ( .A1(n4673), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4267), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U4528 ( .A1(n4645), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U4529 ( .A1(n3773), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U4530 ( .A1(n4231), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4053) );
  NAND4_X1 U4531 ( .A1(n4056), .A2(n4055), .A3(n4054), .A4(n4053), .ZN(n4062)
         );
  AOI22_X1 U4532 ( .A1(n3424), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3582), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U4533 ( .A1(n3444), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U4534 ( .A1(n3719), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U4535 ( .A1(n3448), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4057) );
  NAND4_X1 U4536 ( .A1(n4060), .A2(n4059), .A3(n4058), .A4(n4057), .ZN(n4061)
         );
  NOR2_X1 U4537 ( .A1(n4062), .A2(n4061), .ZN(n4065) );
  INV_X1 U4538 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6930) );
  OAI21_X1 U4539 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6930), .A(n6906), 
        .ZN(n4064) );
  NAND2_X1 U4540 ( .A1(n4691), .A2(EAX_REG_18__SCAN_IN), .ZN(n4063) );
  OAI211_X1 U4541 ( .C1(n4178), .C2(n4065), .A(n4064), .B(n4063), .ZN(n4066)
         );
  OAI21_X1 U4542 ( .B1(n6559), .B2(n4685), .A(n4066), .ZN(n5903) );
  INV_X1 U4543 ( .A(n5903), .ZN(n4083) );
  XNOR2_X1 U4544 ( .A(n4067), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6817)
         );
  AOI22_X1 U4545 ( .A1(n4691), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6906), .ZN(n4082) );
  AOI22_X1 U4546 ( .A1(n4673), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4645), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U4547 ( .A1(n3424), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U4548 ( .A1(n4231), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U4549 ( .A1(n4666), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4068) );
  NAND4_X1 U4550 ( .A1(n4071), .A2(n4070), .A3(n4069), .A4(n4068), .ZN(n4080)
         );
  NAND2_X1 U4551 ( .A1(n3445), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4074)
         );
  NAND2_X1 U4552 ( .A1(n3779), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4073) );
  AND3_X1 U4553 ( .A1(n4074), .A2(n4685), .A3(n4073), .ZN(n4078) );
  AOI22_X1 U4554 ( .A1(n4267), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U4555 ( .A1(n3443), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U4556 ( .A1(n3425), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4075) );
  NAND4_X1 U4557 ( .A1(n4078), .A2(n4077), .A3(n4076), .A4(n4075), .ZN(n4079)
         );
  NAND2_X1 U4558 ( .A1(n4178), .A2(n4685), .ZN(n4133) );
  OAI21_X1 U4559 ( .B1(n4080), .B2(n4079), .A(n4133), .ZN(n4081) );
  AOI22_X1 U4560 ( .A1(n6817), .A2(n3421), .B1(n4082), .B2(n4081), .ZN(n5687)
         );
  NAND2_X1 U4561 ( .A1(n5686), .A2(n4084), .ZN(n5723) );
  AOI22_X1 U4562 ( .A1(n3442), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U4563 ( .A1(n4072), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3423), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U4564 ( .A1(n3612), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3577), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U4565 ( .A1(n4666), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4085) );
  NAND4_X1 U4566 ( .A1(n4088), .A2(n4087), .A3(n4086), .A4(n4085), .ZN(n4096)
         );
  NAND2_X1 U4567 ( .A1(n4231), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4090)
         );
  NAND2_X1 U4568 ( .A1(n4673), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4089) );
  AND3_X1 U4569 ( .A1(n4090), .A2(n4089), .A3(n4685), .ZN(n4094) );
  AOI22_X1 U4570 ( .A1(n3713), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4093) );
  AOI22_X1 U4571 ( .A1(n4650), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4092) );
  AOI22_X1 U4572 ( .A1(n4667), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4091) );
  NAND4_X1 U4573 ( .A1(n4094), .A2(n4093), .A3(n4092), .A4(n4091), .ZN(n4095)
         );
  OAI21_X1 U4574 ( .B1(n4096), .B2(n4095), .A(n4133), .ZN(n4098) );
  AOI22_X1 U4575 ( .A1(n4691), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6906), .ZN(n4097) );
  NAND2_X1 U4576 ( .A1(n4098), .A2(n4097), .ZN(n4100) );
  XNOR2_X1 U4577 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n4102), .ZN(n6054)
         );
  NAND2_X1 U4578 ( .A1(n3421), .A2(n6054), .ZN(n4099) );
  NAND2_X1 U4579 ( .A1(n4100), .A2(n4099), .ZN(n5724) );
  INV_X1 U4580 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4101) );
  INV_X1 U4581 ( .A(n4138), .ZN(n4105) );
  OR2_X1 U4582 ( .A1(n4103), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4104)
         );
  NAND2_X1 U4583 ( .A1(n4105), .A2(n4104), .ZN(n6834) );
  AOI22_X1 U4584 ( .A1(n3444), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4673), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U4585 ( .A1(n4231), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4666), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U4586 ( .A1(n4650), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U4587 ( .A1(n3448), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4106) );
  NAND4_X1 U4588 ( .A1(n4109), .A2(n4108), .A3(n4107), .A4(n4106), .ZN(n4115)
         );
  AOI22_X1 U4589 ( .A1(n4645), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3443), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U4590 ( .A1(n3612), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4112) );
  AOI22_X1 U4591 ( .A1(n3424), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4111) );
  AOI22_X1 U4592 ( .A1(n3577), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4110) );
  NAND4_X1 U4593 ( .A1(n4113), .A2(n4112), .A3(n4111), .A4(n4110), .ZN(n4114)
         );
  NOR2_X1 U4594 ( .A1(n4115), .A2(n4114), .ZN(n4119) );
  NAND2_X1 U4595 ( .A1(n6906), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4116)
         );
  NAND2_X1 U4596 ( .A1(n4685), .A2(n4116), .ZN(n4117) );
  AOI21_X1 U4597 ( .B1(n3870), .B2(EAX_REG_20__SCAN_IN), .A(n4117), .ZN(n4118)
         );
  OAI21_X1 U4598 ( .B1(n4178), .B2(n4119), .A(n4118), .ZN(n4120) );
  INV_X1 U4599 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4122) );
  XNOR2_X1 U4600 ( .A(n4138), .B(n4122), .ZN(n6835) );
  AOI22_X1 U4601 ( .A1(n4691), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6906), .ZN(n4137) );
  AOI22_X1 U4602 ( .A1(n4673), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4645), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U4603 ( .A1(n4650), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U4604 ( .A1(n3423), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U4605 ( .A1(n3445), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4123) );
  NAND4_X1 U4606 ( .A1(n4126), .A2(n4125), .A3(n4124), .A4(n4123), .ZN(n4135)
         );
  NAND2_X1 U4607 ( .A1(n4231), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4128)
         );
  NAND2_X1 U4608 ( .A1(n4268), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4127) );
  AND3_X1 U4609 ( .A1(n4128), .A2(n4127), .A3(n4685), .ZN(n4132) );
  AOI22_X1 U4610 ( .A1(n4267), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3577), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U4611 ( .A1(n3443), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U4612 ( .A1(n4666), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4129) );
  NAND4_X1 U4613 ( .A1(n4132), .A2(n4131), .A3(n4130), .A4(n4129), .ZN(n4134)
         );
  OAI21_X1 U4614 ( .B1(n4135), .B2(n4134), .A(n4133), .ZN(n4136) );
  AOI22_X1 U4615 ( .A1(n6835), .A2(n3421), .B1(n4137), .B2(n4136), .ZN(n5939)
         );
  INV_X1 U4616 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4151) );
  AND2_X1 U4617 ( .A1(n4139), .A2(n4151), .ZN(n4140) );
  OR2_X1 U4618 ( .A1(n4140), .A2(n4188), .ZN(n6040) );
  AOI22_X1 U4619 ( .A1(n4673), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4267), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4144) );
  AOI22_X1 U4620 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4666), .B1(n4231), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4143) );
  AOI22_X1 U4621 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(n4650), .B1(n4268), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4142) );
  AOI22_X1 U4622 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n4645), .B1(n3577), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4141) );
  NAND4_X1 U4623 ( .A1(n4144), .A2(n4143), .A3(n4142), .A4(n4141), .ZN(n4150)
         );
  AOI22_X1 U4624 ( .A1(n3444), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U4625 ( .A1(n3448), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4147) );
  AOI22_X1 U4626 ( .A1(n3425), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4146) );
  AOI22_X1 U4627 ( .A1(n3424), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4145) );
  NAND4_X1 U4628 ( .A1(n4148), .A2(n4147), .A3(n4146), .A4(n4145), .ZN(n4149)
         );
  NOR2_X1 U4629 ( .A1(n4150), .A2(n4149), .ZN(n4154) );
  OAI21_X1 U4630 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4151), .A(n4685), .ZN(
        n4152) );
  AOI21_X1 U4631 ( .B1(n3870), .B2(EAX_REG_22__SCAN_IN), .A(n4152), .ZN(n4153)
         );
  OAI21_X1 U4632 ( .B1(n4178), .B2(n4154), .A(n4153), .ZN(n4155) );
  OAI21_X1 U4633 ( .B1(n6040), .B2(n4685), .A(n4155), .ZN(n5894) );
  INV_X1 U4634 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4157) );
  XNOR2_X1 U4635 ( .A(n4188), .B(n4157), .ZN(n6843) );
  NAND2_X1 U4636 ( .A1(n6843), .A2(n3421), .ZN(n4185) );
  AOI22_X1 U4637 ( .A1(n4645), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4161) );
  AOI22_X1 U4638 ( .A1(n3443), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4160) );
  AOI22_X1 U4639 ( .A1(n4673), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U4640 ( .A1(n4666), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4158) );
  NAND4_X1 U4641 ( .A1(n4161), .A2(n4160), .A3(n4159), .A4(n4158), .ZN(n4167)
         );
  AOI22_X1 U4642 ( .A1(n3423), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4231), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4165) );
  AOI22_X1 U4643 ( .A1(n3445), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4267), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4164) );
  AOI22_X1 U4644 ( .A1(n3773), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4163) );
  AOI22_X1 U4645 ( .A1(n3425), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4162) );
  NAND4_X1 U4646 ( .A1(n4165), .A2(n4164), .A3(n4163), .A4(n4162), .ZN(n4166)
         );
  NOR2_X1 U4647 ( .A1(n4167), .A2(n4166), .ZN(n4189) );
  AOI22_X1 U4648 ( .A1(n4645), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4171) );
  AOI22_X1 U4649 ( .A1(n3445), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U4650 ( .A1(n4666), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U4651 ( .A1(n3773), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4168) );
  NAND4_X1 U4652 ( .A1(n4171), .A2(n4170), .A3(n4169), .A4(n4168), .ZN(n4177)
         );
  AOI22_X1 U4653 ( .A1(n4673), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4267), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4175) );
  AOI22_X1 U4654 ( .A1(n3424), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4231), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U4655 ( .A1(n3443), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4173) );
  AOI22_X1 U4656 ( .A1(n4667), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4172) );
  NAND4_X1 U4657 ( .A1(n4175), .A2(n4174), .A3(n4173), .A4(n4172), .ZN(n4176)
         );
  NOR2_X1 U4658 ( .A1(n4177), .A2(n4176), .ZN(n4190) );
  XOR2_X1 U4659 ( .A(n4189), .B(n4190), .Z(n4179) );
  NAND2_X1 U4660 ( .A1(n4179), .A2(n4682), .ZN(n4183) );
  NAND2_X1 U4661 ( .A1(n6906), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4180)
         );
  NAND2_X1 U4662 ( .A1(n4685), .A2(n4180), .ZN(n4181) );
  AOI21_X1 U4663 ( .B1(n3870), .B2(EAX_REG_23__SCAN_IN), .A(n4181), .ZN(n4182)
         );
  NAND2_X1 U4664 ( .A1(n4183), .A2(n4182), .ZN(n4184) );
  NAND2_X1 U4665 ( .A1(n4185), .A2(n4184), .ZN(n5930) );
  NAND2_X1 U4666 ( .A1(n4187), .A2(n4186), .ZN(n5929) );
  XNOR2_X1 U4667 ( .A(n4221), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6862)
         );
  OR2_X1 U4668 ( .A1(n4190), .A2(n4189), .ZN(n4218) );
  AOI22_X1 U4669 ( .A1(n3424), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4194) );
  AOI22_X1 U4670 ( .A1(n4072), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3713), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4193) );
  AOI22_X1 U4671 ( .A1(n4673), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4267), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4192) );
  AOI22_X1 U4672 ( .A1(n3773), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4191) );
  NAND4_X1 U4673 ( .A1(n4194), .A2(n4193), .A3(n4192), .A4(n4191), .ZN(n4200)
         );
  AOI22_X1 U4674 ( .A1(n4666), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4198) );
  AOI22_X1 U4675 ( .A1(n4231), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4197) );
  AOI22_X1 U4676 ( .A1(n3719), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4196) );
  AOI22_X1 U4677 ( .A1(n3425), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4195) );
  NAND4_X1 U4678 ( .A1(n4198), .A2(n4197), .A3(n4196), .A4(n4195), .ZN(n4199)
         );
  OR2_X1 U4679 ( .A1(n4200), .A2(n4199), .ZN(n4216) );
  XNOR2_X1 U4680 ( .A(n4218), .B(n4216), .ZN(n4203) );
  INV_X1 U4681 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4784) );
  INV_X1 U4682 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6024) );
  OAI22_X1 U4683 ( .A1(n3757), .A2(n4784), .B1(n4201), .B2(n6024), .ZN(n4202)
         );
  AOI21_X1 U4684 ( .B1(n4203), .B2(n4682), .A(n4202), .ZN(n4204) );
  AOI22_X1 U4685 ( .A1(n4072), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4209) );
  AOI22_X1 U4686 ( .A1(n4267), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3441), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4208) );
  AOI22_X1 U4687 ( .A1(n3425), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4668), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4207) );
  AOI22_X1 U4688 ( .A1(n4666), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4206) );
  NAND4_X1 U4689 ( .A1(n4209), .A2(n4208), .A3(n4207), .A4(n4206), .ZN(n4215)
         );
  AOI22_X1 U4690 ( .A1(n4673), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3713), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4213) );
  AOI22_X1 U4691 ( .A1(n3424), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4231), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4212) );
  AOI22_X1 U4692 ( .A1(n3443), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4211) );
  AOI22_X1 U4693 ( .A1(n3448), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4210) );
  NAND4_X1 U4694 ( .A1(n4213), .A2(n4212), .A3(n4211), .A4(n4210), .ZN(n4214)
         );
  NOR2_X1 U4695 ( .A1(n4215), .A2(n4214), .ZN(n4226) );
  INV_X1 U4696 ( .A(n4216), .ZN(n4217) );
  XOR2_X1 U4697 ( .A(n4226), .B(n4225), .Z(n4219) );
  NAND2_X1 U4698 ( .A1(n4219), .A2(n4682), .ZN(n4224) );
  INV_X1 U4699 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6005) );
  OAI21_X1 U4700 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6005), .A(n4685), .ZN(
        n4220) );
  AOI21_X1 U4701 ( .B1(n4691), .B2(EAX_REG_25__SCAN_IN), .A(n4220), .ZN(n4223)
         );
  XNOR2_X1 U4702 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .B(n4242), .ZN(n6007)
         );
  AOI21_X1 U4703 ( .B1(n4224), .B2(n4223), .A(n4222), .ZN(n5881) );
  NOR2_X1 U4704 ( .A1(n4226), .A2(n4225), .ZN(n4260) );
  AOI22_X1 U4705 ( .A1(n4673), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4267), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4230) );
  AOI22_X1 U4706 ( .A1(n3444), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4229) );
  AOI22_X1 U4707 ( .A1(n3713), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4228) );
  AOI22_X1 U4708 ( .A1(n3442), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3773), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4227) );
  NAND4_X1 U4709 ( .A1(n4230), .A2(n4229), .A3(n4228), .A4(n4227), .ZN(n4237)
         );
  AOI22_X1 U4710 ( .A1(n4231), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4666), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4235) );
  AOI22_X1 U4711 ( .A1(n3448), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4234) );
  AOI22_X1 U4712 ( .A1(n3425), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4233) );
  AOI22_X1 U4713 ( .A1(n3423), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4232) );
  NAND4_X1 U4714 ( .A1(n4235), .A2(n4234), .A3(n4233), .A4(n4232), .ZN(n4236)
         );
  OR2_X1 U4715 ( .A1(n4237), .A2(n4236), .ZN(n4259) );
  INV_X1 U4716 ( .A(n4259), .ZN(n4238) );
  XNOR2_X1 U4717 ( .A(n4260), .B(n4238), .ZN(n4241) );
  NAND2_X1 U4718 ( .A1(n6906), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4239)
         );
  OAI211_X1 U4719 ( .C1(n3757), .C2(n4863), .A(n4685), .B(n4239), .ZN(n4240)
         );
  AOI21_X1 U4720 ( .B1(n4241), .B2(n4682), .A(n4240), .ZN(n4248) );
  INV_X1 U4721 ( .A(n4244), .ZN(n4245) );
  INV_X1 U4722 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U4723 ( .A1(n4245), .A2(n5868), .ZN(n4246) );
  NAND2_X1 U4724 ( .A1(n4283), .A2(n4246), .ZN(n6000) );
  NOR2_X1 U4725 ( .A1(n6000), .A2(n4685), .ZN(n4247) );
  AOI22_X1 U4726 ( .A1(n4673), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3612), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4252) );
  AOI22_X1 U4727 ( .A1(n3445), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4251) );
  AOI22_X1 U4728 ( .A1(n3719), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3577), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4250) );
  AOI22_X1 U4729 ( .A1(n3423), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4249) );
  NAND4_X1 U4730 ( .A1(n4252), .A2(n4251), .A3(n4250), .A4(n4249), .ZN(n4258)
         );
  AOI22_X1 U4731 ( .A1(n4666), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4231), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4256) );
  AOI22_X1 U4732 ( .A1(n4645), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3441), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4255) );
  AOI22_X1 U4733 ( .A1(n3448), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4254) );
  AOI22_X1 U4734 ( .A1(n3425), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4253) );
  NAND4_X1 U4735 ( .A1(n4256), .A2(n4255), .A3(n4254), .A4(n4253), .ZN(n4257)
         );
  NOR2_X1 U4736 ( .A1(n4258), .A2(n4257), .ZN(n4280) );
  NAND2_X1 U4737 ( .A1(n4260), .A2(n4259), .ZN(n4279) );
  XOR2_X1 U4738 ( .A(n4280), .B(n4279), .Z(n4261) );
  NAND2_X1 U4739 ( .A1(n4261), .A2(n4682), .ZN(n4264) );
  INV_X1 U4740 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5989) );
  AOI21_X1 U4741 ( .B1(n5989), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4262) );
  AOI21_X1 U4742 ( .B1(n4691), .B2(EAX_REG_27__SCAN_IN), .A(n4262), .ZN(n4263)
         );
  NAND2_X1 U4743 ( .A1(n4264), .A2(n4263), .ZN(n4266) );
  XNOR2_X1 U4744 ( .A(n4283), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5992)
         );
  NAND2_X1 U4745 ( .A1(n5992), .A2(n3421), .ZN(n4265) );
  NAND2_X1 U4746 ( .A1(n4266), .A2(n4265), .ZN(n5855) );
  AOI22_X1 U4747 ( .A1(n4673), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4267), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4272) );
  AOI22_X1 U4748 ( .A1(n3444), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4268), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4271) );
  AOI22_X1 U4749 ( .A1(n3713), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4270) );
  AOI22_X1 U4750 ( .A1(n3443), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3577), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4269) );
  NAND4_X1 U4751 ( .A1(n4272), .A2(n4271), .A3(n4270), .A4(n4269), .ZN(n4278)
         );
  AOI22_X1 U4752 ( .A1(n4231), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3582), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4276) );
  AOI22_X1 U4753 ( .A1(n3448), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3603), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4275) );
  AOI22_X1 U4754 ( .A1(n3425), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4274) );
  AOI22_X1 U4755 ( .A1(n3424), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4273) );
  NAND4_X1 U4756 ( .A1(n4276), .A2(n4275), .A3(n4274), .A4(n4273), .ZN(n4277)
         );
  OR2_X1 U4757 ( .A1(n4278), .A2(n4277), .ZN(n4657) );
  NOR2_X1 U4758 ( .A1(n4280), .A2(n4279), .ZN(n4658) );
  XOR2_X1 U4759 ( .A(n4657), .B(n4658), .Z(n4281) );
  NAND2_X1 U4760 ( .A1(n4281), .A2(n4682), .ZN(n4288) );
  INV_X1 U4761 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5847) );
  NOR2_X1 U4762 ( .A1(n5847), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4282) );
  AOI211_X1 U4763 ( .C1(n4691), .C2(EAX_REG_28__SCAN_IN), .A(n3421), .B(n4282), 
        .ZN(n4287) );
  NAND2_X1 U4764 ( .A1(n4284), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4687)
         );
  INV_X1 U4765 ( .A(n4284), .ZN(n4285) );
  NAND2_X1 U4766 ( .A1(n4285), .A2(n5847), .ZN(n4286) );
  AND2_X1 U4767 ( .A1(n4687), .A2(n4286), .ZN(n5846) );
  AOI22_X1 U4768 ( .A1(n4288), .A2(n4287), .B1(n3421), .B2(n5846), .ZN(n4290)
         );
  INV_X1 U4769 ( .A(n4663), .ZN(n4292) );
  INV_X1 U4770 ( .A(n4289), .ZN(n5857) );
  INV_X1 U4771 ( .A(n4290), .ZN(n4291) );
  MUX2_X1 U4772 ( .A(n5172), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n4299) );
  NAND2_X1 U4773 ( .A1(n7025), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4303) );
  NAND2_X1 U4774 ( .A1(n4299), .A2(n4298), .ZN(n4294) );
  NAND2_X1 U4775 ( .A1(n5172), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4293) );
  NAND2_X1 U4776 ( .A1(n4294), .A2(n4293), .ZN(n4316) );
  XNOR2_X1 U4777 ( .A(n5774), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4315)
         );
  NAND2_X1 U4778 ( .A1(n4316), .A2(n4315), .ZN(n4296) );
  NAND2_X1 U4779 ( .A1(n6883), .A2(n5774), .ZN(n4295) );
  NAND2_X1 U4780 ( .A1(n4296), .A2(n4295), .ZN(n4328) );
  MUX2_X1 U4781 ( .A(n6889), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n4327) );
  XNOR2_X1 U4782 ( .A(n4328), .B(n4327), .ZN(n4566) );
  NAND2_X1 U4783 ( .A1(n4297), .A2(n4566), .ZN(n4325) );
  XNOR2_X1 U4784 ( .A(n4299), .B(n4298), .ZN(n4565) );
  NOR2_X1 U4785 ( .A1(n4565), .A2(n6923), .ZN(n4300) );
  NOR2_X1 U4786 ( .A1(n4343), .A2(n4300), .ZN(n4309) );
  INV_X1 U4787 ( .A(n4309), .ZN(n4314) );
  NAND2_X1 U4788 ( .A1(n4329), .A2(n4565), .ZN(n4302) );
  NAND2_X1 U4789 ( .A1(n4340), .A2(n3659), .ZN(n4301) );
  AND3_X1 U4790 ( .A1(n4302), .A2(n4455), .A3(n4301), .ZN(n4310) );
  INV_X1 U4791 ( .A(n4310), .ZN(n4313) );
  OAI21_X1 U4792 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7025), .A(n4303), 
        .ZN(n4305) );
  INV_X1 U4793 ( .A(n4305), .ZN(n4304) );
  NAND2_X1 U4794 ( .A1(n4340), .A2(n4304), .ZN(n4311) );
  INV_X1 U4795 ( .A(n4343), .ZN(n4330) );
  INV_X1 U4796 ( .A(n3660), .ZN(n4306) );
  OAI21_X1 U4797 ( .B1(n4306), .B2(n4305), .A(n3643), .ZN(n4308) );
  NAND2_X1 U4798 ( .A1(n4913), .A2(n4455), .ZN(n4307) );
  AOI222_X1 U4799 ( .A1(n4311), .A2(n4330), .B1(n4310), .B2(n4309), .C1(n4308), 
        .C2(n4321), .ZN(n4312) );
  AOI21_X1 U4800 ( .B1(n4314), .B2(n4313), .A(n4312), .ZN(n4323) );
  XNOR2_X1 U4801 ( .A(n4316), .B(n4315), .ZN(n4564) );
  INV_X1 U4802 ( .A(n4321), .ZN(n4318) );
  INV_X1 U4803 ( .A(n4340), .ZN(n4317) );
  AOI211_X1 U4804 ( .C1(n4329), .C2(n4564), .A(n4318), .B(n4319), .ZN(n4322)
         );
  INV_X1 U4805 ( .A(n4319), .ZN(n4320) );
  OAI22_X1 U4806 ( .A1(n4323), .A2(n4322), .B1(n4321), .B2(n4320), .ZN(n4324)
         );
  AOI22_X1 U4807 ( .A1(n4325), .A2(n4324), .B1(n4343), .B2(n4566), .ZN(n4332)
         );
  NOR2_X1 U4808 ( .A1(n4950), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4326)
         );
  NAND2_X1 U4809 ( .A1(n4335), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4334) );
  NOR2_X1 U4810 ( .A1(n4329), .A2(n4569), .ZN(n4331) );
  NAND2_X1 U4811 ( .A1(n4334), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4339) );
  INV_X1 U4812 ( .A(n4335), .ZN(n4337) );
  INV_X1 U4813 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4336) );
  NAND2_X1 U4814 ( .A1(n4337), .A2(n4336), .ZN(n4338) );
  NAND2_X1 U4815 ( .A1(n4339), .A2(n4338), .ZN(n4568) );
  NAND2_X1 U4816 ( .A1(n4340), .A2(n4568), .ZN(n4341) );
  NAND2_X1 U4817 ( .A1(n4343), .A2(n4568), .ZN(n4344) );
  NAND2_X1 U4818 ( .A1(n4905), .A2(n3658), .ZN(n4366) );
  INV_X1 U4819 ( .A(n5790), .ZN(n4349) );
  OAI21_X1 U4820 ( .B1(n4357), .B2(n3643), .A(n3676), .ZN(n4348) );
  AND2_X1 U4821 ( .A1(n4886), .A2(n3659), .ZN(n5826) );
  NAND2_X1 U4822 ( .A1(n5826), .A2(n3446), .ZN(n4347) );
  OAI211_X1 U4823 ( .C1(n4556), .C2(n4349), .A(n4348), .B(n4347), .ZN(n4353)
         );
  AND2_X1 U4824 ( .A1(n4350), .A2(n3643), .ZN(n4352) );
  MUX2_X1 U4825 ( .A(n4352), .B(n6581), .S(n4351), .Z(n4563) );
  NOR2_X1 U4826 ( .A1(n4353), .A2(n4563), .ZN(n4603) );
  AND3_X1 U4827 ( .A1(n4354), .A2(n4355), .A3(n4874), .ZN(n4356) );
  AND2_X1 U4828 ( .A1(n4357), .A2(n3643), .ZN(n4580) );
  NAND2_X1 U4829 ( .A1(n4358), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6928) );
  NAND4_X1 U4830 ( .A1(n5160), .A2(n5812), .A3(n5829), .A4(n3634), .ZN(n4873)
         );
  NOR3_X1 U4831 ( .A1(n4360), .A2(n4873), .A3(n4359), .ZN(n4361) );
  MUX2_X1 U4832 ( .A(n4374), .B(n4366), .S(EBX_REG_1__SCAN_IN), .Z(n4365) );
  INV_X1 U4833 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4363) );
  NAND2_X1 U4834 ( .A1(n4365), .A2(n4364), .ZN(n4370) );
  INV_X1 U4835 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4849) );
  NAND2_X1 U4836 ( .A1(n4374), .A2(n4849), .ZN(n4367) );
  NAND2_X1 U4837 ( .A1(n4368), .A2(n4367), .ZN(n4848) );
  XNOR2_X1 U4838 ( .A(n4370), .B(n4848), .ZN(n5368) );
  INV_X1 U4839 ( .A(n4848), .ZN(n4369) );
  NOR2_X1 U4840 ( .A1(n4370), .A2(n4369), .ZN(n4371) );
  AOI21_X1 U4841 ( .B1(n5368), .B2(n4850), .A(n4371), .ZN(n4836) );
  NAND2_X1 U4842 ( .A1(n4359), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4372)
         );
  NAND2_X1 U4843 ( .A1(n4373), .A2(n4372), .ZN(n4835) );
  NAND2_X1 U4844 ( .A1(n4836), .A2(n4835), .ZN(n4834) );
  MUX2_X1 U4845 ( .A(n4440), .B(n4374), .S(EBX_REG_3__SCAN_IN), .Z(n4376) );
  NAND2_X1 U4846 ( .A1(n4376), .A2(n4375), .ZN(n4827) );
  MUX2_X1 U4847 ( .A(n4374), .B(n4444), .S(EBX_REG_4__SCAN_IN), .Z(n4378) );
  NAND2_X1 U4848 ( .A1(n4359), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4377)
         );
  OR2_X1 U4849 ( .A1(n4440), .A2(EBX_REG_5__SCAN_IN), .ZN(n4381) );
  NAND2_X1 U4850 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4379)
         );
  INV_X1 U4851 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6638) );
  NAND2_X1 U4852 ( .A1(n4444), .A2(n6638), .ZN(n4382) );
  OAI211_X1 U4853 ( .C1(n4359), .C2(EBX_REG_6__SCAN_IN), .A(n4382), .B(n4374), 
        .ZN(n4385) );
  INV_X1 U4854 ( .A(n4383), .ZN(n4595) );
  INV_X1 U4855 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6762) );
  NAND2_X1 U4856 ( .A1(n4595), .A2(n6762), .ZN(n4384) );
  NAND2_X1 U4857 ( .A1(n4385), .A2(n4384), .ZN(n5048) );
  OR2_X1 U4858 ( .A1(n4440), .A2(EBX_REG_7__SCAN_IN), .ZN(n4388) );
  NAND2_X1 U4859 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4386)
         );
  OAI211_X1 U4860 ( .C1(n4359), .C2(EBX_REG_7__SCAN_IN), .A(n4444), .B(n4386), 
        .ZN(n4387) );
  NAND2_X1 U4861 ( .A1(n4388), .A2(n4387), .ZN(n6492) );
  NAND2_X1 U4862 ( .A1(n4359), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4389)
         );
  OR2_X1 U4863 ( .A1(n4440), .A2(EBX_REG_9__SCAN_IN), .ZN(n4393) );
  NAND2_X1 U4864 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4391)
         );
  OAI211_X1 U4865 ( .C1(n4359), .C2(EBX_REG_9__SCAN_IN), .A(n4444), .B(n4391), 
        .ZN(n4392) );
  MUX2_X1 U4866 ( .A(n4440), .B(n4374), .S(EBX_REG_11__SCAN_IN), .Z(n4395) );
  OR2_X1 U4867 ( .A1(n5790), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4394)
         );
  NAND2_X1 U4868 ( .A1(n4395), .A2(n4394), .ZN(n5498) );
  NAND2_X1 U4869 ( .A1(n4359), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4396) );
  NAND2_X1 U4870 ( .A1(n4397), .A2(n4396), .ZN(n5496) );
  INV_X1 U4871 ( .A(n5496), .ZN(n4398) );
  NOR2_X1 U4872 ( .A1(n5498), .A2(n4398), .ZN(n4399) );
  INV_X1 U4873 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U4874 ( .A1(n4444), .A2(n5618), .ZN(n4400) );
  OAI211_X1 U4875 ( .C1(n4359), .C2(EBX_REG_12__SCAN_IN), .A(n4400), .B(n4374), 
        .ZN(n4402) );
  INV_X1 U4876 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U4877 ( .A1(n4595), .A2(n5598), .ZN(n4401) );
  MUX2_X1 U4878 ( .A(n4440), .B(n4374), .S(EBX_REG_13__SCAN_IN), .Z(n4404) );
  OR2_X1 U4879 ( .A1(n5790), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4403)
         );
  NAND2_X1 U4880 ( .A1(n4404), .A2(n4403), .ZN(n5644) );
  OR2_X2 U4881 ( .A1(n5645), .A2(n5644), .ZN(n5647) );
  MUX2_X1 U4882 ( .A(n4374), .B(n4444), .S(EBX_REG_14__SCAN_IN), .Z(n4406) );
  NAND2_X1 U4883 ( .A1(n4359), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4405) );
  NAND2_X1 U4884 ( .A1(n4406), .A2(n4405), .ZN(n5641) );
  INV_X1 U4885 ( .A(n5641), .ZN(n4407) );
  NOR2_X2 U4886 ( .A1(n5647), .A2(n4407), .ZN(n5678) );
  OR2_X1 U4887 ( .A1(n4440), .A2(EBX_REG_15__SCAN_IN), .ZN(n4410) );
  NAND2_X1 U4888 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4408) );
  NAND2_X1 U4889 ( .A1(n5678), .A2(n5677), .ZN(n5711) );
  NAND2_X1 U4890 ( .A1(n4359), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4411) );
  AND2_X1 U4891 ( .A1(n4412), .A2(n4411), .ZN(n5710) );
  OR2_X1 U4892 ( .A1(n4440), .A2(EBX_REG_17__SCAN_IN), .ZN(n4415) );
  NAND2_X1 U4893 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4413) );
  OAI211_X1 U4894 ( .C1(n4359), .C2(EBX_REG_17__SCAN_IN), .A(n4444), .B(n4413), 
        .ZN(n4414) );
  NAND2_X1 U4895 ( .A1(n4415), .A2(n4414), .ZN(n5688) );
  MUX2_X1 U4896 ( .A(n4374), .B(n4444), .S(EBX_REG_18__SCAN_IN), .Z(n4417) );
  NAND2_X1 U4897 ( .A1(n4359), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4416) );
  NAND2_X1 U4898 ( .A1(n4417), .A2(n4416), .ZN(n5907) );
  OR2_X1 U4899 ( .A1(n4440), .A2(EBX_REG_19__SCAN_IN), .ZN(n4420) );
  NAND2_X1 U4900 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4418) );
  AND2_X1 U4901 ( .A1(n4420), .A2(n4419), .ZN(n5726) );
  INV_X1 U4902 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U4903 ( .A1(n4444), .A2(n6018), .ZN(n4421) );
  OAI211_X1 U4904 ( .C1(n4359), .C2(EBX_REG_20__SCAN_IN), .A(n4421), .B(n4374), 
        .ZN(n4423) );
  INV_X1 U4905 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U4906 ( .A1(n4595), .A2(n5953), .ZN(n4422) );
  AND2_X1 U4907 ( .A1(n4423), .A2(n4422), .ZN(n5949) );
  OR2_X1 U4908 ( .A1(n4440), .A2(EBX_REG_21__SCAN_IN), .ZN(n4426) );
  NAND2_X1 U4909 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4424) );
  OAI211_X1 U4910 ( .C1(n4359), .C2(EBX_REG_21__SCAN_IN), .A(n4444), .B(n4424), 
        .ZN(n4425) );
  NAND2_X1 U4911 ( .A1(n4426), .A2(n4425), .ZN(n5941) );
  NAND2_X1 U4912 ( .A1(n4359), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4427) );
  NAND2_X1 U4913 ( .A1(n4428), .A2(n4427), .ZN(n5896) );
  INV_X1 U4914 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5935) );
  MUX2_X1 U4915 ( .A(n4374), .B(n4440), .S(n5935), .Z(n4430) );
  OR2_X1 U4916 ( .A1(n5790), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4429)
         );
  NAND2_X1 U4917 ( .A1(n4430), .A2(n4429), .ZN(n5932) );
  MUX2_X1 U4918 ( .A(n4440), .B(n4374), .S(EBX_REG_25__SCAN_IN), .Z(n4432) );
  OR2_X1 U4919 ( .A1(n5790), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4431)
         );
  AND2_X1 U4920 ( .A1(n4432), .A2(n4431), .ZN(n5884) );
  INV_X1 U4921 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U4922 ( .A1(n4444), .A2(n6117), .ZN(n4434) );
  OR2_X1 U4923 ( .A1(n4359), .A2(EBX_REG_24__SCAN_IN), .ZN(n4433) );
  NAND3_X1 U4924 ( .A1(n4434), .A2(n4374), .A3(n4433), .ZN(n4436) );
  INV_X1 U4925 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6502) );
  NAND2_X1 U4926 ( .A1(n4595), .A2(n6502), .ZN(n4435) );
  NAND2_X1 U4927 ( .A1(n4436), .A2(n4435), .ZN(n6111) );
  NAND2_X1 U4928 ( .A1(n4359), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4437) );
  NAND2_X1 U4929 ( .A1(n4438), .A2(n4437), .ZN(n5871) );
  INV_X1 U4930 ( .A(n5871), .ZN(n4439) );
  OR2_X1 U4931 ( .A1(n4440), .A2(EBX_REG_27__SCAN_IN), .ZN(n4443) );
  NAND2_X1 U4932 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4441) );
  AND2_X1 U4933 ( .A1(n4443), .A2(n4442), .ZN(n4628) );
  MUX2_X1 U4934 ( .A(n4374), .B(n4444), .S(EBX_REG_28__SCAN_IN), .Z(n4446) );
  NAND2_X1 U4935 ( .A1(n4359), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4445) );
  NAND2_X1 U4936 ( .A1(n4446), .A2(n4445), .ZN(n4447) );
  NOR2_X1 U4937 ( .A1(n4630), .A2(n4447), .ZN(n4448) );
  INV_X1 U4938 ( .A(EBX_REG_28__SCAN_IN), .ZN(n4449) );
  INV_X1 U4939 ( .A(n6581), .ZN(n4593) );
  AND2_X1 U4940 ( .A1(n4462), .A2(n4454), .ZN(n4469) );
  NOR2_X1 U4941 ( .A1(n4593), .A2(n4469), .ZN(n4471) );
  INV_X1 U4942 ( .A(n4471), .ZN(n4457) );
  NOR2_X1 U4943 ( .A1(n4462), .A2(n4454), .ZN(n4456) );
  OAI211_X1 U4944 ( .C1(n4457), .C2(n4456), .A(n4908), .B(n4455), .ZN(n4458)
         );
  INV_X1 U4945 ( .A(n4574), .ZN(n4519) );
  AND2_X1 U4946 ( .A1(n4886), .A2(n4460), .ZN(n4472) );
  INV_X1 U4947 ( .A(n4472), .ZN(n4461) );
  OAI21_X1 U4948 ( .B1(n4593), .B2(n4462), .A(n4461), .ZN(n4463) );
  INV_X1 U4949 ( .A(n4463), .ZN(n4464) );
  OAI21_X1 U4950 ( .B1(n5746), .B2(n4519), .A(n4464), .ZN(n4811) );
  NAND2_X1 U4951 ( .A1(n4810), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4465)
         );
  NAND2_X1 U4952 ( .A1(n5523), .A2(n4465), .ZN(n4468) );
  INV_X1 U4953 ( .A(n4810), .ZN(n4466) );
  NAND2_X1 U4954 ( .A1(n4466), .A2(n4363), .ZN(n4467) );
  INV_X1 U4955 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6661) );
  INV_X1 U4956 ( .A(n4469), .ZN(n4478) );
  NOR2_X1 U4957 ( .A1(n4593), .A2(n4478), .ZN(n4470) );
  MUX2_X1 U4958 ( .A(n4471), .B(n4470), .S(n4476), .Z(n4473) );
  AOI21_X2 U4959 ( .B1(n4888), .B2(n4574), .A(n3456), .ZN(n6512) );
  NAND2_X1 U4960 ( .A1(n6511), .A2(n6661), .ZN(n4474) );
  NAND2_X1 U4961 ( .A1(n4475), .A2(n4474), .ZN(n4483) );
  INV_X1 U4962 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6620) );
  NAND2_X1 U4963 ( .A1(n4483), .A2(n6620), .ZN(n4820) );
  INV_X1 U4964 ( .A(n4476), .ZN(n4477) );
  NAND2_X1 U4965 ( .A1(n4478), .A2(n4477), .ZN(n4479) );
  NAND2_X1 U4966 ( .A1(n4479), .A2(n4480), .ZN(n4495) );
  OAI211_X1 U4967 ( .C1(n4480), .C2(n4479), .A(n4495), .B(n6581), .ZN(n4481)
         );
  NAND2_X1 U4968 ( .A1(n4820), .A2(n4823), .ZN(n4485) );
  INV_X1 U4969 ( .A(n4483), .ZN(n4484) );
  NAND2_X1 U4970 ( .A1(n4484), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4821)
         );
  NAND2_X1 U4971 ( .A1(n4486), .A2(n4574), .ZN(n4489) );
  XNOR2_X1 U4972 ( .A(n4495), .B(n4493), .ZN(n4487) );
  NAND2_X1 U4973 ( .A1(n4487), .A2(n6581), .ZN(n4488) );
  INV_X1 U4974 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6627) );
  NAND2_X1 U4975 ( .A1(n6520), .A2(n6519), .ZN(n6518) );
  NAND2_X1 U4976 ( .A1(n4490), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4491)
         );
  INV_X1 U4977 ( .A(n4493), .ZN(n4494) );
  OR2_X1 U4978 ( .A1(n4495), .A2(n4494), .ZN(n4502) );
  XNOR2_X1 U4979 ( .A(n4502), .B(n4503), .ZN(n4496) );
  NAND2_X1 U4980 ( .A1(n4496), .A2(n6581), .ZN(n4497) );
  INV_X1 U4981 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6633) );
  XNOR2_X1 U4982 ( .A(n4498), .B(n6633), .ZN(n6525) );
  NAND2_X1 U4983 ( .A1(n4498), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4499)
         );
  NAND3_X1 U4984 ( .A1(n4500), .A2(n4574), .A3(n4501), .ZN(n4507) );
  INV_X1 U4985 ( .A(n4502), .ZN(n4504) );
  NAND2_X1 U4986 ( .A1(n4504), .A2(n4503), .ZN(n4511) );
  XNOR2_X1 U4987 ( .A(n4511), .B(n4512), .ZN(n4505) );
  NAND2_X1 U4988 ( .A1(n4505), .A2(n6581), .ZN(n4506) );
  NAND2_X1 U4989 ( .A1(n4507), .A2(n4506), .ZN(n4508) );
  XNOR2_X1 U4990 ( .A(n4508), .B(n6638), .ZN(n6532) );
  NAND2_X1 U4991 ( .A1(n4508), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4509)
         );
  INV_X1 U4992 ( .A(n4510), .ZN(n4516) );
  INV_X1 U4993 ( .A(n4511), .ZN(n4513) );
  NAND2_X1 U4994 ( .A1(n4513), .A2(n4512), .ZN(n4522) );
  XNOR2_X1 U4995 ( .A(n4523), .B(n4522), .ZN(n4514) );
  NAND2_X1 U4996 ( .A1(n4514), .A2(n6581), .ZN(n4515) );
  INV_X1 U4997 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6667) );
  XNOR2_X1 U4998 ( .A(n4517), .B(n6667), .ZN(n6539) );
  NAND2_X1 U4999 ( .A1(n4517), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4518)
         );
  NOR3_X1 U5000 ( .A1(n4520), .A2(n4519), .A3(n6923), .ZN(n4521) );
  INV_X1 U5001 ( .A(n4522), .ZN(n4524) );
  NAND3_X1 U5002 ( .A1(n4524), .A2(n6581), .A3(n4523), .ZN(n4525) );
  NAND2_X1 U5003 ( .A1(n4540), .A2(n4525), .ZN(n4526) );
  INV_X1 U5004 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5337) );
  XNOR2_X1 U5005 ( .A(n4526), .B(n5337), .ZN(n5332) );
  NAND2_X1 U5006 ( .A1(n5333), .A2(n5332), .ZN(n5331) );
  NAND2_X1 U5007 ( .A1(n4526), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4527)
         );
  XNOR2_X1 U5008 ( .A(n3449), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5591)
         );
  NAND2_X1 U5009 ( .A1(n5592), .A2(n5591), .ZN(n5590) );
  INV_X1 U5010 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6669) );
  OR2_X1 U5011 ( .A1(n3449), .A2(n6669), .ZN(n4528) );
  AND2_X1 U5012 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4530) );
  INV_X1 U5013 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5609) );
  OR2_X1 U5014 ( .A1(n4540), .A2(n5609), .ZN(n5610) );
  OAI21_X1 U5015 ( .B1(n5618), .B2(n4540), .A(n5610), .ZN(n4529) );
  INV_X1 U5016 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4531) );
  NAND2_X1 U5017 ( .A1(n4540), .A2(n4531), .ZN(n4532) );
  INV_X1 U5018 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5635) );
  AND2_X1 U5019 ( .A1(n3449), .A2(n5635), .ZN(n4535) );
  INV_X1 U5020 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6700) );
  NAND2_X1 U5021 ( .A1(n4540), .A2(n6700), .ZN(n5696) );
  INV_X1 U5022 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6707) );
  NOR2_X1 U5023 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4537) );
  NAND2_X1 U5024 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4609) );
  NAND2_X1 U5025 ( .A1(n3449), .A2(n4609), .ZN(n4538) );
  NOR2_X1 U5026 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6132) );
  NOR2_X1 U5027 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6156) );
  NOR2_X1 U5028 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4539) );
  INV_X1 U5029 ( .A(n6014), .ZN(n6029) );
  AND2_X1 U5030 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U5031 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U5032 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4613) );
  NOR2_X1 U5033 ( .A1(n6123), .A2(n4613), .ZN(n4620) );
  XNOR2_X1 U5034 ( .A(n4540), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6010)
         );
  INV_X1 U5035 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U5036 ( .A1(n4540), .A2(n6095), .ZN(n4543) );
  INV_X1 U5037 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6096) );
  AND2_X1 U5038 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5751) );
  NAND2_X1 U5039 ( .A1(n5751), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5786) );
  NAND2_X1 U5040 ( .A1(n4540), .A2(n5786), .ZN(n4545) );
  NAND2_X1 U5041 ( .A1(n4640), .A2(n4545), .ZN(n4548) );
  NOR2_X1 U5042 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4546) );
  OR2_X1 U5043 ( .A1(n4540), .A2(n4546), .ZN(n5978) );
  INV_X1 U5044 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6082) );
  OR2_X1 U5045 ( .A1(n4540), .A2(n6082), .ZN(n4547) );
  NAND2_X1 U5046 ( .A1(n4548), .A2(n5747), .ZN(n4639) );
  NAND2_X1 U5047 ( .A1(n6019), .A2(n4638), .ZN(n4549) );
  OR2_X2 U5048 ( .A1(n4639), .A2(n4549), .ZN(n4551) );
  NAND2_X1 U5049 ( .A1(n4639), .A2(n3449), .ZN(n4550) );
  NAND2_X1 U5050 ( .A1(n4551), .A2(n4550), .ZN(n4552) );
  XNOR2_X1 U5051 ( .A(n4552), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5772)
         );
  OR2_X1 U5052 ( .A1(n6942), .A2(STATE_REG_0__SCAN_IN), .ZN(n6575) );
  INV_X1 U5053 ( .A(n6575), .ZN(n5827) );
  OR2_X1 U5054 ( .A1(n3659), .A2(n5827), .ZN(n5363) );
  INV_X1 U5055 ( .A(READY_N), .ZN(n6943) );
  AND2_X1 U5056 ( .A1(n5363), .A2(n6943), .ZN(n4553) );
  NAND2_X1 U5057 ( .A1(n5817), .A2(n4553), .ZN(n4753) );
  NAND2_X1 U5058 ( .A1(n3654), .A2(n3746), .ZN(n4554) );
  OR2_X1 U5059 ( .A1(n3653), .A2(n4554), .ZN(n4597) );
  NAND2_X1 U5060 ( .A1(n4597), .A2(n4886), .ZN(n4555) );
  NAND2_X1 U5061 ( .A1(n4556), .A2(n4555), .ZN(n4585) );
  INV_X1 U5062 ( .A(n4557), .ZN(n4559) );
  NOR2_X1 U5063 ( .A1(n4559), .A2(n4558), .ZN(n4560) );
  AND2_X1 U5064 ( .A1(n4561), .A2(n4560), .ZN(n5821) );
  INV_X1 U5065 ( .A(n5821), .ZN(n4562) );
  OAI21_X1 U5066 ( .B1(n4563), .B2(n4585), .A(n4562), .ZN(n4755) );
  NAND2_X1 U5067 ( .A1(n3659), .A2(n6575), .ZN(n4572) );
  NOR3_X1 U5068 ( .A1(n4566), .A2(n4565), .A3(n4564), .ZN(n4567) );
  OR2_X1 U5069 ( .A1(n4568), .A2(n4567), .ZN(n4570) );
  NAND2_X1 U5070 ( .A1(n4570), .A2(n4569), .ZN(n5816) );
  NAND2_X1 U5071 ( .A1(n6943), .A2(n5816), .ZN(n4872) );
  INV_X1 U5072 ( .A(n4872), .ZN(n4571) );
  NAND3_X1 U5073 ( .A1(n4572), .A2(n3676), .A3(n4571), .ZN(n4573) );
  AND2_X1 U5074 ( .A1(n4755), .A2(n4573), .ZN(n4578) );
  NAND2_X1 U5075 ( .A1(n4575), .A2(n4574), .ZN(n4576) );
  OR2_X1 U5076 ( .A1(n5817), .A2(n4576), .ZN(n4577) );
  OAI211_X1 U5077 ( .C1(n4753), .C2(n4354), .A(n4578), .B(n4577), .ZN(n4579)
         );
  NAND2_X1 U5078 ( .A1(n4579), .A2(n5829), .ZN(n4582) );
  INV_X1 U5079 ( .A(n4584), .ZN(n4586) );
  OR2_X1 U5080 ( .A1(n4585), .A2(n3673), .ZN(n4879) );
  OR2_X1 U5081 ( .A1(n4585), .A2(n3660), .ZN(n6891) );
  AND2_X1 U5082 ( .A1(n4879), .A2(n6891), .ZN(n5819) );
  OAI211_X1 U5083 ( .C1(n5160), .C2(n4583), .A(n4586), .B(n5819), .ZN(n4587)
         );
  INV_X1 U5084 ( .A(n4590), .ZN(n5756) );
  OAI22_X1 U5085 ( .A1(n5790), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n4359), .ZN(n4591) );
  INV_X1 U5086 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4588) );
  NAND2_X1 U5087 ( .A1(n4595), .A2(n4588), .ZN(n4589) );
  OAI21_X1 U5088 ( .B1(n4591), .B2(n4595), .A(n4589), .ZN(n5754) );
  OAI21_X1 U5089 ( .B1(n5756), .B2(n4591), .A(n5791), .ZN(n4592) );
  OAI22_X1 U5090 ( .A1(n5790), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        EBX_REG_30__SCAN_IN), .B2(n4359), .ZN(n5792) );
  OR2_X1 U5091 ( .A1(n4354), .A2(n4593), .ZN(n6904) );
  OAI21_X1 U5092 ( .B1(n4583), .B2(n3654), .A(n6904), .ZN(n4594) );
  NAND2_X1 U5093 ( .A1(n5920), .A2(n6721), .ZN(n4625) );
  INV_X1 U5094 ( .A(n5786), .ZN(n4615) );
  INV_X1 U5095 ( .A(n3680), .ZN(n4600) );
  NAND2_X1 U5096 ( .A1(n4596), .A2(n4595), .ZN(n4599) );
  INV_X1 U5097 ( .A(n4597), .ZN(n4598) );
  NAND2_X1 U5098 ( .A1(n4598), .A2(n3446), .ZN(n4957) );
  OAI211_X1 U5099 ( .C1(n4874), .C2(n4600), .A(n4599), .B(n4957), .ZN(n4601)
         );
  INV_X1 U5100 ( .A(n4601), .ZN(n4602) );
  NAND3_X1 U5101 ( .A1(n4603), .A2(n4602), .A3(n4747), .ZN(n4604) );
  NAND2_X1 U5102 ( .A1(n4606), .A2(n4604), .ZN(n6594) );
  NAND2_X1 U5103 ( .A1(n6594), .A2(n6651), .ZN(n6725) );
  AND2_X1 U5104 ( .A1(n5821), .A2(n3659), .ZN(n4958) );
  NAND2_X1 U5105 ( .A1(n4606), .A2(n4958), .ZN(n4612) );
  INV_X1 U5106 ( .A(n4612), .ZN(n6727) );
  NAND2_X1 U5107 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4622) );
  NAND2_X1 U5108 ( .A1(n4612), .A2(n6594), .ZN(n6170) );
  NOR2_X1 U5109 ( .A1(n6170), .A2(n6612), .ZN(n4611) );
  NAND2_X1 U5110 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6598) );
  NOR2_X1 U5111 ( .A1(n4531), .A2(n6598), .ZN(n5640) );
  NAND2_X1 U5112 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5640), .ZN(n6695) );
  NOR3_X1 U5113 ( .A1(n6707), .A2(n6700), .A3(n6695), .ZN(n6167) );
  NAND2_X1 U5114 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6167), .ZN(n6154) );
  NAND2_X1 U5115 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6640) );
  NOR3_X1 U5116 ( .A1(n6638), .A2(n6633), .A3(n6640), .ZN(n5334) );
  NOR2_X1 U5117 ( .A1(n5337), .A2(n6667), .ZN(n6673) );
  NAND4_X1 U5118 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n5334), .A4(n6673), .ZN(n4608)
         );
  INV_X1 U5119 ( .A(n4608), .ZN(n4605) );
  INV_X1 U5120 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6611) );
  OAI21_X1 U5121 ( .B1(n4363), .B2(n6611), .A(n6661), .ZN(n6653) );
  NAND2_X1 U5122 ( .A1(n4605), .A2(n6653), .ZN(n4616) );
  NOR2_X1 U5123 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n7031) );
  NAND2_X1 U5124 ( .A1(n7031), .A2(n5348), .ZN(n6571) );
  INV_X2 U5125 ( .A(n6821), .ZN(n6789) );
  OAI22_X1 U5126 ( .A1(n6594), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(n6789), 
        .B2(n4606), .ZN(n6610) );
  AOI21_X1 U5127 ( .B1(n6612), .B2(n4616), .A(n6610), .ZN(n5619) );
  INV_X1 U5128 ( .A(n5619), .ZN(n4607) );
  AOI21_X1 U5129 ( .B1(n6612), .B2(n6154), .A(n4607), .ZN(n6168) );
  NAND2_X1 U5130 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6649) );
  NOR2_X1 U5131 ( .A1(n4608), .A2(n6649), .ZN(n6597) );
  NAND2_X1 U5132 ( .A1(n6167), .A2(n6597), .ZN(n6171) );
  NOR2_X1 U5133 ( .A1(n6171), .A2(n4609), .ZN(n6151) );
  INV_X1 U5134 ( .A(n6151), .ZN(n4618) );
  INV_X1 U5135 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6165) );
  AOI22_X1 U5136 ( .A1(n6170), .A2(n4618), .B1(n6612), .B2(n6165), .ZN(n4610)
         );
  OAI211_X1 U5137 ( .C1(n6155), .C2(n4611), .A(n6168), .B(n4610), .ZN(n6142)
         );
  AOI21_X1 U5138 ( .B1(n6123), .B2(n6694), .A(n6142), .ZN(n6122) );
  NAND2_X1 U5139 ( .A1(n6611), .A2(n4612), .ZN(n6609) );
  NAND2_X1 U5140 ( .A1(n6170), .A2(n6609), .ZN(n4824) );
  INV_X1 U5141 ( .A(n4824), .ZN(n6648) );
  OAI21_X1 U5142 ( .B1(n6648), .B2(n6612), .A(n4613), .ZN(n4614) );
  NAND2_X1 U5143 ( .A1(n6122), .A2(n4614), .ZN(n6114) );
  AOI21_X1 U5144 ( .B1(n6694), .B2(n4622), .A(n6114), .ZN(n6084) );
  OAI21_X1 U5145 ( .B1(n4615), .B2(n6674), .A(n6084), .ZN(n5783) );
  INV_X1 U5146 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6470) );
  NOR2_X1 U5147 ( .A1(n6821), .A2(n6470), .ZN(n5767) );
  NAND2_X1 U5148 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6595), .ZN(n4617) );
  OAI22_X1 U5149 ( .A1(n4824), .A2(n4618), .B1(n6154), .B2(n4617), .ZN(n4619)
         );
  NAND2_X1 U5150 ( .A1(n4619), .A2(n6155), .ZN(n6139) );
  INV_X1 U5151 ( .A(n4620), .ZN(n4621) );
  NOR2_X1 U5152 ( .A1(n6139), .A2(n4621), .ZN(n6093) );
  INV_X1 U5153 ( .A(n4622), .ZN(n6094) );
  NAND2_X1 U5154 ( .A1(n6093), .A2(n6094), .ZN(n6086) );
  NOR3_X1 U5155 ( .A1(n6086), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5786), 
        .ZN(n4623) );
  AOI211_X1 U5156 ( .C1(n5783), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5767), .B(n4623), .ZN(n4624) );
  OAI21_X1 U5157 ( .B1(n5772), .B2(n6702), .A(n3510), .ZN(U2988) );
  NAND2_X1 U5158 ( .A1(n6019), .A2(n6096), .ZN(n4626) );
  MUX2_X1 U5159 ( .A(n4626), .B(n6019), .S(n4640), .Z(n4627) );
  NAND2_X1 U5160 ( .A1(n5988), .A2(n6723), .ZN(n4635) );
  NOR2_X1 U5161 ( .A1(n5869), .A2(n4628), .ZN(n4629) );
  OR2_X1 U5162 ( .A1(n4630), .A2(n4629), .ZN(n5926) );
  INV_X1 U5163 ( .A(n6084), .ZN(n4631) );
  INV_X1 U5164 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6461) );
  NOR2_X1 U5165 ( .A1(n6821), .A2(n6461), .ZN(n5991) );
  NOR2_X1 U5166 ( .A1(n6086), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6081)
         );
  AOI211_X1 U5167 ( .C1(n4631), .C2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5991), .B(n6081), .ZN(n4632) );
  NAND2_X1 U5168 ( .A1(n4635), .A2(n4634), .ZN(U2991) );
  NAND2_X1 U5169 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4636) );
  AND2_X1 U5170 ( .A1(n4636), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4637)
         );
  XNOR2_X1 U5171 ( .A(n3449), .B(n4638), .ZN(n5748) );
  NAND2_X1 U5172 ( .A1(n4642), .A2(n4641), .ZN(n4644) );
  XNOR2_X1 U5173 ( .A(n4644), .B(n4643), .ZN(n5799) );
  INV_X1 U5174 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5839) );
  XNOR2_X1 U5175 ( .A(n4687), .B(n5839), .ZN(n5838) );
  INV_X1 U5176 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4715) );
  AOI22_X1 U5177 ( .A1(n4072), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3612), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4649) );
  AOI22_X1 U5178 ( .A1(n4645), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3577), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4648) );
  AOI22_X1 U5179 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(n3448), .B1(n3425), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4647) );
  AOI22_X1 U5180 ( .A1(n4231), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4646) );
  NAND4_X1 U5181 ( .A1(n4649), .A2(n4648), .A3(n4647), .A4(n4646), .ZN(n4656)
         );
  AOI22_X1 U5182 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n3719), .B1(n4650), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4654) );
  AOI22_X1 U5183 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n4666), .B1(n3423), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4653) );
  AOI22_X1 U5184 ( .A1(n4673), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3441), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4652) );
  AOI22_X1 U5185 ( .A1(n4668), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4651) );
  NAND4_X1 U5186 ( .A1(n4654), .A2(n4653), .A3(n4652), .A4(n4651), .ZN(n4655)
         );
  NOR2_X1 U5187 ( .A1(n4656), .A2(n4655), .ZN(n4665) );
  NAND2_X1 U5188 ( .A1(n4658), .A2(n4657), .ZN(n4664) );
  XOR2_X1 U5189 ( .A(n4665), .B(n4664), .Z(n4659) );
  NAND2_X1 U5190 ( .A1(n4659), .A2(n4682), .ZN(n4661) );
  OAI21_X1 U5191 ( .B1(n6930), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n6906), 
        .ZN(n4660) );
  OAI211_X1 U5192 ( .C1(n3757), .C2(n4715), .A(n4661), .B(n4660), .ZN(n4662)
         );
  OAI21_X1 U5193 ( .B1(n4685), .B2(n5838), .A(n4662), .ZN(n5760) );
  NOR2_X1 U5194 ( .A1(n4665), .A2(n4664), .ZN(n4681) );
  AOI22_X1 U5195 ( .A1(n3445), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4650), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4672) );
  AOI22_X1 U5196 ( .A1(n4666), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4231), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4671) );
  AOI22_X1 U5197 ( .A1(n3713), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3577), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4670) );
  AOI22_X1 U5198 ( .A1(n4668), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4667), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4669) );
  NAND4_X1 U5199 ( .A1(n4672), .A2(n4671), .A3(n4670), .A4(n4669), .ZN(n4679)
         );
  AOI22_X1 U5200 ( .A1(n4673), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3612), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4677) );
  AOI22_X1 U5201 ( .A1(n3443), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4676) );
  AOI22_X1 U5202 ( .A1(n3448), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3425), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4675) );
  AOI22_X1 U5203 ( .A1(n3424), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3779), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4674) );
  NAND4_X1 U5204 ( .A1(n4677), .A2(n4676), .A3(n4675), .A4(n4674), .ZN(n4678)
         );
  NOR2_X1 U5205 ( .A1(n4679), .A2(n4678), .ZN(n4680) );
  XNOR2_X1 U5206 ( .A(n4681), .B(n4680), .ZN(n4683) );
  NAND2_X1 U5207 ( .A1(n4683), .A2(n4682), .ZN(n4690) );
  NAND2_X1 U5208 ( .A1(n6906), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4684)
         );
  NAND2_X1 U5209 ( .A1(n4685), .A2(n4684), .ZN(n4686) );
  AOI21_X1 U5210 ( .B1(n4691), .B2(EAX_REG_30__SCAN_IN), .A(n4686), .ZN(n4689)
         );
  XNOR2_X1 U5211 ( .A(n4698), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5831)
         );
  AOI21_X1 U5212 ( .B1(n4690), .B2(n4689), .A(n4688), .ZN(n5766) );
  AOI22_X1 U5213 ( .A1(n4691), .A2(EAX_REG_31__SCAN_IN), .B1(n3744), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4692) );
  NAND2_X1 U5214 ( .A1(n6923), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4858) );
  INV_X1 U5215 ( .A(n4858), .ZN(n5344) );
  NAND2_X1 U5216 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n5344), .ZN(n6577) );
  INV_X1 U5217 ( .A(n6577), .ZN(n4693) );
  NAND2_X1 U5218 ( .A1(n7031), .A2(n4693), .ZN(n6069) );
  NAND2_X1 U5219 ( .A1(n5813), .A2(n6561), .ZN(n4705) );
  INV_X1 U5220 ( .A(n7031), .ZN(n7052) );
  NAND2_X1 U5221 ( .A1(n7052), .A2(n4694), .ZN(n6584) );
  NAND2_X1 U5222 ( .A1(n6584), .A2(n6923), .ZN(n4695) );
  NAND2_X1 U5223 ( .A1(n6923), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4697) );
  NAND2_X1 U5224 ( .A1(n6930), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4696) );
  AND2_X1 U5225 ( .A1(n4697), .A2(n4696), .ZN(n4813) );
  INV_X1 U5226 ( .A(n4698), .ZN(n4699) );
  NAND2_X1 U5227 ( .A1(n4699), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4700)
         );
  INV_X1 U5228 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5805) );
  XNOR2_X1 U5229 ( .A(n4700), .B(n5805), .ZN(n5353) );
  INV_X1 U5230 ( .A(REIP_REG_31__SCAN_IN), .ZN(n4701) );
  NOR2_X1 U5231 ( .A1(n6821), .A2(n4701), .ZN(n5788) );
  AOI21_X1 U5232 ( .B1(n6560), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5788), 
        .ZN(n4702) );
  OAI21_X1 U5233 ( .B1(n6566), .B2(n5353), .A(n4702), .ZN(n4703) );
  INV_X1 U5234 ( .A(n4703), .ZN(n4704) );
  OAI211_X1 U5235 ( .C1(n5799), .C2(n6869), .A(n4705), .B(n4704), .ZN(U2955)
         );
  INV_X1 U5236 ( .A(n5817), .ZN(n5825) );
  INV_X1 U5237 ( .A(n4710), .ZN(n4707) );
  AOI22_X1 U5238 ( .A1(n5825), .A2(n3673), .B1(n5818), .B2(n4707), .ZN(n5828)
         );
  AND2_X1 U5239 ( .A1(n5828), .A2(n5829), .ZN(n4709) );
  INV_X1 U5240 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6358) );
  NAND2_X1 U5241 ( .A1(n6906), .A2(n5348), .ZN(n6925) );
  OR3_X1 U5242 ( .A1(n6923), .A2(n6925), .A3(STATE2_REG_3__SCAN_IN), .ZN(n4708) );
  OAI21_X1 U5243 ( .B1(n4709), .B2(n6358), .A(n4708), .ZN(U2790) );
  NAND2_X1 U5244 ( .A1(n4710), .A2(n5829), .ZN(n5342) );
  INV_X1 U5245 ( .A(n5342), .ZN(n4711) );
  INV_X1 U5246 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6954) );
  OAI211_X1 U5247 ( .C1(n4711), .C2(n6954), .A(n5343), .B(n6571), .ZN(U2788)
         );
  INV_X1 U5248 ( .A(n5343), .ZN(n4712) );
  OAI21_X2 U5249 ( .B1(n6581), .B2(n6943), .A(n4712), .ZN(n4764) );
  NAND2_X1 U5250 ( .A1(n4764), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4714) );
  INV_X1 U5251 ( .A(DATAI_13_), .ZN(n5634) );
  OR2_X1 U5252 ( .A1(n4877), .A2(n5634), .ZN(n4770) );
  OAI211_X1 U5253 ( .C1(n4856), .C2(n4715), .A(n4714), .B(n4770), .ZN(U2937)
         );
  INV_X1 U5254 ( .A(EAX_REG_11__SCAN_IN), .ZN(n4717) );
  NAND2_X1 U5255 ( .A1(n4764), .A2(LWORD_REG_11__SCAN_IN), .ZN(n4716) );
  NAND2_X1 U5256 ( .A1(n4795), .A2(DATAI_11_), .ZN(n4792) );
  OAI211_X1 U5257 ( .C1(n4856), .C2(n4717), .A(n4716), .B(n4792), .ZN(U2950)
         );
  INV_X1 U5258 ( .A(EAX_REG_9__SCAN_IN), .ZN(n4719) );
  NAND2_X1 U5259 ( .A1(n4764), .A2(LWORD_REG_9__SCAN_IN), .ZN(n4718) );
  NAND2_X1 U5260 ( .A1(n4795), .A2(DATAI_9_), .ZN(n4797) );
  OAI211_X1 U5261 ( .C1(n4856), .C2(n4719), .A(n4718), .B(n4797), .ZN(U2948)
         );
  INV_X1 U5262 ( .A(EAX_REG_1__SCAN_IN), .ZN(n4721) );
  NAND2_X1 U5263 ( .A1(n4764), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4720) );
  NAND2_X1 U5264 ( .A1(n4795), .A2(DATAI_1_), .ZN(n4786) );
  OAI211_X1 U5265 ( .C1(n4856), .C2(n4721), .A(n4720), .B(n4786), .ZN(U2940)
         );
  INV_X1 U5266 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n4723) );
  INV_X1 U5267 ( .A(n4856), .ZN(n4740) );
  INV_X1 U5268 ( .A(DATAI_0_), .ZN(n4916) );
  NOR2_X1 U5269 ( .A1(n4877), .A2(n4916), .ZN(n4736) );
  AOI21_X1 U5270 ( .B1(n4740), .B2(EAX_REG_0__SCAN_IN), .A(n4736), .ZN(n4722)
         );
  OAI21_X1 U5271 ( .B1(n4743), .B2(n4723), .A(n4722), .ZN(U2939) );
  INV_X1 U5272 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n4725) );
  INV_X1 U5273 ( .A(DATAI_12_), .ZN(n6238) );
  NOR2_X1 U5274 ( .A1(n4877), .A2(n6238), .ZN(n4731) );
  AOI21_X1 U5275 ( .B1(n4740), .B2(EAX_REG_28__SCAN_IN), .A(n4731), .ZN(n4724)
         );
  OAI21_X1 U5276 ( .B1(n4743), .B2(n4725), .A(n4724), .ZN(U2936) );
  INV_X1 U5277 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n4727) );
  INV_X1 U5278 ( .A(DATAI_3_), .ZN(n4884) );
  NOR2_X1 U5279 ( .A1(n4877), .A2(n4884), .ZN(n4728) );
  AOI21_X1 U5280 ( .B1(n4740), .B2(EAX_REG_19__SCAN_IN), .A(n4728), .ZN(n4726)
         );
  OAI21_X1 U5281 ( .B1(n4743), .B2(n4727), .A(n4726), .ZN(U2927) );
  INV_X1 U5282 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n4730) );
  AOI21_X1 U5283 ( .B1(n4740), .B2(EAX_REG_3__SCAN_IN), .A(n4728), .ZN(n4729)
         );
  OAI21_X1 U5284 ( .B1(n4743), .B2(n4730), .A(n4729), .ZN(U2942) );
  INV_X1 U5285 ( .A(LWORD_REG_12__SCAN_IN), .ZN(n4733) );
  AOI21_X1 U5286 ( .B1(n4740), .B2(EAX_REG_12__SCAN_IN), .A(n4731), .ZN(n4732)
         );
  OAI21_X1 U5287 ( .B1(n4743), .B2(n4733), .A(n4732), .ZN(U2951) );
  INV_X1 U5288 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n4735) );
  INV_X1 U5289 ( .A(DATAI_5_), .ZN(n5046) );
  NOR2_X1 U5290 ( .A1(n4877), .A2(n5046), .ZN(n4739) );
  AOI21_X1 U5291 ( .B1(n4740), .B2(EAX_REG_21__SCAN_IN), .A(n4739), .ZN(n4734)
         );
  OAI21_X1 U5292 ( .B1(n4743), .B2(n4735), .A(n4734), .ZN(U2929) );
  INV_X1 U5293 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n4738) );
  AOI21_X1 U5294 ( .B1(n4740), .B2(EAX_REG_16__SCAN_IN), .A(n4736), .ZN(n4737)
         );
  OAI21_X1 U5295 ( .B1(n4743), .B2(n4738), .A(n4737), .ZN(U2924) );
  INV_X1 U5296 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n4742) );
  AOI21_X1 U5297 ( .B1(n4740), .B2(EAX_REG_5__SCAN_IN), .A(n4739), .ZN(n4741)
         );
  OAI21_X1 U5298 ( .B1(n4743), .B2(n4742), .A(n4741), .ZN(U2944) );
  INV_X1 U5299 ( .A(EAX_REG_15__SCAN_IN), .ZN(n4745) );
  INV_X1 U5300 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4744) );
  INV_X1 U5301 ( .A(DATAI_15_), .ZN(n6296) );
  OAI222_X1 U5302 ( .A1(n4856), .A2(n4745), .B1(n4744), .B2(n4743), .C1(n4877), 
        .C2(n6296), .ZN(U2954) );
  AND2_X1 U5303 ( .A1(n3432), .A2(n4747), .ZN(n4748) );
  AND2_X1 U5304 ( .A1(n4749), .A2(n4748), .ZN(n4962) );
  OAI22_X1 U5305 ( .A1(n3792), .A2(n4962), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6183), .ZN(n6877) );
  OAI22_X1 U5306 ( .A1(n5348), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6924), .ZN(n4750) );
  AOI21_X1 U5307 ( .B1(n6877), .B2(n5775), .A(n4750), .ZN(n4761) );
  INV_X1 U5308 ( .A(n5818), .ZN(n4751) );
  AOI21_X1 U5309 ( .B1(n4958), .B2(n5827), .A(n4751), .ZN(n4752) );
  OR2_X1 U5310 ( .A1(n4753), .A2(n4752), .ZN(n4759) );
  INV_X1 U5311 ( .A(n4879), .ZN(n4945) );
  NAND2_X1 U5312 ( .A1(n5826), .A2(n4908), .ZN(n4754) );
  OAI211_X1 U5313 ( .C1(n4872), .C2(n4746), .A(n4755), .B(n4754), .ZN(n4756)
         );
  AOI21_X1 U5314 ( .B1(n5817), .B2(n4945), .A(n4756), .ZN(n4758) );
  NAND3_X1 U5315 ( .A1(n4759), .A2(n4758), .A3(n4757), .ZN(n4969) );
  INV_X1 U5316 ( .A(n4969), .ZN(n6880) );
  NAND2_X1 U5317 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n6914) );
  INV_X1 U5318 ( .A(n6914), .ZN(n5739) );
  NAND2_X1 U5319 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5739), .ZN(n6915) );
  INV_X1 U5320 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6894) );
  OAI22_X1 U5321 ( .A1(n6880), .A2(n6928), .B1(n6915), .B2(n6894), .ZN(n6873)
         );
  AOI21_X1 U5322 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6923), .A(n6873), .ZN(
        n6189) );
  AND2_X1 U5323 ( .A1(n4958), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6876)
         );
  AOI22_X1 U5324 ( .A1(n6876), .A2(n5775), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6189), .ZN(n4760) );
  OAI21_X1 U5325 ( .B1(n4761), .B2(n6189), .A(n4760), .ZN(U3461) );
  INV_X1 U5326 ( .A(EAX_REG_4__SCAN_IN), .ZN(n4763) );
  NAND2_X1 U5327 ( .A1(n4764), .A2(LWORD_REG_4__SCAN_IN), .ZN(n4762) );
  NAND2_X1 U5328 ( .A1(n4795), .A2(DATAI_4_), .ZN(n4780) );
  OAI211_X1 U5329 ( .C1(n4856), .C2(n4763), .A(n4762), .B(n4780), .ZN(U2943)
         );
  INV_X1 U5330 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4766) );
  NAND2_X1 U5331 ( .A1(n4806), .A2(UWORD_REG_14__SCAN_IN), .ZN(n4765) );
  NAND2_X1 U5332 ( .A1(n4795), .A2(DATAI_14_), .ZN(n4767) );
  OAI211_X1 U5333 ( .C1(n4856), .C2(n4766), .A(n4765), .B(n4767), .ZN(U2938)
         );
  INV_X1 U5334 ( .A(EAX_REG_14__SCAN_IN), .ZN(n4769) );
  NAND2_X1 U5335 ( .A1(n4764), .A2(LWORD_REG_14__SCAN_IN), .ZN(n4768) );
  OAI211_X1 U5336 ( .C1(n4856), .C2(n4769), .A(n4768), .B(n4767), .ZN(U2953)
         );
  INV_X1 U5337 ( .A(EAX_REG_13__SCAN_IN), .ZN(n4772) );
  NAND2_X1 U5338 ( .A1(n4806), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4771) );
  OAI211_X1 U5339 ( .C1(n4856), .C2(n4772), .A(n4771), .B(n4770), .ZN(U2952)
         );
  INV_X1 U5340 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4774) );
  NAND2_X1 U5341 ( .A1(n4764), .A2(LWORD_REG_7__SCAN_IN), .ZN(n4773) );
  NAND2_X1 U5342 ( .A1(n4795), .A2(DATAI_7_), .ZN(n4803) );
  OAI211_X1 U5343 ( .C1(n4856), .C2(n4774), .A(n4773), .B(n4803), .ZN(U2946)
         );
  INV_X1 U5344 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4776) );
  NAND2_X1 U5345 ( .A1(n4806), .A2(UWORD_REG_6__SCAN_IN), .ZN(n4775) );
  NAND2_X1 U5346 ( .A1(n4795), .A2(DATAI_6_), .ZN(n4777) );
  OAI211_X1 U5347 ( .C1(n4856), .C2(n4776), .A(n4775), .B(n4777), .ZN(U2930)
         );
  INV_X1 U5348 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4779) );
  NAND2_X1 U5349 ( .A1(n4806), .A2(LWORD_REG_6__SCAN_IN), .ZN(n4778) );
  OAI211_X1 U5350 ( .C1(n4856), .C2(n4779), .A(n4778), .B(n4777), .ZN(U2945)
         );
  INV_X1 U5351 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4782) );
  NAND2_X1 U5352 ( .A1(n4806), .A2(UWORD_REG_4__SCAN_IN), .ZN(n4781) );
  OAI211_X1 U5353 ( .C1(n4856), .C2(n4782), .A(n4781), .B(n4780), .ZN(U2928)
         );
  NAND2_X1 U5354 ( .A1(n4764), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4783) );
  NAND2_X1 U5355 ( .A1(n4795), .A2(DATAI_8_), .ZN(n4789) );
  OAI211_X1 U5356 ( .C1(n4856), .C2(n4784), .A(n4783), .B(n4789), .ZN(U2932)
         );
  INV_X1 U5357 ( .A(EAX_REG_18__SCAN_IN), .ZN(n6961) );
  NAND2_X1 U5358 ( .A1(n4764), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4785) );
  NAND2_X1 U5359 ( .A1(n4795), .A2(DATAI_2_), .ZN(n4807) );
  OAI211_X1 U5360 ( .C1(n4856), .C2(n6961), .A(n4785), .B(n4807), .ZN(U2926)
         );
  INV_X1 U5361 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4788) );
  NAND2_X1 U5362 ( .A1(n4764), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4787) );
  OAI211_X1 U5363 ( .C1(n4856), .C2(n4788), .A(n4787), .B(n4786), .ZN(U2925)
         );
  INV_X1 U5364 ( .A(EAX_REG_8__SCAN_IN), .ZN(n4791) );
  NAND2_X1 U5365 ( .A1(n4764), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4790) );
  OAI211_X1 U5366 ( .C1(n4856), .C2(n4791), .A(n4790), .B(n4789), .ZN(U2947)
         );
  INV_X1 U5367 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4794) );
  NAND2_X1 U5368 ( .A1(n4764), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4793) );
  OAI211_X1 U5369 ( .C1(n4856), .C2(n4794), .A(n4793), .B(n4792), .ZN(U2935)
         );
  NAND2_X1 U5370 ( .A1(n4764), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4796) );
  NAND2_X1 U5371 ( .A1(n4795), .A2(DATAI_10_), .ZN(n4800) );
  OAI211_X1 U5372 ( .C1(n4856), .C2(n4863), .A(n4796), .B(n4800), .ZN(U2934)
         );
  INV_X1 U5373 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4799) );
  NAND2_X1 U5374 ( .A1(n4806), .A2(UWORD_REG_9__SCAN_IN), .ZN(n4798) );
  OAI211_X1 U5375 ( .C1(n4856), .C2(n4799), .A(n4798), .B(n4797), .ZN(U2933)
         );
  INV_X1 U5376 ( .A(EAX_REG_10__SCAN_IN), .ZN(n4802) );
  NAND2_X1 U5377 ( .A1(n4806), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4801) );
  OAI211_X1 U5378 ( .C1(n4856), .C2(n4802), .A(n4801), .B(n4800), .ZN(U2949)
         );
  INV_X1 U5379 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4805) );
  NAND2_X1 U5380 ( .A1(n4806), .A2(UWORD_REG_7__SCAN_IN), .ZN(n4804) );
  OAI211_X1 U5381 ( .C1(n4856), .C2(n4805), .A(n4804), .B(n4803), .ZN(U2931)
         );
  INV_X1 U5382 ( .A(EAX_REG_2__SCAN_IN), .ZN(n4809) );
  NAND2_X1 U5383 ( .A1(n4806), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4808) );
  OAI211_X1 U5384 ( .C1(n4856), .C2(n4809), .A(n4808), .B(n4807), .ZN(U2941)
         );
  NOR2_X1 U5385 ( .A1(n4811), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4812)
         );
  OR2_X1 U5386 ( .A1(n4810), .A2(n4812), .ZN(n6718) );
  INV_X1 U5387 ( .A(n4813), .ZN(n4814) );
  OAI21_X1 U5388 ( .B1(n6560), .B2(n4814), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4819) );
  XOR2_X1 U5389 ( .A(n4816), .B(n4815), .Z(n5475) );
  INV_X1 U5390 ( .A(n5475), .ZN(n4817) );
  AOI22_X1 U5391 ( .A1(n4817), .A2(n6561), .B1(n6789), .B2(REIP_REG_0__SCAN_IN), .ZN(n4818) );
  OAI211_X1 U5392 ( .C1(n6718), .C2(n6869), .A(n4819), .B(n4818), .ZN(U2986)
         );
  NAND2_X1 U5393 ( .A1(n4821), .A2(n4820), .ZN(n4822) );
  XOR2_X1 U5394 ( .A(n4823), .B(n4822), .Z(n5487) );
  AOI21_X1 U5395 ( .B1(n6170), .B2(n6649), .A(n6610), .ZN(n6660) );
  OAI21_X1 U5396 ( .B1(n6651), .B2(n6653), .A(n6660), .ZN(n6630) );
  OAI21_X1 U5397 ( .B1(n4824), .B2(n6649), .A(n6651), .ZN(n6632) );
  NAND2_X1 U5398 ( .A1(n6632), .A2(n6653), .ZN(n6639) );
  INV_X1 U5399 ( .A(n6639), .ZN(n4825) );
  AOI22_X1 U5400 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n6630), .B1(n4825), 
        .B2(n6620), .ZN(n4830) );
  INV_X1 U5401 ( .A(n4845), .ZN(n4826) );
  AOI21_X1 U5402 ( .B1(n4834), .B2(n4827), .A(n4826), .ZN(n5456) );
  INV_X1 U5403 ( .A(REIP_REG_3__SCAN_IN), .ZN(n4828) );
  NOR2_X1 U5404 ( .A1(n6821), .A2(n4828), .ZN(n5481) );
  AOI21_X1 U5405 ( .B1(n6721), .B2(n5456), .A(n5481), .ZN(n4829) );
  OAI211_X1 U5406 ( .C1(n5487), .C2(n6702), .A(n4830), .B(n4829), .ZN(U3015)
         );
  AOI21_X1 U5407 ( .B1(n4832), .B2(n4831), .A(n4843), .ZN(n5485) );
  INV_X1 U5408 ( .A(n5485), .ZN(n5458) );
  AOI22_X1 U5409 ( .A1(n6507), .A2(n5456), .B1(n6200), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4833) );
  OAI21_X1 U5410 ( .B1(n5458), .B2(n5958), .A(n4833), .ZN(U2856) );
  OAI21_X1 U5411 ( .B1(n4836), .B2(n4835), .A(n4834), .ZN(n6655) );
  INV_X1 U5412 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4840) );
  INV_X1 U5413 ( .A(n4837), .ZN(n4839) );
  INV_X1 U5414 ( .A(n4831), .ZN(n4838) );
  AOI21_X1 U5415 ( .B1(n4839), .B2(n4851), .A(n4838), .ZN(n6514) );
  INV_X1 U5416 ( .A(n6514), .ZN(n4885) );
  OAI222_X1 U5417 ( .A1(n6655), .A2(n5956), .B1(n4840), .B2(n6510), .C1(n4885), 
        .C2(n5958), .ZN(U2857) );
  INV_X1 U5418 ( .A(n4841), .ZN(n4842) );
  XNOR2_X1 U5419 ( .A(n4843), .B(n4842), .ZN(n6742) );
  INV_X1 U5420 ( .A(n6742), .ZN(n4917) );
  AND2_X1 U5421 ( .A1(n4845), .A2(n4844), .ZN(n4846) );
  NOR2_X1 U5422 ( .A1(n6504), .A2(n4846), .ZN(n6736) );
  AOI22_X1 U5423 ( .A1(n6507), .A2(n6736), .B1(n6200), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4847) );
  OAI21_X1 U5424 ( .B1(n4917), .B2(n5958), .A(n4847), .ZN(U2855) );
  OAI21_X1 U5425 ( .B1(n5790), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4848), 
        .ZN(n6719) );
  OAI222_X1 U5426 ( .A1(n5956), .A2(n6719), .B1(n6510), .B2(n4849), .C1(n5958), 
        .C2(n5475), .ZN(U2859) );
  XNOR2_X1 U5427 ( .A(n5368), .B(n4850), .ZN(n6613) );
  INV_X1 U5428 ( .A(n6613), .ZN(n4854) );
  OAI21_X1 U5429 ( .B1(n4853), .B2(n4852), .A(n4851), .ZN(n5525) );
  OAI222_X1 U5430 ( .A1(n4854), .A2(n5956), .B1(n6510), .B2(n5365), .C1(n5958), 
        .C2(n5525), .ZN(U2858) );
  INV_X1 U5431 ( .A(n4958), .ZN(n4947) );
  OR2_X1 U5432 ( .A1(n4880), .A2(n4947), .ZN(n4855) );
  NAND2_X1 U5433 ( .A1(n4856), .A2(n4855), .ZN(n4857) );
  NAND2_X1 U5434 ( .A1(n6406), .A2(n3643), .ZN(n5301) );
  OR2_X1 U5435 ( .A1(n6906), .A2(n4858), .ZN(n6902) );
  NOR2_X4 U5438 ( .A1(n6585), .A2(n6406), .ZN(n6198) );
  AOI22_X1 U5439 ( .A1(n6585), .A2(UWORD_REG_11__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4859) );
  OAI21_X1 U5440 ( .B1(n4794), .B2(n5301), .A(n4859), .ZN(U2896) );
  AOI22_X1 U5441 ( .A1(n6585), .A2(UWORD_REG_8__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4860) );
  OAI21_X1 U5442 ( .B1(n4784), .B2(n5301), .A(n4860), .ZN(U2899) );
  AOI22_X1 U5443 ( .A1(n6585), .A2(UWORD_REG_9__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4861) );
  OAI21_X1 U5444 ( .B1(n4799), .B2(n5301), .A(n4861), .ZN(U2898) );
  INV_X1 U5445 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4863) );
  AOI22_X1 U5446 ( .A1(n6585), .A2(UWORD_REG_10__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4862) );
  OAI21_X1 U5447 ( .B1(n4863), .B2(n5301), .A(n4862), .ZN(U2897) );
  AOI22_X1 U5448 ( .A1(n6585), .A2(UWORD_REG_13__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4864) );
  OAI21_X1 U5449 ( .B1(n4715), .B2(n5301), .A(n4864), .ZN(U2894) );
  INV_X1 U5450 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4866) );
  AOI22_X1 U5451 ( .A1(n6585), .A2(UWORD_REG_5__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4865) );
  OAI21_X1 U5452 ( .B1(n4866), .B2(n5301), .A(n4865), .ZN(U2902) );
  AOI22_X1 U5453 ( .A1(n6585), .A2(UWORD_REG_4__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4867) );
  OAI21_X1 U5454 ( .B1(n4782), .B2(n5301), .A(n4867), .ZN(U2903) );
  AOI22_X1 U5455 ( .A1(n6585), .A2(UWORD_REG_7__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4868) );
  OAI21_X1 U5456 ( .B1(n4805), .B2(n5301), .A(n4868), .ZN(U2900) );
  AOI22_X1 U5457 ( .A1(n6585), .A2(UWORD_REG_6__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4869) );
  OAI21_X1 U5458 ( .B1(n4776), .B2(n5301), .A(n4869), .ZN(U2901) );
  INV_X1 U5459 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4871) );
  AOI22_X1 U5460 ( .A1(n6585), .A2(UWORD_REG_12__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4870) );
  OAI21_X1 U5461 ( .B1(n4871), .B2(n5301), .A(n4870), .ZN(U2895) );
  OR2_X1 U5462 ( .A1(n6928), .A2(n4872), .ZN(n4875) );
  OAI22_X1 U5463 ( .A1(n3432), .A2(n4875), .B1(n4874), .B2(n4873), .ZN(n4876)
         );
  INV_X1 U5464 ( .A(n4876), .ZN(n4878) );
  NAND2_X1 U5465 ( .A1(n3653), .A2(n3746), .ZN(n4881) );
  INV_X1 U5466 ( .A(n7077), .ZN(n4883) );
  AND2_X1 U5467 ( .A1(n5155), .A2(n3746), .ZN(n4882) );
  NAND2_X1 U5468 ( .A1(n3422), .A2(n4882), .ZN(n6963) );
  INV_X1 U5469 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6412) );
  OAI222_X1 U5470 ( .A1(n5458), .A2(n5976), .B1(n5975), .B2(n4884), .C1(n3422), 
        .C2(n6412), .ZN(U2888) );
  OAI222_X1 U5471 ( .A1(n4885), .A2(n5976), .B1(n5975), .B2(n6962), .C1(n3422), 
        .C2(n4809), .ZN(U2889) );
  INV_X1 U5472 ( .A(DATAI_1_), .ZN(n6290) );
  OAI222_X1 U5473 ( .A1(n5525), .A2(n5976), .B1(n5975), .B2(n6290), .C1(n3422), 
        .C2(n4721), .ZN(U2890) );
  NOR2_X2 U5474 ( .A1(n5161), .A2(n4886), .ZN(n7047) );
  INV_X1 U5475 ( .A(n7047), .ZN(n5415) );
  OAI21_X1 U5476 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6916), .A(n5175), 
        .ZN(n7050) );
  INV_X1 U5477 ( .A(n7050), .ZN(n7029) );
  OR2_X1 U5478 ( .A1(n4889), .A2(n3821), .ZN(n4990) );
  NAND2_X1 U5479 ( .A1(n4890), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5091) );
  NOR2_X1 U5480 ( .A1(n4990), .A2(n5091), .ZN(n4981) );
  NOR2_X1 U5481 ( .A1(n4981), .A2(n7052), .ZN(n4896) );
  OR2_X1 U5482 ( .A1(n5548), .A2(n3792), .ZN(n7044) );
  INV_X1 U5483 ( .A(n7044), .ZN(n7023) );
  NOR2_X1 U5484 ( .A1(n4892), .A2(n5357), .ZN(n5007) );
  INV_X1 U5485 ( .A(n5315), .ZN(n4894) );
  AOI21_X1 U5486 ( .B1(n7023), .B2(n5007), .A(n4894), .ZN(n4898) );
  OR2_X1 U5487 ( .A1(n5172), .A2(n7024), .ZN(n5125) );
  AOI22_X1 U5488 ( .A1(n4896), .A2(n4898), .B1(n7052), .B2(n5125), .ZN(n4895)
         );
  NAND2_X1 U5489 ( .A1(n7029), .A2(n4895), .ZN(n5311) );
  NAND2_X1 U5490 ( .A1(DATAI_0_), .A2(n5175), .ZN(n7059) );
  INV_X1 U5491 ( .A(n4896), .ZN(n4897) );
  OAI22_X1 U5492 ( .A1(n4898), .A2(n4897), .B1(n6906), .B2(n5125), .ZN(n5310)
         );
  AOI22_X1 U5493 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n5311), .B1(n5578), 
        .B2(n5310), .ZN(n4902) );
  AND2_X1 U5494 ( .A1(n6561), .A2(DATAI_24_), .ZN(n7056) );
  NAND2_X1 U5495 ( .A1(n4976), .A2(n5746), .ZN(n4899) );
  NAND2_X1 U5496 ( .A1(n4976), .A2(n6990), .ZN(n4900) );
  AND2_X1 U5497 ( .A1(n6561), .A2(DATAI_16_), .ZN(n7048) );
  AOI22_X1 U5498 ( .A1(n7056), .A2(n5312), .B1(n5372), .B2(n7048), .ZN(n4901)
         );
  OAI211_X1 U5499 ( .C1(n5315), .C2(n5415), .A(n4902), .B(n4901), .ZN(U3076)
         );
  NOR2_X2 U5500 ( .A1(n5161), .A2(n5812), .ZN(n7182) );
  INV_X1 U5501 ( .A(n7182), .ZN(n5397) );
  NAND2_X1 U5502 ( .A1(DATAI_7_), .A2(n5175), .ZN(n7190) );
  AOI22_X1 U5503 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n5311), .B1(n5584), 
        .B2(n5310), .ZN(n4904) );
  AND2_X1 U5504 ( .A1(n6561), .A2(DATAI_31_), .ZN(n7183) );
  AND2_X1 U5505 ( .A1(n6561), .A2(DATAI_23_), .ZN(n7186) );
  AOI22_X1 U5506 ( .A1(n5312), .A2(n7183), .B1(n5372), .B2(n7186), .ZN(n4903)
         );
  OAI211_X1 U5507 ( .C1(n5315), .C2(n5397), .A(n4904), .B(n4903), .ZN(U3083)
         );
  NOR2_X2 U5508 ( .A1(n5161), .A2(n4905), .ZN(n7106) );
  INV_X1 U5509 ( .A(n7106), .ZN(n5403) );
  NAND2_X1 U5510 ( .A1(DATAI_3_), .A2(n5175), .ZN(n7111) );
  AOI22_X1 U5511 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n5311), .B1(n5574), 
        .B2(n5310), .ZN(n4907) );
  AND2_X1 U5512 ( .A1(n6561), .A2(DATAI_27_), .ZN(n7108) );
  AND2_X1 U5513 ( .A1(n6561), .A2(DATAI_19_), .ZN(n7107) );
  AOI22_X1 U5514 ( .A1(n5312), .A2(n7108), .B1(n5372), .B2(n7107), .ZN(n4906)
         );
  OAI211_X1 U5515 ( .C1(n5315), .C2(n5403), .A(n4907), .B(n4906), .ZN(U3079)
         );
  NOR2_X2 U5516 ( .A1(n5161), .A2(n4908), .ZN(n7092) );
  INV_X1 U5517 ( .A(n7092), .ZN(n5409) );
  NAND2_X1 U5518 ( .A1(DATAI_2_), .A2(n5175), .ZN(n7097) );
  AOI22_X1 U5519 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n5311), .B1(n5554), 
        .B2(n5310), .ZN(n4910) );
  AND2_X1 U5520 ( .A1(n6561), .A2(DATAI_26_), .ZN(n7094) );
  AND2_X1 U5521 ( .A1(n6561), .A2(DATAI_18_), .ZN(n7093) );
  AOI22_X1 U5522 ( .A1(n5312), .A2(n7094), .B1(n5372), .B2(n7093), .ZN(n4909)
         );
  OAI211_X1 U5523 ( .C1(n5315), .C2(n5409), .A(n4910), .B(n4909), .ZN(U3078)
         );
  NOR2_X2 U5524 ( .A1(n5161), .A2(n3500), .ZN(n7148) );
  INV_X1 U5525 ( .A(n7148), .ZN(n5391) );
  NAND2_X1 U5526 ( .A1(DATAI_6_), .A2(n5175), .ZN(n7153) );
  AOI22_X1 U5527 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n5311), .B1(n5566), 
        .B2(n5310), .ZN(n4912) );
  AND2_X1 U5528 ( .A1(n6561), .A2(DATAI_30_), .ZN(n7150) );
  AND2_X1 U5529 ( .A1(n6561), .A2(DATAI_22_), .ZN(n7149) );
  AOI22_X1 U5530 ( .A1(n5312), .A2(n7150), .B1(n5372), .B2(n7149), .ZN(n4911)
         );
  OAI211_X1 U5531 ( .C1(n5315), .C2(n5391), .A(n4912), .B(n4911), .ZN(U3082)
         );
  NOR2_X2 U5532 ( .A1(n5161), .A2(n4913), .ZN(n7071) );
  INV_X1 U5533 ( .A(n7071), .ZN(n5430) );
  NAND2_X1 U5534 ( .A1(DATAI_1_), .A2(n5175), .ZN(n7076) );
  AOI22_X1 U5535 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n5311), .B1(n5570), 
        .B2(n5310), .ZN(n4915) );
  AND2_X1 U5536 ( .A1(n6561), .A2(DATAI_25_), .ZN(n7072) );
  AND2_X1 U5537 ( .A1(n6561), .A2(DATAI_17_), .ZN(n7073) );
  AOI22_X1 U5538 ( .A1(n5312), .A2(n7072), .B1(n5372), .B2(n7073), .ZN(n4914)
         );
  OAI211_X1 U5539 ( .C1(n5315), .C2(n5430), .A(n4915), .B(n4914), .ZN(U3077)
         );
  INV_X1 U5540 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6408) );
  OAI222_X1 U5541 ( .A1(n5976), .A2(n5475), .B1(n3422), .B2(n6408), .C1(n4916), 
        .C2(n5975), .ZN(U2891) );
  INV_X1 U5542 ( .A(DATAI_4_), .ZN(n6344) );
  OAI222_X1 U5543 ( .A1(n5976), .A2(n4917), .B1(n3422), .B2(n4763), .C1(n6344), 
        .C2(n5975), .ZN(U2887) );
  NOR2_X1 U5544 ( .A1(n4923), .A2(n4976), .ZN(n4925) );
  AND2_X1 U5545 ( .A1(n7031), .A2(n6930), .ZN(n6991) );
  INV_X1 U5546 ( .A(n6991), .ZN(n7039) );
  OAI21_X1 U5547 ( .B1(n4925), .B2(n6069), .A(n7039), .ZN(n4921) );
  NAND2_X1 U5548 ( .A1(n5548), .A2(n5093), .ZN(n7008) );
  INV_X1 U5549 ( .A(n7008), .ZN(n6982) );
  NOR2_X1 U5550 ( .A1(n4918), .A2(n6889), .ZN(n5276) );
  AOI21_X1 U5551 ( .B1(n6982), .B2(n5007), .A(n5276), .ZN(n4922) );
  NAND3_X1 U5552 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5002) );
  AOI21_X1 U5553 ( .B1(n7052), .B2(n5002), .A(n7050), .ZN(n4919) );
  INV_X1 U5554 ( .A(n4919), .ZN(n4920) );
  AOI21_X1 U5555 ( .B1(n4921), .B2(n4922), .A(n4920), .ZN(n5280) );
  INV_X1 U5556 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4928) );
  OAI22_X1 U5557 ( .A1(n4922), .A2(n7052), .B1(n5002), .B2(n6906), .ZN(n5275)
         );
  INV_X1 U5558 ( .A(n4923), .ZN(n4924) );
  NAND3_X1 U5559 ( .A1(n4924), .A2(n6990), .A3(n3821), .ZN(n5255) );
  AOI22_X1 U5560 ( .A1(n5584), .A2(n5275), .B1(n7186), .B2(n5274), .ZN(n4927)
         );
  NAND2_X1 U5561 ( .A1(n4925), .A2(n5746), .ZN(n5005) );
  AOI22_X1 U5562 ( .A1(n5283), .A2(n7183), .B1(n7182), .B2(n5276), .ZN(n4926)
         );
  OAI211_X1 U5563 ( .C1(n5280), .C2(n4928), .A(n4927), .B(n4926), .ZN(U3147)
         );
  INV_X1 U5564 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4931) );
  AOI22_X1 U5565 ( .A1(n5554), .A2(n5275), .B1(n7093), .B2(n5274), .ZN(n4930)
         );
  AOI22_X1 U5566 ( .A1(n5283), .A2(n7094), .B1(n7092), .B2(n5276), .ZN(n4929)
         );
  OAI211_X1 U5567 ( .C1(n5280), .C2(n4931), .A(n4930), .B(n4929), .ZN(U3142)
         );
  INV_X1 U5568 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4934) );
  AOI22_X1 U5569 ( .A1(n5574), .A2(n5275), .B1(n7107), .B2(n5274), .ZN(n4933)
         );
  AOI22_X1 U5570 ( .A1(n5283), .A2(n7108), .B1(n7106), .B2(n5276), .ZN(n4932)
         );
  OAI211_X1 U5571 ( .C1(n5280), .C2(n4934), .A(n4933), .B(n4932), .ZN(U3143)
         );
  INV_X1 U5572 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4937) );
  AOI22_X1 U5573 ( .A1(n5578), .A2(n5275), .B1(n7048), .B2(n5274), .ZN(n4936)
         );
  AOI22_X1 U5574 ( .A1(n5283), .A2(n7056), .B1(n7047), .B2(n5276), .ZN(n4935)
         );
  OAI211_X1 U5575 ( .C1(n5280), .C2(n4937), .A(n4936), .B(n4935), .ZN(U3140)
         );
  INV_X1 U5576 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4940) );
  AOI22_X1 U5577 ( .A1(n5566), .A2(n5275), .B1(n7149), .B2(n5274), .ZN(n4939)
         );
  AOI22_X1 U5578 ( .A1(n5283), .A2(n7150), .B1(n7148), .B2(n5276), .ZN(n4938)
         );
  OAI211_X1 U5579 ( .C1(n5280), .C2(n4940), .A(n4939), .B(n4938), .ZN(U3146)
         );
  AOI21_X1 U5580 ( .B1(n4941), .B2(n5774), .A(n4950), .ZN(n4942) );
  NOR2_X1 U5581 ( .A1(n3612), .A2(n4942), .ZN(n6192) );
  NAND2_X1 U5582 ( .A1(n4947), .A2(n4941), .ZN(n4944) );
  NAND2_X1 U5583 ( .A1(n4958), .A2(n3513), .ZN(n6182) );
  INV_X1 U5584 ( .A(n6182), .ZN(n4943) );
  AOI21_X1 U5585 ( .B1(n4944), .B2(n5780), .A(n4943), .ZN(n4952) );
  INV_X1 U5586 ( .A(n4941), .ZN(n5779) );
  NOR2_X1 U5587 ( .A1(n4946), .A2(n4945), .ZN(n4956) );
  AOI21_X1 U5588 ( .B1(n5780), .B2(n5779), .A(n4956), .ZN(n4949) );
  NOR3_X1 U5589 ( .A1(n4947), .A2(n5780), .A3(n3513), .ZN(n4948) );
  NOR2_X1 U5590 ( .A1(n4949), .A2(n4948), .ZN(n4951) );
  MUX2_X1 U5591 ( .A(n4952), .B(n4951), .S(n4950), .Z(n4954) );
  INV_X1 U5592 ( .A(n4962), .ZN(n6185) );
  NAND2_X1 U5593 ( .A1(n5548), .A2(n6185), .ZN(n4953) );
  OAI211_X1 U5594 ( .C1(n6192), .C2(n4957), .A(n4954), .B(n4953), .ZN(n6191)
         );
  MUX2_X1 U5595 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6191), .S(n4969), 
        .Z(n6888) );
  NAND2_X1 U5596 ( .A1(n5348), .A2(n6888), .ZN(n4967) );
  XNOR2_X1 U5597 ( .A(n4941), .B(n5774), .ZN(n4955) );
  MUX2_X1 U5598 ( .A(n4957), .B(n4956), .S(n4955), .Z(n4961) );
  NAND2_X1 U5599 ( .A1(n4958), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4959) );
  MUX2_X1 U5600 ( .A(n4959), .B(n6182), .S(n5774), .Z(n4960) );
  OAI211_X1 U5601 ( .C1(n4892), .C2(n4962), .A(n4961), .B(n4960), .ZN(n5776)
         );
  NOR2_X1 U5602 ( .A1(n4969), .A2(n5780), .ZN(n4963) );
  AOI21_X1 U5603 ( .B1(n5776), .B2(n4969), .A(n4963), .ZN(n6886) );
  NAND2_X1 U5604 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6894), .ZN(n4966) );
  INV_X1 U5605 ( .A(n4964), .ZN(n4965) );
  OAI22_X1 U5606 ( .A1(n4967), .A2(n6886), .B1(n4966), .B2(n4965), .ZN(n6898)
         );
  INV_X1 U5607 ( .A(n4968), .ZN(n4975) );
  MUX2_X1 U5608 ( .A(n4969), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n4974) );
  INV_X1 U5609 ( .A(n4971), .ZN(n4972) );
  NOR2_X1 U5610 ( .A1(n3431), .A2(n4972), .ZN(n4973) );
  XNOR2_X1 U5611 ( .A(n4973), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6732)
         );
  OR3_X1 U5612 ( .A1(n6732), .A2(STATE2_REG_1__SCAN_IN), .A3(n3432), .ZN(n6871) );
  OAI21_X1 U5613 ( .B1(n4974), .B2(n3846), .A(n6871), .ZN(n6890) );
  AOI21_X1 U5614 ( .B1(n6898), .B2(n4975), .A(n6890), .ZN(n6921) );
  INV_X1 U5615 ( .A(n6915), .ZN(n6920) );
  AOI21_X1 U5616 ( .B1(n6920), .B2(FLUSH_REG_SCAN_IN), .A(n5175), .ZN(n5738)
         );
  OAI21_X1 U5617 ( .B1(n6921), .B2(n6915), .A(n5738), .ZN(n5150) );
  OAI21_X1 U5618 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5348), .A(n5150), .ZN(
        n5741) );
  INV_X1 U5619 ( .A(n5548), .ZN(n5451) );
  NAND2_X1 U5620 ( .A1(n5150), .A2(n7031), .ZN(n5745) );
  NOR2_X1 U5621 ( .A1(n4889), .A2(n4976), .ZN(n4977) );
  NAND2_X1 U5622 ( .A1(n4978), .A2(n4889), .ZN(n5371) );
  NAND2_X1 U5623 ( .A1(n4978), .A2(n6930), .ZN(n4979) );
  NAND2_X1 U5624 ( .A1(n5371), .A2(n4979), .ZN(n4980) );
  NOR3_X1 U5625 ( .A1(n6980), .A2(n4981), .A3(n4980), .ZN(n4982) );
  OAI222_X1 U5626 ( .A1(n5741), .A2(n5451), .B1(n5150), .B2(n6889), .C1(n5745), 
        .C2(n4982), .ZN(U3462) );
  XNOR2_X1 U5627 ( .A(n5091), .B(n4889), .ZN(n4983) );
  INV_X1 U5628 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4986) );
  AOI22_X1 U5629 ( .A1(n5570), .A2(n5275), .B1(n7073), .B2(n5274), .ZN(n4985)
         );
  AOI22_X1 U5630 ( .A1(n5283), .A2(n7072), .B1(n7071), .B2(n5276), .ZN(n4984)
         );
  OAI211_X1 U5631 ( .C1(n5280), .C2(n4986), .A(n4985), .B(n4984), .ZN(U3141)
         );
  NOR2_X1 U5632 ( .A1(n7024), .A2(n5052), .ZN(n5289) );
  INV_X1 U5633 ( .A(n5289), .ZN(n4987) );
  INV_X1 U5634 ( .A(n5227), .ZN(n5003) );
  OR2_X1 U5635 ( .A1(n5228), .A2(n5003), .ZN(n5059) );
  AND2_X1 U5636 ( .A1(n5059), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U5637 ( .A1(n4993), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6993) );
  NAND2_X1 U5638 ( .A1(n5175), .A2(n6993), .ZN(n5220) );
  AOI211_X1 U5639 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4987), .A(n5053), .B(
        n5220), .ZN(n4992) );
  NOR2_X1 U5640 ( .A1(n4892), .A2(n4893), .ZN(n7022) );
  NOR2_X1 U5641 ( .A1(n7022), .A2(n7052), .ZN(n5223) );
  NOR2_X1 U5642 ( .A1(n5152), .A2(n4988), .ZN(n5097) );
  INV_X1 U5643 ( .A(n5097), .ZN(n4989) );
  NAND2_X1 U5644 ( .A1(n7040), .A2(n6990), .ZN(n4995) );
  NOR2_X1 U5645 ( .A1(n4990), .A2(n4890), .ZN(n7021) );
  NAND2_X1 U5646 ( .A1(n7021), .A2(n5746), .ZN(n4994) );
  OAI211_X1 U5647 ( .C1(n5127), .C2(n5223), .A(n4995), .B(n4994), .ZN(n4991)
         );
  INV_X1 U5648 ( .A(n7022), .ZN(n5230) );
  NAND2_X1 U5649 ( .A1(n5230), .A2(n6991), .ZN(n5225) );
  AND3_X1 U5650 ( .A1(n4992), .A2(n4991), .A3(n5225), .ZN(n5293) );
  INV_X1 U5651 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4998) );
  OR2_X1 U5652 ( .A1(n4993), .A2(n6906), .ZN(n5229) );
  OAI22_X1 U5653 ( .A1(n5230), .A2(n5553), .B1(n5059), .B2(n5229), .ZN(n5288)
         );
  AOI22_X1 U5654 ( .A1(n5574), .A2(n5288), .B1(n7107), .B2(n7176), .ZN(n4997)
         );
  AOI22_X1 U5655 ( .A1(n7185), .A2(n7108), .B1(n7106), .B2(n5289), .ZN(n4996)
         );
  OAI211_X1 U5656 ( .C1(n5293), .C2(n4998), .A(n4997), .B(n4996), .ZN(U3055)
         );
  INV_X1 U5657 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5001) );
  AOI22_X1 U5658 ( .A1(n5554), .A2(n5288), .B1(n7093), .B2(n7176), .ZN(n5000)
         );
  AOI22_X1 U5659 ( .A1(n7185), .A2(n7094), .B1(n7092), .B2(n5289), .ZN(n4999)
         );
  OAI211_X1 U5660 ( .C1(n5293), .C2(n5001), .A(n5000), .B(n4999), .ZN(U3054)
         );
  NOR2_X1 U5661 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5002), .ZN(n5282)
         );
  INV_X1 U5662 ( .A(n5282), .ZN(n5004) );
  NAND2_X1 U5663 ( .A1(n5003), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5010) );
  INV_X1 U5664 ( .A(n5010), .ZN(n6994) );
  NOR2_X1 U5665 ( .A1(n6994), .A2(n6906), .ZN(n6999) );
  AOI211_X1 U5666 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5004), .A(n6999), .B(
        n5220), .ZN(n5009) );
  NOR2_X1 U5667 ( .A1(n5007), .A2(n7052), .ZN(n5126) );
  INV_X1 U5668 ( .A(n7154), .ZN(n5006) );
  OAI211_X1 U5669 ( .C1(n5374), .C2(n5126), .A(n5006), .B(n5005), .ZN(n5008)
         );
  INV_X1 U5670 ( .A(n5007), .ZN(n5131) );
  NAND2_X1 U5671 ( .A1(n5131), .A2(n6991), .ZN(n5129) );
  AND3_X1 U5672 ( .A1(n5009), .A2(n5008), .A3(n5129), .ZN(n5287) );
  INV_X1 U5673 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5013) );
  INV_X1 U5674 ( .A(n5127), .ZN(n5379) );
  OAI22_X1 U5675 ( .A1(n5379), .A2(n5131), .B1(n5229), .B2(n5010), .ZN(n5281)
         );
  AOI22_X1 U5676 ( .A1(n5554), .A2(n5281), .B1(n7094), .B2(n7154), .ZN(n5012)
         );
  AOI22_X1 U5677 ( .A1(n5283), .A2(n7093), .B1(n7092), .B2(n5282), .ZN(n5011)
         );
  OAI211_X1 U5678 ( .C1(n5287), .C2(n5013), .A(n5012), .B(n5011), .ZN(U3134)
         );
  INV_X1 U5679 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5016) );
  AOI22_X1 U5680 ( .A1(n5584), .A2(n5281), .B1(n7183), .B2(n7154), .ZN(n5015)
         );
  AOI22_X1 U5681 ( .A1(n5283), .A2(n7186), .B1(n7182), .B2(n5282), .ZN(n5014)
         );
  OAI211_X1 U5682 ( .C1(n5287), .C2(n5016), .A(n5015), .B(n5014), .ZN(U3139)
         );
  INV_X1 U5683 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5019) );
  AOI22_X1 U5684 ( .A1(n5574), .A2(n5281), .B1(n7108), .B2(n7154), .ZN(n5018)
         );
  AOI22_X1 U5685 ( .A1(n5283), .A2(n7107), .B1(n7106), .B2(n5282), .ZN(n5017)
         );
  OAI211_X1 U5686 ( .C1(n5287), .C2(n5019), .A(n5018), .B(n5017), .ZN(U3135)
         );
  INV_X1 U5687 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5022) );
  AOI22_X1 U5688 ( .A1(n5584), .A2(n5288), .B1(n7186), .B2(n7176), .ZN(n5021)
         );
  AOI22_X1 U5689 ( .A1(n7185), .A2(n7183), .B1(n7182), .B2(n5289), .ZN(n5020)
         );
  OAI211_X1 U5690 ( .C1(n5293), .C2(n5022), .A(n5021), .B(n5020), .ZN(U3059)
         );
  INV_X1 U5691 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5025) );
  AOI22_X1 U5692 ( .A1(n5566), .A2(n5288), .B1(n7149), .B2(n7176), .ZN(n5024)
         );
  AOI22_X1 U5693 ( .A1(n7185), .A2(n7150), .B1(n7148), .B2(n5289), .ZN(n5023)
         );
  OAI211_X1 U5694 ( .C1(n5293), .C2(n5025), .A(n5024), .B(n5023), .ZN(U3058)
         );
  INV_X1 U5695 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5028) );
  AOI22_X1 U5696 ( .A1(n5566), .A2(n5281), .B1(n7150), .B2(n7154), .ZN(n5027)
         );
  AOI22_X1 U5697 ( .A1(n5283), .A2(n7149), .B1(n7148), .B2(n5282), .ZN(n5026)
         );
  OAI211_X1 U5698 ( .C1(n5287), .C2(n5028), .A(n5027), .B(n5026), .ZN(U3138)
         );
  INV_X1 U5699 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5031) );
  AOI22_X1 U5700 ( .A1(n5578), .A2(n5281), .B1(n7056), .B2(n7154), .ZN(n5030)
         );
  AOI22_X1 U5701 ( .A1(n7048), .A2(n5283), .B1(n7047), .B2(n5282), .ZN(n5029)
         );
  OAI211_X1 U5702 ( .C1(n5287), .C2(n5031), .A(n5030), .B(n5029), .ZN(U3132)
         );
  INV_X1 U5703 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5034) );
  AOI22_X1 U5704 ( .A1(n5578), .A2(n5288), .B1(n7048), .B2(n7176), .ZN(n5033)
         );
  AOI22_X1 U5705 ( .A1(n7185), .A2(n7056), .B1(n7047), .B2(n5289), .ZN(n5032)
         );
  OAI211_X1 U5706 ( .C1(n5293), .C2(n5034), .A(n5033), .B(n5032), .ZN(U3052)
         );
  INV_X1 U5707 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5037) );
  AOI22_X1 U5708 ( .A1(n5570), .A2(n5281), .B1(n7072), .B2(n7154), .ZN(n5036)
         );
  AOI22_X1 U5709 ( .A1(n5283), .A2(n7073), .B1(n7071), .B2(n5282), .ZN(n5035)
         );
  OAI211_X1 U5710 ( .C1(n5287), .C2(n5037), .A(n5036), .B(n5035), .ZN(U3133)
         );
  INV_X1 U5711 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5040) );
  AOI22_X1 U5712 ( .A1(n5570), .A2(n5288), .B1(n7073), .B2(n7176), .ZN(n5039)
         );
  AOI22_X1 U5713 ( .A1(n7185), .A2(n7072), .B1(n7071), .B2(n5289), .ZN(n5038)
         );
  OAI211_X1 U5714 ( .C1(n5293), .C2(n5040), .A(n5039), .B(n5038), .ZN(U3053)
         );
  NAND2_X1 U5715 ( .A1(n5044), .A2(n5043), .ZN(n5045) );
  AND2_X1 U5716 ( .A1(n5042), .A2(n5045), .ZN(n6752) );
  INV_X1 U5717 ( .A(n6752), .ZN(n5047) );
  OAI222_X1 U5718 ( .A1(n5047), .A2(n5976), .B1(n5975), .B2(n5046), .C1(n3422), 
        .C2(n3875), .ZN(U2886) );
  XNOR2_X1 U5719 ( .A(n5042), .B(n5085), .ZN(n6535) );
  INV_X1 U5720 ( .A(n6535), .ZN(n6766) );
  OAI21_X1 U5721 ( .B1(n6506), .B2(n5048), .A(n6493), .ZN(n6761) );
  INV_X1 U5722 ( .A(n6761), .ZN(n5049) );
  AOI22_X1 U5723 ( .A1(n6507), .A2(n5049), .B1(n6200), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n5050) );
  OAI21_X1 U5724 ( .B1(n6766), .B2(n5958), .A(n5050), .ZN(U2853) );
  INV_X1 U5725 ( .A(DATAI_6_), .ZN(n6247) );
  OAI222_X1 U5726 ( .A1(n5976), .A2(n6766), .B1(n3422), .B2(n4779), .C1(n6247), 
        .C2(n5975), .ZN(U2885) );
  NOR2_X1 U5727 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n7042) );
  INV_X1 U5728 ( .A(n7042), .ZN(n5051) );
  NOR2_X1 U5729 ( .A1(n5052), .A2(n5051), .ZN(n5259) );
  INV_X1 U5730 ( .A(n5259), .ZN(n5054) );
  NAND2_X1 U5731 ( .A1(n5175), .A2(n5229), .ZN(n7000) );
  AOI211_X1 U5732 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5054), .A(n5053), .B(
        n7000), .ZN(n5058) );
  NOR2_X1 U5733 ( .A1(n5170), .A2(n7052), .ZN(n5373) );
  NOR2_X1 U5734 ( .A1(n4978), .A2(n4888), .ZN(n5055) );
  NAND2_X1 U5735 ( .A1(n5183), .A2(n5746), .ZN(n5256) );
  OAI211_X1 U5736 ( .C1(n5373), .C2(n5127), .A(n5256), .B(n5255), .ZN(n5057)
         );
  INV_X1 U5737 ( .A(n5170), .ZN(n7007) );
  NAND2_X1 U5738 ( .A1(n7007), .A2(n6991), .ZN(n5056) );
  AND3_X1 U5739 ( .A1(n5058), .A2(n5057), .A3(n5056), .ZN(n5263) );
  INV_X1 U5740 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5063) );
  OAI22_X1 U5741 ( .A1(n5553), .A2(n7007), .B1(n6993), .B2(n5059), .ZN(n5258)
         );
  INV_X1 U5742 ( .A(n7073), .ZN(n5425) );
  INV_X1 U5743 ( .A(n7072), .ZN(n5423) );
  OAI22_X1 U5744 ( .A1(n5256), .A2(n5425), .B1(n5423), .B2(n5255), .ZN(n5060)
         );
  AOI21_X1 U5745 ( .B1(n5570), .B2(n5258), .A(n5060), .ZN(n5062) );
  NAND2_X1 U5746 ( .A1(n7071), .A2(n5259), .ZN(n5061) );
  OAI211_X1 U5747 ( .C1(n5263), .C2(n5063), .A(n5062), .B(n5061), .ZN(U3021)
         );
  INV_X1 U5748 ( .A(n7048), .ZN(n5411) );
  INV_X1 U5749 ( .A(n7056), .ZN(n5410) );
  OAI22_X1 U5750 ( .A1(n5256), .A2(n5411), .B1(n5410), .B2(n5255), .ZN(n5064)
         );
  AOI21_X1 U5751 ( .B1(n5578), .B2(n5258), .A(n5064), .ZN(n5066) );
  NAND2_X1 U5752 ( .A1(n7047), .A2(n5259), .ZN(n5065) );
  OAI211_X1 U5753 ( .C1(n5263), .C2(n5067), .A(n5066), .B(n5065), .ZN(U3020)
         );
  INV_X1 U5754 ( .A(n7186), .ZN(n5393) );
  INV_X1 U5755 ( .A(n7183), .ZN(n5392) );
  OAI22_X1 U5756 ( .A1(n5256), .A2(n5393), .B1(n5392), .B2(n5255), .ZN(n5068)
         );
  AOI21_X1 U5757 ( .B1(n5584), .B2(n5258), .A(n5068), .ZN(n5070) );
  NAND2_X1 U5758 ( .A1(n7182), .A2(n5259), .ZN(n5069) );
  OAI211_X1 U5759 ( .C1(n5263), .C2(n5071), .A(n5070), .B(n5069), .ZN(U3027)
         );
  INV_X1 U5760 ( .A(n7149), .ZN(n5387) );
  INV_X1 U5761 ( .A(n7150), .ZN(n5386) );
  OAI22_X1 U5762 ( .A1(n5256), .A2(n5387), .B1(n5386), .B2(n5255), .ZN(n5072)
         );
  AOI21_X1 U5763 ( .B1(n5566), .B2(n5258), .A(n5072), .ZN(n5074) );
  NAND2_X1 U5764 ( .A1(n7148), .A2(n5259), .ZN(n5073) );
  OAI211_X1 U5765 ( .C1(n5263), .C2(n5075), .A(n5074), .B(n5073), .ZN(U3026)
         );
  INV_X1 U5766 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5079) );
  INV_X1 U5767 ( .A(n7093), .ZN(n5405) );
  INV_X1 U5768 ( .A(n7094), .ZN(n5404) );
  OAI22_X1 U5769 ( .A1(n5256), .A2(n5405), .B1(n5404), .B2(n5255), .ZN(n5076)
         );
  AOI21_X1 U5770 ( .B1(n5554), .B2(n5258), .A(n5076), .ZN(n5078) );
  NAND2_X1 U5771 ( .A1(n7092), .A2(n5259), .ZN(n5077) );
  OAI211_X1 U5772 ( .C1(n5263), .C2(n5079), .A(n5078), .B(n5077), .ZN(U3022)
         );
  INV_X1 U5773 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5083) );
  INV_X1 U5774 ( .A(n7107), .ZN(n5399) );
  INV_X1 U5775 ( .A(n7108), .ZN(n5398) );
  OAI22_X1 U5776 ( .A1(n5256), .A2(n5399), .B1(n5398), .B2(n5255), .ZN(n5080)
         );
  AOI21_X1 U5777 ( .B1(n5574), .B2(n5258), .A(n5080), .ZN(n5082) );
  NAND2_X1 U5778 ( .A1(n7106), .A2(n5259), .ZN(n5081) );
  OAI211_X1 U5779 ( .C1(n5263), .C2(n5083), .A(n5082), .B(n5081), .ZN(U3023)
         );
  INV_X1 U5780 ( .A(n5085), .ZN(n5088) );
  INV_X1 U5781 ( .A(n5086), .ZN(n5087) );
  OAI21_X1 U5782 ( .B1(n5042), .B2(n5088), .A(n5087), .ZN(n5089) );
  AND2_X1 U5783 ( .A1(n5084), .A2(n5089), .ZN(n6779) );
  INV_X1 U5784 ( .A(n6779), .ZN(n5090) );
  INV_X1 U5785 ( .A(DATAI_7_), .ZN(n6342) );
  OAI222_X1 U5786 ( .A1(n5090), .A2(n5976), .B1(n5975), .B2(n6342), .C1(n3422), 
        .C2(n4774), .ZN(U2884) );
  INV_X1 U5787 ( .A(n5371), .ZN(n5092) );
  INV_X1 U5788 ( .A(n5091), .ZN(n5151) );
  AOI21_X1 U5789 ( .B1(n5092), .B2(n5151), .A(n7052), .ZN(n5099) );
  AND2_X1 U5790 ( .A1(n4892), .A2(n4893), .ZN(n5546) );
  AND2_X1 U5791 ( .A1(n5546), .A2(n5548), .ZN(n7003) );
  NAND3_X1 U5792 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6883), .ZN(n6998) );
  NOR2_X1 U5793 ( .A1(n7025), .A2(n6998), .ZN(n5164) );
  AOI21_X1 U5794 ( .B1(n7003), .B2(n5093), .A(n5164), .ZN(n5100) );
  INV_X1 U5795 ( .A(n6998), .ZN(n5094) );
  NOR2_X1 U5796 ( .A1(n7031), .A2(n5094), .ZN(n5095) );
  AOI211_X2 U5797 ( .C1(n5099), .C2(n5100), .A(n7050), .B(n5095), .ZN(n5169)
         );
  INV_X1 U5798 ( .A(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n5104) );
  NOR2_X1 U5799 ( .A1(n4988), .A2(n6990), .ZN(n5096) );
  NAND3_X1 U5800 ( .A1(n4978), .A2(n6990), .A3(n5097), .ZN(n5324) );
  OAI22_X1 U5801 ( .A1(n5162), .A2(n5410), .B1(n5411), .B2(n5324), .ZN(n5098)
         );
  AOI21_X1 U5802 ( .B1(n7047), .B2(n5164), .A(n5098), .ZN(n5103) );
  INV_X1 U5803 ( .A(n5099), .ZN(n5101) );
  OAI22_X1 U5804 ( .A1(n5101), .A2(n5100), .B1(n6998), .B2(n6906), .ZN(n5165)
         );
  NAND2_X1 U5805 ( .A1(n5165), .A2(n5578), .ZN(n5102) );
  OAI211_X1 U5806 ( .C1(n5169), .C2(n5104), .A(n5103), .B(n5102), .ZN(U3108)
         );
  INV_X1 U5807 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n5108) );
  OAI22_X1 U5808 ( .A1(n5162), .A2(n5386), .B1(n5387), .B2(n5324), .ZN(n5105)
         );
  AOI21_X1 U5809 ( .B1(n7148), .B2(n5164), .A(n5105), .ZN(n5107) );
  NAND2_X1 U5810 ( .A1(n5165), .A2(n5566), .ZN(n5106) );
  OAI211_X1 U5811 ( .C1(n5169), .C2(n5108), .A(n5107), .B(n5106), .ZN(U3114)
         );
  INV_X1 U5812 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n5112) );
  OAI22_X1 U5813 ( .A1(n5162), .A2(n5398), .B1(n5399), .B2(n5324), .ZN(n5109)
         );
  AOI21_X1 U5814 ( .B1(n7106), .B2(n5164), .A(n5109), .ZN(n5111) );
  NAND2_X1 U5815 ( .A1(n5165), .A2(n5574), .ZN(n5110) );
  OAI211_X1 U5816 ( .C1(n5169), .C2(n5112), .A(n5111), .B(n5110), .ZN(U3111)
         );
  INV_X1 U5817 ( .A(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n5116) );
  OAI22_X1 U5818 ( .A1(n5162), .A2(n5392), .B1(n5393), .B2(n5324), .ZN(n5113)
         );
  AOI21_X1 U5819 ( .B1(n7182), .B2(n5164), .A(n5113), .ZN(n5115) );
  NAND2_X1 U5820 ( .A1(n5165), .A2(n5584), .ZN(n5114) );
  OAI211_X1 U5821 ( .C1(n5169), .C2(n5116), .A(n5115), .B(n5114), .ZN(U3115)
         );
  INV_X1 U5822 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n5120) );
  OAI22_X1 U5823 ( .A1(n5162), .A2(n5404), .B1(n5405), .B2(n5324), .ZN(n5117)
         );
  AOI21_X1 U5824 ( .B1(n7092), .B2(n5164), .A(n5117), .ZN(n5119) );
  NAND2_X1 U5825 ( .A1(n5165), .A2(n5554), .ZN(n5118) );
  OAI211_X1 U5826 ( .C1(n5169), .C2(n5120), .A(n5119), .B(n5118), .ZN(U3110)
         );
  INV_X1 U5827 ( .A(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n5124) );
  OAI22_X1 U5828 ( .A1(n5162), .A2(n5423), .B1(n5425), .B2(n5324), .ZN(n5121)
         );
  AOI21_X1 U5829 ( .B1(n7071), .B2(n5164), .A(n5121), .ZN(n5123) );
  NAND2_X1 U5830 ( .A1(n5165), .A2(n5570), .ZN(n5122) );
  OAI211_X1 U5831 ( .C1(n5169), .C2(n5124), .A(n5123), .B(n5122), .ZN(U3109)
         );
  OR2_X1 U5832 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5125), .ZN(n5322)
         );
  OR2_X1 U5833 ( .A1(n5227), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5552)
         );
  AND2_X1 U5834 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5552), .ZN(n5550) );
  AOI211_X1 U5835 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5322), .A(n5550), .B(
        n5220), .ZN(n5130) );
  NAND2_X1 U5836 ( .A1(n7021), .A2(n6990), .ZN(n7036) );
  OAI211_X1 U5837 ( .C1(n5127), .C2(n5126), .A(n5317), .B(n7036), .ZN(n5128)
         );
  NAND3_X1 U5838 ( .A1(n5130), .A2(n5129), .A3(n5128), .ZN(n5316) );
  NAND2_X1 U5839 ( .A1(n5316), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5134) );
  OAI22_X1 U5840 ( .A1(n5553), .A2(n5131), .B1(n5552), .B2(n5229), .ZN(n5319)
         );
  OAI22_X1 U5841 ( .A1(n5317), .A2(n5399), .B1(n7036), .B2(n5398), .ZN(n5132)
         );
  AOI21_X1 U5842 ( .B1(n5574), .B2(n5319), .A(n5132), .ZN(n5133) );
  OAI211_X1 U5843 ( .C1(n5322), .C2(n5403), .A(n5134), .B(n5133), .ZN(U3071)
         );
  NAND2_X1 U5844 ( .A1(n5316), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5137) );
  OAI22_X1 U5845 ( .A1(n5317), .A2(n5387), .B1(n7036), .B2(n5386), .ZN(n5135)
         );
  AOI21_X1 U5846 ( .B1(n5566), .B2(n5319), .A(n5135), .ZN(n5136) );
  OAI211_X1 U5847 ( .C1(n5322), .C2(n5391), .A(n5137), .B(n5136), .ZN(U3074)
         );
  NAND2_X1 U5848 ( .A1(n5316), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5140) );
  OAI22_X1 U5849 ( .A1(n5317), .A2(n5425), .B1(n7036), .B2(n5423), .ZN(n5138)
         );
  AOI21_X1 U5850 ( .B1(n5570), .B2(n5319), .A(n5138), .ZN(n5139) );
  OAI211_X1 U5851 ( .C1(n5322), .C2(n5430), .A(n5140), .B(n5139), .ZN(U3069)
         );
  NAND2_X1 U5852 ( .A1(n5316), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5143) );
  OAI22_X1 U5853 ( .A1(n5317), .A2(n5411), .B1(n7036), .B2(n5410), .ZN(n5141)
         );
  AOI21_X1 U5854 ( .B1(n5578), .B2(n5319), .A(n5141), .ZN(n5142) );
  OAI211_X1 U5855 ( .C1(n5415), .C2(n5322), .A(n5143), .B(n5142), .ZN(U3068)
         );
  NAND2_X1 U5856 ( .A1(n5316), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5146) );
  OAI22_X1 U5857 ( .A1(n5317), .A2(n5393), .B1(n7036), .B2(n5392), .ZN(n5144)
         );
  AOI21_X1 U5858 ( .B1(n5584), .B2(n5319), .A(n5144), .ZN(n5145) );
  OAI211_X1 U5859 ( .C1(n5322), .C2(n5397), .A(n5146), .B(n5145), .ZN(U3075)
         );
  NAND2_X1 U5860 ( .A1(n5316), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5149) );
  OAI22_X1 U5861 ( .A1(n5317), .A2(n5405), .B1(n7036), .B2(n5404), .ZN(n5147)
         );
  AOI21_X1 U5862 ( .B1(n5554), .B2(n5319), .A(n5147), .ZN(n5148) );
  OAI211_X1 U5863 ( .C1(n5322), .C2(n5409), .A(n5149), .B(n5148), .ZN(U3070)
         );
  INV_X1 U5864 ( .A(n5150), .ZN(n6197) );
  AOI211_X1 U5865 ( .C1(n5152), .C2(n6930), .A(n5151), .B(n5745), .ZN(n5153)
         );
  AOI21_X1 U5866 ( .B1(n6197), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n5153), 
        .ZN(n5154) );
  OAI21_X1 U5867 ( .B1(n5357), .B2(n5741), .A(n5154), .ZN(U3464) );
  INV_X1 U5868 ( .A(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n5159) );
  NOR2_X2 U5869 ( .A1(n5161), .A2(n5155), .ZN(n7134) );
  AND2_X1 U5870 ( .A1(n6561), .A2(DATAI_29_), .ZN(n7136) );
  INV_X1 U5871 ( .A(n7136), .ZN(n5380) );
  AND2_X1 U5872 ( .A1(n6561), .A2(DATAI_21_), .ZN(n7135) );
  INV_X1 U5873 ( .A(n7135), .ZN(n5381) );
  OAI22_X1 U5874 ( .A1(n5162), .A2(n5380), .B1(n5381), .B2(n5324), .ZN(n5156)
         );
  AOI21_X1 U5875 ( .B1(n7134), .B2(n5164), .A(n5156), .ZN(n5158) );
  NAND2_X1 U5876 ( .A1(DATAI_5_), .A2(n5175), .ZN(n7139) );
  NAND2_X1 U5877 ( .A1(n5165), .A2(n5562), .ZN(n5157) );
  OAI211_X1 U5878 ( .C1(n5169), .C2(n5159), .A(n5158), .B(n5157), .ZN(U3113)
         );
  INV_X1 U5879 ( .A(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n5168) );
  NOR2_X2 U5880 ( .A1(n5161), .A2(n5160), .ZN(n7120) );
  AND2_X1 U5881 ( .A1(n6561), .A2(DATAI_28_), .ZN(n7122) );
  INV_X1 U5882 ( .A(n7122), .ZN(n5416) );
  AND2_X1 U5883 ( .A1(n6561), .A2(DATAI_20_), .ZN(n7121) );
  INV_X1 U5884 ( .A(n7121), .ZN(n5417) );
  OAI22_X1 U5885 ( .A1(n5162), .A2(n5416), .B1(n5417), .B2(n5324), .ZN(n5163)
         );
  AOI21_X1 U5886 ( .B1(n7120), .B2(n5164), .A(n5163), .ZN(n5167) );
  NAND2_X1 U5887 ( .A1(DATAI_4_), .A2(n5175), .ZN(n7125) );
  NAND2_X1 U5888 ( .A1(n5165), .A2(n5558), .ZN(n5166) );
  OAI211_X1 U5889 ( .C1(n5169), .C2(n5168), .A(n5167), .B(n5166), .ZN(U3112)
         );
  INV_X1 U5890 ( .A(n5183), .ZN(n5171) );
  NAND2_X1 U5891 ( .A1(n7023), .A2(n5170), .ZN(n5179) );
  OAI21_X1 U5892 ( .B1(n5171), .B2(n6930), .A(n5179), .ZN(n5174) );
  NAND3_X1 U5893 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7042), .A3(n5172), .ZN(
        n5180) );
  NAND3_X1 U5894 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7042), .A3(n5172), .ZN(n5178) );
  OAI21_X1 U5895 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5180), .A(n5178), .ZN(
        n5173) );
  AOI21_X1 U5896 ( .B1(n5174), .B2(n7031), .A(n5173), .ZN(n5177) );
  INV_X1 U5897 ( .A(n5175), .ZN(n5176) );
  INV_X1 U5898 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5187) );
  INV_X1 U5899 ( .A(n5178), .ZN(n5216) );
  AOI21_X1 U5900 ( .B1(n5179), .B2(n5178), .A(n7052), .ZN(n5182) );
  INV_X1 U5901 ( .A(n5180), .ZN(n5181) );
  NOR2_X1 U5902 ( .A1(n5182), .A2(n5181), .ZN(n5214) );
  AOI22_X1 U5903 ( .A1(n5212), .A2(n7183), .B1(n5582), .B2(n7186), .ZN(n5184)
         );
  OAI21_X1 U5904 ( .B1(n7190), .B2(n5214), .A(n5184), .ZN(n5185) );
  AOI21_X1 U5905 ( .B1(n7182), .B2(n5216), .A(n5185), .ZN(n5186) );
  OAI21_X1 U5906 ( .B1(n5219), .B2(n5187), .A(n5186), .ZN(U3035) );
  INV_X1 U5907 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n5191) );
  AOI22_X1 U5908 ( .A1(n5212), .A2(n7072), .B1(n5582), .B2(n7073), .ZN(n5188)
         );
  OAI21_X1 U5909 ( .B1(n7076), .B2(n5214), .A(n5188), .ZN(n5189) );
  AOI21_X1 U5910 ( .B1(n7071), .B2(n5216), .A(n5189), .ZN(n5190) );
  OAI21_X1 U5911 ( .B1(n5219), .B2(n5191), .A(n5190), .ZN(U3029) );
  INV_X1 U5912 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n5195) );
  AOI22_X1 U5913 ( .A1(n5212), .A2(n7056), .B1(n5582), .B2(n7048), .ZN(n5192)
         );
  OAI21_X1 U5914 ( .B1(n7059), .B2(n5214), .A(n5192), .ZN(n5193) );
  AOI21_X1 U5915 ( .B1(n7047), .B2(n5216), .A(n5193), .ZN(n5194) );
  OAI21_X1 U5916 ( .B1(n5219), .B2(n5195), .A(n5194), .ZN(U3028) );
  INV_X1 U5917 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n5199) );
  AOI22_X1 U5918 ( .A1(n5212), .A2(n7108), .B1(n5582), .B2(n7107), .ZN(n5196)
         );
  OAI21_X1 U5919 ( .B1(n7111), .B2(n5214), .A(n5196), .ZN(n5197) );
  AOI21_X1 U5920 ( .B1(n7106), .B2(n5216), .A(n5197), .ZN(n5198) );
  OAI21_X1 U5921 ( .B1(n5219), .B2(n5199), .A(n5198), .ZN(U3031) );
  INV_X1 U5922 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n5203) );
  AOI22_X1 U5923 ( .A1(n5212), .A2(n7094), .B1(n5582), .B2(n7093), .ZN(n5200)
         );
  OAI21_X1 U5924 ( .B1(n7097), .B2(n5214), .A(n5200), .ZN(n5201) );
  AOI21_X1 U5925 ( .B1(n7092), .B2(n5216), .A(n5201), .ZN(n5202) );
  OAI21_X1 U5926 ( .B1(n5219), .B2(n5203), .A(n5202), .ZN(U3030) );
  INV_X1 U5927 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5207) );
  AOI22_X1 U5928 ( .A1(n5212), .A2(n7150), .B1(n5582), .B2(n7149), .ZN(n5204)
         );
  OAI21_X1 U5929 ( .B1(n7153), .B2(n5214), .A(n5204), .ZN(n5205) );
  AOI21_X1 U5930 ( .B1(n7148), .B2(n5216), .A(n5205), .ZN(n5206) );
  OAI21_X1 U5931 ( .B1(n5219), .B2(n5207), .A(n5206), .ZN(U3034) );
  INV_X1 U5932 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5211) );
  AOI22_X1 U5933 ( .A1(n5212), .A2(n7136), .B1(n5582), .B2(n7135), .ZN(n5208)
         );
  OAI21_X1 U5934 ( .B1(n7139), .B2(n5214), .A(n5208), .ZN(n5209) );
  AOI21_X1 U5935 ( .B1(n7134), .B2(n5216), .A(n5209), .ZN(n5210) );
  OAI21_X1 U5936 ( .B1(n5219), .B2(n5211), .A(n5210), .ZN(U3033) );
  INV_X1 U5937 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n5218) );
  AOI22_X1 U5938 ( .A1(n5212), .A2(n7122), .B1(n5582), .B2(n7121), .ZN(n5213)
         );
  OAI21_X1 U5939 ( .B1(n7125), .B2(n5214), .A(n5213), .ZN(n5215) );
  AOI21_X1 U5940 ( .B1(n7120), .B2(n5216), .A(n5215), .ZN(n5217) );
  OAI21_X1 U5941 ( .B1(n5219), .B2(n5218), .A(n5217), .ZN(U3032) );
  NOR3_X1 U5942 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6883), .A3(n6889), 
        .ZN(n6987) );
  INV_X1 U5943 ( .A(n6987), .ZN(n6981) );
  OR2_X1 U5944 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6981), .ZN(n5330)
         );
  AOI21_X1 U5945 ( .B1(n5228), .B2(n5227), .A(n6906), .ZN(n5370) );
  AOI211_X1 U5946 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5330), .A(n5370), .B(
        n5220), .ZN(n5226) );
  INV_X1 U5947 ( .A(n5221), .ZN(n5222) );
  OAI211_X1 U5948 ( .C1(n5374), .C2(n5223), .A(n5325), .B(n5324), .ZN(n5224)
         );
  NAND3_X1 U5949 ( .A1(n5226), .A2(n5225), .A3(n5224), .ZN(n5323) );
  NAND2_X1 U5950 ( .A1(n5323), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5233)
         );
  NAND2_X1 U5951 ( .A1(n5228), .A2(n5227), .ZN(n5378) );
  OAI22_X1 U5952 ( .A1(n5379), .A2(n5230), .B1(n5378), .B2(n5229), .ZN(n5327)
         );
  OAI22_X1 U5953 ( .A1(n5325), .A2(n5425), .B1(n5423), .B2(n5324), .ZN(n5231)
         );
  AOI21_X1 U5954 ( .B1(n5570), .B2(n5327), .A(n5231), .ZN(n5232) );
  OAI211_X1 U5955 ( .C1(n5330), .C2(n5430), .A(n5233), .B(n5232), .ZN(U3117)
         );
  NAND2_X1 U5956 ( .A1(n5323), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5236)
         );
  OAI22_X1 U5957 ( .A1(n5325), .A2(n5387), .B1(n5386), .B2(n5324), .ZN(n5234)
         );
  AOI21_X1 U5958 ( .B1(n5566), .B2(n5327), .A(n5234), .ZN(n5235) );
  OAI211_X1 U5959 ( .C1(n5330), .C2(n5391), .A(n5236), .B(n5235), .ZN(U3122)
         );
  NAND2_X1 U5960 ( .A1(n5323), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5239)
         );
  OAI22_X1 U5961 ( .A1(n5325), .A2(n5411), .B1(n5410), .B2(n5324), .ZN(n5237)
         );
  AOI21_X1 U5962 ( .B1(n5578), .B2(n5327), .A(n5237), .ZN(n5238) );
  OAI211_X1 U5963 ( .C1(n5415), .C2(n5330), .A(n5239), .B(n5238), .ZN(U3116)
         );
  NAND2_X1 U5964 ( .A1(n5323), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5242)
         );
  OAI22_X1 U5965 ( .A1(n5325), .A2(n5405), .B1(n5404), .B2(n5324), .ZN(n5240)
         );
  AOI21_X1 U5966 ( .B1(n5554), .B2(n5327), .A(n5240), .ZN(n5241) );
  OAI211_X1 U5967 ( .C1(n5330), .C2(n5409), .A(n5242), .B(n5241), .ZN(U3118)
         );
  NAND2_X1 U5968 ( .A1(n5323), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5245)
         );
  OAI22_X1 U5969 ( .A1(n5325), .A2(n5399), .B1(n5398), .B2(n5324), .ZN(n5243)
         );
  AOI21_X1 U5970 ( .B1(n5574), .B2(n5327), .A(n5243), .ZN(n5244) );
  OAI211_X1 U5971 ( .C1(n5330), .C2(n5403), .A(n5245), .B(n5244), .ZN(U3119)
         );
  NAND2_X1 U5972 ( .A1(n5323), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5248)
         );
  OAI22_X1 U5973 ( .A1(n5325), .A2(n5393), .B1(n5392), .B2(n5324), .ZN(n5246)
         );
  AOI21_X1 U5974 ( .B1(n5584), .B2(n5327), .A(n5246), .ZN(n5247) );
  OAI211_X1 U5975 ( .C1(n5330), .C2(n5397), .A(n5248), .B(n5247), .ZN(U3123)
         );
  AOI21_X1 U5976 ( .B1(n5250), .B2(n5084), .A(n5249), .ZN(n5491) );
  INV_X1 U5977 ( .A(n5491), .ZN(n5522) );
  INV_X1 U5978 ( .A(DATAI_8_), .ZN(n6341) );
  OAI222_X1 U5979 ( .A1(n5522), .A2(n5976), .B1(n5975), .B2(n6341), .C1(n3422), 
        .C2(n4791), .ZN(U2883) );
  OAI22_X1 U5980 ( .A1(n5256), .A2(n5381), .B1(n5380), .B2(n5255), .ZN(n5251)
         );
  AOI21_X1 U5981 ( .B1(n5562), .B2(n5258), .A(n5251), .ZN(n5253) );
  NAND2_X1 U5982 ( .A1(n7134), .A2(n5259), .ZN(n5252) );
  OAI211_X1 U5983 ( .C1(n5263), .C2(n5254), .A(n5253), .B(n5252), .ZN(U3025)
         );
  OAI22_X1 U5984 ( .A1(n5256), .A2(n5417), .B1(n5416), .B2(n5255), .ZN(n5257)
         );
  AOI21_X1 U5985 ( .B1(n5558), .B2(n5258), .A(n5257), .ZN(n5261) );
  NAND2_X1 U5986 ( .A1(n7120), .A2(n5259), .ZN(n5260) );
  OAI211_X1 U5987 ( .C1(n5263), .C2(n5262), .A(n5261), .B(n5260), .ZN(U3024)
         );
  AOI21_X1 U5988 ( .B1(n5264), .B2(n6495), .A(n5445), .ZN(n5340) );
  INV_X1 U5989 ( .A(n5340), .ZN(n5519) );
  INV_X1 U5990 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5514) );
  OAI222_X1 U5991 ( .A1(n5519), .A2(n5956), .B1(n6510), .B2(n5514), .C1(n5958), 
        .C2(n5522), .ZN(U2851) );
  INV_X1 U5992 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5267) );
  AOI22_X1 U5993 ( .A1(n5558), .A2(n5281), .B1(n7122), .B2(n7154), .ZN(n5266)
         );
  AOI22_X1 U5994 ( .A1(n5283), .A2(n7121), .B1(n7120), .B2(n5282), .ZN(n5265)
         );
  OAI211_X1 U5995 ( .C1(n5287), .C2(n5267), .A(n5266), .B(n5265), .ZN(U3136)
         );
  INV_X1 U5996 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5270) );
  AOI22_X1 U5997 ( .A1(n5562), .A2(n5275), .B1(n7135), .B2(n5274), .ZN(n5269)
         );
  AOI22_X1 U5998 ( .A1(n5283), .A2(n7136), .B1(n7134), .B2(n5276), .ZN(n5268)
         );
  OAI211_X1 U5999 ( .C1(n5280), .C2(n5270), .A(n5269), .B(n5268), .ZN(U3145)
         );
  INV_X1 U6000 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5273) );
  AOI22_X1 U6001 ( .A1(n5562), .A2(n5288), .B1(n7135), .B2(n7176), .ZN(n5272)
         );
  AOI22_X1 U6002 ( .A1(n7185), .A2(n7136), .B1(n7134), .B2(n5289), .ZN(n5271)
         );
  OAI211_X1 U6003 ( .C1(n5293), .C2(n5273), .A(n5272), .B(n5271), .ZN(U3057)
         );
  INV_X1 U6004 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5279) );
  AOI22_X1 U6005 ( .A1(n5558), .A2(n5275), .B1(n7121), .B2(n5274), .ZN(n5278)
         );
  AOI22_X1 U6006 ( .A1(n5283), .A2(n7122), .B1(n7120), .B2(n5276), .ZN(n5277)
         );
  OAI211_X1 U6007 ( .C1(n5280), .C2(n5279), .A(n5278), .B(n5277), .ZN(U3144)
         );
  INV_X1 U6008 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5286) );
  AOI22_X1 U6009 ( .A1(n5562), .A2(n5281), .B1(n7136), .B2(n7154), .ZN(n5285)
         );
  AOI22_X1 U6010 ( .A1(n5283), .A2(n7135), .B1(n7134), .B2(n5282), .ZN(n5284)
         );
  OAI211_X1 U6011 ( .C1(n5287), .C2(n5286), .A(n5285), .B(n5284), .ZN(U3137)
         );
  INV_X1 U6012 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5292) );
  AOI22_X1 U6013 ( .A1(n5558), .A2(n5288), .B1(n7121), .B2(n7176), .ZN(n5291)
         );
  AOI22_X1 U6014 ( .A1(n7185), .A2(n7122), .B1(n7120), .B2(n5289), .ZN(n5290)
         );
  OAI211_X1 U6015 ( .C1(n5293), .C2(n5292), .A(n5291), .B(n5290), .ZN(U3056)
         );
  AOI22_X1 U6016 ( .A1(n6585), .A2(UWORD_REG_14__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n5294) );
  OAI21_X1 U6017 ( .B1(n4766), .B2(n5301), .A(n5294), .ZN(U2893) );
  INV_X1 U6018 ( .A(EAX_REG_16__SCAN_IN), .ZN(n5296) );
  AOI22_X1 U6019 ( .A1(n6585), .A2(UWORD_REG_0__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5295) );
  OAI21_X1 U6020 ( .B1(n5296), .B2(n5301), .A(n5295), .ZN(U2907) );
  INV_X1 U6021 ( .A(EAX_REG_19__SCAN_IN), .ZN(n5298) );
  AOI22_X1 U6022 ( .A1(n6585), .A2(UWORD_REG_3__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n5297) );
  OAI21_X1 U6023 ( .B1(n5298), .B2(n5301), .A(n5297), .ZN(U2904) );
  AOI22_X1 U6024 ( .A1(n6585), .A2(UWORD_REG_1__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n5299) );
  OAI21_X1 U6025 ( .B1(n4788), .B2(n5301), .A(n5299), .ZN(U2906) );
  AOI22_X1 U6026 ( .A1(n6585), .A2(UWORD_REG_2__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5300) );
  OAI21_X1 U6027 ( .B1(n6961), .B2(n5301), .A(n5300), .ZN(U2905) );
  INV_X1 U6028 ( .A(n7120), .ZN(n5421) );
  AOI22_X1 U6029 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n5311), .B1(n5558), 
        .B2(n5310), .ZN(n5303) );
  AOI22_X1 U6030 ( .A1(n5312), .A2(n7122), .B1(n5372), .B2(n7121), .ZN(n5302)
         );
  OAI211_X1 U6031 ( .C1(n5315), .C2(n5421), .A(n5303), .B(n5302), .ZN(U3080)
         );
  INV_X1 U6032 ( .A(n7134), .ZN(n5385) );
  NAND2_X1 U6033 ( .A1(n5323), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5306)
         );
  OAI22_X1 U6034 ( .A1(n5325), .A2(n5381), .B1(n5380), .B2(n5324), .ZN(n5304)
         );
  AOI21_X1 U6035 ( .B1(n5562), .B2(n5327), .A(n5304), .ZN(n5305) );
  OAI211_X1 U6036 ( .C1(n5330), .C2(n5385), .A(n5306), .B(n5305), .ZN(U3121)
         );
  NAND2_X1 U6037 ( .A1(n5316), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5309) );
  OAI22_X1 U6038 ( .A1(n5317), .A2(n5381), .B1(n7036), .B2(n5380), .ZN(n5307)
         );
  AOI21_X1 U6039 ( .B1(n5562), .B2(n5319), .A(n5307), .ZN(n5308) );
  OAI211_X1 U6040 ( .C1(n5322), .C2(n5385), .A(n5309), .B(n5308), .ZN(U3073)
         );
  AOI22_X1 U6041 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n5311), .B1(n5562), 
        .B2(n5310), .ZN(n5314) );
  AOI22_X1 U6042 ( .A1(n5312), .A2(n7136), .B1(n5372), .B2(n7135), .ZN(n5313)
         );
  OAI211_X1 U6043 ( .C1(n5315), .C2(n5385), .A(n5314), .B(n5313), .ZN(U3081)
         );
  NAND2_X1 U6044 ( .A1(n5316), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5321) );
  OAI22_X1 U6045 ( .A1(n5317), .A2(n5417), .B1(n7036), .B2(n5416), .ZN(n5318)
         );
  AOI21_X1 U6046 ( .B1(n5558), .B2(n5319), .A(n5318), .ZN(n5320) );
  OAI211_X1 U6047 ( .C1(n5322), .C2(n5421), .A(n5321), .B(n5320), .ZN(U3072)
         );
  NAND2_X1 U6048 ( .A1(n5323), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5329)
         );
  OAI22_X1 U6049 ( .A1(n5325), .A2(n5417), .B1(n5416), .B2(n5324), .ZN(n5326)
         );
  AOI21_X1 U6050 ( .B1(n5558), .B2(n5327), .A(n5326), .ZN(n5328) );
  OAI211_X1 U6051 ( .C1(n5330), .C2(n5421), .A(n5329), .B(n5328), .ZN(U3120)
         );
  OAI21_X1 U6052 ( .B1(n3435), .B2(n5332), .A(n5331), .ZN(n5493) );
  AND2_X1 U6053 ( .A1(n6789), .A2(REIP_REG_8__SCAN_IN), .ZN(n5488) );
  INV_X1 U6054 ( .A(n5334), .ZN(n5336) );
  NOR2_X1 U6055 ( .A1(n5336), .A2(n6639), .ZN(n6668) );
  OAI21_X1 U6056 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6668), .ZN(n5338) );
  INV_X1 U6057 ( .A(n6660), .ZN(n5335) );
  OAI22_X1 U6058 ( .A1(n5336), .A2(n6630), .B1(n6694), .B2(n5335), .ZN(n6672)
         );
  OAI22_X1 U6059 ( .A1(n6673), .A2(n5338), .B1(n5337), .B2(n6672), .ZN(n5339)
         );
  AOI211_X1 U6060 ( .C1(n6721), .C2(n5340), .A(n5488), .B(n5339), .ZN(n5341)
         );
  OAI21_X1 U6061 ( .B1(n6702), .B2(n5493), .A(n5341), .ZN(U3010) );
  INV_X1 U6062 ( .A(n6583), .ZN(n5350) );
  AND2_X1 U6063 ( .A1(n3421), .A2(n5344), .ZN(n6908) );
  NOR3_X1 U6064 ( .A1(n6923), .A2(n6916), .A3(n6925), .ZN(n6919) );
  NOR2_X1 U6065 ( .A1(n6908), .A2(n6919), .ZN(n5346) );
  NAND2_X1 U6066 ( .A1(n5346), .A2(n6821), .ZN(n5347) );
  NOR2_X1 U6067 ( .A1(n5353), .A2(n5348), .ZN(n5349) );
  OAI21_X1 U6068 ( .B1(n5350), .B2(n3673), .A(n6827), .ZN(n6751) );
  INV_X1 U6069 ( .A(n6751), .ZN(n5476) );
  NAND2_X1 U6070 ( .A1(n6583), .A2(EBX_REG_31__SCAN_IN), .ZN(n5804) );
  INV_X1 U6071 ( .A(n5804), .ZN(n5352) );
  NOR2_X1 U6072 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5361) );
  NOR2_X1 U6073 ( .A1(n4359), .A2(n5361), .ZN(n5351) );
  NAND2_X1 U6074 ( .A1(n6583), .A2(n5826), .ZN(n6731) );
  AOI22_X1 U6075 ( .A1(n6856), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n5658), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5356) );
  AND2_X1 U6076 ( .A1(n5353), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5354) );
  INV_X1 U6077 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U6078 ( .A1(n6861), .A2(n5527), .ZN(n5355) );
  OAI211_X1 U6079 ( .C1(n6731), .C2(n5357), .A(n5356), .B(n5355), .ZN(n5367)
         );
  NAND2_X1 U6080 ( .A1(n5827), .A2(n5361), .ZN(n6905) );
  NAND2_X1 U6081 ( .A1(n6581), .A2(n6905), .ZN(n5803) );
  INV_X1 U6082 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5918) );
  INV_X1 U6083 ( .A(n5361), .ZN(n5358) );
  NAND3_X1 U6084 ( .A1(n3643), .A2(n5918), .A3(n5358), .ZN(n5359) );
  NAND2_X1 U6085 ( .A1(n5803), .A2(n5359), .ZN(n5360) );
  INV_X1 U6086 ( .A(EBX_REG_1__SCAN_IN), .ZN(n5365) );
  AND2_X1 U6087 ( .A1(n3643), .A2(n5361), .ZN(n5362) );
  AND2_X1 U6088 ( .A1(n5363), .A2(n5362), .ZN(n5364) );
  OAI22_X1 U6089 ( .A1(n6796), .A2(n5365), .B1(REIP_REG_1__SCAN_IN), .B2(n6802), .ZN(n5366) );
  AOI211_X1 U6090 ( .C1(n6864), .C2(n5368), .A(n5367), .B(n5366), .ZN(n5369)
         );
  OAI21_X1 U6091 ( .B1(n5476), .B2(n5525), .A(n5369), .ZN(U2826) );
  NOR3_X1 U6092 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6889), .ZN(n7012) );
  INV_X1 U6093 ( .A(n7012), .ZN(n7015) );
  OR2_X1 U6094 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7015), .ZN(n5431)
         );
  AOI211_X1 U6095 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5431), .A(n5370), .B(
        n7000), .ZN(n5377) );
  NAND2_X1 U6096 ( .A1(n5374), .A2(n6930), .ZN(n5376) );
  NOR2_X1 U6097 ( .A1(n5371), .A2(n4890), .ZN(n7011) );
  NAND2_X1 U6098 ( .A1(n7011), .A2(n5746), .ZN(n7013) );
  OAI211_X1 U6099 ( .C1(n5374), .C2(n5373), .A(n7013), .B(n5424), .ZN(n5375)
         );
  NAND3_X1 U6100 ( .A1(n5377), .A2(n5376), .A3(n5375), .ZN(n5422) );
  NAND2_X1 U6101 ( .A1(n5422), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5384) );
  OAI22_X1 U6102 ( .A1(n5379), .A2(n7007), .B1(n6993), .B2(n5378), .ZN(n5427)
         );
  OAI22_X1 U6103 ( .A1(n7013), .A2(n5381), .B1(n5424), .B2(n5380), .ZN(n5382)
         );
  AOI21_X1 U6104 ( .B1(n5562), .B2(n5427), .A(n5382), .ZN(n5383) );
  OAI211_X1 U6105 ( .C1(n5431), .C2(n5385), .A(n5384), .B(n5383), .ZN(U3089)
         );
  NAND2_X1 U6106 ( .A1(n5422), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5390) );
  OAI22_X1 U6107 ( .A1(n7013), .A2(n5387), .B1(n5424), .B2(n5386), .ZN(n5388)
         );
  AOI21_X1 U6108 ( .B1(n5566), .B2(n5427), .A(n5388), .ZN(n5389) );
  OAI211_X1 U6109 ( .C1(n5431), .C2(n5391), .A(n5390), .B(n5389), .ZN(U3090)
         );
  NAND2_X1 U6110 ( .A1(n5422), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5396) );
  OAI22_X1 U6111 ( .A1(n7013), .A2(n5393), .B1(n5424), .B2(n5392), .ZN(n5394)
         );
  AOI21_X1 U6112 ( .B1(n5584), .B2(n5427), .A(n5394), .ZN(n5395) );
  OAI211_X1 U6113 ( .C1(n5431), .C2(n5397), .A(n5396), .B(n5395), .ZN(U3091)
         );
  NAND2_X1 U6114 ( .A1(n5422), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5402) );
  OAI22_X1 U6115 ( .A1(n7013), .A2(n5399), .B1(n5424), .B2(n5398), .ZN(n5400)
         );
  AOI21_X1 U6116 ( .B1(n5574), .B2(n5427), .A(n5400), .ZN(n5401) );
  OAI211_X1 U6117 ( .C1(n5431), .C2(n5403), .A(n5402), .B(n5401), .ZN(U3087)
         );
  NAND2_X1 U6118 ( .A1(n5422), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5408) );
  OAI22_X1 U6119 ( .A1(n7013), .A2(n5405), .B1(n5424), .B2(n5404), .ZN(n5406)
         );
  AOI21_X1 U6120 ( .B1(n5554), .B2(n5427), .A(n5406), .ZN(n5407) );
  OAI211_X1 U6121 ( .C1(n5431), .C2(n5409), .A(n5408), .B(n5407), .ZN(U3086)
         );
  NAND2_X1 U6122 ( .A1(n5422), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5414) );
  OAI22_X1 U6123 ( .A1(n7013), .A2(n5411), .B1(n5410), .B2(n5424), .ZN(n5412)
         );
  AOI21_X1 U6124 ( .B1(n5578), .B2(n5427), .A(n5412), .ZN(n5413) );
  OAI211_X1 U6125 ( .C1(n5415), .C2(n5431), .A(n5414), .B(n5413), .ZN(U3084)
         );
  NAND2_X1 U6126 ( .A1(n5422), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5420) );
  OAI22_X1 U6127 ( .A1(n7013), .A2(n5417), .B1(n5424), .B2(n5416), .ZN(n5418)
         );
  AOI21_X1 U6128 ( .B1(n5558), .B2(n5427), .A(n5418), .ZN(n5419) );
  OAI211_X1 U6129 ( .C1(n5431), .C2(n5421), .A(n5420), .B(n5419), .ZN(U3088)
         );
  NAND2_X1 U6130 ( .A1(n5422), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5429) );
  OAI22_X1 U6131 ( .A1(n7013), .A2(n5425), .B1(n5424), .B2(n5423), .ZN(n5426)
         );
  AOI21_X1 U6132 ( .B1(n5570), .B2(n5427), .A(n5426), .ZN(n5428) );
  OAI211_X1 U6133 ( .C1(n5431), .C2(n5430), .A(n5429), .B(n5428), .ZN(U3085)
         );
  INV_X1 U6134 ( .A(n6517), .ZN(n5432) );
  AOI22_X1 U6135 ( .A1(n6861), .A2(n5432), .B1(n5658), .B2(REIP_REG_2__SCAN_IN), .ZN(n5434) );
  NAND2_X1 U6136 ( .A1(n6856), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5433)
         );
  OAI211_X1 U6137 ( .C1(n6731), .C2(n4892), .A(n5434), .B(n5433), .ZN(n5439)
         );
  NOR2_X1 U6138 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n5435) );
  AOI211_X1 U6139 ( .C1(REIP_REG_1__SCAN_IN), .C2(REIP_REG_2__SCAN_IN), .A(
        n5435), .B(n6802), .ZN(n5436) );
  AOI21_X1 U6140 ( .B1(EBX_REG_2__SCAN_IN), .B2(n6855), .A(n5436), .ZN(n5437)
         );
  OAI21_X1 U6141 ( .B1(n6847), .B2(n6655), .A(n5437), .ZN(n5438) );
  AOI211_X1 U6142 ( .C1(n6514), .C2(n6751), .A(n5439), .B(n5438), .ZN(n5440)
         );
  INV_X1 U6143 ( .A(n5440), .ZN(U2825) );
  INV_X1 U6144 ( .A(n5441), .ZN(n5442) );
  OAI21_X1 U6145 ( .B1(n5249), .B2(n5443), .A(n5442), .ZN(n6791) );
  NOR2_X1 U6146 ( .A1(n5445), .A2(n5444), .ZN(n5446) );
  OR2_X1 U6147 ( .A1(n5497), .A2(n5446), .ZN(n6787) );
  INV_X1 U6148 ( .A(n6787), .ZN(n6681) );
  AOI22_X1 U6149 ( .A1(n6507), .A2(n6681), .B1(n6200), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n5447) );
  OAI21_X1 U6150 ( .B1(n6791), .B2(n5958), .A(n5447), .ZN(U2850) );
  INV_X1 U6151 ( .A(n5483), .ZN(n5448) );
  AOI22_X1 U6152 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n6856), .B1(n6861), 
        .B2(n5448), .ZN(n5450) );
  NAND2_X1 U6153 ( .A1(n6855), .A2(EBX_REG_3__SCAN_IN), .ZN(n5449) );
  OAI211_X1 U6154 ( .C1(n5451), .C2(n6731), .A(n5450), .B(n5449), .ZN(n5455)
         );
  NAND2_X1 U6155 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n5452) );
  OR2_X1 U6156 ( .A1(n5658), .A2(n5452), .ZN(n5453) );
  NAND3_X1 U6157 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .ZN(n6737) );
  NAND2_X1 U6158 ( .A1(n6802), .A2(n6756), .ZN(n6846) );
  OAI21_X1 U6159 ( .B1(n5658), .B2(n6737), .A(n6846), .ZN(n6733) );
  AOI21_X1 U6160 ( .B1(n4828), .B2(n5453), .A(n6733), .ZN(n5454) );
  AOI211_X1 U6161 ( .C1(n5456), .C2(n6864), .A(n5455), .B(n5454), .ZN(n5457)
         );
  OAI21_X1 U6162 ( .B1(n5476), .B2(n5458), .A(n5457), .ZN(U2824) );
  INV_X1 U6163 ( .A(DATAI_9_), .ZN(n6339) );
  OAI222_X1 U6164 ( .A1(n6791), .A2(n5976), .B1(n5975), .B2(n6339), .C1(n3422), 
        .C2(n4719), .ZN(U2882) );
  NOR2_X1 U6165 ( .A1(n5441), .A2(n5460), .ZN(n5461) );
  OR2_X1 U6166 ( .A1(n5459), .A2(n5461), .ZN(n5545) );
  XNOR2_X1 U6167 ( .A(n5497), .B(n5496), .ZN(n5474) );
  INV_X1 U6168 ( .A(n5474), .ZN(n6671) );
  AOI22_X1 U6169 ( .A1(n6864), .A2(n6671), .B1(n6855), .B2(EBX_REG_10__SCAN_IN), .ZN(n5462) );
  OAI211_X1 U6170 ( .C1(n6854), .C2(n5463), .A(n5462), .B(n6821), .ZN(n5471)
         );
  INV_X1 U6171 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6734) );
  NOR2_X1 U6172 ( .A1(n6737), .A2(n6734), .ZN(n6753) );
  NAND2_X1 U6173 ( .A1(n6753), .A2(REIP_REG_5__SCAN_IN), .ZN(n6755) );
  INV_X1 U6174 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6775) );
  INV_X1 U6175 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6435) );
  NOR3_X1 U6176 ( .A1(n6755), .A2(n6775), .A3(n6435), .ZN(n5512) );
  NAND2_X1 U6177 ( .A1(n5512), .A2(REIP_REG_8__SCAN_IN), .ZN(n5466) );
  NOR3_X1 U6178 ( .A1(n6802), .A2(REIP_REG_9__SCAN_IN), .A3(n5466), .ZN(n6785)
         );
  INV_X1 U6179 ( .A(n5466), .ZN(n5464) );
  NAND2_X1 U6180 ( .A1(n6756), .A2(n5464), .ZN(n5465) );
  AND2_X1 U6181 ( .A1(n6846), .A2(n5465), .ZN(n6786) );
  OAI21_X1 U6182 ( .B1(n6785), .B2(n6786), .A(REIP_REG_10__SCAN_IN), .ZN(n5469) );
  INV_X1 U6183 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6438) );
  NOR2_X1 U6184 ( .A1(n5466), .A2(n6438), .ZN(n5505) );
  INV_X1 U6185 ( .A(n5505), .ZN(n5467) );
  OR3_X1 U6186 ( .A1(n6802), .A2(REIP_REG_10__SCAN_IN), .A3(n5467), .ZN(n5468)
         );
  OAI211_X1 U6187 ( .C1(n5541), .C2(n6833), .A(n5469), .B(n5468), .ZN(n5470)
         );
  NOR2_X1 U6188 ( .A1(n5471), .A2(n5470), .ZN(n5472) );
  OAI21_X1 U6189 ( .B1(n5545), .B2(n6827), .A(n5472), .ZN(U2817) );
  INV_X1 U6190 ( .A(DATAI_10_), .ZN(n6335) );
  OAI222_X1 U6191 ( .A1(n5545), .A2(n5976), .B1(n5975), .B2(n6335), .C1(n3422), 
        .C2(n4802), .ZN(U2881) );
  INV_X1 U6192 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5473) );
  OAI222_X1 U6193 ( .A1(n5545), .A2(n5958), .B1(n5956), .B2(n5474), .C1(n6510), 
        .C2(n5473), .ZN(U2849) );
  OAI22_X1 U6194 ( .A1(n5476), .A2(n5475), .B1(n3792), .B2(n6731), .ZN(n5477)
         );
  AOI21_X1 U6195 ( .B1(REIP_REG_0__SCAN_IN), .B2(n6846), .A(n5477), .ZN(n5480)
         );
  NAND2_X1 U6196 ( .A1(n6854), .A2(n6833), .ZN(n5478) );
  AOI22_X1 U6197 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n5478), .B1(n6855), 
        .B2(EBX_REG_0__SCAN_IN), .ZN(n5479) );
  OAI211_X1 U6198 ( .C1(n6847), .C2(n6719), .A(n5480), .B(n5479), .ZN(U2827)
         );
  AOI21_X1 U6199 ( .B1(n6560), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n5481), 
        .ZN(n5482) );
  OAI21_X1 U6200 ( .B1(n6566), .B2(n5483), .A(n5482), .ZN(n5484) );
  AOI21_X1 U6201 ( .B1(n5485), .B2(n6561), .A(n5484), .ZN(n5486) );
  OAI21_X1 U6202 ( .B1(n5487), .B2(n6869), .A(n5486), .ZN(U2983) );
  AOI21_X1 U6203 ( .B1(n6560), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n5488), 
        .ZN(n5489) );
  OAI21_X1 U6204 ( .B1(n6566), .B2(n5511), .A(n5489), .ZN(n5490) );
  AOI21_X1 U6205 ( .B1(n5491), .B2(n6561), .A(n5490), .ZN(n5492) );
  OAI21_X1 U6206 ( .B1(n5493), .B2(n6869), .A(n5492), .ZN(U2978) );
  OR2_X1 U6207 ( .A1(n5459), .A2(n5494), .ZN(n5495) );
  AND2_X1 U6208 ( .A1(n5495), .A2(n3998), .ZN(n6549) );
  INV_X1 U6209 ( .A(n6549), .ZN(n5510) );
  NAND2_X1 U6210 ( .A1(n5497), .A2(n5496), .ZN(n5499) );
  NAND2_X1 U6211 ( .A1(n5499), .A2(n5498), .ZN(n5500) );
  AND2_X1 U6212 ( .A1(n5500), .A2(n5532), .ZN(n6688) );
  INV_X1 U6213 ( .A(n6547), .ZN(n5503) );
  AOI21_X1 U6214 ( .B1(n6856), .B2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6789), 
        .ZN(n5502) );
  NAND2_X1 U6215 ( .A1(n6855), .A2(EBX_REG_11__SCAN_IN), .ZN(n5501) );
  OAI211_X1 U6216 ( .C1(n5503), .C2(n6833), .A(n5502), .B(n5501), .ZN(n5504)
         );
  AOI21_X1 U6217 ( .B1(n6864), .B2(n6688), .A(n5504), .ZN(n5509) );
  NAND2_X1 U6218 ( .A1(n5505), .A2(REIP_REG_10__SCAN_IN), .ZN(n5506) );
  INV_X1 U6219 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6441) );
  NOR2_X1 U6220 ( .A1(n5506), .A2(n6441), .ZN(n5653) );
  OAI21_X1 U6221 ( .B1(n6802), .B2(n5653), .A(n6756), .ZN(n6809) );
  OAI21_X1 U6222 ( .B1(n6802), .B2(n5506), .A(n6441), .ZN(n5507) );
  NAND2_X1 U6223 ( .A1(n6809), .A2(n5507), .ZN(n5508) );
  OAI211_X1 U6224 ( .C1(n5510), .C2(n6827), .A(n5509), .B(n5508), .ZN(U2816)
         );
  INV_X1 U6225 ( .A(DATAI_11_), .ZN(n6333) );
  OAI222_X1 U6226 ( .A1(n5510), .A2(n5976), .B1(n5975), .B2(n6333), .C1(n3422), 
        .C2(n4717), .ZN(U2880) );
  OAI22_X1 U6227 ( .A1(n3920), .A2(n6854), .B1(n6833), .B2(n5511), .ZN(n5517)
         );
  INV_X1 U6228 ( .A(n6802), .ZN(n5513) );
  NAND2_X1 U6229 ( .A1(n5513), .A2(n5512), .ZN(n5515) );
  OAI22_X1 U6230 ( .A1(REIP_REG_8__SCAN_IN), .A2(n5515), .B1(n5514), .B2(n6796), .ZN(n5516) );
  NOR3_X1 U6231 ( .A1(n5517), .A2(n6789), .A3(n5516), .ZN(n5518) );
  OAI21_X1 U6232 ( .B1(n6847), .B2(n5519), .A(n5518), .ZN(n5520) );
  AOI21_X1 U6233 ( .B1(REIP_REG_8__SCAN_IN), .B2(n6786), .A(n5520), .ZN(n5521)
         );
  OAI21_X1 U6234 ( .B1(n5522), .B2(n6827), .A(n5521), .ZN(U2819) );
  XNOR2_X1 U6235 ( .A(n4810), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5524)
         );
  XNOR2_X1 U6236 ( .A(n5523), .B(n5524), .ZN(n6616) );
  NOR2_X1 U6237 ( .A1(n5525), .A2(n6069), .ZN(n5529) );
  INV_X1 U6238 ( .A(n6560), .ZN(n6065) );
  INV_X1 U6239 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5526) );
  OAI22_X1 U6240 ( .A1(n6065), .A2(n5527), .B1(n6821), .B2(n5526), .ZN(n5528)
         );
  AOI211_X1 U6241 ( .C1(n6548), .C2(n5527), .A(n5529), .B(n5528), .ZN(n5530)
         );
  OAI21_X1 U6242 ( .B1(n6616), .B2(n6869), .A(n5530), .ZN(U2985) );
  XNOR2_X1 U6243 ( .A(n3998), .B(n5531), .ZN(n5616) );
  INV_X1 U6244 ( .A(n5616), .ZN(n5604) );
  INV_X1 U6245 ( .A(n5532), .ZN(n5535) );
  INV_X1 U6246 ( .A(n5533), .ZN(n5534) );
  OAI21_X1 U6247 ( .B1(n5535), .B2(n5534), .A(n5645), .ZN(n5622) );
  INV_X1 U6248 ( .A(n5622), .ZN(n5536) );
  AOI22_X1 U6249 ( .A1(n5536), .A2(n6507), .B1(n6200), .B2(EBX_REG_12__SCAN_IN), .ZN(n5537) );
  OAI21_X1 U6250 ( .B1(n5604), .B2(n5958), .A(n5537), .ZN(U2847) );
  XNOR2_X1 U6251 ( .A(n6019), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5539)
         );
  XNOR2_X1 U6252 ( .A(n5538), .B(n5539), .ZN(n6675) );
  NAND2_X1 U6253 ( .A1(n6675), .A2(n6562), .ZN(n5544) );
  INV_X1 U6254 ( .A(REIP_REG_10__SCAN_IN), .ZN(n5540) );
  NOR2_X1 U6255 ( .A1(n6821), .A2(n5540), .ZN(n6670) );
  NOR2_X1 U6256 ( .A1(n6566), .A2(n5541), .ZN(n5542) );
  AOI211_X1 U6257 ( .C1(n6560), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6670), 
        .B(n5542), .ZN(n5543) );
  OAI211_X1 U6258 ( .C1(n6069), .C2(n5545), .A(n5544), .B(n5543), .ZN(U2976)
         );
  OAI21_X1 U6259 ( .B1(n5582), .B2(n7184), .A(n7039), .ZN(n5547) );
  OAI21_X1 U6260 ( .B1(n5548), .B2(n7043), .A(n5547), .ZN(n5549) );
  NAND2_X1 U6261 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n7042), .ZN(n7051) );
  NOR2_X1 U6262 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7051), .ZN(n5585)
         );
  AOI21_X1 U6263 ( .B1(n5549), .B2(n6916), .A(n5585), .ZN(n5551) );
  NOR3_X2 U6264 ( .A1(n5551), .A2(n7000), .A3(n5550), .ZN(n5589) );
  INV_X1 U6265 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5557) );
  OAI22_X1 U6266 ( .A1(n5553), .A2(n7043), .B1(n6993), .B2(n5552), .ZN(n5583)
         );
  AOI22_X1 U6267 ( .A1(n5554), .A2(n5583), .B1(n5582), .B2(n7094), .ZN(n5556)
         );
  AOI22_X1 U6268 ( .A1(n7184), .A2(n7093), .B1(n7092), .B2(n5585), .ZN(n5555)
         );
  OAI211_X1 U6269 ( .C1(n5589), .C2(n5557), .A(n5556), .B(n5555), .ZN(U3038)
         );
  INV_X1 U6270 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5561) );
  AOI22_X1 U6271 ( .A1(n5558), .A2(n5583), .B1(n5582), .B2(n7122), .ZN(n5560)
         );
  AOI22_X1 U6272 ( .A1(n7184), .A2(n7121), .B1(n7120), .B2(n5585), .ZN(n5559)
         );
  OAI211_X1 U6273 ( .C1(n5589), .C2(n5561), .A(n5560), .B(n5559), .ZN(U3040)
         );
  INV_X1 U6274 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5565) );
  AOI22_X1 U6275 ( .A1(n5562), .A2(n5583), .B1(n5582), .B2(n7136), .ZN(n5564)
         );
  AOI22_X1 U6276 ( .A1(n7184), .A2(n7135), .B1(n7134), .B2(n5585), .ZN(n5563)
         );
  OAI211_X1 U6277 ( .C1(n5589), .C2(n5565), .A(n5564), .B(n5563), .ZN(U3041)
         );
  INV_X1 U6278 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5569) );
  AOI22_X1 U6279 ( .A1(n5566), .A2(n5583), .B1(n5582), .B2(n7150), .ZN(n5568)
         );
  AOI22_X1 U6280 ( .A1(n7184), .A2(n7149), .B1(n7148), .B2(n5585), .ZN(n5567)
         );
  OAI211_X1 U6281 ( .C1(n5589), .C2(n5569), .A(n5568), .B(n5567), .ZN(U3042)
         );
  INV_X1 U6282 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5573) );
  AOI22_X1 U6283 ( .A1(n5570), .A2(n5583), .B1(n5582), .B2(n7072), .ZN(n5572)
         );
  AOI22_X1 U6284 ( .A1(n7184), .A2(n7073), .B1(n7071), .B2(n5585), .ZN(n5571)
         );
  OAI211_X1 U6285 ( .C1(n5589), .C2(n5573), .A(n5572), .B(n5571), .ZN(U3037)
         );
  INV_X1 U6286 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5577) );
  AOI22_X1 U6287 ( .A1(n5574), .A2(n5583), .B1(n5582), .B2(n7108), .ZN(n5576)
         );
  AOI22_X1 U6288 ( .A1(n7184), .A2(n7107), .B1(n7106), .B2(n5585), .ZN(n5575)
         );
  OAI211_X1 U6289 ( .C1(n5589), .C2(n5577), .A(n5576), .B(n5575), .ZN(U3039)
         );
  INV_X1 U6290 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5581) );
  AOI22_X1 U6291 ( .A1(n5578), .A2(n5583), .B1(n5582), .B2(n7056), .ZN(n5580)
         );
  AOI22_X1 U6292 ( .A1(n7184), .A2(n7048), .B1(n7047), .B2(n5585), .ZN(n5579)
         );
  OAI211_X1 U6293 ( .C1(n5589), .C2(n5581), .A(n5580), .B(n5579), .ZN(U3036)
         );
  INV_X1 U6294 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5588) );
  AOI22_X1 U6295 ( .A1(n5584), .A2(n5583), .B1(n5582), .B2(n7183), .ZN(n5587)
         );
  AOI22_X1 U6296 ( .A1(n7184), .A2(n7186), .B1(n7182), .B2(n5585), .ZN(n5586)
         );
  OAI211_X1 U6297 ( .C1(n5589), .C2(n5588), .A(n5587), .B(n5586), .ZN(U3043)
         );
  INV_X1 U6298 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6422) );
  OAI222_X1 U6299 ( .A1(n5976), .A2(n5604), .B1(n3422), .B2(n6422), .C1(n6238), 
        .C2(n5975), .ZN(U2879) );
  OAI21_X1 U6300 ( .B1(n5592), .B2(n5591), .A(n5590), .ZN(n6682) );
  INV_X1 U6301 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U6302 ( .A1(n6789), .A2(REIP_REG_9__SCAN_IN), .ZN(n6679) );
  OAI21_X1 U6303 ( .B1(n6065), .B2(n5593), .A(n6679), .ZN(n5595) );
  NOR2_X1 U6304 ( .A1(n6791), .A2(n6069), .ZN(n5594) );
  AOI211_X1 U6305 ( .C1(n6548), .C2(n6793), .A(n5595), .B(n5594), .ZN(n5596)
         );
  OAI21_X1 U6306 ( .B1(n6869), .B2(n6682), .A(n5596), .ZN(U2977) );
  INV_X1 U6307 ( .A(n5653), .ZN(n5597) );
  NOR3_X1 U6308 ( .A1(n6802), .A2(REIP_REG_12__SCAN_IN), .A3(n5597), .ZN(n6810) );
  OAI22_X1 U6309 ( .A1(n5614), .A2(n6833), .B1(n6854), .B2(n3968), .ZN(n5600)
         );
  NOR2_X1 U6310 ( .A1(n5598), .A2(n6796), .ZN(n5599) );
  NOR4_X1 U6311 ( .A1(n6810), .A2(n5600), .A3(n6789), .A4(n5599), .ZN(n5601)
         );
  OAI21_X1 U6312 ( .B1(n6847), .B2(n5622), .A(n5601), .ZN(n5602) );
  AOI21_X1 U6313 ( .B1(REIP_REG_12__SCAN_IN), .B2(n6809), .A(n5602), .ZN(n5603) );
  OAI21_X1 U6314 ( .B1(n5604), .B2(n6827), .A(n5603), .ZN(U2815) );
  INV_X1 U6315 ( .A(n5538), .ZN(n5607) );
  INV_X1 U6316 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5606) );
  OAI21_X1 U6317 ( .B1(n5607), .B2(n5606), .A(n5605), .ZN(n6546) );
  INV_X1 U6318 ( .A(n5610), .ZN(n5608) );
  AOI21_X1 U6319 ( .B1(n4540), .B2(n5609), .A(n5608), .ZN(n6545) );
  NAND2_X1 U6320 ( .A1(n6546), .A2(n6545), .ZN(n6544) );
  NAND2_X1 U6321 ( .A1(n6544), .A2(n5610), .ZN(n5612) );
  XNOR2_X1 U6322 ( .A(n3449), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5611)
         );
  XNOR2_X1 U6323 ( .A(n5612), .B(n5611), .ZN(n5627) );
  NAND2_X1 U6324 ( .A1(n6560), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5613)
         );
  NAND2_X1 U6325 ( .A1(n6789), .A2(REIP_REG_12__SCAN_IN), .ZN(n5621) );
  OAI211_X1 U6326 ( .C1(n6566), .C2(n5614), .A(n5613), .B(n5621), .ZN(n5615)
         );
  AOI21_X1 U6327 ( .B1(n5616), .B2(n6561), .A(n5615), .ZN(n5617) );
  OAI21_X1 U6328 ( .B1(n5627), .B2(n6869), .A(n5617), .ZN(U2974) );
  AOI21_X1 U6329 ( .B1(n6597), .B2(n6648), .A(n6595), .ZN(n6717) );
  OAI21_X1 U6330 ( .B1(n6717), .B2(n5609), .A(n5618), .ZN(n5625) );
  INV_X1 U6331 ( .A(n6598), .ZN(n5620) );
  INV_X1 U6332 ( .A(n6170), .ZN(n6152) );
  OAI21_X1 U6333 ( .B1(n6152), .B2(n6597), .A(n5619), .ZN(n6693) );
  INV_X1 U6334 ( .A(n6693), .ZN(n5638) );
  OAI221_X1 U6335 ( .B1(n5620), .B2(n6651), .C1(n5620), .C2(n4824), .A(n5638), 
        .ZN(n5624) );
  OAI21_X1 U6336 ( .B1(n6709), .B2(n5622), .A(n5621), .ZN(n5623) );
  AOI21_X1 U6337 ( .B1(n5625), .B2(n5624), .A(n5623), .ZN(n5626) );
  OAI21_X1 U6338 ( .B1(n5627), .B2(n6702), .A(n5626), .ZN(U3006) );
  INV_X1 U6339 ( .A(n5628), .ZN(n5631) );
  INV_X1 U6340 ( .A(n5629), .ZN(n5630) );
  NAND2_X1 U6341 ( .A1(n5631), .A2(n5630), .ZN(n5633) );
  AND2_X1 U6342 ( .A1(n5633), .A2(n5632), .ZN(n6808) );
  INV_X1 U6343 ( .A(n6808), .ZN(n5648) );
  OAI222_X1 U6344 ( .A1(n5648), .A2(n5976), .B1(n5975), .B2(n5634), .C1(n3422), 
        .C2(n4772), .ZN(U2878) );
  XNOR2_X1 U6345 ( .A(n3449), .B(n5635), .ZN(n5636) );
  XNOR2_X1 U6346 ( .A(n5637), .B(n5636), .ZN(n5673) );
  OAI21_X1 U6347 ( .B1(n6674), .B2(n5640), .A(n5638), .ZN(n6606) );
  NOR2_X1 U6348 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6717), .ZN(n5639)
         );
  AOI22_X1 U6349 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6606), .B1(n5640), .B2(n5639), .ZN(n5643) );
  XNOR2_X1 U6350 ( .A(n5647), .B(n5641), .ZN(n5664) );
  INV_X1 U6351 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5654) );
  NOR2_X1 U6352 ( .A1(n6821), .A2(n5654), .ZN(n5667) );
  AOI21_X1 U6353 ( .B1(n6721), .B2(n5664), .A(n5667), .ZN(n5642) );
  OAI211_X1 U6354 ( .C1(n5673), .C2(n6702), .A(n5643), .B(n5642), .ZN(U3004)
         );
  NAND2_X1 U6355 ( .A1(n5645), .A2(n5644), .ZN(n5646) );
  NAND2_X1 U6356 ( .A1(n5647), .A2(n5646), .ZN(n6806) );
  INV_X1 U6357 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5649) );
  OAI222_X1 U6358 ( .A1(n6806), .A2(n5956), .B1(n5649), .B2(n6510), .C1(n5648), 
        .C2(n5958), .ZN(U2846) );
  OAI21_X1 U6359 ( .B1(n5652), .B2(n5651), .A(n5650), .ZN(n5669) );
  NAND2_X1 U6360 ( .A1(n5653), .A2(REIP_REG_12__SCAN_IN), .ZN(n6798) );
  INV_X1 U6361 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6601) );
  NOR2_X1 U6362 ( .A1(n6798), .A2(n6601), .ZN(n5657) );
  NAND2_X1 U6363 ( .A1(n5654), .A2(n5657), .ZN(n5655) );
  OAI22_X1 U6364 ( .A1(n6833), .A2(n5656), .B1(n6802), .B2(n5655), .ZN(n5662)
         );
  INV_X1 U6365 ( .A(n6846), .ZN(n6825) );
  NAND2_X1 U6366 ( .A1(n5657), .A2(REIP_REG_14__SCAN_IN), .ZN(n5681) );
  NOR2_X1 U6367 ( .A1(n5658), .A2(n5681), .ZN(n5732) );
  NOR2_X1 U6368 ( .A1(n6825), .A2(n5732), .ZN(n5714) );
  AOI22_X1 U6369 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6855), .B1(
        REIP_REG_14__SCAN_IN), .B2(n5714), .ZN(n5659) );
  OAI211_X1 U6370 ( .C1(n6854), .C2(n5660), .A(n5659), .B(n6821), .ZN(n5661)
         );
  AOI211_X1 U6371 ( .C1(n6864), .C2(n5664), .A(n5662), .B(n5661), .ZN(n5663)
         );
  OAI21_X1 U6372 ( .B1(n5669), .B2(n6827), .A(n5663), .ZN(U2813) );
  AOI22_X1 U6373 ( .A1(n5664), .A2(n6507), .B1(EBX_REG_14__SCAN_IN), .B2(n6200), .ZN(n5665) );
  OAI21_X1 U6374 ( .B1(n5669), .B2(n5958), .A(n5665), .ZN(U2845) );
  INV_X1 U6375 ( .A(DATAI_14_), .ZN(n6295) );
  OAI222_X1 U6376 ( .A1(n5669), .A2(n5976), .B1(n5975), .B2(n6295), .C1(n3422), 
        .C2(n4769), .ZN(U2877) );
  AND2_X1 U6377 ( .A1(n6560), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5666)
         );
  AOI211_X1 U6378 ( .C1(n6548), .C2(n5668), .A(n5667), .B(n5666), .ZN(n5672)
         );
  INV_X1 U6379 ( .A(n5669), .ZN(n5670) );
  NAND2_X1 U6380 ( .A1(n5670), .A2(n6561), .ZN(n5671) );
  OAI211_X1 U6381 ( .C1(n5673), .C2(n6869), .A(n5672), .B(n5671), .ZN(U2972)
         );
  INV_X1 U6382 ( .A(n5674), .ZN(n5675) );
  AOI21_X1 U6383 ( .B1(n5676), .B2(n5650), .A(n5675), .ZN(n5703) );
  INV_X1 U6384 ( .A(n5703), .ZN(n5977) );
  OR2_X1 U6385 ( .A1(n5678), .A2(n5677), .ZN(n5679) );
  AND2_X1 U6386 ( .A1(n5679), .A2(n5711), .ZN(n6696) );
  NAND2_X1 U6387 ( .A1(n6856), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5680)
         );
  OAI211_X1 U6388 ( .C1(n6833), .C2(n5701), .A(n6821), .B(n5680), .ZN(n5684)
         );
  AOI22_X1 U6389 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6855), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5714), .ZN(n5682) );
  OAI21_X1 U6390 ( .B1(REIP_REG_15__SCAN_IN), .B2(n5730), .A(n5682), .ZN(n5683) );
  AOI211_X1 U6391 ( .C1(n6696), .C2(n6864), .A(n5684), .B(n5683), .ZN(n5685)
         );
  OAI21_X1 U6392 ( .B1(n5977), .B2(n6827), .A(n5685), .ZN(U2812) );
  NAND2_X1 U6393 ( .A1(n5686), .A2(n5687), .ZN(n5904) );
  OAI21_X1 U6394 ( .B1(n5686), .B2(n5687), .A(n5904), .ZN(n6815) );
  XNOR2_X1 U6395 ( .A(n3462), .B(n5688), .ZN(n6814) );
  INV_X1 U6396 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5689) );
  OAI22_X1 U6397 ( .A1(n6814), .A2(n5956), .B1(n5689), .B2(n6510), .ZN(n5690)
         );
  INV_X1 U6398 ( .A(n5690), .ZN(n5691) );
  OAI21_X1 U6399 ( .B1(n6815), .B2(n5958), .A(n5691), .ZN(U2842) );
  INV_X1 U6400 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U6401 ( .A1(n5703), .A2(n6508), .ZN(n5693) );
  NAND2_X1 U6402 ( .A1(n6696), .A2(n6507), .ZN(n5692) );
  OAI211_X1 U6403 ( .C1(n5694), .C2(n6510), .A(n5693), .B(n5692), .ZN(U2844)
         );
  INV_X1 U6404 ( .A(n5695), .ZN(n5697) );
  NAND2_X1 U6405 ( .A1(n5697), .A2(n5696), .ZN(n5698) );
  XNOR2_X1 U6406 ( .A(n5699), .B(n5698), .ZN(n6697) );
  INV_X1 U6407 ( .A(n6697), .ZN(n5705) );
  AOI22_X1 U6408 ( .A1(n6560), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6789), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5700) );
  OAI21_X1 U6409 ( .B1(n6566), .B2(n5701), .A(n5700), .ZN(n5702) );
  AOI21_X1 U6410 ( .B1(n5703), .B2(n6561), .A(n5702), .ZN(n5704) );
  OAI21_X1 U6411 ( .B1(n5705), .B2(n6869), .A(n5704), .ZN(U2971) );
  AOI22_X1 U6412 ( .A1(n7077), .A2(DATAI_17_), .B1(n7080), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U6413 ( .A1(n7081), .A2(DATAI_1_), .ZN(n5706) );
  OAI211_X1 U6414 ( .C1(n6815), .C2(n5976), .A(n5707), .B(n5706), .ZN(U2874)
         );
  AND2_X1 U6415 ( .A1(n5674), .A2(n5708), .ZN(n5709) );
  NOR2_X1 U6416 ( .A1(n5686), .A2(n5709), .ZN(n6956) );
  INV_X1 U6417 ( .A(n6956), .ZN(n5722) );
  NAND2_X1 U6418 ( .A1(n5711), .A2(n5710), .ZN(n5712) );
  NAND2_X1 U6419 ( .A1(n3462), .A2(n5712), .ZN(n6701) );
  INV_X1 U6420 ( .A(n6701), .ZN(n5719) );
  AOI21_X1 U6421 ( .B1(n6856), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6789), 
        .ZN(n5713) );
  OAI21_X1 U6422 ( .B1(n6833), .B2(n6077), .A(n5713), .ZN(n5718) );
  NAND2_X1 U6423 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .ZN(
        n5731) );
  OAI21_X1 U6424 ( .B1(REIP_REG_15__SCAN_IN), .B2(REIP_REG_16__SCAN_IN), .A(
        n5731), .ZN(n5716) );
  AOI22_X1 U6425 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6855), .B1(
        REIP_REG_16__SCAN_IN), .B2(n5714), .ZN(n5715) );
  OAI21_X1 U6426 ( .B1(n5730), .B2(n5716), .A(n5715), .ZN(n5717) );
  AOI211_X1 U6427 ( .C1(n5719), .C2(n6864), .A(n5718), .B(n5717), .ZN(n5720)
         );
  OAI21_X1 U6428 ( .B1(n5722), .B2(n6827), .A(n5720), .ZN(U2811) );
  INV_X1 U6429 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5721) );
  OAI222_X1 U6430 ( .A1(n5722), .A2(n5958), .B1(n6510), .B2(n5721), .C1(n6701), 
        .C2(n5956), .ZN(U2843) );
  XNOR2_X1 U6431 ( .A(n5723), .B(n5724), .ZN(n6498) );
  OAI21_X1 U6432 ( .B1(n5725), .B2(n5726), .A(n5950), .ZN(n5727) );
  INV_X1 U6433 ( .A(n5727), .ZN(n6589) );
  NAND2_X1 U6434 ( .A1(n6856), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5729)
         );
  NAND2_X1 U6435 ( .A1(n6861), .A2(n6054), .ZN(n5728) );
  NAND3_X1 U6436 ( .A1(n5729), .A2(n5728), .A3(n6821), .ZN(n5736) );
  NOR2_X1 U6437 ( .A1(n5731), .A2(n5730), .ZN(n6819) );
  NAND2_X1 U6438 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6819), .ZN(n5913) );
  NAND2_X1 U6439 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5806) );
  OAI21_X1 U6440 ( .B1(REIP_REG_19__SCAN_IN), .B2(REIP_REG_18__SCAN_IN), .A(
        n5806), .ZN(n5734) );
  NAND4_X1 U6441 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .A4(n5732), .ZN(n5800) );
  AND2_X1 U6442 ( .A1(n6846), .A2(n5800), .ZN(n6818) );
  AOI22_X1 U6443 ( .A1(EBX_REG_19__SCAN_IN), .A2(n6855), .B1(
        REIP_REG_19__SCAN_IN), .B2(n6818), .ZN(n5733) );
  OAI21_X1 U6444 ( .B1(n5913), .B2(n5734), .A(n5733), .ZN(n5735) );
  AOI211_X1 U6445 ( .C1(n6589), .C2(n6864), .A(n5736), .B(n5735), .ZN(n5737)
         );
  OAI21_X1 U6446 ( .B1(n6498), .B2(n6827), .A(n5737), .ZN(U2808) );
  INV_X1 U6447 ( .A(n5738), .ZN(n5740) );
  AND3_X1 U6448 ( .A1(n6921), .A2(n5740), .A3(n5739), .ZN(n5743) );
  NOR2_X1 U6449 ( .A1(n5741), .A2(n3792), .ZN(n5742) );
  AOI211_X1 U6450 ( .C1(n6197), .C2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n5743), .B(n5742), .ZN(n5744) );
  OAI21_X1 U6451 ( .B1(n5746), .B2(n5745), .A(n5744), .ZN(U3465) );
  INV_X1 U6452 ( .A(n5748), .ZN(n5749) );
  INV_X1 U6453 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6466) );
  NOR2_X1 U6454 ( .A1(n6821), .A2(n6466), .ZN(n5761) );
  INV_X1 U6455 ( .A(n5751), .ZN(n5752) );
  NOR3_X1 U6456 ( .A1(n6086), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5752), 
        .ZN(n5753) );
  AOI211_X1 U6457 ( .C1(n5783), .C2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5761), .B(n5753), .ZN(n5759) );
  INV_X1 U6458 ( .A(n5754), .ZN(n5757) );
  INV_X1 U6459 ( .A(n5793), .ZN(n5755) );
  AOI21_X1 U6460 ( .B1(n5757), .B2(n5756), .A(n5755), .ZN(n5923) );
  NAND2_X1 U6461 ( .A1(n5923), .A2(n6721), .ZN(n5758) );
  OAI211_X1 U6462 ( .C1(n5765), .C2(n6702), .A(n5759), .B(n5758), .ZN(U2989)
         );
  AOI21_X2 U6463 ( .B1(n5760), .B2(n4663), .A(n3451), .ZN(n5963) );
  AOI21_X1 U6464 ( .B1(n6560), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5761), 
        .ZN(n5762) );
  OAI21_X1 U6465 ( .B1(n6566), .B2(n5838), .A(n5762), .ZN(n5763) );
  AOI21_X1 U6466 ( .B1(n5963), .B2(n6561), .A(n5763), .ZN(n5764) );
  OAI21_X1 U6467 ( .B1(n6869), .B2(n5765), .A(n5764), .ZN(U2957) );
  INV_X1 U6468 ( .A(n5831), .ZN(n5769) );
  AOI21_X1 U6469 ( .B1(n6560), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5767), 
        .ZN(n5768) );
  OAI21_X1 U6470 ( .B1(n6566), .B2(n5769), .A(n5768), .ZN(n5770) );
  AOI21_X1 U6471 ( .B1(n5960), .B2(n6561), .A(n5770), .ZN(n5771) );
  OAI21_X1 U6472 ( .B1(n5772), .B2(n6869), .A(n5771), .ZN(U2956) );
  AND2_X1 U6473 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6179) );
  AOI22_X1 U6474 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4643), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4363), .ZN(n5773) );
  INV_X1 U6475 ( .A(n5773), .ZN(n6187) );
  NOR2_X1 U6476 ( .A1(n6924), .A2(n5774), .ZN(n5777) );
  AOI222_X1 U6477 ( .A1(n6179), .A2(n6187), .B1(n4941), .B2(n5777), .C1(n5776), 
        .C2(n5775), .ZN(n5782) );
  AOI21_X1 U6478 ( .B1(n5779), .B2(n5778), .A(n6189), .ZN(n5781) );
  OAI22_X1 U6479 ( .A1(n5782), .A2(n6189), .B1(n5781), .B2(n5780), .ZN(U3459)
         );
  INV_X1 U6480 ( .A(n5783), .ZN(n5784) );
  OAI21_X1 U6481 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n6674), .A(n5784), 
        .ZN(n5789) );
  INV_X1 U6482 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5785) );
  NOR4_X1 U6483 ( .A1(n6086), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5786), 
        .A4(n5785), .ZN(n5787) );
  AOI211_X1 U6484 ( .C1(n5789), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5788), .B(n5787), .ZN(n5798) );
  OAI22_X1 U6485 ( .A1(n5790), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4359), .ZN(n5795) );
  XOR2_X1 U6486 ( .A(n5795), .B(n5794), .Z(n5919) );
  INV_X1 U6487 ( .A(n5919), .ZN(n5796) );
  NAND2_X1 U6488 ( .A1(n5796), .A2(n6721), .ZN(n5797) );
  OAI211_X1 U6489 ( .C1(n5799), .C2(n6702), .A(n5798), .B(n5797), .ZN(U2987)
         );
  NAND2_X1 U6490 ( .A1(n5813), .A2(n6865), .ZN(n5811) );
  NOR2_X1 U6491 ( .A1(n6470), .A2(n6466), .ZN(n5802) );
  AND3_X1 U6492 ( .A1(REIP_REG_27__SCAN_IN), .A2(REIP_REG_28__SCAN_IN), .A3(
        REIP_REG_26__SCAN_IN), .ZN(n5807) );
  INV_X1 U6493 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6859) );
  INV_X1 U6494 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6452) );
  NOR3_X1 U6495 ( .A1(n6452), .A2(n5806), .A3(n5800), .ZN(n6824) );
  NAND4_X1 U6496 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_23__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n6824), .ZN(n6845) );
  NOR2_X1 U6497 ( .A1(n6859), .A2(n6845), .ZN(n5886) );
  NAND3_X1 U6498 ( .A1(n5807), .A2(REIP_REG_25__SCAN_IN), .A3(n5886), .ZN(
        n5801) );
  NAND2_X1 U6499 ( .A1(n6846), .A2(n5801), .ZN(n5849) );
  OAI21_X1 U6500 ( .B1(n5802), .B2(n6802), .A(n5849), .ZN(n5830) );
  OAI22_X1 U6501 ( .A1(n5805), .A2(n6854), .B1(n5804), .B2(n5803), .ZN(n5809)
         );
  INV_X1 U6502 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6454) );
  INV_X1 U6503 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6393) );
  NOR2_X1 U6504 ( .A1(n5806), .A2(n5913), .ZN(n6830) );
  NAND2_X1 U6505 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6830), .ZN(n6838) );
  NOR3_X1 U6506 ( .A1(n6454), .A2(n6393), .A3(n6838), .ZN(n6844) );
  NAND2_X1 U6507 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6844), .ZN(n6868) );
  INV_X1 U6508 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6004) );
  NOR3_X1 U6509 ( .A1(n6868), .A2(n6859), .A3(n6004), .ZN(n5877) );
  NAND2_X1 U6510 ( .A1(n5877), .A2(n5807), .ZN(n5845) );
  NOR4_X1 U6511 ( .A1(n5845), .A2(REIP_REG_31__SCAN_IN), .A3(n6470), .A4(n6466), .ZN(n5808) );
  AOI211_X1 U6512 ( .C1(REIP_REG_31__SCAN_IN), .C2(n5830), .A(n5809), .B(n5808), .ZN(n5810) );
  OAI211_X1 U6513 ( .C1(n5919), .C2(n6847), .A(n5811), .B(n5810), .ZN(U2796)
         );
  NAND3_X1 U6514 ( .A1(n5813), .A2(n5812), .A3(n3422), .ZN(n5815) );
  AOI22_X1 U6515 ( .A1(n7077), .A2(DATAI_31_), .B1(n7080), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U6516 ( .A1(n5815), .A2(n5814), .ZN(U2860) );
  INV_X1 U6517 ( .A(n5816), .ZN(n5822) );
  AOI21_X1 U6518 ( .B1(n5819), .B2(n5818), .A(n5817), .ZN(n5820) );
  AOI21_X1 U6519 ( .B1(n5822), .B2(n5821), .A(n5820), .ZN(n5823) );
  OAI21_X1 U6520 ( .B1(n5825), .B2(n5824), .A(n5823), .ZN(n6895) );
  NOR2_X1 U6521 ( .A1(n5826), .A2(n6581), .ZN(n6569) );
  NOR2_X1 U6522 ( .A1(n6569), .A2(n5827), .ZN(n6579) );
  OAI21_X1 U6523 ( .B1(READY_N), .B2(n6579), .A(n5828), .ZN(n6892) );
  AND2_X1 U6524 ( .A1(n6892), .A2(n5829), .ZN(n6870) );
  MUX2_X1 U6525 ( .A(MORE_REG_SCAN_IN), .B(n6895), .S(n6870), .Z(U3471) );
  INV_X1 U6526 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U6527 ( .A1(n5830), .A2(REIP_REG_30__SCAN_IN), .ZN(n5833) );
  AOI22_X1 U6528 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n6856), .B1(n6861), 
        .B2(n5831), .ZN(n5832) );
  OAI211_X1 U6529 ( .C1(n5834), .C2(n6796), .A(n5833), .B(n5832), .ZN(n5836)
         );
  NOR3_X1 U6530 ( .A1(n5845), .A2(REIP_REG_30__SCAN_IN), .A3(n6466), .ZN(n5835) );
  AOI211_X1 U6531 ( .C1(n6864), .C2(n5920), .A(n5836), .B(n5835), .ZN(n5837)
         );
  OAI21_X1 U6532 ( .B1(n5922), .B2(n6827), .A(n5837), .ZN(U2797) );
  NAND2_X1 U6533 ( .A1(n5963), .A2(n6865), .ZN(n5844) );
  OAI22_X1 U6534 ( .A1(n5839), .A2(n6854), .B1(n6833), .B2(n5838), .ZN(n5840)
         );
  AOI21_X1 U6535 ( .B1(n6855), .B2(EBX_REG_29__SCAN_IN), .A(n5840), .ZN(n5841)
         );
  OAI21_X1 U6536 ( .B1(n6466), .B2(n5849), .A(n5841), .ZN(n5842) );
  AOI21_X1 U6537 ( .B1(n5923), .B2(n6864), .A(n5842), .ZN(n5843) );
  OAI211_X1 U6538 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5845), .A(n5844), .B(n5843), .ZN(U2798) );
  NAND2_X1 U6539 ( .A1(n5986), .A2(n6865), .ZN(n5853) );
  INV_X1 U6540 ( .A(n5846), .ZN(n5984) );
  OAI22_X1 U6541 ( .A1(n5847), .A2(n6854), .B1(n6833), .B2(n5984), .ZN(n5851)
         );
  NAND3_X1 U6542 ( .A1(REIP_REG_26__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .A3(
        n5886), .ZN(n5848) );
  NAND2_X1 U6543 ( .A1(n6846), .A2(n5848), .ZN(n5875) );
  NAND2_X1 U6544 ( .A1(n5875), .A2(REIP_REG_27__SCAN_IN), .ZN(n5862) );
  INV_X1 U6545 ( .A(REIP_REG_28__SCAN_IN), .ZN(n5982) );
  AOI21_X1 U6546 ( .B1(n5862), .B2(n5982), .A(n5849), .ZN(n5850) );
  AOI211_X1 U6547 ( .C1(n6855), .C2(EBX_REG_28__SCAN_IN), .A(n5851), .B(n5850), 
        .ZN(n5852) );
  OAI211_X1 U6548 ( .C1(n6847), .C2(n6080), .A(n5853), .B(n5852), .ZN(U2799)
         );
  NAND2_X1 U6549 ( .A1(n5854), .A2(n5855), .ZN(n5856) );
  NAND2_X1 U6550 ( .A1(n5857), .A2(n5856), .ZN(n5995) );
  INV_X1 U6551 ( .A(n5877), .ZN(n5858) );
  INV_X1 U6552 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5998) );
  OAI21_X1 U6553 ( .B1(n5858), .B2(n5998), .A(n6461), .ZN(n5863) );
  AOI22_X1 U6554 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n6856), .B1(n6861), 
        .B2(n5992), .ZN(n5860) );
  NAND2_X1 U6555 ( .A1(n6855), .A2(EBX_REG_27__SCAN_IN), .ZN(n5859) );
  OAI211_X1 U6556 ( .C1(n5926), .C2(n6847), .A(n5860), .B(n5859), .ZN(n5861)
         );
  AOI21_X1 U6557 ( .B1(n5863), .B2(n5862), .A(n5861), .ZN(n5864) );
  OAI21_X1 U6558 ( .B1(n5995), .B2(n6827), .A(n5864), .ZN(U2800) );
  INV_X1 U6559 ( .A(n5854), .ZN(n5865) );
  AOI21_X1 U6560 ( .B1(n5867), .B2(n5866), .A(n5865), .ZN(n6002) );
  INV_X1 U6561 ( .A(n6002), .ZN(n5972) );
  OAI22_X1 U6562 ( .A1(n5868), .A2(n6854), .B1(n6833), .B2(n6000), .ZN(n5874)
         );
  INV_X1 U6563 ( .A(n5883), .ZN(n5872) );
  INV_X1 U6564 ( .A(n5869), .ZN(n5870) );
  OAI21_X1 U6565 ( .B1(n5872), .B2(n5871), .A(n5870), .ZN(n6099) );
  NOR2_X1 U6566 ( .A1(n6099), .A2(n6847), .ZN(n5873) );
  AOI211_X1 U6567 ( .C1(n6855), .C2(EBX_REG_26__SCAN_IN), .A(n5874), .B(n5873), 
        .ZN(n5879) );
  INV_X1 U6568 ( .A(n5875), .ZN(n5876) );
  OAI21_X1 U6569 ( .B1(n5877), .B2(REIP_REG_26__SCAN_IN), .A(n5876), .ZN(n5878) );
  OAI211_X1 U6570 ( .C1(n5972), .C2(n6827), .A(n5879), .B(n5878), .ZN(U2801)
         );
  XOR2_X1 U6571 ( .A(n5881), .B(n5880), .Z(n7079) );
  NOR3_X1 U6572 ( .A1(n6868), .A2(n6859), .A3(REIP_REG_25__SCAN_IN), .ZN(n5892) );
  INV_X1 U6573 ( .A(n6111), .ZN(n5882) );
  NOR2_X1 U6574 ( .A1(n6112), .A2(n5882), .ZN(n5885) );
  OAI21_X1 U6575 ( .B1(n5885), .B2(n5884), .A(n5883), .ZN(n6110) );
  NOR3_X1 U6576 ( .A1(n6825), .A2(n5886), .A3(n6004), .ZN(n5889) );
  INV_X1 U6577 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5887) );
  OAI22_X1 U6578 ( .A1(n6005), .A2(n6854), .B1(n5887), .B2(n6796), .ZN(n5888)
         );
  AOI211_X1 U6579 ( .C1(n6861), .C2(n6007), .A(n5889), .B(n5888), .ZN(n5890)
         );
  OAI21_X1 U6580 ( .B1(n6110), .B2(n6847), .A(n5890), .ZN(n5891) );
  AOI211_X1 U6581 ( .C1(n7079), .C2(n6865), .A(n5892), .B(n5891), .ZN(n5893)
         );
  INV_X1 U6582 ( .A(n5893), .ZN(U2802) );
  OAI21_X1 U6583 ( .B1(n3453), .B2(n4156), .A(n5895), .ZN(n6976) );
  OAI22_X1 U6584 ( .A1(n6838), .A2(REIP_REG_21__SCAN_IN), .B1(n6825), .B2(
        n6824), .ZN(n5901) );
  OAI22_X1 U6585 ( .A1(n4151), .A2(n6854), .B1(n6040), .B2(n6833), .ZN(n5900)
         );
  OAI21_X1 U6586 ( .B1(n5943), .B2(n5896), .A(n5933), .ZN(n6138) );
  NOR3_X1 U6587 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6393), .A3(n6838), .ZN(n5897) );
  AOI21_X1 U6588 ( .B1(n6855), .B2(EBX_REG_22__SCAN_IN), .A(n5897), .ZN(n5898)
         );
  OAI21_X1 U6589 ( .B1(n6138), .B2(n6847), .A(n5898), .ZN(n5899) );
  AOI211_X1 U6590 ( .C1(n5901), .C2(REIP_REG_22__SCAN_IN), .A(n5900), .B(n5899), .ZN(n5902) );
  OAI21_X1 U6591 ( .B1(n6976), .B2(n6827), .A(n5902), .ZN(U2805) );
  NAND2_X1 U6592 ( .A1(n5904), .A2(n5903), .ZN(n5905) );
  AND2_X1 U6593 ( .A1(n5723), .A2(n5905), .ZN(n6959) );
  INV_X1 U6594 ( .A(n6959), .ZN(n5959) );
  INV_X1 U6595 ( .A(n5725), .ZN(n5906) );
  OAI21_X1 U6596 ( .B1(n5908), .B2(n5907), .A(n5906), .ZN(n6173) );
  INV_X1 U6597 ( .A(n6173), .ZN(n5916) );
  NAND2_X1 U6598 ( .A1(n6856), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5911)
         );
  INV_X1 U6599 ( .A(n6559), .ZN(n5909) );
  NAND2_X1 U6600 ( .A1(n6861), .A2(n5909), .ZN(n5910) );
  NAND3_X1 U6601 ( .A1(n5911), .A2(n5910), .A3(n6821), .ZN(n5915) );
  AOI22_X1 U6602 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6855), .B1(
        REIP_REG_18__SCAN_IN), .B2(n6818), .ZN(n5912) );
  OAI21_X1 U6603 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5913), .A(n5912), .ZN(n5914) );
  AOI211_X1 U6604 ( .C1(n5916), .C2(n6864), .A(n5915), .B(n5914), .ZN(n5917)
         );
  OAI21_X1 U6605 ( .B1(n5959), .B2(n6827), .A(n5917), .ZN(U2809) );
  OAI22_X1 U6606 ( .A1(n5919), .A2(n5956), .B1(n6510), .B2(n5918), .ZN(U2828)
         );
  AOI22_X1 U6607 ( .A1(n5920), .A2(n6507), .B1(EBX_REG_30__SCAN_IN), .B2(n6200), .ZN(n5921) );
  OAI21_X1 U6608 ( .B1(n5922), .B2(n5958), .A(n5921), .ZN(U2829) );
  INV_X1 U6609 ( .A(n5963), .ZN(n5925) );
  AOI22_X1 U6610 ( .A1(n5923), .A2(n6507), .B1(n6200), .B2(EBX_REG_29__SCAN_IN), .ZN(n5924) );
  OAI21_X1 U6611 ( .B1(n5925), .B2(n5958), .A(n5924), .ZN(U2830) );
  INV_X1 U6612 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5927) );
  OAI222_X1 U6613 ( .A1(n5927), .A2(n6510), .B1(n5956), .B2(n5926), .C1(n5995), 
        .C2(n5958), .ZN(U2832) );
  INV_X1 U6614 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5928) );
  OAI222_X1 U6615 ( .A1(n5928), .A2(n6510), .B1(n5956), .B2(n6099), .C1(n5972), 
        .C2(n5958), .ZN(U2833) );
  INV_X1 U6616 ( .A(n7079), .ZN(n6013) );
  OAI222_X1 U6617 ( .A1(n5958), .A2(n6013), .B1(n6510), .B2(n5887), .C1(n6110), 
        .C2(n5956), .ZN(U2834) );
  NAND2_X1 U6618 ( .A1(n5895), .A2(n5930), .ZN(n5931) );
  AND2_X1 U6619 ( .A1(n5929), .A2(n5931), .ZN(n6851) );
  INV_X1 U6620 ( .A(n6851), .ZN(n5936) );
  NAND2_X1 U6621 ( .A1(n5933), .A2(n5932), .ZN(n5934) );
  NAND2_X1 U6622 ( .A1(n6112), .A2(n5934), .ZN(n6848) );
  OAI222_X1 U6623 ( .A1(n5958), .A2(n5936), .B1(n6510), .B2(n5935), .C1(n6848), 
        .C2(n5956), .ZN(U2836) );
  INV_X1 U6624 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5937) );
  OAI222_X1 U6625 ( .A1(n5937), .A2(n6510), .B1(n5956), .B2(n6138), .C1(n6976), 
        .C2(n5958), .ZN(U2837) );
  INV_X1 U6626 ( .A(n5938), .ZN(n5940) );
  INV_X1 U6627 ( .A(n6973), .ZN(n5945) );
  AND2_X1 U6628 ( .A1(n5952), .A2(n5941), .ZN(n5942) );
  NOR2_X1 U6629 ( .A1(n5943), .A2(n5942), .ZN(n6837) );
  AOI22_X1 U6630 ( .A1(n6837), .A2(n6507), .B1(EBX_REG_21__SCAN_IN), .B2(n6200), .ZN(n5944) );
  OAI21_X1 U6631 ( .B1(n5945), .B2(n5958), .A(n5944), .ZN(U2838) );
  NOR2_X1 U6632 ( .A1(n5946), .A2(n5947), .ZN(n5948) );
  OR2_X1 U6633 ( .A1(n5938), .A2(n5948), .ZN(n6828) );
  NAND2_X1 U6634 ( .A1(n5950), .A2(n5949), .ZN(n5951) );
  NAND2_X1 U6635 ( .A1(n5952), .A2(n5951), .ZN(n6826) );
  OAI22_X1 U6636 ( .A1(n6826), .A2(n5956), .B1(n5953), .B2(n6510), .ZN(n5954)
         );
  AOI21_X1 U6637 ( .B1(n6970), .B2(n6508), .A(n5954), .ZN(n5955) );
  INV_X1 U6638 ( .A(n5955), .ZN(U2839) );
  INV_X1 U6639 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5957) );
  OAI222_X1 U6640 ( .A1(n5959), .A2(n5958), .B1(n6510), .B2(n5957), .C1(n5956), 
        .C2(n6173), .ZN(U2841) );
  NAND2_X1 U6641 ( .A1(n5960), .A2(n7078), .ZN(n5962) );
  AOI22_X1 U6642 ( .A1(n7077), .A2(DATAI_30_), .B1(n7080), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5961) );
  OAI211_X1 U6643 ( .C1(n6963), .C2(n6295), .A(n5962), .B(n5961), .ZN(U2861)
         );
  NAND2_X1 U6644 ( .A1(n5963), .A2(n7078), .ZN(n5965) );
  AOI22_X1 U6645 ( .A1(n7077), .A2(DATAI_29_), .B1(n7080), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5964) );
  OAI211_X1 U6646 ( .C1(n6963), .C2(n5634), .A(n5965), .B(n5964), .ZN(U2862)
         );
  NAND2_X1 U6647 ( .A1(n5986), .A2(n7078), .ZN(n5967) );
  AOI22_X1 U6648 ( .A1(n7077), .A2(DATAI_28_), .B1(n7080), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5966) );
  OAI211_X1 U6649 ( .C1(n6963), .C2(n6238), .A(n5967), .B(n5966), .ZN(U2863)
         );
  AOI22_X1 U6650 ( .A1(n7077), .A2(DATAI_27_), .B1(n7080), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U6651 ( .A1(n7081), .A2(DATAI_11_), .ZN(n5968) );
  OAI211_X1 U6652 ( .C1(n5995), .C2(n5976), .A(n5969), .B(n5968), .ZN(U2864)
         );
  AOI22_X1 U6653 ( .A1(n7077), .A2(DATAI_26_), .B1(n7080), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U6654 ( .A1(n7081), .A2(DATAI_10_), .ZN(n5970) );
  OAI211_X1 U6655 ( .C1(n5972), .C2(n5976), .A(n5971), .B(n5970), .ZN(U2865)
         );
  NAND2_X1 U6656 ( .A1(n6851), .A2(n7078), .ZN(n5974) );
  AOI22_X1 U6657 ( .A1(n7077), .A2(DATAI_23_), .B1(n7080), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5973) );
  OAI211_X1 U6658 ( .C1(n6963), .C2(n6342), .A(n5974), .B(n5973), .ZN(U2868)
         );
  OAI222_X1 U6659 ( .A1(n5977), .A2(n5976), .B1(n6296), .B2(n5975), .C1(n3422), 
        .C2(n4745), .ZN(U2876) );
  NAND2_X1 U6660 ( .A1(n5979), .A2(n5978), .ZN(n5981) );
  XNOR2_X1 U6661 ( .A(n3449), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5980)
         );
  XNOR2_X1 U6662 ( .A(n5981), .B(n5980), .ZN(n6092) );
  NOR2_X1 U6663 ( .A1(n6821), .A2(n5982), .ZN(n6088) );
  AOI21_X1 U6664 ( .B1(n6560), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n6088), 
        .ZN(n5983) );
  OAI21_X1 U6665 ( .B1(n6566), .B2(n5984), .A(n5983), .ZN(n5985) );
  AOI21_X1 U6666 ( .B1(n5986), .B2(n6561), .A(n5985), .ZN(n5987) );
  OAI21_X1 U6667 ( .B1(n6092), .B2(n6869), .A(n5987), .ZN(U2958) );
  NAND2_X1 U6668 ( .A1(n5988), .A2(n6562), .ZN(n5994) );
  NOR2_X1 U6669 ( .A1(n6065), .A2(n5989), .ZN(n5990) );
  AOI211_X1 U6670 ( .C1(n6548), .C2(n5992), .A(n5991), .B(n5990), .ZN(n5993)
         );
  OAI211_X1 U6671 ( .C1(n6069), .C2(n5995), .A(n5994), .B(n5993), .ZN(U2959)
         );
  XNOR2_X1 U6672 ( .A(n3449), .B(n6096), .ZN(n5997) );
  XNOR2_X1 U6673 ( .A(n5996), .B(n5997), .ZN(n6103) );
  NOR2_X1 U6674 ( .A1(n6821), .A2(n5998), .ZN(n6098) );
  AOI21_X1 U6675 ( .B1(n6560), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n6098), 
        .ZN(n5999) );
  OAI21_X1 U6676 ( .B1(n6566), .B2(n6000), .A(n5999), .ZN(n6001) );
  AOI21_X1 U6677 ( .B1(n6002), .B2(n6561), .A(n6001), .ZN(n6003) );
  OAI21_X1 U6678 ( .B1(n6869), .B2(n6103), .A(n6003), .ZN(U2960) );
  NOR2_X1 U6679 ( .A1(n6821), .A2(n6004), .ZN(n6107) );
  NOR2_X1 U6680 ( .A1(n6065), .A2(n6005), .ZN(n6006) );
  AOI211_X1 U6681 ( .C1(n6548), .C2(n6007), .A(n6107), .B(n6006), .ZN(n6012)
         );
  OAI21_X1 U6682 ( .B1(n3438), .B2(n6010), .A(n6009), .ZN(n6104) );
  NAND2_X1 U6683 ( .A1(n6104), .A2(n6562), .ZN(n6011) );
  OAI211_X1 U6684 ( .C1(n6013), .C2(n6069), .A(n6012), .B(n6011), .ZN(U2961)
         );
  INV_X1 U6686 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U6687 ( .A1(n4540), .A2(n6016), .ZN(n6146) );
  OR2_X1 U6688 ( .A1(n4540), .A2(n6016), .ZN(n6017) );
  AND2_X1 U6689 ( .A1(n6146), .A2(n6017), .ZN(n6051) );
  AND2_X1 U6690 ( .A1(n6015), .A2(n6051), .ZN(n6050) );
  NAND4_X1 U6691 ( .A1(n6050), .A2(n6019), .A3(n6132), .A4(n6018), .ZN(n6031)
         );
  OAI21_X1 U6692 ( .B1(n6156), .B2(n3449), .A(n6015), .ZN(n6020) );
  OAI21_X1 U6693 ( .B1(n6019), .B2(n6155), .A(n6020), .ZN(n6044) );
  XNOR2_X1 U6694 ( .A(n3449), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6045)
         );
  INV_X1 U6695 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6021) );
  AOI22_X1 U6696 ( .A1(n6044), .A2(n6045), .B1(n3449), .B2(n6021), .ZN(n6039)
         );
  NAND4_X1 U6697 ( .A1(n6039), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .A4(n4540), .ZN(n6022) );
  OAI21_X1 U6698 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n6031), .A(n6022), 
        .ZN(n6023) );
  XNOR2_X1 U6699 ( .A(n6023), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6121)
         );
  NOR2_X1 U6700 ( .A1(n6821), .A2(n6859), .ZN(n6119) );
  NOR2_X1 U6701 ( .A1(n6065), .A2(n6024), .ZN(n6025) );
  AOI211_X1 U6702 ( .C1(n6548), .C2(n6862), .A(n6119), .B(n6025), .ZN(n6028)
         );
  AOI21_X1 U6703 ( .B1(n6026), .B2(n5929), .A(n5880), .ZN(n7060) );
  NAND2_X1 U6704 ( .A1(n7060), .A2(n6561), .ZN(n6027) );
  OAI211_X1 U6705 ( .C1(n6121), .C2(n6869), .A(n6028), .B(n6027), .ZN(U2962)
         );
  INV_X1 U6706 ( .A(n6123), .ZN(n6133) );
  NAND4_X1 U6707 ( .A1(n6029), .A2(n6155), .A3(n6133), .A4(n4540), .ZN(n6030)
         );
  NAND2_X1 U6708 ( .A1(n6031), .A2(n6030), .ZN(n6032) );
  XNOR2_X1 U6709 ( .A(n6032), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6130)
         );
  INV_X1 U6710 ( .A(n6843), .ZN(n6035) );
  INV_X1 U6711 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6033) );
  NOR2_X1 U6712 ( .A1(n6821), .A2(n6033), .ZN(n6125) );
  AOI21_X1 U6713 ( .B1(n6560), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n6125), 
        .ZN(n6034) );
  OAI21_X1 U6714 ( .B1(n6566), .B2(n6035), .A(n6034), .ZN(n6036) );
  AOI21_X1 U6715 ( .B1(n6851), .B2(n6561), .A(n6036), .ZN(n6037) );
  OAI21_X1 U6716 ( .B1(n6130), .B2(n6869), .A(n6037), .ZN(U2963) );
  XNOR2_X1 U6717 ( .A(n6019), .B(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6038)
         );
  XNOR2_X1 U6718 ( .A(n6039), .B(n6038), .ZN(n6131) );
  NAND2_X1 U6719 ( .A1(n6131), .A2(n6562), .ZN(n6043) );
  NOR2_X1 U6720 ( .A1(n6821), .A2(n6454), .ZN(n6135) );
  NOR2_X1 U6721 ( .A1(n6566), .A2(n6040), .ZN(n6041) );
  AOI211_X1 U6722 ( .C1(n6560), .C2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n6135), 
        .B(n6041), .ZN(n6042) );
  OAI211_X1 U6723 ( .C1(n6069), .C2(n6976), .A(n6043), .B(n6042), .ZN(U2964)
         );
  XOR2_X1 U6724 ( .A(n6045), .B(n6044), .Z(n6145) );
  INV_X1 U6725 ( .A(n6835), .ZN(n6047) );
  NOR2_X1 U6726 ( .A1(n6821), .A2(n6393), .ZN(n6141) );
  AOI21_X1 U6727 ( .B1(n6560), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n6141), 
        .ZN(n6046) );
  OAI21_X1 U6728 ( .B1(n6566), .B2(n6047), .A(n6046), .ZN(n6048) );
  AOI21_X1 U6729 ( .B1(n6973), .B2(n6561), .A(n6048), .ZN(n6049) );
  OAI21_X1 U6730 ( .B1(n6145), .B2(n6869), .A(n6049), .ZN(U2965) );
  INV_X1 U6731 ( .A(n6050), .ZN(n6147) );
  OAI21_X1 U6732 ( .B1(n6051), .B2(n6015), .A(n6147), .ZN(n6590) );
  NAND2_X1 U6733 ( .A1(n6590), .A2(n6562), .ZN(n6056) );
  INV_X1 U6734 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6052) );
  OAI22_X1 U6735 ( .A1(n6065), .A2(n4101), .B1(n6821), .B2(n6052), .ZN(n6053)
         );
  AOI21_X1 U6736 ( .B1(n6548), .B2(n6054), .A(n6053), .ZN(n6055) );
  OAI211_X1 U6737 ( .C1(n6069), .C2(n6498), .A(n6056), .B(n6055), .ZN(U2967)
         );
  NAND2_X1 U6738 ( .A1(n4540), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6164) );
  NOR2_X1 U6739 ( .A1(n3449), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6060)
         );
  INV_X1 U6740 ( .A(n6060), .ZN(n6057) );
  NAND2_X1 U6741 ( .A1(n6057), .A2(n6164), .ZN(n6059) );
  MUX2_X1 U6742 ( .A(n6164), .B(n6059), .S(n6058), .Z(n6062) );
  INV_X1 U6743 ( .A(n6058), .ZN(n6061) );
  NAND2_X1 U6744 ( .A1(n6061), .A2(n6060), .ZN(n6163) );
  NAND2_X1 U6745 ( .A1(n6062), .A2(n6163), .ZN(n6713) );
  NAND2_X1 U6746 ( .A1(n6713), .A2(n6562), .ZN(n6068) );
  INV_X1 U6747 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6064) );
  INV_X1 U6748 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6063) );
  OAI22_X1 U6749 ( .A1(n6065), .A2(n6064), .B1(n6821), .B2(n6063), .ZN(n6066)
         );
  AOI21_X1 U6750 ( .B1(n6548), .B2(n6817), .A(n6066), .ZN(n6067) );
  OAI211_X1 U6751 ( .C1(n6069), .C2(n6815), .A(n6068), .B(n6067), .ZN(U2969)
         );
  INV_X1 U6752 ( .A(n6071), .ZN(n6075) );
  OAI21_X1 U6753 ( .B1(n6073), .B2(n6075), .A(n6072), .ZN(n6074) );
  OAI21_X1 U6754 ( .B1(n6070), .B2(n6075), .A(n6074), .ZN(n6703) );
  AOI22_X1 U6755 ( .A1(n6560), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6789), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n6076) );
  OAI21_X1 U6756 ( .B1(n6566), .B2(n6077), .A(n6076), .ZN(n6078) );
  AOI21_X1 U6757 ( .B1(n6956), .B2(n6561), .A(n6078), .ZN(n6079) );
  OAI21_X1 U6758 ( .B1(n6703), .B2(n6869), .A(n6079), .ZN(U2970) );
  NOR2_X1 U6759 ( .A1(n6080), .A2(n6709), .ZN(n6090) );
  INV_X1 U6760 ( .A(n6081), .ZN(n6083) );
  AOI21_X1 U6761 ( .B1(n6084), .B2(n6083), .A(n6082), .ZN(n6089) );
  INV_X1 U6762 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6085) );
  NOR3_X1 U6763 ( .A1(n6086), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n6085), 
        .ZN(n6087) );
  NOR4_X1 U6764 ( .A1(n6090), .A2(n6089), .A3(n6088), .A4(n6087), .ZN(n6091)
         );
  OAI21_X1 U6765 ( .B1(n6092), .B2(n6702), .A(n6091), .ZN(U2990) );
  INV_X1 U6766 ( .A(n6093), .ZN(n6105) );
  AOI211_X1 U6767 ( .C1(n6096), .C2(n6095), .A(n6094), .B(n6105), .ZN(n6097)
         );
  AOI211_X1 U6768 ( .C1(n6114), .C2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n6098), .B(n6097), .ZN(n6102) );
  INV_X1 U6769 ( .A(n6099), .ZN(n6100) );
  NAND2_X1 U6770 ( .A1(n6100), .A2(n6721), .ZN(n6101) );
  OAI211_X1 U6771 ( .C1(n6103), .C2(n6702), .A(n6102), .B(n6101), .ZN(U2992)
         );
  NAND2_X1 U6772 ( .A1(n6104), .A2(n6723), .ZN(n6109) );
  NOR2_X1 U6773 ( .A1(n6105), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6106)
         );
  AOI211_X1 U6774 ( .C1(n6114), .C2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n6107), .B(n6106), .ZN(n6108) );
  OAI211_X1 U6775 ( .C1(n6709), .C2(n6110), .A(n6109), .B(n6108), .ZN(U2993)
         );
  XNOR2_X1 U6776 ( .A(n6112), .B(n6111), .ZN(n6863) );
  INV_X1 U6777 ( .A(n6139), .ZN(n6113) );
  NAND3_X1 U6778 ( .A1(n6113), .A2(n6133), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6116) );
  INV_X1 U6779 ( .A(n6114), .ZN(n6115) );
  AOI21_X1 U6780 ( .B1(n6117), .B2(n6116), .A(n6115), .ZN(n6118) );
  AOI211_X1 U6781 ( .C1(n6721), .C2(n6863), .A(n6119), .B(n6118), .ZN(n6120)
         );
  OAI21_X1 U6782 ( .B1(n6121), .B2(n6702), .A(n6120), .ZN(U2994) );
  INV_X1 U6783 ( .A(n6122), .ZN(n6126) );
  NOR3_X1 U6784 ( .A1(n6139), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n6123), 
        .ZN(n6124) );
  AOI211_X1 U6785 ( .C1(n6126), .C2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n6125), .B(n6124), .ZN(n6129) );
  INV_X1 U6786 ( .A(n6848), .ZN(n6127) );
  NAND2_X1 U6787 ( .A1(n6127), .A2(n6721), .ZN(n6128) );
  OAI211_X1 U6788 ( .C1(n6130), .C2(n6702), .A(n6129), .B(n6128), .ZN(U2995)
         );
  NAND2_X1 U6789 ( .A1(n6131), .A2(n6723), .ZN(n6137) );
  NOR3_X1 U6790 ( .A1(n6139), .A2(n6133), .A3(n6132), .ZN(n6134) );
  AOI211_X1 U6791 ( .C1(n6142), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n6135), .B(n6134), .ZN(n6136) );
  OAI211_X1 U6792 ( .C1(n6709), .C2(n6138), .A(n6137), .B(n6136), .ZN(U2996)
         );
  NOR2_X1 U6793 ( .A1(n6139), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6140)
         );
  AOI211_X1 U6794 ( .C1(n6142), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n6141), .B(n6140), .ZN(n6144) );
  NAND2_X1 U6795 ( .A1(n6837), .A2(n6721), .ZN(n6143) );
  OAI211_X1 U6796 ( .C1(n6145), .C2(n6702), .A(n6144), .B(n6143), .ZN(U2997)
         );
  NAND2_X1 U6797 ( .A1(n6147), .A2(n6146), .ZN(n6149) );
  XNOR2_X1 U6798 ( .A(n4540), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6148)
         );
  XNOR2_X1 U6799 ( .A(n6149), .B(n6148), .ZN(n6563) );
  INV_X1 U6800 ( .A(n6563), .ZN(n6161) );
  NAND2_X1 U6801 ( .A1(n6612), .A2(n6165), .ZN(n6150) );
  OAI211_X1 U6802 ( .C1(n6152), .C2(n6151), .A(n6168), .B(n6150), .ZN(n6588)
         );
  OAI22_X1 U6803 ( .A1(n6826), .A2(n6709), .B1(n6821), .B2(n6452), .ZN(n6153)
         );
  AOI21_X1 U6804 ( .B1(INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n6588), .A(n6153), 
        .ZN(n6160) );
  NOR2_X1 U6805 ( .A1(n6717), .A2(n6154), .ZN(n6162) );
  NAND2_X1 U6806 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6162), .ZN(n6593) );
  NOR2_X1 U6807 ( .A1(n6155), .A2(n6593), .ZN(n6158) );
  INV_X1 U6808 ( .A(n6156), .ZN(n6157) );
  NAND2_X1 U6809 ( .A1(n6158), .A2(n6157), .ZN(n6159) );
  OAI211_X1 U6810 ( .C1(n6161), .C2(n6702), .A(n6160), .B(n6159), .ZN(U2998)
         );
  INV_X1 U6811 ( .A(n6162), .ZN(n6178) );
  OAI21_X1 U6812 ( .B1(n6070), .B2(n6164), .A(n6163), .ZN(n6166) );
  XNOR2_X1 U6813 ( .A(n6166), .B(n6165), .ZN(n6556) );
  NAND2_X1 U6814 ( .A1(n6556), .A2(n6723), .ZN(n6177) );
  INV_X1 U6815 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6710) );
  NAND2_X1 U6816 ( .A1(n6167), .A2(n6710), .ZN(n6716) );
  INV_X1 U6817 ( .A(n6168), .ZN(n6169) );
  AOI21_X1 U6818 ( .B1(n6171), .B2(n6170), .A(n6169), .ZN(n6711) );
  OAI21_X1 U6819 ( .B1(n4824), .B2(n6716), .A(n6711), .ZN(n6175) );
  INV_X1 U6820 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6172) );
  OAI22_X1 U6821 ( .A1(n6173), .A2(n6709), .B1(n6821), .B2(n6172), .ZN(n6174)
         );
  AOI21_X1 U6822 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6175), .A(n6174), 
        .ZN(n6176) );
  OAI211_X1 U6823 ( .C1(INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n6178), .A(n6177), .B(n6176), .ZN(U3000) );
  INV_X1 U6824 ( .A(n6179), .ZN(n6188) );
  NOR2_X1 U6825 ( .A1(n6181), .A2(n6180), .ZN(n6186) );
  OAI21_X1 U6826 ( .B1(n6186), .B2(n6183), .A(n6182), .ZN(n6184) );
  AOI21_X1 U6827 ( .B1(n4893), .B2(n6185), .A(n6184), .ZN(n6879) );
  OAI222_X1 U6828 ( .A1(n6188), .A2(n6187), .B1(n6186), .B2(n6924), .C1(n6910), 
        .C2(n6879), .ZN(n6190) );
  INV_X1 U6829 ( .A(n6189), .ZN(n6875) );
  MUX2_X1 U6830 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n6190), .S(n6875), 
        .Z(U3460) );
  INV_X1 U6831 ( .A(n6191), .ZN(n6193) );
  OAI22_X1 U6832 ( .A1(n6193), .A2(n6910), .B1(n6192), .B2(n6924), .ZN(n6194)
         );
  MUX2_X1 U6833 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6194), .S(n6875), 
        .Z(U3456) );
  INV_X1 U6834 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6944) );
  NAND2_X1 U6835 ( .A1(STATE_REG_1__SCAN_IN), .A2(n6944), .ZN(n6952) );
  INV_X1 U6836 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6574) );
  AOI21_X1 U6837 ( .B1(n6574), .B2(STATE_REG_1__SCAN_IN), .A(n6944), .ZN(n6199) );
  NOR2_X1 U6838 ( .A1(n6955), .A2(n6199), .ZN(n6933) );
  NOR2_X1 U6839 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6567) );
  OAI21_X1 U6840 ( .B1(BS16_N), .B2(n6567), .A(n6933), .ZN(n6931) );
  OAI21_X1 U6841 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6933), .A(n6931), .ZN(
        n6195) );
  INV_X1 U6842 ( .A(n6195), .ZN(U3451) );
  INV_X1 U6843 ( .A(n6933), .ZN(n6196) );
  AND2_X1 U6844 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6196), .ZN(U3180) );
  AND2_X1 U6845 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6196), .ZN(U3179) );
  AND2_X1 U6846 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6196), .ZN(U3178) );
  AND2_X1 U6847 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6196), .ZN(U3177) );
  AND2_X1 U6848 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6196), .ZN(U3176) );
  AND2_X1 U6849 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6196), .ZN(U3175) );
  AND2_X1 U6850 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6196), .ZN(U3174) );
  AND2_X1 U6851 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6196), .ZN(U3173) );
  AND2_X1 U6852 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6196), .ZN(U3172) );
  AND2_X1 U6853 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6196), .ZN(U3171) );
  AND2_X1 U6854 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6196), .ZN(U3170) );
  AND2_X1 U6855 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6196), .ZN(U3169) );
  AND2_X1 U6856 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6196), .ZN(U3168) );
  AND2_X1 U6857 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6196), .ZN(U3167) );
  AND2_X1 U6858 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6196), .ZN(U3166) );
  AND2_X1 U6859 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6196), .ZN(U3165) );
  AND2_X1 U6860 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6196), .ZN(U3164) );
  AND2_X1 U6861 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6196), .ZN(U3163) );
  AND2_X1 U6862 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6196), .ZN(U3162) );
  AND2_X1 U6863 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6196), .ZN(U3161) );
  AND2_X1 U6864 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6196), .ZN(U3160) );
  AND2_X1 U6865 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6196), .ZN(U3159) );
  AND2_X1 U6866 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6196), .ZN(U3158) );
  AND2_X1 U6867 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6196), .ZN(U3157) );
  AND2_X1 U6868 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6196), .ZN(U3156) );
  AND2_X1 U6869 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6196), .ZN(U3155) );
  AND2_X1 U6870 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6196), .ZN(U3154) );
  AND2_X1 U6871 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6196), .ZN(U3153) );
  AND2_X1 U6872 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6196), .ZN(U3152) );
  AND2_X1 U6873 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6196), .ZN(U3151) );
  AND2_X1 U6874 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6197), .ZN(U3019)
         );
  AND2_X1 U6875 ( .A1(n6198), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U6876 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6352) );
  AOI21_X1 U6877 ( .B1(n6199), .B2(n6352), .A(n6955), .ZN(U2789) );
  NAND2_X1 U6878 ( .A1(n6507), .A2(n6688), .ZN(n6202) );
  NAND2_X1 U6879 ( .A1(n6200), .A2(EBX_REG_11__SCAN_IN), .ZN(n6201) );
  NAND2_X1 U6880 ( .A1(n6202), .A2(n6201), .ZN(n6203) );
  AOI21_X1 U6881 ( .B1(n6549), .B2(n6508), .A(n6203), .ZN(n6405) );
  OAI22_X1 U6882 ( .A1(REIP_REG_27__SCAN_IN), .A2(keyinput_119), .B1(
        REIP_REG_26__SCAN_IN), .B2(keyinput_120), .ZN(n6204) );
  AOI221_X1 U6883 ( .B1(REIP_REG_27__SCAN_IN), .B2(keyinput_119), .C1(
        keyinput_120), .C2(REIP_REG_26__SCAN_IN), .A(n6204), .ZN(n6403) );
  INV_X1 U6884 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6206) );
  INV_X1 U6885 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6483) );
  OAI22_X1 U6886 ( .A1(n6206), .A2(keyinput_114), .B1(n6483), .B2(keyinput_113), .ZN(n6205) );
  AOI221_X1 U6887 ( .B1(n6206), .B2(keyinput_114), .C1(keyinput_113), .C2(
        n6483), .A(n6205), .ZN(n6281) );
  INV_X1 U6888 ( .A(keyinput_112), .ZN(n6279) );
  INV_X1 U6889 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6486) );
  INV_X1 U6890 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6489) );
  INV_X1 U6891 ( .A(keyinput_111), .ZN(n6277) );
  INV_X1 U6892 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6573) );
  INV_X1 U6893 ( .A(keyinput_110), .ZN(n6275) );
  OAI22_X1 U6894 ( .A1(n6341), .A2(keyinput_87), .B1(DATAI_7_), .B2(
        keyinput_88), .ZN(n6207) );
  AOI221_X1 U6895 ( .B1(n6341), .B2(keyinput_87), .C1(keyinput_88), .C2(
        DATAI_7_), .A(n6207), .ZN(n6252) );
  INV_X1 U6896 ( .A(keyinput_86), .ZN(n6245) );
  INV_X1 U6897 ( .A(keyinput_85), .ZN(n6243) );
  INV_X1 U6898 ( .A(keyinput_84), .ZN(n6241) );
  INV_X1 U6899 ( .A(keyinput_83), .ZN(n6239) );
  OAI22_X1 U6900 ( .A1(DATAI_17_), .A2(keyinput_78), .B1(DATAI_16_), .B2(
        keyinput_79), .ZN(n6208) );
  AOI221_X1 U6901 ( .B1(DATAI_17_), .B2(keyinput_78), .C1(keyinput_79), .C2(
        DATAI_16_), .A(n6208), .ZN(n6233) );
  INV_X1 U6902 ( .A(DATAI_18_), .ZN(n6231) );
  INV_X1 U6903 ( .A(DATAI_19_), .ZN(n6210) );
  OAI22_X1 U6904 ( .A1(n6210), .A2(keyinput_76), .B1(DATAI_20_), .B2(
        keyinput_75), .ZN(n6209) );
  AOI221_X1 U6905 ( .B1(n6210), .B2(keyinput_76), .C1(keyinput_75), .C2(
        DATAI_20_), .A(n6209), .ZN(n6229) );
  INV_X1 U6906 ( .A(DATAI_21_), .ZN(n6303) );
  INV_X1 U6907 ( .A(DATAI_24_), .ZN(n6212) );
  OAI22_X1 U6908 ( .A1(n6212), .A2(keyinput_71), .B1(keyinput_69), .B2(
        DATAI_26_), .ZN(n6211) );
  AOI221_X1 U6909 ( .B1(n6212), .B2(keyinput_71), .C1(DATAI_26_), .C2(
        keyinput_69), .A(n6211), .ZN(n6221) );
  INV_X1 U6910 ( .A(keyinput_68), .ZN(n6219) );
  INV_X1 U6911 ( .A(DATAI_27_), .ZN(n6312) );
  INV_X1 U6912 ( .A(DATAI_28_), .ZN(n6309) );
  INV_X1 U6913 ( .A(keyinput_67), .ZN(n6217) );
  INV_X1 U6914 ( .A(keyinput_66), .ZN(n6215) );
  INV_X1 U6915 ( .A(DATAI_29_), .ZN(n6307) );
  AOI22_X1 U6916 ( .A1(DATAI_30_), .A2(keyinput_65), .B1(DATAI_31_), .B2(
        keyinput_64), .ZN(n6213) );
  OAI221_X1 U6917 ( .B1(DATAI_30_), .B2(keyinput_65), .C1(DATAI_31_), .C2(
        keyinput_64), .A(n6213), .ZN(n6214) );
  OAI221_X1 U6918 ( .B1(DATAI_29_), .B2(n6215), .C1(n6307), .C2(keyinput_66), 
        .A(n6214), .ZN(n6216) );
  OAI221_X1 U6919 ( .B1(DATAI_28_), .B2(keyinput_67), .C1(n6309), .C2(n6217), 
        .A(n6216), .ZN(n6218) );
  OAI221_X1 U6920 ( .B1(DATAI_27_), .B2(n6219), .C1(n6312), .C2(keyinput_68), 
        .A(n6218), .ZN(n6220) );
  OAI211_X1 U6921 ( .C1(DATAI_25_), .C2(keyinput_70), .A(n6221), .B(n6220), 
        .ZN(n6222) );
  AOI21_X1 U6922 ( .B1(DATAI_25_), .B2(keyinput_70), .A(n6222), .ZN(n6226) );
  INV_X1 U6923 ( .A(DATAI_22_), .ZN(n6224) );
  AOI22_X1 U6924 ( .A1(DATAI_23_), .A2(keyinput_72), .B1(n6224), .B2(
        keyinput_73), .ZN(n6223) );
  OAI221_X1 U6925 ( .B1(DATAI_23_), .B2(keyinput_72), .C1(n6224), .C2(
        keyinput_73), .A(n6223), .ZN(n6225) );
  AOI211_X1 U6926 ( .C1(n6303), .C2(keyinput_74), .A(n6226), .B(n6225), .ZN(
        n6227) );
  OAI21_X1 U6927 ( .B1(n6303), .B2(keyinput_74), .A(n6227), .ZN(n6228) );
  AOI22_X1 U6928 ( .A1(keyinput_77), .A2(n6231), .B1(n6229), .B2(n6228), .ZN(
        n6230) );
  OAI21_X1 U6929 ( .B1(n6231), .B2(keyinput_77), .A(n6230), .ZN(n6232) );
  AOI22_X1 U6930 ( .A1(n6233), .A2(n6232), .B1(DATAI_13_), .B2(keyinput_82), 
        .ZN(n6234) );
  OAI21_X1 U6931 ( .B1(DATAI_13_), .B2(keyinput_82), .A(n6234), .ZN(n6237) );
  AOI22_X1 U6932 ( .A1(DATAI_14_), .A2(keyinput_81), .B1(n6296), .B2(
        keyinput_80), .ZN(n6235) );
  OAI221_X1 U6933 ( .B1(DATAI_14_), .B2(keyinput_81), .C1(n6296), .C2(
        keyinput_80), .A(n6235), .ZN(n6236) );
  OAI222_X1 U6934 ( .A1(DATAI_12_), .A2(n6239), .B1(n6238), .B2(keyinput_83), 
        .C1(n6237), .C2(n6236), .ZN(n6240) );
  OAI221_X1 U6935 ( .B1(DATAI_11_), .B2(keyinput_84), .C1(n6333), .C2(n6241), 
        .A(n6240), .ZN(n6242) );
  OAI221_X1 U6936 ( .B1(DATAI_10_), .B2(keyinput_85), .C1(n6335), .C2(n6243), 
        .A(n6242), .ZN(n6244) );
  OAI221_X1 U6937 ( .B1(DATAI_9_), .B2(keyinput_86), .C1(n6339), .C2(n6245), 
        .A(n6244), .ZN(n6251) );
  AOI22_X1 U6938 ( .A1(n6344), .A2(keyinput_91), .B1(n6247), .B2(keyinput_89), 
        .ZN(n6246) );
  OAI221_X1 U6939 ( .B1(n6344), .B2(keyinput_91), .C1(n6247), .C2(keyinput_89), 
        .A(n6246), .ZN(n6250) );
  AOI22_X1 U6940 ( .A1(DATAI_3_), .A2(keyinput_92), .B1(DATAI_5_), .B2(
        keyinput_90), .ZN(n6248) );
  OAI221_X1 U6941 ( .B1(DATAI_3_), .B2(keyinput_92), .C1(DATAI_5_), .C2(
        keyinput_90), .A(n6248), .ZN(n6249) );
  AOI211_X1 U6942 ( .C1(n6252), .C2(n6251), .A(n6250), .B(n6249), .ZN(n6267)
         );
  INV_X1 U6943 ( .A(HOLD), .ZN(n6935) );
  OAI22_X1 U6944 ( .A1(n6935), .A2(keyinput_100), .B1(BS16_N), .B2(keyinput_98), .ZN(n6253) );
  AOI221_X1 U6945 ( .B1(n6935), .B2(keyinput_100), .C1(keyinput_98), .C2(
        BS16_N), .A(n6253), .ZN(n6256) );
  INV_X1 U6946 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6572) );
  OAI22_X1 U6947 ( .A1(n6572), .A2(keyinput_101), .B1(keyinput_102), .B2(
        ADS_N_REG_SCAN_IN), .ZN(n6254) );
  AOI221_X1 U6948 ( .B1(n6572), .B2(keyinput_101), .C1(ADS_N_REG_SCAN_IN), 
        .C2(keyinput_102), .A(n6254), .ZN(n6255) );
  OAI211_X1 U6949 ( .C1(READY_N), .C2(keyinput_99), .A(n6256), .B(n6255), .ZN(
        n6257) );
  AOI21_X1 U6950 ( .B1(READY_N), .B2(keyinput_99), .A(n6257), .ZN(n6266) );
  INV_X1 U6951 ( .A(NA_N), .ZN(n6946) );
  AOI22_X1 U6952 ( .A1(n6946), .A2(keyinput_97), .B1(n6962), .B2(keyinput_93), 
        .ZN(n6258) );
  OAI221_X1 U6953 ( .B1(n6946), .B2(keyinput_97), .C1(n6962), .C2(keyinput_93), 
        .A(n6258), .ZN(n6261) );
  AOI22_X1 U6954 ( .A1(DATAI_1_), .A2(keyinput_94), .B1(n6954), .B2(
        keyinput_96), .ZN(n6259) );
  OAI221_X1 U6955 ( .B1(DATAI_1_), .B2(keyinput_94), .C1(n6954), .C2(
        keyinput_96), .A(n6259), .ZN(n6260) );
  AOI211_X1 U6956 ( .C1(keyinput_95), .C2(DATAI_0_), .A(n6261), .B(n6260), 
        .ZN(n6262) );
  OAI21_X1 U6957 ( .B1(keyinput_95), .B2(DATAI_0_), .A(n6262), .ZN(n6265) );
  AOI22_X1 U6958 ( .A1(keyinput_104), .A2(M_IO_N_REG_SCAN_IN), .B1(n6358), 
        .B2(keyinput_103), .ZN(n6263) );
  OAI221_X1 U6959 ( .B1(keyinput_104), .B2(M_IO_N_REG_SCAN_IN), .C1(n6358), 
        .C2(keyinput_103), .A(n6263), .ZN(n6264) );
  AOI221_X1 U6960 ( .B1(n6267), .B2(n6266), .C1(n6265), .C2(n6266), .A(n6264), 
        .ZN(n6273) );
  INV_X1 U6961 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6937) );
  AOI22_X1 U6962 ( .A1(keyinput_105), .A2(D_C_N_REG_SCAN_IN), .B1(n6937), .B2(
        keyinput_106), .ZN(n6268) );
  OAI221_X1 U6963 ( .B1(keyinput_105), .B2(D_C_N_REG_SCAN_IN), .C1(n6937), 
        .C2(keyinput_106), .A(n6268), .ZN(n6272) );
  OAI22_X1 U6964 ( .A1(STATEBS16_REG_SCAN_IN), .A2(keyinput_107), .B1(
        FLUSH_REG_SCAN_IN), .B2(keyinput_109), .ZN(n6269) );
  AOI221_X1 U6965 ( .B1(STATEBS16_REG_SCAN_IN), .B2(keyinput_107), .C1(
        keyinput_109), .C2(FLUSH_REG_SCAN_IN), .A(n6269), .ZN(n6271) );
  XNOR2_X1 U6966 ( .A(MORE_REG_SCAN_IN), .B(keyinput_108), .ZN(n6270) );
  OAI211_X1 U6967 ( .C1(n6273), .C2(n6272), .A(n6271), .B(n6270), .ZN(n6274)
         );
  OAI221_X1 U6968 ( .B1(W_R_N_REG_SCAN_IN), .B2(keyinput_110), .C1(n6573), 
        .C2(n6275), .A(n6274), .ZN(n6276) );
  OAI221_X1 U6969 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_111), .C1(
        n6489), .C2(n6277), .A(n6276), .ZN(n6278) );
  OAI221_X1 U6970 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(n6279), .C1(n6486), 
        .C2(keyinput_112), .A(n6278), .ZN(n6280) );
  AOI22_X1 U6971 ( .A1(n6281), .A2(n6280), .B1(REIP_REG_31__SCAN_IN), .B2(
        keyinput_115), .ZN(n6282) );
  OAI21_X1 U6972 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_115), .A(n6282), 
        .ZN(n6285) );
  AOI22_X1 U6973 ( .A1(n6466), .A2(keyinput_117), .B1(n6470), .B2(keyinput_116), .ZN(n6283) );
  OAI221_X1 U6974 ( .B1(n6466), .B2(keyinput_117), .C1(n6470), .C2(
        keyinput_116), .A(n6283), .ZN(n6284) );
  OAI22_X1 U6975 ( .A1(n6285), .A2(n6284), .B1(REIP_REG_28__SCAN_IN), .B2(
        keyinput_118), .ZN(n6286) );
  AOI21_X1 U6976 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput_118), .A(n6286), 
        .ZN(n6402) );
  OAI22_X1 U6977 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_50), .B1(
        BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_49), .ZN(n6287) );
  AOI221_X1 U6978 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_50), .C1(
        keyinput_49), .C2(BYTEENABLE_REG_2__SCAN_IN), .A(n6287), .ZN(n6375) );
  INV_X1 U6979 ( .A(keyinput_48), .ZN(n6373) );
  INV_X1 U6980 ( .A(keyinput_47), .ZN(n6371) );
  INV_X1 U6981 ( .A(keyinput_46), .ZN(n6369) );
  XOR2_X1 U6982 ( .A(READY_N), .B(keyinput_35), .Z(n6361) );
  OAI22_X1 U6983 ( .A1(n6946), .A2(keyinput_33), .B1(DATAI_2_), .B2(
        keyinput_29), .ZN(n6288) );
  AOI221_X1 U6984 ( .B1(n6946), .B2(keyinput_33), .C1(keyinput_29), .C2(
        DATAI_2_), .A(n6288), .ZN(n6292) );
  OAI22_X1 U6985 ( .A1(n6290), .A2(keyinput_30), .B1(keyinput_31), .B2(
        DATAI_0_), .ZN(n6289) );
  AOI221_X1 U6986 ( .B1(n6290), .B2(keyinput_30), .C1(DATAI_0_), .C2(
        keyinput_31), .A(n6289), .ZN(n6291) );
  OAI211_X1 U6987 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_32), .A(n6292), 
        .B(n6291), .ZN(n6293) );
  AOI21_X1 U6988 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_32), .A(n6293), 
        .ZN(n6356) );
  INV_X1 U6989 ( .A(keyinput_22), .ZN(n6338) );
  INV_X1 U6990 ( .A(keyinput_21), .ZN(n6336) );
  INV_X1 U6991 ( .A(keyinput_20), .ZN(n6332) );
  AOI22_X1 U6992 ( .A1(n6296), .A2(keyinput_16), .B1(n6295), .B2(keyinput_17), 
        .ZN(n6294) );
  OAI221_X1 U6993 ( .B1(n6296), .B2(keyinput_16), .C1(n6295), .C2(keyinput_17), 
        .A(n6294), .ZN(n6329) );
  INV_X1 U6994 ( .A(DATAI_16_), .ZN(n6299) );
  INV_X1 U6995 ( .A(DATAI_17_), .ZN(n6298) );
  AOI22_X1 U6996 ( .A1(n6299), .A2(keyinput_15), .B1(n6298), .B2(keyinput_14), 
        .ZN(n6297) );
  OAI221_X1 U6997 ( .B1(n6299), .B2(keyinput_15), .C1(n6298), .C2(keyinput_14), 
        .A(n6297), .ZN(n6327) );
  INV_X1 U6998 ( .A(DATAI_20_), .ZN(n6301) );
  AOI22_X1 U6999 ( .A1(DATAI_19_), .A2(keyinput_12), .B1(n6301), .B2(
        keyinput_11), .ZN(n6300) );
  OAI221_X1 U7000 ( .B1(DATAI_19_), .B2(keyinput_12), .C1(n6301), .C2(
        keyinput_11), .A(n6300), .ZN(n6323) );
  INV_X1 U7001 ( .A(DATAI_23_), .ZN(n6321) );
  OAI22_X1 U7002 ( .A1(n6303), .A2(keyinput_10), .B1(DATAI_22_), .B2(
        keyinput_9), .ZN(n6302) );
  AOI221_X1 U7003 ( .B1(n6303), .B2(keyinput_10), .C1(keyinput_9), .C2(
        DATAI_22_), .A(n6302), .ZN(n6319) );
  INV_X1 U7004 ( .A(keyinput_4), .ZN(n6313) );
  INV_X1 U7005 ( .A(keyinput_3), .ZN(n6310) );
  INV_X1 U7006 ( .A(keyinput_2), .ZN(n6306) );
  OAI22_X1 U7007 ( .A1(DATAI_31_), .A2(keyinput_0), .B1(keyinput_1), .B2(
        DATAI_30_), .ZN(n6304) );
  AOI221_X1 U7008 ( .B1(DATAI_31_), .B2(keyinput_0), .C1(DATAI_30_), .C2(
        keyinput_1), .A(n6304), .ZN(n6305) );
  AOI221_X1 U7009 ( .B1(DATAI_29_), .B2(keyinput_2), .C1(n6307), .C2(n6306), 
        .A(n6305), .ZN(n6308) );
  AOI221_X1 U7010 ( .B1(DATAI_28_), .B2(n6310), .C1(n6309), .C2(keyinput_3), 
        .A(n6308), .ZN(n6311) );
  AOI221_X1 U7011 ( .B1(DATAI_27_), .B2(n6313), .C1(n6312), .C2(keyinput_4), 
        .A(n6311), .ZN(n6316) );
  AOI22_X1 U7012 ( .A1(DATAI_24_), .A2(keyinput_7), .B1(DATAI_26_), .B2(
        keyinput_5), .ZN(n6314) );
  OAI221_X1 U7013 ( .B1(DATAI_24_), .B2(keyinput_7), .C1(DATAI_26_), .C2(
        keyinput_5), .A(n6314), .ZN(n6315) );
  AOI211_X1 U7014 ( .C1(DATAI_25_), .C2(keyinput_6), .A(n6316), .B(n6315), 
        .ZN(n6317) );
  OAI21_X1 U7015 ( .B1(DATAI_25_), .B2(keyinput_6), .A(n6317), .ZN(n6318) );
  OAI211_X1 U7016 ( .C1(n6321), .C2(keyinput_8), .A(n6319), .B(n6318), .ZN(
        n6320) );
  AOI21_X1 U7017 ( .B1(n6321), .B2(keyinput_8), .A(n6320), .ZN(n6322) );
  OAI22_X1 U7018 ( .A1(n6323), .A2(n6322), .B1(keyinput_13), .B2(DATAI_18_), 
        .ZN(n6324) );
  AOI21_X1 U7019 ( .B1(keyinput_13), .B2(DATAI_18_), .A(n6324), .ZN(n6326) );
  NAND2_X1 U7020 ( .A1(keyinput_18), .A2(DATAI_13_), .ZN(n6325) );
  OAI221_X1 U7021 ( .B1(n6327), .B2(n6326), .C1(keyinput_18), .C2(DATAI_13_), 
        .A(n6325), .ZN(n6328) );
  OAI22_X1 U7022 ( .A1(n6329), .A2(n6328), .B1(keyinput_19), .B2(DATAI_12_), 
        .ZN(n6330) );
  AOI21_X1 U7023 ( .B1(keyinput_19), .B2(DATAI_12_), .A(n6330), .ZN(n6331) );
  AOI221_X1 U7024 ( .B1(DATAI_11_), .B2(keyinput_20), .C1(n6333), .C2(n6332), 
        .A(n6331), .ZN(n6334) );
  AOI221_X1 U7025 ( .B1(DATAI_10_), .B2(n6336), .C1(n6335), .C2(keyinput_21), 
        .A(n6334), .ZN(n6337) );
  AOI221_X1 U7026 ( .B1(DATAI_9_), .B2(keyinput_22), .C1(n6339), .C2(n6338), 
        .A(n6337), .ZN(n6349) );
  AOI22_X1 U7027 ( .A1(n6342), .A2(keyinput_24), .B1(n6341), .B2(keyinput_23), 
        .ZN(n6340) );
  OAI221_X1 U7028 ( .B1(n6342), .B2(keyinput_24), .C1(n6341), .C2(keyinput_23), 
        .A(n6340), .ZN(n6348) );
  OAI22_X1 U7029 ( .A1(n6344), .A2(keyinput_27), .B1(keyinput_26), .B2(
        DATAI_5_), .ZN(n6343) );
  AOI221_X1 U7030 ( .B1(n6344), .B2(keyinput_27), .C1(DATAI_5_), .C2(
        keyinput_26), .A(n6343), .ZN(n6347) );
  OAI22_X1 U7031 ( .A1(DATAI_6_), .A2(keyinput_25), .B1(DATAI_3_), .B2(
        keyinput_28), .ZN(n6345) );
  AOI221_X1 U7032 ( .B1(DATAI_6_), .B2(keyinput_25), .C1(keyinput_28), .C2(
        DATAI_3_), .A(n6345), .ZN(n6346) );
  OAI211_X1 U7033 ( .C1(n6349), .C2(n6348), .A(n6347), .B(n6346), .ZN(n6355)
         );
  AOI22_X1 U7034 ( .A1(READREQUEST_REG_SCAN_IN), .A2(keyinput_37), .B1(n6935), 
        .B2(keyinput_36), .ZN(n6350) );
  OAI221_X1 U7035 ( .B1(READREQUEST_REG_SCAN_IN), .B2(keyinput_37), .C1(n6935), 
        .C2(keyinput_36), .A(n6350), .ZN(n6354) );
  AOI22_X1 U7036 ( .A1(BS16_N), .A2(keyinput_34), .B1(n6352), .B2(keyinput_38), 
        .ZN(n6351) );
  OAI221_X1 U7037 ( .B1(BS16_N), .B2(keyinput_34), .C1(n6352), .C2(keyinput_38), .A(n6351), .ZN(n6353) );
  AOI211_X1 U7038 ( .C1(n6356), .C2(n6355), .A(n6354), .B(n6353), .ZN(n6360)
         );
  AOI22_X1 U7039 ( .A1(M_IO_N_REG_SCAN_IN), .A2(keyinput_40), .B1(n6358), .B2(
        keyinput_39), .ZN(n6357) );
  OAI221_X1 U7040 ( .B1(M_IO_N_REG_SCAN_IN), .B2(keyinput_40), .C1(n6358), 
        .C2(keyinput_39), .A(n6357), .ZN(n6359) );
  AOI21_X1 U7041 ( .B1(n6361), .B2(n6360), .A(n6359), .ZN(n6367) );
  AOI22_X1 U7042 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_42), .B1(
        D_C_N_REG_SCAN_IN), .B2(keyinput_41), .ZN(n6362) );
  OAI221_X1 U7043 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_42), .C1(
        D_C_N_REG_SCAN_IN), .C2(keyinput_41), .A(n6362), .ZN(n6366) );
  OAI22_X1 U7044 ( .A1(n6930), .A2(keyinput_43), .B1(keyinput_45), .B2(
        FLUSH_REG_SCAN_IN), .ZN(n6363) );
  AOI221_X1 U7045 ( .B1(n6930), .B2(keyinput_43), .C1(FLUSH_REG_SCAN_IN), .C2(
        keyinput_45), .A(n6363), .ZN(n6365) );
  XNOR2_X1 U7046 ( .A(MORE_REG_SCAN_IN), .B(keyinput_44), .ZN(n6364) );
  OAI211_X1 U7047 ( .C1(n6367), .C2(n6366), .A(n6365), .B(n6364), .ZN(n6368)
         );
  OAI221_X1 U7048 ( .B1(W_R_N_REG_SCAN_IN), .B2(n6369), .C1(n6573), .C2(
        keyinput_46), .A(n6368), .ZN(n6370) );
  OAI221_X1 U7049 ( .B1(BYTEENABLE_REG_0__SCAN_IN), .B2(n6371), .C1(n6489), 
        .C2(keyinput_47), .A(n6370), .ZN(n6372) );
  OAI221_X1 U7050 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_48), .C1(
        n6486), .C2(n6373), .A(n6372), .ZN(n6374) );
  AOI22_X1 U7051 ( .A1(n6375), .A2(n6374), .B1(REIP_REG_31__SCAN_IN), .B2(
        keyinput_51), .ZN(n6376) );
  OAI21_X1 U7052 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_51), .A(n6376), 
        .ZN(n6379) );
  AOI22_X1 U7053 ( .A1(REIP_REG_30__SCAN_IN), .A2(keyinput_52), .B1(n6466), 
        .B2(keyinput_53), .ZN(n6377) );
  OAI221_X1 U7054 ( .B1(REIP_REG_30__SCAN_IN), .B2(keyinput_52), .C1(n6466), 
        .C2(keyinput_53), .A(n6377), .ZN(n6378) );
  OAI22_X1 U7055 ( .A1(n6379), .A2(n6378), .B1(n5982), .B2(keyinput_54), .ZN(
        n6380) );
  AOI21_X1 U7056 ( .B1(n5982), .B2(keyinput_54), .A(n6380), .ZN(n6391) );
  OAI22_X1 U7057 ( .A1(n6461), .A2(keyinput_55), .B1(n5998), .B2(keyinput_56), 
        .ZN(n6381) );
  AOI221_X1 U7058 ( .B1(n6461), .B2(keyinput_55), .C1(keyinput_56), .C2(n5998), 
        .A(n6381), .ZN(n6390) );
  AOI22_X1 U7059 ( .A1(REIP_REG_20__SCAN_IN), .A2(keyinput_62), .B1(n6052), 
        .B2(keyinput_63), .ZN(n6382) );
  OAI221_X1 U7060 ( .B1(REIP_REG_20__SCAN_IN), .B2(keyinput_62), .C1(n6052), 
        .C2(keyinput_63), .A(n6382), .ZN(n6389) );
  AOI22_X1 U7061 ( .A1(n6004), .A2(keyinput_57), .B1(n6033), .B2(keyinput_59), 
        .ZN(n6383) );
  OAI221_X1 U7062 ( .B1(n6004), .B2(keyinput_57), .C1(n6033), .C2(keyinput_59), 
        .A(n6383), .ZN(n6386) );
  AOI22_X1 U7063 ( .A1(REIP_REG_21__SCAN_IN), .A2(keyinput_61), .B1(n6454), 
        .B2(keyinput_60), .ZN(n6384) );
  OAI221_X1 U7064 ( .B1(REIP_REG_21__SCAN_IN), .B2(keyinput_61), .C1(n6454), 
        .C2(keyinput_60), .A(n6384), .ZN(n6385) );
  AOI211_X1 U7065 ( .C1(keyinput_58), .C2(REIP_REG_24__SCAN_IN), .A(n6386), 
        .B(n6385), .ZN(n6387) );
  OAI21_X1 U7066 ( .B1(keyinput_58), .B2(REIP_REG_24__SCAN_IN), .A(n6387), 
        .ZN(n6388) );
  AOI211_X1 U7067 ( .C1(n6391), .C2(n6390), .A(n6389), .B(n6388), .ZN(n6401)
         );
  OAI22_X1 U7068 ( .A1(n6393), .A2(keyinput_125), .B1(keyinput_124), .B2(
        REIP_REG_22__SCAN_IN), .ZN(n6392) );
  AOI221_X1 U7069 ( .B1(n6393), .B2(keyinput_125), .C1(REIP_REG_22__SCAN_IN), 
        .C2(keyinput_124), .A(n6392), .ZN(n6399) );
  OAI22_X1 U7070 ( .A1(n6004), .A2(keyinput_121), .B1(REIP_REG_24__SCAN_IN), 
        .B2(keyinput_122), .ZN(n6394) );
  AOI221_X1 U7071 ( .B1(n6004), .B2(keyinput_121), .C1(keyinput_122), .C2(
        REIP_REG_24__SCAN_IN), .A(n6394), .ZN(n6398) );
  OAI22_X1 U7072 ( .A1(n6452), .A2(keyinput_126), .B1(n6052), .B2(keyinput_127), .ZN(n6395) );
  AOI221_X1 U7073 ( .B1(n6452), .B2(keyinput_126), .C1(keyinput_127), .C2(
        n6052), .A(n6395), .ZN(n6397) );
  XNOR2_X1 U7074 ( .A(REIP_REG_23__SCAN_IN), .B(keyinput_123), .ZN(n6396) );
  NAND4_X1 U7075 ( .A1(n6399), .A2(n6398), .A3(n6397), .A4(n6396), .ZN(n6400)
         );
  AOI211_X1 U7076 ( .C1(n6403), .C2(n6402), .A(n6401), .B(n6400), .ZN(n6404)
         );
  XNOR2_X1 U7077 ( .A(n6405), .B(n6404), .ZN(U2848) );
  AOI22_X1 U7078 ( .A1(n6585), .A2(LWORD_REG_0__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6407) );
  OAI21_X1 U7079 ( .B1(n6408), .B2(n6427), .A(n6407), .ZN(U2923) );
  AOI22_X1 U7080 ( .A1(n6585), .A2(LWORD_REG_1__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6409) );
  OAI21_X1 U7081 ( .B1(n4721), .B2(n6427), .A(n6409), .ZN(U2922) );
  AOI22_X1 U7082 ( .A1(n6585), .A2(LWORD_REG_2__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6410) );
  OAI21_X1 U7083 ( .B1(n4809), .B2(n6427), .A(n6410), .ZN(U2921) );
  AOI22_X1 U7084 ( .A1(n6585), .A2(LWORD_REG_3__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6411) );
  OAI21_X1 U7085 ( .B1(n6412), .B2(n6427), .A(n6411), .ZN(U2920) );
  AOI22_X1 U7086 ( .A1(n6585), .A2(LWORD_REG_4__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6413) );
  OAI21_X1 U7087 ( .B1(n4763), .B2(n6427), .A(n6413), .ZN(U2919) );
  AOI22_X1 U7088 ( .A1(n6585), .A2(LWORD_REG_5__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6414) );
  OAI21_X1 U7089 ( .B1(n3875), .B2(n6427), .A(n6414), .ZN(U2918) );
  AOI22_X1 U7090 ( .A1(n6585), .A2(LWORD_REG_6__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6415) );
  OAI21_X1 U7091 ( .B1(n4779), .B2(n6427), .A(n6415), .ZN(U2917) );
  AOI22_X1 U7092 ( .A1(n6585), .A2(LWORD_REG_7__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6416) );
  OAI21_X1 U7093 ( .B1(n4774), .B2(n6427), .A(n6416), .ZN(U2916) );
  AOI22_X1 U7094 ( .A1(n6585), .A2(LWORD_REG_8__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6417) );
  OAI21_X1 U7095 ( .B1(n4791), .B2(n6427), .A(n6417), .ZN(U2915) );
  AOI22_X1 U7096 ( .A1(n6585), .A2(LWORD_REG_9__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6418) );
  OAI21_X1 U7097 ( .B1(n4719), .B2(n6427), .A(n6418), .ZN(U2914) );
  AOI22_X1 U7098 ( .A1(n6585), .A2(LWORD_REG_10__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6419) );
  OAI21_X1 U7099 ( .B1(n4802), .B2(n6427), .A(n6419), .ZN(U2913) );
  AOI22_X1 U7100 ( .A1(n6585), .A2(LWORD_REG_11__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6420) );
  OAI21_X1 U7101 ( .B1(n4717), .B2(n6427), .A(n6420), .ZN(U2912) );
  AOI22_X1 U7102 ( .A1(n6585), .A2(LWORD_REG_12__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6421) );
  OAI21_X1 U7103 ( .B1(n6422), .B2(n6427), .A(n6421), .ZN(U2911) );
  AOI22_X1 U7104 ( .A1(n6585), .A2(LWORD_REG_13__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6423) );
  OAI21_X1 U7105 ( .B1(n4772), .B2(n6427), .A(n6423), .ZN(U2910) );
  AOI22_X1 U7106 ( .A1(n6585), .A2(LWORD_REG_14__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6424) );
  OAI21_X1 U7107 ( .B1(n4769), .B2(n6427), .A(n6424), .ZN(U2909) );
  AOI22_X1 U7108 ( .A1(n6585), .A2(LWORD_REG_15__SCAN_IN), .B1(n6198), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6426) );
  OAI21_X1 U7109 ( .B1(n4745), .B2(n6427), .A(n6426), .ZN(U2908) );
  INV_X1 U7110 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6654) );
  NAND2_X1 U7111 ( .A1(n6955), .A2(n6574), .ZN(n6464) );
  NOR2_X2 U7112 ( .A1(n6574), .A2(n6938), .ZN(n6462) );
  AOI22_X1 U7113 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6462), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6938), .ZN(n6428) );
  OAI21_X1 U7114 ( .B1(n6654), .B2(n6464), .A(n6428), .ZN(U3184) );
  AOI22_X1 U7115 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6462), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6952), .ZN(n6429) );
  OAI21_X1 U7116 ( .B1(n4828), .B2(n6464), .A(n6429), .ZN(U3185) );
  AOI22_X1 U7117 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6462), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6952), .ZN(n6430) );
  OAI21_X1 U7118 ( .B1(n6734), .B2(n6464), .A(n6430), .ZN(U3186) );
  INV_X1 U7119 ( .A(n6462), .ZN(n6469) );
  INV_X1 U7120 ( .A(n6464), .ZN(n6467) );
  AOI22_X1 U7121 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6467), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6952), .ZN(n6431) );
  OAI21_X1 U7122 ( .B1(n6734), .B2(n6469), .A(n6431), .ZN(U3187) );
  AOI22_X1 U7123 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6462), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6952), .ZN(n6432) );
  OAI21_X1 U7124 ( .B1(n6775), .B2(n6464), .A(n6432), .ZN(U3188) );
  AOI22_X1 U7125 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6462), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6952), .ZN(n6433) );
  OAI21_X1 U7126 ( .B1(n6435), .B2(n6464), .A(n6433), .ZN(U3189) );
  AOI22_X1 U7127 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6467), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6952), .ZN(n6434) );
  OAI21_X1 U7128 ( .B1(n6435), .B2(n6469), .A(n6434), .ZN(U3190) );
  AOI22_X1 U7129 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6462), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6952), .ZN(n6436) );
  OAI21_X1 U7130 ( .B1(n6438), .B2(n6464), .A(n6436), .ZN(U3191) );
  AOI22_X1 U7131 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6467), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6952), .ZN(n6437) );
  OAI21_X1 U7132 ( .B1(n6438), .B2(n6469), .A(n6437), .ZN(U3192) );
  AOI22_X1 U7133 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6462), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6952), .ZN(n6439) );
  OAI21_X1 U7134 ( .B1(n6441), .B2(n6464), .A(n6439), .ZN(U3193) );
  AOI22_X1 U7135 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6467), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6952), .ZN(n6440) );
  OAI21_X1 U7136 ( .B1(n6441), .B2(n6469), .A(n6440), .ZN(U3194) );
  AOI22_X1 U7137 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6462), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6952), .ZN(n6442) );
  OAI21_X1 U7138 ( .B1(n6601), .B2(n6464), .A(n6442), .ZN(U3195) );
  AOI22_X1 U7139 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6467), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6952), .ZN(n6443) );
  OAI21_X1 U7140 ( .B1(n6601), .B2(n6469), .A(n6443), .ZN(U3196) );
  INV_X1 U7141 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6446) );
  AOI22_X1 U7142 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6462), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6938), .ZN(n6444) );
  OAI21_X1 U7143 ( .B1(n6446), .B2(n6464), .A(n6444), .ZN(U3197) );
  AOI22_X1 U7144 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6467), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6952), .ZN(n6445) );
  OAI21_X1 U7145 ( .B1(n6446), .B2(n6469), .A(n6445), .ZN(U3198) );
  AOI22_X1 U7146 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6462), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6938), .ZN(n6447) );
  OAI21_X1 U7147 ( .B1(n6063), .B2(n6464), .A(n6447), .ZN(U3199) );
  AOI22_X1 U7148 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6467), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6952), .ZN(n6448) );
  OAI21_X1 U7149 ( .B1(n6063), .B2(n6469), .A(n6448), .ZN(U3200) );
  AOI22_X1 U7150 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6462), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6938), .ZN(n6449) );
  OAI21_X1 U7151 ( .B1(n6052), .B2(n6464), .A(n6449), .ZN(U3201) );
  AOI22_X1 U7152 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6467), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6952), .ZN(n6450) );
  OAI21_X1 U7153 ( .B1(n6052), .B2(n6469), .A(n6450), .ZN(U3202) );
  AOI22_X1 U7154 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6467), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6952), .ZN(n6451) );
  OAI21_X1 U7155 ( .B1(n6452), .B2(n6469), .A(n6451), .ZN(U3203) );
  AOI22_X1 U7156 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6462), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6938), .ZN(n6453) );
  OAI21_X1 U7157 ( .B1(n6454), .B2(n6464), .A(n6453), .ZN(U3204) );
  AOI22_X1 U7158 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6462), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6938), .ZN(n6455) );
  OAI21_X1 U7159 ( .B1(n6033), .B2(n6464), .A(n6455), .ZN(U3205) );
  AOI22_X1 U7160 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6467), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6952), .ZN(n6456) );
  OAI21_X1 U7161 ( .B1(n6033), .B2(n6469), .A(n6456), .ZN(U3206) );
  AOI22_X1 U7162 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6467), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6938), .ZN(n6457) );
  OAI21_X1 U7163 ( .B1(n6859), .B2(n6469), .A(n6457), .ZN(U3207) );
  AOI22_X1 U7164 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6462), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6938), .ZN(n6458) );
  OAI21_X1 U7165 ( .B1(n5998), .B2(n6464), .A(n6458), .ZN(U3208) );
  AOI22_X1 U7166 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6467), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6938), .ZN(n6459) );
  OAI21_X1 U7167 ( .B1(n5998), .B2(n6469), .A(n6459), .ZN(U3209) );
  AOI22_X1 U7168 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6467), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6938), .ZN(n6460) );
  OAI21_X1 U7169 ( .B1(n6461), .B2(n6469), .A(n6460), .ZN(U3210) );
  AOI22_X1 U7170 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6462), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6938), .ZN(n6463) );
  OAI21_X1 U7171 ( .B1(n6466), .B2(n6464), .A(n6463), .ZN(U3211) );
  AOI22_X1 U7172 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6467), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6938), .ZN(n6465) );
  OAI21_X1 U7173 ( .B1(n6466), .B2(n6469), .A(n6465), .ZN(U3212) );
  AOI22_X1 U7174 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6467), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6938), .ZN(n6468) );
  OAI21_X1 U7175 ( .B1(n6470), .B2(n6469), .A(n6468), .ZN(U3213) );
  MUX2_X1 U7176 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6955), .Z(U3445) );
  AOI221_X1 U7177 ( .B1(REIP_REG_0__SCAN_IN), .B2(REIP_REG_1__SCAN_IN), .C1(
        DATAWIDTH_REG_0__SCAN_IN), .C2(REIP_REG_1__SCAN_IN), .A(
        DATAWIDTH_REG_1__SCAN_IN), .ZN(n6481) );
  NOR4_X1 U7178 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(
        DATAWIDTH_REG_10__SCAN_IN), .ZN(n6474) );
  NOR4_X1 U7179 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6473) );
  NOR4_X1 U7180 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_2__SCAN_IN), .ZN(
        n6472) );
  NOR4_X1 U7181 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n6471) );
  NAND4_X1 U7182 ( .A1(n6474), .A2(n6473), .A3(n6472), .A4(n6471), .ZN(n6480)
         );
  NOR4_X1 U7183 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_27__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6478) );
  AOI211_X1 U7184 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_31__SCAN_IN), .B(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6477) );
  NOR4_X1 U7185 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6476) );
  NOR4_X1 U7186 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6475) );
  NAND4_X1 U7187 ( .A1(n6478), .A2(n6477), .A3(n6476), .A4(n6475), .ZN(n6479)
         );
  NOR2_X1 U7188 ( .A1(n6480), .A2(n6479), .ZN(n6491) );
  MUX2_X1 U7189 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(n6481), .S(n6491), .Z(
        U2795) );
  MUX2_X1 U7190 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6955), .Z(U3446) );
  AOI211_X1 U7191 ( .C1(REIP_REG_0__SCAN_IN), .C2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(REIP_REG_1__SCAN_IN), .B(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6482) );
  AOI21_X1 U7192 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6482), .ZN(n6484) );
  INV_X1 U7193 ( .A(n6491), .ZN(n6488) );
  AOI22_X1 U7194 ( .A1(n6491), .A2(n6484), .B1(n6483), .B2(n6488), .ZN(U3468)
         );
  MUX2_X1 U7195 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6955), .Z(U3447) );
  NOR3_X1 U7196 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6485) );
  NOR2_X1 U7197 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6485), .ZN(n6487) );
  AOI22_X1 U7198 ( .A1(n6491), .A2(n6487), .B1(n6486), .B2(n6488), .ZN(U2794)
         );
  MUX2_X1 U7199 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6955), .Z(U3448) );
  NOR2_X1 U7200 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6490) );
  AOI22_X1 U7201 ( .A1(n6491), .A2(n6490), .B1(n6489), .B2(n6488), .ZN(U3469)
         );
  INV_X1 U7202 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6497) );
  NAND2_X1 U7203 ( .A1(n6493), .A2(n6492), .ZN(n6494) );
  NAND2_X1 U7204 ( .A1(n6495), .A2(n6494), .ZN(n6774) );
  INV_X1 U7205 ( .A(n6774), .ZN(n6663) );
  AOI22_X1 U7206 ( .A1(n6779), .A2(n6508), .B1(n6507), .B2(n6663), .ZN(n6496)
         );
  OAI21_X1 U7207 ( .B1(n6510), .B2(n6497), .A(n6496), .ZN(U2852) );
  INV_X1 U7208 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6500) );
  INV_X1 U7209 ( .A(n6498), .ZN(n6967) );
  AOI22_X1 U7210 ( .A1(n6967), .A2(n6508), .B1(n6507), .B2(n6589), .ZN(n6499)
         );
  OAI21_X1 U7211 ( .B1(n6510), .B2(n6500), .A(n6499), .ZN(U2840) );
  AOI22_X1 U7212 ( .A1(n7060), .A2(n6508), .B1(n6507), .B2(n6863), .ZN(n6501)
         );
  OAI21_X1 U7213 ( .B1(n6510), .B2(n6502), .A(n6501), .ZN(U2835) );
  INV_X1 U7214 ( .A(EBX_REG_5__SCAN_IN), .ZN(n6746) );
  NOR2_X1 U7215 ( .A1(n6504), .A2(n6503), .ZN(n6505) );
  OR2_X1 U7216 ( .A1(n6506), .A2(n6505), .ZN(n6749) );
  INV_X1 U7217 ( .A(n6749), .ZN(n6642) );
  AOI22_X1 U7218 ( .A1(n6752), .A2(n6508), .B1(n6507), .B2(n6642), .ZN(n6509)
         );
  OAI21_X1 U7219 ( .B1(n6510), .B2(n6746), .A(n6509), .ZN(U2854) );
  AOI22_X1 U7220 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6560), .B1(n6789), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6516) );
  XNOR2_X1 U7221 ( .A(n6512), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6513)
         );
  XNOR2_X1 U7222 ( .A(n6511), .B(n6513), .ZN(n6658) );
  AOI22_X1 U7223 ( .A1(n6514), .A2(n6561), .B1(n6562), .B2(n6658), .ZN(n6515)
         );
  OAI211_X1 U7224 ( .C1(n6566), .C2(n6517), .A(n6516), .B(n6515), .ZN(U2984)
         );
  AOI22_X1 U7225 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n6560), .B1(n6789), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n6524) );
  OR2_X1 U7226 ( .A1(n6520), .A2(n6519), .ZN(n6521) );
  NAND2_X1 U7227 ( .A1(n6518), .A2(n6521), .ZN(n6621) );
  INV_X1 U7228 ( .A(n6621), .ZN(n6522) );
  AOI22_X1 U7229 ( .A1(n6522), .A2(n6562), .B1(n6561), .B2(n6742), .ZN(n6523)
         );
  OAI211_X1 U7230 ( .C1(n6566), .C2(n6745), .A(n6524), .B(n6523), .ZN(U2982)
         );
  AOI22_X1 U7231 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n6560), .B1(n6789), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n6530) );
  OAI21_X1 U7232 ( .B1(n6527), .B2(n6525), .A(n6526), .ZN(n6528) );
  INV_X1 U7233 ( .A(n6528), .ZN(n6643) );
  AOI22_X1 U7234 ( .A1(n6643), .A2(n6562), .B1(n6561), .B2(n6752), .ZN(n6529)
         );
  OAI211_X1 U7235 ( .C1(n6566), .C2(n6760), .A(n6530), .B(n6529), .ZN(U2981)
         );
  AOI22_X1 U7236 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6560), .B1(n6789), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n6537) );
  OAI21_X1 U7237 ( .B1(n6533), .B2(n6532), .A(n6531), .ZN(n6534) );
  INV_X1 U7238 ( .A(n6534), .ZN(n6636) );
  AOI22_X1 U7239 ( .A1(n6636), .A2(n6562), .B1(n6561), .B2(n6535), .ZN(n6536)
         );
  OAI211_X1 U7240 ( .C1(n6566), .C2(n6765), .A(n6537), .B(n6536), .ZN(U2980)
         );
  AOI22_X1 U7241 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n6560), .B1(n6789), 
        .B2(REIP_REG_7__SCAN_IN), .ZN(n6543) );
  OAI21_X1 U7242 ( .B1(n6540), .B2(n6539), .A(n3437), .ZN(n6541) );
  INV_X1 U7243 ( .A(n6541), .ZN(n6664) );
  AOI22_X1 U7244 ( .A1(n6664), .A2(n6562), .B1(n6561), .B2(n6779), .ZN(n6542)
         );
  OAI211_X1 U7245 ( .C1(n6566), .C2(n6784), .A(n6543), .B(n6542), .ZN(U2979)
         );
  OAI21_X1 U7246 ( .B1(n6546), .B2(n6545), .A(n6544), .ZN(n6692) );
  AOI22_X1 U7247 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6560), .B1(n6789), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n6551) );
  AOI22_X1 U7248 ( .A1(n6549), .A2(n6561), .B1(n6548), .B2(n6547), .ZN(n6550)
         );
  OAI211_X1 U7249 ( .C1(n6869), .C2(n6692), .A(n6551), .B(n6550), .ZN(U2975)
         );
  AOI22_X1 U7250 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n6560), .B1(n6789), 
        .B2(REIP_REG_13__SCAN_IN), .ZN(n6555) );
  XNOR2_X1 U7251 ( .A(n6552), .B(n6553), .ZN(n6604) );
  AOI22_X1 U7252 ( .A1(n6604), .A2(n6562), .B1(n6561), .B2(n6808), .ZN(n6554)
         );
  OAI211_X1 U7253 ( .C1(n6566), .C2(n6813), .A(n6555), .B(n6554), .ZN(U2973)
         );
  AOI22_X1 U7254 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n6560), .B1(n6789), 
        .B2(REIP_REG_18__SCAN_IN), .ZN(n6558) );
  AOI22_X1 U7255 ( .A1(n6556), .A2(n6562), .B1(n6561), .B2(n6959), .ZN(n6557)
         );
  OAI211_X1 U7256 ( .C1(n6566), .C2(n6559), .A(n6558), .B(n6557), .ZN(U2968)
         );
  AOI22_X1 U7257 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n6560), .B1(n6789), 
        .B2(REIP_REG_20__SCAN_IN), .ZN(n6565) );
  AOI22_X1 U7258 ( .A1(n6563), .A2(n6562), .B1(n6561), .B2(n6970), .ZN(n6564)
         );
  OAI211_X1 U7259 ( .C1(n6566), .C2(n6834), .A(n6565), .B(n6564), .ZN(U2966)
         );
  OAI21_X1 U7260 ( .B1(n6567), .B2(D_C_N_REG_SCAN_IN), .A(n6938), .ZN(n6568)
         );
  OAI21_X1 U7261 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6952), .A(n6568), .ZN(
        U2791) );
  NAND2_X1 U7262 ( .A1(n6583), .A2(n6569), .ZN(n6570) );
  OAI211_X1 U7263 ( .C1(n6583), .C2(n6572), .A(n6571), .B(n6570), .ZN(U3474)
         );
  AOI22_X1 U7264 ( .A1(n6955), .A2(READREQUEST_REG_SCAN_IN), .B1(n6573), .B2(
        n6938), .ZN(U3470) );
  NOR2_X1 U7265 ( .A1(n6574), .A2(n6935), .ZN(n6934) );
  NOR2_X1 U7266 ( .A1(n6944), .A2(n6937), .ZN(n6947) );
  AOI21_X1 U7267 ( .B1(HOLD), .B2(STATE_REG_1__SCAN_IN), .A(n6947), .ZN(n6576)
         );
  NAND2_X1 U7268 ( .A1(STATE_REG_1__SCAN_IN), .A2(READY_N), .ZN(n6948) );
  OAI211_X1 U7269 ( .C1(n6934), .C2(n6576), .A(n6575), .B(n6948), .ZN(U3182)
         );
  NAND2_X1 U7270 ( .A1(n6925), .A2(n6915), .ZN(n6578) );
  NAND2_X1 U7271 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6943), .ZN(n6909) );
  OAI221_X1 U7272 ( .B1(n6578), .B2(n6906), .C1(n6578), .C2(n6909), .A(n6577), 
        .ZN(U3150) );
  NAND2_X1 U7273 ( .A1(n6943), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6580) );
  AOI211_X1 U7274 ( .C1(n6581), .C2(n6930), .A(n6580), .B(n6579), .ZN(n6582)
         );
  OAI21_X1 U7275 ( .B1(n6582), .B2(n6923), .A(n6925), .ZN(n6587) );
  AOI211_X1 U7276 ( .C1(n6585), .C2(n6943), .A(n6584), .B(n6583), .ZN(n6586)
         );
  MUX2_X1 U7277 ( .A(n6587), .B(REQUESTPENDING_REG_SCAN_IN), .S(n6586), .Z(
        U3472) );
  AOI22_X1 U7278 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n6588), .B1(n6789), .B2(REIP_REG_19__SCAN_IN), .ZN(n6592) );
  AOI22_X1 U7279 ( .A1(n6590), .A2(n6723), .B1(n6721), .B2(n6589), .ZN(n6591)
         );
  OAI211_X1 U7280 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n6593), .A(n6592), .B(n6591), .ZN(U2999) );
  NOR2_X1 U7281 ( .A1(n6611), .A2(n6594), .ZN(n6596) );
  AOI21_X1 U7282 ( .B1(n6597), .B2(n6596), .A(n6595), .ZN(n6600) );
  NAND2_X1 U7283 ( .A1(n6727), .A2(n6597), .ZN(n6599) );
  AOI211_X1 U7284 ( .C1(n6600), .C2(n6599), .A(INSTADDRPOINTER_REG_13__SCAN_IN), .B(n6598), .ZN(n6603) );
  NOR2_X1 U7285 ( .A1(n6821), .A2(n6601), .ZN(n6602) );
  AOI211_X1 U7286 ( .C1(n6604), .C2(n6723), .A(n6603), .B(n6602), .ZN(n6608)
         );
  INV_X1 U7287 ( .A(n6806), .ZN(n6605) );
  AOI22_X1 U7288 ( .A1(n6606), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .B1(n6721), .B2(n6605), .ZN(n6607) );
  NAND2_X1 U7289 ( .A1(n6608), .A2(n6607), .ZN(U3005) );
  NAND2_X1 U7290 ( .A1(n6609), .A2(n6694), .ZN(n6619) );
  AOI21_X1 U7291 ( .B1(n6612), .B2(n6611), .A(n6610), .ZN(n6724) );
  NAND2_X1 U7292 ( .A1(n6721), .A2(n6613), .ZN(n6615) );
  OR2_X1 U7293 ( .A1(n6821), .A2(n5526), .ZN(n6614) );
  OAI211_X1 U7294 ( .C1(n6616), .C2(n6702), .A(n6615), .B(n6614), .ZN(n6617)
         );
  INV_X1 U7295 ( .A(n6617), .ZN(n6618) );
  OAI221_X1 U7296 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n6619), .C1(n4363), .C2(n6724), .A(n6618), .ZN(U3017) );
  INV_X1 U7297 ( .A(n6630), .ZN(n6628) );
  INV_X1 U7298 ( .A(n6640), .ZN(n6629) );
  AOI211_X1 U7299 ( .C1(n6627), .C2(n6620), .A(n6629), .B(n6639), .ZN(n6625)
         );
  NOR2_X1 U7300 ( .A1(n6621), .A2(n6702), .ZN(n6624) );
  NAND2_X1 U7301 ( .A1(n6721), .A2(n6736), .ZN(n6622) );
  OAI21_X1 U7302 ( .B1(n6734), .B2(n6821), .A(n6622), .ZN(n6623) );
  NOR3_X1 U7303 ( .A1(n6625), .A2(n6624), .A3(n6623), .ZN(n6626) );
  OAI21_X1 U7304 ( .B1(n6628), .B2(n6627), .A(n6626), .ZN(U3014) );
  NOR2_X1 U7305 ( .A1(n6629), .A2(n6674), .ZN(n6631) );
  AOI211_X1 U7306 ( .C1(n6632), .C2(n6633), .A(n6631), .B(n6630), .ZN(n6647)
         );
  OAI22_X1 U7307 ( .A1(n6709), .A2(n6761), .B1(n6775), .B2(n6821), .ZN(n6635)
         );
  NOR4_X1 U7308 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6633), .A3(n6640), 
        .A4(n6639), .ZN(n6634) );
  AOI211_X1 U7309 ( .C1(n6636), .C2(n6723), .A(n6635), .B(n6634), .ZN(n6637)
         );
  OAI21_X1 U7310 ( .B1(n6647), .B2(n6638), .A(n6637), .ZN(U3012) );
  NOR2_X1 U7311 ( .A1(n6640), .A2(n6639), .ZN(n6641) );
  NOR2_X1 U7312 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6641), .ZN(n6646)
         );
  AOI22_X1 U7313 ( .A1(n6643), .A2(n6723), .B1(n6721), .B2(n6642), .ZN(n6645)
         );
  NAND2_X1 U7314 ( .A1(n6789), .A2(REIP_REG_5__SCAN_IN), .ZN(n6644) );
  OAI211_X1 U7315 ( .C1(n6647), .C2(n6646), .A(n6645), .B(n6644), .ZN(U3013)
         );
  NAND2_X1 U7316 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6648), .ZN(n6662)
         );
  INV_X1 U7317 ( .A(n6649), .ZN(n6650) );
  NAND2_X1 U7318 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n6650), .ZN(n6652)
         );
  AOI21_X1 U7319 ( .B1(n6653), .B2(n6652), .A(n6651), .ZN(n6657) );
  OAI22_X1 U7320 ( .A1(n6709), .A2(n6655), .B1(n6654), .B2(n6821), .ZN(n6656)
         );
  AOI211_X1 U7321 ( .C1(n6723), .C2(n6658), .A(n6657), .B(n6656), .ZN(n6659)
         );
  OAI221_X1 U7322 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6662), .C1(n6661), .C2(n6660), .A(n6659), .ZN(U3016) );
  AOI22_X1 U7323 ( .A1(n6721), .A2(n6663), .B1(n6789), .B2(REIP_REG_7__SCAN_IN), .ZN(n6666) );
  AOI22_X1 U7324 ( .A1(n6664), .A2(n6723), .B1(n6668), .B2(n6667), .ZN(n6665)
         );
  OAI211_X1 U7325 ( .C1(n6667), .C2(n6672), .A(n6666), .B(n6665), .ZN(U3011)
         );
  NAND2_X1 U7326 ( .A1(n6673), .A2(n6668), .ZN(n6687) );
  AOI22_X1 U7327 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n5606), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6669), .ZN(n6678) );
  AOI21_X1 U7328 ( .B1(n6721), .B2(n6671), .A(n6670), .ZN(n6677) );
  OAI21_X1 U7329 ( .B1(n6674), .B2(n6673), .A(n6672), .ZN(n6683) );
  AOI22_X1 U7330 ( .A1(n6675), .A2(n6723), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6683), .ZN(n6676) );
  OAI211_X1 U7331 ( .C1(n6687), .C2(n6678), .A(n6677), .B(n6676), .ZN(U3008)
         );
  INV_X1 U7332 ( .A(n6679), .ZN(n6680) );
  AOI21_X1 U7333 ( .B1(n6721), .B2(n6681), .A(n6680), .ZN(n6686) );
  INV_X1 U7334 ( .A(n6682), .ZN(n6684) );
  AOI22_X1 U7335 ( .A1(n6684), .A2(n6723), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6683), .ZN(n6685) );
  OAI211_X1 U7336 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6687), .A(n6686), 
        .B(n6685), .ZN(U3009) );
  AOI22_X1 U7337 ( .A1(n6721), .A2(n6688), .B1(n6789), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n6691) );
  INV_X1 U7338 ( .A(n6717), .ZN(n6689) );
  AOI22_X1 U7339 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6693), .B1(n6689), .B2(n5609), .ZN(n6690) );
  OAI211_X1 U7340 ( .C1(n6702), .C2(n6692), .A(n6691), .B(n6690), .ZN(U3007)
         );
  OR2_X1 U7341 ( .A1(n6717), .A2(n6695), .ZN(n6699) );
  AOI21_X1 U7342 ( .B1(n6695), .B2(n6694), .A(n6693), .ZN(n6708) );
  AOI222_X1 U7343 ( .A1(n6697), .A2(n6723), .B1(n6721), .B2(n6696), .C1(
        REIP_REG_15__SCAN_IN), .C2(n6789), .ZN(n6698) );
  OAI221_X1 U7344 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n6699), .C1(
        n6700), .C2(n6708), .A(n6698), .ZN(U3003) );
  AOI221_X1 U7345 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .C1(n6707), .C2(n6700), .A(n6699), 
        .ZN(n6705) );
  OAI22_X1 U7346 ( .A1(n6703), .A2(n6702), .B1(n6709), .B2(n6701), .ZN(n6704)
         );
  AOI211_X1 U7347 ( .C1(REIP_REG_16__SCAN_IN), .C2(n6789), .A(n6705), .B(n6704), .ZN(n6706) );
  OAI21_X1 U7348 ( .B1(n6708), .B2(n6707), .A(n6706), .ZN(U3002) );
  OAI22_X1 U7349 ( .A1(n6711), .A2(n6710), .B1(n6814), .B2(n6709), .ZN(n6712)
         );
  AOI21_X1 U7350 ( .B1(n6713), .B2(n6723), .A(n6712), .ZN(n6715) );
  NAND2_X1 U7351 ( .A1(n6789), .A2(REIP_REG_17__SCAN_IN), .ZN(n6714) );
  OAI211_X1 U7352 ( .C1(n6717), .C2(n6716), .A(n6715), .B(n6714), .ZN(U3001)
         );
  INV_X1 U7353 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6730) );
  INV_X1 U7354 ( .A(n6718), .ZN(n6722) );
  INV_X1 U7355 ( .A(n6719), .ZN(n6720) );
  AOI22_X1 U7356 ( .A1(n6723), .A2(n6722), .B1(n6721), .B2(n6720), .ZN(n6729)
         );
  INV_X1 U7357 ( .A(n6724), .ZN(n6726) );
  OAI22_X1 U7358 ( .A1(n6727), .A2(n6726), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6725), .ZN(n6728) );
  OAI211_X1 U7359 ( .C1(n6730), .C2(n6821), .A(n6729), .B(n6728), .ZN(U3018)
         );
  OAI22_X1 U7360 ( .A1(n6734), .A2(n6733), .B1(n6732), .B2(n6731), .ZN(n6735)
         );
  AOI211_X1 U7361 ( .C1(n6856), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6789), 
        .B(n6735), .ZN(n6744) );
  INV_X1 U7362 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6740) );
  NAND2_X1 U7363 ( .A1(n6864), .A2(n6736), .ZN(n6739) );
  OR3_X1 U7364 ( .A1(n6802), .A2(n6737), .A3(REIP_REG_4__SCAN_IN), .ZN(n6738)
         );
  OAI211_X1 U7365 ( .C1(n6740), .C2(n6796), .A(n6739), .B(n6738), .ZN(n6741)
         );
  AOI21_X1 U7366 ( .B1(n6742), .B2(n6751), .A(n6741), .ZN(n6743) );
  OAI211_X1 U7367 ( .C1(n6745), .C2(n6833), .A(n6744), .B(n6743), .ZN(U2823)
         );
  NOR2_X1 U7368 ( .A1(n6796), .A2(n6746), .ZN(n6747) );
  AOI211_X1 U7369 ( .C1(n6856), .C2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n6789), 
        .B(n6747), .ZN(n6748) );
  OAI21_X1 U7370 ( .B1(n6847), .B2(n6749), .A(n6748), .ZN(n6750) );
  AOI21_X1 U7371 ( .B1(n6752), .B2(n6751), .A(n6750), .ZN(n6759) );
  INV_X1 U7372 ( .A(n6753), .ZN(n6754) );
  NOR2_X1 U7373 ( .A1(n6802), .A2(n6754), .ZN(n6764) );
  INV_X1 U7374 ( .A(n6755), .ZN(n6757) );
  OAI21_X1 U7375 ( .B1(n6802), .B2(n6757), .A(n6756), .ZN(n6780) );
  OAI21_X1 U7376 ( .B1(n6764), .B2(REIP_REG_5__SCAN_IN), .A(n6780), .ZN(n6758)
         );
  OAI211_X1 U7377 ( .C1(n6833), .C2(n6760), .A(n6759), .B(n6758), .ZN(U2822)
         );
  OAI22_X1 U7378 ( .A1(n6762), .A2(n6796), .B1(n6847), .B2(n6761), .ZN(n6763)
         );
  AOI211_X1 U7379 ( .C1(n6856), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6789), 
        .B(n6763), .ZN(n6769) );
  NAND2_X1 U7380 ( .A1(n6764), .A2(REIP_REG_5__SCAN_IN), .ZN(n6776) );
  NOR2_X1 U7381 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6776), .ZN(n6781) );
  OAI22_X1 U7382 ( .A1(n6766), .A2(n6827), .B1(n6765), .B2(n6833), .ZN(n6767)
         );
  AOI211_X1 U7383 ( .C1(REIP_REG_6__SCAN_IN), .C2(n6780), .A(n6781), .B(n6767), 
        .ZN(n6768) );
  NAND2_X1 U7384 ( .A1(n6769), .A2(n6768), .ZN(U2821) );
  INV_X1 U7385 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6771) );
  NAND2_X1 U7386 ( .A1(n6855), .A2(EBX_REG_7__SCAN_IN), .ZN(n6770) );
  OAI211_X1 U7387 ( .C1(n6771), .C2(n6854), .A(n6770), .B(n6821), .ZN(n6772)
         );
  INV_X1 U7388 ( .A(n6772), .ZN(n6773) );
  OAI21_X1 U7389 ( .B1(n6847), .B2(n6774), .A(n6773), .ZN(n6778) );
  NOR3_X1 U7390 ( .A1(n6776), .A2(n6775), .A3(REIP_REG_7__SCAN_IN), .ZN(n6777)
         );
  AOI211_X1 U7391 ( .C1(n6779), .C2(n6865), .A(n6778), .B(n6777), .ZN(n6783)
         );
  OAI21_X1 U7392 ( .B1(n6781), .B2(n6780), .A(REIP_REG_7__SCAN_IN), .ZN(n6782)
         );
  OAI211_X1 U7393 ( .C1(n6833), .C2(n6784), .A(n6783), .B(n6782), .ZN(U2820)
         );
  INV_X1 U7394 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6797) );
  AOI21_X1 U7395 ( .B1(REIP_REG_9__SCAN_IN), .B2(n6786), .A(n6785), .ZN(n6795)
         );
  NOR2_X1 U7396 ( .A1(n6847), .A2(n6787), .ZN(n6788) );
  AOI211_X1 U7397 ( .C1(n6856), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6789), 
        .B(n6788), .ZN(n6790) );
  OAI21_X1 U7398 ( .B1(n6791), .B2(n6827), .A(n6790), .ZN(n6792) );
  AOI21_X1 U7399 ( .B1(n6793), .B2(n6861), .A(n6792), .ZN(n6794) );
  OAI211_X1 U7400 ( .C1(n6797), .C2(n6796), .A(n6795), .B(n6794), .ZN(U2818)
         );
  INV_X1 U7401 ( .A(n6798), .ZN(n6799) );
  NAND2_X1 U7402 ( .A1(n6601), .A2(n6799), .ZN(n6801) );
  NAND2_X1 U7403 ( .A1(n6856), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6800)
         );
  OAI211_X1 U7404 ( .C1(n6802), .C2(n6801), .A(n6821), .B(n6800), .ZN(n6803)
         );
  INV_X1 U7405 ( .A(n6803), .ZN(n6805) );
  NAND2_X1 U7406 ( .A1(n6855), .A2(EBX_REG_13__SCAN_IN), .ZN(n6804) );
  OAI211_X1 U7407 ( .C1(n6847), .C2(n6806), .A(n6805), .B(n6804), .ZN(n6807)
         );
  AOI21_X1 U7408 ( .B1(n6808), .B2(n6865), .A(n6807), .ZN(n6812) );
  OAI21_X1 U7409 ( .B1(n6810), .B2(n6809), .A(REIP_REG_13__SCAN_IN), .ZN(n6811) );
  OAI211_X1 U7410 ( .C1(n6833), .C2(n6813), .A(n6812), .B(n6811), .ZN(U2814)
         );
  AOI22_X1 U7411 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n6856), .B1(
        EBX_REG_17__SCAN_IN), .B2(n6855), .ZN(n6823) );
  OAI22_X1 U7412 ( .A1(n6815), .A2(n6827), .B1(n6847), .B2(n6814), .ZN(n6816)
         );
  AOI21_X1 U7413 ( .B1(n6817), .B2(n6861), .A(n6816), .ZN(n6822) );
  OAI21_X1 U7414 ( .B1(REIP_REG_17__SCAN_IN), .B2(n6819), .A(n6818), .ZN(n6820) );
  NAND4_X1 U7415 ( .A1(n6823), .A2(n6822), .A3(n6821), .A4(n6820), .ZN(U2810)
         );
  AOI22_X1 U7416 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n6856), .B1(
        EBX_REG_20__SCAN_IN), .B2(n6855), .ZN(n6832) );
  NOR2_X1 U7417 ( .A1(n6825), .A2(n6824), .ZN(n6836) );
  OAI22_X1 U7418 ( .A1(n6828), .A2(n6827), .B1(n6826), .B2(n6847), .ZN(n6829)
         );
  AOI221_X1 U7419 ( .B1(REIP_REG_20__SCAN_IN), .B2(n6836), .C1(n6830), .C2(
        n6836), .A(n6829), .ZN(n6831) );
  OAI211_X1 U7420 ( .C1(n6834), .C2(n6833), .A(n6832), .B(n6831), .ZN(U2807)
         );
  AOI22_X1 U7421 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n6856), .B1(n6835), 
        .B2(n6861), .ZN(n6842) );
  AOI22_X1 U7422 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6855), .B1(
        REIP_REG_21__SCAN_IN), .B2(n6836), .ZN(n6841) );
  AOI22_X1 U7423 ( .A1(n6973), .A2(n6865), .B1(n6837), .B2(n6864), .ZN(n6840)
         );
  OR2_X1 U7424 ( .A1(n6838), .A2(REIP_REG_21__SCAN_IN), .ZN(n6839) );
  NAND4_X1 U7425 ( .A1(n6842), .A2(n6841), .A3(n6840), .A4(n6839), .ZN(U2806)
         );
  AOI22_X1 U7426 ( .A1(n6843), .A2(n6861), .B1(EBX_REG_23__SCAN_IN), .B2(n6855), .ZN(n6853) );
  NOR2_X1 U7427 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6844), .ZN(n6849) );
  NAND2_X1 U7428 ( .A1(n6846), .A2(n6845), .ZN(n6858) );
  OAI22_X1 U7429 ( .A1(n6849), .A2(n6858), .B1(n6848), .B2(n6847), .ZN(n6850)
         );
  AOI21_X1 U7430 ( .B1(n6851), .B2(n6865), .A(n6850), .ZN(n6852) );
  OAI211_X1 U7431 ( .C1(n4157), .C2(n6854), .A(n6853), .B(n6852), .ZN(U2804)
         );
  AOI22_X1 U7432 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n6856), .B1(
        EBX_REG_24__SCAN_IN), .B2(n6855), .ZN(n6857) );
  OAI21_X1 U7433 ( .B1(n6859), .B2(n6858), .A(n6857), .ZN(n6860) );
  AOI21_X1 U7434 ( .B1(n6862), .B2(n6861), .A(n6860), .ZN(n6867) );
  AOI22_X1 U7435 ( .A1(n7060), .A2(n6865), .B1(n6864), .B2(n6863), .ZN(n6866)
         );
  OAI211_X1 U7436 ( .C1(REIP_REG_24__SCAN_IN), .C2(n6868), .A(n6867), .B(n6866), .ZN(U2803) );
  OAI21_X1 U7437 ( .B1(n6870), .B2(n6894), .A(n6869), .ZN(U2793) );
  INV_X1 U7438 ( .A(n6871), .ZN(n6872) );
  NAND3_X1 U7439 ( .A1(n6873), .A2(n6872), .A3(n6916), .ZN(n6874) );
  OAI21_X1 U7440 ( .B1(n6875), .B2(n3846), .A(n6874), .ZN(U3455) );
  INV_X1 U7441 ( .A(n6886), .ZN(n6884) );
  NOR3_X1 U7442 ( .A1(n6877), .A2(n7025), .A3(n6876), .ZN(n6878) );
  NAND2_X1 U7443 ( .A1(n6878), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6882) );
  OAI22_X1 U7444 ( .A1(n6880), .A2(n6879), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6878), .ZN(n6881) );
  OAI211_X1 U7445 ( .C1(n6884), .C2(n6883), .A(n6882), .B(n6881), .ZN(n6885)
         );
  OAI21_X1 U7446 ( .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6886), .A(n6885), 
        .ZN(n6887) );
  AOI222_X1 U7447 ( .A1(n6889), .A2(n6888), .B1(n6889), .B2(n6887), .C1(n6888), 
        .C2(n6887), .ZN(n6901) );
  INV_X1 U7448 ( .A(n6890), .ZN(n6900) );
  INV_X1 U7449 ( .A(n6891), .ZN(n6897) );
  INV_X1 U7450 ( .A(MORE_REG_SCAN_IN), .ZN(n6893) );
  AOI21_X1 U7451 ( .B1(n6894), .B2(n6893), .A(n6892), .ZN(n6896) );
  NOR4_X1 U7452 ( .A1(n6898), .A2(n6897), .A3(n6896), .A4(n6895), .ZN(n6899)
         );
  OAI211_X1 U7453 ( .C1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n6901), .A(n6900), .B(n6899), .ZN(n6917) );
  OAI22_X1 U7454 ( .A1(n6917), .A2(n6928), .B1(n6902), .B2(n6943), .ZN(n6903)
         );
  OAI21_X1 U7455 ( .B1(n6905), .B2(n6904), .A(n6903), .ZN(n6922) );
  NAND2_X1 U7456 ( .A1(n6906), .A2(READY_N), .ZN(n6907) );
  AOI21_X1 U7457 ( .B1(n6922), .B2(n6907), .A(n6923), .ZN(n6918) );
  AOI21_X1 U7458 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n6918), .A(n6908), .ZN(
        n6913) );
  OAI21_X1 U7459 ( .B1(n6910), .B2(n6909), .A(n6928), .ZN(n6911) );
  NAND2_X1 U7460 ( .A1(n6922), .A2(n6911), .ZN(n6912) );
  OAI211_X1 U7461 ( .C1(n6914), .C2(n6922), .A(n6913), .B(n6912), .ZN(U3149)
         );
  OAI221_X1 U7462 ( .B1(n6916), .B2(STATE2_REG_0__SCAN_IN), .C1(n6916), .C2(
        n6922), .A(n6915), .ZN(U3453) );
  INV_X1 U7463 ( .A(n6917), .ZN(n6929) );
  AOI211_X1 U7464 ( .C1(n6921), .C2(n6920), .A(n6919), .B(n6918), .ZN(n6927)
         );
  OAI211_X1 U7465 ( .C1(n6925), .C2(n6924), .A(n6923), .B(n6922), .ZN(n6926)
         );
  OAI211_X1 U7466 ( .C1(n6929), .C2(n6928), .A(n6927), .B(n6926), .ZN(U3148)
         );
  OAI21_X1 U7467 ( .B1(n6933), .B2(n6930), .A(n6931), .ZN(U2792) );
  INV_X1 U7468 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6932) );
  OAI21_X1 U7469 ( .B1(n6933), .B2(n6932), .A(n6931), .ZN(U3452) );
  INV_X1 U7470 ( .A(n6934), .ZN(n6941) );
  INV_X1 U7471 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6936) );
  NOR2_X1 U7472 ( .A1(n6936), .A2(n6935), .ZN(n6939) );
  AOI221_X1 U7473 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6946), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6950) );
  AOI221_X1 U7474 ( .B1(n6939), .B2(n6938), .C1(n6937), .C2(n6938), .A(n6950), 
        .ZN(n6940) );
  OAI221_X1 U7475 ( .B1(n6942), .B2(n6948), .C1(n6942), .C2(n6941), .A(n6940), 
        .ZN(U3181) );
  AOI221_X1 U7476 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6943), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6945) );
  AOI221_X1 U7477 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6945), .C2(HOLD), .A(n6944), .ZN(n6951) );
  AOI21_X1 U7478 ( .B1(n6947), .B2(n6946), .A(STATE_REG_2__SCAN_IN), .ZN(n6949) );
  OAI22_X1 U7479 ( .A1(n6951), .A2(n6950), .B1(n6949), .B2(n6948), .ZN(U3183)
         );
  INV_X1 U7480 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6953) );
  AOI22_X1 U7481 ( .A1(n6955), .A2(n6954), .B1(n6953), .B2(n6952), .ZN(U3473)
         );
  AOI22_X1 U7482 ( .A1(n6956), .A2(n7078), .B1(n7077), .B2(DATAI_16_), .ZN(
        n6958) );
  AOI22_X1 U7483 ( .A1(n7081), .A2(DATAI_0_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n7080), .ZN(n6957) );
  NAND2_X1 U7484 ( .A1(n6958), .A2(n6957), .ZN(U2875) );
  AOI22_X1 U7485 ( .A1(n6959), .A2(n7078), .B1(n7077), .B2(DATAI_18_), .ZN(
        n6966) );
  INV_X1 U7486 ( .A(DATAI_2_), .ZN(n6962) );
  OAI22_X1 U7487 ( .A1(n6963), .A2(n6962), .B1(n6961), .B2(n3422), .ZN(n6964)
         );
  INV_X1 U7488 ( .A(n6964), .ZN(n6965) );
  NAND2_X1 U7489 ( .A1(n6966), .A2(n6965), .ZN(U2873) );
  AOI22_X1 U7490 ( .A1(n6967), .A2(n7078), .B1(n7077), .B2(DATAI_19_), .ZN(
        n6969) );
  AOI22_X1 U7491 ( .A1(n7081), .A2(DATAI_3_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n7080), .ZN(n6968) );
  NAND2_X1 U7492 ( .A1(n6969), .A2(n6968), .ZN(U2872) );
  AOI22_X1 U7493 ( .A1(n6970), .A2(n7078), .B1(n7077), .B2(DATAI_20_), .ZN(
        n6972) );
  AOI22_X1 U7494 ( .A1(n7081), .A2(DATAI_4_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n7080), .ZN(n6971) );
  NAND2_X1 U7495 ( .A1(n6972), .A2(n6971), .ZN(U2871) );
  AOI22_X1 U7496 ( .A1(n6973), .A2(n7078), .B1(n7077), .B2(DATAI_21_), .ZN(
        n6975) );
  AOI22_X1 U7497 ( .A1(n7081), .A2(DATAI_5_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n7080), .ZN(n6974) );
  NAND2_X1 U7498 ( .A1(n6975), .A2(n6974), .ZN(U2870) );
  INV_X1 U7499 ( .A(n6976), .ZN(n6977) );
  AOI22_X1 U7500 ( .A1(n6977), .A2(n7078), .B1(n7077), .B2(DATAI_22_), .ZN(
        n6979) );
  AOI22_X1 U7501 ( .A1(n7081), .A2(DATAI_6_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n7080), .ZN(n6978) );
  NAND2_X1 U7502 ( .A1(n6979), .A2(n6978), .ZN(U2869) );
  NOR2_X1 U7503 ( .A1(n6980), .A2(n7052), .ZN(n6984) );
  NOR2_X1 U7504 ( .A1(n7025), .A2(n6981), .ZN(n7155) );
  AOI21_X1 U7505 ( .B1(n6982), .B2(n7022), .A(n7155), .ZN(n6985) );
  INV_X1 U7506 ( .A(n6985), .ZN(n6983) );
  AOI22_X1 U7507 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6987), .B1(n6984), .B2(
        n6983), .ZN(n7160) );
  AOI22_X1 U7508 ( .A1(n7156), .A2(n7056), .B1(n7047), .B2(n7155), .ZN(n6989)
         );
  AOI21_X1 U7509 ( .B1(n6985), .B2(n6984), .A(n7050), .ZN(n6986) );
  OAI21_X1 U7510 ( .B1(n7031), .B2(n6987), .A(n6986), .ZN(n7157) );
  AOI22_X1 U7511 ( .A1(n7157), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n7048), 
        .B2(n7154), .ZN(n6988) );
  OAI211_X1 U7512 ( .C1(n7160), .C2(n7059), .A(n6989), .B(n6988), .ZN(U3124)
         );
  NAND2_X1 U7513 ( .A1(n7011), .A2(n6990), .ZN(n6997) );
  NOR2_X1 U7514 ( .A1(n7162), .A2(n7052), .ZN(n6992) );
  AOI21_X1 U7515 ( .B1(n6997), .B2(n6992), .A(n6991), .ZN(n7004) );
  INV_X1 U7516 ( .A(n7004), .ZN(n6996) );
  INV_X1 U7517 ( .A(n6993), .ZN(n6995) );
  AOI22_X1 U7518 ( .A1(n6996), .A2(n7003), .B1(n6995), .B2(n6994), .ZN(n7166)
         );
  NOR2_X1 U7519 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6998), .ZN(n7161)
         );
  AOI22_X1 U7520 ( .A1(n7168), .A2(n7056), .B1(n7047), .B2(n7161), .ZN(n7006)
         );
  INV_X1 U7521 ( .A(n7161), .ZN(n7001) );
  AOI211_X1 U7522 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n7001), .A(n7000), .B(
        n6999), .ZN(n7002) );
  OAI21_X1 U7523 ( .B1(n7004), .B2(n7003), .A(n7002), .ZN(n7163) );
  AOI22_X1 U7524 ( .A1(n7163), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n7048), 
        .B2(n7162), .ZN(n7005) );
  OAI211_X1 U7525 ( .C1(n7166), .C2(n7059), .A(n7006), .B(n7005), .ZN(U3100)
         );
  OR2_X1 U7526 ( .A1(n7008), .A2(n7007), .ZN(n7010) );
  NOR2_X1 U7527 ( .A1(n7025), .A2(n7015), .ZN(n7167) );
  INV_X1 U7528 ( .A(n7167), .ZN(n7009) );
  NAND2_X1 U7529 ( .A1(n7010), .A2(n7009), .ZN(n7017) );
  AOI21_X1 U7530 ( .B1(n7011), .B2(STATEBS16_REG_SCAN_IN), .A(n7052), .ZN(
        n7014) );
  AOI22_X1 U7531 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7012), .B1(n7017), .B2(
        n7014), .ZN(n7173) );
  AOI22_X1 U7532 ( .A1(n7169), .A2(n7056), .B1(n7047), .B2(n7167), .ZN(n7020)
         );
  INV_X1 U7533 ( .A(n7014), .ZN(n7018) );
  AOI21_X1 U7534 ( .B1(n7052), .B2(n7015), .A(n7050), .ZN(n7016) );
  OAI21_X1 U7535 ( .B1(n7018), .B2(n7017), .A(n7016), .ZN(n7170) );
  AOI22_X1 U7536 ( .A1(n7170), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n7048), 
        .B2(n7168), .ZN(n7019) );
  OAI211_X1 U7537 ( .C1(n7173), .C2(n7059), .A(n7020), .B(n7019), .ZN(U3092)
         );
  NOR2_X1 U7538 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n7024), .ZN(n7030)
         );
  OAI21_X1 U7539 ( .B1(n7021), .B2(n7052), .A(n7039), .ZN(n7033) );
  NAND2_X1 U7540 ( .A1(n7023), .A2(n7022), .ZN(n7027) );
  NOR3_X2 U7541 ( .A1(n7025), .A2(n7024), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n7174) );
  INV_X1 U7542 ( .A(n7174), .ZN(n7026) );
  NAND2_X1 U7543 ( .A1(n7027), .A2(n7026), .ZN(n7028) );
  AOI22_X1 U7544 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7030), .B1(n7033), .B2(
        n7028), .ZN(n7180) );
  AOI22_X1 U7545 ( .A1(n7176), .A2(n7056), .B1(n7047), .B2(n7174), .ZN(n7038)
         );
  INV_X1 U7546 ( .A(n7028), .ZN(n7034) );
  OAI21_X1 U7547 ( .B1(n7031), .B2(n7030), .A(n7029), .ZN(n7032) );
  AOI21_X1 U7548 ( .B1(n7034), .B2(n7033), .A(n7032), .ZN(n7035) );
  AOI22_X1 U7549 ( .A1(n7177), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n7048), 
        .B2(n7175), .ZN(n7037) );
  OAI211_X1 U7550 ( .C1(n7180), .C2(n7059), .A(n7038), .B(n7037), .ZN(U3060)
         );
  INV_X1 U7551 ( .A(n7051), .ZN(n7045) );
  OAI21_X1 U7552 ( .B1(n7040), .B2(n7052), .A(n7039), .ZN(n7049) );
  NAND2_X1 U7553 ( .A1(n7042), .A2(n7041), .ZN(n7046) );
  OAI21_X1 U7554 ( .B1(n7044), .B2(n7043), .A(n7046), .ZN(n7054) );
  AOI22_X1 U7555 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7045), .B1(n7049), .B2(
        n7054), .ZN(n7191) );
  INV_X1 U7556 ( .A(n7046), .ZN(n7181) );
  AOI22_X1 U7557 ( .A1(n7185), .A2(n7048), .B1(n7047), .B2(n7181), .ZN(n7058)
         );
  INV_X1 U7558 ( .A(n7049), .ZN(n7055) );
  AOI21_X1 U7559 ( .B1(n7052), .B2(n7051), .A(n7050), .ZN(n7053) );
  OAI21_X1 U7560 ( .B1(n7055), .B2(n7054), .A(n7053), .ZN(n7187) );
  AOI22_X1 U7561 ( .A1(n7187), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n7056), 
        .B2(n7184), .ZN(n7057) );
  OAI211_X1 U7562 ( .C1(n7191), .C2(n7059), .A(n7058), .B(n7057), .ZN(U3044)
         );
  AOI22_X1 U7563 ( .A1(n7060), .A2(n7078), .B1(n7077), .B2(DATAI_24_), .ZN(
        n7062) );
  AOI22_X1 U7564 ( .A1(n7081), .A2(DATAI_8_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n7080), .ZN(n7061) );
  NAND2_X1 U7565 ( .A1(n7062), .A2(n7061), .ZN(U2867) );
  AOI22_X1 U7566 ( .A1(n7156), .A2(n7072), .B1(n7071), .B2(n7155), .ZN(n7064)
         );
  AOI22_X1 U7567 ( .A1(n7157), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n7073), 
        .B2(n7154), .ZN(n7063) );
  OAI211_X1 U7568 ( .C1(n7160), .C2(n7076), .A(n7064), .B(n7063), .ZN(U3125)
         );
  AOI22_X1 U7569 ( .A1(n7168), .A2(n7072), .B1(n7071), .B2(n7161), .ZN(n7066)
         );
  AOI22_X1 U7570 ( .A1(n7163), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n7073), 
        .B2(n7162), .ZN(n7065) );
  OAI211_X1 U7571 ( .C1(n7166), .C2(n7076), .A(n7066), .B(n7065), .ZN(U3101)
         );
  AOI22_X1 U7572 ( .A1(n7169), .A2(n7072), .B1(n7071), .B2(n7167), .ZN(n7068)
         );
  AOI22_X1 U7573 ( .A1(n7170), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n7073), 
        .B2(n7168), .ZN(n7067) );
  OAI211_X1 U7574 ( .C1(n7173), .C2(n7076), .A(n7068), .B(n7067), .ZN(U3093)
         );
  AOI22_X1 U7575 ( .A1(n7175), .A2(n7073), .B1(n7071), .B2(n7174), .ZN(n7070)
         );
  AOI22_X1 U7576 ( .A1(n7177), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n7072), 
        .B2(n7176), .ZN(n7069) );
  OAI211_X1 U7577 ( .C1(n7180), .C2(n7076), .A(n7070), .B(n7069), .ZN(U3061)
         );
  AOI22_X1 U7578 ( .A1(n7184), .A2(n7072), .B1(n7071), .B2(n7181), .ZN(n7075)
         );
  AOI22_X1 U7579 ( .A1(n7187), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n7073), 
        .B2(n7185), .ZN(n7074) );
  OAI211_X1 U7580 ( .C1(n7191), .C2(n7076), .A(n7075), .B(n7074), .ZN(U3045)
         );
  AOI22_X1 U7581 ( .A1(n7079), .A2(n7078), .B1(n7077), .B2(DATAI_25_), .ZN(
        n7083) );
  AOI22_X1 U7582 ( .A1(n7081), .A2(DATAI_9_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n7080), .ZN(n7082) );
  NAND2_X1 U7583 ( .A1(n7083), .A2(n7082), .ZN(U2866) );
  AOI22_X1 U7584 ( .A1(n7092), .A2(n7155), .B1(n7154), .B2(n7093), .ZN(n7085)
         );
  AOI22_X1 U7585 ( .A1(n7157), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n7094), 
        .B2(n7156), .ZN(n7084) );
  OAI211_X1 U7586 ( .C1(n7160), .C2(n7097), .A(n7085), .B(n7084), .ZN(U3126)
         );
  AOI22_X1 U7587 ( .A1(n7168), .A2(n7094), .B1(n7092), .B2(n7161), .ZN(n7087)
         );
  AOI22_X1 U7588 ( .A1(n7163), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n7093), 
        .B2(n7162), .ZN(n7086) );
  OAI211_X1 U7589 ( .C1(n7166), .C2(n7097), .A(n7087), .B(n7086), .ZN(U3102)
         );
  AOI22_X1 U7590 ( .A1(n7169), .A2(n7094), .B1(n7092), .B2(n7167), .ZN(n7089)
         );
  AOI22_X1 U7591 ( .A1(n7170), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n7093), 
        .B2(n7168), .ZN(n7088) );
  OAI211_X1 U7592 ( .C1(n7173), .C2(n7097), .A(n7089), .B(n7088), .ZN(U3094)
         );
  AOI22_X1 U7593 ( .A1(n7175), .A2(n7093), .B1(n7092), .B2(n7174), .ZN(n7091)
         );
  AOI22_X1 U7594 ( .A1(n7177), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n7094), 
        .B2(n7176), .ZN(n7090) );
  OAI211_X1 U7595 ( .C1(n7180), .C2(n7097), .A(n7091), .B(n7090), .ZN(U3062)
         );
  AOI22_X1 U7596 ( .A1(n7185), .A2(n7093), .B1(n7092), .B2(n7181), .ZN(n7096)
         );
  AOI22_X1 U7597 ( .A1(n7187), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n7094), 
        .B2(n7184), .ZN(n7095) );
  OAI211_X1 U7598 ( .C1(n7191), .C2(n7097), .A(n7096), .B(n7095), .ZN(U3046)
         );
  AOI22_X1 U7599 ( .A1(n7106), .A2(n7155), .B1(n7154), .B2(n7107), .ZN(n7099)
         );
  AOI22_X1 U7600 ( .A1(n7157), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n7108), 
        .B2(n7156), .ZN(n7098) );
  OAI211_X1 U7601 ( .C1(n7160), .C2(n7111), .A(n7099), .B(n7098), .ZN(U3127)
         );
  AOI22_X1 U7602 ( .A1(n7168), .A2(n7108), .B1(n7106), .B2(n7161), .ZN(n7101)
         );
  AOI22_X1 U7603 ( .A1(n7163), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n7107), 
        .B2(n7162), .ZN(n7100) );
  OAI211_X1 U7604 ( .C1(n7166), .C2(n7111), .A(n7101), .B(n7100), .ZN(U3103)
         );
  AOI22_X1 U7605 ( .A1(n7169), .A2(n7108), .B1(n7106), .B2(n7167), .ZN(n7103)
         );
  AOI22_X1 U7606 ( .A1(n7170), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n7107), 
        .B2(n7168), .ZN(n7102) );
  OAI211_X1 U7607 ( .C1(n7173), .C2(n7111), .A(n7103), .B(n7102), .ZN(U3095)
         );
  AOI22_X1 U7608 ( .A1(n7176), .A2(n7108), .B1(n7106), .B2(n7174), .ZN(n7105)
         );
  AOI22_X1 U7609 ( .A1(n7177), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n7107), 
        .B2(n7175), .ZN(n7104) );
  OAI211_X1 U7610 ( .C1(n7180), .C2(n7111), .A(n7105), .B(n7104), .ZN(U3063)
         );
  AOI22_X1 U7611 ( .A1(n7185), .A2(n7107), .B1(n7106), .B2(n7181), .ZN(n7110)
         );
  AOI22_X1 U7612 ( .A1(n7187), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n7108), 
        .B2(n7184), .ZN(n7109) );
  OAI211_X1 U7613 ( .C1(n7191), .C2(n7111), .A(n7110), .B(n7109), .ZN(U3047)
         );
  AOI22_X1 U7614 ( .A1(n7156), .A2(n7122), .B1(n7120), .B2(n7155), .ZN(n7113)
         );
  AOI22_X1 U7615 ( .A1(n7157), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n7121), 
        .B2(n7154), .ZN(n7112) );
  OAI211_X1 U7616 ( .C1(n7160), .C2(n7125), .A(n7113), .B(n7112), .ZN(U3128)
         );
  AOI22_X1 U7617 ( .A1(n7168), .A2(n7122), .B1(n7120), .B2(n7161), .ZN(n7115)
         );
  AOI22_X1 U7618 ( .A1(n7163), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n7121), 
        .B2(n7162), .ZN(n7114) );
  OAI211_X1 U7619 ( .C1(n7166), .C2(n7125), .A(n7115), .B(n7114), .ZN(U3104)
         );
  AOI22_X1 U7620 ( .A1(n7169), .A2(n7122), .B1(n7120), .B2(n7167), .ZN(n7117)
         );
  AOI22_X1 U7621 ( .A1(n7170), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n7121), 
        .B2(n7168), .ZN(n7116) );
  OAI211_X1 U7622 ( .C1(n7173), .C2(n7125), .A(n7117), .B(n7116), .ZN(U3096)
         );
  AOI22_X1 U7623 ( .A1(n7176), .A2(n7122), .B1(n7120), .B2(n7174), .ZN(n7119)
         );
  AOI22_X1 U7624 ( .A1(n7177), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n7121), 
        .B2(n7175), .ZN(n7118) );
  OAI211_X1 U7625 ( .C1(n7180), .C2(n7125), .A(n7119), .B(n7118), .ZN(U3064)
         );
  AOI22_X1 U7626 ( .A1(n7185), .A2(n7121), .B1(n7120), .B2(n7181), .ZN(n7124)
         );
  AOI22_X1 U7627 ( .A1(n7187), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n7122), 
        .B2(n7184), .ZN(n7123) );
  OAI211_X1 U7628 ( .C1(n7191), .C2(n7125), .A(n7124), .B(n7123), .ZN(U3048)
         );
  AOI22_X1 U7629 ( .A1(n7156), .A2(n7136), .B1(n7134), .B2(n7155), .ZN(n7127)
         );
  AOI22_X1 U7630 ( .A1(n7157), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n7135), 
        .B2(n7154), .ZN(n7126) );
  OAI211_X1 U7631 ( .C1(n7160), .C2(n7139), .A(n7127), .B(n7126), .ZN(U3129)
         );
  AOI22_X1 U7632 ( .A1(n7168), .A2(n7136), .B1(n7134), .B2(n7161), .ZN(n7129)
         );
  AOI22_X1 U7633 ( .A1(n7163), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n7135), 
        .B2(n7162), .ZN(n7128) );
  OAI211_X1 U7634 ( .C1(n7166), .C2(n7139), .A(n7129), .B(n7128), .ZN(U3105)
         );
  AOI22_X1 U7635 ( .A1(n7168), .A2(n7135), .B1(n7134), .B2(n7167), .ZN(n7131)
         );
  AOI22_X1 U7636 ( .A1(n7170), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n7136), 
        .B2(n7169), .ZN(n7130) );
  OAI211_X1 U7637 ( .C1(n7173), .C2(n7139), .A(n7131), .B(n7130), .ZN(U3097)
         );
  AOI22_X1 U7638 ( .A1(n7176), .A2(n7136), .B1(n7134), .B2(n7174), .ZN(n7133)
         );
  AOI22_X1 U7639 ( .A1(n7177), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n7135), 
        .B2(n7175), .ZN(n7132) );
  OAI211_X1 U7640 ( .C1(n7180), .C2(n7139), .A(n7133), .B(n7132), .ZN(U3065)
         );
  AOI22_X1 U7641 ( .A1(n7185), .A2(n7135), .B1(n7134), .B2(n7181), .ZN(n7138)
         );
  AOI22_X1 U7642 ( .A1(n7187), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n7136), 
        .B2(n7184), .ZN(n7137) );
  OAI211_X1 U7643 ( .C1(n7191), .C2(n7139), .A(n7138), .B(n7137), .ZN(U3049)
         );
  AOI22_X1 U7644 ( .A1(n7156), .A2(n7150), .B1(n7148), .B2(n7155), .ZN(n7141)
         );
  AOI22_X1 U7645 ( .A1(n7157), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n7149), 
        .B2(n7154), .ZN(n7140) );
  OAI211_X1 U7646 ( .C1(n7160), .C2(n7153), .A(n7141), .B(n7140), .ZN(U3130)
         );
  AOI22_X1 U7647 ( .A1(n7168), .A2(n7150), .B1(n7148), .B2(n7161), .ZN(n7143)
         );
  AOI22_X1 U7648 ( .A1(n7163), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n7149), 
        .B2(n7162), .ZN(n7142) );
  OAI211_X1 U7649 ( .C1(n7166), .C2(n7153), .A(n7143), .B(n7142), .ZN(U3106)
         );
  AOI22_X1 U7650 ( .A1(n7169), .A2(n7150), .B1(n7148), .B2(n7167), .ZN(n7145)
         );
  AOI22_X1 U7651 ( .A1(n7170), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n7149), 
        .B2(n7168), .ZN(n7144) );
  OAI211_X1 U7652 ( .C1(n7173), .C2(n7153), .A(n7145), .B(n7144), .ZN(U3098)
         );
  AOI22_X1 U7653 ( .A1(n7175), .A2(n7149), .B1(n7148), .B2(n7174), .ZN(n7147)
         );
  AOI22_X1 U7654 ( .A1(n7177), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n7150), 
        .B2(n7176), .ZN(n7146) );
  OAI211_X1 U7655 ( .C1(n7180), .C2(n7153), .A(n7147), .B(n7146), .ZN(U3066)
         );
  AOI22_X1 U7656 ( .A1(n7185), .A2(n7149), .B1(n7148), .B2(n7181), .ZN(n7152)
         );
  AOI22_X1 U7657 ( .A1(n7187), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n7150), 
        .B2(n7184), .ZN(n7151) );
  OAI211_X1 U7658 ( .C1(n7191), .C2(n7153), .A(n7152), .B(n7151), .ZN(U3050)
         );
  AOI22_X1 U7659 ( .A1(n7182), .A2(n7155), .B1(n7154), .B2(n7186), .ZN(n7159)
         );
  AOI22_X1 U7660 ( .A1(n7157), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n7183), 
        .B2(n7156), .ZN(n7158) );
  OAI211_X1 U7661 ( .C1(n7160), .C2(n7190), .A(n7159), .B(n7158), .ZN(U3131)
         );
  AOI22_X1 U7662 ( .A1(n7168), .A2(n7183), .B1(n7182), .B2(n7161), .ZN(n7165)
         );
  AOI22_X1 U7663 ( .A1(n7163), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n7186), 
        .B2(n7162), .ZN(n7164) );
  OAI211_X1 U7664 ( .C1(n7166), .C2(n7190), .A(n7165), .B(n7164), .ZN(U3107)
         );
  AOI22_X1 U7665 ( .A1(n7168), .A2(n7186), .B1(n7182), .B2(n7167), .ZN(n7172)
         );
  AOI22_X1 U7666 ( .A1(n7170), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n7183), 
        .B2(n7169), .ZN(n7171) );
  OAI211_X1 U7667 ( .C1(n7173), .C2(n7190), .A(n7172), .B(n7171), .ZN(U3099)
         );
  AOI22_X1 U7668 ( .A1(n7175), .A2(n7186), .B1(n7182), .B2(n7174), .ZN(n7179)
         );
  AOI22_X1 U7669 ( .A1(n7177), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n7183), 
        .B2(n7176), .ZN(n7178) );
  OAI211_X1 U7670 ( .C1(n7180), .C2(n7190), .A(n7179), .B(n7178), .ZN(U3067)
         );
  AOI22_X1 U7671 ( .A1(n7184), .A2(n7183), .B1(n7182), .B2(n7181), .ZN(n7189)
         );
  AOI22_X1 U7672 ( .A1(n7187), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n7186), 
        .B2(n7185), .ZN(n7188) );
  OAI211_X1 U7673 ( .C1(n7191), .C2(n7190), .A(n7189), .B(n7188), .ZN(U3051)
         );
  CLKBUF_X1 U3477 ( .A(n3603), .Z(n4668) );
  CLKBUF_X1 U3513 ( .A(n3441), .Z(n4268) );
  NOR2_X2 U4196 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4968) );
  CLKBUF_X1 U5436 ( .A(n6014), .Z(n6015) );
  INV_X2 U5437 ( .A(n6902), .ZN(n6585) );
endmodule

