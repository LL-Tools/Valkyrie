

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, 
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, 
        keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, 
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, 
        keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, 
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, 
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994;

  AOI21_X1 U2372 ( .B1(n2833), .B2(n4906), .A(n2832), .ZN(n4431) );
  OR2_X1 U2373 ( .A1(n3109), .A2(n3091), .ZN(n3110) );
  AND4_X1 U2374 ( .A1(n2583), .A2(n2582), .A3(n2581), .A4(n2580), .ZN(n3294)
         );
  NAND2_X1 U2375 ( .A1(n2879), .A2(n3078), .ZN(n2986) );
  INV_X1 U2376 ( .A(n3055), .ZN(n3059) );
  AND2_X1 U2377 ( .A1(n2350), .A2(n2137), .ZN(n4438) );
  NAND2_X1 U2378 ( .A1(n2855), .A2(n4327), .ZN(n3300) );
  NOR2_X1 U2379 ( .A1(n3139), .A2(n3135), .ZN(n2852) );
  AOI21_X1 U2380 ( .B1(n3107), .B2(n4906), .A(n3106), .ZN(n3738) );
  AOI21_X1 U2381 ( .B1(n4638), .B2(n2711), .A(n2710), .ZN(n4613) );
  INV_X1 U2382 ( .A(n3336), .ZN(n4136) );
  INV_X2 U2383 ( .A(n3150), .ZN(n4177) );
  AND4_X1 U2384 ( .A1(n2598), .A2(n2597), .A3(n2596), .A4(n2595), .ZN(n3420)
         );
  XNOR2_X1 U2385 ( .A(n3241), .B(n3243), .ZN(n3244) );
  AND2_X1 U2386 ( .A1(n4901), .A2(n2855), .ZN(n4972) );
  XNOR2_X1 U2387 ( .A(n2456), .B(IR_REG_2__SCAN_IN), .ZN(n3164) );
  INV_X1 U2388 ( .A(n3294), .ZN(n4347) );
  XNOR2_X1 U2389 ( .A(n3102), .B(n4248), .ZN(n3743) );
  INV_X1 U2390 ( .A(n4896), .ZN(n4600) );
  INV_X2 U2391 ( .A(n4643), .ZN(n4668) );
  OR2_X2 U2392 ( .A1(n2837), .A2(IR_REG_22__SCAN_IN), .ZN(n2141) );
  OAI21_X2 U2393 ( .B1(n2140), .B2(n4842), .A(n2374), .ZN(n4858) );
  XNOR2_X2 U2394 ( .A(n4398), .B(n4397), .ZN(n4842) );
  NAND2_X2 U2395 ( .A1(n3194), .A2(n3193), .ZN(n3196) );
  XNOR2_X2 U2396 ( .A(n2545), .B(n3961), .ZN(n2551) );
  XNOR2_X2 U2397 ( .A(n4378), .B(n4794), .ZN(n4376) );
  INV_X4 U2398 ( .A(n2285), .ZN(n2585) );
  XNOR2_X2 U2399 ( .A(n3374), .B(n3383), .ZN(n3376) );
  OR2_X1 U2400 ( .A1(n2812), .A2(n2354), .ZN(n2350) );
  OR2_X1 U2401 ( .A1(n4378), .A2(n4377), .ZN(n4379) );
  NAND2_X1 U2402 ( .A1(n2793), .A2(n4191), .ZN(n3418) );
  AND2_X1 U2403 ( .A1(n4191), .A2(n4189), .ZN(n4272) );
  INV_X1 U2404 ( .A(n2578), .ZN(n2885) );
  INV_X1 U2405 ( .A(n2881), .ZN(n2880) );
  AND4_X1 U2406 ( .A1(n2664), .A2(n2663), .A3(n2662), .A4(n2661), .ZN(n3727)
         );
  AND2_X2 U2407 ( .A1(n3136), .A2(n4789), .ZN(n2781) );
  AOI211_X1 U2409 ( .C1(n4896), .C2(n3741), .A(n3740), .B(n3739), .ZN(n3742)
         );
  NAND2_X1 U2410 ( .A1(n4387), .A2(n4388), .ZN(n4801) );
  NAND2_X1 U2411 ( .A1(n4531), .A2(n4532), .ZN(n4530) );
  OAI21_X1 U2412 ( .B1(n4147), .B2(n2226), .A(n2223), .ZN(n3706) );
  NAND2_X1 U2413 ( .A1(n4613), .A2(n4612), .ZN(n4611) );
  NAND2_X1 U2414 ( .A1(n2305), .A2(n2304), .ZN(n4381) );
  NAND2_X1 U2415 ( .A1(n4380), .A2(n2144), .ZN(n2305) );
  NAND2_X1 U2416 ( .A1(n3690), .A2(n2701), .ZN(n4638) );
  NAND2_X1 U2417 ( .A1(n2194), .A2(n2193), .ZN(n3690) );
  AND2_X1 U2418 ( .A1(n2221), .A2(n2220), .ZN(n3446) );
  NAND2_X1 U2419 ( .A1(n2301), .A2(n2300), .ZN(n2303) );
  NAND2_X1 U2420 ( .A1(n3524), .A2(n2279), .ZN(n2276) );
  NAND2_X1 U2421 ( .A1(n2339), .A2(n2347), .ZN(n2344) );
  OAI21_X1 U2422 ( .B1(n3385), .B2(n2376), .A(n2378), .ZN(n3556) );
  NAND2_X1 U2423 ( .A1(n3434), .A2(n3433), .ZN(n3547) );
  NOR2_X1 U2424 ( .A1(n3323), .A2(n4054), .ZN(n3385) );
  NAND2_X1 U2425 ( .A1(n2212), .A2(n3383), .ZN(n2377) );
  OR2_X1 U2426 ( .A1(n3402), .A2(n3470), .ZN(n3526) );
  AOI21_X1 U2427 ( .B1(n2329), .B2(n2332), .A(n2169), .ZN(n2327) );
  NAND2_X1 U2428 ( .A1(n3321), .A2(n2154), .ZN(n3382) );
  NOR2_X2 U2429 ( .A1(n3089), .A2(n4912), .ZN(n3090) );
  AND2_X1 U2430 ( .A1(n2373), .A2(n2372), .ZN(n2370) );
  NOR2_X1 U2431 ( .A1(n2792), .A2(n2319), .ZN(n2318) );
  AND2_X1 U2432 ( .A1(n4188), .A2(n4185), .ZN(n4271) );
  XNOR2_X1 U2433 ( .A(n3235), .B(n3243), .ZN(n3237) );
  AND2_X2 U2434 ( .A1(n3119), .A2(n4931), .ZN(U4043) );
  NOR2_X1 U2435 ( .A1(n3207), .A2(n3206), .ZN(n3235) );
  NAND2_X2 U2436 ( .A1(n3300), .A2(n3077), .ZN(n3055) );
  AND4_X1 U2437 ( .A1(n2616), .A2(n2615), .A3(n2614), .A4(n2613), .ZN(n3353)
         );
  INV_X1 U2438 ( .A(n2606), .ZN(n3717) );
  INV_X1 U2439 ( .A(n2869), .ZN(n4327) );
  XNOR2_X1 U2440 ( .A(n3187), .B(n3195), .ZN(n2206) );
  NAND2_X1 U2442 ( .A1(n4840), .A2(n4667), .ZN(n2304) );
  BUF_X2 U2443 ( .A(n2142), .Z(n3215) );
  NAND2_X1 U2444 ( .A1(n2532), .A2(n2837), .ZN(n2869) );
  NAND2_X1 U2445 ( .A1(n3186), .A2(n3185), .ZN(n3187) );
  NAND3_X1 U2446 ( .A1(n2141), .A2(IR_REG_31__SCAN_IN), .A3(IR_REG_24__SCAN_IN), .ZN(n2842) );
  NAND2_X1 U2447 ( .A1(n2443), .A2(n2444), .ZN(n2844) );
  AND3_X1 U2448 ( .A1(n2150), .A2(n2337), .A3(n2336), .ZN(n2338) );
  NOR2_X1 U2449 ( .A1(n2525), .A2(n2442), .ZN(n2443) );
  NAND2_X1 U2450 ( .A1(n2441), .A2(n2262), .ZN(n2442) );
  NAND2_X1 U2451 ( .A1(n2460), .A2(n2261), .ZN(n2472) );
  NAND2_X1 U2452 ( .A1(n2147), .A2(n2519), .ZN(n2525) );
  NAND2_X1 U2453 ( .A1(n2454), .A2(n2379), .ZN(n3169) );
  AND2_X1 U2454 ( .A1(n2440), .A2(n2439), .ZN(n2519) );
  AND2_X1 U2455 ( .A1(n2433), .A2(n2434), .ZN(n2261) );
  AND4_X1 U2456 ( .A1(n2437), .A2(n2436), .A3(n2435), .A4(n2478), .ZN(n2438)
         );
  NAND2_X1 U2457 ( .A1(n2853), .A2(n2840), .ZN(n2843) );
  INV_X1 U2458 ( .A(IR_REG_19__SCAN_IN), .ZN(n2522) );
  NOR2_X1 U2459 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2434)
         );
  NOR2_X1 U2460 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2433)
         );
  INV_X1 U2461 ( .A(IR_REG_24__SCAN_IN), .ZN(n2840) );
  INV_X1 U2462 ( .A(IR_REG_23__SCAN_IN), .ZN(n2853) );
  NOR2_X1 U2463 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2435)
         );
  NOR2_X1 U2464 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2437)
         );
  INV_X1 U2465 ( .A(IR_REG_8__SCAN_IN), .ZN(n2478) );
  NOR2_X1 U2466 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2436)
         );
  XNOR2_X1 U2467 ( .A(n3556), .B(n3438), .ZN(n3439) );
  BUF_X8 U2468 ( .A(n2986), .Z(n2131) );
  NOR2_X2 U2469 ( .A1(n4521), .A2(n2752), .ZN(n4501) );
  NOR2_X1 U2470 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2544)
         );
  INV_X1 U2471 ( .A(IR_REG_28__SCAN_IN), .ZN(n3850) );
  INV_X1 U2472 ( .A(n2472), .ZN(n2205) );
  NAND2_X1 U2473 ( .A1(n2201), .A2(n2788), .ZN(n3102) );
  OR2_X1 U2474 ( .A1(n3057), .A2(n4447), .ZN(n2788) );
  NAND2_X1 U2475 ( .A1(n2200), .A2(n2175), .ZN(n2201) );
  NAND2_X1 U2476 ( .A1(n3648), .A2(n2694), .ZN(n2194) );
  NOR2_X1 U2477 ( .A1(n4840), .A2(n4736), .ZN(n4396) );
  INV_X1 U2478 ( .A(n3524), .ZN(n2283) );
  INV_X1 U2479 ( .A(IR_REG_9__SCAN_IN), .ZN(n3918) );
  AND2_X1 U2480 ( .A1(n4286), .A2(n2624), .ZN(n2625) );
  NAND2_X1 U2481 ( .A1(n4346), .A2(n3717), .ZN(n4191) );
  AND2_X1 U2482 ( .A1(n2192), .A2(n2191), .ZN(n2665) );
  NAND2_X1 U2483 ( .A1(n4178), .A2(n3959), .ZN(n2191) );
  NAND2_X1 U2484 ( .A1(n3502), .A2(n3255), .ZN(n2392) );
  INV_X1 U2485 ( .A(IR_REG_27__SCAN_IN), .ZN(n2543) );
  NAND2_X1 U2486 ( .A1(n2135), .A2(n3254), .ZN(n2216) );
  AND2_X1 U2487 ( .A1(n4177), .A2(DATAI_21_), .ZN(n2810) );
  INV_X1 U2488 ( .A(n3694), .ZN(n3805) );
  INV_X1 U2489 ( .A(n3707), .ZN(n3031) );
  INV_X1 U2490 ( .A(n3215), .ZN(n2784) );
  INV_X1 U2491 ( .A(n2586), .ZN(n2748) );
  INV_X1 U2492 ( .A(n2781), .ZN(n2771) );
  AND4_X1 U2493 ( .A1(n2605), .A2(n2604), .A3(n2603), .A4(n2602), .ZN(n3716)
         );
  INV_X1 U2494 ( .A(n3136), .ZN(n2552) );
  NAND2_X1 U2495 ( .A1(n3171), .A2(n3170), .ZN(n4350) );
  OR2_X1 U2496 ( .A1(n3169), .A2(REG1_REG_1__SCAN_IN), .ZN(n3171) );
  NAND2_X1 U2497 ( .A1(n2363), .A2(n2362), .ZN(n3207) );
  NAND2_X1 U2498 ( .A1(n3188), .A2(n2367), .ZN(n2362) );
  NAND2_X1 U2499 ( .A1(n2206), .A2(n2157), .ZN(n2363) );
  AND2_X1 U2500 ( .A1(n3187), .A2(n4820), .ZN(n3188) );
  AOI21_X1 U2501 ( .B1(n3195), .B2(REG2_REG_4__SCAN_IN), .A(n4820), .ZN(n2293)
         );
  NAND2_X1 U2502 ( .A1(n2298), .A2(n2187), .ZN(n2301) );
  NAND2_X1 U2503 ( .A1(n3547), .A2(n2299), .ZN(n2298) );
  NAND2_X1 U2504 ( .A1(n2188), .A2(n2176), .ZN(n2187) );
  OR2_X1 U2505 ( .A1(n3438), .A2(n2302), .ZN(n2299) );
  NAND2_X1 U2506 ( .A1(n4795), .A2(REG1_REG_11__SCAN_IN), .ZN(n3642) );
  NAND2_X1 U2507 ( .A1(n4866), .A2(n4386), .ZN(n4387) );
  NAND2_X1 U2508 ( .A1(n4437), .A2(n4467), .ZN(n2777) );
  NAND2_X1 U2509 ( .A1(n4455), .A2(n2431), .ZN(n2200) );
  NOR2_X1 U2510 ( .A1(n4090), .A2(n2241), .ZN(n2238) );
  OR2_X1 U2511 ( .A1(n2737), .A2(n2566), .ZN(n2744) );
  OAI21_X1 U2512 ( .B1(n2804), .B2(n2324), .A(n2322), .ZN(n3692) );
  INV_X1 U2513 ( .A(n2323), .ZN(n2322) );
  OAI21_X1 U2514 ( .B1(n2145), .B2(n2324), .A(n4288), .ZN(n2323) );
  INV_X1 U2515 ( .A(n4209), .ZN(n2324) );
  AND2_X1 U2516 ( .A1(n4302), .A2(n4298), .ZN(n4288) );
  NAND2_X1 U2517 ( .A1(n2535), .A2(n2245), .ZN(n2703) );
  NOR2_X1 U2518 ( .A1(n2246), .A2(n2679), .ZN(n2245) );
  NAND2_X1 U2519 ( .A1(n2276), .A2(n2274), .ZN(n3648) );
  NOR2_X1 U2520 ( .A1(n2275), .A2(n2156), .ZN(n2274) );
  NAND2_X1 U2521 ( .A1(n2549), .A2(IR_REG_31__SCAN_IN), .ZN(n2545) );
  INV_X1 U2522 ( .A(IR_REG_3__SCAN_IN), .ZN(n2464) );
  INV_X1 U2523 ( .A(IR_REG_1__SCAN_IN), .ZN(n2316) );
  INV_X1 U2524 ( .A(IR_REG_0__SCAN_IN), .ZN(n2317) );
  NOR2_X1 U2525 ( .A1(n4313), .A2(n2357), .ZN(n2355) );
  NOR2_X1 U2526 ( .A1(n2672), .A2(n2280), .ZN(n2203) );
  INV_X1 U2527 ( .A(n4273), .ZN(n2204) );
  NOR2_X1 U2528 ( .A1(n3569), .A2(n3449), .ZN(n2280) );
  NOR2_X1 U2529 ( .A1(n3724), .A2(n2409), .ZN(n2408) );
  INV_X1 U2530 ( .A(n2411), .ZN(n2409) );
  INV_X1 U2531 ( .A(n2814), .ZN(n4313) );
  AND2_X1 U2532 ( .A1(n4429), .A2(n2427), .ZN(n4262) );
  AND2_X1 U2533 ( .A1(n2252), .A2(n2248), .ZN(n2247) );
  INV_X1 U2534 ( .A(n4496), .ZN(n2252) );
  NOR2_X1 U2535 ( .A1(n4514), .A2(n2249), .ZN(n2248) );
  NAND2_X1 U2536 ( .A1(n2160), .A2(n4394), .ZN(n2208) );
  INV_X1 U2537 ( .A(n4396), .ZN(n2211) );
  NAND2_X1 U2538 ( .A1(n4401), .A2(n2422), .ZN(n4403) );
  AND2_X1 U2539 ( .A1(n4937), .A2(REG2_REG_15__SCAN_IN), .ZN(n4383) );
  OAI21_X1 U2540 ( .B1(n2270), .B2(n2268), .A(n2760), .ZN(n2267) );
  NAND2_X1 U2541 ( .A1(n4480), .A2(n4502), .ZN(n2271) );
  INV_X1 U2542 ( .A(n2753), .ZN(n2539) );
  NAND2_X1 U2543 ( .A1(n4340), .A2(n2752), .ZN(n2272) );
  OR2_X1 U2544 ( .A1(n2675), .A2(n3853), .ZN(n2680) );
  NAND2_X1 U2545 ( .A1(n4342), .A2(n2190), .ZN(n3587) );
  AOI21_X1 U2546 ( .B1(n2333), .B2(n2331), .A(n2330), .ZN(n2329) );
  INV_X1 U2547 ( .A(n4199), .ZN(n2331) );
  INV_X1 U2548 ( .A(n2333), .ZN(n2332) );
  NAND2_X1 U2549 ( .A1(n2347), .A2(n2346), .ZN(n2343) );
  INV_X1 U2550 ( .A(n4204), .ZN(n2346) );
  INV_X1 U2551 ( .A(n3418), .ZN(n2339) );
  INV_X1 U2552 ( .A(n2592), .ZN(n2255) );
  INV_X1 U2553 ( .A(n2607), .ZN(n2256) );
  NAND2_X1 U2554 ( .A1(n3360), .A2(n2591), .ZN(n2257) );
  INV_X1 U2555 ( .A(n4188), .ZN(n2319) );
  NAND2_X1 U2556 ( .A1(n4186), .A2(n4183), .ZN(n2258) );
  NOR2_X1 U2557 ( .A1(n2415), .A2(n4155), .ZN(n2414) );
  INV_X1 U2558 ( .A(n2416), .ZN(n2415) );
  NOR2_X1 U2559 ( .A1(n2810), .A2(n4577), .ZN(n2420) );
  AND2_X1 U2560 ( .A1(n4268), .A2(n4267), .ZN(n4571) );
  NOR2_X1 U2561 ( .A1(n2521), .A2(n2525), .ZN(n2529) );
  NAND2_X1 U2562 ( .A1(n3486), .A2(n2948), .ZN(n2411) );
  OR2_X1 U2563 ( .A1(n3486), .A2(n2948), .ZN(n2412) );
  XNOR2_X1 U2564 ( .A(n2900), .B(n3059), .ZN(n2906) );
  OAI22_X1 U2565 ( .A1(n3420), .A2(n2131), .B1(n3717), .B2(n3058), .ZN(n2900)
         );
  NAND2_X1 U2566 ( .A1(n2229), .A2(n2227), .ZN(n3838) );
  INV_X1 U2567 ( .A(n2230), .ZN(n2227) );
  NAND2_X1 U2568 ( .A1(n4147), .A2(n2232), .ZN(n2229) );
  OAI21_X1 U2569 ( .B1(n2975), .B2(n2974), .A(n3680), .ZN(n2976) );
  NAND2_X1 U2570 ( .A1(n3792), .A2(n3793), .ZN(n2397) );
  OR2_X1 U2571 ( .A1(n4802), .A2(n2883), .ZN(n3077) );
  NAND2_X1 U2572 ( .A1(n4350), .A2(n4351), .ZN(n4364) );
  OAI211_X1 U2573 ( .C1(n2146), .C2(n3196), .A(n2295), .B(n2290), .ZN(n2297)
         );
  INV_X1 U2574 ( .A(n3198), .ZN(n2295) );
  NAND2_X1 U2575 ( .A1(n2485), .A2(n3918), .ZN(n2489) );
  NAND2_X1 U2576 ( .A1(n3432), .A2(REG2_REG_9__SCAN_IN), .ZN(n3433) );
  NAND2_X1 U2577 ( .A1(n3386), .A2(n2166), .ZN(n2378) );
  NAND2_X1 U2578 ( .A1(n2377), .A2(n2166), .ZN(n2376) );
  INV_X1 U2579 ( .A(n3550), .ZN(n2300) );
  NAND2_X1 U2580 ( .A1(n4376), .A2(REG2_REG_12__SCAN_IN), .ZN(n4380) );
  NAND2_X1 U2581 ( .A1(n4392), .A2(n4794), .ZN(n4393) );
  INV_X1 U2582 ( .A(n4939), .ZN(n4397) );
  XNOR2_X1 U2583 ( .A(n4403), .B(n4936), .ZN(n4871) );
  NAND2_X1 U2584 ( .A1(n4805), .A2(n2182), .ZN(n2380) );
  AND2_X1 U2585 ( .A1(n2767), .A2(n2766), .ZN(n4461) );
  OR2_X1 U2586 ( .A1(n2744), .A2(n3773), .ZN(n2753) );
  AND2_X1 U2587 ( .A1(n2272), .A2(n2273), .ZN(n2270) );
  AND2_X1 U2588 ( .A1(n4512), .A2(n4511), .ZN(n4533) );
  AND2_X1 U2589 ( .A1(n2198), .A2(n2197), .ZN(n4531) );
  NAND2_X1 U2590 ( .A1(n4570), .A2(n4557), .ZN(n2197) );
  AND2_X1 U2591 ( .A1(n2138), .A2(REG3_REG_21__SCAN_IN), .ZN(n2234) );
  NAND2_X1 U2592 ( .A1(n2199), .A2(n4267), .ZN(n4547) );
  NAND2_X1 U2593 ( .A1(n2728), .A2(n2195), .ZN(n2199) );
  NOR2_X1 U2594 ( .A1(n4266), .A2(n2196), .ZN(n2195) );
  AND2_X1 U2595 ( .A1(n2718), .A2(n2717), .ZN(n4624) );
  AND2_X1 U2596 ( .A1(n2709), .A2(n2708), .ZN(n4605) );
  AND2_X1 U2597 ( .A1(n2700), .A2(n2149), .ZN(n2193) );
  NAND2_X1 U2598 ( .A1(n2535), .A2(REG3_REG_14__SCAN_IN), .ZN(n2685) );
  NAND2_X1 U2599 ( .A1(n2804), .A2(n2145), .ZN(n3654) );
  AND2_X1 U2600 ( .A1(n3584), .A2(n3587), .ZN(n4273) );
  OR2_X1 U2601 ( .A1(n2647), .A2(n2646), .ZN(n2648) );
  NAND2_X1 U2602 ( .A1(n2244), .A2(REG3_REG_8__SCAN_IN), .ZN(n2636) );
  NAND2_X1 U2603 ( .A1(n3418), .A2(n4204), .ZN(n2348) );
  INV_X1 U2604 ( .A(n4647), .ZN(n4630) );
  AND2_X1 U2605 ( .A1(n3175), .A2(n3152), .ZN(n4660) );
  INV_X1 U2606 ( .A(n4906), .ZN(n4655) );
  INV_X1 U2607 ( .A(n2258), .ZN(n4276) );
  AND2_X1 U2608 ( .A1(n2883), .A2(n2869), .ZN(n4901) );
  NOR2_X2 U2609 ( .A1(n3110), .A2(n4237), .ZN(n4418) );
  AND2_X1 U2610 ( .A1(n2564), .A2(n4429), .ZN(n2565) );
  INV_X1 U2611 ( .A(n2665), .ZN(n2190) );
  AND2_X1 U2612 ( .A1(n3577), .A2(n2190), .ZN(n3599) );
  INV_X1 U2613 ( .A(n3449), .ZN(n3525) );
  INV_X1 U2614 ( .A(n4967), .ZN(n4975) );
  INV_X1 U2615 ( .A(n3281), .ZN(n3067) );
  NAND2_X1 U2616 ( .A1(n2879), .A2(n4931), .ZN(n3149) );
  NAND2_X1 U2617 ( .A1(n2338), .A2(n2444), .ZN(n2549) );
  NOR2_X1 U2618 ( .A1(n2442), .A2(IR_REG_29__SCAN_IN), .ZN(n2336) );
  INV_X1 U2619 ( .A(n2525), .ZN(n2337) );
  AND4_X1 U2620 ( .A1(n2260), .A2(n2150), .A3(n2438), .A4(n2259), .ZN(n2824)
         );
  INV_X1 U2621 ( .A(n2442), .ZN(n2259) );
  NOR2_X1 U2622 ( .A1(n2525), .A2(n2472), .ZN(n2260) );
  XNOR2_X1 U2623 ( .A(n2215), .B(n2253), .ZN(n2855) );
  NAND2_X1 U2624 ( .A1(n2533), .A2(IR_REG_31__SCAN_IN), .ZN(n2215) );
  OAI21_X1 U2625 ( .B1(n2521), .B2(n2520), .A(IR_REG_31__SCAN_IN), .ZN(n2523)
         );
  NAND2_X1 U2626 ( .A1(n2523), .A2(n2522), .ZN(n2533) );
  INV_X1 U2627 ( .A(IR_REG_15__SCAN_IN), .ZN(n4022) );
  INV_X1 U2628 ( .A(n2444), .ZN(n2521) );
  MUX2_X1 U2629 ( .A(IR_REG_31__SCAN_IN), .B(n2453), .S(IR_REG_1__SCAN_IN), 
        .Z(n2454) );
  OR2_X1 U2630 ( .A1(n4470), .A2(n2771), .ZN(n2776) );
  INV_X1 U2631 ( .A(n4552), .ZN(n4516) );
  OAI21_X1 U2632 ( .B1(n2385), .B2(n2384), .A(n2159), .ZN(n2382) );
  NAND2_X1 U2633 ( .A1(n2410), .A2(n2411), .ZN(n3726) );
  NAND2_X1 U2634 ( .A1(n3484), .A2(n2412), .ZN(n2410) );
  XNOR2_X1 U2635 ( .A(n2906), .B(n2907), .ZN(n3714) );
  AOI21_X1 U2636 ( .B1(n2228), .B2(n2225), .A(n2224), .ZN(n2223) );
  INV_X1 U2637 ( .A(n2228), .ZN(n2226) );
  INV_X1 U2638 ( .A(n2398), .ZN(n2224) );
  INV_X1 U2639 ( .A(n3222), .ZN(n3569) );
  NAND2_X1 U2640 ( .A1(n2189), .A2(n3552), .ZN(n3488) );
  OR2_X1 U2641 ( .A1(n3090), .A2(n2190), .ZN(n2189) );
  AND2_X1 U2642 ( .A1(n3084), .A2(STATE_REG_SCAN_IN), .ZN(n3845) );
  NAND2_X1 U2643 ( .A1(n2397), .A2(n2396), .ZN(n2222) );
  INV_X1 U2644 ( .A(n3090), .ZN(n4171) );
  INV_X1 U2645 ( .A(n4135), .ZN(n4167) );
  NAND2_X1 U2646 ( .A1(n2563), .A2(n2562), .ZN(n4240) );
  INV_X1 U2647 ( .A(n3062), .ZN(n4444) );
  NAND2_X1 U2648 ( .A1(n2787), .A2(n2786), .ZN(n4463) );
  INV_X1 U2649 ( .A(n4461), .ZN(n4498) );
  NAND2_X1 U2650 ( .A1(n2691), .A2(n2690), .ZN(n3694) );
  NAND2_X1 U2651 ( .A1(n2286), .A2(n2552), .ZN(n2284) );
  NAND2_X1 U2652 ( .A1(n2142), .A2(REG2_REG_0__SCAN_IN), .ZN(n2574) );
  NAND2_X1 U2653 ( .A1(n2364), .A2(n2369), .ZN(n2368) );
  INV_X1 U2654 ( .A(n3188), .ZN(n2369) );
  OAI21_X1 U2655 ( .B1(n2292), .B2(n2293), .A(n2291), .ZN(n2296) );
  NAND2_X1 U2656 ( .A1(n2292), .A2(n2146), .ZN(n2291) );
  INV_X1 U2657 ( .A(n3196), .ZN(n2292) );
  INV_X1 U2658 ( .A(n2297), .ZN(n3205) );
  NAND2_X1 U2659 ( .A1(n2495), .A2(n2496), .ZN(n3640) );
  AND2_X1 U2660 ( .A1(n2380), .A2(n4873), .ZN(n2213) );
  NAND2_X1 U2661 ( .A1(n2180), .A2(n2312), .ZN(n2311) );
  OAI22_X1 U2662 ( .A1(n2139), .A2(n2311), .B1(n2180), .B2(n2312), .ZN(n2309)
         );
  INV_X1 U2663 ( .A(n4875), .ZN(n4878) );
  AND2_X1 U2664 ( .A1(n2139), .A2(n2186), .ZN(n2310) );
  XNOR2_X1 U2665 ( .A(n4240), .B(n4237), .ZN(n4429) );
  INV_X1 U2666 ( .A(n3175), .ZN(n4790) );
  NAND2_X1 U2667 ( .A1(n2469), .A2(n2472), .ZN(n3204) );
  AND2_X1 U2668 ( .A1(n2813), .A2(n4456), .ZN(n2814) );
  NOR2_X1 U2669 ( .A1(n4612), .A2(n2251), .ZN(n2250) );
  NAND2_X1 U2670 ( .A1(n3322), .A2(REG1_REG_7__SCAN_IN), .ZN(n2372) );
  OR2_X1 U2671 ( .A1(n2642), .A2(n2641), .ZN(n2644) );
  NAND2_X1 U2672 ( .A1(n4347), .A2(n2458), .ZN(n4186) );
  INV_X1 U2673 ( .A(IR_REG_17__SCAN_IN), .ZN(n3852) );
  INV_X1 U2674 ( .A(n3058), .ZN(n3010) );
  OAI22_X1 U2675 ( .A1(n3779), .A2(n2231), .B1(n3015), .B2(n3016), .ZN(n2230)
         );
  NOR2_X1 U2676 ( .A1(n3779), .A2(n2233), .ZN(n2232) );
  INV_X1 U2677 ( .A(n4145), .ZN(n2233) );
  AND2_X1 U2678 ( .A1(n2404), .A2(n2969), .ZN(n2403) );
  AND2_X1 U2679 ( .A1(n2968), .A2(n3681), .ZN(n2969) );
  NAND2_X1 U2680 ( .A1(n2405), .A2(n2407), .ZN(n2404) );
  NOR2_X1 U2681 ( .A1(n2617), .A2(n2534), .ZN(n2610) );
  INV_X1 U2682 ( .A(n3300), .ZN(n3078) );
  AND2_X1 U2683 ( .A1(n3555), .A2(REG2_REG_10__SCAN_IN), .ZN(n2302) );
  INV_X1 U2684 ( .A(n3547), .ZN(n2188) );
  INV_X1 U2685 ( .A(n4834), .ZN(n2306) );
  INV_X1 U2686 ( .A(n4463), .ZN(n3057) );
  AND2_X1 U2687 ( .A1(n4233), .A2(n2352), .ZN(n2351) );
  NAND2_X1 U2688 ( .A1(n2355), .A2(n2353), .ZN(n2352) );
  INV_X1 U2689 ( .A(n4307), .ZN(n2353) );
  INV_X1 U2690 ( .A(n2355), .ZN(n2354) );
  AND2_X1 U2691 ( .A1(REG3_REG_25__SCAN_IN), .A2(n2240), .ZN(n2239) );
  NOR2_X1 U2692 ( .A1(n2242), .A2(n2241), .ZN(n2240) );
  NAND2_X1 U2693 ( .A1(n2358), .A2(n2356), .ZN(n4477) );
  INV_X1 U2694 ( .A(n4252), .ZN(n2359) );
  AND2_X1 U2695 ( .A1(n4593), .A2(n4577), .ZN(n4266) );
  AND2_X1 U2696 ( .A1(n2809), .A2(n4299), .ZN(n4304) );
  NOR2_X1 U2697 ( .A1(n4046), .A2(n2236), .ZN(n2235) );
  INV_X1 U2698 ( .A(n2712), .ZN(n2538) );
  INV_X1 U2699 ( .A(n2680), .ZN(n2535) );
  NAND2_X1 U2700 ( .A1(n2161), .A2(n2202), .ZN(n2275) );
  NAND2_X1 U2701 ( .A1(n2279), .A2(n2657), .ZN(n2202) );
  INV_X1 U2702 ( .A(n2659), .ZN(n2243) );
  NAND2_X1 U2703 ( .A1(n2281), .A2(n2278), .ZN(n3571) );
  INV_X1 U2704 ( .A(n2280), .ZN(n2278) );
  NAND2_X1 U2705 ( .A1(n2283), .A2(n2282), .ZN(n2281) );
  INV_X1 U2706 ( .A(n2634), .ZN(n2244) );
  AND2_X1 U2707 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n3869) );
  NOR2_X1 U2708 ( .A1(n3047), .A2(n3831), .ZN(n2416) );
  NOR2_X1 U2709 ( .A1(n3651), .A2(n4172), .ZN(n3697) );
  NOR2_X1 U2710 ( .A1(n2392), .A2(n2389), .ZN(n3401) );
  INV_X1 U2711 ( .A(IR_REG_22__SCAN_IN), .ZN(n2527) );
  INV_X1 U2712 ( .A(IR_REG_20__SCAN_IN), .ZN(n2253) );
  NOR2_X1 U2713 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2440)
         );
  NOR2_X1 U2714 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2439)
         );
  OR2_X1 U2715 ( .A1(n2513), .A2(IR_REG_17__SCAN_IN), .ZN(n2516) );
  OR2_X1 U2716 ( .A1(n2489), .A2(IR_REG_10__SCAN_IN), .ZN(n2491) );
  AND2_X1 U2717 ( .A1(n2480), .A2(IR_REG_31__SCAN_IN), .ZN(n2473) );
  INV_X1 U2718 ( .A(IR_REG_2__SCAN_IN), .ZN(n3851) );
  INV_X1 U2719 ( .A(n3406), .ZN(n2384) );
  NAND2_X1 U2720 ( .A1(n2136), .A2(n2183), .ZN(n2217) );
  INV_X1 U2721 ( .A(n3272), .ZN(n2218) );
  INV_X1 U2722 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2650) );
  INV_X1 U2723 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4046) );
  NAND2_X1 U2724 ( .A1(n2397), .A2(n2174), .ZN(n2395) );
  AND2_X1 U2725 ( .A1(n2954), .A2(n2955), .ZN(n3724) );
  NAND2_X1 U2726 ( .A1(n2388), .A2(n2928), .ZN(n2387) );
  INV_X1 U2727 ( .A(n3349), .ZN(n2388) );
  INV_X1 U2728 ( .A(n2386), .ZN(n2385) );
  OAI21_X1 U2729 ( .B1(n3751), .B2(n2387), .A(n3348), .ZN(n2386) );
  NAND2_X1 U2730 ( .A1(n2452), .A2(n2451), .ZN(n2457) );
  NAND2_X1 U2731 ( .A1(n3838), .A2(n3839), .ZN(n3837) );
  INV_X1 U2732 ( .A(n2408), .ZN(n2407) );
  AOI21_X1 U2733 ( .B1(n2408), .B2(n2406), .A(n2181), .ZN(n2405) );
  INV_X1 U2734 ( .A(n2412), .ZN(n2406) );
  AOI21_X1 U2735 ( .B1(n2400), .B2(n2399), .A(n2158), .ZN(n2398) );
  INV_X1 U2736 ( .A(n3839), .ZN(n2399) );
  NOR2_X1 U2737 ( .A1(n2230), .A2(n2401), .ZN(n2228) );
  INV_X1 U2738 ( .A(n2232), .ZN(n2225) );
  OAI22_X1 U2739 ( .A1(n2131), .A2(n3727), .B1(n3058), .B2(n2190), .ZN(n2947)
         );
  OR2_X1 U2740 ( .A1(n2651), .A2(n2650), .ZN(n2659) );
  INV_X1 U2741 ( .A(n3314), .ZN(n2458) );
  AOI21_X1 U2742 ( .B1(n3229), .B2(n3228), .A(n2890), .ZN(n4131) );
  AND2_X1 U2743 ( .A1(n3152), .A2(n3068), .ZN(n3081) );
  INV_X1 U2744 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2534) );
  AND2_X1 U2745 ( .A1(n4262), .A2(n2247), .ZN(n4293) );
  AND2_X1 U2746 ( .A1(n2557), .A2(n2556), .ZN(n3062) );
  OR2_X1 U2747 ( .A1(n3737), .A2(n2771), .ZN(n2557) );
  NAND2_X1 U2748 ( .A1(n2288), .A2(n2287), .ZN(n2286) );
  NAND2_X1 U2749 ( .A1(n2361), .A2(n3174), .ZN(n3184) );
  NOR2_X1 U2750 ( .A1(n3204), .A2(n4989), .ZN(n3206) );
  AND2_X2 U2751 ( .A1(n2297), .A2(n2151), .ZN(n3241) );
  INV_X1 U2752 ( .A(n3382), .ZN(n2212) );
  NAND2_X1 U2753 ( .A1(n2315), .A2(n2314), .ZN(n3378) );
  NAND2_X1 U2754 ( .A1(n3375), .A2(n3383), .ZN(n2314) );
  AND2_X1 U2755 ( .A1(n2491), .A2(IR_REG_31__SCAN_IN), .ZN(n2492) );
  NAND2_X1 U2756 ( .A1(n2208), .A2(n2209), .ZN(n4398) );
  AND2_X1 U2757 ( .A1(n2208), .A2(n2207), .ZN(n4399) );
  NOR2_X1 U2758 ( .A1(n2210), .A2(n4397), .ZN(n2207) );
  NOR2_X1 U2759 ( .A1(n4842), .A2(n4843), .ZN(n4841) );
  INV_X1 U2760 ( .A(n4403), .ZN(n4402) );
  INV_X1 U2761 ( .A(n2186), .ZN(n2312) );
  AND2_X1 U2762 ( .A1(n2780), .A2(n2779), .ZN(n4448) );
  NAND2_X1 U2763 ( .A1(n2350), .A2(n2351), .ZN(n4439) );
  AND2_X1 U2764 ( .A1(n2143), .A2(n2762), .ZN(n4489) );
  NAND2_X1 U2765 ( .A1(n2269), .A2(n2271), .ZN(n2264) );
  INV_X1 U2766 ( .A(n2271), .ZN(n2263) );
  INV_X1 U2767 ( .A(n2267), .ZN(n2266) );
  AND2_X1 U2768 ( .A1(n4456), .A2(n4258), .ZN(n4478) );
  AND2_X1 U2769 ( .A1(n2358), .A2(n2359), .ZN(n4495) );
  AND2_X1 U2770 ( .A1(n2751), .A2(n2750), .ZN(n4536) );
  AND2_X1 U2771 ( .A1(n2734), .A2(n2733), .ZN(n4550) );
  NAND2_X1 U2772 ( .A1(n2538), .A2(n2138), .ZN(n2735) );
  NAND2_X1 U2773 ( .A1(n2538), .A2(REG3_REG_18__SCAN_IN), .ZN(n2720) );
  INV_X1 U2774 ( .A(REG3_REG_17__SCAN_IN), .ZN(n3821) );
  INV_X1 U2775 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2702) );
  NAND2_X1 U2776 ( .A1(n2537), .A2(n2536), .ZN(n2712) );
  NOR2_X1 U2777 ( .A1(n2702), .A2(n3821), .ZN(n2536) );
  INV_X1 U2778 ( .A(n2703), .ZN(n2537) );
  NOR2_X1 U2779 ( .A1(n2326), .A2(n2325), .ZN(n2429) );
  INV_X1 U2780 ( .A(n4215), .ZN(n2325) );
  INV_X1 U2781 ( .A(n2804), .ZN(n2326) );
  NAND2_X1 U2782 ( .A1(n2276), .A2(n2277), .ZN(n4644) );
  INV_X1 U2783 ( .A(n2275), .ZN(n2277) );
  NAND2_X1 U2784 ( .A1(n3727), .A2(n2190), .ZN(n3595) );
  NAND2_X1 U2785 ( .A1(n2243), .A2(REG3_REG_11__SCAN_IN), .ZN(n2666) );
  AND2_X1 U2786 ( .A1(n2343), .A2(n2342), .ZN(n2341) );
  NOR2_X1 U2787 ( .A1(n2345), .A2(n2795), .ZN(n2342) );
  NAND2_X1 U2788 ( .A1(n2344), .A2(n2340), .ZN(n3492) );
  AND2_X1 U2789 ( .A1(n2343), .A2(n4193), .ZN(n2340) );
  AND4_X1 U2790 ( .A1(n2640), .A2(n2639), .A3(n2638), .A4(n2637), .ZN(n3495)
         );
  NOR2_X1 U2791 ( .A1(n2432), .A2(n2424), .ZN(n2608) );
  NAND2_X1 U2792 ( .A1(n3869), .A2(REG3_REG_5__SCAN_IN), .ZN(n2617) );
  NAND2_X1 U2793 ( .A1(n2791), .A2(n2318), .ZN(n2793) );
  INV_X1 U2794 ( .A(n3869), .ZN(n2600) );
  NAND2_X1 U2795 ( .A1(n2791), .A2(n4188), .ZN(n2321) );
  NOR2_X1 U2796 ( .A1(n3367), .A2(n3368), .ZN(n3366) );
  INV_X1 U2797 ( .A(n3291), .ZN(n3286) );
  INV_X1 U2798 ( .A(n3747), .ZN(n4903) );
  AND2_X1 U2799 ( .A1(n2414), .A2(n4447), .ZN(n2413) );
  NAND2_X1 U2800 ( .A1(n4501), .A2(n2416), .ZN(n4486) );
  NAND2_X1 U2801 ( .A1(n4501), .A2(n4502), .ZN(n4485) );
  AND2_X1 U2802 ( .A1(n3030), .A2(n2420), .ZN(n2419) );
  NAND2_X1 U2803 ( .A1(n4576), .A2(n2420), .ZN(n4556) );
  NAND2_X1 U2804 ( .A1(n2728), .A2(n4269), .ZN(n4572) );
  NOR2_X1 U2805 ( .A1(n4631), .A2(n4149), .ZN(n4614) );
  OR2_X1 U2806 ( .A1(n3698), .A2(n3823), .ZN(n4631) );
  NAND2_X1 U2807 ( .A1(n3577), .A2(n2418), .ZN(n3651) );
  AND2_X1 U2808 ( .A1(n2132), .A2(n3684), .ZN(n2418) );
  NAND2_X1 U2809 ( .A1(n3577), .A2(n2132), .ZN(n4664) );
  INV_X1 U2810 ( .A(n3466), .ZN(n3470) );
  INV_X1 U2811 ( .A(n2392), .ZN(n2391) );
  NAND2_X1 U2812 ( .A1(n3290), .A2(n2579), .ZN(n3307) );
  OR2_X1 U2813 ( .A1(n3280), .A2(n2870), .ZN(n2874) );
  AND2_X1 U2814 ( .A1(n4904), .A2(n2883), .ZN(n4963) );
  INV_X1 U2815 ( .A(IR_REG_25__SCAN_IN), .ZN(n2846) );
  OR2_X1 U2816 ( .A1(n2844), .A2(IR_REG_25__SCAN_IN), .ZN(n2850) );
  XNOR2_X1 U2817 ( .A(n2854), .B(n2853), .ZN(n3151) );
  XNOR2_X1 U2818 ( .A(n2528), .B(n2527), .ZN(n2883) );
  NAND2_X1 U2819 ( .A1(n2837), .A2(IR_REG_31__SCAN_IN), .ZN(n2528) );
  INV_X1 U2820 ( .A(IR_REG_16__SCAN_IN), .ZN(n2509) );
  NOR2_X1 U2821 ( .A1(n2521), .A2(IR_REG_13__SCAN_IN), .ZN(n2511) );
  XNOR2_X1 U2822 ( .A(n2471), .B(IR_REG_6__SCAN_IN), .ZN(n3243) );
  NAND2_X1 U2823 ( .A1(n2216), .A2(n2217), .ZN(n3752) );
  NAND2_X1 U2824 ( .A1(n3752), .A2(n3751), .ZN(n3750) );
  NAND2_X1 U2825 ( .A1(n2395), .A2(n4154), .ZN(n3762) );
  NAND2_X1 U2826 ( .A1(n2395), .A2(n2393), .ZN(n3101) );
  NOR2_X1 U2827 ( .A1(n3761), .A2(n2394), .ZN(n2393) );
  INV_X1 U2828 ( .A(n4154), .ZN(n2394) );
  NAND2_X1 U2829 ( .A1(n3750), .A2(n2928), .ZN(n3352) );
  INV_X1 U2830 ( .A(n2810), .ZN(n4557) );
  INV_X1 U2831 ( .A(n4632), .ZN(n3823) );
  CLKBUF_X1 U2832 ( .A(n3263), .Z(n3264) );
  AND2_X1 U2833 ( .A1(n3714), .A2(n3715), .ZN(n2905) );
  OAI21_X1 U2834 ( .B1(n3752), .B2(n2387), .A(n2385), .ZN(n3407) );
  NAND2_X1 U2835 ( .A1(n2943), .A2(n2945), .ZN(n2946) );
  INV_X1 U2836 ( .A(n2999), .ZN(n3001) );
  AND2_X1 U2837 ( .A1(n2219), .A2(n2914), .ZN(n3274) );
  NAND2_X1 U2838 ( .A1(n3254), .A2(n3253), .ZN(n2219) );
  INV_X1 U2839 ( .A(n4536), .ZN(n4340) );
  NAND2_X1 U2840 ( .A1(n2572), .A2(n2571), .ZN(n4552) );
  NAND2_X1 U2841 ( .A1(n2742), .A2(n2741), .ZN(n4534) );
  OR2_X1 U2842 ( .A1(n4559), .A2(n2771), .ZN(n2742) );
  INV_X1 U2843 ( .A(n4550), .ZN(n4593) );
  INV_X1 U2844 ( .A(n4624), .ZN(n3820) );
  NAND2_X1 U2845 ( .A1(n2699), .A2(n2698), .ZN(n4629) );
  OAI211_X1 U2846 ( .C1(n3617), .C2(n2771), .A(n2683), .B(n2682), .ZN(n4659)
         );
  OR2_X1 U2847 ( .A1(n2678), .A2(n2677), .ZN(n3589) );
  INV_X1 U2848 ( .A(n3495), .ZN(n4344) );
  INV_X1 U2849 ( .A(n3353), .ZN(n3397) );
  INV_X1 U2850 ( .A(n3716), .ZN(n4345) );
  INV_X1 U2851 ( .A(n3420), .ZN(n4346) );
  CLKBUF_X1 U2852 ( .A(U4043), .Z(n3562) );
  NAND2_X1 U2853 ( .A1(n3162), .A2(n3161), .ZN(n4349) );
  OR2_X1 U2854 ( .A1(n3169), .A2(REG2_REG_1__SCAN_IN), .ZN(n3162) );
  NAND2_X1 U2855 ( .A1(n4873), .A2(n2360), .ZN(n4367) );
  XNOR2_X1 U2856 ( .A(n3196), .B(n3195), .ZN(n4818) );
  AND2_X1 U2857 ( .A1(n2371), .A2(n2373), .ZN(n3239) );
  NOR2_X1 U2858 ( .A1(n3385), .A2(n3384), .ZN(n3387) );
  INV_X1 U2859 ( .A(n2377), .ZN(n3384) );
  INV_X1 U2860 ( .A(n3378), .ZN(n3381) );
  NAND2_X1 U2861 ( .A1(n2486), .A2(n2489), .ZN(n3437) );
  XNOR2_X1 U2862 ( .A(n3547), .B(n3555), .ZN(n3548) );
  INV_X1 U2863 ( .A(n2301), .ZN(n3549) );
  NAND2_X1 U2864 ( .A1(n4380), .A2(n4379), .ZN(n4835) );
  NAND2_X1 U2865 ( .A1(n4394), .A2(n4393), .ZN(n4829) );
  AND2_X1 U2866 ( .A1(n3176), .A2(n3175), .ZN(n4849) );
  AND2_X1 U2867 ( .A1(n3176), .A2(n4333), .ZN(n4875) );
  NAND2_X1 U2868 ( .A1(n2200), .A2(n2777), .ZN(n4446) );
  NAND2_X1 U2869 ( .A1(n2265), .A2(n2269), .ZN(n4494) );
  NAND2_X1 U2870 ( .A1(n4530), .A2(n2270), .ZN(n2265) );
  NAND2_X1 U2871 ( .A1(n4530), .A2(n2273), .ZN(n4509) );
  NAND2_X1 U2872 ( .A1(n4611), .A2(n2719), .ZN(n4584) );
  NAND2_X1 U2873 ( .A1(n3654), .A2(n4209), .ZN(n3693) );
  AND2_X1 U2874 ( .A1(n2194), .A2(n2149), .ZN(n3691) );
  OAI22_X1 U2875 ( .A1(n3569), .A2(n4647), .B1(n4645), .B2(n2190), .ZN(n3573)
         );
  AND2_X1 U2876 ( .A1(n4668), .A2(n4812), .ZN(n4618) );
  AND2_X1 U2877 ( .A1(n4618), .A2(n4972), .ZN(n4896) );
  INV_X1 U2878 ( .A(n4665), .ZN(n4912) );
  AOI21_X1 U2879 ( .B1(n4430), .B2(n4972), .A(n2565), .ZN(n2836) );
  NOR2_X1 U2880 ( .A1(n3577), .A2(n2190), .ZN(n3578) );
  INV_X1 U2881 ( .A(IR_REG_30__SCAN_IN), .ZN(n3961) );
  INV_X1 U2882 ( .A(n2551), .ZN(n4789) );
  AND2_X2 U2883 ( .A1(n2550), .A2(n2549), .ZN(n3136) );
  NAND2_X1 U2884 ( .A1(n2548), .A2(n2547), .ZN(n2550) );
  NAND2_X1 U2885 ( .A1(IR_REG_31__SCAN_IN), .A2(n2546), .ZN(n2547) );
  XNOR2_X1 U2886 ( .A(n2851), .B(IR_REG_26__SCAN_IN), .ZN(n4791) );
  NAND2_X1 U2887 ( .A1(n2850), .A2(IR_REG_31__SCAN_IN), .ZN(n2851) );
  NAND2_X1 U2888 ( .A1(n2849), .A2(n2850), .ZN(n3135) );
  NAND2_X1 U2889 ( .A1(n2848), .A2(n2847), .ZN(n2849) );
  NAND2_X1 U2890 ( .A1(IR_REG_31__SCAN_IN), .A2(n2846), .ZN(n2847) );
  NAND2_X1 U2891 ( .A1(n2845), .A2(IR_REG_25__SCAN_IN), .ZN(n2848) );
  AND2_X1 U2892 ( .A1(n3151), .A2(STATE_REG_SCAN_IN), .ZN(n4931) );
  INV_X1 U2893 ( .A(n2883), .ZN(n4792) );
  AND2_X1 U2894 ( .A1(n2533), .A2(n2524), .ZN(n4802) );
  AND2_X1 U2895 ( .A1(n2506), .A2(n2505), .ZN(n4937) );
  XNOR2_X1 U2896 ( .A(n2497), .B(IR_REG_12__SCAN_IN), .ZN(n4794) );
  XNOR2_X1 U2897 ( .A(n2463), .B(IR_REG_4__SCAN_IN), .ZN(n4820) );
  INV_X1 U2898 ( .A(n3191), .ZN(n3178) );
  INV_X1 U2899 ( .A(n3169), .ZN(n4798) );
  XNOR2_X1 U2900 ( .A(n2222), .B(n2168), .ZN(n4160) );
  NOR2_X1 U2901 ( .A1(n4887), .A2(n2365), .ZN(n3202) );
  NAND2_X1 U2902 ( .A1(n2214), .A2(n2213), .ZN(n4890) );
  NAND2_X1 U2903 ( .A1(n4888), .A2(n4889), .ZN(n2214) );
  INV_X1 U2904 ( .A(n2309), .ZN(n2308) );
  OR2_X1 U2905 ( .A1(n3736), .A2(n4738), .ZN(n3113) );
  OR2_X1 U2906 ( .A1(n3736), .A2(n4787), .ZN(n3117) );
  AND2_X1 U2907 ( .A1(n2134), .A2(n4646), .ZN(n2132) );
  AND2_X1 U2908 ( .A1(n2391), .A2(n2390), .ZN(n2133) );
  AND2_X1 U2909 ( .A1(n3730), .A2(n2190), .ZN(n2134) );
  AND2_X1 U2910 ( .A1(n2183), .A2(n3253), .ZN(n2135) );
  AND2_X1 U2911 ( .A1(n2167), .A2(n4202), .ZN(n2347) );
  OR2_X1 U2912 ( .A1(n2218), .A2(n2915), .ZN(n2136) );
  AND2_X1 U2913 ( .A1(n2351), .A2(n2349), .ZN(n2137) );
  AND2_X1 U2914 ( .A1(n2235), .A2(REG3_REG_20__SCAN_IN), .ZN(n2138) );
  NOR2_X1 U2915 ( .A1(n4879), .A2(n2313), .ZN(n2139) );
  OR2_X1 U2916 ( .A1(n4859), .A2(n4843), .ZN(n2140) );
  INV_X2 U2917 ( .A(n3061), .ZN(n2919) );
  OAI21_X1 U2918 ( .B1(n3484), .B2(n2407), .A(n2405), .ZN(n3622) );
  NAND2_X1 U2919 ( .A1(n4576), .A2(n3843), .ZN(n4555) );
  AND2_X1 U2920 ( .A1(n2552), .A2(n4789), .ZN(n2142) );
  NAND2_X1 U2921 ( .A1(n2539), .A2(n2238), .ZN(n2143) );
  AND2_X1 U2922 ( .A1(n4379), .A2(n2306), .ZN(n2144) );
  AND2_X1 U2923 ( .A1(n2428), .A2(n4215), .ZN(n2145) );
  NOR2_X1 U2924 ( .A1(n3195), .A2(n2294), .ZN(n2146) );
  AND4_X1 U2925 ( .A1(n2522), .A2(n3852), .A3(n2509), .A4(n2253), .ZN(n2147)
         );
  NAND2_X1 U2926 ( .A1(n2538), .A2(n2235), .ZN(n2148) );
  AOI21_X1 U2927 ( .B1(n4147), .B2(n4145), .A(n4144), .ZN(n3778) );
  AND2_X1 U2928 ( .A1(n3837), .A2(n3841), .ZN(n3784) );
  NAND4_X1 U2929 ( .A1(n2577), .A2(n2576), .A3(n2575), .A4(n2574), .ZN(n2881)
         );
  NAND2_X1 U2930 ( .A1(n2317), .A2(n2316), .ZN(n2379) );
  NAND2_X1 U2931 ( .A1(n3805), .A2(n3650), .ZN(n2149) );
  OAI22_X1 U2932 ( .A1(n2131), .A2(n2190), .B1(n3727), .B2(n3061), .ZN(n2948)
         );
  AND3_X1 U2933 ( .A1(n2544), .A2(n3850), .A3(n2543), .ZN(n2150) );
  OR2_X1 U2934 ( .A1(n3204), .A2(n4030), .ZN(n2151) );
  NOR2_X1 U2935 ( .A1(n4841), .A2(n4399), .ZN(n2152) );
  AND2_X1 U2936 ( .A1(n3322), .A2(REG2_REG_7__SCAN_IN), .ZN(n2153) );
  OR2_X1 U2937 ( .A1(n3322), .A2(REG1_REG_7__SCAN_IN), .ZN(n2154) );
  INV_X1 U2938 ( .A(n2457), .ZN(n3150) );
  NAND2_X1 U2939 ( .A1(n4801), .A2(n2139), .ZN(n2155) );
  INV_X1 U2940 ( .A(n2657), .ZN(n2282) );
  OR2_X1 U2941 ( .A1(n3608), .A2(n2684), .ZN(n2156) );
  NAND2_X1 U2942 ( .A1(n4501), .A2(n2414), .ZN(n2417) );
  AND2_X1 U2943 ( .A1(n2367), .A2(REG1_REG_4__SCAN_IN), .ZN(n2157) );
  INV_X1 U2944 ( .A(n3189), .ZN(n2367) );
  AND2_X1 U2945 ( .A1(n2204), .A2(n2203), .ZN(n2279) );
  INV_X1 U2946 ( .A(IR_REG_31__SCAN_IN), .ZN(n2455) );
  INV_X1 U2947 ( .A(n2357), .ZN(n2356) );
  NAND2_X1 U2948 ( .A1(n4249), .A2(n2359), .ZN(n2357) );
  INV_X1 U2949 ( .A(IR_REG_29__SCAN_IN), .ZN(n2546) );
  INV_X1 U2950 ( .A(n2401), .ZN(n2400) );
  NAND2_X1 U2951 ( .A1(n3026), .A2(n3841), .ZN(n2401) );
  AND2_X1 U2952 ( .A1(n3028), .A2(n3785), .ZN(n2158) );
  NAND2_X1 U2953 ( .A1(n2940), .A2(n2939), .ZN(n2159) );
  AND2_X1 U2954 ( .A1(n4393), .A2(n2211), .ZN(n2160) );
  AND2_X1 U2955 ( .A1(n2674), .A2(n2673), .ZN(n2161) );
  NAND2_X1 U2956 ( .A1(n4343), .A2(n3470), .ZN(n2162) );
  AND2_X1 U2957 ( .A1(n2727), .A2(n2719), .ZN(n2163) );
  AND2_X1 U2958 ( .A1(n4829), .A2(n4395), .ZN(n2164) );
  NOR2_X1 U2959 ( .A1(n2384), .A2(n2387), .ZN(n2383) );
  AND2_X1 U2960 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2165) );
  NAND2_X1 U2961 ( .A1(n3577), .A2(n2134), .ZN(n3598) );
  NAND2_X1 U2962 ( .A1(n3432), .A2(REG1_REG_9__SCAN_IN), .ZN(n2166) );
  NAND2_X1 U2963 ( .A1(n2257), .A2(n2592), .ZN(n3338) );
  INV_X1 U2964 ( .A(n4203), .ZN(n2335) );
  NAND2_X1 U2965 ( .A1(n4345), .A2(n3255), .ZN(n2167) );
  INV_X1 U2966 ( .A(n4269), .ZN(n2196) );
  INV_X1 U2967 ( .A(n4445), .ZN(n2349) );
  AND2_X1 U2968 ( .A1(n4154), .A2(n4153), .ZN(n2168) );
  OR2_X1 U2969 ( .A1(n2799), .A2(n2798), .ZN(n2169) );
  INV_X1 U2970 ( .A(n4212), .ZN(n2334) );
  INV_X1 U2971 ( .A(n4207), .ZN(n2330) );
  AND2_X1 U2972 ( .A1(n4536), .A2(n4523), .ZN(n2170) );
  AND2_X1 U2973 ( .A1(n3041), .A2(n3042), .ZN(n2171) );
  NOR2_X1 U2974 ( .A1(n3387), .A2(n3386), .ZN(n2172) );
  OR2_X1 U2975 ( .A1(n4463), .A2(n2815), .ZN(n2173) );
  AND2_X1 U2976 ( .A1(n4153), .A2(n2396), .ZN(n2174) );
  AND2_X1 U2977 ( .A1(n2777), .A2(n2173), .ZN(n2175) );
  INV_X1 U2978 ( .A(n2210), .ZN(n2209) );
  NOR2_X1 U2979 ( .A1(n4395), .A2(n4396), .ZN(n2210) );
  AND2_X1 U2980 ( .A1(n3438), .A2(REG2_REG_10__SCAN_IN), .ZN(n2176) );
  AND2_X1 U2981 ( .A1(n2776), .A2(n2775), .ZN(n4437) );
  INV_X1 U2982 ( .A(n2269), .ZN(n2268) );
  NAND2_X1 U2983 ( .A1(n2272), .A2(n2170), .ZN(n2269) );
  INV_X1 U2984 ( .A(n3030), .ZN(n4542) );
  AND2_X1 U2985 ( .A1(n2348), .A2(n2167), .ZN(n2177) );
  INV_X1 U2986 ( .A(n3684), .ZN(n3615) );
  NAND2_X1 U2987 ( .A1(n4795), .A2(REG2_REG_11__SCAN_IN), .ZN(n2178) );
  INV_X1 U2988 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4077) );
  AND2_X1 U2989 ( .A1(REG3_REG_11__SCAN_IN), .A2(REG3_REG_12__SCAN_IN), .ZN(
        n2179) );
  INV_X1 U2990 ( .A(REG3_REG_20__SCAN_IN), .ZN(n2237) );
  INV_X1 U2991 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2236) );
  NAND2_X1 U2992 ( .A1(n4807), .A2(REG2_REG_18__SCAN_IN), .ZN(n2180) );
  XNOR2_X1 U2993 ( .A(n2887), .B(n2888), .ZN(n3228) );
  AND2_X1 U2994 ( .A1(n3176), .A2(n4358), .ZN(n4873) );
  AND2_X1 U2995 ( .A1(n2957), .A2(n2956), .ZN(n2181) );
  INV_X1 U2996 ( .A(n4859), .ZN(n2375) );
  NOR2_X1 U2997 ( .A1(n4889), .A2(n2381), .ZN(n2182) );
  INV_X1 U2998 ( .A(REG3_REG_24__SCAN_IN), .ZN(n2241) );
  INV_X1 U2999 ( .A(n4144), .ZN(n2231) );
  INV_X1 U3000 ( .A(n3831), .ZN(n4502) );
  AND2_X1 U3001 ( .A1(n4177), .A2(DATAI_24_), .ZN(n3831) );
  NAND2_X1 U3002 ( .A1(n2924), .A2(n2923), .ZN(n2183) );
  INV_X1 U3003 ( .A(n4193), .ZN(n2345) );
  INV_X1 U3004 ( .A(n2815), .ZN(n4447) );
  AND2_X1 U3005 ( .A1(n2239), .A2(REG3_REG_27__SCAN_IN), .ZN(n2184) );
  OR2_X1 U3006 ( .A1(n3424), .A2(n3425), .ZN(n2185) );
  XOR2_X1 U3007 ( .A(n4802), .B(REG2_REG_19__SCAN_IN), .Z(n2186) );
  INV_X1 U3008 ( .A(n2296), .ZN(n3197) );
  INV_X1 U3009 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2294) );
  NOR2_X2 U3010 ( .A1(n3246), .A2(n3245), .ZN(n3318) );
  NAND2_X1 U3011 ( .A1(n3376), .A2(REG2_REG_8__SCAN_IN), .ZN(n2315) );
  AOI21_X1 U3012 ( .B1(n4880), .B2(n4879), .A(n4878), .ZN(n4886) );
  NAND2_X1 U3013 ( .A1(n3150), .A2(n3640), .ZN(n2192) );
  NAND2_X1 U3014 ( .A1(n4547), .A2(n2743), .ZN(n2198) );
  AND2_X2 U3015 ( .A1(n2205), .A2(n2438), .ZN(n2444) );
  NAND2_X1 U3016 ( .A1(n2206), .A2(REG1_REG_4__SCAN_IN), .ZN(n2364) );
  XNOR2_X1 U3017 ( .A(n2206), .B(n4987), .ZN(n4817) );
  INV_X1 U3018 ( .A(n2382), .ZN(n2220) );
  NAND3_X1 U3019 ( .A1(n2216), .A2(n2217), .A3(n2383), .ZN(n2221) );
  INV_X1 U3020 ( .A(n3706), .ZN(n3032) );
  NAND2_X1 U3021 ( .A1(n2538), .A2(n2234), .ZN(n2737) );
  NAND2_X1 U3022 ( .A1(n2539), .A2(n2239), .ZN(n2778) );
  NAND2_X1 U3023 ( .A1(n2539), .A2(n2184), .ZN(n2780) );
  NAND2_X1 U3024 ( .A1(n2539), .A2(REG3_REG_24__SCAN_IN), .ZN(n2761) );
  INV_X1 U3025 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2242) );
  NAND2_X1 U3026 ( .A1(n2243), .A2(n2179), .ZN(n2675) );
  NAND2_X1 U3027 ( .A1(n2244), .A2(n2165), .ZN(n2651) );
  INV_X1 U3028 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2246) );
  NAND4_X1 U3029 ( .A1(n4291), .A2(n4292), .A3(n4290), .A4(n2250), .ZN(n2249)
         );
  NAND3_X1 U3030 ( .A1(n4264), .A2(n4911), .A3(n4263), .ZN(n2251) );
  NAND3_X1 U3031 ( .A1(n2257), .A2(n2254), .A3(n2256), .ZN(n2609) );
  NOR2_X1 U3032 ( .A1(n4272), .A2(n2255), .ZN(n2254) );
  NAND3_X1 U3033 ( .A1(n3290), .A2(n2579), .A3(n2258), .ZN(n3305) );
  NAND2_X1 U3034 ( .A1(n3287), .A2(n3288), .ZN(n3290) );
  AND2_X1 U3035 ( .A1(n2527), .A2(n2526), .ZN(n2262) );
  NAND2_X1 U3036 ( .A1(n4611), .A2(n2163), .ZN(n2728) );
  OAI22_X2 U3037 ( .A1(n4530), .A2(n2264), .B1(n2266), .B2(n2263), .ZN(n4475)
         );
  AOI21_X2 U3038 ( .B1(n4475), .B2(n2769), .A(n2768), .ZN(n4455) );
  OR2_X1 U3039 ( .A1(n4516), .A2(n3030), .ZN(n2273) );
  NAND2_X1 U3040 ( .A1(n2551), .A2(REG0_REG_1__SCAN_IN), .ZN(n2288) );
  NAND3_X1 U3041 ( .A1(n2573), .A2(n2289), .A3(n2284), .ZN(n2578) );
  NAND2_X1 U3042 ( .A1(n2552), .A2(n2551), .ZN(n2285) );
  NAND2_X1 U3043 ( .A1(n4789), .A2(REG2_REG_1__SCAN_IN), .ZN(n2287) );
  NAND3_X1 U3044 ( .A1(n3136), .A2(n4789), .A3(REG3_REG_1__SCAN_IN), .ZN(n2289) );
  NAND2_X1 U3045 ( .A1(n3196), .A2(n2293), .ZN(n2290) );
  INV_X1 U3046 ( .A(n2303), .ZN(n3636) );
  AND2_X2 U3047 ( .A1(n2303), .A2(n2178), .ZN(n4378) );
  NOR2_X2 U3048 ( .A1(n4845), .A2(n4846), .ZN(n4844) );
  XNOR2_X2 U3049 ( .A(n4381), .B(n4397), .ZN(n4845) );
  NAND2_X1 U3050 ( .A1(n4801), .A2(n2310), .ZN(n2307) );
  OAI211_X1 U3051 ( .C1(n4801), .C2(n2311), .A(n2307), .B(n2308), .ZN(n4816)
         );
  NAND2_X1 U3052 ( .A1(n4801), .A2(n4800), .ZN(n4880) );
  INV_X1 U3053 ( .A(n4800), .ZN(n2313) );
  NOR2_X2 U3054 ( .A1(n3318), .A2(n2153), .ZN(n3374) );
  NAND2_X1 U3055 ( .A1(n2649), .A2(n2648), .ZN(n3524) );
  NAND2_X1 U3056 ( .A1(n3305), .A2(n2584), .ZN(n3360) );
  NAND2_X1 U3057 ( .A1(n2578), .A2(n3286), .ZN(n4180) );
  NAND2_X1 U3058 ( .A1(n4372), .A2(n3166), .ZN(n3192) );
  NAND2_X1 U3059 ( .A1(n4180), .A2(n4182), .ZN(n3287) );
  NAND2_X1 U3060 ( .A1(n3328), .A2(n2625), .ZN(n3393) );
  XNOR2_X1 U3061 ( .A(n2321), .B(n2320), .ZN(n3343) );
  INV_X1 U3062 ( .A(n4272), .ZN(n2320) );
  OAI21_X1 U3063 ( .B1(n3465), .B2(n2332), .A(n2329), .ZN(n3586) );
  NAND2_X1 U3064 ( .A1(n2328), .A2(n2327), .ZN(n2803) );
  NAND2_X1 U3065 ( .A1(n3465), .A2(n2329), .ZN(n2328) );
  OAI21_X1 U3066 ( .B1(n3465), .B2(n4203), .A(n4199), .ZN(n3520) );
  AOI21_X1 U3067 ( .B1(n4203), .B2(n4199), .A(n2334), .ZN(n2333) );
  NAND2_X1 U3068 ( .A1(n2344), .A2(n2341), .ZN(n2796) );
  NAND2_X1 U3069 ( .A1(n2812), .A2(n4307), .ZN(n2358) );
  AND2_X1 U3070 ( .A1(n2361), .A2(n4365), .ZN(n2360) );
  NAND2_X1 U3071 ( .A1(n3172), .A2(n3173), .ZN(n2361) );
  OR2_X1 U3072 ( .A1(n3207), .A2(n2366), .ZN(n2365) );
  NOR2_X1 U3073 ( .A1(n2368), .A2(n2367), .ZN(n2366) );
  NAND2_X1 U3074 ( .A1(n3237), .A2(REG1_REG_6__SCAN_IN), .ZN(n2371) );
  NAND2_X1 U3075 ( .A1(n2371), .A2(n2370), .ZN(n3321) );
  NAND2_X1 U3076 ( .A1(n3236), .A2(n3243), .ZN(n2373) );
  NAND2_X1 U3077 ( .A1(n4399), .A2(n2375), .ZN(n2374) );
  NAND2_X1 U3078 ( .A1(n2379), .A2(IR_REG_31__SCAN_IN), .ZN(n2456) );
  INV_X1 U3079 ( .A(n2379), .ZN(n2460) );
  NAND2_X1 U3080 ( .A1(n2380), .A2(n4808), .ZN(n4809) );
  NAND2_X1 U3081 ( .A1(n4805), .A2(n4804), .ZN(n4888) );
  INV_X1 U3082 ( .A(n4804), .ZN(n2381) );
  NAND2_X1 U3083 ( .A1(n3366), .A2(n3717), .ZN(n3424) );
  INV_X1 U3084 ( .A(n3424), .ZN(n2390) );
  NAND2_X1 U3085 ( .A1(n3754), .A2(n2390), .ZN(n2389) );
  INV_X1 U3086 ( .A(n3255), .ZN(n3425) );
  INV_X1 U3087 ( .A(n3795), .ZN(n2396) );
  NAND2_X1 U3088 ( .A1(n3484), .A2(n2405), .ZN(n2402) );
  NAND2_X1 U3089 ( .A1(n2402), .A2(n2403), .ZN(n2978) );
  NAND2_X1 U3090 ( .A1(n4501), .A2(n2413), .ZN(n3109) );
  INV_X1 U3091 ( .A(n2417), .ZN(n4466) );
  NAND2_X1 U3092 ( .A1(n4576), .A2(n2419), .ZN(n4521) );
  NAND2_X1 U3093 ( .A1(n4871), .A2(n4870), .ZN(n4869) );
  NAND2_X1 U3094 ( .A1(n3644), .A2(REG1_REG_12__SCAN_IN), .ZN(n4394) );
  XNOR2_X1 U3095 ( .A(n4392), .B(n4377), .ZN(n3644) );
  AOI21_X1 U3096 ( .B1(n4814), .B2(n4873), .A(n4813), .ZN(n4815) );
  NOR2_X2 U3097 ( .A1(n4853), .A2(n4383), .ZN(n4385) );
  XNOR2_X1 U3098 ( .A(n2886), .B(n3055), .ZN(n2888) );
  INV_X1 U3099 ( .A(n4858), .ZN(n4401) );
  NAND2_X1 U3100 ( .A1(n3705), .A2(n3036), .ZN(n3771) );
  NAND2_X1 U3101 ( .A1(n2459), .A2(n2458), .ZN(n3367) );
  NAND2_X1 U3102 ( .A1(n3771), .A2(n2171), .ZN(n3828) );
  AND2_X1 U3103 ( .A1(n2889), .A2(n2888), .ZN(n2890) );
  INV_X1 U3104 ( .A(n2889), .ZN(n2887) );
  NAND2_X1 U3105 ( .A1(n2844), .A2(IR_REG_31__SCAN_IN), .ZN(n2845) );
  NAND2_X1 U3106 ( .A1(n3444), .A2(n2946), .ZN(n3484) );
  INV_X1 U3107 ( .A(n3285), .ZN(n2459) );
  AOI22_X2 U3108 ( .A1(n3244), .A2(REG2_REG_6__SCAN_IN), .B1(n3243), .B2(n3242), .ZN(n3246) );
  INV_X1 U3109 ( .A(n4438), .ZN(n4441) );
  NOR2_X2 U3110 ( .A1(n4438), .A2(n2816), .ZN(n3103) );
  OAI22_X1 U3111 ( .A1(n2880), .A2(n2986), .B1(n3058), .B2(n4903), .ZN(n2884)
         );
  OAI22_X1 U3112 ( .A1(n2885), .A2(n3061), .B1(n3286), .B2(n2131), .ZN(n2889)
         );
  NAND2_X1 U3113 ( .A1(n2885), .A2(n3291), .ZN(n4182) );
  AOI21_X2 U3114 ( .B1(n3002), .B2(n3001), .A(n3000), .ZN(n4147) );
  INV_X2 U3115 ( .A(n4991), .ZN(n4994) );
  AND2_X2 U3116 ( .A1(n3284), .A2(n4665), .ZN(n4643) );
  OR2_X1 U3117 ( .A1(n3556), .A2(n3555), .ZN(n2421) );
  NAND2_X1 U3118 ( .A1(n4937), .A2(REG1_REG_15__SCAN_IN), .ZN(n2422) );
  AND3_X1 U3119 ( .A1(n4288), .A2(n4287), .A3(n2428), .ZN(n2423) );
  AND2_X1 U3120 ( .A1(n4345), .A2(n3425), .ZN(n2424) );
  XOR2_X1 U3121 ( .A(n4812), .B(REG1_REG_19__SCAN_IN), .Z(n2425) );
  INV_X1 U3122 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2679) );
  NOR2_X1 U3123 ( .A1(n2500), .A2(n2511), .ZN(n4941) );
  INV_X1 U3124 ( .A(n3555), .ZN(n3438) );
  AND2_X1 U3125 ( .A1(n3094), .A2(n4140), .ZN(n2426) );
  AND4_X1 U3126 ( .A1(n4460), .A2(n4478), .A3(n4261), .A4(n4260), .ZN(n2427)
         );
  AND2_X1 U3127 ( .A1(n4216), .A2(n4209), .ZN(n2428) );
  NAND2_X1 U3128 ( .A1(n2692), .A2(n3610), .ZN(n2430) );
  OR2_X1 U3129 ( .A1(n4437), .A2(n4467), .ZN(n2431) );
  INV_X1 U3130 ( .A(n4467), .ZN(n4155) );
  NOR2_X1 U3131 ( .A1(n2607), .A2(n3415), .ZN(n2432) );
  INV_X1 U3132 ( .A(n4259), .ZN(n4260) );
  OR2_X1 U3133 ( .A1(n3676), .A2(n3675), .ZN(n2968) );
  AND2_X1 U3134 ( .A1(n4289), .A2(n2423), .ZN(n4290) );
  OR2_X1 U3135 ( .A1(n3753), .A2(n3332), .ZN(n2624) );
  INV_X1 U3136 ( .A(IR_REG_21__SCAN_IN), .ZN(n2526) );
  OAI22_X1 U3137 ( .A1(n2885), .A2(n2986), .B1(n3286), .B2(n3058), .ZN(n2886)
         );
  INV_X1 U3138 ( .A(n2944), .ZN(n2945) );
  INV_X1 U3139 ( .A(n2976), .ZN(n2977) );
  INV_X1 U3140 ( .A(n3437), .ZN(n3432) );
  OR2_X1 U3141 ( .A1(n4579), .A2(n2771), .ZN(n2734) );
  XNOR2_X1 U3142 ( .A(n3184), .B(n3178), .ZN(n3183) );
  NAND2_X1 U3143 ( .A1(n4807), .A2(REG1_REG_18__SCAN_IN), .ZN(n4808) );
  INV_X1 U3144 ( .A(n4645), .ZN(n4568) );
  INV_X1 U3145 ( .A(n4523), .ZN(n2752) );
  NAND2_X1 U3146 ( .A1(n2610), .A2(REG3_REG_7__SCAN_IN), .ZN(n2634) );
  INV_X1 U3147 ( .A(n4343), .ZN(n3447) );
  NAND2_X1 U31480 ( .A1(n2908), .A2(n2907), .ZN(n2909) );
  AND2_X1 U31490 ( .A1(n3816), .A2(n3817), .ZN(n3000) );
  INV_X1 U3150 ( .A(n3845), .ZN(n4169) );
  OR2_X1 U3151 ( .A1(n4504), .A2(n2771), .ZN(n2759) );
  NAND2_X1 U3152 ( .A1(n3169), .A2(REG1_REG_1__SCAN_IN), .ZN(n3170) );
  INV_X1 U3153 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3853) );
  INV_X1 U3154 ( .A(n4882), .ZN(n4883) );
  INV_X1 U3155 ( .A(n4534), .ZN(n4570) );
  AND2_X1 U3156 ( .A1(n4327), .A2(n4792), .ZN(n3152) );
  INV_X1 U3157 ( .A(n4288), .ZN(n2700) );
  OAI21_X1 U3158 ( .B1(n3287), .B2(n4257), .A(n4182), .ZN(n3309) );
  INV_X1 U3159 ( .A(REG1_REG_2__SCAN_IN), .ZN(n4018) );
  INV_X1 U3160 ( .A(n3590), .ZN(n3730) );
  INV_X1 U3161 ( .A(n2626), .ZN(n3754) );
  INV_X1 U3162 ( .A(n4660), .ZN(n4908) );
  AND2_X1 U3163 ( .A1(n2476), .A2(n2477), .ZN(n3322) );
  AND2_X1 U3164 ( .A1(n3095), .A2(n2426), .ZN(n3076) );
  NAND2_X1 U3165 ( .A1(n3713), .A2(n2909), .ZN(n3254) );
  INV_X1 U3166 ( .A(n4175), .ZN(n4140) );
  INV_X1 U3167 ( .A(n4802), .ZN(n4812) );
  NAND2_X1 U3168 ( .A1(n2759), .A2(n2758), .ZN(n4518) );
  AND2_X1 U3169 ( .A1(n3155), .A2(n3154), .ZN(n3176) );
  NAND2_X1 U3170 ( .A1(n4884), .A2(n4883), .ZN(n4885) );
  NAND2_X1 U3171 ( .A1(n2726), .A2(n2725), .ZN(n4610) );
  INV_X1 U3172 ( .A(n4603), .ZN(n4640) );
  OR2_X1 U3173 ( .A1(n3088), .A2(n3149), .ZN(n4665) );
  NAND2_X1 U3174 ( .A1(n2820), .A2(n2819), .ZN(n4906) );
  AND2_X1 U3175 ( .A1(n4668), .A2(n3301), .ZN(n4913) );
  OAI21_X1 U3176 ( .B1(n3141), .B2(D_REG_0__SCAN_IN), .A(n3143), .ZN(n3281) );
  INV_X1 U3177 ( .A(n3009), .ZN(n4597) );
  AND2_X1 U3178 ( .A1(n4905), .A2(n4954), .ZN(n4967) );
  NAND2_X1 U3179 ( .A1(n4791), .A2(n2857), .ZN(n3141) );
  XNOR2_X1 U3180 ( .A(n2479), .B(n2478), .ZN(n3373) );
  AND2_X1 U3181 ( .A1(n3155), .A2(n3153), .ZN(n4881) );
  INV_X1 U3182 ( .A(n4518), .ZN(n4480) );
  INV_X1 U3183 ( .A(n4166), .ZN(n4137) );
  OR2_X1 U3184 ( .A1(n3087), .A2(n3072), .ZN(n4175) );
  INV_X1 U3185 ( .A(n4437), .ZN(n4482) );
  INV_X1 U3186 ( .A(n4605), .ZN(n4341) );
  AOI21_X1 U3187 ( .B1(n4886), .B2(n2155), .A(n4885), .ZN(n4891) );
  NAND2_X1 U3188 ( .A1(n4668), .A2(n3414), .ZN(n4603) );
  NAND2_X1 U3189 ( .A1(n4994), .A2(n4972), .ZN(n4738) );
  OR2_X1 U3190 ( .A1(n2874), .A2(n3281), .ZN(n4991) );
  OR2_X1 U3191 ( .A1(n4777), .A2(n2876), .ZN(n2877) );
  NAND2_X1 U3192 ( .A1(n4777), .A2(n4972), .ZN(n4787) );
  INV_X1 U3193 ( .A(n4777), .ZN(n4980) );
  INV_X1 U3194 ( .A(n4928), .ZN(n4930) );
  NAND2_X1 U3195 ( .A1(n3142), .A2(n3141), .ZN(n4928) );
  INV_X1 U3196 ( .A(n2843), .ZN(n2441) );
  NAND2_X1 U3197 ( .A1(n2544), .A2(n3850), .ZN(n2450) );
  NAND3_X1 U3198 ( .A1(n2844), .A2(IR_REG_27__SCAN_IN), .A3(IR_REG_31__SCAN_IN), .ZN(n2449) );
  INV_X1 U3199 ( .A(n2544), .ZN(n2445) );
  NAND2_X1 U3200 ( .A1(n2445), .A2(IR_REG_27__SCAN_IN), .ZN(n2446) );
  NAND2_X1 U3201 ( .A1(n2446), .A2(IR_REG_31__SCAN_IN), .ZN(n2447) );
  OAI21_X1 U3202 ( .B1(IR_REG_31__SCAN_IN), .B2(n3850), .A(n2447), .ZN(n2448)
         );
  OAI211_X1 U3203 ( .C1(n2844), .C2(n2450), .A(n2449), .B(n2448), .ZN(n2452)
         );
  NAND2_X1 U3204 ( .A1(n3850), .A2(IR_REG_27__SCAN_IN), .ZN(n2451) );
  AND2_X1 U3205 ( .A1(n4177), .A2(DATAI_29_), .ZN(n4237) );
  NAND2_X1 U3206 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2453)
         );
  MUX2_X1 U3207 ( .A(n4798), .B(DATAI_1_), .S(n2457), .Z(n3291) );
  MUX2_X1 U3208 ( .A(IR_REG_0__SCAN_IN), .B(DATAI_0_), .S(n2457), .Z(n3747) );
  NAND2_X1 U3209 ( .A1(n3286), .A2(n4903), .ZN(n3285) );
  MUX2_X1 U32100 ( .A(n2130), .B(DATAI_2_), .S(n2457), .Z(n3314) );
  NAND2_X1 U32110 ( .A1(n2460), .A2(n3851), .ZN(n2467) );
  NAND2_X1 U32120 ( .A1(n2467), .A2(IR_REG_31__SCAN_IN), .ZN(n2461) );
  XNOR2_X1 U32130 ( .A(n2461), .B(IR_REG_3__SCAN_IN), .ZN(n3191) );
  MUX2_X1 U32140 ( .A(n3191), .B(DATAI_3_), .S(n4177), .Z(n3368) );
  NAND2_X1 U32150 ( .A1(n2461), .A2(n2464), .ZN(n2462) );
  NAND2_X1 U32160 ( .A1(n2462), .A2(IR_REG_31__SCAN_IN), .ZN(n2463) );
  MUX2_X1 U32170 ( .A(n4820), .B(DATAI_4_), .S(n4177), .Z(n2606) );
  INV_X1 U32180 ( .A(IR_REG_4__SCAN_IN), .ZN(n2465) );
  NAND2_X1 U32190 ( .A1(n2465), .A2(n2464), .ZN(n2466) );
  OAI21_X1 U32200 ( .B1(n2467), .B2(n2466), .A(IR_REG_31__SCAN_IN), .ZN(n2468)
         );
  MUX2_X1 U32210 ( .A(IR_REG_31__SCAN_IN), .B(n2468), .S(IR_REG_5__SCAN_IN), 
        .Z(n2469) );
  INV_X1 U32220 ( .A(DATAI_5_), .ZN(n2470) );
  MUX2_X1 U32230 ( .A(n3204), .B(n2470), .S(n4178), .Z(n3255) );
  NAND2_X1 U32240 ( .A1(n2472), .A2(IR_REG_31__SCAN_IN), .ZN(n2471) );
  MUX2_X1 U32250 ( .A(n3243), .B(DATAI_6_), .S(n4178), .Z(n3332) );
  OR2_X1 U32260 ( .A1(n2472), .A2(IR_REG_6__SCAN_IN), .ZN(n2480) );
  NAND2_X1 U32270 ( .A1(n2473), .A2(IR_REG_7__SCAN_IN), .ZN(n2476) );
  INV_X1 U32280 ( .A(n2473), .ZN(n2475) );
  INV_X1 U32290 ( .A(IR_REG_7__SCAN_IN), .ZN(n2474) );
  NAND2_X1 U32300 ( .A1(n2475), .A2(n2474), .ZN(n2477) );
  MUX2_X1 U32310 ( .A(n3322), .B(DATAI_7_), .S(n4177), .Z(n2626) );
  NAND2_X1 U32320 ( .A1(n2477), .A2(IR_REG_31__SCAN_IN), .ZN(n2479) );
  INV_X1 U32330 ( .A(DATAI_8_), .ZN(n3130) );
  MUX2_X1 U32340 ( .A(n3373), .B(n3130), .S(n4177), .Z(n3395) );
  NAND2_X1 U32350 ( .A1(n3401), .A2(n3395), .ZN(n3402) );
  INV_X1 U32360 ( .A(n2480), .ZN(n2482) );
  NOR2_X1 U32370 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2481)
         );
  NAND2_X1 U32380 ( .A1(n2482), .A2(n2481), .ZN(n2484) );
  NAND2_X1 U32390 ( .A1(n2484), .A2(IR_REG_31__SCAN_IN), .ZN(n2483) );
  MUX2_X1 U32400 ( .A(IR_REG_31__SCAN_IN), .B(n2483), .S(IR_REG_9__SCAN_IN), 
        .Z(n2486) );
  INV_X1 U32410 ( .A(n2484), .ZN(n2485) );
  INV_X1 U32420 ( .A(DATAI_9_), .ZN(n2487) );
  MUX2_X1 U32430 ( .A(n3437), .B(n2487), .S(n4177), .Z(n3466) );
  NAND2_X1 U32440 ( .A1(n2489), .A2(IR_REG_31__SCAN_IN), .ZN(n2488) );
  MUX2_X1 U32450 ( .A(IR_REG_31__SCAN_IN), .B(n2488), .S(IR_REG_10__SCAN_IN), 
        .Z(n2490) );
  NAND2_X1 U32460 ( .A1(n2490), .A2(n2491), .ZN(n3555) );
  INV_X1 U32470 ( .A(DATAI_10_), .ZN(n3933) );
  MUX2_X1 U32480 ( .A(n3555), .B(n3933), .S(n4178), .Z(n3449) );
  NOR2_X4 U32490 ( .A1(n3526), .A2(n3525), .ZN(n3577) );
  NAND2_X1 U32500 ( .A1(n2492), .A2(IR_REG_11__SCAN_IN), .ZN(n2495) );
  INV_X1 U32510 ( .A(n2492), .ZN(n2494) );
  INV_X1 U32520 ( .A(IR_REG_11__SCAN_IN), .ZN(n2493) );
  NAND2_X1 U32530 ( .A1(n2494), .A2(n2493), .ZN(n2496) );
  INV_X1 U32540 ( .A(DATAI_11_), .ZN(n3959) );
  NAND2_X1 U32550 ( .A1(n2496), .A2(IR_REG_31__SCAN_IN), .ZN(n2497) );
  MUX2_X1 U32560 ( .A(DATAI_12_), .B(n4794), .S(n3150), .Z(n3590) );
  NAND2_X1 U32570 ( .A1(n2521), .A2(IR_REG_31__SCAN_IN), .ZN(n2498) );
  MUX2_X1 U32580 ( .A(IR_REG_31__SCAN_IN), .B(n2498), .S(IR_REG_13__SCAN_IN), 
        .Z(n2499) );
  INV_X1 U32590 ( .A(n2499), .ZN(n2500) );
  MUX2_X1 U32600 ( .A(n4941), .B(DATAI_13_), .S(n4178), .Z(n4662) );
  OR2_X1 U32610 ( .A1(n2511), .A2(n2455), .ZN(n2501) );
  XNOR2_X1 U32620 ( .A(n2501), .B(IR_REG_14__SCAN_IN), .ZN(n4939) );
  INV_X1 U32630 ( .A(DATAI_14_), .ZN(n2502) );
  MUX2_X1 U32640 ( .A(n4397), .B(n2502), .S(n4177), .Z(n3684) );
  INV_X1 U32650 ( .A(IR_REG_14__SCAN_IN), .ZN(n2508) );
  NAND2_X1 U32660 ( .A1(n2511), .A2(n2508), .ZN(n2503) );
  NAND2_X1 U32670 ( .A1(n2503), .A2(IR_REG_31__SCAN_IN), .ZN(n2504) );
  NAND2_X1 U32680 ( .A1(n2504), .A2(n4022), .ZN(n2506) );
  OR2_X1 U32690 ( .A1(n2504), .A2(n4022), .ZN(n2505) );
  MUX2_X1 U32700 ( .A(n4937), .B(DATAI_15_), .S(n4178), .Z(n4172) );
  INV_X1 U32710 ( .A(DATAI_16_), .ZN(n4935) );
  NAND2_X1 U32720 ( .A1(n2506), .A2(IR_REG_31__SCAN_IN), .ZN(n2507) );
  XNOR2_X1 U32730 ( .A(n2509), .B(n2507), .ZN(n4936) );
  MUX2_X1 U32740 ( .A(n4935), .B(n4936), .S(n3150), .Z(n3806) );
  NAND2_X1 U32750 ( .A1(n3697), .A2(n3806), .ZN(n3698) );
  AND3_X1 U32760 ( .A1(n4022), .A2(n2509), .A3(n2508), .ZN(n2510) );
  NAND2_X1 U32770 ( .A1(n2511), .A2(n2510), .ZN(n2513) );
  NAND2_X1 U32780 ( .A1(n2513), .A2(IR_REG_31__SCAN_IN), .ZN(n2512) );
  MUX2_X1 U32790 ( .A(IR_REG_31__SCAN_IN), .B(n2512), .S(IR_REG_17__SCAN_IN), 
        .Z(n2514) );
  NAND2_X1 U32800 ( .A1(n2514), .A2(n2516), .ZN(n4391) );
  INV_X1 U32810 ( .A(DATAI_17_), .ZN(n2515) );
  MUX2_X1 U32820 ( .A(n4391), .B(n2515), .S(n4178), .Z(n4632) );
  NAND2_X1 U32830 ( .A1(n2516), .A2(IR_REG_31__SCAN_IN), .ZN(n2517) );
  XNOR2_X1 U32840 ( .A(n2517), .B(IR_REG_18__SCAN_IN), .ZN(n4807) );
  MUX2_X1 U32850 ( .A(n4807), .B(DATAI_18_), .S(n4178), .Z(n4149) );
  NOR2_X1 U32860 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U32870 ( .A1(n2519), .A2(n2518), .ZN(n2520) );
  OR2_X1 U32880 ( .A1(n2523), .A2(n2522), .ZN(n2524) );
  MUX2_X1 U32890 ( .A(n4802), .B(DATAI_19_), .S(n4178), .Z(n3009) );
  AND2_X2 U32900 ( .A1(n4614), .A2(n4597), .ZN(n4576) );
  NAND2_X1 U32910 ( .A1(n4177), .A2(DATAI_20_), .ZN(n3843) );
  NAND2_X1 U32920 ( .A1(n4178), .A2(DATAI_22_), .ZN(n3030) );
  NAND2_X1 U32930 ( .A1(n4177), .A2(DATAI_23_), .ZN(n4523) );
  NAND2_X1 U32940 ( .A1(n4177), .A2(DATAI_25_), .ZN(n4487) );
  INV_X1 U32950 ( .A(n4487), .ZN(n3047) );
  NAND2_X1 U32960 ( .A1(n4178), .A2(DATAI_26_), .ZN(n4467) );
  AND2_X1 U32970 ( .A1(n4178), .A2(DATAI_27_), .ZN(n2815) );
  AND2_X1 U32980 ( .A1(n4177), .A2(DATAI_28_), .ZN(n3091) );
  AOI21_X1 U32990 ( .B1(n4237), .B2(n3110), .A(n4418), .ZN(n4430) );
  NAND2_X1 U33000 ( .A1(n2529), .A2(n2526), .ZN(n2837) );
  INV_X1 U33010 ( .A(n2529), .ZN(n2530) );
  NAND2_X1 U33020 ( .A1(n2530), .A2(IR_REG_31__SCAN_IN), .ZN(n2531) );
  MUX2_X1 U33030 ( .A(IR_REG_31__SCAN_IN), .B(n2531), .S(IR_REG_21__SCAN_IN), 
        .Z(n2532) );
  INV_X1 U33040 ( .A(REG3_REG_22__SCAN_IN), .ZN(n2566) );
  INV_X1 U33050 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3773) );
  INV_X1 U33060 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4090) );
  INV_X1 U33070 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4072) );
  INV_X1 U33080 ( .A(n2780), .ZN(n2540) );
  NAND2_X1 U33090 ( .A1(n2540), .A2(REG3_REG_28__SCAN_IN), .ZN(n4432) );
  INV_X1 U33100 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2541) );
  NAND2_X1 U33110 ( .A1(n2780), .A2(n2541), .ZN(n2542) );
  NAND2_X1 U33120 ( .A1(n4432), .A2(n2542), .ZN(n3737) );
  OAI21_X1 U33130 ( .B1(n2824), .B2(n2455), .A(IR_REG_29__SCAN_IN), .ZN(n2548)
         );
  INV_X1 U33140 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4085) );
  NAND2_X1 U33150 ( .A1(n2585), .A2(REG0_REG_28__SCAN_IN), .ZN(n2554) );
  AND2_X4 U33160 ( .A1(n3136), .A2(n2551), .ZN(n2586) );
  NAND2_X1 U33170 ( .A1(n2586), .A2(REG1_REG_28__SCAN_IN), .ZN(n2553) );
  OAI211_X1 U33180 ( .C1(n4085), .C2(n2784), .A(n2554), .B(n2553), .ZN(n2555)
         );
  INV_X1 U33190 ( .A(n2555), .ZN(n2556) );
  NAND2_X1 U33200 ( .A1(n4444), .A2(n3091), .ZN(n4426) );
  XNOR2_X1 U33210 ( .A(n3300), .B(n4792), .ZN(n2558) );
  NAND2_X1 U33220 ( .A1(n2558), .A2(n4812), .ZN(n4905) );
  AND2_X1 U33230 ( .A1(n2855), .A2(n4802), .ZN(n4904) );
  INV_X1 U33240 ( .A(n4963), .ZN(n4954) );
  NOR2_X1 U33250 ( .A1(n4426), .A2(n4967), .ZN(n2564) );
  OR2_X1 U33260 ( .A1(n4432), .A2(n2771), .ZN(n2563) );
  INV_X1 U33270 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3905) );
  NAND2_X1 U33280 ( .A1(n3215), .A2(REG2_REG_29__SCAN_IN), .ZN(n2560) );
  NAND2_X1 U33290 ( .A1(n2585), .A2(REG0_REG_29__SCAN_IN), .ZN(n2559) );
  OAI211_X1 U33300 ( .C1(n2748), .C2(n3905), .A(n2560), .B(n2559), .ZN(n2561)
         );
  INV_X1 U33310 ( .A(n2561), .ZN(n2562) );
  NAND2_X1 U33320 ( .A1(n2737), .A2(n2566), .ZN(n2567) );
  AND2_X1 U33330 ( .A1(n2744), .A2(n2567), .ZN(n4541) );
  NAND2_X1 U33340 ( .A1(n4541), .A2(n2781), .ZN(n2572) );
  INV_X1 U33350 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4539) );
  NAND2_X1 U33360 ( .A1(n2586), .A2(REG1_REG_22__SCAN_IN), .ZN(n2569) );
  NAND2_X1 U33370 ( .A1(n2585), .A2(REG0_REG_22__SCAN_IN), .ZN(n2568) );
  OAI211_X1 U33380 ( .C1(n4539), .C2(n2784), .A(n2569), .B(n2568), .ZN(n2570)
         );
  INV_X1 U33390 ( .A(n2570), .ZN(n2571) );
  NAND2_X1 U33400 ( .A1(n2586), .A2(REG1_REG_1__SCAN_IN), .ZN(n2573) );
  NAND2_X1 U33410 ( .A1(n2585), .A2(REG0_REG_0__SCAN_IN), .ZN(n2577) );
  NAND2_X1 U33420 ( .A1(n2586), .A2(REG1_REG_0__SCAN_IN), .ZN(n2576) );
  NAND2_X1 U33430 ( .A1(n2781), .A2(REG3_REG_0__SCAN_IN), .ZN(n2575) );
  AND2_X1 U33440 ( .A1(n2881), .A2(n3747), .ZN(n3288) );
  NAND2_X1 U33450 ( .A1(n2578), .A2(n3291), .ZN(n2579) );
  NAND2_X1 U33460 ( .A1(n2585), .A2(REG0_REG_2__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U33470 ( .A1(n2586), .A2(REG1_REG_2__SCAN_IN), .ZN(n2582) );
  NAND2_X1 U33480 ( .A1(n2142), .A2(REG2_REG_2__SCAN_IN), .ZN(n2581) );
  NAND2_X1 U33490 ( .A1(n2781), .A2(REG3_REG_2__SCAN_IN), .ZN(n2580) );
  NAND2_X1 U33500 ( .A1(n3294), .A2(n3314), .ZN(n4183) );
  NAND2_X1 U33510 ( .A1(n3294), .A2(n2458), .ZN(n2584) );
  INV_X1 U33520 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3266) );
  NAND2_X1 U3353 ( .A1(n2781), .A2(n3266), .ZN(n2590) );
  NAND2_X1 U33540 ( .A1(n2585), .A2(REG0_REG_3__SCAN_IN), .ZN(n2589) );
  NAND2_X1 U3355 ( .A1(n2586), .A2(REG1_REG_3__SCAN_IN), .ZN(n2588) );
  NAND2_X1 U3356 ( .A1(n2142), .A2(REG2_REG_3__SCAN_IN), .ZN(n2587) );
  NAND4_X1 U3357 ( .A1(n2590), .A2(n2589), .A3(n2588), .A4(n2587), .ZN(n3336)
         );
  NAND2_X1 U3358 ( .A1(n3336), .A2(n3368), .ZN(n2591) );
  INV_X1 U3359 ( .A(n3368), .ZN(n2896) );
  NAND2_X1 U3360 ( .A1(n4136), .A2(n2896), .ZN(n2592) );
  NAND2_X1 U3361 ( .A1(n2586), .A2(REG1_REG_4__SCAN_IN), .ZN(n2598) );
  NAND2_X1 U3362 ( .A1(n2585), .A2(REG0_REG_4__SCAN_IN), .ZN(n2597) );
  INV_X1 U3363 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2593) );
  NAND2_X1 U3364 ( .A1(n3266), .A2(n2593), .ZN(n2594) );
  AND2_X1 U3365 ( .A1(n2594), .A2(n2600), .ZN(n3720) );
  NAND2_X1 U3366 ( .A1(n2781), .A2(n3720), .ZN(n2596) );
  NAND2_X1 U3367 ( .A1(n3215), .A2(REG2_REG_4__SCAN_IN), .ZN(n2595) );
  NAND2_X1 U3368 ( .A1(n3420), .A2(n2606), .ZN(n4189) );
  NAND2_X1 U3369 ( .A1(n2585), .A2(REG0_REG_5__SCAN_IN), .ZN(n2605) );
  NAND2_X1 U3370 ( .A1(n2586), .A2(REG1_REG_5__SCAN_IN), .ZN(n2604) );
  INV_X1 U3371 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2599) );
  NAND2_X1 U3372 ( .A1(n2600), .A2(n2599), .ZN(n2601) );
  AND2_X1 U3373 ( .A1(n2617), .A2(n2601), .ZN(n3426) );
  NAND2_X1 U3374 ( .A1(n2781), .A2(n3426), .ZN(n2603) );
  NAND2_X1 U3375 ( .A1(n3215), .A2(REG2_REG_5__SCAN_IN), .ZN(n2602) );
  AND2_X1 U3376 ( .A1(n3716), .A2(n3255), .ZN(n2607) );
  NAND2_X1 U3377 ( .A1(n4346), .A2(n2606), .ZN(n3415) );
  NAND2_X1 U3378 ( .A1(n2609), .A2(n2608), .ZN(n3328) );
  NAND2_X1 U3379 ( .A1(n2586), .A2(REG1_REG_7__SCAN_IN), .ZN(n2616) );
  NAND2_X1 U3380 ( .A1(n2585), .A2(REG0_REG_7__SCAN_IN), .ZN(n2615) );
  INV_X1 U3381 ( .A(n2610), .ZN(n2619) );
  INV_X1 U3382 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2611) );
  NAND2_X1 U3383 ( .A1(n2619), .A2(n2611), .ZN(n2612) );
  AND2_X1 U3384 ( .A1(n2634), .A2(n2612), .ZN(n3757) );
  NAND2_X1 U3385 ( .A1(n2781), .A2(n3757), .ZN(n2614) );
  NAND2_X1 U3386 ( .A1(n3215), .A2(REG2_REG_7__SCAN_IN), .ZN(n2613) );
  NAND2_X1 U3387 ( .A1(n3353), .A2(n2626), .ZN(n4194) );
  NAND2_X1 U3388 ( .A1(n3397), .A2(n3754), .ZN(n4197) );
  NAND2_X1 U3389 ( .A1(n4194), .A2(n4197), .ZN(n4286) );
  NAND2_X1 U3390 ( .A1(n2586), .A2(REG1_REG_6__SCAN_IN), .ZN(n2623) );
  NAND2_X1 U3391 ( .A1(n2585), .A2(REG0_REG_6__SCAN_IN), .ZN(n2622) );
  NAND2_X1 U3392 ( .A1(n2617), .A2(n2534), .ZN(n2618) );
  AND2_X1 U3393 ( .A1(n2619), .A2(n2618), .ZN(n3511) );
  NAND2_X1 U3394 ( .A1(n2781), .A2(n3511), .ZN(n2621) );
  NAND2_X1 U3395 ( .A1(n3215), .A2(REG2_REG_6__SCAN_IN), .ZN(n2620) );
  NAND4_X1 U3396 ( .A1(n2623), .A2(n2622), .A3(n2621), .A4(n2620), .ZN(n3753)
         );
  AND2_X1 U3397 ( .A1(n3753), .A2(n3332), .ZN(n2627) );
  AOI22_X1 U3398 ( .A1(n4286), .A2(n2627), .B1(n2626), .B2(n3397), .ZN(n3392)
         );
  NAND2_X1 U3399 ( .A1(n2586), .A2(REG1_REG_9__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U3400 ( .A1(n2585), .A2(REG0_REG_9__SCAN_IN), .ZN(n2632) );
  INV_X1 U3401 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2628) );
  NAND2_X1 U3402 ( .A1(n2636), .A2(n2628), .ZN(n2629) );
  AND2_X1 U3403 ( .A1(n2651), .A2(n2629), .ZN(n3478) );
  NAND2_X1 U3404 ( .A1(n2781), .A2(n3478), .ZN(n2631) );
  NAND2_X1 U3405 ( .A1(n3215), .A2(REG2_REG_9__SCAN_IN), .ZN(n2630) );
  NAND4_X1 U3406 ( .A1(n2633), .A2(n2632), .A3(n2631), .A4(n2630), .ZN(n4343)
         );
  NAND2_X1 U3407 ( .A1(n3447), .A2(n3466), .ZN(n2645) );
  INV_X1 U3408 ( .A(n2645), .ZN(n2642) );
  NAND2_X1 U3409 ( .A1(n2585), .A2(REG0_REG_8__SCAN_IN), .ZN(n2640) );
  NAND2_X1 U3410 ( .A1(n2586), .A2(REG1_REG_8__SCAN_IN), .ZN(n2639) );
  INV_X1 U3411 ( .A(REG3_REG_8__SCAN_IN), .ZN(n3988) );
  NAND2_X1 U3412 ( .A1(n2634), .A2(n3988), .ZN(n2635) );
  AND2_X1 U3413 ( .A1(n2636), .A2(n2635), .ZN(n3536) );
  NAND2_X1 U3414 ( .A1(n2781), .A2(n3536), .ZN(n2638) );
  NAND2_X1 U3415 ( .A1(n3215), .A2(REG2_REG_8__SCAN_IN), .ZN(n2637) );
  INV_X1 U3416 ( .A(n3395), .ZN(n3404) );
  NAND2_X1 U3417 ( .A1(n4344), .A2(n3404), .ZN(n3462) );
  AND2_X1 U3418 ( .A1(n2162), .A2(n3462), .ZN(n2641) );
  AND2_X1 U3419 ( .A1(n3392), .A2(n2644), .ZN(n2643) );
  NAND2_X1 U3420 ( .A1(n3393), .A2(n2643), .ZN(n2649) );
  INV_X1 U3421 ( .A(n2644), .ZN(n2647) );
  NAND2_X1 U3422 ( .A1(n3495), .A2(n3395), .ZN(n3460) );
  AND2_X1 U3423 ( .A1(n3460), .A2(n2645), .ZN(n2646) );
  NAND2_X1 U3424 ( .A1(n2585), .A2(REG0_REG_10__SCAN_IN), .ZN(n2656) );
  NAND2_X1 U3425 ( .A1(n2586), .A2(REG1_REG_10__SCAN_IN), .ZN(n2655) );
  NAND2_X1 U3426 ( .A1(n2651), .A2(n2650), .ZN(n2652) );
  AND2_X1 U3427 ( .A1(n2659), .A2(n2652), .ZN(n3528) );
  NAND2_X1 U3428 ( .A1(n2781), .A2(n3528), .ZN(n2654) );
  NAND2_X1 U3429 ( .A1(n3215), .A2(REG2_REG_10__SCAN_IN), .ZN(n2653) );
  NAND4_X1 U3430 ( .A1(n2656), .A2(n2655), .A3(n2654), .A4(n2653), .ZN(n3222)
         );
  NOR2_X1 U3431 ( .A1(n3222), .A2(n3525), .ZN(n2657) );
  NAND2_X1 U3432 ( .A1(n2585), .A2(REG0_REG_11__SCAN_IN), .ZN(n2664) );
  NAND2_X1 U3433 ( .A1(n2586), .A2(REG1_REG_11__SCAN_IN), .ZN(n2663) );
  INV_X1 U3434 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2658) );
  NAND2_X1 U3435 ( .A1(n2659), .A2(n2658), .ZN(n2660) );
  AND2_X1 U3436 ( .A1(n2666), .A2(n2660), .ZN(n3579) );
  NAND2_X1 U3437 ( .A1(n2781), .A2(n3579), .ZN(n2662) );
  NAND2_X1 U3438 ( .A1(n3215), .A2(REG2_REG_11__SCAN_IN), .ZN(n2661) );
  NAND2_X1 U3439 ( .A1(n3727), .A2(n2665), .ZN(n3584) );
  INV_X1 U3440 ( .A(n3727), .ZN(n4342) );
  NAND2_X1 U3441 ( .A1(n2586), .A2(REG1_REG_12__SCAN_IN), .ZN(n2671) );
  NAND2_X1 U3442 ( .A1(n2585), .A2(REG0_REG_12__SCAN_IN), .ZN(n2670) );
  INV_X1 U3443 ( .A(REG3_REG_12__SCAN_IN), .ZN(n3854) );
  NAND2_X1 U3444 ( .A1(n2666), .A2(n3854), .ZN(n2667) );
  AND2_X1 U3445 ( .A1(n2675), .A2(n2667), .ZN(n3733) );
  NAND2_X1 U3446 ( .A1(n2781), .A2(n3733), .ZN(n2669) );
  NAND2_X1 U3447 ( .A1(n3215), .A2(REG2_REG_12__SCAN_IN), .ZN(n2668) );
  NAND4_X1 U3448 ( .A1(n2671), .A2(n2670), .A3(n2669), .A4(n2668), .ZN(n3624)
         );
  AND2_X1 U3449 ( .A1(n3624), .A2(n3590), .ZN(n2672) );
  OR2_X1 U3450 ( .A1(n2672), .A2(n3595), .ZN(n2674) );
  INV_X1 U3451 ( .A(n3624), .ZN(n4648) );
  NAND2_X1 U3452 ( .A1(n4648), .A2(n3730), .ZN(n2673) );
  NAND2_X1 U3453 ( .A1(n2675), .A2(n3853), .ZN(n2676) );
  NAND2_X1 U3454 ( .A1(n2680), .A2(n2676), .ZN(n4666) );
  INV_X1 U3455 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4667) );
  OAI22_X1 U3456 ( .A1(n4666), .A2(n2771), .B1(n2784), .B2(n4667), .ZN(n2678)
         );
  INV_X1 U3457 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4736) );
  INV_X1 U34580 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4785) );
  OAI22_X1 U34590 ( .A1(n2748), .A2(n4736), .B1(n2285), .B2(n4785), .ZN(n2677)
         );
  NOR2_X1 U3460 ( .A1(n3589), .A2(n4662), .ZN(n3608) );
  NAND2_X1 U3461 ( .A1(n2680), .A2(n2679), .ZN(n2681) );
  NAND2_X1 U3462 ( .A1(n2685), .A2(n2681), .ZN(n3617) );
  AOI22_X1 U3463 ( .A1(n2585), .A2(REG0_REG_14__SCAN_IN), .B1(n2586), .B2(
        REG1_REG_14__SCAN_IN), .ZN(n2683) );
  NAND2_X1 U3464 ( .A1(n3215), .A2(REG2_REG_14__SCAN_IN), .ZN(n2682) );
  OR2_X1 U3465 ( .A1(n4659), .A2(n3615), .ZN(n2692) );
  INV_X1 U3466 ( .A(n2692), .ZN(n2684) );
  NAND2_X1 U34670 ( .A1(n2685), .A2(n2246), .ZN(n2686) );
  NAND2_X1 U3468 ( .A1(n2703), .A2(n2686), .ZN(n4168) );
  OR2_X1 U34690 ( .A1(n4168), .A2(n2771), .ZN(n2691) );
  INV_X1 U3470 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4400) );
  NAND2_X1 U34710 ( .A1(n3215), .A2(REG2_REG_15__SCAN_IN), .ZN(n2688) );
  NAND2_X1 U3472 ( .A1(n2585), .A2(REG0_REG_15__SCAN_IN), .ZN(n2687) );
  OAI211_X1 U34730 ( .C1(n2748), .C2(n4400), .A(n2688), .B(n2687), .ZN(n2689)
         );
  INV_X1 U3474 ( .A(n2689), .ZN(n2690) );
  NAND2_X1 U34750 ( .A1(n3694), .A2(n4172), .ZN(n2693) );
  OR2_X1 U3476 ( .A1(n4659), .A2(n3684), .ZN(n4215) );
  NAND2_X1 U34770 ( .A1(n4659), .A2(n3684), .ZN(n4208) );
  NAND2_X1 U3478 ( .A1(n4215), .A2(n4208), .ZN(n3613) );
  INV_X1 U34790 ( .A(n3613), .ZN(n4274) );
  AND2_X1 U3480 ( .A1(n3589), .A2(n4662), .ZN(n3609) );
  OR2_X1 U34810 ( .A1(n4274), .A2(n3609), .ZN(n3610) );
  AND2_X1 U3482 ( .A1(n2693), .A2(n2430), .ZN(n2694) );
  INV_X1 U34830 ( .A(n4172), .ZN(n3650) );
  XNOR2_X1 U3484 ( .A(n2703), .B(REG3_REG_16__SCAN_IN), .ZN(n3809) );
  NAND2_X1 U34850 ( .A1(n3809), .A2(n2781), .ZN(n2699) );
  INV_X1 U3486 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4870) );
  NAND2_X1 U34870 ( .A1(n3215), .A2(REG2_REG_16__SCAN_IN), .ZN(n2696) );
  NAND2_X1 U3488 ( .A1(n2585), .A2(REG0_REG_16__SCAN_IN), .ZN(n2695) );
  OAI211_X1 U34890 ( .C1(n2748), .C2(n4870), .A(n2696), .B(n2695), .ZN(n2697)
         );
  INV_X1 U3490 ( .A(n2697), .ZN(n2698) );
  OR2_X1 U34910 ( .A1(n4629), .A2(n3806), .ZN(n4302) );
  NAND2_X1 U3492 ( .A1(n4629), .A2(n3806), .ZN(n4298) );
  INV_X1 U34930 ( .A(n3806), .ZN(n3700) );
  NAND2_X1 U3494 ( .A1(n4629), .A2(n3700), .ZN(n2701) );
  OAI21_X1 U34950 ( .B1(n2703), .B2(n2702), .A(n3821), .ZN(n2704) );
  NAND2_X1 U3496 ( .A1(n2704), .A2(n2712), .ZN(n4634) );
  OR2_X1 U34970 ( .A1(n4634), .A2(n2771), .ZN(n2709) );
  INV_X1 U3498 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4635) );
  NAND2_X1 U34990 ( .A1(n2585), .A2(REG0_REG_17__SCAN_IN), .ZN(n2706) );
  NAND2_X1 U3500 ( .A1(n2586), .A2(REG1_REG_17__SCAN_IN), .ZN(n2705) );
  OAI211_X1 U35010 ( .C1(n4635), .C2(n2784), .A(n2706), .B(n2705), .ZN(n2707)
         );
  INV_X1 U3502 ( .A(n2707), .ZN(n2708) );
  NAND2_X1 U35030 ( .A1(n4605), .A2(n4632), .ZN(n2711) );
  AND2_X1 U3504 ( .A1(n4341), .A2(n3823), .ZN(n2710) );
  NAND2_X1 U35050 ( .A1(n2712), .A2(n2236), .ZN(n2713) );
  NAND2_X1 U35060 ( .A1(n2720), .A2(n2713), .ZN(n4620) );
  OR2_X1 U35070 ( .A1(n4620), .A2(n2771), .ZN(n2718) );
  INV_X1 U35080 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4806) );
  NAND2_X1 U35090 ( .A1(n2585), .A2(REG0_REG_18__SCAN_IN), .ZN(n2715) );
  NAND2_X1 U35100 ( .A1(n3215), .A2(REG2_REG_18__SCAN_IN), .ZN(n2714) );
  OAI211_X1 U35110 ( .C1(n2748), .C2(n4806), .A(n2715), .B(n2714), .ZN(n2716)
         );
  INV_X1 U35120 ( .A(n2716), .ZN(n2717) );
  NAND2_X1 U35130 ( .A1(n4624), .A2(n4149), .ZN(n4587) );
  INV_X1 U35140 ( .A(n4149), .ZN(n4616) );
  NAND2_X1 U35150 ( .A1(n3820), .A2(n4616), .ZN(n4588) );
  NAND2_X1 U35160 ( .A1(n4587), .A2(n4588), .ZN(n4612) );
  NAND2_X1 U35170 ( .A1(n4624), .A2(n4616), .ZN(n2719) );
  NAND2_X1 U35180 ( .A1(n2720), .A2(n4046), .ZN(n2721) );
  AND2_X1 U35190 ( .A1(n2148), .A2(n2721), .ZN(n4598) );
  NAND2_X1 U35200 ( .A1(n4598), .A2(n2781), .ZN(n2726) );
  INV_X1 U35210 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4087) );
  NAND2_X1 U35220 ( .A1(n2585), .A2(REG0_REG_19__SCAN_IN), .ZN(n2723) );
  NAND2_X1 U35230 ( .A1(n2586), .A2(REG1_REG_19__SCAN_IN), .ZN(n2722) );
  OAI211_X1 U35240 ( .C1(n4087), .C2(n2784), .A(n2723), .B(n2722), .ZN(n2724)
         );
  INV_X1 U35250 ( .A(n2724), .ZN(n2725) );
  NOR2_X1 U35260 ( .A1(n4610), .A2(n3009), .ZN(n4270) );
  INV_X1 U35270 ( .A(n4270), .ZN(n2727) );
  NAND2_X1 U35280 ( .A1(n4610), .A2(n3009), .ZN(n4269) );
  NAND2_X1 U35290 ( .A1(n2148), .A2(n2237), .ZN(n2729) );
  NAND2_X1 U35300 ( .A1(n2735), .A2(n2729), .ZN(n4579) );
  INV_X1 U35310 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4578) );
  NAND2_X1 U35320 ( .A1(n2586), .A2(REG1_REG_20__SCAN_IN), .ZN(n2731) );
  NAND2_X1 U35330 ( .A1(n2585), .A2(REG0_REG_20__SCAN_IN), .ZN(n2730) );
  OAI211_X1 U35340 ( .C1(n4578), .C2(n2784), .A(n2731), .B(n2730), .ZN(n2732)
         );
  INV_X1 U35350 ( .A(n2732), .ZN(n2733) );
  INV_X1 U35360 ( .A(n3843), .ZN(n4577) );
  NAND2_X1 U35370 ( .A1(n4550), .A2(n3843), .ZN(n4267) );
  NAND2_X1 U35380 ( .A1(n2735), .A2(n4077), .ZN(n2736) );
  NAND2_X1 U35390 ( .A1(n2737), .A2(n2736), .ZN(n4559) );
  INV_X1 U35400 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4768) );
  NAND2_X1 U35410 ( .A1(n2586), .A2(REG1_REG_21__SCAN_IN), .ZN(n2739) );
  NAND2_X1 U35420 ( .A1(n3215), .A2(REG2_REG_21__SCAN_IN), .ZN(n2738) );
  OAI211_X1 U35430 ( .C1(n2285), .C2(n4768), .A(n2739), .B(n2738), .ZN(n2740)
         );
  INV_X1 U35440 ( .A(n2740), .ZN(n2741) );
  NAND2_X1 U35450 ( .A1(n4534), .A2(n2810), .ZN(n2743) );
  XNOR2_X1 U35460 ( .A(n4552), .B(n3030), .ZN(n4532) );
  NAND2_X1 U35470 ( .A1(n2744), .A2(n3773), .ZN(n2745) );
  AND2_X1 U35480 ( .A1(n2753), .A2(n2745), .ZN(n4525) );
  NAND2_X1 U35490 ( .A1(n4525), .A2(n2781), .ZN(n2751) );
  INV_X1 U35500 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4698) );
  NAND2_X1 U35510 ( .A1(n2585), .A2(REG0_REG_23__SCAN_IN), .ZN(n2747) );
  NAND2_X1 U35520 ( .A1(n3215), .A2(REG2_REG_23__SCAN_IN), .ZN(n2746) );
  OAI211_X1 U35530 ( .C1(n2748), .C2(n4698), .A(n2747), .B(n2746), .ZN(n2749)
         );
  INV_X1 U35540 ( .A(n2749), .ZN(n2750) );
  NAND2_X1 U35550 ( .A1(n2753), .A2(n2241), .ZN(n2754) );
  NAND2_X1 U35560 ( .A1(n2761), .A2(n2754), .ZN(n4504) );
  INV_X1 U35570 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4503) );
  NAND2_X1 U35580 ( .A1(n2586), .A2(REG1_REG_24__SCAN_IN), .ZN(n2756) );
  NAND2_X1 U35590 ( .A1(n2585), .A2(REG0_REG_24__SCAN_IN), .ZN(n2755) );
  OAI211_X1 U35600 ( .C1(n4503), .C2(n2784), .A(n2756), .B(n2755), .ZN(n2757)
         );
  INV_X1 U35610 ( .A(n2757), .ZN(n2758) );
  NAND2_X1 U35620 ( .A1(n4518), .A2(n3831), .ZN(n2760) );
  NAND2_X1 U35630 ( .A1(n2761), .A2(n4090), .ZN(n2762) );
  NAND2_X1 U35640 ( .A1(n4489), .A2(n2781), .ZN(n2767) );
  INV_X1 U35650 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4755) );
  NAND2_X1 U35660 ( .A1(n3215), .A2(REG2_REG_25__SCAN_IN), .ZN(n2764) );
  NAND2_X1 U35670 ( .A1(n2586), .A2(REG1_REG_25__SCAN_IN), .ZN(n2763) );
  OAI211_X1 U35680 ( .C1(n2285), .C2(n4755), .A(n2764), .B(n2763), .ZN(n2765)
         );
  INV_X1 U35690 ( .A(n2765), .ZN(n2766) );
  NAND2_X1 U35700 ( .A1(n4461), .A2(n4487), .ZN(n2769) );
  NOR2_X1 U35710 ( .A1(n4461), .A2(n4487), .ZN(n2768) );
  NAND2_X1 U35720 ( .A1(n2143), .A2(n2242), .ZN(n2770) );
  NAND2_X1 U35730 ( .A1(n2778), .A2(n2770), .ZN(n4470) );
  INV_X1 U35740 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4469) );
  NAND2_X1 U35750 ( .A1(n2585), .A2(REG0_REG_26__SCAN_IN), .ZN(n2773) );
  NAND2_X1 U35760 ( .A1(n2586), .A2(REG1_REG_26__SCAN_IN), .ZN(n2772) );
  OAI211_X1 U35770 ( .C1(n4469), .C2(n2784), .A(n2773), .B(n2772), .ZN(n2774)
         );
  INV_X1 U35780 ( .A(n2774), .ZN(n2775) );
  NAND2_X1 U35790 ( .A1(n2778), .A2(n4072), .ZN(n2779) );
  NAND2_X1 U35800 ( .A1(n4448), .A2(n2781), .ZN(n2787) );
  INV_X1 U35810 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4449) );
  NAND2_X1 U3582 ( .A1(n2585), .A2(REG0_REG_27__SCAN_IN), .ZN(n2783) );
  NAND2_X1 U3583 ( .A1(n2586), .A2(REG1_REG_27__SCAN_IN), .ZN(n2782) );
  OAI211_X1 U3584 ( .C1(n4449), .C2(n2784), .A(n2783), .B(n2782), .ZN(n2785)
         );
  INV_X1 U3585 ( .A(n2785), .ZN(n2786) );
  NAND2_X1 U3586 ( .A1(n3062), .A2(n3091), .ZN(n4236) );
  INV_X1 U3587 ( .A(n3091), .ZN(n3111) );
  NAND2_X1 U3588 ( .A1(n4444), .A2(n3111), .ZN(n4230) );
  NAND2_X1 U3589 ( .A1(n4236), .A2(n4230), .ZN(n4248) );
  NAND2_X1 U3590 ( .A1(n3102), .A2(n4248), .ZN(n4427) );
  INV_X1 U3591 ( .A(n4427), .ZN(n2789) );
  NAND3_X1 U3592 ( .A1(n2789), .A2(n4429), .A3(n4975), .ZN(n2835) );
  INV_X1 U3593 ( .A(n4429), .ZN(n2790) );
  NAND4_X1 U3594 ( .A1(n4427), .A2(n4975), .A3(n2790), .A4(n4426), .ZN(n2834)
         );
  NAND2_X1 U3595 ( .A1(n2880), .A2(n3747), .ZN(n4257) );
  NAND2_X1 U3596 ( .A1(n3309), .A2(n4276), .ZN(n3308) );
  NAND2_X1 U3597 ( .A1(n3308), .A2(n4183), .ZN(n3361) );
  NAND2_X1 U3598 ( .A1(n4136), .A2(n3368), .ZN(n4188) );
  NAND2_X1 U3599 ( .A1(n3336), .A2(n2896), .ZN(n4185) );
  NAND2_X1 U3600 ( .A1(n3361), .A2(n4271), .ZN(n2791) );
  INV_X1 U3601 ( .A(n4189), .ZN(n2792) );
  NAND2_X1 U3602 ( .A1(n3716), .A2(n3425), .ZN(n4204) );
  INV_X1 U3603 ( .A(n3332), .ZN(n3502) );
  NAND2_X1 U3604 ( .A1(n3753), .A2(n3502), .ZN(n4202) );
  INV_X1 U3605 ( .A(n3753), .ZN(n2794) );
  NAND2_X1 U3606 ( .A1(n2794), .A2(n3332), .ZN(n4193) );
  INV_X1 U3607 ( .A(n4194), .ZN(n2795) );
  NAND2_X1 U3608 ( .A1(n2796), .A2(n4197), .ZN(n3394) );
  NAND2_X1 U3609 ( .A1(n3495), .A2(n3404), .ZN(n4198) );
  NAND2_X1 U3610 ( .A1(n3394), .A2(n4198), .ZN(n2797) );
  NAND2_X1 U3611 ( .A1(n4344), .A2(n3395), .ZN(n4196) );
  NAND2_X1 U3612 ( .A1(n2797), .A2(n4196), .ZN(n3465) );
  AND2_X1 U3613 ( .A1(n4343), .A2(n3466), .ZN(n4203) );
  NAND2_X1 U3614 ( .A1(n3447), .A2(n3470), .ZN(n4199) );
  NAND2_X1 U3615 ( .A1(n3222), .A2(n3449), .ZN(n4212) );
  NAND2_X1 U3616 ( .A1(n3569), .A2(n3525), .ZN(n4207) );
  INV_X1 U3617 ( .A(n4662), .ZN(n4646) );
  NAND2_X1 U3618 ( .A1(n3589), .A2(n4646), .ZN(n4253) );
  NAND2_X1 U3619 ( .A1(n3624), .A2(n3730), .ZN(n4649) );
  NAND2_X1 U3620 ( .A1(n4253), .A2(n4649), .ZN(n2799) );
  INV_X1 U3621 ( .A(n3587), .ZN(n2798) );
  INV_X1 U3622 ( .A(n2799), .ZN(n2801) );
  NAND2_X1 U3623 ( .A1(n4648), .A2(n3590), .ZN(n4651) );
  NAND2_X1 U3624 ( .A1(n3584), .A2(n4651), .ZN(n2800) );
  NAND2_X1 U3625 ( .A1(n2801), .A2(n2800), .ZN(n2802) );
  INV_X1 U3626 ( .A(n3589), .ZN(n3728) );
  NAND2_X1 U3627 ( .A1(n3728), .A2(n4662), .ZN(n4254) );
  AND2_X1 U3628 ( .A1(n2802), .A2(n4254), .ZN(n4219) );
  NAND2_X1 U3629 ( .A1(n2803), .A2(n4219), .ZN(n3604) );
  NAND2_X1 U3630 ( .A1(n3604), .A2(n4274), .ZN(n2804) );
  NAND2_X1 U3631 ( .A1(n3805), .A2(n4172), .ZN(n4216) );
  NAND2_X1 U3632 ( .A1(n3694), .A2(n3650), .ZN(n4209) );
  NAND2_X1 U3633 ( .A1(n3692), .A2(n4298), .ZN(n4625) );
  NAND2_X1 U3634 ( .A1(n4610), .A2(n4597), .ZN(n2805) );
  NAND2_X1 U3635 ( .A1(n2805), .A2(n4588), .ZN(n2807) );
  AND2_X1 U3636 ( .A1(n4341), .A2(n4632), .ZN(n4586) );
  OR2_X1 U3637 ( .A1(n2807), .A2(n4586), .ZN(n4301) );
  NOR2_X1 U3638 ( .A1(n4625), .A2(n4301), .ZN(n4565) );
  NAND2_X1 U3639 ( .A1(n4593), .A2(n3843), .ZN(n4299) );
  NAND2_X1 U3640 ( .A1(n4605), .A2(n3823), .ZN(n4585) );
  AND2_X1 U3641 ( .A1(n4587), .A2(n4585), .ZN(n2806) );
  OAI22_X1 U3642 ( .A1(n2807), .A2(n2806), .B1(n4610), .B2(n4597), .ZN(n4564)
         );
  NOR2_X1 U3643 ( .A1(n4593), .A2(n3843), .ZN(n2808) );
  OR2_X1 U3644 ( .A1(n4564), .A2(n2808), .ZN(n2809) );
  AOI21_X1 U3645 ( .B1(n4565), .B2(n4299), .A(n4304), .ZN(n4548) );
  NAND2_X1 U3646 ( .A1(n4516), .A2(n4542), .ZN(n4513) );
  NAND2_X1 U3647 ( .A1(n4570), .A2(n2810), .ZN(n4511) );
  AND2_X1 U3648 ( .A1(n4513), .A2(n4511), .ZN(n4306) );
  NAND2_X1 U3649 ( .A1(n4548), .A2(n4306), .ZN(n2812) );
  AND2_X1 U3650 ( .A1(n4534), .A2(n4557), .ZN(n4510) );
  NAND2_X1 U3651 ( .A1(n4340), .A2(n4523), .ZN(n4250) );
  NAND2_X1 U3652 ( .A1(n4552), .A2(n3030), .ZN(n2811) );
  NAND2_X1 U3653 ( .A1(n4250), .A2(n2811), .ZN(n4225) );
  AOI21_X1 U3654 ( .B1(n4510), .B2(n4513), .A(n4225), .ZN(n4307) );
  NOR2_X1 U3655 ( .A1(n4340), .A2(n4523), .ZN(n4252) );
  NAND2_X1 U3656 ( .A1(n4480), .A2(n3831), .ZN(n4249) );
  NAND2_X1 U3657 ( .A1(n4437), .A2(n4155), .ZN(n2813) );
  NAND2_X1 U3658 ( .A1(n4461), .A2(n3047), .ZN(n4456) );
  NAND2_X1 U3659 ( .A1(n4498), .A2(n4487), .ZN(n4258) );
  NAND2_X1 U3660 ( .A1(n4518), .A2(n4502), .ZN(n4476) );
  NAND2_X1 U3661 ( .A1(n4258), .A2(n4476), .ZN(n4457) );
  AND2_X1 U3662 ( .A1(n4482), .A2(n4467), .ZN(n4316) );
  AOI21_X1 U3663 ( .B1(n2814), .B2(n4457), .A(n4316), .ZN(n4233) );
  NAND2_X1 U3664 ( .A1(n3057), .A2(n2815), .ZN(n4235) );
  NAND2_X1 U3665 ( .A1(n4463), .A2(n4447), .ZN(n4232) );
  NAND2_X1 U3666 ( .A1(n4235), .A2(n4232), .ZN(n4445) );
  INV_X1 U3667 ( .A(n4235), .ZN(n2816) );
  INV_X1 U3668 ( .A(n4230), .ZN(n2817) );
  OAI21_X1 U3669 ( .B1(n3103), .B2(n2817), .A(n4236), .ZN(n2818) );
  XNOR2_X1 U3670 ( .A(n2818), .B(n4429), .ZN(n2833) );
  INV_X1 U3671 ( .A(n2855), .ZN(n4793) );
  NAND2_X1 U3672 ( .A1(n4793), .A2(n4327), .ZN(n2820) );
  NAND2_X1 U3673 ( .A1(n4792), .A2(n4802), .ZN(n2819) );
  INV_X1 U3674 ( .A(n2850), .ZN(n2822) );
  NOR2_X1 U3675 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .ZN(n2821)
         );
  AOI21_X1 U3676 ( .B1(n2822), .B2(n2821), .A(n2455), .ZN(n2823) );
  MUX2_X1 U3677 ( .A(n2455), .B(n2823), .S(IR_REG_28__SCAN_IN), .Z(n2825) );
  OR2_X1 U3678 ( .A1(n2825), .A2(n2824), .ZN(n3175) );
  NAND2_X1 U3679 ( .A1(n4790), .A2(n3152), .ZN(n4647) );
  NAND2_X1 U3680 ( .A1(n2586), .A2(REG1_REG_30__SCAN_IN), .ZN(n2828) );
  NAND2_X1 U3681 ( .A1(n3215), .A2(REG2_REG_30__SCAN_IN), .ZN(n2827) );
  NAND2_X1 U3682 ( .A1(n2585), .A2(REG0_REG_30__SCAN_IN), .ZN(n2826) );
  NAND3_X1 U3683 ( .A1(n2828), .A2(n2827), .A3(n2826), .ZN(n4339) );
  OAI21_X1 U3684 ( .B1(n2850), .B2(IR_REG_26__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2829) );
  XNOR2_X1 U3685 ( .A(n2829), .B(IR_REG_27__SCAN_IN), .ZN(n3167) );
  NAND2_X1 U3686 ( .A1(n3167), .A2(B_REG_SCAN_IN), .ZN(n2830) );
  AND2_X1 U3687 ( .A1(n4660), .A2(n2830), .ZN(n4411) );
  NAND2_X1 U3688 ( .A1(n4901), .A2(n4793), .ZN(n4645) );
  AOI22_X1 U3689 ( .A1(n4339), .A2(n4411), .B1(n4568), .B2(n4237), .ZN(n2831)
         );
  OAI21_X1 U3690 ( .B1(n3062), .B2(n4647), .A(n2831), .ZN(n2832) );
  NAND4_X1 U3691 ( .A1(n2836), .A2(n2835), .A3(n2834), .A4(n4431), .ZN(n2875)
         );
  NAND2_X1 U3692 ( .A1(IR_REG_23__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2838) );
  NAND2_X1 U3693 ( .A1(n2838), .A2(IR_REG_31__SCAN_IN), .ZN(n2839) );
  OAI21_X1 U3694 ( .B1(n2840), .B2(IR_REG_31__SCAN_IN), .A(n2839), .ZN(n2841)
         );
  OAI211_X2 U3695 ( .C1(n2141), .C2(n2843), .A(n2842), .B(n2841), .ZN(n3139)
         );
  NAND2_X2 U3696 ( .A1(n2852), .A2(n4791), .ZN(n2879) );
  NAND2_X1 U3697 ( .A1(n2141), .A2(IR_REG_31__SCAN_IN), .ZN(n2854) );
  NAND2_X1 U3698 ( .A1(n2855), .A2(n4812), .ZN(n3068) );
  NOR2_X1 U3699 ( .A1(n3149), .A2(n3081), .ZN(n3230) );
  NAND2_X1 U3700 ( .A1(n3139), .A2(n3135), .ZN(n2856) );
  MUX2_X1 U3701 ( .A(n3139), .B(n2856), .S(B_REG_SCAN_IN), .Z(n2857) );
  INV_X1 U3702 ( .A(n3141), .ZN(n2868) );
  NOR4_X1 U3703 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_7__SCAN_IN), .ZN(n2858) );
  INV_X1 U3704 ( .A(D_REG_5__SCAN_IN), .ZN(n4927) );
  INV_X1 U3705 ( .A(D_REG_26__SCAN_IN), .ZN(n4918) );
  NAND3_X1 U3706 ( .A1(n2858), .A2(n4927), .A3(n4918), .ZN(n2864) );
  NOR4_X1 U3707 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2862) );
  NOR4_X1 U3708 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2861) );
  NOR4_X1 U3709 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2860) );
  NOR4_X1 U3710 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n2859) );
  NAND4_X1 U3711 ( .A1(n2862), .A2(n2861), .A3(n2860), .A4(n2859), .ZN(n2863)
         );
  NOR4_X1 U3712 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(n2864), 
        .A4(n2863), .ZN(n2866) );
  INV_X1 U3713 ( .A(D_REG_19__SCAN_IN), .ZN(n4922) );
  INV_X1 U3714 ( .A(D_REG_20__SCAN_IN), .ZN(n4921) );
  INV_X1 U3715 ( .A(D_REG_2__SCAN_IN), .ZN(n4929) );
  INV_X1 U3716 ( .A(D_REG_30__SCAN_IN), .ZN(n4917) );
  NAND4_X1 U3717 ( .A1(n4922), .A2(n4921), .A3(n4929), .A4(n4917), .ZN(n2865)
         );
  NOR3_X1 U3718 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(n2865), 
        .ZN(n3874) );
  NAND2_X1 U3719 ( .A1(n2866), .A2(n3874), .ZN(n2867) );
  NAND2_X1 U3720 ( .A1(n2868), .A2(n2867), .ZN(n3066) );
  NAND2_X1 U3721 ( .A1(n3230), .A2(n3066), .ZN(n3280) );
  INV_X1 U3722 ( .A(n4791), .ZN(n2871) );
  NAND2_X1 U3723 ( .A1(n2871), .A2(n3135), .ZN(n3145) );
  OAI21_X1 U3724 ( .B1(n3141), .B2(D_REG_1__SCAN_IN), .A(n3145), .ZN(n3065) );
  NAND2_X1 U3725 ( .A1(n4963), .A2(n2869), .ZN(n3088) );
  NAND2_X1 U3726 ( .A1(n3065), .A2(n3088), .ZN(n2870) );
  NAND2_X1 U3727 ( .A1(n3139), .A2(n2871), .ZN(n3143) );
  NAND2_X1 U3728 ( .A1(n2875), .A2(n4994), .ZN(n2873) );
  NAND2_X1 U3729 ( .A1(n4991), .A2(REG1_REG_29__SCAN_IN), .ZN(n2872) );
  NAND2_X1 U3730 ( .A1(n2873), .A2(n2872), .ZN(U3547) );
  NOR2_X4 U3731 ( .A1(n2874), .A2(n3067), .ZN(n4777) );
  NAND2_X1 U3732 ( .A1(n2875), .A2(n4777), .ZN(n2878) );
  INV_X1 U3733 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2876) );
  NAND2_X1 U3734 ( .A1(n2878), .A2(n2877), .ZN(U3515) );
  INV_X2 U3735 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3736 ( .A(n2879), .ZN(n3119) );
  NAND2_X4 U3737 ( .A1(n2879), .A2(n3300), .ZN(n3058) );
  AOI21_X1 U3738 ( .B1(REG1_REG_0__SCAN_IN), .B2(n3119), .A(n2884), .ZN(n3744)
         );
  OR2_X4 U3739 ( .A1(n3058), .A2(n4972), .ZN(n3061) );
  INV_X1 U3740 ( .A(IR_REG_0__SCAN_IN), .ZN(n4943) );
  OAI22_X1 U3741 ( .A1(n2131), .A2(n4903), .B1(n4943), .B2(n2879), .ZN(n2882)
         );
  AOI21_X2 U3742 ( .B1(n2919), .B2(n2881), .A(n2882), .ZN(n3745) );
  OAI22_X1 U3743 ( .A1(n3744), .A2(n3745), .B1(n3055), .B2(n2884), .ZN(n3229)
         );
  OAI22_X1 U3744 ( .A1(n3294), .A2(n2131), .B1(n3058), .B2(n2458), .ZN(n2891)
         );
  XNOR2_X1 U3745 ( .A(n2891), .B(n3055), .ZN(n2893) );
  OAI22_X1 U3746 ( .A1(n3294), .A2(n3061), .B1(n2131), .B2(n2458), .ZN(n2892)
         );
  NOR2_X1 U3747 ( .A1(n2893), .A2(n2892), .ZN(n2894) );
  AOI21_X1 U3748 ( .B1(n2893), .B2(n2892), .A(n2894), .ZN(n4132) );
  NAND2_X1 U3749 ( .A1(n4131), .A2(n4132), .ZN(n4130) );
  INV_X1 U3750 ( .A(n2894), .ZN(n2895) );
  NAND2_X1 U3751 ( .A1(n4130), .A2(n2895), .ZN(n3262) );
  OAI22_X1 U3752 ( .A1(n4136), .A2(n3061), .B1(n2131), .B2(n2896), .ZN(n2902)
         );
  NAND2_X1 U3753 ( .A1(n3336), .A2(n2962), .ZN(n2898) );
  OR2_X1 U3754 ( .A1(n3058), .A2(n2896), .ZN(n2897) );
  NAND2_X1 U3755 ( .A1(n2898), .A2(n2897), .ZN(n2899) );
  XNOR2_X1 U3756 ( .A(n2899), .B(n3055), .ZN(n2901) );
  XOR2_X1 U3757 ( .A(n2902), .B(n2901), .Z(n3265) );
  NAND2_X1 U3758 ( .A1(n3262), .A2(n3265), .ZN(n3263) );
  OAI22_X1 U3759 ( .A1(n3420), .A2(n3061), .B1(n3717), .B2(n2131), .ZN(n2907)
         );
  INV_X1 U3760 ( .A(n2901), .ZN(n2904) );
  INV_X1 U3761 ( .A(n2902), .ZN(n2903) );
  NAND2_X1 U3762 ( .A1(n2904), .A2(n2903), .ZN(n3715) );
  NAND2_X1 U3763 ( .A1(n3263), .A2(n2905), .ZN(n3713) );
  INV_X1 U3764 ( .A(n2906), .ZN(n2908) );
  OAI22_X1 U3765 ( .A1(n3716), .A2(n2131), .B1(n3255), .B2(n3058), .ZN(n2910)
         );
  XNOR2_X1 U3766 ( .A(n2910), .B(n3059), .ZN(n2911) );
  OAI22_X1 U3767 ( .A1(n3716), .A2(n3061), .B1(n3255), .B2(n2131), .ZN(n2912)
         );
  XNOR2_X1 U3768 ( .A(n2911), .B(n2912), .ZN(n3253) );
  INV_X1 U3769 ( .A(n2911), .ZN(n2913) );
  NAND2_X1 U3770 ( .A1(n2913), .A2(n2912), .ZN(n2914) );
  INV_X1 U3771 ( .A(n2914), .ZN(n2915) );
  INV_X2 U3772 ( .A(n2131), .ZN(n2962) );
  NAND2_X1 U3773 ( .A1(n3753), .A2(n2962), .ZN(n2917) );
  OR2_X1 U3774 ( .A1(n3058), .A2(n3502), .ZN(n2916) );
  NAND2_X1 U3775 ( .A1(n2917), .A2(n2916), .ZN(n2918) );
  XNOR2_X1 U3776 ( .A(n2918), .B(n3059), .ZN(n2924) );
  INV_X1 U3777 ( .A(n2924), .ZN(n2922) );
  NOR2_X1 U3778 ( .A1(n2131), .A2(n3502), .ZN(n2920) );
  AOI21_X1 U3779 ( .B1(n3753), .B2(n2919), .A(n2920), .ZN(n2923) );
  INV_X1 U3780 ( .A(n2923), .ZN(n2921) );
  NAND2_X1 U3781 ( .A1(n2922), .A2(n2921), .ZN(n3272) );
  OAI22_X1 U3782 ( .A1(n3353), .A2(n3061), .B1(n3754), .B2(n2131), .ZN(n2927)
         );
  OAI22_X1 U3783 ( .A1(n3353), .A2(n2131), .B1(n3754), .B2(n3058), .ZN(n2925)
         );
  XNOR2_X1 U3784 ( .A(n2925), .B(n3055), .ZN(n2926) );
  XOR2_X1 U3785 ( .A(n2927), .B(n2926), .Z(n3751) );
  NAND2_X1 U3786 ( .A1(n2926), .A2(n2927), .ZN(n2928) );
  OAI22_X1 U3787 ( .A1(n3495), .A2(n2131), .B1(n3395), .B2(n3058), .ZN(n2929)
         );
  XNOR2_X1 U3788 ( .A(n2929), .B(n3055), .ZN(n2930) );
  OAI22_X1 U3789 ( .A1(n3495), .A2(n3061), .B1(n3395), .B2(n2131), .ZN(n2931)
         );
  AND2_X1 U3790 ( .A1(n2930), .A2(n2931), .ZN(n3349) );
  INV_X1 U3791 ( .A(n2930), .ZN(n2933) );
  INV_X1 U3792 ( .A(n2931), .ZN(n2932) );
  NAND2_X1 U3793 ( .A1(n2933), .A2(n2932), .ZN(n3348) );
  OAI22_X1 U3794 ( .A1(n3447), .A2(n3061), .B1(n2131), .B2(n3466), .ZN(n2938)
         );
  NAND2_X1 U3795 ( .A1(n4343), .A2(n2962), .ZN(n2935) );
  NAND2_X1 U3796 ( .A1(n3010), .A2(n3470), .ZN(n2934) );
  NAND2_X1 U3797 ( .A1(n2935), .A2(n2934), .ZN(n2936) );
  XNOR2_X1 U3798 ( .A(n2936), .B(n3055), .ZN(n2937) );
  XOR2_X1 U3799 ( .A(n2938), .B(n2937), .Z(n3406) );
  INV_X1 U3800 ( .A(n2937), .ZN(n2940) );
  INV_X1 U3801 ( .A(n2938), .ZN(n2939) );
  OAI22_X1 U3802 ( .A1(n3569), .A2(n2131), .B1(n3058), .B2(n3449), .ZN(n2941)
         );
  XNOR2_X1 U3803 ( .A(n2941), .B(n3055), .ZN(n2943) );
  NOR2_X1 U3804 ( .A1(n2131), .A2(n3449), .ZN(n2942) );
  AOI21_X1 U3805 ( .B1(n3222), .B2(n2919), .A(n2942), .ZN(n2944) );
  XNOR2_X1 U3806 ( .A(n2943), .B(n2944), .ZN(n3445) );
  NAND2_X1 U3807 ( .A1(n3446), .A2(n3445), .ZN(n3444) );
  INV_X1 U3808 ( .A(n2948), .ZN(n3485) );
  XNOR2_X1 U3809 ( .A(n2947), .B(n3055), .ZN(n3486) );
  NAND2_X1 U3810 ( .A1(n3624), .A2(n2962), .ZN(n2950) );
  NAND2_X1 U3811 ( .A1(n3590), .A2(n3010), .ZN(n2949) );
  NAND2_X1 U3812 ( .A1(n2950), .A2(n2949), .ZN(n2951) );
  XNOR2_X1 U3813 ( .A(n2951), .B(n3055), .ZN(n2954) );
  NAND2_X1 U3814 ( .A1(n3624), .A2(n2919), .ZN(n2953) );
  NAND2_X1 U3815 ( .A1(n3590), .A2(n2962), .ZN(n2952) );
  NAND2_X1 U3816 ( .A1(n2953), .A2(n2952), .ZN(n2955) );
  INV_X1 U3817 ( .A(n2954), .ZN(n2957) );
  INV_X1 U3818 ( .A(n2955), .ZN(n2956) );
  NAND2_X1 U3819 ( .A1(n3589), .A2(n2962), .ZN(n2959) );
  NAND2_X1 U3820 ( .A1(n3010), .A2(n4662), .ZN(n2958) );
  NAND2_X1 U3821 ( .A1(n2959), .A2(n2958), .ZN(n2960) );
  XNOR2_X1 U3822 ( .A(n2960), .B(n3059), .ZN(n3676) );
  NOR2_X1 U3823 ( .A1(n2131), .A2(n4646), .ZN(n2961) );
  AOI21_X1 U3824 ( .B1(n3589), .B2(n2919), .A(n2961), .ZN(n3675) );
  NAND2_X1 U3825 ( .A1(n4659), .A2(n2962), .ZN(n2964) );
  NAND2_X1 U3826 ( .A1(n3010), .A2(n3615), .ZN(n2963) );
  NAND2_X1 U3827 ( .A1(n2964), .A2(n2963), .ZN(n2965) );
  XNOR2_X1 U3828 ( .A(n2965), .B(n3055), .ZN(n2970) );
  NAND2_X1 U3829 ( .A1(n4659), .A2(n2919), .ZN(n2967) );
  NAND2_X1 U3830 ( .A1(n2962), .A2(n3615), .ZN(n2966) );
  NAND2_X1 U3831 ( .A1(n2967), .A2(n2966), .ZN(n2971) );
  NAND2_X1 U3832 ( .A1(n2970), .A2(n2971), .ZN(n3681) );
  INV_X1 U3833 ( .A(n3681), .ZN(n2975) );
  NAND2_X1 U3834 ( .A1(n3676), .A2(n3675), .ZN(n2974) );
  INV_X1 U3835 ( .A(n2970), .ZN(n2973) );
  INV_X1 U3836 ( .A(n2971), .ZN(n2972) );
  NAND2_X1 U3837 ( .A1(n2973), .A2(n2972), .ZN(n3680) );
  NAND2_X1 U3838 ( .A1(n2978), .A2(n2977), .ZN(n3802) );
  NAND2_X1 U3839 ( .A1(n4629), .A2(n2962), .ZN(n2980) );
  OR2_X1 U3840 ( .A1(n3806), .A2(n3058), .ZN(n2979) );
  NAND2_X1 U3841 ( .A1(n2980), .A2(n2979), .ZN(n2981) );
  XNOR2_X1 U3842 ( .A(n2981), .B(n3059), .ZN(n3815) );
  INV_X1 U3843 ( .A(n3815), .ZN(n2990) );
  NAND2_X1 U3844 ( .A1(n4629), .A2(n2919), .ZN(n2983) );
  OR2_X1 U3845 ( .A1(n3806), .A2(n2131), .ZN(n2982) );
  NAND2_X1 U3846 ( .A1(n2983), .A2(n2982), .ZN(n2995) );
  NAND2_X1 U3847 ( .A1(n3694), .A2(n2919), .ZN(n2985) );
  NAND2_X1 U3848 ( .A1(n2962), .A2(n4172), .ZN(n2984) );
  NAND2_X1 U3849 ( .A1(n2985), .A2(n2984), .ZN(n4164) );
  NAND2_X1 U3850 ( .A1(n3694), .A2(n2962), .ZN(n2988) );
  NAND2_X1 U3851 ( .A1(n3010), .A2(n4172), .ZN(n2987) );
  NAND2_X1 U3852 ( .A1(n2988), .A2(n2987), .ZN(n2989) );
  XNOR2_X1 U3853 ( .A(n2989), .B(n3055), .ZN(n2994) );
  AOI22_X1 U3854 ( .A1(n2990), .A2(n2995), .B1(n4164), .B2(n2994), .ZN(n2991)
         );
  NAND2_X1 U3855 ( .A1(n3802), .A2(n2991), .ZN(n3002) );
  OAI22_X1 U3856 ( .A1(n4605), .A2(n2131), .B1(n3058), .B2(n4632), .ZN(n2992)
         );
  XNOR2_X1 U3857 ( .A(n2992), .B(n3055), .ZN(n3816) );
  OAI22_X1 U3858 ( .A1(n4605), .A2(n3061), .B1(n2131), .B2(n4632), .ZN(n3817)
         );
  OAI21_X1 U3859 ( .B1(n2994), .B2(n4164), .A(n2995), .ZN(n2993) );
  NAND2_X1 U3860 ( .A1(n2993), .A2(n3815), .ZN(n2998) );
  INV_X1 U3861 ( .A(n2994), .ZN(n3803) );
  INV_X1 U3862 ( .A(n2995), .ZN(n3814) );
  INV_X1 U3863 ( .A(n4164), .ZN(n2996) );
  NAND3_X1 U3864 ( .A1(n3803), .A2(n3814), .A3(n2996), .ZN(n2997) );
  OAI211_X1 U3865 ( .C1(n3816), .C2(n3817), .A(n2998), .B(n2997), .ZN(n2999)
         );
  OAI22_X1 U3866 ( .A1(n4624), .A2(n2131), .B1(n3058), .B2(n4616), .ZN(n3003)
         );
  XNOR2_X1 U3867 ( .A(n3003), .B(n3059), .ZN(n3008) );
  INV_X1 U3868 ( .A(n3008), .ZN(n3006) );
  AND2_X1 U3869 ( .A1(n2962), .A2(n4149), .ZN(n3004) );
  AOI21_X1 U3870 ( .B1(n3820), .B2(n2919), .A(n3004), .ZN(n3007) );
  INV_X1 U3871 ( .A(n3007), .ZN(n3005) );
  NAND2_X1 U3872 ( .A1(n3006), .A2(n3005), .ZN(n4145) );
  AND2_X1 U3873 ( .A1(n3008), .A2(n3007), .ZN(n4144) );
  AOI22_X1 U3874 ( .A1(n4610), .A2(n2919), .B1(n2962), .B2(n3009), .ZN(n3014)
         );
  NAND2_X1 U3875 ( .A1(n4610), .A2(n2962), .ZN(n3012) );
  NAND2_X1 U3876 ( .A1(n3010), .A2(n3009), .ZN(n3011) );
  NAND2_X1 U3877 ( .A1(n3012), .A2(n3011), .ZN(n3013) );
  XNOR2_X1 U3878 ( .A(n3013), .B(n3055), .ZN(n3016) );
  XOR2_X1 U3879 ( .A(n3014), .B(n3016), .Z(n3779) );
  INV_X1 U3880 ( .A(n3014), .ZN(n3015) );
  OAI22_X1 U3881 ( .A1(n4550), .A2(n2131), .B1(n3058), .B2(n3843), .ZN(n3017)
         );
  XNOR2_X1 U3882 ( .A(n3017), .B(n3055), .ZN(n3018) );
  OAI22_X1 U3883 ( .A1(n4550), .A2(n3061), .B1(n2131), .B2(n3843), .ZN(n3019)
         );
  NAND2_X1 U3884 ( .A1(n3018), .A2(n3019), .ZN(n3839) );
  INV_X1 U3885 ( .A(n3018), .ZN(n3021) );
  INV_X1 U3886 ( .A(n3019), .ZN(n3020) );
  NAND2_X1 U3887 ( .A1(n3021), .A2(n3020), .ZN(n3841) );
  NAND2_X1 U3888 ( .A1(n4534), .A2(n2962), .ZN(n3023) );
  OR2_X1 U3889 ( .A1(n3058), .A2(n4557), .ZN(n3022) );
  NAND2_X1 U3890 ( .A1(n3023), .A2(n3022), .ZN(n3024) );
  XNOR2_X1 U3891 ( .A(n3024), .B(n3059), .ZN(n3786) );
  NOR2_X1 U3892 ( .A1(n2131), .A2(n4557), .ZN(n3025) );
  AOI21_X1 U3893 ( .B1(n4534), .B2(n2919), .A(n3025), .ZN(n3027) );
  NAND2_X1 U3894 ( .A1(n3786), .A2(n3027), .ZN(n3026) );
  INV_X1 U3895 ( .A(n3786), .ZN(n3028) );
  INV_X1 U3896 ( .A(n3027), .ZN(n3785) );
  OAI22_X1 U3897 ( .A1(n4516), .A2(n2131), .B1(n3058), .B2(n3030), .ZN(n3029)
         );
  XNOR2_X1 U3898 ( .A(n3029), .B(n3055), .ZN(n3035) );
  OAI22_X1 U3899 ( .A1(n4516), .A2(n3061), .B1(n2131), .B2(n3030), .ZN(n3034)
         );
  XNOR2_X1 U3900 ( .A(n3035), .B(n3034), .ZN(n3707) );
  NAND2_X1 U3901 ( .A1(n3032), .A2(n3031), .ZN(n3705) );
  OAI22_X1 U3902 ( .A1(n4536), .A2(n2131), .B1(n4523), .B2(n3058), .ZN(n3033)
         );
  XNOR2_X1 U3903 ( .A(n3033), .B(n3055), .ZN(n3038) );
  OAI22_X1 U3904 ( .A1(n4536), .A2(n3061), .B1(n4523), .B2(n2131), .ZN(n3037)
         );
  XNOR2_X1 U3905 ( .A(n3038), .B(n3037), .ZN(n3768) );
  NOR2_X1 U3906 ( .A1(n3035), .A2(n3034), .ZN(n3769) );
  NOR2_X1 U3907 ( .A1(n3768), .A2(n3769), .ZN(n3036) );
  NAND2_X1 U3908 ( .A1(n3038), .A2(n3037), .ZN(n3041) );
  NOR2_X1 U3909 ( .A1(n2131), .A2(n4502), .ZN(n3039) );
  AOI21_X1 U3910 ( .B1(n4518), .B2(n2919), .A(n3039), .ZN(n3042) );
  OAI22_X1 U3911 ( .A1(n4480), .A2(n2131), .B1(n4502), .B2(n3058), .ZN(n3040)
         );
  XNOR2_X1 U3912 ( .A(n3040), .B(n3055), .ZN(n3830) );
  NAND2_X1 U3913 ( .A1(n3828), .A2(n3830), .ZN(n3045) );
  NAND2_X1 U3914 ( .A1(n3771), .A2(n3041), .ZN(n3044) );
  INV_X1 U3915 ( .A(n3042), .ZN(n3043) );
  NAND2_X1 U3916 ( .A1(n3044), .A2(n3043), .ZN(n3827) );
  NAND2_X1 U3917 ( .A1(n3045), .A2(n3827), .ZN(n3792) );
  OAI22_X1 U3918 ( .A1(n4461), .A2(n2131), .B1(n3058), .B2(n4487), .ZN(n3046)
         );
  XOR2_X1 U3919 ( .A(n3046), .B(n3055), .Z(n3049) );
  AOI22_X1 U3920 ( .A1(n4498), .A2(n2919), .B1(n2962), .B2(n3047), .ZN(n3048)
         );
  NAND2_X1 U3921 ( .A1(n3049), .A2(n3048), .ZN(n3793) );
  NOR2_X1 U3922 ( .A1(n3049), .A2(n3048), .ZN(n3795) );
  OAI22_X1 U3923 ( .A1(n4437), .A2(n2131), .B1(n3058), .B2(n4467), .ZN(n3050)
         );
  XNOR2_X1 U3924 ( .A(n3050), .B(n3055), .ZN(n3051) );
  OAI22_X1 U3925 ( .A1(n4437), .A2(n3061), .B1(n2131), .B2(n4467), .ZN(n3052)
         );
  NAND2_X1 U3926 ( .A1(n3051), .A2(n3052), .ZN(n4153) );
  INV_X1 U3927 ( .A(n3051), .ZN(n3054) );
  INV_X1 U3928 ( .A(n3052), .ZN(n3053) );
  NAND2_X1 U3929 ( .A1(n3054), .A2(n3053), .ZN(n4154) );
  OAI22_X1 U3930 ( .A1(n3057), .A2(n2131), .B1(n3058), .B2(n4447), .ZN(n3056)
         );
  XNOR2_X1 U3931 ( .A(n3056), .B(n3055), .ZN(n3075) );
  OAI22_X1 U3932 ( .A1(n3057), .A2(n3061), .B1(n2131), .B2(n4447), .ZN(n3074)
         );
  XNOR2_X1 U3933 ( .A(n3075), .B(n3074), .ZN(n3761) );
  OAI22_X1 U3934 ( .A1(n3062), .A2(n2131), .B1(n3111), .B2(n3058), .ZN(n3060)
         );
  XNOR2_X1 U3935 ( .A(n3060), .B(n3059), .ZN(n3064) );
  OAI22_X1 U3936 ( .A1(n3062), .A2(n3061), .B1(n3111), .B2(n2131), .ZN(n3063)
         );
  XNOR2_X1 U3937 ( .A(n3064), .B(n3063), .ZN(n3095) );
  INV_X1 U3938 ( .A(n3095), .ZN(n3073) );
  INV_X1 U3939 ( .A(n3065), .ZN(n3282) );
  NAND3_X1 U3940 ( .A1(n3067), .A2(n3282), .A3(n3066), .ZN(n3087) );
  INV_X1 U3941 ( .A(n3152), .ZN(n3070) );
  NAND2_X1 U3942 ( .A1(n4901), .A2(n3068), .ZN(n3069) );
  NAND2_X1 U3943 ( .A1(n3070), .A2(n3069), .ZN(n3071) );
  OR2_X1 U3944 ( .A1(n3149), .A2(n3071), .ZN(n3072) );
  NAND2_X1 U3945 ( .A1(n3073), .A2(n4140), .ZN(n3100) );
  NAND2_X1 U3946 ( .A1(n3075), .A2(n3074), .ZN(n3094) );
  NAND2_X1 U3947 ( .A1(n3101), .A2(n3076), .ZN(n3099) );
  INV_X1 U3948 ( .A(n3077), .ZN(n4334) );
  NAND2_X1 U3949 ( .A1(n3078), .A2(n4334), .ZN(n3079) );
  OR2_X1 U3950 ( .A1(n3149), .A2(n3079), .ZN(n3080) );
  NOR2_X1 U3951 ( .A1(n3087), .A2(n3080), .ZN(n3085) );
  NAND2_X1 U3952 ( .A1(n3085), .A2(n4790), .ZN(n4135) );
  NAND2_X1 U3953 ( .A1(n3087), .A2(n3088), .ZN(n3231) );
  NAND2_X1 U3954 ( .A1(n2879), .A2(n3151), .ZN(n3082) );
  NOR2_X1 U3955 ( .A1(n3082), .A2(n3081), .ZN(n3083) );
  NAND2_X1 U3956 ( .A1(n3231), .A2(n3083), .ZN(n3084) );
  INV_X1 U3957 ( .A(n3085), .ZN(n3086) );
  NOR2_X2 U3958 ( .A1(n3086), .A2(n4790), .ZN(n4166) );
  NAND2_X1 U3959 ( .A1(n4240), .A2(n4166), .ZN(n3093) );
  NOR3_X1 U3960 ( .A1(n3087), .A2(n4645), .A3(n3149), .ZN(n3089) );
  AOI22_X1 U3961 ( .A1(n4171), .A2(n3091), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3092) );
  OAI211_X1 U3962 ( .C1(n4169), .C2(n3737), .A(n3093), .B(n3092), .ZN(n3097)
         );
  NOR3_X1 U3963 ( .A1(n3095), .A2(n4175), .A3(n3094), .ZN(n3096) );
  AOI211_X1 U3964 ( .C1(n4167), .C2(n4463), .A(n3097), .B(n3096), .ZN(n3098)
         );
  OAI211_X1 U3965 ( .C1(n3101), .C2(n3100), .A(n3099), .B(n3098), .ZN(U3217)
         );
  XNOR2_X1 U3966 ( .A(n3103), .B(n4248), .ZN(n3107) );
  NAND2_X1 U3967 ( .A1(n4240), .A2(n4660), .ZN(n3105) );
  NAND2_X1 U3968 ( .A1(n4463), .A2(n4630), .ZN(n3104) );
  OAI211_X1 U3969 ( .C1(n3111), .C2(n4645), .A(n3105), .B(n3104), .ZN(n3106)
         );
  OAI21_X1 U3970 ( .B1(n3743), .B2(n4967), .A(n3738), .ZN(n3115) );
  MUX2_X1 U3971 ( .A(REG1_REG_28__SCAN_IN), .B(n3115), .S(n4994), .Z(n3108) );
  INV_X1 U3972 ( .A(n3108), .ZN(n3114) );
  INV_X1 U3973 ( .A(n3109), .ZN(n3112) );
  OAI21_X1 U3974 ( .B1(n3112), .B2(n3111), .A(n3110), .ZN(n3736) );
  NAND2_X1 U3975 ( .A1(n3114), .A2(n3113), .ZN(U3546) );
  MUX2_X1 U3976 ( .A(REG0_REG_28__SCAN_IN), .B(n3115), .S(n4777), .Z(n3116) );
  INV_X1 U3977 ( .A(n3116), .ZN(n3118) );
  NAND2_X1 U3978 ( .A1(n3118), .A2(n3117), .ZN(U3514) );
  INV_X1 U3979 ( .A(DATAI_6_), .ZN(n3120) );
  INV_X1 U3980 ( .A(n3243), .ZN(n3209) );
  MUX2_X1 U3981 ( .A(n3120), .B(n3209), .S(STATE_REG_SCAN_IN), .Z(n3121) );
  INV_X1 U3982 ( .A(n3121), .ZN(U3346) );
  INV_X1 U3983 ( .A(DATAI_3_), .ZN(n3122) );
  MUX2_X1 U3984 ( .A(n3122), .B(n3178), .S(STATE_REG_SCAN_IN), .Z(n3123) );
  INV_X1 U3985 ( .A(n3123), .ZN(U3349) );
  NAND3_X1 U3986 ( .A1(n3961), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3125) );
  INV_X1 U3987 ( .A(DATAI_31_), .ZN(n3124) );
  OAI22_X1 U3988 ( .A1(n2549), .A2(n3125), .B1(STATE_REG_SCAN_IN), .B2(n3124), 
        .ZN(U3321) );
  INV_X1 U3989 ( .A(n3322), .ZN(n3320) );
  INV_X1 U3990 ( .A(DATAI_7_), .ZN(n3126) );
  MUX2_X1 U3991 ( .A(n3320), .B(n3126), .S(U3149), .Z(n3127) );
  INV_X1 U3992 ( .A(n3127), .ZN(U3345) );
  INV_X1 U3993 ( .A(DATAI_21_), .ZN(n3129) );
  NAND2_X1 U3994 ( .A1(n4327), .A2(STATE_REG_SCAN_IN), .ZN(n3128) );
  OAI21_X1 U3995 ( .B1(STATE_REG_SCAN_IN), .B2(n3129), .A(n3128), .ZN(U3331)
         );
  MUX2_X1 U3996 ( .A(n3373), .B(n3130), .S(U3149), .Z(n3131) );
  INV_X1 U3997 ( .A(n3131), .ZN(U3344) );
  INV_X1 U3998 ( .A(DATAI_27_), .ZN(n3133) );
  NAND2_X1 U3999 ( .A1(n3167), .A2(STATE_REG_SCAN_IN), .ZN(n3132) );
  OAI21_X1 U4000 ( .B1(STATE_REG_SCAN_IN), .B2(n3133), .A(n3132), .ZN(U3325)
         );
  NAND2_X1 U4001 ( .A1(U3149), .A2(DATAI_25_), .ZN(n3134) );
  OAI21_X1 U4002 ( .B1(n3135), .B2(U3149), .A(n3134), .ZN(U3327) );
  INV_X1 U4003 ( .A(DATAI_29_), .ZN(n3138) );
  NAND2_X1 U4004 ( .A1(n3136), .A2(STATE_REG_SCAN_IN), .ZN(n3137) );
  OAI21_X1 U4005 ( .B1(STATE_REG_SCAN_IN), .B2(n3138), .A(n3137), .ZN(U3323)
         );
  INV_X1 U4006 ( .A(DATAI_24_), .ZN(n3945) );
  MUX2_X1 U4007 ( .A(n3139), .B(n3945), .S(U3149), .Z(n3140) );
  INV_X1 U4008 ( .A(n3140), .ZN(U3328) );
  INV_X1 U4009 ( .A(n3149), .ZN(n3142) );
  INV_X1 U4010 ( .A(D_REG_0__SCAN_IN), .ZN(n3994) );
  INV_X1 U4011 ( .A(n3143), .ZN(n3144) );
  AOI22_X1 U4012 ( .A1(n4928), .A2(n3994), .B1(n3144), .B2(n4931), .ZN(U3458)
         );
  INV_X1 U4013 ( .A(D_REG_1__SCAN_IN), .ZN(n3147) );
  INV_X1 U4014 ( .A(n3145), .ZN(n3146) );
  AOI22_X1 U4015 ( .A1(n4928), .A2(n3147), .B1(n4931), .B2(n3146), .ZN(U3459)
         );
  INV_X1 U4016 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n3969) );
  NAND2_X1 U4017 ( .A1(n3624), .A2(U4043), .ZN(n3148) );
  OAI21_X1 U4018 ( .B1(U4043), .B2(n3969), .A(n3148), .ZN(U3562) );
  OR2_X1 U4019 ( .A1(n3151), .A2(U3149), .ZN(n4337) );
  NAND2_X1 U4020 ( .A1(n3149), .A2(n4337), .ZN(n3155) );
  AOI21_X1 U4021 ( .B1(n3152), .B2(n3151), .A(n3150), .ZN(n3154) );
  INV_X1 U4022 ( .A(n3154), .ZN(n3153) );
  INV_X1 U4023 ( .A(n4881), .ZN(n3638) );
  INV_X1 U4024 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n3159) );
  INV_X1 U4025 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4915) );
  AOI21_X1 U4026 ( .B1(n3167), .B2(n4915), .A(n3175), .ZN(n4361) );
  OAI21_X1 U4027 ( .B1(REG1_REG_0__SCAN_IN), .B2(n3167), .A(n4361), .ZN(n3156)
         );
  XOR2_X1 U4028 ( .A(n4943), .B(n3156), .Z(n3157) );
  AOI22_X1 U4029 ( .A1(n3176), .A2(n3157), .B1(REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n3158) );
  OAI21_X1 U4030 ( .B1(n3638), .B2(n3159), .A(n3158), .ZN(U3240) );
  INV_X1 U4031 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n3917) );
  NAND2_X1 U4032 ( .A1(n3397), .A2(U4043), .ZN(n3160) );
  OAI21_X1 U4033 ( .B1(U4043), .B2(n3917), .A(n3160), .ZN(U3557) );
  NAND2_X1 U4034 ( .A1(n3169), .A2(REG2_REG_1__SCAN_IN), .ZN(n3161) );
  AND2_X1 U4035 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4359)
         );
  NAND2_X1 U4036 ( .A1(n4349), .A2(n4359), .ZN(n4348) );
  NAND2_X1 U4037 ( .A1(n4798), .A2(REG2_REG_1__SCAN_IN), .ZN(n4370) );
  NAND2_X1 U4038 ( .A1(n4348), .A2(n4370), .ZN(n3165) );
  INV_X1 U4039 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3163) );
  MUX2_X1 U4040 ( .A(REG2_REG_2__SCAN_IN), .B(n3163), .S(n2130), .Z(n4368) );
  NAND2_X1 U4041 ( .A1(n3165), .A2(n4368), .ZN(n4372) );
  NAND2_X1 U4042 ( .A1(n2130), .A2(REG2_REG_2__SCAN_IN), .ZN(n3166) );
  XNOR2_X1 U40430 ( .A(n3192), .B(n3178), .ZN(n3190) );
  XNOR2_X1 U4044 ( .A(n3190), .B(REG2_REG_3__SCAN_IN), .ZN(n3182) );
  INV_X1 U4045 ( .A(n3167), .ZN(n4358) );
  NOR2_X1 U4046 ( .A1(n4358), .A2(n3175), .ZN(n4333) );
  INV_X1 U4047 ( .A(REG1_REG_1__SCAN_IN), .ZN(n3168) );
  INV_X1 U4048 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4982) );
  NOR2_X1 U4049 ( .A1(n4943), .A2(n4982), .ZN(n4351) );
  NAND2_X1 U4050 ( .A1(n4798), .A2(REG1_REG_1__SCAN_IN), .ZN(n4363) );
  NAND2_X1 U4051 ( .A1(n4364), .A2(n4363), .ZN(n3173) );
  MUX2_X1 U4052 ( .A(n4018), .B(REG1_REG_2__SCAN_IN), .S(n3164), .Z(n4362) );
  INV_X1 U4053 ( .A(n4362), .ZN(n3172) );
  NAND2_X1 U4054 ( .A1(n2130), .A2(REG1_REG_2__SCAN_IN), .ZN(n3174) );
  XOR2_X1 U4055 ( .A(n3183), .B(REG1_REG_3__SCAN_IN), .Z(n3180) );
  INV_X1 U4056 ( .A(n4849), .ZN(n4892) );
  AOI22_X1 U4057 ( .A1(n4881), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3177) );
  OAI21_X1 U4058 ( .B1(n4892), .B2(n3178), .A(n3177), .ZN(n3179) );
  AOI21_X1 U4059 ( .B1(n4873), .B2(n3180), .A(n3179), .ZN(n3181) );
  OAI21_X1 U4060 ( .B1(n3182), .B2(n4878), .A(n3181), .ZN(U3243) );
  NAND2_X1 U4061 ( .A1(n3183), .A2(REG1_REG_3__SCAN_IN), .ZN(n3186) );
  NAND2_X1 U4062 ( .A1(n3184), .A2(n3191), .ZN(n3185) );
  INV_X1 U4063 ( .A(n4820), .ZN(n3195) );
  INV_X1 U4064 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4989) );
  MUX2_X1 U4065 ( .A(REG1_REG_5__SCAN_IN), .B(n4989), .S(n3204), .Z(n3189) );
  INV_X1 U4066 ( .A(n4873), .ZN(n4887) );
  NAND2_X1 U4067 ( .A1(n3190), .A2(REG2_REG_3__SCAN_IN), .ZN(n3194) );
  NAND2_X1 U4068 ( .A1(n3192), .A2(n3191), .ZN(n3193) );
  INV_X1 U4069 ( .A(REG2_REG_5__SCAN_IN), .ZN(n4030) );
  MUX2_X1 U4070 ( .A(REG2_REG_5__SCAN_IN), .B(n4030), .S(n3204), .Z(n3198) );
  AOI211_X1 U4071 ( .C1(n3197), .C2(n3198), .A(n4878), .B(n3205), .ZN(n3201)
         );
  AND2_X1 U4072 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3257) );
  AOI21_X1 U4073 ( .B1(n4881), .B2(ADDR_REG_5__SCAN_IN), .A(n3257), .ZN(n3199)
         );
  OAI21_X1 U4074 ( .B1(n4892), .B2(n3204), .A(n3199), .ZN(n3200) );
  OR3_X1 U4075 ( .A1(n3202), .A2(n3201), .A3(n3200), .ZN(U3245) );
  NOR2_X1 U4076 ( .A1(n4881), .A2(n3562), .ZN(U3148) );
  INV_X1 U4077 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n3934) );
  NAND2_X1 U4078 ( .A1(n3694), .A2(U4043), .ZN(n3203) );
  OAI21_X1 U4079 ( .B1(n3562), .B2(n3934), .A(n3203), .ZN(U3565) );
  INV_X1 U4080 ( .A(n3204), .ZN(n4796) );
  XNOR2_X1 U4081 ( .A(n3244), .B(REG2_REG_6__SCAN_IN), .ZN(n3213) );
  XOR2_X1 U4082 ( .A(n3237), .B(REG1_REG_6__SCAN_IN), .Z(n3211) );
  NAND2_X1 U4083 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3275) );
  NAND2_X1 U4084 ( .A1(n4881), .A2(ADDR_REG_6__SCAN_IN), .ZN(n3208) );
  OAI211_X1 U4085 ( .C1(n4892), .C2(n3209), .A(n3275), .B(n3208), .ZN(n3210)
         );
  AOI21_X1 U4086 ( .B1(n3211), .B2(n4873), .A(n3210), .ZN(n3212) );
  OAI21_X1 U4087 ( .B1(n3213), .B2(n4878), .A(n3212), .ZN(U3246) );
  INV_X1 U4088 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n4003) );
  NAND2_X1 U4089 ( .A1(n3753), .A2(n3562), .ZN(n3214) );
  OAI21_X1 U4090 ( .B1(U4043), .B2(n4003), .A(n3214), .ZN(U3556) );
  INV_X1 U4091 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n4000) );
  NAND2_X1 U4092 ( .A1(n2586), .A2(REG1_REG_31__SCAN_IN), .ZN(n3218) );
  NAND2_X1 U4093 ( .A1(n2585), .A2(REG0_REG_31__SCAN_IN), .ZN(n3217) );
  NAND2_X1 U4094 ( .A1(n3215), .A2(REG2_REG_31__SCAN_IN), .ZN(n3216) );
  NAND3_X1 U4095 ( .A1(n3218), .A2(n3217), .A3(n3216), .ZN(n4412) );
  NAND2_X1 U4096 ( .A1(n4412), .A2(n3562), .ZN(n3219) );
  OAI21_X1 U4097 ( .B1(n4000), .B2(U4043), .A(n3219), .ZN(U3581) );
  INV_X1 U4098 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n3974) );
  NAND2_X1 U4099 ( .A1(n4629), .A2(n3562), .ZN(n3220) );
  OAI21_X1 U4100 ( .B1(n3562), .B2(n3974), .A(n3220), .ZN(U3566) );
  INV_X1 U4101 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n3935) );
  NAND2_X1 U4102 ( .A1(n3820), .A2(n3562), .ZN(n3221) );
  OAI21_X1 U4103 ( .B1(U4043), .B2(n3935), .A(n3221), .ZN(U3568) );
  INV_X1 U4104 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n4006) );
  NAND2_X1 U4105 ( .A1(n3222), .A2(n3562), .ZN(n3223) );
  OAI21_X1 U4106 ( .B1(U4043), .B2(n4006), .A(n3223), .ZN(U3560) );
  INV_X1 U4107 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n3916) );
  NAND2_X1 U4108 ( .A1(n3336), .A2(n3562), .ZN(n3224) );
  OAI21_X1 U4109 ( .B1(U4043), .B2(n3916), .A(n3224), .ZN(U3553) );
  INV_X1 U4110 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n3968) );
  NAND2_X1 U4111 ( .A1(n3589), .A2(n3562), .ZN(n3225) );
  OAI21_X1 U4112 ( .B1(n3562), .B2(n3968), .A(n3225), .ZN(U3563) );
  INV_X1 U4113 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n3931) );
  NAND2_X1 U4114 ( .A1(n2578), .A2(n3562), .ZN(n3226) );
  OAI21_X1 U4115 ( .B1(U4043), .B2(n3931), .A(n3226), .ZN(U3551) );
  INV_X1 U4116 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4002) );
  NAND2_X1 U4117 ( .A1(n4610), .A2(n3562), .ZN(n3227) );
  OAI21_X1 U4118 ( .B1(U4043), .B2(n4002), .A(n3227), .ZN(U3569) );
  XNOR2_X1 U4119 ( .A(n3228), .B(n3229), .ZN(n3234) );
  AND2_X1 U4120 ( .A1(n3231), .A2(n3230), .ZN(n4134) );
  INV_X1 U4121 ( .A(n4134), .ZN(n3746) );
  AOI22_X1 U4122 ( .A1(n4171), .A2(n3291), .B1(REG3_REG_1__SCAN_IN), .B2(n3746), .ZN(n3233) );
  AOI22_X1 U4123 ( .A1(n4167), .A2(n2881), .B1(n4166), .B2(n4347), .ZN(n3232)
         );
  OAI211_X1 U4124 ( .C1(n3234), .C2(n4175), .A(n3233), .B(n3232), .ZN(U3219)
         );
  INV_X1 U4125 ( .A(n3235), .ZN(n3236) );
  INV_X1 U4126 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4992) );
  XNOR2_X1 U4127 ( .A(n3322), .B(n4992), .ZN(n3238) );
  XNOR2_X1 U4128 ( .A(n3239), .B(n3238), .ZN(n3249) );
  NOR2_X1 U4129 ( .A1(STATE_REG_SCAN_IN), .A2(n2611), .ZN(n3756) );
  AOI21_X1 U4130 ( .B1(n4881), .B2(ADDR_REG_7__SCAN_IN), .A(n3756), .ZN(n3240)
         );
  OAI21_X1 U4131 ( .B1(n4892), .B2(n3320), .A(n3240), .ZN(n3248) );
  INV_X1 U4132 ( .A(n3241), .ZN(n3242) );
  INV_X1 U4133 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4037) );
  MUX2_X1 U4134 ( .A(n4037), .B(REG2_REG_7__SCAN_IN), .S(n3322), .Z(n3245) );
  AOI211_X1 U4135 ( .C1(n3246), .C2(n3245), .A(n4878), .B(n3318), .ZN(n3247)
         );
  AOI211_X1 U4136 ( .C1(n3249), .C2(n4873), .A(n3248), .B(n3247), .ZN(n3250)
         );
  INV_X1 U4137 ( .A(n3250), .ZN(U3247) );
  INV_X1 U4138 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n3977) );
  NAND2_X1 U4139 ( .A1(n4593), .A2(n3562), .ZN(n3251) );
  OAI21_X1 U4140 ( .B1(U4043), .B2(n3977), .A(n3251), .ZN(U3570) );
  INV_X1 U4141 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n3928) );
  NAND2_X1 U4142 ( .A1(n4534), .A2(n3562), .ZN(n3252) );
  OAI21_X1 U4143 ( .B1(U4043), .B2(n3928), .A(n3252), .ZN(U3571) );
  XNOR2_X1 U4144 ( .A(n3254), .B(n3253), .ZN(n3260) );
  AOI22_X1 U4145 ( .A1(n4167), .A2(n4346), .B1(n4166), .B2(n3753), .ZN(n3259)
         );
  NOR2_X1 U4146 ( .A1(n3090), .A2(n3255), .ZN(n3256) );
  AOI211_X1 U4147 ( .C1(n3845), .C2(n3426), .A(n3257), .B(n3256), .ZN(n3258)
         );
  OAI211_X1 U4148 ( .C1(n3260), .C2(n4175), .A(n3259), .B(n3258), .ZN(U3224)
         );
  INV_X1 U4149 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n3908) );
  NAND2_X1 U4150 ( .A1(n4552), .A2(n3562), .ZN(n3261) );
  OAI21_X1 U4151 ( .B1(U4043), .B2(n3908), .A(n3261), .ZN(U3572) );
  OAI21_X1 U4152 ( .B1(n3265), .B2(n3262), .A(n3264), .ZN(n3270) );
  MUX2_X1 U4153 ( .A(U3149), .B(n3845), .S(n3266), .Z(n3269) );
  AOI22_X1 U4154 ( .A1(n4171), .A2(n3368), .B1(n4167), .B2(n4347), .ZN(n3267)
         );
  OAI21_X1 U4155 ( .B1(n3420), .B2(n4137), .A(n3267), .ZN(n3268) );
  AOI211_X1 U4156 ( .C1(n3270), .C2(n4140), .A(n3269), .B(n3268), .ZN(n3271)
         );
  INV_X1 U4157 ( .A(n3271), .ZN(U3215) );
  NAND2_X1 U4158 ( .A1(n2183), .A2(n3272), .ZN(n3273) );
  XNOR2_X1 U4159 ( .A(n3274), .B(n3273), .ZN(n3279) );
  OAI22_X1 U4160 ( .A1(n4137), .A2(n3353), .B1(n3716), .B2(n4135), .ZN(n3277)
         );
  OAI21_X1 U4161 ( .B1(n3090), .B2(n3502), .A(n3275), .ZN(n3276) );
  AOI211_X1 U4162 ( .C1(n3511), .C2(n3845), .A(n3277), .B(n3276), .ZN(n3278)
         );
  OAI21_X1 U4163 ( .B1(n3279), .B2(n4175), .A(n3278), .ZN(U3236) );
  INV_X1 U4164 ( .A(n3280), .ZN(n3283) );
  NAND3_X1 U4165 ( .A1(n3283), .A2(n3282), .A3(n3281), .ZN(n3284) );
  OAI21_X1 U4166 ( .B1(n4903), .B2(n3286), .A(n3285), .ZN(n4948) );
  OR2_X1 U4167 ( .A1(n3288), .A2(n3287), .ZN(n3289) );
  NAND2_X1 U4168 ( .A1(n3290), .A2(n3289), .ZN(n4950) );
  NAND2_X1 U4169 ( .A1(n4568), .A2(n3291), .ZN(n3293) );
  NAND2_X1 U4170 ( .A1(n2881), .A2(n4630), .ZN(n3292) );
  OAI211_X1 U4171 ( .C1(n3294), .C2(n4908), .A(n3293), .B(n3292), .ZN(n3295)
         );
  INV_X1 U4172 ( .A(n3295), .ZN(n3298) );
  XNOR2_X1 U4173 ( .A(n3287), .B(n4257), .ZN(n3296) );
  NAND2_X1 U4174 ( .A1(n3296), .A2(n4906), .ZN(n3297) );
  OAI211_X1 U4175 ( .C1(n4950), .C2(n4905), .A(n3298), .B(n3297), .ZN(n4952)
         );
  MUX2_X1 U4176 ( .A(n4952), .B(REG2_REG_1__SCAN_IN), .S(n4643), .Z(n3299) );
  INV_X1 U4177 ( .A(n3299), .ZN(n3304) );
  INV_X1 U4178 ( .A(n4950), .ZN(n3302) );
  OR2_X1 U4179 ( .A1(n3300), .A2(n4812), .ZN(n3413) );
  INV_X1 U4180 ( .A(n3413), .ZN(n3301) );
  AOI22_X1 U4181 ( .A1(n3302), .A2(n4913), .B1(REG3_REG_1__SCAN_IN), .B2(n4912), .ZN(n3303) );
  OAI211_X1 U4182 ( .C1(n4600), .C2(n4948), .A(n3304), .B(n3303), .ZN(U3289)
         );
  INV_X1 U4183 ( .A(n3305), .ZN(n3306) );
  AOI21_X1 U4184 ( .B1(n4276), .B2(n3307), .A(n3306), .ZN(n4893) );
  OAI21_X1 U4185 ( .B1(n4276), .B2(n3309), .A(n3308), .ZN(n3313) );
  AOI22_X1 U4186 ( .A1(n2578), .A2(n4630), .B1(n3314), .B2(n4568), .ZN(n3310)
         );
  OAI21_X1 U4187 ( .B1(n4136), .B2(n4908), .A(n3310), .ZN(n3312) );
  NOR2_X1 U4188 ( .A1(n4893), .A2(n4905), .ZN(n3311) );
  AOI211_X1 U4189 ( .C1(n4906), .C2(n3313), .A(n3312), .B(n3311), .ZN(n4900)
         );
  OAI21_X1 U4190 ( .B1(n4893), .B2(n4954), .A(n4900), .ZN(n3430) );
  NAND2_X1 U4191 ( .A1(n3285), .A2(n3314), .ZN(n3315) );
  NAND2_X1 U4192 ( .A1(n3367), .A2(n3315), .ZN(n4894) );
  OAI22_X1 U4193 ( .A1(n4738), .A2(n4894), .B1(n4994), .B2(n4018), .ZN(n3316)
         );
  AOI21_X1 U4194 ( .B1(n3430), .B2(n4994), .A(n3316), .ZN(n3317) );
  INV_X1 U4195 ( .A(n3317), .ZN(U3520) );
  XOR2_X1 U4196 ( .A(REG2_REG_8__SCAN_IN), .B(n3376), .Z(n3326) );
  NAND2_X1 U4197 ( .A1(U3149), .A2(REG3_REG_8__SCAN_IN), .ZN(n3354) );
  NAND2_X1 U4198 ( .A1(n4881), .A2(ADDR_REG_8__SCAN_IN), .ZN(n3319) );
  OAI211_X1 U4199 ( .C1(n4892), .C2(n3373), .A(n3354), .B(n3319), .ZN(n3325)
         );
  INV_X1 U4200 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4054) );
  XNOR2_X1 U4201 ( .A(n3382), .B(n3373), .ZN(n3323) );
  AOI211_X1 U4202 ( .C1(n4054), .C2(n3323), .A(n4887), .B(n3385), .ZN(n3324)
         );
  AOI211_X1 U4203 ( .C1(n4875), .C2(n3326), .A(n3325), .B(n3324), .ZN(n3327)
         );
  INV_X1 U4204 ( .A(n3327), .ZN(U3248) );
  INV_X1 U4205 ( .A(REG1_REG_6__SCAN_IN), .ZN(n4099) );
  NAND2_X1 U4206 ( .A1(n4193), .A2(n4202), .ZN(n4285) );
  XNOR2_X1 U4207 ( .A(n3328), .B(n4285), .ZN(n3514) );
  XOR2_X1 U4208 ( .A(n2177), .B(n4285), .Z(n3331) );
  AOI22_X1 U4209 ( .A1(n4345), .A2(n4630), .B1(n4568), .B2(n3332), .ZN(n3329)
         );
  OAI21_X1 U4210 ( .B1(n3353), .B2(n4908), .A(n3329), .ZN(n3330) );
  AOI21_X1 U4211 ( .B1(n3331), .B2(n4906), .A(n3330), .ZN(n3519) );
  OAI21_X1 U4212 ( .B1(n4967), .B2(n3514), .A(n3519), .ZN(n3454) );
  NAND2_X1 U4213 ( .A1(n3454), .A2(n4994), .ZN(n3335) );
  AND2_X1 U4214 ( .A1(n2185), .A2(n3332), .ZN(n3333) );
  NOR2_X1 U4215 ( .A1(n2133), .A2(n3333), .ZN(n3517) );
  INV_X1 U4216 ( .A(n4738), .ZN(n4676) );
  NAND2_X1 U4217 ( .A1(n3517), .A2(n4676), .ZN(n3334) );
  OAI211_X1 U4218 ( .C1(n4994), .C2(n4099), .A(n3335), .B(n3334), .ZN(U3524)
         );
  OAI211_X1 U4219 ( .C1(n3366), .C2(n3717), .A(n3424), .B(n4972), .ZN(n4960)
         );
  NOR2_X1 U4220 ( .A1(n4960), .A2(n4802), .ZN(n3344) );
  NAND2_X1 U4221 ( .A1(n3336), .A2(n4630), .ZN(n3337) );
  OAI21_X1 U4222 ( .B1(n4645), .B2(n3717), .A(n3337), .ZN(n3341) );
  OR2_X1 U4223 ( .A1(n3338), .A2(n4272), .ZN(n3416) );
  NAND2_X1 U4224 ( .A1(n3338), .A2(n4272), .ZN(n3339) );
  NAND2_X1 U4225 ( .A1(n3416), .A2(n3339), .ZN(n3345) );
  NOR2_X1 U4226 ( .A1(n3345), .A2(n4905), .ZN(n3340) );
  AOI211_X1 U4227 ( .C1(n4660), .C2(n4345), .A(n3341), .B(n3340), .ZN(n3342)
         );
  OAI21_X1 U4228 ( .B1(n4655), .B2(n3343), .A(n3342), .ZN(n4961) );
  AOI211_X1 U4229 ( .C1(n4912), .C2(n3720), .A(n3344), .B(n4961), .ZN(n3347)
         );
  INV_X1 U4230 ( .A(n3345), .ZN(n4964) );
  AOI22_X1 U4231 ( .A1(n4964), .A2(n4913), .B1(REG2_REG_4__SCAN_IN), .B2(n4643), .ZN(n3346) );
  OAI21_X1 U4232 ( .B1(n3347), .B2(n4643), .A(n3346), .ZN(U3286) );
  INV_X1 U4233 ( .A(n3348), .ZN(n3350) );
  NOR2_X1 U4234 ( .A1(n3350), .A2(n3349), .ZN(n3351) );
  XNOR2_X1 U4235 ( .A(n3352), .B(n3351), .ZN(n3358) );
  OAI22_X1 U4236 ( .A1(n4137), .A2(n3447), .B1(n3353), .B2(n4135), .ZN(n3356)
         );
  OAI21_X1 U4237 ( .B1(n3090), .B2(n3395), .A(n3354), .ZN(n3355) );
  AOI211_X1 U4238 ( .C1(n3536), .C2(n3845), .A(n3356), .B(n3355), .ZN(n3357)
         );
  OAI21_X1 U4239 ( .B1(n3358), .B2(n4175), .A(n3357), .ZN(U3218) );
  INV_X1 U4240 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n3995) );
  NAND2_X1 U4241 ( .A1(n4518), .A2(n3562), .ZN(n3359) );
  OAI21_X1 U4242 ( .B1(U4043), .B2(n3995), .A(n3359), .ZN(U3574) );
  XNOR2_X1 U4243 ( .A(n3360), .B(n4271), .ZN(n4955) );
  INV_X1 U4244 ( .A(n4913), .ZN(n4673) );
  XNOR2_X1 U4245 ( .A(n3361), .B(n4271), .ZN(n3364) );
  AOI22_X1 U4246 ( .A1(n4347), .A2(n4630), .B1(n4568), .B2(n3368), .ZN(n3362)
         );
  OAI21_X1 U4247 ( .B1(n3420), .B2(n4908), .A(n3362), .ZN(n3363) );
  AOI21_X1 U4248 ( .B1(n3364), .B2(n4906), .A(n3363), .ZN(n3365) );
  OAI21_X1 U4249 ( .B1(n4955), .B2(n4905), .A(n3365), .ZN(n4956) );
  NAND2_X1 U4250 ( .A1(n4956), .A2(n4668), .ZN(n3372) );
  AOI21_X1 U4251 ( .B1(n3368), .B2(n3367), .A(n3366), .ZN(n4958) );
  INV_X1 U4252 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3369) );
  OAI22_X1 U4253 ( .A1(n4668), .A2(n3369), .B1(REG3_REG_3__SCAN_IN), .B2(n4665), .ZN(n3370) );
  AOI21_X1 U4254 ( .B1(n4896), .B2(n4958), .A(n3370), .ZN(n3371) );
  OAI211_X1 U4255 ( .C1(n4955), .C2(n4673), .A(n3372), .B(n3371), .ZN(U3287)
         );
  INV_X1 U4256 ( .A(n3373), .ZN(n3383) );
  INV_X1 U4257 ( .A(n3374), .ZN(n3375) );
  INV_X1 U4258 ( .A(REG2_REG_9__SCAN_IN), .ZN(n4036) );
  MUX2_X1 U4259 ( .A(REG2_REG_9__SCAN_IN), .B(n4036), .S(n3437), .Z(n3380) );
  INV_X1 U4260 ( .A(n3380), .ZN(n3377) );
  NAND2_X1 U4261 ( .A1(n3378), .A2(n3377), .ZN(n3434) );
  INV_X1 U4262 ( .A(n3434), .ZN(n3379) );
  AOI211_X1 U4263 ( .C1(n3381), .C2(n3380), .A(n4878), .B(n3379), .ZN(n3391)
         );
  XOR2_X1 U4264 ( .A(REG1_REG_9__SCAN_IN), .B(n3437), .Z(n3386) );
  AOI211_X1 U4265 ( .C1(n3387), .C2(n3386), .A(n4887), .B(n2172), .ZN(n3390)
         );
  NAND2_X1 U4266 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n3408) );
  NAND2_X1 U4267 ( .A1(n4881), .A2(ADDR_REG_9__SCAN_IN), .ZN(n3388) );
  OAI211_X1 U4268 ( .C1(n4892), .C2(n3437), .A(n3408), .B(n3388), .ZN(n3389)
         );
  OR3_X1 U4269 ( .A1(n3391), .A2(n3390), .A3(n3389), .ZN(U3249) );
  NAND2_X1 U4270 ( .A1(n3393), .A2(n3392), .ZN(n3461) );
  AND2_X1 U4271 ( .A1(n4198), .A2(n4196), .ZN(n4275) );
  XNOR2_X1 U4272 ( .A(n3461), .B(n4275), .ZN(n3540) );
  XNOR2_X1 U4273 ( .A(n3394), .B(n4275), .ZN(n3400) );
  NOR2_X1 U4274 ( .A1(n4645), .A2(n3395), .ZN(n3396) );
  AOI21_X1 U4275 ( .B1(n4343), .B2(n4660), .A(n3396), .ZN(n3399) );
  NAND2_X1 U4276 ( .A1(n3397), .A2(n4630), .ZN(n3398) );
  OAI211_X1 U4277 ( .C1(n3400), .C2(n4655), .A(n3399), .B(n3398), .ZN(n3534)
         );
  AOI21_X1 U4278 ( .B1(n3540), .B2(n4975), .A(n3534), .ZN(n3459) );
  INV_X1 U4279 ( .A(n3401), .ZN(n3498) );
  INV_X1 U4280 ( .A(n3402), .ZN(n3403) );
  AOI21_X1 U4281 ( .B1(n3404), .B2(n3498), .A(n3403), .ZN(n3535) );
  AOI22_X1 U4282 ( .A1(n3535), .A2(n4676), .B1(REG1_REG_8__SCAN_IN), .B2(n4991), .ZN(n3405) );
  OAI21_X1 U4283 ( .B1(n3459), .B2(n4991), .A(n3405), .ZN(U3526) );
  XOR2_X1 U4284 ( .A(n3407), .B(n3406), .Z(n3412) );
  OAI22_X1 U4285 ( .A1(n4137), .A2(n3569), .B1(n3495), .B2(n4135), .ZN(n3410)
         );
  OAI21_X1 U4286 ( .B1(n3090), .B2(n3466), .A(n3408), .ZN(n3409) );
  AOI211_X1 U4287 ( .C1(n3478), .C2(n3845), .A(n3410), .B(n3409), .ZN(n3411)
         );
  OAI21_X1 U4288 ( .B1(n3412), .B2(n4175), .A(n3411), .ZN(U3228) );
  NAND2_X1 U4289 ( .A1(n4905), .A2(n3413), .ZN(n3414) );
  AND2_X1 U4290 ( .A1(n2167), .A2(n4204), .ZN(n4277) );
  NAND2_X1 U4291 ( .A1(n3416), .A2(n3415), .ZN(n3417) );
  XOR2_X1 U4292 ( .A(n4277), .B(n3417), .Z(n4968) );
  XOR2_X1 U4293 ( .A(n4277), .B(n3418), .Z(n3422) );
  AOI22_X1 U4294 ( .A1(n3753), .A2(n4660), .B1(n3425), .B2(n4568), .ZN(n3419)
         );
  OAI21_X1 U4295 ( .B1(n3420), .B2(n4647), .A(n3419), .ZN(n3421) );
  AOI21_X1 U4296 ( .B1(n3422), .B2(n4906), .A(n3421), .ZN(n4966) );
  MUX2_X1 U4297 ( .A(n4966), .B(n4030), .S(n4643), .Z(n3428) );
  INV_X1 U4298 ( .A(n2185), .ZN(n3423) );
  AOI21_X1 U4299 ( .B1(n3425), .B2(n3424), .A(n3423), .ZN(n4971) );
  AOI22_X1 U4300 ( .A1(n4896), .A2(n4971), .B1(n3426), .B2(n4912), .ZN(n3427)
         );
  OAI211_X1 U4301 ( .C1(n4603), .C2(n4968), .A(n3428), .B(n3427), .ZN(U3285)
         );
  INV_X1 U4302 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3943) );
  OAI22_X1 U4303 ( .A1(n4787), .A2(n4894), .B1(n4777), .B2(n3943), .ZN(n3429)
         );
  AOI21_X1 U4304 ( .B1(n3430), .B2(n4777), .A(n3429), .ZN(n3431) );
  INV_X1 U4305 ( .A(n3431), .ZN(U3471) );
  XNOR2_X1 U4306 ( .A(n3548), .B(REG2_REG_10__SCAN_IN), .ZN(n3442) );
  NAND2_X1 U4307 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n3448) );
  INV_X1 U4308 ( .A(n3448), .ZN(n3436) );
  NOR2_X1 U4309 ( .A1(n4892), .A2(n3555), .ZN(n3435) );
  AOI211_X1 U4310 ( .C1(n4881), .C2(ADDR_REG_10__SCAN_IN), .A(n3436), .B(n3435), .ZN(n3441) );
  NAND2_X1 U4311 ( .A1(n3439), .A2(REG1_REG_10__SCAN_IN), .ZN(n3557) );
  OAI211_X1 U4312 ( .C1(n3439), .C2(REG1_REG_10__SCAN_IN), .A(n3557), .B(n4873), .ZN(n3440) );
  OAI211_X1 U4313 ( .C1(n3442), .C2(n4878), .A(n3441), .B(n3440), .ZN(U3250)
         );
  INV_X1 U4314 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n3966) );
  NAND2_X1 U4315 ( .A1(n4498), .A2(n3562), .ZN(n3443) );
  OAI21_X1 U4316 ( .B1(U4043), .B2(n3966), .A(n3443), .ZN(U3575) );
  OAI211_X1 U4317 ( .C1(n3446), .C2(n3445), .A(n3444), .B(n4140), .ZN(n3453)
         );
  OAI22_X1 U4318 ( .A1(n4137), .A2(n3727), .B1(n3447), .B2(n4135), .ZN(n3451)
         );
  OAI21_X1 U4319 ( .B1(n3090), .B2(n3449), .A(n3448), .ZN(n3450) );
  AOI211_X1 U4320 ( .C1(n3528), .C2(n3845), .A(n3451), .B(n3450), .ZN(n3452)
         );
  NAND2_X1 U4321 ( .A1(n3453), .A2(n3452), .ZN(U3214) );
  INV_X1 U4322 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3457) );
  NAND2_X1 U4323 ( .A1(n3454), .A2(n4777), .ZN(n3456) );
  INV_X1 U4324 ( .A(n4787), .ZN(n4743) );
  NAND2_X1 U4325 ( .A1(n3517), .A2(n4743), .ZN(n3455) );
  OAI211_X1 U4326 ( .C1(n4777), .C2(n3457), .A(n3456), .B(n3455), .ZN(U3479)
         );
  AOI22_X1 U4327 ( .A1(n3535), .A2(n4743), .B1(REG0_REG_8__SCAN_IN), .B2(n4980), .ZN(n3458) );
  OAI21_X1 U4328 ( .B1(n3459), .B2(n4980), .A(n3458), .ZN(U3483) );
  NAND2_X1 U4329 ( .A1(n3461), .A2(n3460), .ZN(n3463) );
  NAND2_X1 U4330 ( .A1(n3463), .A2(n3462), .ZN(n3464) );
  AND2_X1 U4331 ( .A1(n2335), .A2(n4199), .ZN(n4263) );
  XNOR2_X1 U4332 ( .A(n3464), .B(n4263), .ZN(n3475) );
  XNOR2_X1 U4333 ( .A(n3465), .B(n4263), .ZN(n3469) );
  OAI22_X1 U4334 ( .A1(n3569), .A2(n4908), .B1(n4645), .B2(n3466), .ZN(n3467)
         );
  AOI21_X1 U4335 ( .B1(n4630), .B2(n4344), .A(n3467), .ZN(n3468) );
  OAI21_X1 U4336 ( .B1(n3469), .B2(n4655), .A(n3468), .ZN(n3476) );
  AOI21_X1 U4337 ( .B1(n3475), .B2(n4975), .A(n3476), .ZN(n3474) );
  NAND2_X1 U4338 ( .A1(n3402), .A2(n3470), .ZN(n3471) );
  AND2_X1 U4339 ( .A1(n3526), .A2(n3471), .ZN(n3479) );
  AOI22_X1 U4340 ( .A1(n3479), .A2(n4743), .B1(REG0_REG_9__SCAN_IN), .B2(n4980), .ZN(n3472) );
  OAI21_X1 U4341 ( .B1(n3474), .B2(n4980), .A(n3472), .ZN(U3485) );
  AOI22_X1 U4342 ( .A1(n3479), .A2(n4676), .B1(REG1_REG_9__SCAN_IN), .B2(n4991), .ZN(n3473) );
  OAI21_X1 U4343 ( .B1(n3474), .B2(n4991), .A(n3473), .ZN(U3527) );
  INV_X1 U4344 ( .A(n3475), .ZN(n3482) );
  INV_X1 U4345 ( .A(n3476), .ZN(n3477) );
  MUX2_X1 U4346 ( .A(n4036), .B(n3477), .S(n4668), .Z(n3481) );
  AOI22_X1 U4347 ( .A1(n3479), .A2(n4896), .B1(n3478), .B2(n4912), .ZN(n3480)
         );
  OAI211_X1 U4348 ( .C1(n4603), .C2(n3482), .A(n3481), .B(n3480), .ZN(U3281)
         );
  INV_X1 U4349 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n3946) );
  NAND2_X1 U4350 ( .A1(n4463), .A2(n3562), .ZN(n3483) );
  OAI21_X1 U4351 ( .B1(U4043), .B2(n3946), .A(n3483), .ZN(U3577) );
  XNOR2_X1 U4352 ( .A(n3486), .B(n3485), .ZN(n3487) );
  XNOR2_X1 U4353 ( .A(n3484), .B(n3487), .ZN(n3491) );
  OAI22_X1 U4354 ( .A1(n4137), .A2(n4648), .B1(n3569), .B2(n4135), .ZN(n3489)
         );
  NAND2_X1 U4355 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n3552) );
  AOI211_X1 U4356 ( .C1(n3579), .C2(n3845), .A(n3489), .B(n3488), .ZN(n3490)
         );
  OAI21_X1 U4357 ( .B1(n3491), .B2(n4175), .A(n3490), .ZN(U3233) );
  INV_X1 U4358 ( .A(n4286), .ZN(n3507) );
  XNOR2_X1 U4359 ( .A(n3492), .B(n3507), .ZN(n3497) );
  NOR2_X1 U4360 ( .A1(n3754), .A2(n4645), .ZN(n3493) );
  AOI21_X1 U4361 ( .B1(n3753), .B2(n4630), .A(n3493), .ZN(n3494) );
  OAI21_X1 U4362 ( .B1(n3495), .B2(n4908), .A(n3494), .ZN(n3496) );
  AOI21_X1 U4363 ( .B1(n3497), .B2(n4906), .A(n3496), .ZN(n4979) );
  OAI211_X1 U4364 ( .C1(n2133), .C2(n3754), .A(n3498), .B(n4972), .ZN(n4978)
         );
  INV_X1 U4365 ( .A(n4978), .ZN(n3501) );
  INV_X1 U4366 ( .A(n3757), .ZN(n3499) );
  OAI22_X1 U4367 ( .A1(n4668), .A2(n4037), .B1(n3499), .B2(n4665), .ZN(n3500)
         );
  AOI21_X1 U4368 ( .B1(n3501), .B2(n4618), .A(n3500), .ZN(n3510) );
  OR2_X1 U4369 ( .A1(n3328), .A2(n3753), .ZN(n3505) );
  NAND2_X1 U4370 ( .A1(n3328), .A2(n3753), .ZN(n3503) );
  NAND2_X1 U4371 ( .A1(n3503), .A2(n3502), .ZN(n3504) );
  AND2_X1 U4372 ( .A1(n3505), .A2(n3504), .ZN(n3506) );
  NAND2_X1 U4373 ( .A1(n3506), .A2(n4286), .ZN(n4976) );
  INV_X1 U4374 ( .A(n3506), .ZN(n3508) );
  NAND2_X1 U4375 ( .A1(n3508), .A2(n3507), .ZN(n4974) );
  NAND3_X1 U4376 ( .A1(n4976), .A2(n4640), .A3(n4974), .ZN(n3509) );
  OAI211_X1 U4377 ( .C1(n4979), .C2(n4643), .A(n3510), .B(n3509), .ZN(U3283)
         );
  INV_X1 U4378 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3513) );
  INV_X1 U4379 ( .A(n3511), .ZN(n3512) );
  OAI22_X1 U4380 ( .A1(n4668), .A2(n3513), .B1(n3512), .B2(n4665), .ZN(n3516)
         );
  NOR2_X1 U4381 ( .A1(n3514), .A2(n4603), .ZN(n3515) );
  AOI211_X1 U4382 ( .C1(n3517), .C2(n4896), .A(n3516), .B(n3515), .ZN(n3518)
         );
  OAI21_X1 U4383 ( .B1(n4643), .B2(n3519), .A(n3518), .ZN(U3284) );
  NAND2_X1 U4384 ( .A1(n4207), .A2(n4212), .ZN(n4255) );
  XOR2_X1 U4385 ( .A(n4255), .B(n3520), .Z(n3523) );
  AOI22_X1 U4386 ( .A1(n4343), .A2(n4630), .B1(n3525), .B2(n4568), .ZN(n3521)
         );
  OAI21_X1 U4387 ( .B1(n3727), .B2(n4908), .A(n3521), .ZN(n3522) );
  AOI21_X1 U4388 ( .B1(n3523), .B2(n4906), .A(n3522), .ZN(n3543) );
  XOR2_X1 U4389 ( .A(n4255), .B(n3524), .Z(n3544) );
  INV_X1 U4390 ( .A(n3544), .ZN(n3532) );
  AND2_X1 U4391 ( .A1(n3526), .A2(n3525), .ZN(n3527) );
  NOR2_X1 U4392 ( .A1(n3577), .A2(n3527), .ZN(n3566) );
  INV_X1 U4393 ( .A(n3566), .ZN(n3530) );
  AOI22_X1 U4394 ( .A1(n4643), .A2(REG2_REG_10__SCAN_IN), .B1(n3528), .B2(
        n4912), .ZN(n3529) );
  OAI21_X1 U4395 ( .B1(n3530), .B2(n4600), .A(n3529), .ZN(n3531) );
  AOI21_X1 U4396 ( .B1(n3532), .B2(n4640), .A(n3531), .ZN(n3533) );
  OAI21_X1 U4397 ( .B1(n3543), .B2(n4643), .A(n3533), .ZN(U3280) );
  INV_X1 U4398 ( .A(n3534), .ZN(n3542) );
  INV_X1 U4399 ( .A(n3535), .ZN(n3538) );
  AOI22_X1 U4400 ( .A1(n4643), .A2(REG2_REG_8__SCAN_IN), .B1(n3536), .B2(n4912), .ZN(n3537) );
  OAI21_X1 U4401 ( .B1(n3538), .B2(n4600), .A(n3537), .ZN(n3539) );
  AOI21_X1 U4402 ( .B1(n3540), .B2(n4640), .A(n3539), .ZN(n3541) );
  OAI21_X1 U4403 ( .B1(n3542), .B2(n4643), .A(n3541), .ZN(U3282) );
  OAI21_X1 U4404 ( .B1(n4967), .B2(n3544), .A(n3543), .ZN(n3565) );
  INV_X1 U4405 ( .A(n3565), .ZN(n3546) );
  AOI22_X1 U4406 ( .A1(n3566), .A2(n4743), .B1(REG0_REG_10__SCAN_IN), .B2(
        n4980), .ZN(n3545) );
  OAI21_X1 U4407 ( .B1(n3546), .B2(n4980), .A(n3545), .ZN(U3487) );
  INV_X1 U4408 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4034) );
  MUX2_X1 U4409 ( .A(REG2_REG_11__SCAN_IN), .B(n4034), .S(n3640), .Z(n3550) );
  AOI211_X1 U4410 ( .C1(n3549), .C2(n3550), .A(n4878), .B(n3636), .ZN(n3554)
         );
  NAND2_X1 U4411 ( .A1(n4881), .A2(ADDR_REG_11__SCAN_IN), .ZN(n3551) );
  OAI211_X1 U4412 ( .C1(n4892), .C2(n3640), .A(n3552), .B(n3551), .ZN(n3553)
         );
  NOR2_X1 U4413 ( .A1(n3554), .A2(n3553), .ZN(n3561) );
  NAND2_X1 U4414 ( .A1(n3557), .A2(n2421), .ZN(n3559) );
  XNOR2_X1 U4415 ( .A(n3640), .B(REG1_REG_11__SCAN_IN), .ZN(n3558) );
  NAND2_X1 U4416 ( .A1(n3559), .A2(n3558), .ZN(n3643) );
  OAI211_X1 U4417 ( .C1(n3559), .C2(n3558), .A(n3643), .B(n4873), .ZN(n3560)
         );
  NAND2_X1 U4418 ( .A1(n3561), .A2(n3560), .ZN(U3251) );
  INV_X1 U4419 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n3987) );
  NAND2_X1 U4420 ( .A1(n4240), .A2(n3562), .ZN(n3563) );
  OAI21_X1 U4421 ( .B1(U4043), .B2(n3987), .A(n3563), .ZN(U3579) );
  INV_X1 U4422 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4059) );
  NAND2_X1 U4423 ( .A1(n3565), .A2(n4994), .ZN(n3568) );
  NAND2_X1 U4424 ( .A1(n3566), .A2(n4676), .ZN(n3567) );
  OAI211_X1 U4425 ( .C1(n4994), .C2(n4059), .A(n3568), .B(n3567), .ZN(U3528)
         );
  XOR2_X1 U4426 ( .A(n3586), .B(n4273), .Z(n3575) );
  OR2_X1 U4427 ( .A1(n3571), .A2(n4273), .ZN(n3596) );
  INV_X1 U4428 ( .A(n3596), .ZN(n3570) );
  AOI21_X1 U4429 ( .B1(n4273), .B2(n3571), .A(n3570), .ZN(n3576) );
  NOR2_X1 U4430 ( .A1(n3576), .A2(n4905), .ZN(n3572) );
  AOI211_X1 U4431 ( .C1(n4660), .C2(n3624), .A(n3573), .B(n3572), .ZN(n3574)
         );
  OAI21_X1 U4432 ( .B1(n4655), .B2(n3575), .A(n3574), .ZN(n3629) );
  INV_X1 U4433 ( .A(n3629), .ZN(n3583) );
  INV_X1 U4434 ( .A(n3576), .ZN(n3630) );
  OR2_X1 U4435 ( .A1(n3599), .A2(n3578), .ZN(n3635) );
  AOI22_X1 U4436 ( .A1(n4643), .A2(REG2_REG_11__SCAN_IN), .B1(n3579), .B2(
        n4912), .ZN(n3580) );
  OAI21_X1 U4437 ( .B1(n3635), .B2(n4600), .A(n3580), .ZN(n3581) );
  AOI21_X1 U4438 ( .B1(n3630), .B2(n4913), .A(n3581), .ZN(n3582) );
  OAI21_X1 U4439 ( .B1(n3583), .B2(n4643), .A(n3582), .ZN(U3279) );
  INV_X1 U4440 ( .A(n3584), .ZN(n3585) );
  OR2_X1 U4441 ( .A1(n3586), .A2(n3585), .ZN(n3588) );
  NAND2_X1 U4442 ( .A1(n3588), .A2(n3587), .ZN(n4652) );
  NAND2_X1 U4443 ( .A1(n4651), .A2(n4649), .ZN(n4279) );
  XNOR2_X1 U4444 ( .A(n4652), .B(n4279), .ZN(n3594) );
  NAND2_X1 U4445 ( .A1(n3589), .A2(n4660), .ZN(n3592) );
  NAND2_X1 U4446 ( .A1(n3590), .A2(n4568), .ZN(n3591) );
  OAI211_X1 U4447 ( .C1(n3727), .C2(n4647), .A(n3592), .B(n3591), .ZN(n3593)
         );
  AOI21_X1 U4448 ( .B1(n3594), .B2(n4906), .A(n3593), .ZN(n3668) );
  NAND2_X1 U4449 ( .A1(n3596), .A2(n3595), .ZN(n3597) );
  XNOR2_X1 U4450 ( .A(n3597), .B(n4279), .ZN(n3666) );
  OR2_X1 U4451 ( .A1(n3599), .A2(n3730), .ZN(n3600) );
  NAND2_X1 U4452 ( .A1(n3598), .A2(n3600), .ZN(n3674) );
  AOI22_X1 U4453 ( .A1(n4643), .A2(REG2_REG_12__SCAN_IN), .B1(n3733), .B2(
        n4912), .ZN(n3601) );
  OAI21_X1 U4454 ( .B1(n3674), .B2(n4600), .A(n3601), .ZN(n3602) );
  AOI21_X1 U4455 ( .B1(n3666), .B2(n4640), .A(n3602), .ZN(n3603) );
  OAI21_X1 U4456 ( .B1(n3668), .B2(n4643), .A(n3603), .ZN(U3278) );
  XNOR2_X1 U4457 ( .A(n3604), .B(n3613), .ZN(n3607) );
  OAI22_X1 U4458 ( .A1(n3728), .A2(n4647), .B1(n3684), .B2(n4645), .ZN(n3605)
         );
  AOI21_X1 U4459 ( .B1(n4660), .B2(n3694), .A(n3605), .ZN(n3606) );
  OAI21_X1 U4460 ( .B1(n3607), .B2(n4655), .A(n3606), .ZN(n3660) );
  INV_X1 U4461 ( .A(n3660), .ZN(n3621) );
  NOR2_X1 U4462 ( .A1(n4644), .A2(n3608), .ZN(n3611) );
  NOR2_X1 U4463 ( .A1(n3611), .A2(n3609), .ZN(n3614) );
  OR2_X1 U4464 ( .A1(n3611), .A2(n3610), .ZN(n3612) );
  OAI21_X1 U4465 ( .B1(n3614), .B2(n3613), .A(n3612), .ZN(n3661) );
  NAND2_X1 U4466 ( .A1(n4664), .A2(n3615), .ZN(n3616) );
  NAND2_X1 U4467 ( .A1(n3651), .A2(n3616), .ZN(n3665) );
  INV_X1 U4468 ( .A(n3617), .ZN(n3687) );
  AOI22_X1 U4469 ( .A1(n4643), .A2(REG2_REG_14__SCAN_IN), .B1(n3687), .B2(
        n4912), .ZN(n3618) );
  OAI21_X1 U4470 ( .B1(n3665), .B2(n4600), .A(n3618), .ZN(n3619) );
  AOI21_X1 U4471 ( .B1(n3661), .B2(n4640), .A(n3619), .ZN(n3620) );
  OAI21_X1 U4472 ( .B1(n4643), .B2(n3621), .A(n3620), .ZN(U3276) );
  XNOR2_X1 U4473 ( .A(n3676), .B(n3675), .ZN(n3623) );
  XNOR2_X1 U4474 ( .A(n3622), .B(n3623), .ZN(n3628) );
  AOI22_X1 U4475 ( .A1(n4167), .A2(n3624), .B1(n4166), .B2(n4659), .ZN(n3627)
         );
  NOR2_X1 U4476 ( .A1(n3853), .A2(STATE_REG_SCAN_IN), .ZN(n4833) );
  NOR2_X1 U4477 ( .A1(n4169), .A2(n4666), .ZN(n3625) );
  AOI211_X1 U4478 ( .C1(n4662), .C2(n4171), .A(n4833), .B(n3625), .ZN(n3626)
         );
  OAI211_X1 U4479 ( .C1(n3628), .C2(n4175), .A(n3627), .B(n3626), .ZN(U3231)
         );
  INV_X1 U4480 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3631) );
  AOI21_X1 U4481 ( .B1(n4963), .B2(n3630), .A(n3629), .ZN(n3633) );
  MUX2_X1 U4482 ( .A(n3631), .B(n3633), .S(n4777), .Z(n3632) );
  OAI21_X1 U4483 ( .B1(n3635), .B2(n4787), .A(n3632), .ZN(U3489) );
  INV_X1 U4484 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3641) );
  MUX2_X1 U4485 ( .A(n3641), .B(n3633), .S(n4994), .Z(n3634) );
  OAI21_X1 U4486 ( .B1(n4738), .B2(n3635), .A(n3634), .ZN(U3529) );
  INV_X1 U4487 ( .A(n3640), .ZN(n4795) );
  XNOR2_X1 U4488 ( .A(n4376), .B(REG2_REG_12__SCAN_IN), .ZN(n3647) );
  INV_X1 U4489 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n3637) );
  NAND2_X1 U4490 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n3729) );
  OAI21_X1 U4491 ( .B1(n3638), .B2(n3637), .A(n3729), .ZN(n3639) );
  AOI21_X1 U4492 ( .B1(n4794), .B2(n4849), .A(n3639), .ZN(n3646) );
  NAND2_X1 U4493 ( .A1(n3643), .A2(n3642), .ZN(n4392) );
  INV_X1 U4494 ( .A(n4794), .ZN(n4377) );
  OAI211_X1 U4495 ( .C1(n3644), .C2(REG1_REG_12__SCAN_IN), .A(n4394), .B(n4873), .ZN(n3645) );
  OAI211_X1 U4496 ( .C1(n3647), .C2(n4878), .A(n3646), .B(n3645), .ZN(U3252)
         );
  AND2_X1 U4497 ( .A1(n3648), .A2(n2430), .ZN(n3649) );
  XNOR2_X1 U4498 ( .A(n3649), .B(n2428), .ZN(n4732) );
  XNOR2_X1 U4499 ( .A(n3651), .B(n3650), .ZN(n4730) );
  INV_X1 U4500 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3652) );
  OAI22_X1 U4501 ( .A1(n4668), .A2(n3652), .B1(n4168), .B2(n4665), .ZN(n3653)
         );
  AOI21_X1 U4502 ( .B1(n4730), .B2(n4896), .A(n3653), .ZN(n3659) );
  INV_X1 U4503 ( .A(n4629), .ZN(n3657) );
  OAI211_X1 U4504 ( .C1(n2429), .C2(n2428), .A(n4906), .B(n3654), .ZN(n3656)
         );
  AOI22_X1 U4505 ( .A1(n4659), .A2(n4630), .B1(n4568), .B2(n4172), .ZN(n3655)
         );
  OAI211_X1 U4506 ( .C1(n3657), .C2(n4908), .A(n3656), .B(n3655), .ZN(n4729)
         );
  NAND2_X1 U4507 ( .A1(n4729), .A2(n4668), .ZN(n3658) );
  OAI211_X1 U4508 ( .C1(n4732), .C2(n4603), .A(n3659), .B(n3658), .ZN(U3275)
         );
  AOI21_X1 U4509 ( .B1(n3661), .B2(n4975), .A(n3660), .ZN(n3663) );
  INV_X1 U4510 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4843) );
  MUX2_X1 U4511 ( .A(n3663), .B(n4843), .S(n4991), .Z(n3662) );
  OAI21_X1 U4512 ( .B1(n4738), .B2(n3665), .A(n3662), .ZN(U3532) );
  INV_X1 U4513 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4057) );
  MUX2_X1 U4514 ( .A(n3663), .B(n4057), .S(n4980), .Z(n3664) );
  OAI21_X1 U4515 ( .B1(n3665), .B2(n4787), .A(n3664), .ZN(U3495) );
  NAND2_X1 U4516 ( .A1(n3666), .A2(n4975), .ZN(n3667) );
  NAND2_X1 U4517 ( .A1(n3668), .A2(n3667), .ZN(n3671) );
  MUX2_X1 U4518 ( .A(REG0_REG_12__SCAN_IN), .B(n3671), .S(n4777), .Z(n3669) );
  INV_X1 U4519 ( .A(n3669), .ZN(n3670) );
  OAI21_X1 U4520 ( .B1(n3674), .B2(n4787), .A(n3670), .ZN(U3491) );
  MUX2_X1 U4521 ( .A(REG1_REG_12__SCAN_IN), .B(n3671), .S(n4994), .Z(n3672) );
  INV_X1 U4522 ( .A(n3672), .ZN(n3673) );
  OAI21_X1 U4523 ( .B1(n4738), .B2(n3674), .A(n3673), .ZN(U3530) );
  INV_X1 U4524 ( .A(n3622), .ZN(n3679) );
  INV_X1 U4525 ( .A(n3676), .ZN(n3678) );
  AOI21_X1 U4526 ( .B1(n3622), .B2(n3676), .A(n3675), .ZN(n3677) );
  AOI21_X1 U4527 ( .B1(n3679), .B2(n3678), .A(n3677), .ZN(n3683) );
  NAND2_X1 U4528 ( .A1(n3681), .A2(n3680), .ZN(n3682) );
  XNOR2_X1 U4529 ( .A(n3683), .B(n3682), .ZN(n3689) );
  OAI22_X1 U4530 ( .A1(n4137), .A2(n3805), .B1(n3728), .B2(n4135), .ZN(n3686)
         );
  NAND2_X1 U4531 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n4850) );
  OAI21_X1 U4532 ( .B1(n3090), .B2(n3684), .A(n4850), .ZN(n3685) );
  AOI211_X1 U4533 ( .C1(n3687), .C2(n3845), .A(n3686), .B(n3685), .ZN(n3688)
         );
  OAI21_X1 U4534 ( .B1(n3689), .B2(n4175), .A(n3688), .ZN(U3212) );
  OAI21_X1 U4535 ( .B1(n3691), .B2(n2700), .A(n3690), .ZN(n4728) );
  OAI211_X1 U4536 ( .C1(n3693), .C2(n4288), .A(n3692), .B(n4906), .ZN(n3696)
         );
  AOI22_X1 U4537 ( .A1(n3694), .A2(n4630), .B1(n3700), .B2(n4568), .ZN(n3695)
         );
  OAI211_X1 U4538 ( .C1(n4605), .C2(n4908), .A(n3696), .B(n3695), .ZN(n4725)
         );
  INV_X1 U4539 ( .A(n3697), .ZN(n3699) );
  INV_X1 U4540 ( .A(n3698), .ZN(n4633) );
  AOI21_X1 U4541 ( .B1(n3700), .B2(n3699), .A(n4633), .ZN(n4726) );
  INV_X1 U4542 ( .A(n4726), .ZN(n3702) );
  AOI22_X1 U4543 ( .A1(n4643), .A2(REG2_REG_16__SCAN_IN), .B1(n3809), .B2(
        n4912), .ZN(n3701) );
  OAI21_X1 U4544 ( .B1(n3702), .B2(n4600), .A(n3701), .ZN(n3703) );
  AOI21_X1 U4545 ( .B1(n4725), .B2(n4668), .A(n3703), .ZN(n3704) );
  OAI21_X1 U4546 ( .B1(n4728), .B2(n4603), .A(n3704), .ZN(U3274) );
  INV_X1 U4547 ( .A(n3705), .ZN(n3770) );
  AOI21_X1 U4548 ( .B1(n3707), .B2(n3706), .A(n3770), .ZN(n3712) );
  AOI22_X1 U4549 ( .A1(n4171), .A2(n4542), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3709) );
  NAND2_X1 U4550 ( .A1(n4541), .A2(n3845), .ZN(n3708) );
  OAI211_X1 U4551 ( .C1(n4570), .C2(n4135), .A(n3709), .B(n3708), .ZN(n3710)
         );
  AOI21_X1 U4552 ( .B1(n4340), .B2(n4166), .A(n3710), .ZN(n3711) );
  OAI21_X1 U4553 ( .B1(n3712), .B2(n4175), .A(n3711), .ZN(U3232) );
  NAND2_X1 U4554 ( .A1(n3713), .A2(n4140), .ZN(n3723) );
  AOI21_X1 U4555 ( .B1(n3264), .B2(n3715), .A(n3714), .ZN(n3722) );
  OAI22_X1 U4556 ( .A1(n4137), .A2(n3716), .B1(n4136), .B2(n4135), .ZN(n3719)
         );
  NAND2_X1 U4557 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4821) );
  OAI21_X1 U4558 ( .B1(n3090), .B2(n3717), .A(n4821), .ZN(n3718) );
  AOI211_X1 U4559 ( .C1(n3720), .C2(n3845), .A(n3719), .B(n3718), .ZN(n3721)
         );
  OAI21_X1 U4560 ( .B1(n3723), .B2(n3722), .A(n3721), .ZN(U3227) );
  NOR2_X1 U4561 ( .A1(n2181), .A2(n3724), .ZN(n3725) );
  XNOR2_X1 U4562 ( .A(n3726), .B(n3725), .ZN(n3735) );
  OAI22_X1 U4563 ( .A1(n4137), .A2(n3728), .B1(n3727), .B2(n4135), .ZN(n3732)
         );
  OAI21_X1 U4564 ( .B1(n3090), .B2(n3730), .A(n3729), .ZN(n3731) );
  AOI211_X1 U4565 ( .C1(n3733), .C2(n3845), .A(n3732), .B(n3731), .ZN(n3734)
         );
  OAI21_X1 U4566 ( .B1(n3735), .B2(n4175), .A(n3734), .ZN(U3221) );
  INV_X1 U4567 ( .A(n3736), .ZN(n3741) );
  OAI22_X1 U4568 ( .A1(n3737), .A2(n4665), .B1(n4085), .B2(n4668), .ZN(n3740)
         );
  NOR2_X1 U4569 ( .A1(n3738), .A2(n4643), .ZN(n3739) );
  OAI21_X1 U4570 ( .B1(n3743), .B2(n4603), .A(n3742), .ZN(U3262) );
  XOR2_X1 U4571 ( .A(n3745), .B(n3744), .Z(n4356) );
  NAND2_X1 U4572 ( .A1(n4356), .A2(n4140), .ZN(n3749) );
  AOI22_X1 U4573 ( .A1(n4171), .A2(n3747), .B1(REG3_REG_0__SCAN_IN), .B2(n3746), .ZN(n3748) );
  OAI211_X1 U4574 ( .C1(n2885), .C2(n4137), .A(n3749), .B(n3748), .ZN(U3229)
         );
  OAI211_X1 U4575 ( .C1(n3752), .C2(n3751), .A(n3750), .B(n4140), .ZN(n3760)
         );
  AOI22_X1 U4576 ( .A1(n4167), .A2(n3753), .B1(n4166), .B2(n4344), .ZN(n3759)
         );
  NOR2_X1 U4577 ( .A1(n3090), .A2(n3754), .ZN(n3755) );
  AOI211_X1 U4578 ( .C1(n3845), .C2(n3757), .A(n3756), .B(n3755), .ZN(n3758)
         );
  NAND3_X1 U4579 ( .A1(n3760), .A2(n3759), .A3(n3758), .ZN(U3210) );
  XNOR2_X1 U4580 ( .A(n3762), .B(n3761), .ZN(n3767) );
  OAI22_X1 U4581 ( .A1(n3090), .A2(n4447), .B1(STATE_REG_SCAN_IN), .B2(n4072), 
        .ZN(n3763) );
  AOI21_X1 U4582 ( .B1(n4448), .B2(n3845), .A(n3763), .ZN(n3764) );
  OAI21_X1 U4583 ( .B1(n4437), .B2(n4135), .A(n3764), .ZN(n3765) );
  AOI21_X1 U4584 ( .B1(n4444), .B2(n4166), .A(n3765), .ZN(n3766) );
  OAI21_X1 U4585 ( .B1(n3767), .B2(n4175), .A(n3766), .ZN(U3211) );
  OAI21_X1 U4586 ( .B1(n3770), .B2(n3769), .A(n3768), .ZN(n3772) );
  NAND3_X1 U4587 ( .A1(n3772), .A2(n4140), .A3(n3771), .ZN(n3777) );
  OAI22_X1 U4588 ( .A1(n3090), .A2(n4523), .B1(STATE_REG_SCAN_IN), .B2(n3773), 
        .ZN(n3775) );
  NOR2_X1 U4589 ( .A1(n4516), .A2(n4135), .ZN(n3774) );
  AOI211_X1 U4590 ( .C1(n3845), .C2(n4525), .A(n3775), .B(n3774), .ZN(n3776)
         );
  OAI211_X1 U4591 ( .C1(n4480), .C2(n4137), .A(n3777), .B(n3776), .ZN(U3213)
         );
  XOR2_X1 U4592 ( .A(n3779), .B(n3778), .Z(n3783) );
  AOI22_X1 U4593 ( .A1(n4593), .A2(n4166), .B1(n4167), .B2(n3820), .ZN(n3782)
         );
  NOR2_X1 U4594 ( .A1(n4046), .A2(STATE_REG_SCAN_IN), .ZN(n4810) );
  NOR2_X1 U4595 ( .A1(n3090), .A2(n4597), .ZN(n3780) );
  AOI211_X1 U4596 ( .C1(n3845), .C2(n4598), .A(n4810), .B(n3780), .ZN(n3781)
         );
  OAI211_X1 U4597 ( .C1(n3783), .C2(n4175), .A(n3782), .B(n3781), .ZN(U3216)
         );
  XNOR2_X1 U4598 ( .A(n3786), .B(n3785), .ZN(n3787) );
  XNOR2_X1 U4599 ( .A(n3784), .B(n3787), .ZN(n3791) );
  OAI22_X1 U4600 ( .A1(n3090), .A2(n4557), .B1(STATE_REG_SCAN_IN), .B2(n4077), 
        .ZN(n3789) );
  OAI22_X1 U4601 ( .A1(n4516), .A2(n4137), .B1(n4169), .B2(n4559), .ZN(n3788)
         );
  AOI211_X1 U4602 ( .C1(n4167), .C2(n4593), .A(n3789), .B(n3788), .ZN(n3790)
         );
  OAI21_X1 U4603 ( .B1(n3791), .B2(n4175), .A(n3790), .ZN(U3220) );
  INV_X1 U4604 ( .A(n3793), .ZN(n3794) );
  NOR2_X1 U4605 ( .A1(n3795), .A2(n3794), .ZN(n3796) );
  XNOR2_X1 U4606 ( .A(n3792), .B(n3796), .ZN(n3801) );
  OAI22_X1 U4607 ( .A1(n3090), .A2(n4487), .B1(STATE_REG_SCAN_IN), .B2(n4090), 
        .ZN(n3797) );
  AOI21_X1 U4608 ( .B1(n4489), .B2(n3845), .A(n3797), .ZN(n3798) );
  OAI21_X1 U4609 ( .B1(n4480), .B2(n4135), .A(n3798), .ZN(n3799) );
  AOI21_X1 U4610 ( .B1(n4482), .B2(n4166), .A(n3799), .ZN(n3800) );
  OAI21_X1 U4611 ( .B1(n3801), .B2(n4175), .A(n3800), .ZN(U3222) );
  NOR2_X1 U4612 ( .A1(n3802), .A2(n3803), .ZN(n4163) );
  NAND2_X1 U4613 ( .A1(n3802), .A2(n3803), .ZN(n4161) );
  OAI21_X1 U4614 ( .B1(n4163), .B2(n4164), .A(n4161), .ZN(n3804) );
  XNOR2_X1 U4615 ( .A(n3815), .B(n3814), .ZN(n3812) );
  XNOR2_X1 U4616 ( .A(n3804), .B(n3812), .ZN(n3811) );
  OAI22_X1 U4617 ( .A1(n4137), .A2(n4605), .B1(n3805), .B2(n4135), .ZN(n3808)
         );
  NAND2_X1 U4618 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4864) );
  OAI21_X1 U4619 ( .B1(n3090), .B2(n3806), .A(n4864), .ZN(n3807) );
  AOI211_X1 U4620 ( .C1(n3809), .C2(n3845), .A(n3808), .B(n3807), .ZN(n3810)
         );
  OAI21_X1 U4621 ( .B1(n3811), .B2(n4175), .A(n3810), .ZN(U3223) );
  AOI211_X1 U4622 ( .C1(n4164), .C2(n4161), .A(n3812), .B(n4163), .ZN(n3813)
         );
  AOI21_X1 U4623 ( .B1(n3815), .B2(n3814), .A(n3813), .ZN(n3819) );
  XOR2_X1 U4624 ( .A(n3817), .B(n3816), .Z(n3818) );
  XNOR2_X1 U4625 ( .A(n3819), .B(n3818), .ZN(n3826) );
  AOI22_X1 U4626 ( .A1(n4166), .A2(n3820), .B1(n4167), .B2(n4629), .ZN(n3825)
         );
  NOR2_X1 U4627 ( .A1(n3821), .A2(STATE_REG_SCAN_IN), .ZN(n4390) );
  NOR2_X1 U4628 ( .A1(n4169), .A2(n4634), .ZN(n3822) );
  AOI211_X1 U4629 ( .C1(n3823), .C2(n4171), .A(n4390), .B(n3822), .ZN(n3824)
         );
  OAI211_X1 U4630 ( .C1(n3826), .C2(n4175), .A(n3825), .B(n3824), .ZN(U3225)
         );
  NAND2_X1 U4631 ( .A1(n3827), .A2(n3828), .ZN(n3829) );
  XOR2_X1 U4632 ( .A(n3830), .B(n3829), .Z(n3836) );
  NAND2_X1 U4633 ( .A1(n4340), .A2(n4167), .ZN(n3833) );
  AOI22_X1 U4634 ( .A1(n4171), .A2(n3831), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3832) );
  OAI211_X1 U4635 ( .C1(n4169), .C2(n4504), .A(n3833), .B(n3832), .ZN(n3834)
         );
  AOI21_X1 U4636 ( .B1(n4498), .B2(n4166), .A(n3834), .ZN(n3835) );
  OAI21_X1 U4637 ( .B1(n3836), .B2(n4175), .A(n3835), .ZN(U3226) );
  INV_X1 U4638 ( .A(n3837), .ZN(n3842) );
  AOI21_X1 U4639 ( .B1(n3841), .B2(n3839), .A(n3838), .ZN(n3840) );
  AOI21_X1 U4640 ( .B1(n3842), .B2(n3841), .A(n3840), .ZN(n3849) );
  AOI22_X1 U4641 ( .A1(n4534), .A2(n4166), .B1(n4167), .B2(n4610), .ZN(n3848)
         );
  INV_X1 U4642 ( .A(n4579), .ZN(n3846) );
  OAI22_X1 U4643 ( .A1(n3090), .A2(n3843), .B1(STATE_REG_SCAN_IN), .B2(n2237), 
        .ZN(n3844) );
  AOI21_X1 U4644 ( .B1(n3846), .B2(n3845), .A(n3844), .ZN(n3847) );
  OAI211_X1 U4645 ( .C1(n3849), .C2(n4175), .A(n3848), .B(n3847), .ZN(U3230)
         );
  INV_X1 U4646 ( .A(keyinput108), .ZN(n4129) );
  INV_X1 U4647 ( .A(IR_REG_13__SCAN_IN), .ZN(n3975) );
  NAND4_X1 U4648 ( .A1(n3852), .A2(n3975), .A3(n3851), .A4(n3850), .ZN(n3860)
         );
  NAND4_X1 U4649 ( .A1(n2846), .A2(n3854), .A3(n3853), .A4(REG3_REG_8__SCAN_IN), .ZN(n3859) );
  INV_X1 U4650 ( .A(REG3_REG_2__SCAN_IN), .ZN(n4133) );
  INV_X1 U4651 ( .A(DATAI_0_), .ZN(n3855) );
  NAND4_X1 U4652 ( .A1(n4133), .A2(n3855), .A3(IR_REG_19__SCAN_IN), .A4(
        REG3_REG_0__SCAN_IN), .ZN(n3858) );
  NOR4_X1 U4653 ( .A1(REG2_REG_29__SCAN_IN), .A2(n4072), .A3(n4077), .A4(n2237), .ZN(n3856) );
  NAND4_X1 U4654 ( .A1(ADDR_REG_0__SCAN_IN), .A2(IR_REG_30__SCAN_IN), .A3(
        n3856), .A4(REG1_REG_3__SCAN_IN), .ZN(n3857) );
  NOR4_X1 U4655 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3863)
         );
  NOR4_X1 U4656 ( .A1(REG2_REG_19__SCAN_IN), .A2(REG3_REG_1__SCAN_IN), .A3(
        ADDR_REG_3__SCAN_IN), .A4(DATAO_REG_12__SCAN_IN), .ZN(n3862) );
  NOR4_X1 U4657 ( .A1(DATAO_REG_13__SCAN_IN), .A2(DATAO_REG_16__SCAN_IN), .A3(
        DATAO_REG_19__SCAN_IN), .A4(DATAO_REG_20__SCAN_IN), .ZN(n3861) );
  NAND4_X1 U4658 ( .A1(n3863), .A2(n3862), .A3(n3861), .A4(D_REG_24__SCAN_IN), 
        .ZN(n3873) );
  INV_X1 U4659 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4060) );
  INV_X1 U4660 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4055) );
  NOR4_X1 U4661 ( .A1(n2611), .A2(n4060), .A3(n4054), .A4(n4055), .ZN(n3868)
         );
  INV_X1 U4662 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3864) );
  INV_X1 U4663 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4021) );
  INV_X1 U4664 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4973) );
  NOR4_X1 U4665 ( .A1(IR_REG_15__SCAN_IN), .A2(n3864), .A3(n4021), .A4(n4973), 
        .ZN(n3867) );
  NOR4_X1 U4666 ( .A1(IR_REG_11__SCAN_IN), .A2(REG0_REG_19__SCAN_IN), .A3(
        REG0_REG_16__SCAN_IN), .A4(DATAI_9_), .ZN(n3866) );
  NOR4_X1 U4667 ( .A1(IR_REG_7__SCAN_IN), .A2(REG2_REG_14__SCAN_IN), .A3(n4057), .A4(n4059), .ZN(n3865) );
  NAND4_X1 U4668 ( .A1(n3868), .A2(n3867), .A3(n3866), .A4(n3865), .ZN(n3872)
         );
  INV_X1 U4669 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4867) );
  NAND4_X1 U4670 ( .A1(REG3_REG_18__SCAN_IN), .A2(REG2_REG_24__SCAN_IN), .A3(
        n4867), .A4(n4578), .ZN(n3871) );
  NAND4_X1 U4671 ( .A1(n4000), .A2(n3869), .A3(DATAO_REG_6__SCAN_IN), .A4(
        DATAO_REG_10__SCAN_IN), .ZN(n3870) );
  OR4_X1 U4672 ( .A1(n3873), .A2(n3872), .A3(n3871), .A4(n3870), .ZN(n3876) );
  NAND3_X1 U4673 ( .A1(n3874), .A2(D_REG_17__SCAN_IN), .A3(DATAI_22_), .ZN(
        n3875) );
  NOR2_X1 U4674 ( .A1(n3876), .A2(n3875), .ZN(n3888) );
  INV_X1 U4675 ( .A(DATAI_12_), .ZN(n3960) );
  NOR4_X1 U4676 ( .A1(DATAI_11_), .A2(n3960), .A3(n4927), .A4(n3966), .ZN(
        n3887) );
  INV_X1 U4677 ( .A(DATAI_20_), .ZN(n3986) );
  NAND4_X1 U4678 ( .A1(D_REG_26__SCAN_IN), .A2(DATAO_REG_24__SCAN_IN), .A3(
        DATAO_REG_29__SCAN_IN), .A4(n3994), .ZN(n3877) );
  NOR3_X1 U4679 ( .A1(DATAI_23_), .A2(n3986), .A3(n3877), .ZN(n3886) );
  NOR4_X1 U4680 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4667), .A3(n3652), .A4(n4099), 
        .ZN(n3881) );
  INV_X1 U4681 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4101) );
  INV_X1 U4682 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n4103) );
  NOR4_X1 U4683 ( .A1(n3637), .A2(n4101), .A3(n4103), .A4(REG1_REG_4__SCAN_IN), 
        .ZN(n3880) );
  NOR4_X1 U4684 ( .A1(REG1_REG_2__SCAN_IN), .A2(n4989), .A3(n4034), .A4(n3168), 
        .ZN(n3879) );
  INV_X1 U4685 ( .A(REG2_REG_1__SCAN_IN), .ZN(n4031) );
  NOR4_X1 U4686 ( .A1(n4036), .A2(n4037), .A3(n4030), .A4(n4031), .ZN(n3878)
         );
  NAND4_X1 U4687 ( .A1(n3881), .A2(n3880), .A3(n3879), .A4(n3878), .ZN(n3884)
         );
  INV_X1 U4688 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4093) );
  INV_X1 U4689 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4088) );
  NOR4_X1 U4690 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG2_REG_17__SCAN_IN), .A3(
        n4093), .A4(n4088), .ZN(n3882) );
  NAND4_X1 U4691 ( .A1(REG2_REG_28__SCAN_IN), .A2(REG2_REG_27__SCAN_IN), .A3(
        n4351), .A4(n3882), .ZN(n3883) );
  NOR2_X1 U4692 ( .A1(n3884), .A2(n3883), .ZN(n3885) );
  NAND4_X1 U4693 ( .A1(n3888), .A2(n3887), .A3(n3886), .A4(n3885), .ZN(n3900)
         );
  INV_X1 U4694 ( .A(D_REG_11__SCAN_IN), .ZN(n4926) );
  INV_X1 U4695 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3906) );
  INV_X1 U4696 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4690) );
  NAND4_X1 U4697 ( .A1(DATAI_19_), .A2(DATAO_REG_3__SCAN_IN), .A3(n3906), .A4(
        n4690), .ZN(n3889) );
  NOR3_X1 U4698 ( .A1(DATAO_REG_22__SCAN_IN), .A2(n4926), .A3(n3889), .ZN(
        n3898) );
  NAND3_X1 U4699 ( .A1(IR_REG_4__SCAN_IN), .A2(DATAI_4_), .A3(
        DATAO_REG_1__SCAN_IN), .ZN(n3890) );
  OR4_X1 U4700 ( .A1(n3928), .A2(n3890), .A3(DATAO_REG_15__SCAN_IN), .A4(
        DATAO_REG_18__SCAN_IN), .ZN(n3896) );
  INV_X1 U4701 ( .A(D_REG_12__SCAN_IN), .ZN(n4925) );
  NOR4_X1 U4702 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .A3(
        REG0_REG_2__SCAN_IN), .A4(n3933), .ZN(n3893) );
  NOR4_X1 U4703 ( .A1(REG1_REG_21__SCAN_IN), .A2(REG2_REG_21__SCAN_IN), .A3(
        n4046), .A4(n4768), .ZN(n3892) );
  NOR4_X1 U4704 ( .A1(REG0_REG_25__SCAN_IN), .A2(REG1_REG_23__SCAN_IN), .A3(
        REG2_REG_22__SCAN_IN), .A4(REG1_REG_24__SCAN_IN), .ZN(n3891) );
  NAND4_X1 U4705 ( .A1(IR_REG_22__SCAN_IN), .A2(n3893), .A3(n3892), .A4(n3891), 
        .ZN(n3894) );
  OR4_X1 U4706 ( .A1(n4925), .A2(n3894), .A3(DATAI_24_), .A4(
        DATAO_REG_27__SCAN_IN), .ZN(n3895) );
  NOR4_X1 U4707 ( .A1(IR_REG_9__SCAN_IN), .A2(DATAO_REG_7__SCAN_IN), .A3(n3896), .A4(n3895), .ZN(n3897) );
  INV_X1 U4708 ( .A(REG0_REG_31__SCAN_IN), .ZN(n3909) );
  NAND4_X1 U4709 ( .A1(n3898), .A2(n3897), .A3(n3905), .A4(n3909), .ZN(n3899)
         );
  OAI21_X1 U4710 ( .B1(n3900), .B2(n3899), .A(IR_REG_21__SCAN_IN), .ZN(n3901)
         );
  INV_X1 U4711 ( .A(n3901), .ZN(n4128) );
  INV_X1 U4712 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4694) );
  AOI22_X1 U4713 ( .A1(n4698), .A2(keyinput92), .B1(keyinput46), .B2(n4694), 
        .ZN(n3902) );
  OAI221_X1 U4714 ( .B1(n4698), .B2(keyinput92), .C1(n4694), .C2(keyinput46), 
        .A(n3902), .ZN(n3913) );
  AOI22_X1 U4715 ( .A1(n4755), .A2(keyinput87), .B1(n4690), .B2(keyinput127), 
        .ZN(n3903) );
  OAI221_X1 U4716 ( .B1(n4755), .B2(keyinput87), .C1(n4690), .C2(keyinput127), 
        .A(n3903), .ZN(n3912) );
  AOI22_X1 U4717 ( .A1(n3906), .A2(keyinput17), .B1(n3905), .B2(keyinput126), 
        .ZN(n3904) );
  OAI221_X1 U4718 ( .B1(n3906), .B2(keyinput17), .C1(n3905), .C2(keyinput126), 
        .A(n3904), .ZN(n3911) );
  AOI22_X1 U4719 ( .A1(n3909), .A2(keyinput90), .B1(keyinput27), .B2(n3908), 
        .ZN(n3907) );
  OAI221_X1 U4720 ( .B1(n3909), .B2(keyinput90), .C1(n3908), .C2(keyinput27), 
        .A(n3907), .ZN(n3910) );
  NOR4_X1 U4721 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3957)
         );
  INV_X1 U4722 ( .A(DATAI_19_), .ZN(n3915) );
  AOI22_X1 U4723 ( .A1(n3916), .A2(keyinput15), .B1(n3915), .B2(keyinput103), 
        .ZN(n3914) );
  OAI221_X1 U4724 ( .B1(n3916), .B2(keyinput15), .C1(n3915), .C2(keyinput103), 
        .A(n3914), .ZN(n3921) );
  XNOR2_X1 U4725 ( .A(n3917), .B(keyinput83), .ZN(n3920) );
  XNOR2_X1 U4726 ( .A(n3918), .B(keyinput51), .ZN(n3919) );
  OR3_X1 U4727 ( .A1(n3921), .A2(n3920), .A3(n3919), .ZN(n3926) );
  AOI22_X1 U4728 ( .A1(n4921), .A2(keyinput115), .B1(keyinput75), .B2(n4929), 
        .ZN(n3922) );
  OAI221_X1 U4729 ( .B1(n4921), .B2(keyinput115), .C1(n4929), .C2(keyinput75), 
        .A(n3922), .ZN(n3925) );
  AOI22_X1 U4730 ( .A1(n4926), .A2(keyinput111), .B1(n4922), .B2(keyinput79), 
        .ZN(n3923) );
  OAI221_X1 U4731 ( .B1(n4926), .B2(keyinput111), .C1(n4922), .C2(keyinput79), 
        .A(n3923), .ZN(n3924) );
  NOR3_X1 U4732 ( .A1(n3926), .A2(n3925), .A3(n3924), .ZN(n3956) );
  AOI22_X1 U4733 ( .A1(n3928), .A2(keyinput26), .B1(n4917), .B2(keyinput29), 
        .ZN(n3927) );
  OAI221_X1 U4734 ( .B1(n3928), .B2(keyinput26), .C1(n4917), .C2(keyinput29), 
        .A(n3927), .ZN(n3941) );
  INV_X1 U4735 ( .A(DATAI_4_), .ZN(n3930) );
  AOI22_X1 U4736 ( .A1(n3931), .A2(keyinput35), .B1(n3930), .B2(keyinput67), 
        .ZN(n3929) );
  OAI221_X1 U4737 ( .B1(n3931), .B2(keyinput35), .C1(n3930), .C2(keyinput67), 
        .A(n3929), .ZN(n3940) );
  AOI22_X1 U4738 ( .A1(n3934), .A2(keyinput30), .B1(n3933), .B2(keyinput20), 
        .ZN(n3932) );
  OAI221_X1 U4739 ( .B1(n3934), .B2(keyinput30), .C1(n3933), .C2(keyinput20), 
        .A(n3932), .ZN(n3939) );
  XOR2_X1 U4740 ( .A(n3935), .B(keyinput59), .Z(n3937) );
  XNOR2_X1 U4741 ( .A(IR_REG_4__SCAN_IN), .B(keyinput71), .ZN(n3936) );
  NAND2_X1 U4742 ( .A1(n3937), .A2(n3936), .ZN(n3938) );
  NOR4_X1 U4743 ( .A1(n3941), .A2(n3940), .A3(n3939), .A4(n3938), .ZN(n3955)
         );
  INV_X1 U4744 ( .A(D_REG_21__SCAN_IN), .ZN(n4920) );
  AOI22_X1 U4745 ( .A1(n4920), .A2(keyinput25), .B1(keyinput24), .B2(n3943), 
        .ZN(n3942) );
  OAI221_X1 U4746 ( .B1(n4920), .B2(keyinput25), .C1(n3943), .C2(keyinput24), 
        .A(n3942), .ZN(n3953) );
  AOI22_X1 U4747 ( .A1(n3946), .A2(keyinput34), .B1(n3945), .B2(keyinput4), 
        .ZN(n3944) );
  OAI221_X1 U4748 ( .B1(n3946), .B2(keyinput34), .C1(n3945), .C2(keyinput4), 
        .A(n3944), .ZN(n3952) );
  XNOR2_X1 U4749 ( .A(IR_REG_22__SCAN_IN), .B(keyinput6), .ZN(n3949) );
  XNOR2_X1 U4750 ( .A(IR_REG_5__SCAN_IN), .B(keyinput32), .ZN(n3948) );
  XNOR2_X1 U4751 ( .A(IR_REG_12__SCAN_IN), .B(keyinput40), .ZN(n3947) );
  NAND3_X1 U4752 ( .A1(n3949), .A2(n3948), .A3(n3947), .ZN(n3951) );
  XNOR2_X1 U4753 ( .A(n4925), .B(keyinput0), .ZN(n3950) );
  NOR4_X1 U4754 ( .A1(n3953), .A2(n3952), .A3(n3951), .A4(n3950), .ZN(n3954)
         );
  NAND4_X1 U4755 ( .A1(n3957), .A2(n3956), .A3(n3955), .A4(n3954), .ZN(n4126)
         );
  AOI22_X1 U4756 ( .A1(n3960), .A2(keyinput21), .B1(keyinput10), .B2(n3959), 
        .ZN(n3958) );
  OAI221_X1 U4757 ( .B1(n3960), .B2(keyinput21), .C1(n3959), .C2(keyinput10), 
        .A(n3958), .ZN(n3964) );
  INV_X1 U4758 ( .A(D_REG_14__SCAN_IN), .ZN(n4924) );
  XNOR2_X1 U4759 ( .A(n4924), .B(keyinput117), .ZN(n3963) );
  XNOR2_X1 U4760 ( .A(n3961), .B(keyinput118), .ZN(n3962) );
  OR3_X1 U4761 ( .A1(n3964), .A2(n3963), .A3(n3962), .ZN(n3972) );
  AOI22_X1 U4762 ( .A1(n4927), .A2(keyinput124), .B1(keyinput121), .B2(n3966), 
        .ZN(n3965) );
  OAI221_X1 U4763 ( .B1(n4927), .B2(keyinput124), .C1(n3966), .C2(keyinput121), 
        .A(n3965), .ZN(n3971) );
  AOI22_X1 U4764 ( .A1(n3969), .A2(keyinput112), .B1(keyinput110), .B2(n3968), 
        .ZN(n3967) );
  OAI221_X1 U4765 ( .B1(n3969), .B2(keyinput112), .C1(n3968), .C2(keyinput110), 
        .A(n3967), .ZN(n3970) );
  NOR3_X1 U4766 ( .A1(n3972), .A2(n3971), .A3(n3970), .ZN(n4016) );
  AOI22_X1 U4767 ( .A1(n3975), .A2(keyinput102), .B1(keyinput98), .B2(n3974), 
        .ZN(n3973) );
  OAI221_X1 U4768 ( .B1(n3975), .B2(keyinput102), .C1(n3974), .C2(keyinput98), 
        .A(n3973), .ZN(n3984) );
  AOI22_X1 U4769 ( .A1(n3977), .A2(keyinput84), .B1(n3855), .B2(keyinput86), 
        .ZN(n3976) );
  OAI221_X1 U4770 ( .B1(n3977), .B2(keyinput84), .C1(n3855), .C2(keyinput86), 
        .A(n3976), .ZN(n3983) );
  XNOR2_X1 U4771 ( .A(IR_REG_2__SCAN_IN), .B(keyinput89), .ZN(n3981) );
  XNOR2_X1 U4772 ( .A(IR_REG_19__SCAN_IN), .B(keyinput96), .ZN(n3980) );
  XNOR2_X1 U4773 ( .A(IR_REG_28__SCAN_IN), .B(keyinput82), .ZN(n3979) );
  XNOR2_X1 U4774 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput81), .ZN(n3978) );
  NAND4_X1 U4775 ( .A1(n3981), .A2(n3980), .A3(n3979), .A4(n3978), .ZN(n3982)
         );
  NOR3_X1 U4776 ( .A1(n3984), .A2(n3983), .A3(n3982), .ZN(n4015) );
  AOI22_X1 U4777 ( .A1(n4918), .A2(keyinput74), .B1(keyinput73), .B2(n3986), 
        .ZN(n3985) );
  OAI221_X1 U4778 ( .B1(n4918), .B2(keyinput74), .C1(n3986), .C2(keyinput73), 
        .A(n3985), .ZN(n3992) );
  XNOR2_X1 U4779 ( .A(n3987), .B(keyinput70), .ZN(n3991) );
  XNOR2_X1 U4780 ( .A(n3988), .B(keyinput80), .ZN(n3990) );
  XNOR2_X1 U4781 ( .A(n2846), .B(keyinput66), .ZN(n3989) );
  OR4_X1 U4782 ( .A1(n3992), .A2(n3991), .A3(n3990), .A4(n3989), .ZN(n3998) );
  INV_X1 U4783 ( .A(DATAI_23_), .ZN(n4932) );
  AOI22_X1 U4784 ( .A1(n4932), .A2(keyinput72), .B1(n3994), .B2(keyinput68), 
        .ZN(n3993) );
  OAI221_X1 U4785 ( .B1(n4932), .B2(keyinput72), .C1(n3994), .C2(keyinput68), 
        .A(n3993), .ZN(n3997) );
  XNOR2_X1 U4786 ( .A(n3995), .B(keyinput78), .ZN(n3996) );
  NOR3_X1 U4787 ( .A1(n3998), .A2(n3997), .A3(n3996), .ZN(n4014) );
  INV_X1 U4788 ( .A(D_REG_17__SCAN_IN), .ZN(n4923) );
  AOI22_X1 U4789 ( .A1(n4923), .A2(keyinput54), .B1(keyinput49), .B2(n4000), 
        .ZN(n3999) );
  OAI221_X1 U4790 ( .B1(n4923), .B2(keyinput54), .C1(n4000), .C2(keyinput49), 
        .A(n3999), .ZN(n4012) );
  AOI22_X1 U4791 ( .A1(n4003), .A2(keyinput64), .B1(keyinput58), .B2(n4002), 
        .ZN(n4001) );
  OAI221_X1 U4792 ( .B1(n4003), .B2(keyinput64), .C1(n4002), .C2(keyinput58), 
        .A(n4001), .ZN(n4011) );
  INV_X1 U4793 ( .A(D_REG_24__SCAN_IN), .ZN(n4919) );
  INV_X1 U4794 ( .A(DATAI_22_), .ZN(n4005) );
  AOI22_X1 U4795 ( .A1(n4919), .A2(keyinput61), .B1(keyinput56), .B2(n4005), 
        .ZN(n4004) );
  OAI221_X1 U4796 ( .B1(n4919), .B2(keyinput61), .C1(n4005), .C2(keyinput56), 
        .A(n4004), .ZN(n4010) );
  XOR2_X1 U4797 ( .A(n4006), .B(keyinput42), .Z(n4008) );
  XNOR2_X1 U4798 ( .A(IR_REG_17__SCAN_IN), .B(keyinput44), .ZN(n4007) );
  NAND2_X1 U4799 ( .A1(n4008), .A2(n4007), .ZN(n4009) );
  NOR4_X1 U4800 ( .A1(n4012), .A2(n4011), .A3(n4010), .A4(n4009), .ZN(n4013)
         );
  NAND4_X1 U4801 ( .A1(n4016), .A2(n4015), .A3(n4014), .A4(n4013), .ZN(n4125)
         );
  AOI22_X1 U4802 ( .A1(n4018), .A2(keyinput31), .B1(n4989), .B2(keyinput57), 
        .ZN(n4017) );
  OAI221_X1 U4803 ( .B1(n4018), .B2(keyinput31), .C1(n4989), .C2(keyinput57), 
        .A(n4017), .ZN(n4028) );
  AOI22_X1 U4804 ( .A1(n4973), .A2(keyinput36), .B1(n2611), .B2(keyinput53), 
        .ZN(n4019) );
  OAI221_X1 U4805 ( .B1(n4973), .B2(keyinput36), .C1(n2611), .C2(keyinput53), 
        .A(n4019), .ZN(n4027) );
  AOI22_X1 U4806 ( .A1(n4022), .A2(keyinput63), .B1(keyinput47), .B2(n4021), 
        .ZN(n4020) );
  OAI221_X1 U4807 ( .B1(n4022), .B2(keyinput63), .C1(n4021), .C2(keyinput47), 
        .A(n4020), .ZN(n4026) );
  XNOR2_X1 U4808 ( .A(REG1_REG_12__SCAN_IN), .B(keyinput107), .ZN(n4024) );
  XNOR2_X1 U4809 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput12), .ZN(n4023) );
  NAND2_X1 U4810 ( .A1(n4024), .A2(n4023), .ZN(n4025) );
  NOR4_X1 U4811 ( .A1(n4028), .A2(n4027), .A3(n4026), .A4(n4025), .ZN(n4070)
         );
  AOI22_X1 U4812 ( .A1(n4031), .A2(keyinput52), .B1(n4030), .B2(keyinput88), 
        .ZN(n4029) );
  OAI221_X1 U4813 ( .B1(n4031), .B2(keyinput52), .C1(n4030), .C2(keyinput88), 
        .A(n4029), .ZN(n4041) );
  AOI22_X1 U4814 ( .A1(n3652), .A2(keyinput114), .B1(keyinput23), .B2(n4667), 
        .ZN(n4032) );
  OAI221_X1 U4815 ( .B1(n3652), .B2(keyinput114), .C1(n4667), .C2(keyinput23), 
        .A(n4032), .ZN(n4040) );
  AOI22_X1 U4816 ( .A1(n4034), .A2(keyinput33), .B1(keyinput77), .B2(n3168), 
        .ZN(n4033) );
  OAI221_X1 U4817 ( .B1(n4034), .B2(keyinput33), .C1(n3168), .C2(keyinput77), 
        .A(n4033), .ZN(n4039) );
  AOI22_X1 U4818 ( .A1(n4037), .A2(keyinput39), .B1(n4036), .B2(keyinput48), 
        .ZN(n4035) );
  OAI221_X1 U4819 ( .B1(n4037), .B2(keyinput39), .C1(n4036), .C2(keyinput48), 
        .A(n4035), .ZN(n4038) );
  NOR4_X1 U4820 ( .A1(n4041), .A2(n4040), .A3(n4039), .A4(n4038), .ZN(n4069)
         );
  INV_X1 U4821 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U4822 ( .A1(n4043), .A2(keyinput106), .B1(n4768), .B2(keyinput116), 
        .ZN(n4042) );
  OAI221_X1 U4823 ( .B1(n4043), .B2(keyinput106), .C1(n4768), .C2(keyinput116), 
        .A(n4042), .ZN(n4052) );
  INV_X1 U4824 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4706) );
  AOI22_X1 U4825 ( .A1(n4706), .A2(keyinput1), .B1(n4539), .B2(keyinput99), 
        .ZN(n4044) );
  OAI221_X1 U4826 ( .B1(n4706), .B2(keyinput1), .C1(n4539), .C2(keyinput99), 
        .A(n4044), .ZN(n4051) );
  INV_X1 U4827 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4773) );
  AOI22_X1 U4828 ( .A1(n4773), .A2(keyinput50), .B1(n4046), .B2(keyinput76), 
        .ZN(n4045) );
  OAI221_X1 U4829 ( .B1(n4773), .B2(keyinput50), .C1(n4046), .C2(keyinput76), 
        .A(n4045), .ZN(n4050) );
  XNOR2_X1 U4830 ( .A(REG0_REG_16__SCAN_IN), .B(keyinput113), .ZN(n4048) );
  XNOR2_X1 U4831 ( .A(IR_REG_11__SCAN_IN), .B(keyinput65), .ZN(n4047) );
  NAND2_X1 U4832 ( .A1(n4048), .A2(n4047), .ZN(n4049) );
  NOR4_X1 U4833 ( .A1(n4052), .A2(n4051), .A3(n4050), .A4(n4049), .ZN(n4068)
         );
  AOI22_X1 U4834 ( .A1(n4055), .A2(keyinput16), .B1(n4054), .B2(keyinput93), 
        .ZN(n4053) );
  OAI221_X1 U4835 ( .B1(n4055), .B2(keyinput16), .C1(n4054), .C2(keyinput93), 
        .A(n4053), .ZN(n4066) );
  INV_X1 U4836 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4846) );
  AOI22_X1 U4837 ( .A1(n4846), .A2(keyinput91), .B1(n4057), .B2(keyinput8), 
        .ZN(n4056) );
  OAI221_X1 U4838 ( .B1(n4846), .B2(keyinput91), .C1(n4057), .C2(keyinput8), 
        .A(n4056), .ZN(n4065) );
  AOI22_X1 U4839 ( .A1(n4060), .A2(keyinput45), .B1(n4059), .B2(keyinput19), 
        .ZN(n4058) );
  OAI221_X1 U4840 ( .B1(n4060), .B2(keyinput45), .C1(n4059), .C2(keyinput19), 
        .A(n4058), .ZN(n4064) );
  XNOR2_X1 U4841 ( .A(IR_REG_7__SCAN_IN), .B(keyinput60), .ZN(n4062) );
  XNOR2_X1 U4842 ( .A(keyinput5), .B(DATAI_9_), .ZN(n4061) );
  NAND2_X1 U4843 ( .A1(n4062), .A2(n4061), .ZN(n4063) );
  NOR4_X1 U4844 ( .A1(n4066), .A2(n4065), .A3(n4064), .A4(n4063), .ZN(n4067)
         );
  NAND4_X1 U4845 ( .A1(n4070), .A2(n4069), .A3(n4068), .A4(n4067), .ZN(n4124)
         );
  INV_X1 U4846 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U4847 ( .A1(n4073), .A2(keyinput97), .B1(keyinput9), .B2(n4072), 
        .ZN(n4071) );
  OAI221_X1 U4848 ( .B1(n4073), .B2(keyinput97), .C1(n4072), .C2(keyinput9), 
        .A(n4071), .ZN(n4083) );
  INV_X1 U4849 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4985) );
  INV_X1 U4850 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n4075) );
  AOI22_X1 U4851 ( .A1(n4985), .A2(keyinput94), .B1(keyinput69), .B2(n4075), 
        .ZN(n4074) );
  OAI221_X1 U4852 ( .B1(n4985), .B2(keyinput94), .C1(n4075), .C2(keyinput69), 
        .A(n4074), .ZN(n4082) );
  AOI22_X1 U4853 ( .A1(n4077), .A2(keyinput125), .B1(keyinput105), .B2(n2237), 
        .ZN(n4076) );
  OAI221_X1 U4854 ( .B1(n4077), .B2(keyinput125), .C1(n2237), .C2(keyinput105), 
        .A(n4076), .ZN(n4081) );
  XNOR2_X1 U4855 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput41), .ZN(n4079) );
  XNOR2_X1 U4856 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput28), .ZN(n4078) );
  NAND2_X1 U4857 ( .A1(n4079), .A2(n4078), .ZN(n4080) );
  NOR4_X1 U4858 ( .A1(n4083), .A2(n4082), .A3(n4081), .A4(n4080), .ZN(n4122)
         );
  AOI22_X1 U4859 ( .A1(n4085), .A2(keyinput123), .B1(keyinput38), .B2(n4449), 
        .ZN(n4084) );
  OAI221_X1 U4860 ( .B1(n4085), .B2(keyinput123), .C1(n4449), .C2(keyinput38), 
        .A(n4084), .ZN(n4097) );
  AOI22_X1 U4861 ( .A1(n4088), .A2(keyinput109), .B1(n4087), .B2(keyinput37), 
        .ZN(n4086) );
  OAI221_X1 U4862 ( .B1(n4088), .B2(keyinput109), .C1(n4087), .C2(keyinput37), 
        .A(n4086), .ZN(n4096) );
  AOI22_X1 U4863 ( .A1(n4635), .A2(keyinput2), .B1(n4090), .B2(keyinput119), 
        .ZN(n4089) );
  OAI221_X1 U4864 ( .B1(n4635), .B2(keyinput2), .C1(n4090), .C2(keyinput119), 
        .A(n4089), .ZN(n4095) );
  NAND2_X1 U4865 ( .A1(n4129), .A2(IR_REG_21__SCAN_IN), .ZN(n4092) );
  NAND2_X1 U4866 ( .A1(n4093), .A2(keyinput120), .ZN(n4091) );
  OAI211_X1 U4867 ( .C1(keyinput120), .C2(n4093), .A(n4092), .B(n4091), .ZN(
        n4094) );
  NOR4_X1 U4868 ( .A1(n4097), .A2(n4096), .A3(n4095), .A4(n4094), .ZN(n4121)
         );
  AOI22_X1 U4869 ( .A1(n3513), .A2(keyinput85), .B1(n4099), .B2(keyinput22), 
        .ZN(n4098) );
  OAI221_X1 U4870 ( .B1(n3513), .B2(keyinput85), .C1(n4099), .C2(keyinput22), 
        .A(n4098), .ZN(n4109) );
  INV_X1 U4871 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4987) );
  AOI22_X1 U4872 ( .A1(n4101), .A2(keyinput13), .B1(n4987), .B2(keyinput11), 
        .ZN(n4100) );
  OAI221_X1 U4873 ( .B1(n4101), .B2(keyinput13), .C1(n4987), .C2(keyinput11), 
        .A(n4100), .ZN(n4108) );
  AOI22_X1 U4874 ( .A1(n4103), .A2(keyinput104), .B1(n3637), .B2(keyinput55), 
        .ZN(n4102) );
  OAI221_X1 U4875 ( .B1(n4103), .B2(keyinput104), .C1(n3637), .C2(keyinput55), 
        .A(n4102), .ZN(n4107) );
  XNOR2_X1 U4876 ( .A(REG3_REG_2__SCAN_IN), .B(keyinput100), .ZN(n4105) );
  XNOR2_X1 U4877 ( .A(IR_REG_0__SCAN_IN), .B(keyinput14), .ZN(n4104) );
  NAND2_X1 U4878 ( .A1(n4105), .A2(n4104), .ZN(n4106) );
  NOR4_X1 U4879 ( .A1(n4109), .A2(n4108), .A3(n4107), .A4(n4106), .ZN(n4120)
         );
  AOI22_X1 U4880 ( .A1(n4578), .A2(keyinput3), .B1(keyinput18), .B2(n4867), 
        .ZN(n4110) );
  OAI221_X1 U4881 ( .B1(n4578), .B2(keyinput3), .C1(n4867), .C2(keyinput18), 
        .A(n4110), .ZN(n4118) );
  AOI22_X1 U4882 ( .A1(n3159), .A2(keyinput122), .B1(n4982), .B2(keyinput62), 
        .ZN(n4111) );
  OAI221_X1 U4883 ( .B1(n3159), .B2(keyinput122), .C1(n4982), .C2(keyinput62), 
        .A(n4111), .ZN(n4117) );
  AOI22_X1 U4884 ( .A1(n2236), .A2(keyinput101), .B1(keyinput43), .B2(n4503), 
        .ZN(n4112) );
  OAI221_X1 U4885 ( .B1(n2236), .B2(keyinput101), .C1(n4503), .C2(keyinput43), 
        .A(n4112), .ZN(n4116) );
  XNOR2_X1 U4886 ( .A(REG3_REG_12__SCAN_IN), .B(keyinput95), .ZN(n4114) );
  XNOR2_X1 U4887 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput7), .ZN(n4113) );
  NAND2_X1 U4888 ( .A1(n4114), .A2(n4113), .ZN(n4115) );
  NOR4_X1 U4889 ( .A1(n4118), .A2(n4117), .A3(n4116), .A4(n4115), .ZN(n4119)
         );
  NAND4_X1 U4890 ( .A1(n4122), .A2(n4121), .A3(n4120), .A4(n4119), .ZN(n4123)
         );
  NOR4_X1 U4891 ( .A1(n4126), .A2(n4125), .A3(n4124), .A4(n4123), .ZN(n4127)
         );
  OAI21_X1 U4892 ( .B1(n4129), .B2(n4128), .A(n4127), .ZN(n4143) );
  OAI21_X1 U4893 ( .B1(n4132), .B2(n4131), .A(n4130), .ZN(n4141) );
  OAI22_X1 U4894 ( .A1(n3090), .A2(n2458), .B1(n4134), .B2(n4133), .ZN(n4139)
         );
  OAI22_X1 U4895 ( .A1(n4137), .A2(n4136), .B1(n2885), .B2(n4135), .ZN(n4138)
         );
  AOI211_X1 U4896 ( .C1(n4141), .C2(n4140), .A(n4139), .B(n4138), .ZN(n4142)
         );
  XOR2_X1 U4897 ( .A(n4143), .B(n4142), .Z(U3234) );
  NAND2_X1 U4898 ( .A1(n2231), .A2(n4145), .ZN(n4146) );
  XNOR2_X1 U4899 ( .A(n4147), .B(n4146), .ZN(n4152) );
  AOI22_X1 U4900 ( .A1(n4166), .A2(n4610), .B1(n4167), .B2(n4341), .ZN(n4151)
         );
  NOR2_X1 U4901 ( .A1(n2236), .A2(STATE_REG_SCAN_IN), .ZN(n4882) );
  NOR2_X1 U4902 ( .A1(n4169), .A2(n4620), .ZN(n4148) );
  AOI211_X1 U4903 ( .C1(n4149), .C2(n4171), .A(n4882), .B(n4148), .ZN(n4150)
         );
  OAI211_X1 U4904 ( .C1(n4152), .C2(n4175), .A(n4151), .B(n4150), .ZN(U3235)
         );
  NAND2_X1 U4905 ( .A1(n4498), .A2(n4167), .ZN(n4157) );
  AOI22_X1 U4906 ( .A1(n4171), .A2(n4155), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n4156) );
  OAI211_X1 U4907 ( .C1(n4169), .C2(n4470), .A(n4157), .B(n4156), .ZN(n4158)
         );
  AOI21_X1 U4908 ( .B1(n4166), .B2(n4463), .A(n4158), .ZN(n4159) );
  OAI21_X1 U4909 ( .B1(n4160), .B2(n4175), .A(n4159), .ZN(U3237) );
  INV_X1 U4910 ( .A(n4161), .ZN(n4162) );
  NOR2_X1 U4911 ( .A1(n4163), .A2(n4162), .ZN(n4165) );
  XNOR2_X1 U4912 ( .A(n4165), .B(n4164), .ZN(n4176) );
  AOI22_X1 U4913 ( .A1(n4167), .A2(n4659), .B1(n4166), .B2(n4629), .ZN(n4174)
         );
  AND2_X1 U4914 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4857) );
  NOR2_X1 U4915 ( .A1(n4169), .A2(n4168), .ZN(n4170) );
  AOI211_X1 U4916 ( .C1(n4172), .C2(n4171), .A(n4857), .B(n4170), .ZN(n4173)
         );
  OAI211_X1 U4917 ( .C1(n4176), .C2(n4175), .A(n4174), .B(n4173), .ZN(U3238)
         );
  INV_X1 U4918 ( .A(n4412), .ZN(n4323) );
  NAND2_X1 U4919 ( .A1(n4177), .A2(DATAI_31_), .ZN(n4413) );
  INV_X1 U4920 ( .A(n4413), .ZN(n4322) );
  NOR2_X1 U4921 ( .A1(n4323), .A2(n4322), .ZN(n4247) );
  NAND2_X1 U4922 ( .A1(n4178), .A2(DATAI_30_), .ZN(n4417) );
  AND2_X1 U4923 ( .A1(n4339), .A2(n4417), .ZN(n4324) );
  INV_X1 U4924 ( .A(n4324), .ZN(n4179) );
  OAI21_X1 U4925 ( .B1(n4412), .B2(n4413), .A(n4179), .ZN(n4259) );
  INV_X1 U4926 ( .A(n4257), .ZN(n4181) );
  NAND2_X1 U4927 ( .A1(n2881), .A2(n4903), .ZN(n4256) );
  OAI211_X1 U4928 ( .C1(n4181), .C2(n4327), .A(n4256), .B(n4180), .ZN(n4184)
         );
  NAND3_X1 U4929 ( .A1(n4184), .A2(n4183), .A3(n4182), .ZN(n4187) );
  NAND3_X1 U4930 ( .A1(n4187), .A2(n4186), .A3(n4185), .ZN(n4190) );
  NAND3_X1 U4931 ( .A1(n4190), .A2(n4189), .A3(n4188), .ZN(n4192) );
  NAND4_X1 U4932 ( .A1(n4192), .A2(n4191), .A3(n4202), .A4(n2167), .ZN(n4195)
         );
  AND3_X1 U4933 ( .A1(n4195), .A2(n4194), .A3(n4193), .ZN(n4200) );
  NAND2_X1 U4934 ( .A1(n4197), .A2(n4196), .ZN(n4205) );
  OAI211_X1 U4935 ( .C1(n4200), .C2(n4205), .A(n4199), .B(n4198), .ZN(n4201)
         );
  NAND4_X1 U4936 ( .A1(n4201), .A2(n4208), .A3(n4209), .A4(n2335), .ZN(n4214)
         );
  INV_X1 U4937 ( .A(n4202), .ZN(n4206) );
  NOR4_X1 U4938 ( .A1(n4206), .A2(n4205), .A3(n4204), .A4(n4203), .ZN(n4211)
         );
  NAND2_X1 U4939 ( .A1(n4209), .A2(n4208), .ZN(n4210) );
  NAND2_X1 U4940 ( .A1(n4210), .A2(n4216), .ZN(n4296) );
  OAI21_X1 U4941 ( .B1(n4211), .B2(n2330), .A(n4296), .ZN(n4213) );
  AOI211_X1 U4942 ( .C1(n4214), .C2(n4213), .A(n2334), .B(n2169), .ZN(n4221)
         );
  NAND2_X1 U4943 ( .A1(n4216), .A2(n4215), .ZN(n4297) );
  INV_X1 U4944 ( .A(n4297), .ZN(n4218) );
  INV_X1 U4945 ( .A(n4296), .ZN(n4217) );
  AOI21_X1 U4946 ( .B1(n4219), .B2(n4218), .A(n4217), .ZN(n4220) );
  OAI21_X1 U4947 ( .B1(n4221), .B2(n4220), .A(n4298), .ZN(n4223) );
  INV_X1 U4948 ( .A(n4299), .ZN(n4222) );
  AOI211_X1 U4949 ( .C1(n4223), .C2(n4302), .A(n4222), .B(n4301), .ZN(n4224)
         );
  INV_X1 U4950 ( .A(n4510), .ZN(n4265) );
  OAI21_X1 U4951 ( .B1(n4224), .B2(n4304), .A(n4265), .ZN(n4226) );
  AOI21_X1 U4952 ( .B1(n4226), .B2(n4306), .A(n4225), .ZN(n4229) );
  INV_X1 U4953 ( .A(n4249), .ZN(n4227) );
  NOR2_X1 U4954 ( .A1(n4227), .A2(n4252), .ZN(n4310) );
  INV_X1 U4955 ( .A(n4310), .ZN(n4228) );
  NOR3_X1 U4956 ( .A1(n4229), .A2(n4313), .A3(n4228), .ZN(n4245) );
  INV_X1 U4957 ( .A(n4240), .ZN(n4231) );
  OAI21_X1 U4958 ( .B1(n4231), .B2(n4237), .A(n4230), .ZN(n4317) );
  INV_X1 U4959 ( .A(n4317), .ZN(n4234) );
  NAND3_X1 U4960 ( .A1(n4234), .A2(n4233), .A3(n4232), .ZN(n4244) );
  NAND2_X1 U4961 ( .A1(n4236), .A2(n4235), .ZN(n4314) );
  INV_X1 U4962 ( .A(n4314), .ZN(n4242) );
  INV_X1 U4963 ( .A(n4237), .ZN(n4239) );
  INV_X1 U4964 ( .A(n4339), .ZN(n4238) );
  INV_X1 U4965 ( .A(n4417), .ZN(n4420) );
  AOI21_X1 U4966 ( .B1(n4238), .B2(n4420), .A(n4247), .ZN(n4261) );
  OAI21_X1 U4967 ( .B1(n4240), .B2(n4239), .A(n4261), .ZN(n4312) );
  INV_X1 U4968 ( .A(n4312), .ZN(n4241) );
  OAI21_X1 U4969 ( .B1(n4242), .B2(n4317), .A(n4241), .ZN(n4319) );
  INV_X1 U4970 ( .A(n4319), .ZN(n4243) );
  OAI21_X1 U4971 ( .B1(n4245), .B2(n4244), .A(n4243), .ZN(n4246) );
  OAI21_X1 U4972 ( .B1(n4247), .B2(n4260), .A(n4246), .ZN(n4331) );
  INV_X1 U4973 ( .A(n4248), .ZN(n4295) );
  INV_X1 U4974 ( .A(n4532), .ZN(n4294) );
  NAND2_X1 U4975 ( .A1(n4249), .A2(n4476), .ZN(n4496) );
  INV_X1 U4976 ( .A(n4250), .ZN(n4251) );
  OR2_X1 U4977 ( .A1(n4252), .A2(n4251), .ZN(n4514) );
  NAND2_X1 U4978 ( .A1(n4254), .A2(n4253), .ZN(n4653) );
  NOR2_X1 U4979 ( .A1(n4653), .A2(n4255), .ZN(n4264) );
  AND2_X1 U4980 ( .A1(n4257), .A2(n4256), .ZN(n4911) );
  XNOR2_X1 U4981 ( .A(n4437), .B(n4467), .ZN(n4460) );
  NAND2_X1 U4982 ( .A1(n4265), .A2(n4511), .ZN(n4549) );
  INV_X1 U4983 ( .A(n4549), .ZN(n4292) );
  INV_X1 U4984 ( .A(n4266), .ZN(n4268) );
  OR2_X1 U4985 ( .A1(n4270), .A2(n2196), .ZN(n4590) );
  NAND4_X1 U4986 ( .A1(n4274), .A2(n4273), .A3(n4272), .A4(n4271), .ZN(n4281)
         );
  INV_X1 U4987 ( .A(n3287), .ZN(n4278) );
  NAND4_X1 U4988 ( .A1(n4278), .A2(n4277), .A3(n4276), .A4(n4275), .ZN(n4280)
         );
  NOR3_X1 U4989 ( .A1(n4281), .A2(n4280), .A3(n4279), .ZN(n4282) );
  NAND2_X1 U4990 ( .A1(n4590), .A2(n4282), .ZN(n4283) );
  NOR2_X1 U4991 ( .A1(n4571), .A2(n4283), .ZN(n4291) );
  INV_X1 U4992 ( .A(n4586), .ZN(n4284) );
  NAND2_X1 U4993 ( .A1(n4284), .A2(n4585), .ZN(n4639) );
  INV_X1 U4994 ( .A(n4639), .ZN(n4289) );
  NOR2_X1 U4995 ( .A1(n4286), .A2(n4285), .ZN(n4287) );
  NAND4_X1 U4996 ( .A1(n4295), .A2(n4294), .A3(n2349), .A4(n4293), .ZN(n4329)
         );
  OAI21_X1 U4997 ( .B1(n3604), .B2(n4297), .A(n4296), .ZN(n4303) );
  NAND2_X1 U4998 ( .A1(n4299), .A2(n4298), .ZN(n4300) );
  AOI211_X1 U4999 ( .C1(n4303), .C2(n4302), .A(n4301), .B(n4300), .ZN(n4309)
         );
  INV_X1 U5000 ( .A(n4304), .ZN(n4305) );
  NAND2_X1 U5001 ( .A1(n4306), .A2(n4305), .ZN(n4308) );
  OAI21_X1 U5002 ( .B1(n4309), .B2(n4308), .A(n4307), .ZN(n4311) );
  AOI21_X1 U5003 ( .B1(n4311), .B2(n4310), .A(n4457), .ZN(n4315) );
  NOR4_X1 U5004 ( .A1(n4315), .A2(n4314), .A3(n4313), .A4(n4312), .ZN(n4321)
         );
  NOR3_X1 U5005 ( .A1(n4317), .A2(n4445), .A3(n4316), .ZN(n4318) );
  NOR2_X1 U5006 ( .A1(n4319), .A2(n4318), .ZN(n4320) );
  OAI22_X1 U5007 ( .A1(n4321), .A2(n4320), .B1(n4412), .B2(n4417), .ZN(n4326)
         );
  OAI21_X1 U5008 ( .B1(n4324), .B2(n4323), .A(n4322), .ZN(n4325) );
  NAND2_X1 U5009 ( .A1(n4326), .A2(n4325), .ZN(n4328) );
  MUX2_X1 U5010 ( .A(n4329), .B(n4328), .S(n4327), .Z(n4330) );
  MUX2_X1 U5011 ( .A(n4331), .B(n4330), .S(n4793), .Z(n4332) );
  XNOR2_X1 U5012 ( .A(n4332), .B(n4812), .ZN(n4338) );
  NAND4_X1 U5013 ( .A1(n2962), .A2(n4931), .A3(n4334), .A4(n4333), .ZN(n4335)
         );
  OAI211_X1 U5014 ( .C1(n4792), .C2(n4337), .A(n4335), .B(B_REG_SCAN_IN), .ZN(
        n4336) );
  OAI21_X1 U5015 ( .B1(n4338), .B2(n4337), .A(n4336), .ZN(U3239) );
  MUX2_X1 U5016 ( .A(DATAO_REG_30__SCAN_IN), .B(n4339), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U5017 ( .A(DATAO_REG_28__SCAN_IN), .B(n4444), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U5018 ( .A(DATAO_REG_26__SCAN_IN), .B(n4482), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U5019 ( .A(DATAO_REG_23__SCAN_IN), .B(n4340), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U5020 ( .A(DATAO_REG_17__SCAN_IN), .B(n4341), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U5021 ( .A(DATAO_REG_14__SCAN_IN), .B(n4659), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U5022 ( .A(DATAO_REG_11__SCAN_IN), .B(n4342), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U5023 ( .A(DATAO_REG_9__SCAN_IN), .B(n4343), .S(U4043), .Z(U3559) );
  MUX2_X1 U5024 ( .A(DATAO_REG_8__SCAN_IN), .B(n4344), .S(U4043), .Z(U3558) );
  MUX2_X1 U5025 ( .A(DATAO_REG_5__SCAN_IN), .B(n4345), .S(U4043), .Z(U3555) );
  MUX2_X1 U5026 ( .A(DATAO_REG_4__SCAN_IN), .B(n4346), .S(U4043), .Z(U3554) );
  MUX2_X1 U5027 ( .A(DATAO_REG_2__SCAN_IN), .B(n4347), .S(U4043), .Z(U3552) );
  MUX2_X1 U5028 ( .A(DATAO_REG_0__SCAN_IN), .B(n2881), .S(U4043), .Z(U3550) );
  OAI211_X1 U5029 ( .C1(n4359), .C2(n4349), .A(n4875), .B(n4348), .ZN(n4355)
         );
  OAI211_X1 U5030 ( .C1(n4351), .C2(n4350), .A(n4873), .B(n4364), .ZN(n4354)
         );
  AOI22_X1 U5031 ( .A1(n4881), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4353) );
  NAND2_X1 U5032 ( .A1(n4849), .A2(n4798), .ZN(n4352) );
  NAND4_X1 U5033 ( .A1(n4355), .A2(n4354), .A3(n4353), .A4(n4352), .ZN(U3241)
         );
  NAND2_X1 U5034 ( .A1(n4356), .A2(n4358), .ZN(n4357) );
  OAI211_X1 U5035 ( .C1(n4359), .C2(n4358), .A(n4357), .B(n4790), .ZN(n4360)
         );
  OAI211_X1 U5036 ( .C1(IR_REG_0__SCAN_IN), .C2(n4361), .A(n4360), .B(n3562), 
        .ZN(n4827) );
  AOI22_X1 U5037 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4881), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4375) );
  NAND3_X1 U5038 ( .A1(n4364), .A2(n4363), .A3(n4362), .ZN(n4365) );
  NAND2_X1 U5039 ( .A1(n4849), .A2(n2130), .ZN(n4366) );
  AND2_X1 U5040 ( .A1(n4367), .A2(n4366), .ZN(n4374) );
  INV_X1 U5041 ( .A(n4368), .ZN(n4369) );
  NAND3_X1 U5042 ( .A1(n4348), .A2(n4370), .A3(n4369), .ZN(n4371) );
  NAND3_X1 U5043 ( .A1(n4875), .A2(n4372), .A3(n4371), .ZN(n4373) );
  NAND4_X1 U5044 ( .A1(n4827), .A2(n4375), .A3(n4374), .A4(n4373), .ZN(U3242)
         );
  INV_X1 U5045 ( .A(n4391), .ZN(n4803) );
  XNOR2_X1 U5046 ( .A(n4391), .B(REG2_REG_17__SCAN_IN), .ZN(n4388) );
  INV_X1 U5047 ( .A(n4941), .ZN(n4840) );
  NOR2_X1 U5048 ( .A1(n4667), .A2(n4840), .ZN(n4834) );
  NOR2_X1 U5049 ( .A1(n4397), .A2(n4381), .ZN(n4382) );
  NOR2_X1 U5050 ( .A1(n4382), .A2(n4844), .ZN(n4855) );
  INV_X1 U5051 ( .A(n4937), .ZN(n4863) );
  AOI22_X1 U5052 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4863), .B1(n4937), .B2(
        n3652), .ZN(n4854) );
  NOR2_X1 U5053 ( .A1(n4855), .A2(n4854), .ZN(n4853) );
  INV_X1 U5054 ( .A(n4936), .ZN(n4384) );
  XNOR2_X1 U5055 ( .A(n4385), .B(n4384), .ZN(n4868) );
  NAND2_X1 U5056 ( .A1(n4868), .A2(n4867), .ZN(n4866) );
  NAND2_X1 U5057 ( .A1(n4385), .A2(n4936), .ZN(n4386) );
  OAI21_X1 U5058 ( .B1(n4388), .B2(n4387), .A(n4801), .ZN(n4389) );
  AOI22_X1 U5059 ( .A1(n4803), .A2(n4849), .B1(n4875), .B2(n4389), .ZN(n4410)
         );
  AOI21_X1 U5060 ( .B1(n4881), .B2(ADDR_REG_17__SCAN_IN), .A(n4390), .ZN(n4409) );
  XNOR2_X1 U5061 ( .A(n4391), .B(REG1_REG_17__SCAN_IN), .ZN(n4406) );
  AOI22_X1 U5062 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4840), .B1(n4941), .B2(
        n4736), .ZN(n4830) );
  INV_X1 U5063 ( .A(n4830), .ZN(n4395) );
  AOI22_X1 U5064 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4863), .B1(n4937), .B2(
        n4400), .ZN(n4859) );
  NAND2_X1 U5065 ( .A1(n4402), .A2(n4936), .ZN(n4404) );
  NAND2_X1 U5066 ( .A1(n4404), .A2(n4869), .ZN(n4405) );
  NAND2_X1 U5067 ( .A1(n4405), .A2(n4406), .ZN(n4805) );
  OAI21_X1 U5068 ( .B1(n4406), .B2(n4405), .A(n4805), .ZN(n4407) );
  NAND2_X1 U5069 ( .A1(n4873), .A2(n4407), .ZN(n4408) );
  NAND3_X1 U5070 ( .A1(n4410), .A2(n4409), .A3(n4408), .ZN(U3257) );
  NAND2_X1 U5071 ( .A1(n4418), .A2(n4417), .ZN(n4416) );
  XOR2_X1 U5072 ( .A(n4413), .B(n4416), .Z(n4742) );
  NAND2_X1 U5073 ( .A1(n4412), .A2(n4411), .ZN(n4422) );
  OAI21_X1 U5074 ( .B1(n4413), .B2(n4645), .A(n4422), .ZN(n4739) );
  NAND2_X1 U5075 ( .A1(n4668), .A2(n4739), .ZN(n4415) );
  NAND2_X1 U5076 ( .A1(n4643), .A2(REG2_REG_31__SCAN_IN), .ZN(n4414) );
  OAI211_X1 U5077 ( .C1(n4742), .C2(n4600), .A(n4415), .B(n4414), .ZN(U3260)
         );
  INV_X1 U5078 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4425) );
  OAI21_X1 U5079 ( .B1(n4418), .B2(n4417), .A(n4416), .ZN(n4419) );
  INV_X1 U5080 ( .A(n4419), .ZN(n4744) );
  NAND2_X1 U5081 ( .A1(n4744), .A2(n4896), .ZN(n4424) );
  NAND2_X1 U5082 ( .A1(n4568), .A2(n4420), .ZN(n4421) );
  NAND2_X1 U5083 ( .A1(n4422), .A2(n4421), .ZN(n4745) );
  NAND2_X1 U5084 ( .A1(n4668), .A2(n4745), .ZN(n4423) );
  OAI211_X1 U5085 ( .C1(n4668), .C2(n4425), .A(n4424), .B(n4423), .ZN(U3261)
         );
  NAND2_X1 U5086 ( .A1(n4427), .A2(n4426), .ZN(n4428) );
  XOR2_X1 U5087 ( .A(n4429), .B(n4428), .Z(n4436) );
  AOI22_X1 U5088 ( .A1(n4430), .A2(n4896), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4643), .ZN(n4435) );
  OAI21_X1 U5089 ( .B1(n4432), .B2(n4665), .A(n4431), .ZN(n4433) );
  NAND2_X1 U5090 ( .A1(n4433), .A2(n4668), .ZN(n4434) );
  OAI211_X1 U5091 ( .C1(n4436), .C2(n4603), .A(n4435), .B(n4434), .ZN(U3354)
         );
  OAI22_X1 U5092 ( .A1(n4437), .A2(n4647), .B1(n4447), .B2(n4645), .ZN(n4443)
         );
  NAND2_X1 U5093 ( .A1(n4439), .A2(n4445), .ZN(n4440) );
  AOI21_X1 U5094 ( .B1(n4441), .B2(n4440), .A(n4655), .ZN(n4442) );
  AOI211_X2 U5095 ( .C1(n4660), .C2(n4444), .A(n4443), .B(n4442), .ZN(n4681)
         );
  XNOR2_X1 U5096 ( .A(n4446), .B(n4445), .ZN(n4680) );
  NAND2_X1 U5097 ( .A1(n4680), .A2(n4640), .ZN(n4454) );
  OAI21_X1 U5098 ( .B1(n4466), .B2(n4447), .A(n3109), .ZN(n4683) );
  INV_X1 U5099 ( .A(n4683), .ZN(n4452) );
  INV_X1 U5100 ( .A(n4448), .ZN(n4450) );
  OAI22_X1 U5101 ( .A1(n4450), .A2(n4665), .B1(n4449), .B2(n4668), .ZN(n4451)
         );
  AOI21_X1 U5102 ( .B1(n4452), .B2(n4896), .A(n4451), .ZN(n4453) );
  OAI211_X1 U5103 ( .C1(n4681), .C2(n4643), .A(n4454), .B(n4453), .ZN(U3263)
         );
  XOR2_X1 U5104 ( .A(n4460), .B(n4455), .Z(n4685) );
  INV_X1 U5105 ( .A(n4685), .ZN(n4474) );
  INV_X1 U5106 ( .A(n4477), .ZN(n4458) );
  OAI21_X1 U5107 ( .B1(n4458), .B2(n4457), .A(n4456), .ZN(n4459) );
  XOR2_X1 U5108 ( .A(n4460), .B(n4459), .Z(n4465) );
  OAI22_X1 U5109 ( .A1(n4461), .A2(n4647), .B1(n4467), .B2(n4645), .ZN(n4462)
         );
  AOI21_X1 U5110 ( .B1(n4463), .B2(n4660), .A(n4462), .ZN(n4464) );
  OAI21_X1 U5111 ( .B1(n4465), .B2(n4655), .A(n4464), .ZN(n4684) );
  INV_X1 U5112 ( .A(n4486), .ZN(n4468) );
  OAI21_X1 U5113 ( .B1(n4468), .B2(n4467), .A(n2417), .ZN(n4753) );
  NOR2_X1 U5114 ( .A1(n4753), .A2(n4600), .ZN(n4472) );
  OAI22_X1 U5115 ( .A1(n4470), .A2(n4665), .B1(n4469), .B2(n4668), .ZN(n4471)
         );
  AOI211_X1 U5116 ( .C1(n4684), .C2(n4668), .A(n4472), .B(n4471), .ZN(n4473)
         );
  OAI21_X1 U5117 ( .B1(n4474), .B2(n4603), .A(n4473), .ZN(U3264) );
  XNOR2_X1 U5118 ( .A(n4475), .B(n4478), .ZN(n4689) );
  INV_X1 U5119 ( .A(n4689), .ZN(n4493) );
  NAND2_X1 U5120 ( .A1(n4477), .A2(n4476), .ZN(n4479) );
  XNOR2_X1 U5121 ( .A(n4479), .B(n4478), .ZN(n4484) );
  OAI22_X1 U5122 ( .A1(n4480), .A2(n4647), .B1(n4487), .B2(n4645), .ZN(n4481)
         );
  AOI21_X1 U5123 ( .B1(n4482), .B2(n4660), .A(n4481), .ZN(n4483) );
  OAI21_X1 U5124 ( .B1(n4484), .B2(n4655), .A(n4483), .ZN(n4688) );
  INV_X1 U5125 ( .A(n4485), .ZN(n4488) );
  OAI21_X1 U5126 ( .B1(n4488), .B2(n4487), .A(n4486), .ZN(n4757) );
  AOI22_X1 U5127 ( .A1(n4489), .A2(n4912), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4643), .ZN(n4490) );
  OAI21_X1 U5128 ( .B1(n4757), .B2(n4600), .A(n4490), .ZN(n4491) );
  AOI21_X1 U5129 ( .B1(n4688), .B2(n4668), .A(n4491), .ZN(n4492) );
  OAI21_X1 U5130 ( .B1(n4493), .B2(n4603), .A(n4492), .ZN(U3265) );
  XNOR2_X1 U5131 ( .A(n4494), .B(n4496), .ZN(n4693) );
  INV_X1 U5132 ( .A(n4693), .ZN(n4508) );
  XOR2_X1 U5133 ( .A(n4496), .B(n4495), .Z(n4500) );
  OAI22_X1 U5134 ( .A1(n4536), .A2(n4647), .B1(n4502), .B2(n4645), .ZN(n4497)
         );
  AOI21_X1 U5135 ( .B1(n4498), .B2(n4660), .A(n4497), .ZN(n4499) );
  OAI21_X1 U5136 ( .B1(n4500), .B2(n4655), .A(n4499), .ZN(n4692) );
  OAI21_X1 U5137 ( .B1(n4501), .B2(n4502), .A(n4485), .ZN(n4761) );
  NOR2_X1 U5138 ( .A1(n4761), .A2(n4600), .ZN(n4506) );
  OAI22_X1 U5139 ( .A1(n4504), .A2(n4665), .B1(n4503), .B2(n4668), .ZN(n4505)
         );
  AOI211_X1 U5140 ( .C1(n4692), .C2(n4668), .A(n4506), .B(n4505), .ZN(n4507)
         );
  OAI21_X1 U5141 ( .B1(n4508), .B2(n4603), .A(n4507), .ZN(U3266) );
  XOR2_X1 U5142 ( .A(n4514), .B(n4509), .Z(n4697) );
  INV_X1 U5143 ( .A(n4697), .ZN(n4529) );
  OR2_X1 U5144 ( .A1(n4548), .A2(n4510), .ZN(n4512) );
  OAI21_X1 U5145 ( .B1(n4533), .B2(n4532), .A(n4513), .ZN(n4515) );
  XNOR2_X1 U5146 ( .A(n4515), .B(n4514), .ZN(n4520) );
  OAI22_X1 U5147 ( .A1(n4516), .A2(n4647), .B1(n4645), .B2(n4523), .ZN(n4517)
         );
  AOI21_X1 U5148 ( .B1(n4660), .B2(n4518), .A(n4517), .ZN(n4519) );
  OAI21_X1 U5149 ( .B1(n4520), .B2(n4655), .A(n4519), .ZN(n4696) );
  INV_X1 U5150 ( .A(n4521), .ZN(n4524) );
  INV_X1 U5151 ( .A(n4501), .ZN(n4522) );
  OAI21_X1 U5152 ( .B1(n4524), .B2(n4523), .A(n4522), .ZN(n4765) );
  AOI22_X1 U5153 ( .A1(n4525), .A2(n4912), .B1(REG2_REG_23__SCAN_IN), .B2(
        n4643), .ZN(n4526) );
  OAI21_X1 U5154 ( .B1(n4765), .B2(n4600), .A(n4526), .ZN(n4527) );
  AOI21_X1 U5155 ( .B1(n4696), .B2(n4668), .A(n4527), .ZN(n4528) );
  OAI21_X1 U5156 ( .B1(n4529), .B2(n4603), .A(n4528), .ZN(U3267) );
  OAI21_X1 U5157 ( .B1(n4531), .B2(n4532), .A(n4530), .ZN(n4703) );
  XNOR2_X1 U5158 ( .A(n4533), .B(n4532), .ZN(n4538) );
  AOI22_X1 U5159 ( .A1(n4534), .A2(n4630), .B1(n4542), .B2(n4568), .ZN(n4535)
         );
  OAI21_X1 U5160 ( .B1(n4536), .B2(n4908), .A(n4535), .ZN(n4537) );
  AOI21_X1 U5161 ( .B1(n4538), .B2(n4906), .A(n4537), .ZN(n4702) );
  NOR2_X1 U5162 ( .A1(n4668), .A2(n4539), .ZN(n4540) );
  AOI21_X1 U5163 ( .B1(n4541), .B2(n4912), .A(n4540), .ZN(n4544) );
  NAND2_X1 U5164 ( .A1(n4556), .A2(n4542), .ZN(n4700) );
  NAND3_X1 U5165 ( .A1(n4521), .A2(n4896), .A3(n4700), .ZN(n4543) );
  OAI211_X1 U5166 ( .C1(n4702), .C2(n4643), .A(n4544), .B(n4543), .ZN(n4545)
         );
  INV_X1 U5167 ( .A(n4545), .ZN(n4546) );
  OAI21_X1 U5168 ( .B1(n4703), .B2(n4603), .A(n4546), .ZN(U3268) );
  XNOR2_X1 U5169 ( .A(n4547), .B(n4549), .ZN(n4705) );
  INV_X1 U5170 ( .A(n4705), .ZN(n4563) );
  XOR2_X1 U5171 ( .A(n4549), .B(n4548), .Z(n4554) );
  OAI22_X1 U5172 ( .A1(n4550), .A2(n4647), .B1(n4645), .B2(n4557), .ZN(n4551)
         );
  AOI21_X1 U5173 ( .B1(n4552), .B2(n4660), .A(n4551), .ZN(n4553) );
  OAI21_X1 U5174 ( .B1(n4554), .B2(n4655), .A(n4553), .ZN(n4704) );
  INV_X1 U5175 ( .A(n4555), .ZN(n4558) );
  OAI21_X1 U5176 ( .B1(n4558), .B2(n4557), .A(n4556), .ZN(n4770) );
  NOR2_X1 U5177 ( .A1(n4770), .A2(n4600), .ZN(n4561) );
  OAI22_X1 U5178 ( .A1(n4559), .A2(n4665), .B1(n4043), .B2(n4668), .ZN(n4560)
         );
  AOI211_X1 U5179 ( .C1(n4704), .C2(n4668), .A(n4561), .B(n4560), .ZN(n4562)
         );
  OAI21_X1 U5180 ( .B1(n4563), .B2(n4603), .A(n4562), .ZN(U3269) );
  INV_X1 U5181 ( .A(n4571), .ZN(n4567) );
  NOR2_X1 U5182 ( .A1(n4565), .A2(n4564), .ZN(n4566) );
  XOR2_X1 U5183 ( .A(n4567), .B(n4566), .Z(n4575) );
  AOI22_X1 U5184 ( .A1(n4610), .A2(n4630), .B1(n4577), .B2(n4568), .ZN(n4569)
         );
  OAI21_X1 U5185 ( .B1(n4570), .B2(n4908), .A(n4569), .ZN(n4574) );
  XNOR2_X1 U5186 ( .A(n4572), .B(n4571), .ZN(n4711) );
  NOR2_X1 U5187 ( .A1(n4711), .A2(n4905), .ZN(n4573) );
  AOI211_X1 U5188 ( .C1(n4906), .C2(n4575), .A(n4574), .B(n4573), .ZN(n4710)
         );
  INV_X1 U5189 ( .A(n4711), .ZN(n4582) );
  INV_X1 U5190 ( .A(n4576), .ZN(n4596) );
  NAND2_X1 U5191 ( .A1(n4596), .A2(n4577), .ZN(n4708) );
  AND3_X1 U5192 ( .A1(n4708), .A2(n4896), .A3(n4555), .ZN(n4581) );
  OAI22_X1 U5193 ( .A1(n4579), .A2(n4665), .B1(n4578), .B2(n4668), .ZN(n4580)
         );
  AOI211_X1 U5194 ( .C1(n4582), .C2(n4913), .A(n4581), .B(n4580), .ZN(n4583)
         );
  OAI21_X1 U5195 ( .B1(n4710), .B2(n4643), .A(n4583), .ZN(U3270) );
  XOR2_X1 U5196 ( .A(n4590), .B(n4584), .Z(n4713) );
  INV_X1 U5197 ( .A(n4713), .ZN(n4604) );
  OAI21_X1 U5198 ( .B1(n4625), .B2(n4586), .A(n4585), .ZN(n4606) );
  INV_X1 U5199 ( .A(n4587), .ZN(n4589) );
  OAI21_X1 U5200 ( .B1(n4606), .B2(n4589), .A(n4588), .ZN(n4591) );
  XNOR2_X1 U5201 ( .A(n4591), .B(n4590), .ZN(n4595) );
  OAI22_X1 U5202 ( .A1(n4624), .A2(n4647), .B1(n4597), .B2(n4645), .ZN(n4592)
         );
  AOI21_X1 U5203 ( .B1(n4593), .B2(n4660), .A(n4592), .ZN(n4594) );
  OAI21_X1 U5204 ( .B1(n4595), .B2(n4655), .A(n4594), .ZN(n4712) );
  OAI21_X1 U5205 ( .B1(n4614), .B2(n4597), .A(n4596), .ZN(n4775) );
  AOI22_X1 U5206 ( .A1(n4598), .A2(n4912), .B1(n4643), .B2(
        REG2_REG_19__SCAN_IN), .ZN(n4599) );
  OAI21_X1 U5207 ( .B1(n4775), .B2(n4600), .A(n4599), .ZN(n4601) );
  AOI21_X1 U5208 ( .B1(n4712), .B2(n4668), .A(n4601), .ZN(n4602) );
  OAI21_X1 U5209 ( .B1(n4604), .B2(n4603), .A(n4602), .ZN(U3271) );
  OAI22_X1 U5210 ( .A1(n4605), .A2(n4647), .B1(n4616), .B2(n4645), .ZN(n4609)
         );
  XNOR2_X1 U5211 ( .A(n4606), .B(n4612), .ZN(n4607) );
  NOR2_X1 U5212 ( .A1(n4607), .A2(n4655), .ZN(n4608) );
  AOI211_X1 U5213 ( .C1(n4660), .C2(n4610), .A(n4609), .B(n4608), .ZN(n4718)
         );
  OAI21_X1 U5214 ( .B1(n4613), .B2(n4612), .A(n4611), .ZN(n4716) );
  INV_X1 U5215 ( .A(n4631), .ZN(n4617) );
  INV_X1 U5216 ( .A(n4614), .ZN(n4615) );
  OAI211_X1 U5217 ( .C1(n4617), .C2(n4616), .A(n4615), .B(n4972), .ZN(n4717)
         );
  INV_X1 U5218 ( .A(n4618), .ZN(n4619) );
  NOR2_X1 U5219 ( .A1(n4717), .A2(n4619), .ZN(n4622) );
  OAI22_X1 U5220 ( .A1(n4088), .A2(n4668), .B1(n4620), .B2(n4665), .ZN(n4621)
         );
  AOI211_X1 U5221 ( .C1(n4716), .C2(n4640), .A(n4622), .B(n4621), .ZN(n4623)
         );
  OAI21_X1 U5222 ( .B1(n4718), .B2(n4643), .A(n4623), .ZN(U3272) );
  OAI22_X1 U5223 ( .A1(n4624), .A2(n4908), .B1(n4645), .B2(n4632), .ZN(n4628)
         );
  XOR2_X1 U5224 ( .A(n4639), .B(n4625), .Z(n4626) );
  NOR2_X1 U5225 ( .A1(n4626), .A2(n4655), .ZN(n4627) );
  AOI211_X1 U5226 ( .C1(n4630), .C2(n4629), .A(n4628), .B(n4627), .ZN(n4720)
         );
  OAI21_X1 U5227 ( .B1(n4633), .B2(n4632), .A(n4631), .ZN(n4781) );
  INV_X1 U5228 ( .A(n4781), .ZN(n4637) );
  OAI22_X1 U5229 ( .A1(n4668), .A2(n4635), .B1(n4634), .B2(n4665), .ZN(n4636)
         );
  AOI21_X1 U5230 ( .B1(n4637), .B2(n4896), .A(n4636), .ZN(n4642) );
  XOR2_X1 U5231 ( .A(n4639), .B(n4638), .Z(n4722) );
  NAND2_X1 U5232 ( .A1(n4722), .A2(n4640), .ZN(n4641) );
  OAI211_X1 U5233 ( .C1(n4720), .C2(n4643), .A(n4642), .B(n4641), .ZN(U3273)
         );
  XOR2_X1 U5234 ( .A(n4653), .B(n4644), .Z(n4733) );
  OAI22_X1 U5235 ( .A1(n4648), .A2(n4647), .B1(n4646), .B2(n4645), .ZN(n4658)
         );
  INV_X1 U5236 ( .A(n4649), .ZN(n4650) );
  AOI21_X1 U5237 ( .B1(n4652), .B2(n4651), .A(n4650), .ZN(n4654) );
  XNOR2_X1 U5238 ( .A(n4654), .B(n4653), .ZN(n4656) );
  NOR2_X1 U5239 ( .A1(n4656), .A2(n4655), .ZN(n4657) );
  AOI211_X1 U5240 ( .C1(n4660), .C2(n4659), .A(n4658), .B(n4657), .ZN(n4661)
         );
  OAI21_X1 U5241 ( .B1(n4733), .B2(n4905), .A(n4661), .ZN(n4734) );
  NAND2_X1 U5242 ( .A1(n4734), .A2(n4668), .ZN(n4672) );
  NAND2_X1 U5243 ( .A1(n3598), .A2(n4662), .ZN(n4663) );
  NAND2_X1 U5244 ( .A1(n4664), .A2(n4663), .ZN(n4788) );
  INV_X1 U5245 ( .A(n4788), .ZN(n4670) );
  OAI22_X1 U5246 ( .A1(n4668), .A2(n4667), .B1(n4666), .B2(n4665), .ZN(n4669)
         );
  AOI21_X1 U5247 ( .B1(n4670), .B2(n4896), .A(n4669), .ZN(n4671) );
  OAI211_X1 U5248 ( .C1(n4733), .C2(n4673), .A(n4672), .B(n4671), .ZN(U3277)
         );
  NAND2_X1 U5249 ( .A1(n4994), .A2(n4739), .ZN(n4675) );
  NAND2_X1 U5250 ( .A1(n4991), .A2(REG1_REG_31__SCAN_IN), .ZN(n4674) );
  OAI211_X1 U5251 ( .C1(n4742), .C2(n4738), .A(n4675), .B(n4674), .ZN(U3549)
         );
  INV_X1 U5252 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4679) );
  NAND2_X1 U5253 ( .A1(n4744), .A2(n4676), .ZN(n4678) );
  NAND2_X1 U5254 ( .A1(n4994), .A2(n4745), .ZN(n4677) );
  OAI211_X1 U5255 ( .C1(n4994), .C2(n4679), .A(n4678), .B(n4677), .ZN(U3548)
         );
  INV_X1 U5256 ( .A(n4972), .ZN(n4949) );
  NAND2_X1 U5257 ( .A1(n4680), .A2(n4975), .ZN(n4682) );
  OAI211_X1 U5258 ( .C1(n4949), .C2(n4683), .A(n4682), .B(n4681), .ZN(n4749)
         );
  MUX2_X1 U5259 ( .A(REG1_REG_27__SCAN_IN), .B(n4749), .S(n4994), .Z(U3545) );
  INV_X1 U5260 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4686) );
  AOI21_X1 U5261 ( .B1(n4685), .B2(n4975), .A(n4684), .ZN(n4750) );
  MUX2_X1 U5262 ( .A(n4686), .B(n4750), .S(n4994), .Z(n4687) );
  OAI21_X1 U5263 ( .B1(n4738), .B2(n4753), .A(n4687), .ZN(U3544) );
  AOI21_X1 U5264 ( .B1(n4689), .B2(n4975), .A(n4688), .ZN(n4754) );
  MUX2_X1 U5265 ( .A(n4690), .B(n4754), .S(n4994), .Z(n4691) );
  OAI21_X1 U5266 ( .B1(n4738), .B2(n4757), .A(n4691), .ZN(U3543) );
  AOI21_X1 U5267 ( .B1(n4693), .B2(n4975), .A(n4692), .ZN(n4758) );
  MUX2_X1 U5268 ( .A(n4694), .B(n4758), .S(n4994), .Z(n4695) );
  OAI21_X1 U5269 ( .B1(n4738), .B2(n4761), .A(n4695), .ZN(U3542) );
  AOI21_X1 U5270 ( .B1(n4697), .B2(n4975), .A(n4696), .ZN(n4762) );
  MUX2_X1 U5271 ( .A(n4698), .B(n4762), .S(n4994), .Z(n4699) );
  OAI21_X1 U5272 ( .B1(n4738), .B2(n4765), .A(n4699), .ZN(U3541) );
  NAND3_X1 U5273 ( .A1(n4521), .A2(n4972), .A3(n4700), .ZN(n4701) );
  OAI211_X1 U5274 ( .C1(n4703), .C2(n4967), .A(n4702), .B(n4701), .ZN(n4766)
         );
  MUX2_X1 U5275 ( .A(REG1_REG_22__SCAN_IN), .B(n4766), .S(n4994), .Z(U3540) );
  AOI21_X1 U5276 ( .B1(n4705), .B2(n4975), .A(n4704), .ZN(n4767) );
  MUX2_X1 U5277 ( .A(n4706), .B(n4767), .S(n4994), .Z(n4707) );
  OAI21_X1 U5278 ( .B1(n4738), .B2(n4770), .A(n4707), .ZN(U3539) );
  NAND3_X1 U5279 ( .A1(n4708), .A2(n4972), .A3(n4555), .ZN(n4709) );
  OAI211_X1 U5280 ( .C1(n4711), .C2(n4954), .A(n4710), .B(n4709), .ZN(n4771)
         );
  MUX2_X1 U5281 ( .A(REG1_REG_20__SCAN_IN), .B(n4771), .S(n4994), .Z(U3538) );
  INV_X1 U5282 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4714) );
  AOI21_X1 U5283 ( .B1(n4713), .B2(n4975), .A(n4712), .ZN(n4772) );
  MUX2_X1 U5284 ( .A(n4714), .B(n4772), .S(n4994), .Z(n4715) );
  OAI21_X1 U5285 ( .B1(n4738), .B2(n4775), .A(n4715), .ZN(U3537) );
  INV_X1 U5286 ( .A(n4716), .ZN(n4719) );
  OAI211_X1 U5287 ( .C1(n4967), .C2(n4719), .A(n4718), .B(n4717), .ZN(n4776)
         );
  MUX2_X1 U5288 ( .A(REG1_REG_18__SCAN_IN), .B(n4776), .S(n4994), .Z(U3536) );
  INV_X1 U5289 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4723) );
  INV_X1 U5290 ( .A(n4720), .ZN(n4721) );
  AOI21_X1 U5291 ( .B1(n4722), .B2(n4975), .A(n4721), .ZN(n4778) );
  MUX2_X1 U5292 ( .A(n4723), .B(n4778), .S(n4994), .Z(n4724) );
  OAI21_X1 U5293 ( .B1(n4738), .B2(n4781), .A(n4724), .ZN(U3535) );
  AOI21_X1 U5294 ( .B1(n4972), .B2(n4726), .A(n4725), .ZN(n4727) );
  OAI21_X1 U5295 ( .B1(n4728), .B2(n4967), .A(n4727), .ZN(n4782) );
  MUX2_X1 U5296 ( .A(REG1_REG_16__SCAN_IN), .B(n4782), .S(n4994), .Z(U3534) );
  AOI21_X1 U5297 ( .B1(n4972), .B2(n4730), .A(n4729), .ZN(n4731) );
  OAI21_X1 U5298 ( .B1(n4732), .B2(n4967), .A(n4731), .ZN(n4783) );
  MUX2_X1 U5299 ( .A(REG1_REG_15__SCAN_IN), .B(n4783), .S(n4994), .Z(U3533) );
  INV_X1 U5300 ( .A(n4733), .ZN(n4735) );
  AOI21_X1 U5301 ( .B1(n4963), .B2(n4735), .A(n4734), .ZN(n4784) );
  MUX2_X1 U5302 ( .A(n4736), .B(n4784), .S(n4994), .Z(n4737) );
  OAI21_X1 U5303 ( .B1(n4738), .B2(n4788), .A(n4737), .ZN(U3531) );
  NAND2_X1 U5304 ( .A1(n4777), .A2(n4739), .ZN(n4741) );
  NAND2_X1 U5305 ( .A1(n4980), .A2(REG0_REG_31__SCAN_IN), .ZN(n4740) );
  OAI211_X1 U5306 ( .C1(n4742), .C2(n4787), .A(n4741), .B(n4740), .ZN(U3517)
         );
  INV_X1 U5307 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4748) );
  NAND2_X1 U5308 ( .A1(n4744), .A2(n4743), .ZN(n4747) );
  NAND2_X1 U5309 ( .A1(n4777), .A2(n4745), .ZN(n4746) );
  OAI211_X1 U5310 ( .C1(n4777), .C2(n4748), .A(n4747), .B(n4746), .ZN(U3516)
         );
  MUX2_X1 U5311 ( .A(REG0_REG_27__SCAN_IN), .B(n4749), .S(n4777), .Z(U3513) );
  INV_X1 U5312 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4751) );
  MUX2_X1 U5313 ( .A(n4751), .B(n4750), .S(n4777), .Z(n4752) );
  OAI21_X1 U5314 ( .B1(n4753), .B2(n4787), .A(n4752), .ZN(U3512) );
  MUX2_X1 U5315 ( .A(n4755), .B(n4754), .S(n4777), .Z(n4756) );
  OAI21_X1 U5316 ( .B1(n4757), .B2(n4787), .A(n4756), .ZN(U3511) );
  INV_X1 U5317 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4759) );
  MUX2_X1 U5318 ( .A(n4759), .B(n4758), .S(n4777), .Z(n4760) );
  OAI21_X1 U5319 ( .B1(n4761), .B2(n4787), .A(n4760), .ZN(U3510) );
  INV_X1 U5320 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4763) );
  MUX2_X1 U5321 ( .A(n4763), .B(n4762), .S(n4777), .Z(n4764) );
  OAI21_X1 U5322 ( .B1(n4765), .B2(n4787), .A(n4764), .ZN(U3509) );
  MUX2_X1 U5323 ( .A(REG0_REG_22__SCAN_IN), .B(n4766), .S(n4777), .Z(U3508) );
  MUX2_X1 U5324 ( .A(n4768), .B(n4767), .S(n4777), .Z(n4769) );
  OAI21_X1 U5325 ( .B1(n4770), .B2(n4787), .A(n4769), .ZN(U3507) );
  MUX2_X1 U5326 ( .A(REG0_REG_20__SCAN_IN), .B(n4771), .S(n4777), .Z(U3506) );
  MUX2_X1 U5327 ( .A(n4773), .B(n4772), .S(n4777), .Z(n4774) );
  OAI21_X1 U5328 ( .B1(n4775), .B2(n4787), .A(n4774), .ZN(U3505) );
  MUX2_X1 U5329 ( .A(REG0_REG_18__SCAN_IN), .B(n4776), .S(n4777), .Z(U3503) );
  INV_X1 U5330 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4779) );
  MUX2_X1 U5331 ( .A(n4779), .B(n4778), .S(n4777), .Z(n4780) );
  OAI21_X1 U5332 ( .B1(n4781), .B2(n4787), .A(n4780), .ZN(U3501) );
  MUX2_X1 U5333 ( .A(REG0_REG_16__SCAN_IN), .B(n4782), .S(n4777), .Z(U3499) );
  MUX2_X1 U5334 ( .A(REG0_REG_15__SCAN_IN), .B(n4783), .S(n4777), .Z(U3497) );
  MUX2_X1 U5335 ( .A(n4785), .B(n4784), .S(n4777), .Z(n4786) );
  OAI21_X1 U5336 ( .B1(n4788), .B2(n4787), .A(n4786), .ZN(U3493) );
  MUX2_X1 U5337 ( .A(DATAI_30_), .B(n4789), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U5338 ( .A(n4790), .B(DATAI_28_), .S(U3149), .Z(U3324) );
  MUX2_X1 U5339 ( .A(n4791), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5340 ( .A(DATAI_22_), .B(n4792), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U5341 ( .A(DATAI_20_), .B(n4793), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5342 ( .A(n4802), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5343 ( .A(n4803), .B(DATAI_17_), .S(U3149), .Z(U3335) );
  MUX2_X1 U5344 ( .A(DATAI_12_), .B(n4794), .S(STATE_REG_SCAN_IN), .Z(U3340)
         );
  MUX2_X1 U5345 ( .A(DATAI_11_), .B(n4795), .S(STATE_REG_SCAN_IN), .Z(U3341)
         );
  MUX2_X1 U5346 ( .A(n3438), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U5347 ( .A(n3432), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5348 ( .A(DATAI_5_), .B(n4796), .S(STATE_REG_SCAN_IN), .Z(U3347) );
  MUX2_X1 U5349 ( .A(DATAI_4_), .B(n4820), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5350 ( .A(n2130), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5351 ( .A(n4798), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  NAND2_X1 U5352 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4807), .ZN(n4799) );
  OAI21_X1 U5353 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4807), .A(n4799), .ZN(n4879) );
  NAND2_X1 U5354 ( .A1(n4391), .A2(n4635), .ZN(n4800) );
  NAND2_X1 U5355 ( .A1(n4391), .A2(n4723), .ZN(n4804) );
  INV_X1 U5356 ( .A(n4807), .ZN(n4934) );
  AOI22_X1 U5357 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4934), .B1(n4807), .B2(
        n4806), .ZN(n4889) );
  XNOR2_X1 U5358 ( .A(n4809), .B(n2425), .ZN(n4814) );
  AOI21_X1 U5359 ( .B1(n4881), .B2(ADDR_REG_19__SCAN_IN), .A(n4810), .ZN(n4811) );
  OAI21_X1 U5360 ( .B1(n4892), .B2(n4812), .A(n4811), .ZN(n4813) );
  OAI21_X1 U5361 ( .B1(n4816), .B2(n4878), .A(n4815), .ZN(U3259) );
  NAND2_X1 U5362 ( .A1(n4873), .A2(n4817), .ZN(n4826) );
  XNOR2_X1 U5363 ( .A(n4818), .B(n2294), .ZN(n4819) );
  NAND2_X1 U5364 ( .A1(n4875), .A2(n4819), .ZN(n4825) );
  NAND2_X1 U5365 ( .A1(n4849), .A2(n4820), .ZN(n4824) );
  INV_X1 U5366 ( .A(n4821), .ZN(n4822) );
  AOI21_X1 U5367 ( .B1(n4881), .B2(ADDR_REG_4__SCAN_IN), .A(n4822), .ZN(n4823)
         );
  AND4_X1 U5368 ( .A1(n4826), .A2(n4825), .A3(n4824), .A4(n4823), .ZN(n4828)
         );
  NAND2_X1 U5369 ( .A1(n4828), .A2(n4827), .ZN(U3244) );
  INV_X1 U5370 ( .A(n4829), .ZN(n4831) );
  AOI211_X1 U5371 ( .C1(n4831), .C2(n4830), .A(n2164), .B(n4887), .ZN(n4832)
         );
  AOI211_X1 U5372 ( .C1(n4881), .C2(ADDR_REG_13__SCAN_IN), .A(n4833), .B(n4832), .ZN(n4839) );
  AOI21_X1 U5373 ( .B1(n4667), .B2(n4840), .A(n4834), .ZN(n4837) );
  AOI21_X1 U5374 ( .B1(n4837), .B2(n4835), .A(n4878), .ZN(n4836) );
  OAI21_X1 U5375 ( .B1(n4837), .B2(n4835), .A(n4836), .ZN(n4838) );
  OAI211_X1 U5376 ( .C1(n4892), .C2(n4840), .A(n4839), .B(n4838), .ZN(U3253)
         );
  NAND2_X1 U5377 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4881), .ZN(n4852) );
  AOI211_X1 U5378 ( .C1(n4843), .C2(n4842), .A(n4841), .B(n4887), .ZN(n4848)
         );
  AOI211_X1 U5379 ( .C1(n4846), .C2(n4845), .A(n4844), .B(n4878), .ZN(n4847)
         );
  AOI211_X1 U5380 ( .C1(n4849), .C2(n4939), .A(n4848), .B(n4847), .ZN(n4851)
         );
  NAND3_X1 U5381 ( .A1(n4852), .A2(n4851), .A3(n4850), .ZN(U3254) );
  AOI211_X1 U5382 ( .C1(n4855), .C2(n4854), .A(n4853), .B(n4878), .ZN(n4856)
         );
  AOI211_X1 U5383 ( .C1(n4881), .C2(ADDR_REG_15__SCAN_IN), .A(n4857), .B(n4856), .ZN(n4862) );
  AOI21_X1 U5384 ( .B1(n4859), .B2(n2152), .A(n4858), .ZN(n4860) );
  NAND2_X1 U5385 ( .A1(n4873), .A2(n4860), .ZN(n4861) );
  OAI211_X1 U5386 ( .C1(n4892), .C2(n4863), .A(n4862), .B(n4861), .ZN(U3255)
         );
  INV_X1 U5387 ( .A(n4864), .ZN(n4865) );
  AOI21_X1 U5388 ( .B1(n4881), .B2(ADDR_REG_16__SCAN_IN), .A(n4865), .ZN(n4877) );
  OAI21_X1 U5389 ( .B1(n4868), .B2(n4867), .A(n4866), .ZN(n4874) );
  OAI21_X1 U5390 ( .B1(n4871), .B2(n4870), .A(n4869), .ZN(n4872) );
  AOI22_X1 U5391 ( .A1(n4875), .A2(n4874), .B1(n4873), .B2(n4872), .ZN(n4876)
         );
  OAI211_X1 U5392 ( .C1(n4936), .C2(n4892), .A(n4877), .B(n4876), .ZN(U3256)
         );
  NAND2_X1 U5393 ( .A1(n4881), .A2(ADDR_REG_18__SCAN_IN), .ZN(n4884) );
  OAI211_X1 U5394 ( .C1(n4892), .C2(n4934), .A(n4891), .B(n4890), .ZN(U3258)
         );
  AOI22_X1 U5395 ( .A1(REG3_REG_2__SCAN_IN), .A2(n4912), .B1(
        REG2_REG_2__SCAN_IN), .B2(n4643), .ZN(n4899) );
  INV_X1 U5396 ( .A(n4893), .ZN(n4897) );
  INV_X1 U5397 ( .A(n4894), .ZN(n4895) );
  AOI22_X1 U5398 ( .A1(n4897), .A2(n4913), .B1(n4896), .B2(n4895), .ZN(n4898)
         );
  OAI211_X1 U5399 ( .C1(n4643), .C2(n4900), .A(n4899), .B(n4898), .ZN(U3288)
         );
  INV_X1 U5400 ( .A(n4901), .ZN(n4902) );
  NOR2_X1 U5401 ( .A1(n4903), .A2(n4902), .ZN(n4945) );
  INV_X1 U5402 ( .A(n4904), .ZN(n4910) );
  INV_X1 U5403 ( .A(n4905), .ZN(n4907) );
  NOR2_X1 U5404 ( .A1(n4907), .A2(n4906), .ZN(n4909) );
  OAI22_X1 U5405 ( .A1(n4911), .A2(n4909), .B1(n2885), .B2(n4908), .ZN(n4944)
         );
  AOI21_X1 U5406 ( .B1(n4945), .B2(n4910), .A(n4944), .ZN(n4916) );
  INV_X1 U5407 ( .A(n4911), .ZN(n4946) );
  AOI22_X1 U5408 ( .A1(n4913), .A2(n4946), .B1(REG3_REG_0__SCAN_IN), .B2(n4912), .ZN(n4914) );
  OAI221_X1 U5409 ( .B1(n4643), .B2(n4916), .C1(n4668), .C2(n4915), .A(n4914), 
        .ZN(U3290) );
  AND2_X1 U5410 ( .A1(D_REG_31__SCAN_IN), .A2(n4928), .ZN(U3291) );
  NOR2_X1 U5411 ( .A1(n4930), .A2(n4917), .ZN(U3292) );
  AND2_X1 U5412 ( .A1(D_REG_29__SCAN_IN), .A2(n4928), .ZN(U3293) );
  AND2_X1 U5413 ( .A1(D_REG_28__SCAN_IN), .A2(n4928), .ZN(U3294) );
  AND2_X1 U5414 ( .A1(D_REG_27__SCAN_IN), .A2(n4928), .ZN(U3295) );
  NOR2_X1 U5415 ( .A1(n4930), .A2(n4918), .ZN(U3296) );
  AND2_X1 U5416 ( .A1(D_REG_25__SCAN_IN), .A2(n4928), .ZN(U3297) );
  NOR2_X1 U5417 ( .A1(n4930), .A2(n4919), .ZN(U3298) );
  AND2_X1 U5418 ( .A1(D_REG_23__SCAN_IN), .A2(n4928), .ZN(U3299) );
  AND2_X1 U5419 ( .A1(D_REG_22__SCAN_IN), .A2(n4928), .ZN(U3300) );
  NOR2_X1 U5420 ( .A1(n4930), .A2(n4920), .ZN(U3301) );
  NOR2_X1 U5421 ( .A1(n4930), .A2(n4921), .ZN(U3302) );
  NOR2_X1 U5422 ( .A1(n4930), .A2(n4922), .ZN(U3303) );
  AND2_X1 U5423 ( .A1(D_REG_18__SCAN_IN), .A2(n4928), .ZN(U3304) );
  NOR2_X1 U5424 ( .A1(n4930), .A2(n4923), .ZN(U3305) );
  AND2_X1 U5425 ( .A1(D_REG_16__SCAN_IN), .A2(n4928), .ZN(U3306) );
  AND2_X1 U5426 ( .A1(D_REG_15__SCAN_IN), .A2(n4928), .ZN(U3307) );
  NOR2_X1 U5427 ( .A1(n4930), .A2(n4924), .ZN(U3308) );
  AND2_X1 U5428 ( .A1(D_REG_13__SCAN_IN), .A2(n4928), .ZN(U3309) );
  NOR2_X1 U5429 ( .A1(n4930), .A2(n4925), .ZN(U3310) );
  NOR2_X1 U5430 ( .A1(n4930), .A2(n4926), .ZN(U3311) );
  AND2_X1 U5431 ( .A1(D_REG_10__SCAN_IN), .A2(n4928), .ZN(U3312) );
  AND2_X1 U5432 ( .A1(D_REG_9__SCAN_IN), .A2(n4928), .ZN(U3313) );
  AND2_X1 U5433 ( .A1(D_REG_8__SCAN_IN), .A2(n4928), .ZN(U3314) );
  AND2_X1 U5434 ( .A1(D_REG_7__SCAN_IN), .A2(n4928), .ZN(U3315) );
  AND2_X1 U5435 ( .A1(D_REG_6__SCAN_IN), .A2(n4928), .ZN(U3316) );
  NOR2_X1 U5436 ( .A1(n4930), .A2(n4927), .ZN(U3317) );
  AND2_X1 U5437 ( .A1(D_REG_4__SCAN_IN), .A2(n4928), .ZN(U3318) );
  AND2_X1 U5438 ( .A1(D_REG_3__SCAN_IN), .A2(n4928), .ZN(U3319) );
  NOR2_X1 U5439 ( .A1(n4930), .A2(n4929), .ZN(U3320) );
  AOI21_X1 U5440 ( .B1(U3149), .B2(n4932), .A(n4931), .ZN(U3329) );
  INV_X1 U5441 ( .A(DATAI_18_), .ZN(n4933) );
  AOI22_X1 U5442 ( .A1(STATE_REG_SCAN_IN), .A2(n4934), .B1(n4933), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5443 ( .A1(STATE_REG_SCAN_IN), .A2(n4936), .B1(n4935), .B2(U3149), 
        .ZN(U3336) );
  OAI22_X1 U5444 ( .A1(U3149), .A2(n4937), .B1(DATAI_15_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4938) );
  INV_X1 U5445 ( .A(n4938), .ZN(U3337) );
  OAI22_X1 U5446 ( .A1(U3149), .A2(n4939), .B1(DATAI_14_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4940) );
  INV_X1 U5447 ( .A(n4940), .ZN(U3338) );
  OAI22_X1 U5448 ( .A1(U3149), .A2(n4941), .B1(DATAI_13_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4942) );
  INV_X1 U5449 ( .A(n4942), .ZN(U3339) );
  AOI22_X1 U5450 ( .A1(STATE_REG_SCAN_IN), .A2(n4943), .B1(n3855), .B2(U3149), 
        .ZN(U3352) );
  AOI211_X1 U5451 ( .C1(n4963), .C2(n4946), .A(n4945), .B(n4944), .ZN(n4983)
         );
  INV_X1 U5452 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4947) );
  AOI22_X1 U5453 ( .A1(n4777), .A2(n4983), .B1(n4947), .B2(n4980), .ZN(U3467)
         );
  OAI22_X1 U5454 ( .A1(n4950), .A2(n4954), .B1(n4949), .B2(n4948), .ZN(n4951)
         );
  NOR2_X1 U5455 ( .A1(n4952), .A2(n4951), .ZN(n4984) );
  INV_X1 U5456 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4953) );
  AOI22_X1 U5457 ( .A1(n4777), .A2(n4984), .B1(n4953), .B2(n4980), .ZN(U3469)
         );
  NOR2_X1 U5458 ( .A1(n4955), .A2(n4954), .ZN(n4957) );
  AOI211_X1 U5459 ( .C1(n4972), .C2(n4958), .A(n4957), .B(n4956), .ZN(n4986)
         );
  INV_X1 U5460 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4959) );
  AOI22_X1 U5461 ( .A1(n4777), .A2(n4986), .B1(n4959), .B2(n4980), .ZN(U3473)
         );
  INV_X1 U5462 ( .A(n4960), .ZN(n4962) );
  AOI211_X1 U5463 ( .C1(n4964), .C2(n4963), .A(n4962), .B(n4961), .ZN(n4988)
         );
  INV_X1 U5464 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4965) );
  AOI22_X1 U5465 ( .A1(n4777), .A2(n4988), .B1(n4965), .B2(n4980), .ZN(U3475)
         );
  INV_X1 U5466 ( .A(n4966), .ZN(n4970) );
  NOR2_X1 U5467 ( .A1(n4968), .A2(n4967), .ZN(n4969) );
  AOI211_X1 U5468 ( .C1(n4972), .C2(n4971), .A(n4970), .B(n4969), .ZN(n4990)
         );
  AOI22_X1 U5469 ( .A1(n4777), .A2(n4990), .B1(n4973), .B2(n4980), .ZN(U3477)
         );
  NAND3_X1 U5470 ( .A1(n4976), .A2(n4975), .A3(n4974), .ZN(n4977) );
  AND3_X1 U5471 ( .A1(n4979), .A2(n4978), .A3(n4977), .ZN(n4993) );
  INV_X1 U5472 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4981) );
  AOI22_X1 U5473 ( .A1(n4777), .A2(n4993), .B1(n4981), .B2(n4980), .ZN(U3481)
         );
  AOI22_X1 U5474 ( .A1(n4994), .A2(n4983), .B1(n4982), .B2(n4991), .ZN(U3518)
         );
  AOI22_X1 U5475 ( .A1(n4994), .A2(n4984), .B1(n3168), .B2(n4991), .ZN(U3519)
         );
  AOI22_X1 U5476 ( .A1(n4994), .A2(n4986), .B1(n4985), .B2(n4991), .ZN(U3521)
         );
  AOI22_X1 U5477 ( .A1(n4994), .A2(n4988), .B1(n4987), .B2(n4991), .ZN(U3522)
         );
  AOI22_X1 U5478 ( .A1(n4994), .A2(n4990), .B1(n4989), .B2(n4991), .ZN(U3523)
         );
  AOI22_X1 U5479 ( .A1(n4994), .A2(n4993), .B1(n4992), .B2(n4991), .ZN(U3525)
         );
  CLKBUF_X2 U2408 ( .A(n4177), .Z(n4178) );
  CLKBUF_X2 U2441 ( .A(n3164), .Z(n2130) );
endmodule

