

module b22_C_AntiSAT_k_256_3 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, SUB_1596_U4, SUB_1596_U62, 
        SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, 
        SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, 
        SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, 
        SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, 
        P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, 
        P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, 
        P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, 
        P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, 
        P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, 
        P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, 
        P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, 
        P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, 
        P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, 
        P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, 
        P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, 
        P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, 
        P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, 
        P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, 
        P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, 
        P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, 
        P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, 
        P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, 
        P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, 
        P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, 
        P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, 
        P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, 
        P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, 
        P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, 
        P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, 
        P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, 
        P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, 
        P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, 
        P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, 
        P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, 
        P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, 
        P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, 
        P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, 
        P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, 
        P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, 
        P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, 
        P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, 
        P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, 
        P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, 
        P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, 
        P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, 
        P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, 
        P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, 
        P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, 
        P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, 
        P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, 
        P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, 
        P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, 
        P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, 
        P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, 
        P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, 
        P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, 
        P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, 
        P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, 
        P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, 
        P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, 
        P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, 
        P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, 
        P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, 
        P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, 
        P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, 
        P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, 
        P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, 
        P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, 
        P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, 
        P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, 
        P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, 
        P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, 
        P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, 
        P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, 
        P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, 
        P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, 
        P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, 
        P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, 
        P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, 
        P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, 
        P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, 
        P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127,
         keyinput128, keyinput129, keyinput130, keyinput131, keyinput132,
         keyinput133, keyinput134, keyinput135, keyinput136, keyinput137,
         keyinput138, keyinput139, keyinput140, keyinput141, keyinput142,
         keyinput143, keyinput144, keyinput145, keyinput146, keyinput147,
         keyinput148, keyinput149, keyinput150, keyinput151, keyinput152,
         keyinput153, keyinput154, keyinput155, keyinput156, keyinput157,
         keyinput158, keyinput159, keyinput160, keyinput161, keyinput162,
         keyinput163, keyinput164, keyinput165, keyinput166, keyinput167,
         keyinput168, keyinput169, keyinput170, keyinput171, keyinput172,
         keyinput173, keyinput174, keyinput175, keyinput176, keyinput177,
         keyinput178, keyinput179, keyinput180, keyinput181, keyinput182,
         keyinput183, keyinput184, keyinput185, keyinput186, keyinput187,
         keyinput188, keyinput189, keyinput190, keyinput191, keyinput192,
         keyinput193, keyinput194, keyinput195, keyinput196, keyinput197,
         keyinput198, keyinput199, keyinput200, keyinput201, keyinput202,
         keyinput203, keyinput204, keyinput205, keyinput206, keyinput207,
         keyinput208, keyinput209, keyinput210, keyinput211, keyinput212,
         keyinput213, keyinput214, keyinput215, keyinput216, keyinput217,
         keyinput218, keyinput219, keyinput220, keyinput221, keyinput222,
         keyinput223, keyinput224, keyinput225, keyinput226, keyinput227,
         keyinput228, keyinput229, keyinput230, keyinput231, keyinput232,
         keyinput233, keyinput234, keyinput235, keyinput236, keyinput237,
         keyinput238, keyinput239, keyinput240, keyinput241, keyinput242,
         keyinput243, keyinput244, keyinput245, keyinput246, keyinput247,
         keyinput248, keyinput249, keyinput250, keyinput251, keyinput252,
         keyinput253, keyinput254, keyinput255;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526;

  NAND2_X1 U7367 ( .A1(n7044), .A2(n7045), .ZN(n14321) );
  OR2_X1 U7369 ( .A1(n13431), .A2(n13334), .ZN(n13320) );
  AND2_X1 U7370 ( .A1(n12964), .A2(n8669), .ZN(n13036) );
  CLKBUF_X3 U7371 ( .A(n7589), .Z(n7810) );
  AND2_X2 U7372 ( .A1(n10343), .A2(n10344), .ZN(n10603) );
  NAND2_X1 U7373 ( .A1(n7438), .A2(n7437), .ZN(n12505) );
  INV_X1 U7374 ( .A(n11983), .ZN(n6770) );
  NAND2_X2 U7375 ( .A1(n8074), .A2(n8075), .ZN(n7585) );
  AND2_X1 U7376 ( .A1(n9403), .A2(n9402), .ZN(n10959) );
  INV_X1 U7377 ( .A(n8797), .ZN(n9028) );
  BUF_X2 U7378 ( .A(n8835), .Z(n6619) );
  NAND2_X1 U7379 ( .A1(n9719), .A2(n11201), .ZN(n10342) );
  INV_X2 U7380 ( .A(n8313), .ZN(n8797) );
  NAND2_X2 U7381 ( .A1(n10176), .A2(n7311), .ZN(n10046) );
  NAND2_X1 U7382 ( .A1(n8217), .A2(n8216), .ZN(n12214) );
  NOR2_X1 U7383 ( .A1(n8235), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n13476) );
  INV_X1 U7384 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8381) );
  NOR2_X1 U7386 ( .A1(n8201), .A2(n8200), .ZN(n8496) );
  XNOR2_X1 U7387 ( .A(n15060), .B(n15050), .ZN(n15041) );
  INV_X1 U7388 ( .A(n8457), .ZN(n9021) );
  INV_X2 U7389 ( .A(n10612), .ZN(n12322) );
  INV_X1 U7390 ( .A(n10046), .ZN(n10071) );
  NAND2_X1 U7391 ( .A1(n14169), .A2(n14170), .ZN(n14171) );
  INV_X1 U7392 ( .A(n9774), .ZN(n12335) );
  BUF_X1 U7393 ( .A(n7622), .Z(n8076) );
  AND3_X1 U7394 ( .A1(n7576), .A2(n7575), .A3(n7574), .ZN(n15057) );
  MUX2_X1 U7395 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8215), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n8217) );
  INV_X2 U7396 ( .A(n12130), .ZN(n9027) );
  AND2_X1 U7397 ( .A1(n6624), .A2(n6730), .ZN(n8865) );
  INV_X2 U7398 ( .A(n6772), .ZN(n9589) );
  INV_X1 U7400 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14138) );
  AND2_X1 U7401 ( .A1(n8350), .A2(n8329), .ZN(n8330) );
  XNOR2_X1 U7402 ( .A(n14171), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n14205) );
  BUF_X2 U7403 ( .A(n7610), .Z(n9106) );
  CLKBUF_X2 U7404 ( .A(n7987), .Z(n7735) );
  NAND2_X1 U7405 ( .A1(n8288), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8260) );
  BUF_X1 U7406 ( .A(n8244), .Z(n12201) );
  AOI21_X1 U7407 ( .B1(n13858), .B2(n13868), .A(n6896), .ZN(n13842) );
  AND2_X1 U7408 ( .A1(n8969), .A2(n8968), .ZN(n12635) );
  MUX2_X1 U7409 ( .A(n12824), .B(n12823), .S(n15132), .Z(n12825) );
  INV_X1 U7410 ( .A(n7562), .ZN(n12938) );
  XNOR2_X1 U7411 ( .A(n8237), .B(n8236), .ZN(n13488) );
  INV_X1 U7412 ( .A(n12201), .ZN(n11284) );
  INV_X1 U7413 ( .A(n14414), .ZN(n9532) );
  XNOR2_X1 U7414 ( .A(n14321), .B(n14320), .ZN(n14319) );
  INV_X1 U7415 ( .A(n7675), .ZN(n8046) );
  NAND2_X1 U7416 ( .A1(n7448), .A2(n7449), .ZN(n12696) );
  NAND2_X2 U7417 ( .A1(n10048), .A2(n10047), .ZN(n13808) );
  XNOR2_X2 U7418 ( .A(n8742), .B(n8740), .ZN(n13052) );
  NAND2_X2 U7419 ( .A1(n12974), .A2(n8722), .ZN(n8742) );
  OR2_X1 U7420 ( .A1(n8545), .A2(n8267), .ZN(n7543) );
  NAND4_X2 U7421 ( .A1(n8343), .A2(n8342), .A3(n8341), .A4(n8340), .ZN(n13109)
         );
  INV_X2 U7422 ( .A(n12130), .ZN(n8794) );
  OAI21_X2 U7423 ( .B1(n14245), .B2(n14244), .A(n14283), .ZN(n14442) );
  INV_X1 U7424 ( .A(n8545), .ZN(n8835) );
  NOR2_X2 U7425 ( .A1(n7972), .A2(n7971), .ZN(n7983) );
  AND3_X2 U7426 ( .A1(n7223), .A2(n7221), .A3(n7222), .ZN(n9575) );
  XNOR2_X2 U7427 ( .A(n6870), .B(P3_IR_REG_2__SCAN_IN), .ZN(n10773) );
  NOR2_X4 U7428 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9370) );
  AND2_X2 U7429 ( .A1(n10342), .A2(n10344), .ZN(n12313) );
  INV_X2 U7430 ( .A(n12313), .ZN(n10348) );
  NAND2_X2 U7431 ( .A1(n7128), .A2(n7127), .ZN(n13509) );
  INV_X1 U7433 ( .A(n10603), .ZN(n12284) );
  XNOR2_X2 U7434 ( .A(n13671), .B(n14585), .ZN(n10892) );
  OAI21_X2 U7435 ( .B1(n7439), .B2(n7440), .A(n7641), .ZN(n11824) );
  NOR2_X2 U7436 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n14211), .ZN(n14210) );
  OAI21_X1 U7437 ( .B1(n12984), .B2(n6940), .A(n6938), .ZN(n8863) );
  OAI21_X1 U7438 ( .B1(n9836), .B2(n6830), .A(n6828), .ZN(n12471) );
  NAND2_X1 U7439 ( .A1(n12299), .A2(n12298), .ZN(n13570) );
  NAND2_X1 U7440 ( .A1(n12732), .A2(n7916), .ZN(n12720) );
  NAND2_X1 U7441 ( .A1(n7881), .A2(n7880), .ZN(n12760) );
  AND2_X1 U7442 ( .A1(n14416), .A2(n9533), .ZN(n14370) );
  NAND2_X1 U7443 ( .A1(n9517), .A2(n6639), .ZN(n14416) );
  OAI21_X1 U7444 ( .B1(n11501), .B2(n9054), .A(n9055), .ZN(n11645) );
  OR2_X1 U7445 ( .A1(n14366), .A2(n11651), .ZN(n14371) );
  INV_X1 U7446 ( .A(n12052), .ZN(n9080) );
  NAND2_X1 U7447 ( .A1(n8459), .A2(n8458), .ZN(n12022) );
  NAND2_X1 U7448 ( .A1(n9145), .A2(n9141), .ZN(n15028) );
  OAI211_X1 U7449 ( .C1(n7987), .C2(SI_2_), .A(n7602), .B(n7601), .ZN(n15050)
         );
  NAND2_X1 U7450 ( .A1(n7962), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7626) );
  INV_X1 U7451 ( .A(n11987), .ZN(n7498) );
  NAND2_X1 U7452 ( .A1(n9889), .A2(n9888), .ZN(n10707) );
  BUF_X2 U7453 ( .A(n7622), .Z(n6620) );
  INV_X4 U7455 ( .A(n9904), .ZN(n9899) );
  INV_X2 U7456 ( .A(n14558), .ZN(n10703) );
  NAND2_X2 U7458 ( .A1(n7585), .A2(n7572), .ZN(n7987) );
  NAND2_X4 U7459 ( .A1(n7002), .A2(n7567), .ZN(n7675) );
  INV_X2 U7460 ( .A(n13359), .ZN(n8272) );
  CLKBUF_X3 U7461 ( .A(n11978), .Z(n6622) );
  NAND4_X1 U7463 ( .A1(n9384), .A2(n9383), .A3(n9382), .A4(n9381), .ZN(n14583)
         );
  INV_X4 U7464 ( .A(n9729), .ZN(n10050) );
  INV_X4 U7465 ( .A(n10053), .ZN(n9725) );
  INV_X2 U7466 ( .A(n9379), .ZN(n9729) );
  XNOR2_X1 U7467 ( .A(n9326), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9327) );
  NAND3_X1 U7468 ( .A1(n8381), .A2(n15356), .A3(n8183), .ZN(n8200) );
  NAND3_X1 U7469 ( .A1(n6790), .A2(n6887), .A3(n15343), .ZN(n6793) );
  AND2_X1 U7470 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n6790) );
  OAI211_X1 U7471 ( .C1(n12210), .C2(n12132), .A(n11284), .B(n6633), .ZN(
        n12200) );
  NOR2_X1 U7472 ( .A1(n12636), .A2(n7545), .ZN(n8958) );
  NAND2_X1 U7473 ( .A1(n8942), .A2(n8941), .ZN(n12648) );
  XNOR2_X1 U7474 ( .A(n8062), .B(n8061), .ZN(n8087) );
  NAND2_X1 U7475 ( .A1(n9846), .A2(n9845), .ZN(n12349) );
  AND2_X1 U7476 ( .A1(n7217), .A2(n7216), .ZN(n6969) );
  OR2_X1 U7477 ( .A1(n13230), .A2(n13229), .ZN(n13232) );
  NAND2_X1 U7478 ( .A1(n13050), .A2(n8743), .ZN(n8759) );
  NAND2_X1 U7479 ( .A1(n12678), .A2(n7968), .ZN(n12666) );
  NAND2_X1 U7480 ( .A1(n12679), .A2(n12680), .ZN(n12678) );
  OR2_X1 U7481 ( .A1(n8014), .A2(n8013), .ZN(n8016) );
  NAND2_X1 U7482 ( .A1(n13926), .A2(n13925), .ZN(n13924) );
  XNOR2_X1 U7483 ( .A(n12396), .B(n12671), .ZN(n12654) );
  NAND2_X1 U7484 ( .A1(n7989), .A2(n7988), .ZN(n9838) );
  NAND2_X1 U7485 ( .A1(n8772), .A2(n8771), .ZN(n13398) );
  INV_X1 U7486 ( .A(n12675), .ZN(n12831) );
  NAND2_X1 U7487 ( .A1(n8647), .A2(n7404), .ZN(n12964) );
  AND2_X1 U7488 ( .A1(n8101), .A2(n9218), .ZN(n7546) );
  NAND2_X1 U7489 ( .A1(n12760), .A2(n7459), .ZN(n12745) );
  NAND2_X1 U7490 ( .A1(n13009), .A2(n6685), .ZN(n8647) );
  NAND2_X1 U7491 ( .A1(n8100), .A2(n12748), .ZN(n12742) );
  INV_X1 U7492 ( .A(n12757), .ZN(n7881) );
  OAI21_X1 U7493 ( .B1(n7984), .B2(n7113), .A(n6758), .ZN(n7112) );
  NAND2_X1 U7494 ( .A1(n14362), .A2(n14367), .ZN(n14361) );
  NAND2_X1 U7495 ( .A1(n13518), .A2(n13519), .ZN(n13517) );
  NAND2_X1 U7496 ( .A1(n6871), .A2(n11856), .ZN(n12508) );
  NAND2_X1 U7497 ( .A1(n7935), .A2(n7934), .ZN(n7945) );
  NOR2_X1 U7498 ( .A1(n14309), .A2(n14310), .ZN(n7220) );
  AOI21_X1 U7499 ( .B1(n6859), .B2(n6857), .A(n6856), .ZN(n6855) );
  NAND2_X1 U7500 ( .A1(n7055), .A2(n14243), .ZN(n14285) );
  NAND2_X1 U7501 ( .A1(n11684), .A2(n9782), .ZN(n11762) );
  NAND2_X1 U7502 ( .A1(n8557), .A2(n8538), .ZN(n10807) );
  NAND2_X1 U7503 ( .A1(n9492), .A2(n9491), .ZN(n14290) );
  NAND2_X1 U7504 ( .A1(n7997), .A2(n7996), .ZN(n12656) );
  NAND2_X1 U7505 ( .A1(n9482), .A2(n9481), .ZN(n14383) );
  NAND2_X2 U7506 ( .A1(n8479), .A2(n8478), .ZN(n12031) );
  NAND2_X1 U7507 ( .A1(n9467), .A2(n9466), .ZN(n14636) );
  NAND2_X1 U7508 ( .A1(n8436), .A2(n8435), .ZN(n12019) );
  INV_X2 U7509 ( .A(n15074), .ZN(n15056) );
  AND3_X1 U7510 ( .A1(n7727), .A2(n7726), .A3(n7725), .ZN(n11888) );
  NAND2_X1 U7511 ( .A1(n9777), .A2(n11495), .ZN(n7537) );
  INV_X2 U7512 ( .A(n14829), .ZN(n6621) );
  NAND2_X1 U7513 ( .A1(n9417), .A2(n9416), .ZN(n11180) );
  AND3_X1 U7514 ( .A1(n7672), .A2(n7671), .A3(n7670), .ZN(n15006) );
  XNOR2_X1 U7515 ( .A(n10958), .B(n11040), .ZN(n14516) );
  OR2_X1 U7516 ( .A1(n15001), .A2(n15097), .ZN(n11705) );
  NAND4_X2 U7517 ( .A1(n7626), .A2(n7625), .A3(n7624), .A4(n7623), .ZN(n15026)
         );
  NAND2_X1 U7518 ( .A1(n8312), .A2(n8311), .ZN(n13031) );
  OAI211_X1 U7519 ( .C1(n7987), .C2(n10132), .A(n7587), .B(n7586), .ZN(n11947)
         );
  NAND4_X2 U7520 ( .A1(n7593), .A2(n7592), .A3(n7591), .A4(n7590), .ZN(n15060)
         );
  AND2_X1 U7521 ( .A1(n9411), .A2(n9410), .ZN(n10958) );
  NAND2_X1 U7522 ( .A1(n8351), .A2(n8350), .ZN(n8356) );
  INV_X1 U7523 ( .A(n7715), .ZN(n7622) );
  NAND2_X1 U7524 ( .A1(n8331), .A2(n8330), .ZN(n8351) );
  NAND4_X2 U7525 ( .A1(n8270), .A2(n8269), .A3(n8268), .A4(n7543), .ZN(n13114)
         );
  CLKBUF_X1 U7526 ( .A(n8834), .Z(n6776) );
  OAI21_X1 U7527 ( .B1(n7681), .B2(n7680), .A(n7682), .ZN(n7700) );
  CLKBUF_X2 U7528 ( .A(n7589), .Z(n6627) );
  INV_X1 U7529 ( .A(n10706), .ZN(n10709) );
  INV_X1 U7530 ( .A(n8657), .ZN(n8288) );
  AND2_X1 U7531 ( .A1(n12131), .A2(n11284), .ZN(n10502) );
  OR2_X1 U7532 ( .A1(n8545), .A2(n8257), .ZN(n8258) );
  NAND2_X2 U7533 ( .A1(n8433), .A2(n7572), .ZN(n12125) );
  INV_X1 U7534 ( .A(n8912), .ZN(n8904) );
  XNOR2_X1 U7535 ( .A(n7560), .B(P3_IR_REG_30__SCAN_IN), .ZN(n7565) );
  INV_X4 U7536 ( .A(n9607), .ZN(n9665) );
  XNOR2_X1 U7537 ( .A(n7571), .B(n7043), .ZN(n8075) );
  BUF_X4 U7538 ( .A(n9390), .Z(n6623) );
  AND2_X1 U7539 ( .A1(n9328), .A2(n14146), .ZN(n9568) );
  NAND2_X1 U7540 ( .A1(n9327), .A2(n9328), .ZN(n9607) );
  OR2_X1 U7541 ( .A1(n12927), .A2(n8127), .ZN(n7560) );
  NAND2_X1 U7542 ( .A1(n8244), .A2(n11208), .ZN(n12203) );
  CLKBUF_X1 U7543 ( .A(n8917), .Z(n13491) );
  AND2_X1 U7544 ( .A1(n8397), .A2(n8379), .ZN(n8380) );
  NAND2_X1 U7545 ( .A1(n9680), .A2(n9679), .ZN(n14158) );
  XNOR2_X1 U7546 ( .A(n9588), .B(n9702), .ZN(n13930) );
  XNOR2_X1 U7547 ( .A(n7346), .B(n9321), .ZN(n9722) );
  XNOR2_X1 U7548 ( .A(n9684), .B(n9683), .ZN(n14152) );
  XNOR2_X1 U7549 ( .A(n8194), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8244) );
  INV_X2 U7550 ( .A(n12933), .ZN(n11943) );
  OR2_X1 U7551 ( .A1(n8865), .A2(n13478), .ZN(n8193) );
  INV_X1 U7552 ( .A(n12163), .ZN(n11208) );
  XNOR2_X1 U7553 ( .A(n8195), .B(P2_IR_REG_20__SCAN_IN), .ZN(n12163) );
  AND2_X1 U7554 ( .A1(n9676), .A2(n7369), .ZN(n9325) );
  OR2_X1 U7555 ( .A1(n9678), .A2(n14138), .ZN(n6765) );
  NAND2_X1 U7556 ( .A1(n7052), .A2(n7050), .ZN(n14167) );
  AND2_X2 U7557 ( .A1(n9575), .A2(n7539), .ZN(n9676) );
  AND2_X1 U7558 ( .A1(n9586), .A2(n9673), .ZN(n9678) );
  NAND2_X2 U7559 ( .A1(n7572), .A2(P3_U3151), .ZN(n12944) );
  INV_X2 U7560 ( .A(n8213), .ZN(n6624) );
  AND3_X2 U7561 ( .A1(n7157), .A2(n7222), .A3(n7221), .ZN(n9586) );
  INV_X4 U7562 ( .A(n8226), .ZN(n7572) );
  NOR2_X1 U7563 ( .A1(n9311), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n7222) );
  AND2_X1 U7564 ( .A1(n9314), .A2(n9388), .ZN(n7223) );
  AND2_X1 U7565 ( .A1(n7373), .A2(n9683), .ZN(n7369) );
  NOR2_X1 U7566 ( .A1(n8200), .A2(n8202), .ZN(n8190) );
  AND3_X1 U7567 ( .A1(n8198), .A2(n8218), .A3(n7526), .ZN(n8309) );
  AND3_X1 U7568 ( .A1(n9314), .A2(n9388), .A3(n9574), .ZN(n7157) );
  NAND3_X1 U7569 ( .A1(n8406), .A2(n8430), .A3(n6902), .ZN(n8201) );
  AND2_X2 U7570 ( .A1(n9370), .A2(n9313), .ZN(n9388) );
  AND4_X1 U7571 ( .A1(n7889), .A2(n7831), .A3(n7888), .A4(n7554), .ZN(n7536)
         );
  NAND4_X1 U7572 ( .A1(n6890), .A2(n6889), .A3(n6888), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n6794) );
  AND2_X1 U7573 ( .A1(n7551), .A2(n15392), .ZN(n6760) );
  AND3_X1 U7574 ( .A1(n15219), .A2(n8187), .A3(n8186), .ZN(n8204) );
  INV_X1 U7575 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9503) );
  NOR3_X1 U7576 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .A3(
        P1_IR_REG_4__SCAN_IN), .ZN(n9314) );
  INV_X1 U7577 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7801) );
  INV_X1 U7578 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9574) );
  INV_X1 U7579 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7831) );
  INV_X1 U7580 ( .A(P1_RD_REG_SCAN_IN), .ZN(n6888) );
  INV_X4 U7581 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X4 U7582 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X4 U7583 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7584 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n7552) );
  NOR2_X1 U7585 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n7553) );
  INV_X1 U7586 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8181) );
  INV_X1 U7587 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8180) );
  INV_X1 U7588 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8179) );
  INV_X1 U7589 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8185) );
  INV_X1 U7590 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8184) );
  INV_X1 U7591 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6775) );
  INV_X1 U7592 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6902) );
  INV_X1 U7593 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n8183) );
  INV_X1 U7594 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8430) );
  INV_X1 U7595 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8406) );
  INV_X1 U7596 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7888) );
  INV_X1 U7597 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n15392) );
  INV_X1 U7598 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7853) );
  OAI21_X2 U7599 ( .B1(n11798), .B2(n8596), .A(n8595), .ZN(n12997) );
  NAND2_X2 U7600 ( .A1(n11576), .A2(n8555), .ZN(n11798) );
  NAND2_X1 U7601 ( .A1(n8396), .A2(n8395), .ZN(n10828) );
  NAND2_X1 U7602 ( .A1(n8129), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7571) );
  OR2_X2 U7603 ( .A1(n8129), .A2(n7042), .ZN(n6703) );
  NAND2_X2 U7604 ( .A1(n8152), .A2(n7462), .ZN(n8129) );
  NOR2_X4 U7605 ( .A1(n8063), .A2(P3_IR_REG_22__SCAN_IN), .ZN(n8152) );
  NAND2_X2 U7606 ( .A1(n8068), .A2(n8072), .ZN(n8063) );
  OAI21_X2 U7607 ( .B1(n14247), .B2(n14246), .A(n14441), .ZN(n14446) );
  OAI21_X2 U7608 ( .B1(n12696), .B2(n6715), .A(n6630), .ZN(n6761) );
  NAND2_X1 U7609 ( .A1(n7585), .A2(n7572), .ZN(n6625) );
  MUX2_X1 U7610 ( .A(n8943), .B(n12823), .S(n15119), .Z(n8946) );
  NAND2_X2 U7611 ( .A1(n6703), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7561) );
  OAI22_X2 U7612 ( .A1(n11786), .A2(n7133), .B1(n7134), .B2(n12224), .ZN(
        n13518) );
  OAI211_X1 U7613 ( .C1(n10124), .C2(n10046), .A(n9392), .B(n9391), .ZN(n13538) );
  OAI211_X2 U7614 ( .C1(n11824), .C2(n7689), .A(n11828), .B(n7688), .ZN(n7691)
         );
  NOR2_X4 U7615 ( .A1(n13997), .A2(n14116), .ZN(n14000) );
  NAND2_X1 U7616 ( .A1(n10176), .A2(n7572), .ZN(n9390) );
  NOR2_X4 U7617 ( .A1(n7633), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n7635) );
  NAND2_X2 U7618 ( .A1(n7158), .A2(n6827), .ZN(n7633) );
  NAND2_X1 U7619 ( .A1(n7179), .A2(n9790), .ZN(n7178) );
  INV_X1 U7620 ( .A(n12364), .ZN(n7179) );
  AOI21_X1 U7621 ( .B1(n7493), .B2(n7491), .A(n7490), .ZN(n7489) );
  INV_X1 U7622 ( .A(n12055), .ZN(n7490) );
  NOR2_X1 U7623 ( .A1(n7494), .A2(n9004), .ZN(n7491) );
  OR2_X1 U7624 ( .A1(n12417), .A2(n7169), .ZN(n7168) );
  INV_X1 U7625 ( .A(n9798), .ZN(n6860) );
  OR2_X1 U7626 ( .A1(n12901), .A2(n12721), .ZN(n9218) );
  INV_X1 U7627 ( .A(n6822), .ZN(n6819) );
  AND2_X1 U7628 ( .A1(n8218), .A2(n8188), .ZN(n8189) );
  NAND2_X1 U7629 ( .A1(n7278), .A2(n7277), .ZN(n7275) );
  AOI21_X1 U7630 ( .B1(n6983), .B2(n8575), .A(n6704), .ZN(n6982) );
  NAND2_X1 U7631 ( .A1(n8535), .A2(n8534), .ZN(n8576) );
  OR2_X1 U7632 ( .A1(n12751), .A2(n12758), .ZN(n9208) );
  AOI21_X1 U7633 ( .B1(n7088), .B2(n7090), .A(n6712), .ZN(n7086) );
  XNOR2_X1 U7634 ( .A(n13388), .B(n13089), .ZN(n13205) );
  NAND2_X1 U7635 ( .A1(n13298), .A2(n12187), .ZN(n9067) );
  NAND2_X1 U7636 ( .A1(n7262), .A2(n7258), .ZN(n7257) );
  NOR2_X1 U7637 ( .A1(n7260), .A2(n9956), .ZN(n7258) );
  INV_X1 U7638 ( .A(n9954), .ZN(n7260) );
  OAI22_X1 U7639 ( .A1(n12046), .A2(n7514), .B1(n12047), .B2(n7513), .ZN(
        n12060) );
  INV_X1 U7640 ( .A(n12045), .ZN(n7513) );
  NOR2_X1 U7641 ( .A1(n12045), .A2(n12048), .ZN(n7514) );
  INV_X1 U7642 ( .A(n7868), .ZN(n7110) );
  NAND2_X1 U7643 ( .A1(n7493), .A2(n12056), .ZN(n7492) );
  AND2_X1 U7644 ( .A1(n6674), .A2(n7322), .ZN(n7321) );
  INV_X1 U7645 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n6889) );
  NAND2_X1 U7646 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n7051), .ZN(n7050) );
  NAND2_X1 U7647 ( .A1(n14207), .A2(n14208), .ZN(n7052) );
  INV_X1 U7648 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7051) );
  INV_X1 U7649 ( .A(n7177), .ZN(n7176) );
  NOR2_X1 U7650 ( .A1(n7178), .A2(n6863), .ZN(n6862) );
  INV_X1 U7651 ( .A(n11761), .ZN(n6863) );
  INV_X1 U7652 ( .A(n7028), .ZN(n7027) );
  OAI21_X1 U7653 ( .B1(n8102), .B2(n7029), .A(n8103), .ZN(n7028) );
  OAI21_X1 U7654 ( .B1(n7034), .B2(n7033), .A(n14337), .ZN(n7032) );
  OR2_X1 U7655 ( .A1(n12455), .A2(n14339), .ZN(n9186) );
  INV_X2 U7656 ( .A(n9854), .ZN(n10752) );
  NAND2_X1 U7657 ( .A1(n9301), .A2(n11451), .ZN(n9854) );
  AND2_X1 U7658 ( .A1(n7463), .A2(n7559), .ZN(n7462) );
  INV_X1 U7659 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7458) );
  OAI21_X1 U7660 ( .B1(n7756), .B2(n7095), .A(n7091), .ZN(n7798) );
  AOI21_X1 U7661 ( .B1(n7093), .B2(n7094), .A(n7092), .ZN(n7091) );
  INV_X1 U7662 ( .A(n7796), .ZN(n7092) );
  INV_X1 U7663 ( .A(n7097), .ZN(n7093) );
  OR2_X1 U7664 ( .A1(n7798), .A2(n10683), .ZN(n7799) );
  NOR2_X1 U7665 ( .A1(n7775), .A2(n7098), .ZN(n7097) );
  AND2_X1 U7666 ( .A1(n10494), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7775) );
  INV_X1 U7667 ( .A(n7755), .ZN(n7098) );
  OR2_X1 U7668 ( .A1(n13370), .A2(n13152), .ZN(n12158) );
  NAND2_X1 U7669 ( .A1(n13484), .A2(n8239), .ZN(n8657) );
  NAND2_X1 U7670 ( .A1(n7480), .A2(n7478), .ZN(n9015) );
  NOR2_X1 U7671 ( .A1(n13171), .A2(n7479), .ZN(n7478) );
  INV_X1 U7672 ( .A(n7481), .ZN(n7479) );
  OAI21_X1 U7673 ( .B1(n9059), .B2(n7306), .A(n9061), .ZN(n7305) );
  AND2_X1 U7674 ( .A1(n6802), .A2(n9000), .ZN(n6801) );
  NAND2_X1 U7675 ( .A1(n8999), .A2(n6803), .ZN(n6802) );
  INV_X1 U7676 ( .A(n8998), .ZN(n6803) );
  NOR2_X1 U7677 ( .A1(n12035), .A2(n12044), .ZN(n7076) );
  INV_X1 U7678 ( .A(n10063), .ZN(n7277) );
  NOR2_X1 U7679 ( .A1(n13925), .A2(n7378), .ZN(n7377) );
  INV_X1 U7680 ( .A(n9614), .ZN(n7378) );
  NAND2_X1 U7681 ( .A1(n7321), .A2(n9747), .ZN(n6883) );
  INV_X1 U7682 ( .A(n8810), .ZN(n6997) );
  AND2_X1 U7683 ( .A1(n6945), .A2(n7409), .ZN(n6944) );
  AOI21_X1 U7684 ( .B1(n7411), .B2(n7413), .A(n6706), .ZN(n7409) );
  AOI21_X1 U7685 ( .B1(n7166), .B2(n7169), .A(n6696), .ZN(n7164) );
  NOR2_X1 U7686 ( .A1(n12379), .A2(n7171), .ZN(n7170) );
  INV_X1 U7687 ( .A(n9812), .ZN(n7171) );
  NAND2_X1 U7688 ( .A1(n12434), .A2(n12435), .ZN(n7172) );
  NAND2_X1 U7689 ( .A1(n9768), .A2(n7578), .ZN(n9771) );
  NAND2_X1 U7690 ( .A1(n6875), .A2(n6874), .ZN(n7201) );
  INV_X1 U7691 ( .A(n11518), .ZN(n6874) );
  AND2_X1 U7692 ( .A1(n12631), .A2(n12498), .ZN(n8051) );
  AND2_X1 U7693 ( .A1(n8961), .A2(n8035), .ZN(n9257) );
  AND2_X1 U7694 ( .A1(n9219), .A2(n9208), .ZN(n7039) );
  NOR2_X1 U7695 ( .A1(n12748), .A2(n7460), .ZN(n7459) );
  INV_X1 U7696 ( .A(n7882), .ZN(n7460) );
  NAND2_X1 U7697 ( .A1(n11053), .A2(n10980), .ZN(n15103) );
  INV_X1 U7698 ( .A(n15103), .ZN(n14345) );
  AND2_X1 U7699 ( .A1(n10751), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11046) );
  AOI22_X1 U7700 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n15324), .B1(n8039), 
        .B2(n8038), .ZN(n8052) );
  OAI21_X1 U7701 ( .B1(n7945), .B2(n7079), .A(n7077), .ZN(n7083) );
  INV_X1 U7702 ( .A(n7080), .ZN(n7079) );
  AOI21_X1 U7703 ( .B1(n7080), .B2(n7078), .A(n6650), .ZN(n7077) );
  INV_X1 U7704 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8072) );
  XNOR2_X1 U7705 ( .A(n7905), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12595) );
  OAI21_X1 U7706 ( .B1(n7851), .B2(n7183), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n7905) );
  NAND2_X1 U7707 ( .A1(n7184), .A2(n7889), .ZN(n7183) );
  INV_X1 U7708 ( .A(n7186), .ZN(n7184) );
  NAND2_X1 U7709 ( .A1(n7702), .A2(n7701), .ZN(n7721) );
  NAND2_X1 U7710 ( .A1(n7700), .A2(n7699), .ZN(n7702) );
  NOR4_X1 U7711 ( .A1(n12195), .A2(n13186), .A3(n13171), .A4(n12194), .ZN(
        n12198) );
  NOR2_X1 U7712 ( .A1(n8212), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n7507) );
  NOR2_X1 U7713 ( .A1(n6816), .A2(n6822), .ZN(n13210) );
  OAI21_X1 U7714 ( .B1(n13284), .B2(n9007), .A(n12162), .ZN(n9008) );
  NAND2_X1 U7715 ( .A1(n13313), .A2(n9066), .ZN(n13298) );
  NOR2_X1 U7716 ( .A1(n7495), .A2(n9003), .ZN(n7494) );
  INV_X1 U7717 ( .A(n9001), .ZN(n7495) );
  OR2_X1 U7718 ( .A1(n12035), .A2(n13102), .ZN(n7312) );
  NAND2_X1 U7719 ( .A1(n11003), .A2(n8989), .ZN(n10878) );
  OR2_X1 U7720 ( .A1(n13476), .A2(n13478), .ZN(n8234) );
  OAI21_X1 U7721 ( .B1(n8629), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8207) );
  INV_X1 U7722 ( .A(n10342), .ZN(n10343) );
  NAND2_X2 U7723 ( .A1(n9720), .A2(n9722), .ZN(n10176) );
  NOR2_X1 U7724 ( .A1(n13592), .A2(n7156), .ZN(n7155) );
  INV_X1 U7725 ( .A(n13581), .ZN(n7156) );
  AOI21_X1 U7726 ( .B1(n7272), .B2(n7274), .A(n6711), .ZN(n7270) );
  INV_X1 U7727 ( .A(n9568), .ZN(n9552) );
  INV_X1 U7728 ( .A(n9380), .ZN(n10053) );
  INV_X1 U7729 ( .A(n14028), .ZN(n10061) );
  NAND2_X1 U7730 ( .A1(n7368), .A2(n7366), .ZN(n13812) );
  AND2_X1 U7731 ( .A1(n13813), .A2(n7367), .ZN(n7366) );
  NAND2_X1 U7732 ( .A1(n13895), .A2(n7361), .ZN(n7360) );
  NOR2_X1 U7733 ( .A1(n13871), .A2(n7362), .ZN(n7361) );
  INV_X1 U7734 ( .A(n9641), .ZN(n7362) );
  XNOR2_X1 U7735 ( .A(n14106), .B(n13665), .ZN(n13954) );
  NOR2_X1 U7736 ( .A1(n13991), .A2(n7338), .ZN(n7337) );
  INV_X1 U7737 ( .A(n9754), .ZN(n7338) );
  NAND2_X1 U7738 ( .A1(n9551), .A2(n9550), .ZN(n12244) );
  OR2_X1 U7739 ( .A1(n14366), .A2(n14409), .ZN(n9962) );
  OR2_X1 U7740 ( .A1(n8627), .A2(n8672), .ZN(n8649) );
  NAND2_X1 U7741 ( .A1(n6977), .A2(n6976), .ZN(n8625) );
  AOI21_X1 U7742 ( .B1(n6979), .B2(n6981), .A(n6723), .ZN(n6976) );
  NAND2_X1 U7743 ( .A1(n8356), .A2(n8355), .ZN(n8376) );
  INV_X1 U7744 ( .A(n7160), .ZN(n7159) );
  OAI21_X1 U7745 ( .B1(n11493), .B2(n7161), .A(n11685), .ZN(n7160) );
  INV_X1 U7746 ( .A(n11053), .ZN(n9301) );
  NAND2_X1 U7747 ( .A1(n8814), .A2(n8813), .ZN(n13388) );
  NAND2_X1 U7748 ( .A1(n6970), .A2(n14376), .ZN(n14029) );
  NAND2_X1 U7749 ( .A1(n7518), .A2(n7517), .ZN(n11990) );
  OR2_X1 U7750 ( .A1(n11985), .A2(n7519), .ZN(n7517) );
  INV_X1 U7751 ( .A(n11984), .ZN(n7519) );
  NOR2_X1 U7752 ( .A1(n9918), .A2(n9921), .ZN(n7227) );
  NAND2_X1 U7753 ( .A1(n9918), .A2(n9921), .ZN(n7228) );
  NAND2_X1 U7754 ( .A1(n11996), .A2(n6923), .ZN(n6922) );
  AND2_X1 U7755 ( .A1(n11998), .A2(n6925), .ZN(n6924) );
  INV_X1 U7756 ( .A(n11996), .ZN(n6925) );
  NAND2_X1 U7757 ( .A1(n12012), .A2(n12014), .ZN(n7510) );
  NAND2_X1 U7758 ( .A1(n12016), .A2(n6920), .ZN(n6919) );
  INV_X1 U7759 ( .A(n7249), .ZN(n7245) );
  NOR2_X1 U7760 ( .A1(n7249), .A2(n7247), .ZN(n7246) );
  NAND2_X1 U7761 ( .A1(n12032), .A2(n12034), .ZN(n7512) );
  NOR2_X1 U7762 ( .A1(n9965), .A2(n7253), .ZN(n7251) );
  INV_X1 U7763 ( .A(n7257), .ZN(n7253) );
  AND2_X1 U7764 ( .A1(n7257), .A2(n7259), .ZN(n7256) );
  NAND2_X1 U7765 ( .A1(n7262), .A2(n6690), .ZN(n7259) );
  INV_X1 U7766 ( .A(n9965), .ZN(n7261) );
  OR2_X1 U7767 ( .A1(n12060), .A2(n6907), .ZN(n6906) );
  NAND2_X1 U7768 ( .A1(n12060), .A2(n6907), .ZN(n12062) );
  INV_X1 U7769 ( .A(n12058), .ZN(n6905) );
  INV_X1 U7770 ( .A(n7242), .ZN(n7238) );
  NOR2_X1 U7771 ( .A1(n7242), .A2(n7240), .ZN(n7239) );
  NAND2_X1 U7772 ( .A1(n12092), .A2(n7524), .ZN(n7523) );
  NOR2_X1 U7773 ( .A1(n6693), .A2(n6915), .ZN(n6914) );
  INV_X1 U7774 ( .A(n6801), .ZN(n6799) );
  INV_X1 U7775 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n15219) );
  OAI22_X1 U7776 ( .A1(n6929), .A2(n6692), .B1(n6931), .B2(n12116), .ZN(n12121) );
  NAND2_X1 U7777 ( .A1(n12114), .A2(n6930), .ZN(n6929) );
  NAND2_X1 U7778 ( .A1(n12116), .A2(n6931), .ZN(n6930) );
  NOR2_X1 U7779 ( .A1(n7492), .A2(n6799), .ZN(n6795) );
  INV_X1 U7780 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9306) );
  NOR2_X1 U7781 ( .A1(n7212), .A2(n13946), .ZN(n7211) );
  INV_X1 U7782 ( .A(n7213), .ZN(n7212) );
  INV_X1 U7783 ( .A(n9312), .ZN(n7221) );
  INV_X1 U7784 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14168) );
  INV_X1 U7785 ( .A(n9807), .ZN(n7169) );
  INV_X1 U7786 ( .A(n12425), .ZN(n9830) );
  XNOR2_X1 U7787 ( .A(n9774), .B(n15033), .ZN(n6826) );
  INV_X1 U7788 ( .A(n7022), .ZN(n7021) );
  INV_X1 U7789 ( .A(n7020), .ZN(n7019) );
  OAI21_X1 U7790 ( .B1(n6669), .B2(n7021), .A(n9265), .ZN(n7020) );
  AND2_X1 U7791 ( .A1(n9271), .A2(n7533), .ZN(n7024) );
  OR2_X1 U7792 ( .A1(n12618), .A2(n12614), .ZN(n7533) );
  NAND2_X1 U7793 ( .A1(n6968), .A2(n6966), .ZN(n6965) );
  INV_X1 U7794 ( .A(n10780), .ZN(n6968) );
  NAND2_X1 U7795 ( .A1(n6965), .A2(n6964), .ZN(n11427) );
  NAND2_X1 U7796 ( .A1(n7599), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n6964) );
  NAND4_X1 U7797 ( .A1(n11376), .A2(n14861), .A3(n14862), .A4(
        P3_REG2_REG_3__SCAN_IN), .ZN(n6872) );
  NAND2_X1 U7798 ( .A1(n14975), .A2(n6952), .ZN(n11527) );
  OR2_X1 U7799 ( .A1(n11441), .A2(n11440), .ZN(n6952) );
  AOI21_X1 U7800 ( .B1(n12558), .B2(n12557), .A(n6954), .ZN(n12576) );
  AND2_X1 U7801 ( .A1(n12556), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n6954) );
  INV_X1 U7802 ( .A(n9242), .ZN(n7038) );
  OR2_X1 U7803 ( .A1(n9838), .A2(n8107), .ZN(n9253) );
  NOR2_X1 U7804 ( .A1(n11893), .A2(n8094), .ZN(n7034) );
  NOR2_X1 U7805 ( .A1(n7712), .A2(n7456), .ZN(n7455) );
  INV_X1 U7806 ( .A(n7620), .ZN(n7441) );
  NAND2_X1 U7807 ( .A1(n9140), .A2(n9138), .ZN(n9129) );
  NAND2_X1 U7808 ( .A1(n8132), .A2(n6852), .ZN(n6851) );
  INV_X1 U7809 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n6852) );
  NAND2_X1 U7810 ( .A1(n7043), .A2(n7569), .ZN(n7042) );
  AND2_X1 U7811 ( .A1(n7464), .A2(n7558), .ZN(n7463) );
  AND2_X1 U7812 ( .A1(n7556), .A2(n7557), .ZN(n7464) );
  OAI21_X1 U7813 ( .B1(n7866), .B2(n7110), .A(n7883), .ZN(n7109) );
  NOR2_X1 U7814 ( .A1(n7110), .A2(n7106), .ZN(n7105) );
  INV_X1 U7815 ( .A(n7847), .ZN(n7106) );
  INV_X1 U7816 ( .A(n7799), .ZN(n7100) );
  AOI21_X1 U7817 ( .B1(n7817), .B2(n7103), .A(n6751), .ZN(n7101) );
  INV_X1 U7818 ( .A(n7778), .ZN(n7099) );
  AND2_X1 U7819 ( .A1(n8749), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8773) );
  INV_X1 U7820 ( .A(n7301), .ZN(n7300) );
  OAI21_X1 U7821 ( .B1(n6632), .B2(n7302), .A(n13270), .ZN(n7301) );
  INV_X1 U7822 ( .A(n9068), .ZN(n7302) );
  NAND2_X1 U7823 ( .A1(n6671), .A2(n9042), .ZN(n7316) );
  NAND2_X1 U7824 ( .A1(n8984), .A2(n7500), .ZN(n7499) );
  NOR2_X1 U7825 ( .A1(n8987), .A2(n7501), .ZN(n7500) );
  INV_X1 U7826 ( .A(n8983), .ZN(n7501) );
  OR2_X1 U7827 ( .A1(n7473), .A2(n7470), .ZN(n7469) );
  AND2_X1 U7828 ( .A1(n13254), .A2(n7474), .ZN(n7473) );
  INV_X1 U7829 ( .A(n7475), .ZN(n7470) );
  NAND2_X1 U7830 ( .A1(n9009), .A2(n7476), .ZN(n7474) );
  NOR2_X1 U7831 ( .A1(n13358), .A2(n13440), .ZN(n13362) );
  NAND2_X1 U7832 ( .A1(n11258), .A2(n7508), .ZN(n11296) );
  AND2_X1 U7833 ( .A1(n8996), .A2(n8994), .ZN(n7508) );
  NAND2_X1 U7834 ( .A1(n8433), .A2(n7309), .ZN(n7308) );
  NOR2_X1 U7835 ( .A1(n10129), .A2(n7311), .ZN(n7309) );
  AND2_X1 U7836 ( .A1(n8197), .A2(n7528), .ZN(n7526) );
  INV_X1 U7837 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7528) );
  OR2_X1 U7838 ( .A1(n11785), .A2(n7136), .ZN(n7135) );
  NAND2_X1 U7839 ( .A1(n7330), .A2(n7329), .ZN(n7328) );
  NOR2_X1 U7840 ( .A1(n7208), .A2(n13851), .ZN(n7206) );
  NOR2_X1 U7841 ( .A1(n13906), .A2(n7344), .ZN(n7343) );
  INV_X1 U7842 ( .A(n9758), .ZN(n7344) );
  NOR2_X1 U7843 ( .A1(n7358), .A2(n7355), .ZN(n7354) );
  INV_X1 U7844 ( .A(n9475), .ZN(n7357) );
  AND2_X1 U7845 ( .A1(n6884), .A2(n6883), .ZN(n6885) );
  AND2_X1 U7846 ( .A1(n11103), .A2(n6734), .ZN(n6884) );
  NAND2_X1 U7847 ( .A1(n10899), .A2(n7321), .ZN(n7319) );
  NAND2_X1 U7848 ( .A1(n6994), .A2(n8809), .ZN(n8829) );
  AND2_X1 U7849 ( .A1(n8787), .A2(n6997), .ZN(n6992) );
  OAI22_X1 U7850 ( .A1(n8764), .A2(n8763), .B1(SI_23_), .B2(n8762), .ZN(n8765)
         );
  NOR2_X1 U7851 ( .A1(n8682), .A2(SI_20_), .ZN(n6989) );
  INV_X1 U7852 ( .A(n8679), .ZN(n6987) );
  NAND2_X1 U7853 ( .A1(n8680), .A2(n8679), .ZN(n6990) );
  AND2_X1 U7854 ( .A1(n9702), .A2(n7282), .ZN(n7281) );
  INV_X1 U7855 ( .A(n6982), .ZN(n6981) );
  INV_X1 U7856 ( .A(n8299), .ZN(n6789) );
  OAI211_X1 U7857 ( .C1(n6794), .C2(n10128), .A(n6792), .B(n6791), .ZN(n8220)
         );
  NOR2_X1 U7858 ( .A1(n14455), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7062) );
  NAND2_X1 U7859 ( .A1(n12471), .A2(n9841), .ZN(n9846) );
  AND2_X1 U7860 ( .A1(n9837), .A2(n9835), .ZN(n12399) );
  NAND2_X1 U7861 ( .A1(n7173), .A2(n11275), .ZN(n6832) );
  AND2_X1 U7862 ( .A1(n11240), .A2(n6675), .ZN(n7173) );
  OR2_X1 U7863 ( .A1(n11239), .A2(n11240), .ZN(n7175) );
  NAND2_X1 U7864 ( .A1(n11762), .A2(n6862), .ZN(n6861) );
  XNOR2_X1 U7865 ( .A(n15050), .B(n9774), .ZN(n9773) );
  OR2_X1 U7866 ( .A1(n9806), .A2(n12778), .ZN(n9807) );
  NAND2_X1 U7867 ( .A1(n7567), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7436) );
  NAND2_X1 U7868 ( .A1(n12938), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7435) );
  NAND2_X1 U7869 ( .A1(n7002), .A2(n12938), .ZN(n7715) );
  OR2_X1 U7870 ( .A1(n10912), .A2(n6967), .ZN(n6966) );
  AND2_X1 U7871 ( .A1(n10777), .A2(n10778), .ZN(n6967) );
  NAND2_X1 U7872 ( .A1(n7188), .A2(n11426), .ZN(n14862) );
  XNOR2_X1 U7873 ( .A(n11434), .B(n11401), .ZN(n14931) );
  NAND2_X1 U7874 ( .A1(n14902), .A2(n6953), .ZN(n11434) );
  NAND2_X1 U7875 ( .A1(n11424), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n6953) );
  NAND2_X1 U7876 ( .A1(n14931), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n14930) );
  AND2_X1 U7877 ( .A1(n10754), .A2(n10753), .ZN(n10782) );
  NAND2_X1 U7878 ( .A1(n14966), .A2(n11439), .ZN(n14977) );
  AND2_X1 U7879 ( .A1(n7190), .A2(n7189), .ZN(n11514) );
  NAND2_X1 U7880 ( .A1(n14981), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7189) );
  XNOR2_X1 U7881 ( .A(n11527), .B(n11521), .ZN(n11442) );
  NAND2_X1 U7882 ( .A1(n11442), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n11529) );
  XNOR2_X1 U7883 ( .A(n12532), .B(n6955), .ZN(n12512) );
  NAND2_X1 U7884 ( .A1(n12512), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n12534) );
  NAND2_X1 U7885 ( .A1(n7192), .A2(n7191), .ZN(n12553) );
  INV_X1 U7886 ( .A(n12530), .ZN(n7191) );
  AND2_X1 U7887 ( .A1(n9253), .A2(n9252), .ZN(n9128) );
  INV_X1 U7888 ( .A(n12654), .ZN(n12651) );
  NAND2_X1 U7889 ( .A1(n12692), .A2(n6660), .ZN(n12664) );
  AOI21_X1 U7890 ( .B1(n7027), .B2(n7029), .A(n6691), .ZN(n7026) );
  AOI21_X1 U7891 ( .B1(n6668), .B2(n7452), .A(n7450), .ZN(n7449) );
  INV_X1 U7892 ( .A(n9224), .ZN(n7450) );
  NAND2_X1 U7893 ( .A1(n12720), .A2(n12719), .ZN(n12718) );
  NAND2_X1 U7894 ( .A1(n7546), .A2(n8102), .ZN(n12717) );
  AND2_X1 U7895 ( .A1(n9208), .A2(n9213), .ZN(n12748) );
  OR2_X1 U7896 ( .A1(n7865), .A2(n7447), .ZN(n7446) );
  AOI21_X1 U7897 ( .B1(n7445), .B2(n7444), .A(n6749), .ZN(n7443) );
  INV_X1 U7898 ( .A(n7003), .ZN(n12774) );
  AND2_X1 U7899 ( .A1(n9203), .A2(n9202), .ZN(n12776) );
  NOR2_X1 U7900 ( .A1(n7011), .A2(n7008), .ZN(n7007) );
  INV_X1 U7901 ( .A(n9194), .ZN(n7011) );
  INV_X1 U7902 ( .A(n9188), .ZN(n7008) );
  NAND2_X1 U7903 ( .A1(n7010), .A2(n9189), .ZN(n7009) );
  INV_X1 U7904 ( .A(n12810), .ZN(n7010) );
  INV_X1 U7905 ( .A(n12501), .ZN(n12802) );
  INV_X1 U7906 ( .A(n8096), .ZN(n14337) );
  AND3_X1 U7907 ( .A1(n7784), .A2(n7783), .A3(n7782), .ZN(n14339) );
  NAND2_X1 U7908 ( .A1(n7035), .A2(n7034), .ZN(n11896) );
  INV_X1 U7909 ( .A(n10980), .ZN(n11451) );
  INV_X1 U7910 ( .A(n15059), .ZN(n15043) );
  NAND2_X1 U7911 ( .A1(n8025), .A2(n8024), .ZN(n9842) );
  NAND2_X1 U7912 ( .A1(n7836), .A2(n7835), .ZN(n12484) );
  NAND2_X1 U7913 ( .A1(n6847), .A2(n8132), .ZN(n8134) );
  NAND2_X1 U7914 ( .A1(n8126), .A2(n11740), .ZN(n6847) );
  OR2_X1 U7915 ( .A1(n8126), .A2(n6851), .ZN(n6846) );
  NAND2_X1 U7916 ( .A1(n6850), .A2(n6849), .ZN(n6848) );
  INV_X1 U7917 ( .A(n6851), .ZN(n6849) );
  AOI21_X1 U7918 ( .B1(n7982), .B2(n6757), .A(n7112), .ZN(n8021) );
  OAI21_X1 U7919 ( .B1(n8063), .B2(n6865), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n6864) );
  NAND2_X1 U7920 ( .A1(n7556), .A2(n8064), .ZN(n6865) );
  XNOR2_X1 U7921 ( .A(n7983), .B(n13504), .ZN(n7982) );
  NAND2_X1 U7922 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n11282), .ZN(n7084) );
  CLKBUF_X1 U7923 ( .A(n8068), .Z(n8069) );
  NAND2_X1 U7924 ( .A1(n7933), .A2(n11202), .ZN(n7934) );
  OAI21_X1 U7925 ( .B1(P2_DATAO_REG_18__SCAN_IN), .B2(n11140), .A(n7904), .ZN(
        n7917) );
  INV_X1 U7926 ( .A(n7187), .ZN(n7185) );
  NAND2_X1 U7927 ( .A1(n7848), .A2(n7847), .ZN(n7867) );
  NAND2_X1 U7928 ( .A1(n7798), .A2(n10683), .ZN(n7817) );
  NAND2_X1 U7929 ( .A1(n6653), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7818) );
  NAND2_X1 U7930 ( .A1(n7756), .A2(n7097), .ZN(n7096) );
  INV_X1 U7931 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7754) );
  INV_X1 U7932 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7722) );
  AND2_X1 U7933 ( .A1(n10173), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7680) );
  NAND2_X1 U7934 ( .A1(n7198), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6870) );
  INV_X1 U7935 ( .A(n7158), .ZN(n7198) );
  XNOR2_X1 U7936 ( .A(n13452), .B(n8860), .ZN(n8550) );
  AND2_X1 U7937 ( .A1(n6950), .A2(n8530), .ZN(n6778) );
  INV_X1 U7938 ( .A(n11578), .ZN(n6950) );
  AND2_X1 U7939 ( .A1(n13377), .A2(n8914), .ZN(n8915) );
  INV_X1 U7940 ( .A(n10825), .ZN(n7406) );
  NOR2_X1 U7941 ( .A1(n7408), .A2(n10825), .ZN(n7407) );
  XNOR2_X1 U7942 ( .A(n12031), .B(n6776), .ZN(n8489) );
  INV_X1 U7943 ( .A(n13060), .ZN(n13075) );
  NAND2_X1 U7944 ( .A1(n12158), .A2(n12140), .ZN(n12197) );
  NAND2_X1 U7945 ( .A1(n12160), .A2(n12159), .ZN(n12210) );
  AND2_X1 U7946 ( .A1(n12215), .A2(n12201), .ZN(n10183) );
  AND2_X1 U7947 ( .A1(n8756), .A2(n8755), .ZN(n13019) );
  NAND2_X1 U7948 ( .A1(n13170), .A2(n13171), .ZN(n13169) );
  INV_X1 U7949 ( .A(n6814), .ZN(n6813) );
  OAI21_X1 U7950 ( .B1(n6818), .B2(n6821), .A(n7482), .ZN(n6814) );
  AOI21_X1 U7951 ( .B1(n7291), .B2(n7293), .A(n7482), .ZN(n7290) );
  INV_X1 U7952 ( .A(n7294), .ZN(n7291) );
  NAND2_X1 U7953 ( .A1(n13213), .A2(n13204), .ZN(n13199) );
  NAND2_X1 U7954 ( .A1(n13279), .A2(n13093), .ZN(n7476) );
  NOR2_X1 U7955 ( .A1(n13279), .A2(n13093), .ZN(n9009) );
  INV_X1 U7956 ( .A(n13268), .ZN(n13285) );
  AOI21_X1 U7957 ( .B1(n6661), .B2(n7494), .A(n7496), .ZN(n7493) );
  NOR2_X1 U7958 ( .A1(n13440), .A2(n9002), .ZN(n7496) );
  NAND2_X1 U7959 ( .A1(n7307), .A2(n9059), .ZN(n13347) );
  INV_X1 U7960 ( .A(n13345), .ZN(n7307) );
  NAND2_X1 U7961 ( .A1(n6800), .A2(n6801), .ZN(n11693) );
  OR2_X1 U7962 ( .A1(n11502), .A2(n6804), .ZN(n6800) );
  AND2_X1 U7963 ( .A1(n7074), .A2(n11298), .ZN(n11640) );
  NOR2_X1 U7964 ( .A1(n13452), .A2(n7075), .ZN(n7074) );
  INV_X1 U7965 ( .A(n7076), .ZN(n7075) );
  NAND2_X1 U7966 ( .A1(n9051), .A2(n9050), .ZN(n11293) );
  NAND2_X1 U7967 ( .A1(n6786), .A2(n12179), .ZN(n11258) );
  INV_X1 U7968 ( .A(n11260), .ZN(n6786) );
  NAND2_X1 U7969 ( .A1(n12011), .A2(n10829), .ZN(n7504) );
  NAND2_X1 U7970 ( .A1(n10878), .A2(n7505), .ZN(n7503) );
  NAND2_X1 U7971 ( .A1(n14765), .A2(n13107), .ZN(n7505) );
  NAND2_X1 U7972 ( .A1(n7503), .A2(n7502), .ZN(n10932) );
  AND2_X1 U7973 ( .A1(n12173), .A2(n7504), .ZN(n7502) );
  NAND2_X1 U7974 ( .A1(n7068), .A2(n7498), .ZN(n10988) );
  NAND2_X1 U7975 ( .A1(n8748), .A2(n8747), .ZN(n13404) );
  OR2_X1 U7976 ( .A1(n11574), .A2(n12125), .ZN(n8732) );
  NAND2_X1 U7977 ( .A1(n8687), .A2(n8686), .ZN(n13419) );
  NAND2_X1 U7978 ( .A1(n8611), .A2(n8610), .ZN(n13437) );
  NOR3_X1 U7979 ( .A1(n8212), .A2(P2_IR_REG_27__SCAN_IN), .A3(
        P2_IR_REG_28__SCAN_IN), .ZN(n7506) );
  NAND2_X1 U7980 ( .A1(n8216), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8214) );
  NAND2_X1 U7981 ( .A1(n6624), .A2(n7285), .ZN(n8870) );
  INV_X1 U7982 ( .A(n8212), .ZN(n7285) );
  AND2_X1 U7983 ( .A1(n8867), .A2(n8866), .ZN(n8877) );
  NAND2_X1 U7984 ( .A1(n8877), .A2(n8868), .ZN(n8880) );
  INV_X1 U7985 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8868) );
  INV_X1 U7986 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8901) );
  XNOR2_X1 U7987 ( .A(n8902), .B(n8901), .ZN(n11770) );
  OR2_X1 U7988 ( .A1(n8498), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8539) );
  OR2_X1 U7989 ( .A1(n8405), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8408) );
  INV_X1 U7990 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8198) );
  INV_X1 U7991 ( .A(n8286), .ZN(n7527) );
  NAND2_X1 U7992 ( .A1(n8218), .A2(n8197), .ZN(n8286) );
  AND2_X1 U7993 ( .A1(n13642), .A2(n7131), .ZN(n7130) );
  OR2_X1 U7994 ( .A1(n13571), .A2(n7132), .ZN(n7131) );
  INV_X1 U7995 ( .A(n12306), .ZN(n7132) );
  INV_X2 U7996 ( .A(n10348), .ZN(n12320) );
  AOI21_X1 U7997 ( .B1(n7141), .B2(n7140), .A(n7139), .ZN(n7138) );
  INV_X1 U7998 ( .A(n11603), .ZN(n7139) );
  INV_X1 U7999 ( .A(n7148), .ZN(n7140) );
  OR2_X1 U8000 ( .A1(n9454), .A2(n9453), .ZN(n9468) );
  AOI21_X1 U8001 ( .B1(n10603), .B2(n14013), .A(n10345), .ZN(n10346) );
  NAND2_X1 U8002 ( .A1(n12321), .A2(n10709), .ZN(n10347) );
  AND2_X1 U8003 ( .A1(n10365), .A2(n6762), .ZN(n10345) );
  AND2_X1 U8004 ( .A1(n13633), .A2(n7152), .ZN(n7151) );
  OR2_X1 U8005 ( .A1(n7154), .A2(n7155), .ZN(n7152) );
  AOI21_X1 U8006 ( .B1(n7273), .B2(n7276), .A(n6710), .ZN(n7272) );
  NOR2_X1 U8007 ( .A1(n7278), .A2(n7277), .ZN(n7276) );
  AOI21_X1 U8008 ( .B1(n7270), .B2(n7271), .A(n7266), .ZN(n7265) );
  INV_X1 U8009 ( .A(n7272), .ZN(n7271) );
  NAND2_X1 U8010 ( .A1(n7267), .A2(n10084), .ZN(n7266) );
  INV_X1 U8011 ( .A(n10083), .ZN(n10084) );
  OR2_X1 U8012 ( .A1(n13485), .A2(n10046), .ZN(n10048) );
  AOI21_X1 U8013 ( .B1(n7330), .B2(n7327), .A(n6700), .ZN(n7326) );
  NOR2_X1 U8014 ( .A1(n7332), .A2(n13813), .ZN(n7327) );
  AOI21_X1 U8015 ( .B1(n14093), .B2(n6665), .A(n7374), .ZN(n13893) );
  NAND2_X1 U8016 ( .A1(n7375), .A2(n6672), .ZN(n7374) );
  AND2_X1 U8017 ( .A1(n14162), .A2(n6772), .ZN(n13913) );
  INV_X1 U8018 ( .A(n10100), .ZN(n13925) );
  NAND2_X1 U8019 ( .A1(n14093), .A2(n7377), .ZN(n13921) );
  NAND2_X1 U8020 ( .A1(n13974), .A2(n6899), .ZN(n13953) );
  AND2_X1 U8021 ( .A1(n13954), .A2(n9756), .ZN(n6899) );
  AND3_X1 U8022 ( .A1(n9571), .A2(n9570), .A3(n9569), .ZN(n13584) );
  NAND2_X1 U8023 ( .A1(n14361), .A2(n6684), .ZN(n11907) );
  AND2_X1 U8024 ( .A1(n9962), .A2(n9963), .ZN(n14367) );
  NAND2_X1 U8025 ( .A1(n14308), .A2(n14307), .ZN(n9517) );
  NAND2_X1 U8026 ( .A1(n6877), .A2(n6880), .ZN(n14301) );
  INV_X1 U8027 ( .A(n6881), .ZN(n6880) );
  OAI21_X1 U8028 ( .B1(n11465), .B2(n6882), .A(n14302), .ZN(n6881) );
  INV_X1 U8029 ( .A(n14288), .ZN(n11792) );
  NAND2_X1 U8030 ( .A1(n14377), .A2(n9750), .ZN(n11466) );
  NAND2_X1 U8031 ( .A1(n11466), .A2(n11465), .ZN(n11464) );
  INV_X1 U8032 ( .A(n10092), .ZN(n11465) );
  AND2_X1 U8033 ( .A1(n11109), .A2(n9930), .ZN(n11156) );
  AND2_X1 U8034 ( .A1(n9930), .A2(n9929), .ZN(n11103) );
  AND2_X1 U8035 ( .A1(n9634), .A2(n9633), .ZN(n14071) );
  NAND2_X1 U8036 ( .A1(n9761), .A2(n9760), .ZN(n14376) );
  INV_X1 U8037 ( .A(n14634), .ZN(n14410) );
  INV_X1 U8038 ( .A(n14635), .ZN(n14626) );
  XNOR2_X1 U8039 ( .A(n10070), .B(n10069), .ZN(n13475) );
  NAND2_X1 U8040 ( .A1(n7419), .A2(n7416), .ZN(n10070) );
  NOR2_X1 U8041 ( .A1(n10043), .A2(n7422), .ZN(n7421) );
  INV_X1 U8042 ( .A(n10041), .ZN(n7422) );
  NAND2_X1 U8043 ( .A1(n8828), .A2(SI_26_), .ZN(n7430) );
  NAND2_X1 U8044 ( .A1(n6996), .A2(n8809), .ZN(n6995) );
  INV_X1 U8045 ( .A(n7431), .ZN(n6996) );
  AND2_X1 U8046 ( .A1(n9677), .A2(n9682), .ZN(n9706) );
  OR2_X1 U8047 ( .A1(n8765), .A2(n11661), .ZN(n8787) );
  NAND2_X1 U8048 ( .A1(n8766), .A2(n8767), .ZN(n7433) );
  INV_X1 U8049 ( .A(n8768), .ZN(n8767) );
  NAND2_X1 U8050 ( .A1(n6990), .A2(n10873), .ZN(n8681) );
  INV_X1 U8051 ( .A(n8683), .ZN(n8682) );
  NAND2_X1 U8052 ( .A1(n8701), .A2(n8681), .ZN(n8684) );
  OR2_X1 U8053 ( .A1(n6990), .A2(n10873), .ZN(n8701) );
  OR2_X1 U8054 ( .A1(n8576), .A2(n6981), .ZN(n6975) );
  AOI21_X1 U8055 ( .B1(n6982), .B2(n6984), .A(n6980), .ZN(n6979) );
  INV_X1 U8056 ( .A(n8598), .ZN(n6980) );
  NAND2_X1 U8057 ( .A1(n6978), .A2(n6982), .ZN(n8599) );
  NAND2_X1 U8058 ( .A1(n8576), .A2(n6983), .ZN(n6978) );
  NAND2_X1 U8059 ( .A1(n8475), .A2(n7414), .ZN(n7410) );
  NAND2_X1 U8060 ( .A1(n8283), .A2(n8282), .ZN(n8300) );
  NAND2_X1 U8061 ( .A1(n6937), .A2(n10160), .ZN(n8221) );
  INV_X1 U8062 ( .A(n8220), .ZN(n6937) );
  NAND2_X1 U8063 ( .A1(n8220), .A2(SI_1_), .ZN(n8225) );
  NAND2_X1 U8064 ( .A1(n14175), .A2(n14174), .ZN(n14228) );
  OR2_X1 U8065 ( .A1(n14222), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n14174) );
  AOI21_X1 U8066 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n14184), .A(n14183), .ZN(
        n14202) );
  AND2_X1 U8067 ( .A1(n14240), .A2(n14239), .ZN(n14183) );
  OAI22_X1 U8068 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14193), .B1(n14253), 
        .B2(n14192), .ZN(n14256) );
  NAND2_X1 U8069 ( .A1(n14317), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n7045) );
  OR2_X1 U8070 ( .A1(n14317), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n7046) );
  AOI21_X1 U8071 ( .B1(n6713), .B2(n6855), .A(n6637), .ZN(n6853) );
  NAND2_X1 U8072 ( .A1(n12335), .A2(n7163), .ZN(n7162) );
  AND2_X1 U8073 ( .A1(n7577), .A2(n12505), .ZN(n7163) );
  INV_X1 U8074 ( .A(n12733), .ZN(n12710) );
  AOI21_X1 U8075 ( .B1(n6842), .B2(n6844), .A(n6670), .ZN(n6839) );
  NAND2_X1 U8076 ( .A1(n7922), .A2(n7921), .ZN(n12848) );
  OR2_X1 U8077 ( .A1(n7735), .A2(n10873), .ZN(n7921) );
  NAND2_X1 U8078 ( .A1(n7949), .A2(n7948), .ZN(n12447) );
  OR2_X1 U8079 ( .A1(n7735), .A2(n7947), .ZN(n7948) );
  INV_X1 U8080 ( .A(n12500), .ZN(n12778) );
  NAND2_X1 U8081 ( .A1(n7893), .A2(n7892), .ZN(n12751) );
  INV_X1 U8082 ( .A(n12490), .ZN(n12462) );
  AND2_X1 U8083 ( .A1(n8034), .A2(n8033), .ZN(n12477) );
  AND2_X1 U8084 ( .A1(n9848), .A2(n10749), .ZN(n12473) );
  AND2_X1 U8085 ( .A1(n9853), .A2(n12766), .ZN(n12485) );
  OR2_X1 U8086 ( .A1(n14974), .A2(n14973), .ZN(n7190) );
  OR2_X1 U8087 ( .A1(n11839), .A2(n11840), .ZN(n6871) );
  INV_X1 U8088 ( .A(n12508), .ZN(n12507) );
  OR2_X1 U8089 ( .A1(n12509), .A2(n12510), .ZN(n6866) );
  XNOR2_X1 U8090 ( .A(n12527), .B(n12533), .ZN(n12509) );
  OAI211_X1 U8091 ( .C1(n7196), .C2(n7195), .A(n7194), .B(n12593), .ZN(n12594)
         );
  INV_X1 U8092 ( .A(n12586), .ZN(n7195) );
  AND2_X1 U8093 ( .A1(n6957), .A2(n6956), .ZN(n6781) );
  INV_X1 U8094 ( .A(n12608), .ZN(n6956) );
  NAND2_X1 U8095 ( .A1(n6958), .A2(n14992), .ZN(n6957) );
  XNOR2_X1 U8096 ( .A(n6782), .B(n12599), .ZN(n12609) );
  NAND2_X1 U8097 ( .A1(n6784), .A2(n6783), .ZN(n6782) );
  AOI21_X1 U8098 ( .B1(n12934), .B2(n9106), .A(n9105), .ZN(n14343) );
  NAND2_X1 U8099 ( .A1(n7018), .A2(n7022), .ZN(n9097) );
  NOR2_X1 U8100 ( .A1(n8085), .A2(n8084), .ZN(n8086) );
  NOR2_X1 U8101 ( .A1(n9868), .A2(n15045), .ZN(n8085) );
  NAND2_X1 U8102 ( .A1(n7873), .A2(n7872), .ZN(n12860) );
  INV_X1 U8103 ( .A(n9842), .ZN(n12639) );
  OAI211_X1 U8104 ( .C1(n7735), .C2(SI_11_), .A(n7762), .B(n7761), .ZN(n12925)
         );
  NOR2_X1 U8105 ( .A1(n8129), .A2(P3_IR_REG_27__SCAN_IN), .ZN(n7568) );
  XNOR2_X1 U8106 ( .A(n8065), .B(n8064), .ZN(n11053) );
  INV_X1 U8107 ( .A(SI_16_), .ZN(n10456) );
  NAND2_X1 U8108 ( .A1(n8652), .A2(n8651), .ZN(n13425) );
  INV_X1 U8109 ( .A(n6939), .ZN(n6938) );
  OAI21_X1 U8110 ( .B1(n6941), .B2(n6940), .A(n8848), .ZN(n6939) );
  INV_X1 U8111 ( .A(n7405), .ZN(n6940) );
  NAND2_X1 U8112 ( .A1(n8519), .A2(n8518), .ZN(n12044) );
  NAND2_X1 U8113 ( .A1(n6769), .A2(n6768), .ZN(n8247) );
  INV_X1 U8114 ( .A(n8245), .ZN(n6768) );
  INV_X1 U8115 ( .A(n13079), .ZN(n13065) );
  OR2_X1 U8116 ( .A1(n11141), .A2(n12125), .ZN(n8632) );
  AOI21_X1 U8117 ( .B1(n10628), .B2(n7391), .A(n7390), .ZN(n7389) );
  INV_X1 U8118 ( .A(n8349), .ZN(n7390) );
  INV_X1 U8119 ( .A(n8324), .ZN(n7391) );
  INV_X1 U8120 ( .A(n10628), .ZN(n7392) );
  NAND2_X1 U8121 ( .A1(n6812), .A2(n12137), .ZN(n6811) );
  INV_X1 U8122 ( .A(n10172), .ZN(n6812) );
  INV_X1 U8123 ( .A(n13019), .ZN(n13092) );
  NAND2_X1 U8124 ( .A1(n8288), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8269) );
  OAI21_X1 U8125 ( .B1(n13485), .B2(n12125), .A(n12124), .ZN(n13161) );
  AOI21_X1 U8126 ( .B1(n9036), .B2(n13350), .A(n9035), .ZN(n11967) );
  NAND2_X1 U8127 ( .A1(n9034), .A2(n9033), .ZN(n9035) );
  NAND2_X1 U8128 ( .A1(n13218), .A2(n7294), .ZN(n7289) );
  NAND2_X1 U8129 ( .A1(n7286), .A2(n7290), .ZN(n13381) );
  OR2_X1 U8130 ( .A1(n13218), .A2(n7292), .ZN(n7286) );
  OAI21_X1 U8131 ( .B1(n7465), .B2(n6820), .A(n6817), .ZN(n7483) );
  AND2_X1 U8132 ( .A1(n7295), .A2(n7296), .ZN(n13206) );
  OAI21_X1 U8133 ( .B1(n13210), .B2(n13219), .A(n7486), .ZN(n13195) );
  NAND2_X1 U8134 ( .A1(n14781), .A2(n9091), .ZN(n13354) );
  NOR2_X1 U8135 ( .A1(n14761), .A2(n8912), .ZN(n13338) );
  INV_X2 U8136 ( .A(n14770), .ZN(n13357) );
  INV_X1 U8137 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11140) );
  NAND2_X1 U8138 ( .A1(n14149), .A2(n10071), .ZN(n6974) );
  INV_X1 U8139 ( .A(n14071), .ZN(n13899) );
  OAI211_X2 U8140 ( .C1(n10046), .C2(n10129), .A(n7203), .B(n7202), .ZN(n14558) );
  NAND2_X1 U8141 ( .A1(n9564), .A2(n9563), .ZN(n14116) );
  NAND2_X1 U8142 ( .A1(n9643), .A2(n9642), .ZN(n14066) );
  OR2_X1 U8143 ( .A1(n14159), .A2(n10046), .ZN(n9643) );
  NOR2_X1 U8144 ( .A1(n7535), .A2(n7547), .ZN(n9409) );
  AND2_X1 U8145 ( .A1(n9452), .A2(n9451), .ZN(n14627) );
  AND2_X1 U8146 ( .A1(n10357), .A2(n10523), .ZN(n14634) );
  OR2_X1 U8147 ( .A1(n9558), .A2(n9557), .ZN(n13666) );
  NAND2_X1 U8148 ( .A1(n9654), .A2(n9653), .ZN(n13821) );
  AOI21_X1 U8149 ( .B1(n14052), .B2(n6640), .A(n6718), .ZN(n7365) );
  XNOR2_X1 U8150 ( .A(n6897), .B(n7329), .ZN(n14037) );
  AND2_X1 U8151 ( .A1(n7330), .A2(n6893), .ZN(n6892) );
  NAND2_X1 U8152 ( .A1(n9592), .A2(n9591), .ZN(n14106) );
  NAND2_X1 U8153 ( .A1(n9718), .A2(n10515), .ZN(n13962) );
  OAI211_X1 U8154 ( .C1(n14563), .C2(n14030), .A(n14029), .B(n6969), .ZN(
        n14124) );
  AOI21_X1 U8155 ( .B1(n14028), .B2(n14635), .A(n14027), .ZN(n7216) );
  OR2_X1 U8156 ( .A1(n14026), .A2(n10341), .ZN(n7217) );
  XNOR2_X1 U8157 ( .A(n9704), .B(P1_IR_REG_23__SCAN_IN), .ZN(n10366) );
  INV_X1 U8158 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11202) );
  INV_X1 U8159 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11142) );
  XNOR2_X1 U8160 ( .A(n14212), .B(n6771), .ZN(n15525) );
  NAND2_X1 U8161 ( .A1(n14282), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7055) );
  INV_X1 U8162 ( .A(n14451), .ZN(n7064) );
  AND2_X1 U8163 ( .A1(n9891), .A2(n9890), .ZN(n9892) );
  OAI21_X1 U8164 ( .B1(n9919), .B2(n7227), .A(n7228), .ZN(n9924) );
  NAND2_X1 U8165 ( .A1(n7225), .A2(n7224), .ZN(n9923) );
  NOR2_X1 U8166 ( .A1(n7227), .A2(n7226), .ZN(n7225) );
  NAND2_X1 U8167 ( .A1(n6926), .A2(n7520), .ZN(n12005) );
  OR2_X1 U8168 ( .A1(n7521), .A2(n12001), .ZN(n7520) );
  INV_X1 U8169 ( .A(n12000), .ZN(n7521) );
  NOR2_X1 U8170 ( .A1(n9936), .A2(n9937), .ZN(n7249) );
  NAND2_X1 U8171 ( .A1(n9935), .A2(n7250), .ZN(n7248) );
  AOI21_X1 U8172 ( .B1(n9936), .B2(n9937), .A(n6709), .ZN(n7250) );
  NAND2_X1 U8173 ( .A1(n6918), .A2(n6917), .ZN(n12025) );
  AOI21_X1 U8174 ( .B1(n6636), .B2(n6921), .A(n6705), .ZN(n6917) );
  NOR2_X1 U8175 ( .A1(n6920), .A2(n12016), .ZN(n6921) );
  NAND2_X1 U8176 ( .A1(n9943), .A2(n9945), .ZN(n7237) );
  AOI21_X1 U8177 ( .B1(n7261), .B2(n7256), .A(n7255), .ZN(n7254) );
  INV_X1 U8178 ( .A(n9964), .ZN(n7255) );
  NAND2_X1 U8179 ( .A1(n6903), .A2(n6904), .ZN(n12078) );
  INV_X1 U8180 ( .A(n12073), .ZN(n6904) );
  NOR2_X1 U8181 ( .A1(n9991), .A2(n9992), .ZN(n7242) );
  NOR2_X1 U8182 ( .A1(n6683), .A2(n7244), .ZN(n7243) );
  INV_X1 U8183 ( .A(n9989), .ZN(n7244) );
  NOR2_X1 U8184 ( .A1(n6916), .A2(n12091), .ZN(n6915) );
  NAND2_X1 U8185 ( .A1(n12091), .A2(n6916), .ZN(n6913) );
  NAND2_X1 U8186 ( .A1(n9998), .A2(n10000), .ZN(n7233) );
  NAND2_X1 U8187 ( .A1(n10009), .A2(n10011), .ZN(n7235) );
  NAND2_X1 U8188 ( .A1(n12103), .A2(n6911), .ZN(n6910) );
  NAND2_X1 U8189 ( .A1(n7231), .A2(n10020), .ZN(n7230) );
  INV_X1 U8190 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7551) );
  NAND2_X1 U8191 ( .A1(n9881), .A2(n9880), .ZN(n9883) );
  OR2_X1 U8192 ( .A1(n9879), .A2(n13930), .ZN(n9881) );
  INV_X1 U8193 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7554) );
  MUX2_X1 U8194 ( .A(n12136), .B(n12135), .S(n12155), .Z(n12146) );
  NAND2_X1 U8195 ( .A1(n13205), .A2(n12192), .ZN(n7477) );
  INV_X1 U8196 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8187) );
  INV_X1 U8197 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8186) );
  NAND2_X1 U8198 ( .A1(n8496), .A2(n8203), .ZN(n8559) );
  INV_X1 U8199 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8199) );
  NAND2_X1 U8200 ( .A1(n9883), .A2(n9882), .ZN(n10058) );
  NOR2_X1 U8201 ( .A1(n14106), .A2(n14110), .ZN(n7213) );
  NAND2_X1 U8202 ( .A1(n7431), .A2(n7430), .ZN(n7426) );
  NOR2_X1 U8203 ( .A1(n8909), .A2(n7429), .ZN(n7428) );
  INV_X1 U8204 ( .A(n7430), .ZN(n7429) );
  INV_X1 U8205 ( .A(n8570), .ZN(n8572) );
  INV_X1 U8206 ( .A(n7412), .ZN(n7411) );
  OAI21_X1 U8207 ( .B1(n7414), .B2(n7413), .A(n8514), .ZN(n7412) );
  INV_X1 U8208 ( .A(n8493), .ZN(n7413) );
  AND2_X1 U8209 ( .A1(n7411), .A2(n6947), .ZN(n6946) );
  NAND2_X1 U8210 ( .A1(n8453), .A2(n6948), .ZN(n6947) );
  INV_X1 U8211 ( .A(n8448), .ZN(n6948) );
  NAND2_X1 U8212 ( .A1(n6946), .A2(n6949), .ZN(n6945) );
  INV_X1 U8213 ( .A(n8453), .ZN(n6949) );
  INV_X1 U8214 ( .A(P2_RD_REG_SCAN_IN), .ZN(n6887) );
  NOR2_X1 U8215 ( .A1(n11884), .A2(n7181), .ZN(n7180) );
  INV_X1 U8216 ( .A(n9785), .ZN(n7181) );
  NAND2_X1 U8217 ( .A1(n11374), .A2(n11373), .ZN(n7188) );
  NAND2_X1 U8218 ( .A1(n14936), .A2(n6951), .ZN(n11438) );
  NAND2_X1 U8219 ( .A1(n14942), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n6951) );
  NAND2_X1 U8220 ( .A1(n12666), .A2(n8015), .ZN(n7457) );
  OR2_X1 U8221 ( .A1(n7950), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n7960) );
  INV_X1 U8222 ( .A(n9222), .ZN(n7029) );
  OR2_X1 U8223 ( .A1(n12719), .A2(n7452), .ZN(n7451) );
  INV_X1 U8224 ( .A(n7931), .ZN(n7452) );
  OR2_X1 U8225 ( .A1(n12447), .A2(n12711), .ZN(n9229) );
  NAND2_X1 U8226 ( .A1(n7874), .A2(n12418), .ZN(n7894) );
  INV_X1 U8227 ( .A(n7844), .ZN(n7447) );
  NOR2_X1 U8228 ( .A1(n12790), .A2(n7447), .ZN(n7444) );
  INV_X1 U8229 ( .A(n7865), .ZN(n7445) );
  NOR2_X1 U8230 ( .A1(n7007), .A2(n7005), .ZN(n7004) );
  INV_X1 U8231 ( .A(n8099), .ZN(n7005) );
  INV_X1 U8232 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n7692) );
  OR2_X1 U8233 ( .A1(n12503), .A2(n15006), .ZN(n9163) );
  AOI21_X1 U8234 ( .B1(n7117), .B2(n7120), .A(n7119), .ZN(n7116) );
  INV_X1 U8235 ( .A(n9113), .ZN(n7119) );
  INV_X1 U8236 ( .A(n7985), .ZN(n7113) );
  AND2_X1 U8237 ( .A1(n11772), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7971) );
  NOR2_X1 U8238 ( .A1(n7957), .A2(n7081), .ZN(n7080) );
  INV_X1 U8239 ( .A(n7084), .ZN(n7081) );
  OAI21_X1 U8240 ( .B1(P2_DATAO_REG_19__SCAN_IN), .B2(n11226), .A(n7919), .ZN(
        n7932) );
  AND2_X1 U8241 ( .A1(n7853), .A2(n7850), .ZN(n7187) );
  NAND2_X1 U8242 ( .A1(n6629), .A2(n7635), .ZN(n7800) );
  INV_X1 U8243 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7738) );
  INV_X1 U8244 ( .A(n7089), .ZN(n7088) );
  OAI21_X1 U8245 ( .B1(n7720), .B2(n7090), .A(n7736), .ZN(n7089) );
  INV_X1 U8246 ( .A(n7723), .ZN(n7090) );
  INV_X1 U8247 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7549) );
  NAND2_X1 U8248 ( .A1(n9077), .A2(n12203), .ZN(n8834) );
  NOR2_X1 U8249 ( .A1(n8634), .A2(n8633), .ZN(n8653) );
  NOR2_X1 U8250 ( .A1(n7477), .A2(n6825), .ZN(n6821) );
  NAND2_X1 U8251 ( .A1(n6824), .A2(n6823), .ZN(n6822) );
  NAND2_X1 U8252 ( .A1(n13398), .A2(n12987), .ZN(n6823) );
  INV_X1 U8253 ( .A(n13230), .ZN(n6825) );
  NOR2_X1 U8254 ( .A1(n13289), .A2(n13415), .ZN(n7073) );
  INV_X1 U8255 ( .A(n13303), .ZN(n6808) );
  NOR2_X1 U8256 ( .A1(n8481), .A2(n8480), .ZN(n8502) );
  INV_X1 U8257 ( .A(n7073), .ZN(n13274) );
  NAND2_X1 U8258 ( .A1(n6797), .A2(n6796), .ZN(n13315) );
  INV_X1 U8259 ( .A(n6798), .ZN(n6797) );
  OAI21_X1 U8260 ( .B1(n7492), .B2(n6716), .A(n7489), .ZN(n6798) );
  NAND2_X1 U8261 ( .A1(n10881), .A2(n14765), .ZN(n10934) );
  INV_X1 U8262 ( .A(n11213), .ZN(n7149) );
  INV_X1 U8263 ( .A(n11332), .ZN(n7143) );
  NOR2_X1 U8264 ( .A1(n9604), .A2(n13615), .ZN(n9605) );
  INV_X1 U8265 ( .A(n10062), .ZN(n7278) );
  OAI21_X1 U8266 ( .B1(n10082), .B2(n10081), .A(n10174), .ZN(n10083) );
  NAND2_X1 U8267 ( .A1(n7272), .A2(n7268), .ZN(n7267) );
  NOR2_X1 U8268 ( .A1(n10081), .A2(n7273), .ZN(n7268) );
  NOR2_X1 U8269 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n9308) );
  INV_X1 U8270 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9307) );
  INV_X1 U8271 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9310) );
  NAND2_X1 U8272 ( .A1(n14042), .A2(n13845), .ZN(n7334) );
  NOR2_X1 U8273 ( .A1(n7336), .A2(n7333), .ZN(n7332) );
  INV_X1 U8274 ( .A(n7334), .ZN(n7333) );
  INV_X1 U8275 ( .A(n9636), .ZN(n9627) );
  NOR2_X1 U8276 ( .A1(n7342), .A2(n13892), .ZN(n7341) );
  INV_X1 U8277 ( .A(n7343), .ZN(n7342) );
  NAND2_X1 U8278 ( .A1(n13906), .A2(n7376), .ZN(n7375) );
  INV_X1 U8279 ( .A(n9624), .ZN(n7376) );
  NAND2_X1 U8280 ( .A1(n9554), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9566) );
  OR2_X1 U8281 ( .A1(n9566), .A2(n9565), .ZN(n9580) );
  NAND2_X1 U8282 ( .A1(n9532), .A2(n9531), .ZN(n9959) );
  NAND2_X1 U8283 ( .A1(n7220), .A2(n9532), .ZN(n11651) );
  INV_X1 U8284 ( .A(n9751), .ZN(n6882) );
  NOR2_X1 U8285 ( .A1(n6882), .A2(n6879), .ZN(n6878) );
  INV_X1 U8286 ( .A(n9750), .ZN(n6879) );
  NAND2_X1 U8287 ( .A1(n9879), .A2(n13930), .ZN(n9880) );
  NAND2_X1 U8288 ( .A1(n10703), .A2(n10605), .ZN(n9889) );
  NAND2_X1 U8289 ( .A1(n14000), .A2(n6641), .ZN(n13927) );
  NAND2_X1 U8290 ( .A1(n14000), .A2(n7211), .ZN(n13942) );
  NAND2_X1 U8291 ( .A1(n14510), .A2(n14609), .ZN(n14509) );
  AND3_X1 U8292 ( .A1(n9317), .A2(n9316), .A3(n9315), .ZN(n9673) );
  OR2_X1 U8293 ( .A1(n10039), .A2(n7420), .ZN(n7419) );
  INV_X1 U8294 ( .A(n7421), .ZN(n7420) );
  AOI21_X1 U8295 ( .B1(n7421), .B2(n7418), .A(n7417), .ZN(n7416) );
  INV_X1 U8296 ( .A(n10065), .ZN(n7417) );
  INV_X1 U8297 ( .A(n10038), .ZN(n7418) );
  NAND2_X1 U8298 ( .A1(n7427), .A2(n7424), .ZN(n9017) );
  INV_X1 U8299 ( .A(n7425), .ZN(n7424) );
  NAND2_X1 U8300 ( .A1(n8829), .A2(n7428), .ZN(n7427) );
  OAI22_X1 U8301 ( .A1(n8909), .A2(n7426), .B1(n8908), .B2(SI_27_), .ZN(n7425)
         );
  NOR2_X1 U8302 ( .A1(n8828), .A2(SI_26_), .ZN(n7431) );
  NAND2_X1 U8303 ( .A1(n8725), .A2(n7947), .ZN(n8727) );
  NAND2_X1 U8304 ( .A1(n8726), .A2(SI_22_), .ZN(n8744) );
  NAND2_X1 U8305 ( .A1(n8625), .A2(n8624), .ZN(n8671) );
  INV_X1 U8306 ( .A(n8605), .ZN(n8604) );
  OR2_X1 U8307 ( .A1(n8576), .A2(n10328), .ZN(n8556) );
  INV_X1 U8308 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9518) );
  NOR2_X1 U8309 ( .A1(n8494), .A2(n7415), .ZN(n7414) );
  INV_X1 U8310 ( .A(n8474), .ZN(n7415) );
  NOR2_X1 U8311 ( .A1(n9450), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n9477) );
  OAI21_X1 U8312 ( .B1(n10067), .B2(n10173), .A(n6773), .ZN(n8352) );
  NAND2_X1 U8313 ( .A1(n10067), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n6773) );
  OAI21_X1 U8314 ( .B1(n8226), .B2(n10122), .A(n6886), .ZN(n8227) );
  XNOR2_X1 U8315 ( .A(n14167), .B(n7049), .ZN(n14216) );
  OAI21_X1 U8316 ( .B1(n14205), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n14172), .ZN(
        n14173) );
  XNOR2_X1 U8317 ( .A(P3_ADDR_REG_5__SCAN_IN), .B(n14173), .ZN(n14222) );
  AOI22_X1 U8318 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14177), .B1(n14228), .B2(
        n14176), .ZN(n14179) );
  AOI21_X1 U8319 ( .B1(n14953), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n14182), .ZN(
        n14240) );
  AND2_X1 U8320 ( .A1(n14203), .A2(n14204), .ZN(n14182) );
  AOI21_X1 U8321 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n14191), .A(n14190), .ZN(
        n14253) );
  NOR2_X1 U8322 ( .A1(n14249), .A2(n14248), .ZN(n14190) );
  OR2_X1 U8323 ( .A1(n7894), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7909) );
  AND2_X1 U8324 ( .A1(n12398), .A2(n9828), .ZN(n12425) );
  NAND2_X1 U8325 ( .A1(n11760), .A2(n7180), .ZN(n11881) );
  AOI21_X1 U8326 ( .B1(n7164), .B2(n7167), .A(n6843), .ZN(n6842) );
  INV_X1 U8327 ( .A(n12370), .ZN(n6843) );
  INV_X1 U8328 ( .A(n7164), .ZN(n6844) );
  INV_X1 U8329 ( .A(n6859), .ZN(n6858) );
  INV_X1 U8330 ( .A(n9797), .ZN(n6856) );
  INV_X1 U8331 ( .A(n6862), .ZN(n6857) );
  NAND2_X1 U8332 ( .A1(n7537), .A2(n6834), .ZN(n6833) );
  INV_X1 U8333 ( .A(n11342), .ZN(n6834) );
  NAND2_X1 U8334 ( .A1(n6838), .A2(n6657), .ZN(n6835) );
  AND2_X1 U8335 ( .A1(n6677), .A2(n7537), .ZN(n6831) );
  INV_X1 U8336 ( .A(n6829), .ZN(n6828) );
  OAI21_X1 U8337 ( .B1(n12399), .B2(n6830), .A(n12472), .ZN(n6829) );
  INV_X1 U8338 ( .A(n9837), .ZN(n6830) );
  OR2_X1 U8339 ( .A1(n8005), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8028) );
  OR2_X1 U8340 ( .A1(n7811), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7837) );
  AND2_X1 U8341 ( .A1(n7024), .A2(n7017), .ZN(n7016) );
  NAND2_X1 U8342 ( .A1(n7019), .A2(n7021), .ZN(n7017) );
  OR2_X1 U8343 ( .A1(n10909), .A2(n10755), .ZN(n10911) );
  INV_X1 U8344 ( .A(n6965), .ZN(n11425) );
  NAND2_X1 U8345 ( .A1(n11376), .A2(n14862), .ZN(n14838) );
  INV_X1 U8346 ( .A(n11427), .ZN(n11428) );
  NAND3_X1 U8347 ( .A1(n6872), .A2(n6873), .A3(n6676), .ZN(n11378) );
  AOI21_X1 U8348 ( .B1(n14887), .B2(n14886), .A(n14885), .ZN(n14910) );
  NOR2_X1 U8349 ( .A1(n14899), .A2(n7199), .ZN(n11379) );
  NOR2_X1 U8350 ( .A1(n14914), .A2(n15009), .ZN(n7199) );
  OAI21_X1 U8351 ( .B1(n14920), .B2(n6868), .A(n6867), .ZN(n14939) );
  NAND2_X1 U8352 ( .A1(n6869), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n6868) );
  NAND2_X1 U8353 ( .A1(n11380), .A2(n6869), .ZN(n6867) );
  INV_X1 U8354 ( .A(n14940), .ZN(n6869) );
  XNOR2_X1 U8355 ( .A(n11438), .B(n11410), .ZN(n14967) );
  NAND2_X1 U8356 ( .A1(n14967), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n14966) );
  AOI21_X1 U8357 ( .B1(n14959), .B2(n14958), .A(n14957), .ZN(n14985) );
  AOI21_X1 U8358 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n14942), .A(n14939), .ZN(
        n11381) );
  OR2_X1 U8359 ( .A1(n11515), .A2(n11516), .ZN(n6875) );
  NAND2_X1 U8360 ( .A1(n11529), .A2(n11530), .ZN(n11531) );
  AND2_X1 U8361 ( .A1(n7201), .A2(n7200), .ZN(n11838) );
  NAND2_X1 U8362 ( .A1(n11586), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7200) );
  NAND2_X1 U8363 ( .A1(n6866), .A2(n6687), .ZN(n7192) );
  NAND2_X1 U8364 ( .A1(n12534), .A2(n12535), .ZN(n12558) );
  OAI21_X1 U8365 ( .B1(n12563), .B2(n12562), .A(n12561), .ZN(n12564) );
  NAND3_X1 U8366 ( .A1(n7197), .A2(n12584), .A3(P3_REG2_REG_17__SCAN_IN), .ZN(
        n7196) );
  XNOR2_X1 U8367 ( .A(n6960), .B(n6959), .ZN(n6958) );
  INV_X1 U8368 ( .A(n12603), .ZN(n6959) );
  AOI21_X1 U8369 ( .B1(n12602), .B2(n12601), .A(n6961), .ZN(n6960) );
  NOR2_X1 U8370 ( .A1(n6962), .A2(n12858), .ZN(n6961) );
  NAND2_X1 U8371 ( .A1(n9262), .A2(n7023), .ZN(n7022) );
  INV_X1 U8372 ( .A(n9261), .ZN(n7023) );
  NAND2_X1 U8373 ( .A1(n8055), .A2(n8054), .ZN(n9118) );
  OR2_X1 U8374 ( .A1(n7987), .A2(n12939), .ZN(n8054) );
  INV_X1 U8375 ( .A(n9291), .ZN(n8061) );
  AND2_X1 U8376 ( .A1(n9262), .A2(n8109), .ZN(n12336) );
  INV_X1 U8377 ( .A(n7037), .ZN(n7036) );
  OAI21_X1 U8378 ( .B1(n6660), .B2(n7038), .A(n12651), .ZN(n7037) );
  NOR2_X1 U8379 ( .A1(n7960), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7976) );
  NAND2_X1 U8380 ( .A1(n9240), .A2(n9242), .ZN(n12667) );
  AND2_X1 U8381 ( .A1(n7924), .A2(n7923), .ZN(n7939) );
  NAND2_X1 U8382 ( .A1(n12745), .A2(n6689), .ZN(n12732) );
  NAND2_X1 U8383 ( .A1(n12762), .A2(n9206), .ZN(n12744) );
  AND2_X1 U8384 ( .A1(n9207), .A2(n9206), .ZN(n12763) );
  INV_X1 U8385 ( .A(n7032), .ZN(n7031) );
  NAND2_X1 U8386 ( .A1(n7012), .A2(n9173), .ZN(n11807) );
  INV_X1 U8387 ( .A(n11723), .ZN(n7012) );
  OR2_X1 U8388 ( .A1(n7729), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7745) );
  AND2_X1 U8389 ( .A1(n11707), .A2(n9169), .ZN(n11723) );
  AND2_X1 U8390 ( .A1(n7693), .A2(n7692), .ZN(n7713) );
  NAND2_X1 U8391 ( .A1(n7713), .A2(n11885), .ZN(n7729) );
  INV_X1 U8392 ( .A(n7711), .ZN(n7453) );
  NAND2_X1 U8393 ( .A1(n7454), .A2(n7711), .ZN(n11728) );
  NAND2_X1 U8394 ( .A1(n7014), .A2(n7013), .ZN(n11707) );
  INV_X1 U8395 ( .A(n11705), .ZN(n7013) );
  NOR2_X1 U8396 ( .A1(n7673), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7693) );
  INV_X1 U8397 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n11344) );
  OAI21_X1 U8398 ( .B1(n15028), .B2(n7441), .A(n11452), .ZN(n7440) );
  NOR2_X1 U8399 ( .A1(n15029), .A2(n7441), .ZN(n7439) );
  INV_X1 U8400 ( .A(n8091), .ZN(n15014) );
  NAND2_X1 U8401 ( .A1(n8090), .A2(n9151), .ZN(n15012) );
  NAND2_X1 U8402 ( .A1(n7620), .A2(n15027), .ZN(n11453) );
  NAND2_X1 U8403 ( .A1(n15029), .A2(n15028), .ZN(n15027) );
  NAND2_X1 U8404 ( .A1(n11067), .A2(n11066), .ZN(n11069) );
  AND2_X1 U8405 ( .A1(n15058), .A2(n11053), .ZN(n15115) );
  AOI21_X1 U8406 ( .B1(n7116), .B2(n7118), .A(n6759), .ZN(n7115) );
  AND2_X1 U8407 ( .A1(n7462), .A2(n7041), .ZN(n7040) );
  NOR2_X1 U8408 ( .A1(n7042), .A2(P3_IR_REG_29__SCAN_IN), .ZN(n7041) );
  OAI22_X1 U8409 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n13490), .B1(n8053), 
        .B2(n8052), .ZN(n9098) );
  INV_X1 U8410 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7569) );
  NAND2_X1 U8411 ( .A1(n8127), .A2(n7559), .ZN(n8128) );
  XNOR2_X1 U8412 ( .A(n8154), .B(n7556), .ZN(n10751) );
  XNOR2_X1 U8413 ( .A(n7932), .B(n7920), .ZN(n7933) );
  NAND2_X1 U8414 ( .A1(n7187), .A2(n7888), .ZN(n7186) );
  INV_X1 U8415 ( .A(n7109), .ZN(n7108) );
  NAND2_X1 U8416 ( .A1(n7100), .A2(n7817), .ZN(n7102) );
  NAND2_X1 U8417 ( .A1(n7832), .A2(n7831), .ZN(n7851) );
  INV_X1 U8418 ( .A(n7830), .ZN(n7832) );
  NAND2_X1 U8419 ( .A1(n7182), .A2(n7555), .ZN(n7803) );
  INV_X1 U8420 ( .A(n7800), .ZN(n7182) );
  OR2_X1 U8421 ( .A1(n7803), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n7830) );
  OR2_X1 U8422 ( .A1(n7704), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n7705) );
  NOR2_X1 U8423 ( .A1(n7705), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7740) );
  XNOR2_X1 U8424 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n7699) );
  NAND2_X1 U8425 ( .A1(n7666), .A2(n7665), .ZN(n7681) );
  XNOR2_X1 U8426 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n7663) );
  XNOR2_X1 U8427 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n7649) );
  XNOR2_X1 U8428 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n7627) );
  XNOR2_X1 U8429 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n7611) );
  AND2_X1 U8430 ( .A1(n8271), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7594) );
  INV_X1 U8431 ( .A(n10670), .ZN(n7388) );
  AND2_X1 U8432 ( .A1(n8668), .A2(n8646), .ZN(n7404) );
  INV_X1 U8433 ( .A(n12966), .ZN(n8668) );
  AND2_X1 U8434 ( .A1(n8847), .A2(n8826), .ZN(n7405) );
  INV_X1 U8435 ( .A(n12948), .ZN(n8847) );
  NOR2_X1 U8436 ( .A1(n13074), .A2(n6942), .ZN(n6941) );
  INV_X1 U8437 ( .A(n8806), .ZN(n6942) );
  NAND2_X1 U8438 ( .A1(n8791), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n8816) );
  OR2_X1 U8439 ( .A1(n8437), .A2(n11022), .ZN(n8461) );
  OR2_X1 U8440 ( .A1(n8521), .A2(n8520), .ZN(n8543) );
  NAND2_X1 U8441 ( .A1(n8447), .A2(n8446), .ZN(n11119) );
  AND2_X1 U8442 ( .A1(n10183), .A2(n13491), .ZN(n13076) );
  AND2_X1 U8443 ( .A1(n8695), .A2(n8694), .ZN(n12969) );
  OR2_X1 U8444 ( .A1(n8579), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n8608) );
  AOI21_X1 U8445 ( .B1(n7290), .B2(n7292), .A(n6686), .ZN(n7287) );
  AND2_X1 U8446 ( .A1(n9075), .A2(n9013), .ZN(n13171) );
  NAND2_X1 U8447 ( .A1(n13189), .A2(n9012), .ZN(n7481) );
  INV_X1 U8448 ( .A(n9015), .ZN(n13164) );
  AND2_X1 U8449 ( .A1(n6634), .A2(n9074), .ZN(n7294) );
  NAND2_X1 U8450 ( .A1(n6724), .A2(n6634), .ZN(n7293) );
  INV_X1 U8451 ( .A(n7293), .ZN(n7292) );
  INV_X1 U8452 ( .A(n6821), .ZN(n6820) );
  OAI21_X1 U8453 ( .B1(n13239), .B2(n6714), .A(n9071), .ZN(n13229) );
  AND2_X1 U8454 ( .A1(n8792), .A2(n8775), .ZN(n13233) );
  NAND2_X1 U8455 ( .A1(n9010), .A2(n6643), .ZN(n7465) );
  NAND2_X1 U8456 ( .A1(n7073), .A2(n13264), .ZN(n13258) );
  AOI21_X1 U8457 ( .B1(n7300), .B2(n7302), .A(n6746), .ZN(n7297) );
  AND2_X1 U8458 ( .A1(n6806), .A2(n6805), .ZN(n13284) );
  NAND2_X1 U8459 ( .A1(n13301), .A2(n13095), .ZN(n6805) );
  NAND2_X1 U8460 ( .A1(n6808), .A2(n6807), .ZN(n6806) );
  NAND2_X1 U8461 ( .A1(n13425), .A2(n13041), .ZN(n6807) );
  NOR2_X1 U8462 ( .A1(n9006), .A2(n6809), .ZN(n13303) );
  NOR2_X1 U8463 ( .A1(n13431), .A2(n12968), .ZN(n6809) );
  NOR2_X1 U8464 ( .A1(n13315), .A2(n9005), .ZN(n9006) );
  AND2_X1 U8465 ( .A1(n13431), .A2(n12968), .ZN(n9005) );
  INV_X1 U8466 ( .A(n7305), .ZN(n7304) );
  OAI22_X1 U8467 ( .A1(n11645), .A2(n9056), .B1(n13452), .B2(n13100), .ZN(
        n11691) );
  NAND2_X1 U8468 ( .A1(n11298), .A2(n7076), .ZN(n11641) );
  NAND2_X1 U8469 ( .A1(n11298), .A2(n11486), .ZN(n11506) );
  NAND2_X1 U8470 ( .A1(n11128), .A2(n8993), .ZN(n11260) );
  OR2_X1 U8471 ( .A1(n8461), .A2(n8460), .ZN(n8481) );
  NAND2_X1 U8472 ( .A1(n11091), .A2(n8991), .ZN(n11129) );
  NAND2_X1 U8473 ( .A1(n11129), .A2(n12176), .ZN(n11128) );
  NAND2_X1 U8474 ( .A1(n10881), .A2(n7069), .ZN(n11096) );
  AND2_X1 U8475 ( .A1(n14765), .A2(n7070), .ZN(n7069) );
  NAND2_X1 U8476 ( .A1(n7316), .A2(n6667), .ZN(n7315) );
  NAND2_X1 U8477 ( .A1(n8988), .A2(n6785), .ZN(n11003) );
  AND2_X1 U8478 ( .A1(n7499), .A2(n8986), .ZN(n6785) );
  NAND2_X1 U8479 ( .A1(n7499), .A2(n8986), .ZN(n11001) );
  NAND2_X1 U8480 ( .A1(n10973), .A2(n14812), .ZN(n10996) );
  NAND2_X1 U8481 ( .A1(n7283), .A2(n9038), .ZN(n10986) );
  NAND2_X1 U8482 ( .A1(n10844), .A2(n10845), .ZN(n7283) );
  XNOR2_X1 U8483 ( .A(n7498), .B(n7497), .ZN(n12167) );
  NAND2_X1 U8484 ( .A1(n8285), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6928) );
  NAND2_X1 U8485 ( .A1(n10181), .A2(n10242), .ZN(n6927) );
  NAND2_X1 U8486 ( .A1(n10737), .A2(n8977), .ZN(n10841) );
  INV_X1 U8487 ( .A(n10845), .ZN(n12165) );
  NAND2_X1 U8488 ( .A1(n9026), .A2(n12206), .ZN(n13350) );
  INV_X1 U8489 ( .A(n8273), .ZN(n10734) );
  INV_X1 U8490 ( .A(n13350), .ZN(n13332) );
  NAND2_X1 U8491 ( .A1(n8790), .A2(n8789), .ZN(n13393) );
  NAND2_X1 U8492 ( .A1(n7471), .A2(n7469), .ZN(n13240) );
  NAND2_X1 U8493 ( .A1(n9010), .A2(n6631), .ZN(n7471) );
  NAND2_X1 U8494 ( .A1(n11258), .A2(n8994), .ZN(n11294) );
  CLKBUF_X1 U8495 ( .A(n9077), .Z(n14815) );
  AND2_X1 U8496 ( .A1(n12161), .A2(n12131), .ZN(n14822) );
  INV_X1 U8497 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7379) );
  INV_X1 U8498 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8864) );
  NAND3_X1 U8499 ( .A1(n8727), .A2(n8728), .A3(n8744), .ZN(n8745) );
  INV_X1 U8500 ( .A(n8729), .ZN(n8728) );
  NAND2_X1 U8501 ( .A1(n11872), .A2(n7137), .ZN(n7133) );
  AND2_X1 U8502 ( .A1(n7135), .A2(n12225), .ZN(n7134) );
  NOR2_X1 U8503 ( .A1(n9580), .A2(n15330), .ZN(n9593) );
  AOI21_X1 U8504 ( .B1(n7147), .B2(n6658), .A(n7146), .ZN(n7145) );
  NOR2_X1 U8505 ( .A1(n11321), .A2(n11322), .ZN(n7146) );
  INV_X1 U8506 ( .A(n11323), .ZN(n7147) );
  NAND2_X1 U8507 ( .A1(n6774), .A2(n7148), .ZN(n7144) );
  NAND2_X1 U8508 ( .A1(n13562), .A2(n13563), .ZN(n13561) );
  INV_X1 U8509 ( .A(n9628), .ZN(n9618) );
  AND2_X1 U8510 ( .A1(n11787), .A2(n11788), .ZN(n11785) );
  NAND2_X1 U8511 ( .A1(n13580), .A2(n13581), .ZN(n13579) );
  CLKBUF_X1 U8512 ( .A(n11674), .Z(n11667) );
  AOI21_X1 U8513 ( .B1(n12313), .B2(n14013), .A(n10349), .ZN(n10350) );
  AND2_X1 U8514 ( .A1(n10365), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10349) );
  NAND2_X1 U8515 ( .A1(n9593), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9604) );
  OR2_X1 U8516 ( .A1(n11173), .A2(n11170), .ZN(n11174) );
  INV_X1 U8517 ( .A(n10175), .ZN(n10357) );
  AND4_X1 U8518 ( .A1(n9530), .A2(n9529), .A3(n9528), .A4(n9527), .ZN(n12229)
         );
  INV_X1 U8519 ( .A(n6972), .ZN(n6971) );
  OAI21_X1 U8520 ( .B1(n6717), .B2(n13842), .A(n6973), .ZN(n6972) );
  NAND2_X1 U8521 ( .A1(n6722), .A2(n7326), .ZN(n6973) );
  AND2_X1 U8522 ( .A1(n10105), .A2(n6638), .ZN(n7364) );
  INV_X1 U8523 ( .A(n7367), .ZN(n7363) );
  NAND2_X1 U8524 ( .A1(n7332), .A2(n6898), .ZN(n6895) );
  NAND2_X1 U8525 ( .A1(n7331), .A2(n7334), .ZN(n7330) );
  OAI21_X1 U8526 ( .B1(n13841), .B2(n7336), .A(n13837), .ZN(n7331) );
  NAND2_X1 U8527 ( .A1(n7332), .A2(n6894), .ZN(n6893) );
  NOR2_X1 U8528 ( .A1(n13868), .A2(n6896), .ZN(n6894) );
  AND2_X1 U8529 ( .A1(n9656), .A2(n9330), .ZN(n13830) );
  NAND2_X1 U8530 ( .A1(n13896), .A2(n7204), .ZN(n13827) );
  NOR2_X1 U8531 ( .A1(n14042), .A2(n7205), .ZN(n7204) );
  INV_X1 U8532 ( .A(n7206), .ZN(n7205) );
  NAND2_X1 U8533 ( .A1(n13896), .A2(n7207), .ZN(n13863) );
  NAND2_X1 U8534 ( .A1(n13896), .A2(n13885), .ZN(n13879) );
  NAND2_X1 U8535 ( .A1(n6876), .A2(n7339), .ZN(n13875) );
  INV_X1 U8536 ( .A(n7340), .ZN(n7339) );
  NAND2_X1 U8537 ( .A1(n13924), .A2(n7341), .ZN(n6876) );
  OAI22_X1 U8538 ( .A1(n13892), .A2(n6666), .B1(n14077), .B2(n14071), .ZN(
        n7340) );
  NOR2_X1 U8539 ( .A1(n13875), .A2(n13876), .ZN(n13874) );
  NOR2_X1 U8540 ( .A1(n13913), .A2(n13927), .ZN(n13910) );
  AND2_X1 U8541 ( .A1(n14071), .A2(n13910), .ZN(n13896) );
  INV_X1 U8542 ( .A(n9645), .ZN(n9635) );
  NAND2_X1 U8543 ( .A1(n14000), .A2(n13985), .ZN(n13980) );
  NAND2_X1 U8544 ( .A1(n9560), .A2(n9559), .ZN(n13990) );
  OR2_X1 U8545 ( .A1(n14371), .A2(n12244), .ZN(n13997) );
  NOR2_X1 U8546 ( .A1(n9525), .A2(n9524), .ZN(n9540) );
  INV_X1 U8547 ( .A(n7220), .ZN(n14311) );
  NAND2_X1 U8548 ( .A1(n14386), .A2(n11467), .ZN(n14309) );
  AOI21_X1 U8549 ( .B1(n14384), .B2(n7357), .A(n6694), .ZN(n7356) );
  NAND2_X1 U8550 ( .A1(n11307), .A2(n9749), .ZN(n14378) );
  NOR2_X1 U8551 ( .A1(n11311), .A2(n14383), .ZN(n14386) );
  OR2_X1 U8552 ( .A1(n9468), .A2(n11677), .ZN(n9484) );
  NAND2_X1 U8553 ( .A1(n14510), .A2(n7218), .ZN(n11312) );
  AND2_X1 U8554 ( .A1(n6635), .A2(n14627), .ZN(n7218) );
  NAND2_X1 U8555 ( .A1(n14510), .A2(n6635), .ZN(n11106) );
  AND4_X1 U8556 ( .A1(n9448), .A2(n9447), .A3(n9446), .A4(n9445), .ZN(n11607)
         );
  AND4_X1 U8557 ( .A1(n9459), .A2(n9458), .A3(n9457), .A4(n9456), .ZN(n11678)
         );
  NAND2_X1 U8558 ( .A1(n13670), .A2(n7323), .ZN(n7322) );
  OR2_X1 U8559 ( .A1(n10899), .A2(n9747), .ZN(n7320) );
  AND3_X1 U8560 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n9418) );
  INV_X1 U8561 ( .A(n9405), .ZN(n7351) );
  NOR2_X1 U8562 ( .A1(n14524), .A2(n11180), .ZN(n14510) );
  NAND2_X1 U8563 ( .A1(n14530), .A2(n10086), .ZN(n9742) );
  NOR2_X1 U8564 ( .A1(n14543), .A2(n6626), .ZN(n14544) );
  NAND2_X1 U8565 ( .A1(n9378), .A2(n9377), .ZN(n14529) );
  OR2_X1 U8566 ( .A1(n14558), .A2(n14013), .ZN(n10723) );
  OR2_X1 U8567 ( .A1(n10341), .A2(n13930), .ZN(n10516) );
  AND2_X1 U8568 ( .A1(n11945), .A2(n9327), .ZN(n9380) );
  NAND2_X1 U8569 ( .A1(n10706), .A2(n14013), .ZN(n9884) );
  NAND2_X1 U8570 ( .A1(n9671), .A2(n9670), .ZN(n14028) );
  NAND2_X1 U8571 ( .A1(n13924), .A2(n9758), .ZN(n13907) );
  NAND2_X1 U8572 ( .A1(n9523), .A2(n9522), .ZN(n14414) );
  NAND2_X1 U8573 ( .A1(n7319), .A2(n7318), .ZN(n11108) );
  AND2_X1 U8574 ( .A1(n6883), .A2(n6734), .ZN(n7318) );
  INV_X1 U8575 ( .A(n10341), .ZN(n14559) );
  INV_X1 U8576 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n15343) );
  AND2_X1 U8577 ( .A1(n9321), .A2(n9319), .ZN(n7373) );
  XNOR2_X1 U8578 ( .A(n9324), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9328) );
  NAND2_X1 U8579 ( .A1(n14139), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9324) );
  XNOR2_X1 U8580 ( .A(n9320), .B(n9319), .ZN(n9720) );
  NAND2_X1 U8581 ( .A1(n9323), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9320) );
  AND2_X1 U8582 ( .A1(n9683), .A2(n9321), .ZN(n7372) );
  NAND2_X1 U8583 ( .A1(n7347), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7346) );
  NAND2_X1 U8584 ( .A1(n8745), .A2(n8744), .ZN(n8764) );
  NAND2_X1 U8585 ( .A1(n8727), .A2(n8744), .ZN(n9625) );
  AND2_X1 U8586 ( .A1(n7281), .A2(n7280), .ZN(n7279) );
  NOR2_X1 U8587 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n7280) );
  NAND2_X1 U8588 ( .A1(n8682), .A2(SI_20_), .ZN(n6988) );
  NOR2_X1 U8589 ( .A1(n6989), .A2(n6987), .ZN(n6986) );
  AND2_X1 U8590 ( .A1(n8723), .A2(n8705), .ZN(n8706) );
  NAND2_X1 U8591 ( .A1(n9716), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9713) );
  INV_X1 U8592 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9702) );
  XNOR2_X1 U8593 ( .A(n8495), .B(n8494), .ZN(n10490) );
  NAND2_X1 U8594 ( .A1(n8475), .A2(n8474), .ZN(n8495) );
  NAND2_X1 U8595 ( .A1(n8454), .A2(n8453), .ZN(n8475) );
  INV_X1 U8596 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9462) );
  AND2_X1 U8597 ( .A1(n8448), .A2(n8424), .ZN(n8425) );
  NAND2_X1 U8598 ( .A1(n8426), .A2(n8425), .ZN(n8449) );
  AND2_X1 U8599 ( .A1(n8420), .A2(n8401), .ZN(n8402) );
  OR2_X1 U8600 ( .A1(n9439), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9450) );
  OR2_X1 U8601 ( .A1(n9400), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9536) );
  NAND2_X1 U8602 ( .A1(n8300), .A2(n8299), .ZN(n8305) );
  NAND2_X1 U8603 ( .A1(n8252), .A2(n8225), .ZN(n8231) );
  NAND2_X1 U8604 ( .A1(n14166), .A2(n7053), .ZN(n14207) );
  NAND2_X1 U8605 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n7054), .ZN(n7053) );
  INV_X1 U8606 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7054) );
  XNOR2_X1 U8607 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n14208) );
  NAND2_X1 U8608 ( .A1(n7058), .A2(n14230), .ZN(n14232) );
  NAND2_X1 U8609 ( .A1(n14280), .A2(n14279), .ZN(n7058) );
  NOR2_X1 U8610 ( .A1(n14237), .A2(n14238), .ZN(n14241) );
  OAI21_X1 U8611 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n14186), .A(n14185), .ZN(
        n14199) );
  AOI21_X1 U8612 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n14188), .A(n14187), .ZN(
        n14249) );
  NOR2_X1 U8613 ( .A1(n14200), .A2(n14199), .ZN(n14187) );
  NAND2_X1 U8614 ( .A1(n14455), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7063) );
  NAND2_X1 U8615 ( .A1(n11492), .A2(n9781), .ZN(n11686) );
  XOR2_X1 U8616 ( .A(n12721), .B(n9809), .Z(n12370) );
  NAND2_X1 U8617 ( .A1(n12416), .A2(n7166), .ZN(n6841) );
  OR2_X1 U8618 ( .A1(n11685), .A2(n11763), .ZN(n9782) );
  NAND2_X1 U8619 ( .A1(n11762), .A2(n11761), .ZN(n11760) );
  NAND2_X1 U8620 ( .A1(n7937), .A2(n7936), .ZN(n12383) );
  OR2_X1 U8621 ( .A1(n7735), .A2(n10981), .ZN(n7936) );
  NAND2_X1 U8622 ( .A1(n7857), .A2(n7856), .ZN(n12779) );
  AND2_X1 U8623 ( .A1(n6832), .A2(n6677), .ZN(n6837) );
  INV_X1 U8624 ( .A(n10685), .ZN(n12792) );
  INV_X1 U8625 ( .A(n12397), .ZN(n12428) );
  NAND2_X1 U8626 ( .A1(n7175), .A2(n7174), .ZN(n11273) );
  AND2_X1 U8627 ( .A1(n7175), .A2(n6675), .ZN(n11274) );
  NAND2_X1 U8628 ( .A1(n11760), .A2(n9785), .ZN(n11883) );
  XNOR2_X1 U8629 ( .A(n9810), .B(n12733), .ZN(n12435) );
  NOR2_X1 U8630 ( .A1(n11073), .A2(n9772), .ZN(n11044) );
  NAND2_X1 U8631 ( .A1(n7600), .A2(n7599), .ZN(n7601) );
  NAND2_X1 U8632 ( .A1(n12416), .A2(n12417), .ZN(n7165) );
  INV_X1 U8633 ( .A(n12485), .ZN(n12467) );
  NAND2_X1 U8634 ( .A1(n11494), .A2(n11493), .ZN(n11492) );
  NAND2_X1 U8635 ( .A1(n6835), .A2(n6833), .ZN(n11494) );
  NAND2_X1 U8636 ( .A1(n9865), .A2(n15059), .ZN(n12490) );
  INV_X1 U8637 ( .A(n12473), .ZN(n12495) );
  AND2_X1 U8638 ( .A1(n9112), .A2(n8080), .ZN(n11014) );
  INV_X1 U8639 ( .A(n12477), .ZN(n12499) );
  INV_X1 U8640 ( .A(n12699), .ZN(n12668) );
  NAND2_X1 U8641 ( .A1(n7622), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7590) );
  NAND2_X1 U8642 ( .A1(n7434), .A2(n7002), .ZN(n7437) );
  NAND2_X1 U8643 ( .A1(n7436), .A2(n7435), .ZN(n7434) );
  OR2_X1 U8644 ( .A1(n7675), .A2(n10757), .ZN(n7581) );
  INV_X2 U8645 ( .A(P3_U3897), .ZN(n12506) );
  NOR2_X1 U8646 ( .A1(n10922), .A2(n10923), .ZN(n10921) );
  INV_X1 U8647 ( .A(n6966), .ZN(n10779) );
  NOR2_X1 U8648 ( .A1(n14838), .A2(n15036), .ZN(n14866) );
  NOR2_X1 U8649 ( .A1(n14920), .A2(n14921), .ZN(n14919) );
  NAND2_X1 U8650 ( .A1(n14930), .A2(n11435), .ZN(n14938) );
  XNOR2_X1 U8651 ( .A(n11514), .B(n11521), .ZN(n11383) );
  INV_X1 U8652 ( .A(n7201), .ZN(n11584) );
  INV_X1 U8653 ( .A(n6875), .ZN(n11519) );
  XNOR2_X1 U8654 ( .A(n11838), .B(n11852), .ZN(n11585) );
  INV_X1 U8655 ( .A(n7192), .ZN(n12531) );
  INV_X1 U8656 ( .A(n7196), .ZN(n12588) );
  NAND2_X1 U8657 ( .A1(n8043), .A2(n8042), .ZN(n12631) );
  INV_X1 U8658 ( .A(n8953), .ZN(n8954) );
  NAND2_X1 U8659 ( .A1(n8939), .A2(n8938), .ZN(n8942) );
  NAND2_X1 U8660 ( .A1(n12664), .A2(n9242), .ZN(n12652) );
  AND2_X1 U8661 ( .A1(n7974), .A2(n7973), .ZN(n12675) );
  NAND2_X1 U8662 ( .A1(n7959), .A2(n7958), .ZN(n12689) );
  OR2_X1 U8663 ( .A1(n7987), .A2(n11206), .ZN(n7958) );
  NAND2_X1 U8664 ( .A1(n12717), .A2(n9222), .ZN(n12706) );
  NAND2_X1 U8665 ( .A1(n12718), .A2(n7931), .ZN(n12707) );
  NAND2_X1 U8666 ( .A1(n12742), .A2(n9208), .ZN(n12731) );
  NAND2_X1 U8667 ( .A1(n12760), .A2(n7882), .ZN(n12747) );
  NAND2_X1 U8668 ( .A1(n7442), .A2(n7844), .ZN(n12775) );
  NAND2_X1 U8669 ( .A1(n12789), .A2(n12790), .ZN(n7442) );
  NAND2_X1 U8670 ( .A1(n7009), .A2(n7007), .ZN(n12786) );
  NAND2_X1 U8671 ( .A1(n7009), .A2(n9188), .ZN(n12798) );
  NAND2_X1 U8672 ( .A1(n11896), .A2(n9178), .ZN(n14338) );
  NAND2_X1 U8673 ( .A1(n15034), .A2(n14345), .ZN(n12818) );
  AND2_X1 U8674 ( .A1(n7035), .A2(n9172), .ZN(n11898) );
  INV_X1 U8675 ( .A(n12822), .ZN(n14340) );
  NOR2_X1 U8676 ( .A1(n11069), .A2(n15058), .ZN(n15034) );
  AND2_X1 U8677 ( .A1(n12595), .A2(n10875), .ZN(n15058) );
  AND2_X2 U8678 ( .A1(n10749), .A2(n9852), .ZN(n15071) );
  AND2_X1 U8679 ( .A1(n15058), .A2(n14345), .ZN(n9852) );
  AND2_X1 U8680 ( .A1(n14344), .A2(n14348), .ZN(n14354) );
  AND2_X1 U8681 ( .A1(n14348), .A2(n14347), .ZN(n14356) );
  AND2_X1 U8682 ( .A1(n12619), .A2(n15101), .ZN(n8115) );
  OR2_X1 U8683 ( .A1(n7735), .A2(n11941), .ZN(n7988) );
  INV_X1 U8684 ( .A(n12396), .ZN(n12886) );
  INV_X1 U8685 ( .A(n12383), .ZN(n12896) );
  NAND2_X1 U8686 ( .A1(n7908), .A2(n7907), .ZN(n12901) );
  NAND2_X1 U8687 ( .A1(n7807), .A2(n7806), .ZN(n12922) );
  NAND2_X1 U8688 ( .A1(n15119), .A2(n14345), .ZN(n12926) );
  INV_X1 U8689 ( .A(n11046), .ZN(n11938) );
  AOI21_X1 U8690 ( .B1(n8123), .B2(P3_IR_REG_25__SCAN_IN), .A(n8122), .ZN(
        n8124) );
  AND2_X1 U8691 ( .A1(n8127), .A2(n7558), .ZN(n8122) );
  AOI21_X1 U8692 ( .B1(n8118), .B2(P3_IR_REG_24__SCAN_IN), .A(n8117), .ZN(
        n8119) );
  AND2_X1 U8693 ( .A1(n8127), .A2(n7557), .ZN(n8117) );
  INV_X1 U8694 ( .A(SI_23_), .ZN(n11206) );
  NAND2_X1 U8695 ( .A1(n7082), .A2(n7084), .ZN(n7956) );
  NAND2_X1 U8696 ( .A1(n7945), .A2(n7946), .ZN(n7082) );
  XNOR2_X1 U8697 ( .A(n8073), .B(n8072), .ZN(n10980) );
  INV_X1 U8698 ( .A(SI_19_), .ZN(n10596) );
  INV_X1 U8699 ( .A(SI_18_), .ZN(n10595) );
  NAND2_X1 U8700 ( .A1(n7107), .A2(n7868), .ZN(n7884) );
  NAND2_X1 U8701 ( .A1(n7867), .A2(n7866), .ZN(n7107) );
  NAND2_X1 U8702 ( .A1(n7818), .A2(n7817), .ZN(n7826) );
  INV_X1 U8703 ( .A(SI_13_), .ZN(n10301) );
  INV_X1 U8704 ( .A(SI_12_), .ZN(n10169) );
  NAND2_X1 U8705 ( .A1(n7096), .A2(n7094), .ZN(n7797) );
  NAND2_X1 U8706 ( .A1(n7096), .A2(n7774), .ZN(n7779) );
  INV_X1 U8707 ( .A(n11594), .ZN(n11586) );
  INV_X1 U8708 ( .A(SI_11_), .ZN(n10151) );
  NAND2_X1 U8709 ( .A1(n7756), .A2(n7755), .ZN(n7776) );
  NAND2_X1 U8710 ( .A1(n7087), .A2(n7723), .ZN(n7737) );
  NAND2_X1 U8711 ( .A1(n7721), .A2(n7720), .ZN(n7087) );
  INV_X1 U8712 ( .A(n14892), .ZN(n11431) );
  NAND2_X1 U8713 ( .A1(n13071), .A2(n7405), .ZN(n12947) );
  NAND2_X1 U8714 ( .A1(n8554), .A2(n8555), .ZN(n11578) );
  NAND2_X1 U8715 ( .A1(n7402), .A2(n8530), .ZN(n11575) );
  XNOR2_X1 U8716 ( .A(n8759), .B(n8757), .ZN(n12957) );
  NAND2_X1 U8717 ( .A1(n7385), .A2(n8472), .ZN(n11120) );
  INV_X1 U8718 ( .A(n11119), .ZN(n7385) );
  NAND2_X1 U8719 ( .A1(n8647), .A2(n8646), .ZN(n12967) );
  OAI21_X1 U8720 ( .B1(n13377), .B2(n7401), .A(n7395), .ZN(n7394) );
  NAND2_X1 U8721 ( .A1(n8915), .A2(n7401), .ZN(n7395) );
  AND2_X1 U8722 ( .A1(n7398), .A2(n7397), .ZN(n7396) );
  OR2_X1 U8723 ( .A1(n13377), .A2(n8862), .ZN(n7398) );
  NAND2_X1 U8724 ( .A1(n8915), .A2(n8862), .ZN(n7397) );
  AOI21_X1 U8725 ( .B1(n8915), .B2(n13083), .A(n7400), .ZN(n7399) );
  NOR2_X1 U8726 ( .A1(n13377), .A2(n13049), .ZN(n7400) );
  NAND2_X1 U8727 ( .A1(n8501), .A2(n8500), .ZN(n12035) );
  NAND2_X1 U8728 ( .A1(n13027), .A2(n8324), .ZN(n10627) );
  NAND2_X1 U8729 ( .A1(n10627), .A2(n10628), .ZN(n10626) );
  INV_X1 U8730 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n11022) );
  CLKBUF_X1 U8731 ( .A(n11019), .Z(n11021) );
  NAND2_X1 U8732 ( .A1(n8273), .A2(n8272), .ZN(n10321) );
  CLKBUF_X1 U8733 ( .A(n11286), .Z(n11287) );
  NAND2_X1 U8734 ( .A1(n11120), .A2(n8473), .ZN(n11196) );
  OR2_X1 U8735 ( .A1(n8925), .A2(n12213), .ZN(n13079) );
  NAND2_X1 U8736 ( .A1(n12984), .A2(n8806), .ZN(n13073) );
  NAND2_X1 U8737 ( .A1(n8870), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8215) );
  NAND2_X1 U8738 ( .A1(n10183), .A2(n8918), .ZN(n13060) );
  INV_X1 U8739 ( .A(n12131), .ZN(n12215) );
  NAND4_X1 U8740 ( .A1(n8243), .A2(n8242), .A3(n8241), .A4(n8240), .ZN(n13111)
         );
  OR2_X1 U8741 ( .A1(n8545), .A2(n6767), .ZN(n8243) );
  OR2_X2 U8742 ( .A1(n10182), .A2(P2_U3088), .ZN(n13113) );
  NAND2_X1 U8743 ( .A1(n12139), .A2(n12138), .ZN(n13370) );
  NAND2_X1 U8744 ( .A1(n7472), .A2(n7476), .ZN(n13255) );
  OR2_X1 U8745 ( .A1(n9010), .A2(n9009), .ZN(n7472) );
  NAND2_X1 U8746 ( .A1(n7299), .A2(n9068), .ZN(n13267) );
  NAND2_X1 U8747 ( .A1(n9067), .A2(n6632), .ZN(n7299) );
  NAND2_X1 U8748 ( .A1(n9067), .A2(n12188), .ZN(n13282) );
  NAND2_X1 U8749 ( .A1(n7488), .A2(n7493), .ZN(n13330) );
  NAND2_X1 U8750 ( .A1(n11693), .A2(n7494), .ZN(n7488) );
  NAND2_X1 U8751 ( .A1(n13347), .A2(n9060), .ZN(n13328) );
  NAND2_X1 U8752 ( .A1(n8582), .A2(n8581), .ZN(n13440) );
  NAND2_X1 U8753 ( .A1(n8563), .A2(n8562), .ZN(n12052) );
  NAND2_X1 U8754 ( .A1(n11502), .A2(n8998), .ZN(n11637) );
  NAND2_X1 U8755 ( .A1(n7503), .A2(n7504), .ZN(n10930) );
  NAND2_X1 U8756 ( .A1(n7317), .A2(n9042), .ZN(n10968) );
  NAND2_X1 U8757 ( .A1(n10584), .A2(n9041), .ZN(n7317) );
  NAND2_X1 U8758 ( .A1(n8984), .A2(n8983), .ZN(n10969) );
  CLKBUF_X1 U8759 ( .A(n13338), .Z(n14757) );
  NAND2_X1 U8760 ( .A1(n10181), .A2(n14679), .ZN(n7067) );
  OR2_X1 U8761 ( .A1(n10124), .A2(n12125), .ZN(n7066) );
  INV_X2 U8762 ( .A(n13357), .ZN(n14761) );
  OR2_X1 U8763 ( .A1(n11964), .A2(n13456), .ZN(n7313) );
  NAND2_X1 U8764 ( .A1(n13384), .A2(n6682), .ZN(n13461) );
  NAND2_X1 U8765 ( .A1(n13383), .A2(n6745), .ZN(n6777) );
  AND2_X1 U8766 ( .A1(n10184), .A2(n8903), .ZN(n14781) );
  CLKBUF_X1 U8767 ( .A(n13476), .Z(n13477) );
  INV_X1 U8768 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8236) );
  INV_X1 U8769 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13490) );
  NAND2_X1 U8770 ( .A1(n8881), .A2(n8880), .ZN(n13502) );
  XNOR2_X1 U8771 ( .A(n8875), .B(n8874), .ZN(n13506) );
  INV_X1 U8772 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8874) );
  INV_X1 U8773 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n15235) );
  INV_X1 U8774 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11226) );
  INV_X1 U8775 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10838) );
  INV_X1 U8776 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10808) );
  INV_X1 U8777 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10625) );
  INV_X1 U8778 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10492) );
  AND2_X1 U8779 ( .A1(n8409), .A2(n8428), .ZN(n10309) );
  INV_X1 U8780 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10147) );
  INV_X1 U8781 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10141) );
  NAND2_X1 U8782 ( .A1(n7527), .A2(n8198), .ZN(n8307) );
  CLKBUF_X1 U8783 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n13507) );
  AOI21_X1 U8784 ( .B1(n7130), .B2(n7132), .A(n6695), .ZN(n7127) );
  CLKBUF_X1 U8785 ( .A(n11749), .Z(n11753) );
  NAND2_X1 U8786 ( .A1(n7144), .A2(n7145), .ZN(n11333) );
  NAND2_X1 U8787 ( .A1(n11750), .A2(n11785), .ZN(n11873) );
  CLKBUF_X1 U8788 ( .A(n11786), .Z(n11750) );
  AND2_X1 U8789 ( .A1(n13579), .A2(n12250), .ZN(n13594) );
  OR2_X1 U8790 ( .A1(n13656), .A2(n14408), .ZN(n13647) );
  OR2_X1 U8791 ( .A1(n13656), .A2(n14410), .ZN(n13646) );
  OR2_X1 U8792 ( .A1(n12269), .A2(n12268), .ZN(n7542) );
  NAND2_X1 U8793 ( .A1(n11873), .A2(n11872), .ZN(n12226) );
  NAND2_X1 U8794 ( .A1(n7150), .A2(n7153), .ZN(n13632) );
  NAND2_X1 U8795 ( .A1(n13580), .A2(n7155), .ZN(n7150) );
  CLKBUF_X1 U8796 ( .A(n11214), .Z(n6774) );
  NAND2_X1 U8797 ( .A1(n10960), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13645) );
  NAND2_X1 U8798 ( .A1(n7129), .A2(n12306), .ZN(n13641) );
  NAND2_X1 U8799 ( .A1(n13570), .A2(n13571), .ZN(n7129) );
  NAND2_X1 U8800 ( .A1(n9343), .A2(n9342), .ZN(n13851) );
  NAND2_X1 U8801 ( .A1(n7272), .A2(n10085), .ZN(n7269) );
  INV_X1 U8802 ( .A(n10958), .ZN(n14584) );
  NAND4_X1 U8803 ( .A1(n9398), .A2(n9397), .A3(n9396), .A4(n9395), .ZN(n13671)
         );
  NAND2_X1 U8804 ( .A1(n10073), .A2(n10072), .ZN(n14019) );
  NAND2_X1 U8805 ( .A1(n7360), .A2(n6688), .ZN(n14060) );
  NAND2_X1 U8806 ( .A1(n7360), .A2(n9650), .ZN(n13867) );
  INV_X1 U8807 ( .A(n14066), .ZN(n13885) );
  NAND2_X1 U8808 ( .A1(n13895), .A2(n9641), .ZN(n13872) );
  AND2_X1 U8809 ( .A1(n7345), .A2(n6666), .ZN(n13888) );
  NAND2_X1 U8810 ( .A1(n13921), .A2(n9624), .ZN(n13905) );
  NAND2_X1 U8811 ( .A1(n14093), .A2(n9614), .ZN(n13923) );
  AND2_X1 U8812 ( .A1(n13953), .A2(n9987), .ZN(n13939) );
  AND2_X1 U8813 ( .A1(n13974), .A2(n9756), .ZN(n13955) );
  NAND2_X1 U8814 ( .A1(n11907), .A2(n9754), .ZN(n13992) );
  NAND2_X1 U8815 ( .A1(n14361), .A2(n9962), .ZN(n11905) );
  NAND2_X1 U8816 ( .A1(n9539), .A2(n9538), .ZN(n14366) );
  NAND2_X1 U8817 ( .A1(n9517), .A2(n9516), .ZN(n11656) );
  NAND2_X1 U8818 ( .A1(n11464), .A2(n9751), .ZN(n14303) );
  NAND2_X1 U8819 ( .A1(n9508), .A2(n9507), .ZN(n14310) );
  NAND2_X1 U8820 ( .A1(n7359), .A2(n9475), .ZN(n14385) );
  NAND2_X1 U8821 ( .A1(n11306), .A2(n11310), .ZN(n7359) );
  NAND2_X1 U8822 ( .A1(n11154), .A2(n9748), .ZN(n11309) );
  NAND2_X1 U8823 ( .A1(n9406), .A2(n9405), .ZN(n14514) );
  OR2_X1 U8824 ( .A1(n14552), .A2(n10355), .ZN(n14541) );
  INV_X1 U8825 ( .A(n14541), .ZN(n14382) );
  INV_X1 U8826 ( .A(n14009), .ZN(n14390) );
  INV_X1 U8827 ( .A(n14006), .ZN(n14552) );
  INV_X1 U8828 ( .A(n13962), .ZN(n14538) );
  INV_X1 U8829 ( .A(n14665), .ZN(n14662) );
  AOI21_X1 U8830 ( .B1(n6652), .B2(n14642), .A(n14035), .ZN(n14036) );
  AND2_X1 U8831 ( .A1(n9708), .A2(n9707), .ZN(n10515) );
  AND2_X1 U8832 ( .A1(n10344), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9707) );
  NAND2_X1 U8833 ( .A1(n9676), .A2(n7370), .ZN(n14139) );
  AND2_X1 U8834 ( .A1(n7373), .A2(n7371), .ZN(n7370) );
  NOR2_X1 U8835 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n7371) );
  NAND2_X1 U8836 ( .A1(n10066), .A2(n10045), .ZN(n13485) );
  NAND2_X1 U8837 ( .A1(n7423), .A2(n7421), .ZN(n10066) );
  NAND2_X1 U8838 ( .A1(n7423), .A2(n10041), .ZN(n10044) );
  INV_X1 U8839 ( .A(n9328), .ZN(n11945) );
  INV_X1 U8840 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14144) );
  CLKBUF_X1 U8841 ( .A(n9720), .Z(n9721) );
  CLKBUF_X1 U8842 ( .A(n9722), .Z(n14150) );
  XNOR2_X1 U8843 ( .A(n8831), .B(n8830), .ZN(n14149) );
  AND2_X1 U8844 ( .A1(n6991), .A2(n6993), .ZN(n8831) );
  NAND2_X1 U8845 ( .A1(n6995), .A2(n7430), .ZN(n6993) );
  INV_X1 U8846 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15324) );
  INV_X1 U8847 ( .A(n9706), .ZN(n14155) );
  NAND2_X1 U8848 ( .A1(n7432), .A2(n8787), .ZN(n8788) );
  NAND2_X1 U8849 ( .A1(n6764), .A2(n6763), .ZN(n9680) );
  NAND2_X1 U8850 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n9674), .ZN(n6763) );
  NAND2_X1 U8851 ( .A1(n6765), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n6764) );
  NAND2_X1 U8852 ( .A1(n6721), .A2(n8701), .ZN(n8702) );
  NOR2_X1 U8853 ( .A1(n9712), .A2(n7125), .ZN(n7124) );
  OR2_X1 U8854 ( .A1(n9715), .A2(n7282), .ZN(n7126) );
  NOR2_X1 U8855 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n7125) );
  NAND2_X1 U8856 ( .A1(n8649), .A2(n8628), .ZN(n11141) );
  NAND2_X1 U8857 ( .A1(n8602), .A2(n8601), .ZN(n8606) );
  NAND2_X1 U8858 ( .A1(n6975), .A2(n6979), .ZN(n8602) );
  INV_X1 U8859 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10840) );
  INV_X1 U8860 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n11016) );
  INV_X1 U8861 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10683) );
  INV_X1 U8862 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10622) );
  INV_X1 U8863 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10494) );
  INV_X1 U8864 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10180) );
  NAND2_X1 U8865 ( .A1(n8398), .A2(n6900), .ZN(n10179) );
  NAND2_X1 U8866 ( .A1(n8376), .A2(n6901), .ZN(n6900) );
  NOR2_X1 U8867 ( .A1(n8380), .A2(n6936), .ZN(n6901) );
  INV_X1 U8868 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10171) );
  NAND2_X1 U8869 ( .A1(n8221), .A2(n8225), .ZN(n8250) );
  NAND2_X1 U8870 ( .A1(n7311), .A2(SI_0_), .ZN(n9362) );
  CLKBUF_X1 U8871 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n6762) );
  NAND2_X1 U8872 ( .A1(n14213), .A2(n14214), .ZN(n14276) );
  NAND2_X1 U8873 ( .A1(n15525), .A2(n15526), .ZN(n14213) );
  NOR2_X1 U8874 ( .A1(n14219), .A2(n15522), .ZN(n15515) );
  XNOR2_X1 U8875 ( .A(n14227), .B(n7059), .ZN(n14280) );
  INV_X1 U8876 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7059) );
  XNOR2_X1 U8877 ( .A(n14232), .B(n7057), .ZN(n15520) );
  INV_X1 U8878 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7057) );
  XNOR2_X1 U8879 ( .A(n14241), .B(n7056), .ZN(n14282) );
  INV_X1 U8880 ( .A(n14242), .ZN(n7056) );
  AND2_X1 U8881 ( .A1(n14261), .A2(n14260), .ZN(n14457) );
  NOR2_X1 U8882 ( .A1(n14461), .A2(n14462), .ZN(n14460) );
  NAND2_X1 U8883 ( .A1(n14263), .A2(n14463), .ZN(n7048) );
  OAI21_X1 U8884 ( .B1(n12639), .B2(n12485), .A(n9870), .ZN(n9871) );
  OAI21_X1 U8885 ( .B1(n7121), .B2(n9299), .A(n9298), .ZN(n9305) );
  INV_X1 U8886 ( .A(n7190), .ZN(n14972) );
  INV_X1 U8887 ( .A(n6871), .ZN(n11843) );
  INV_X1 U8888 ( .A(n6866), .ZN(n12528) );
  INV_X1 U8889 ( .A(n6780), .ZN(n6779) );
  NAND2_X1 U8890 ( .A1(n12609), .A2(n14960), .ZN(n6963) );
  OAI21_X1 U8891 ( .B1(n13027), .B2(n7392), .A(n7389), .ZN(n10671) );
  AOI211_X1 U8892 ( .C1(n13387), .C2(n13338), .A(n13208), .B(n13207), .ZN(
        n13209) );
  OR2_X1 U8893 ( .A1(n10344), .A2(P1_U3086), .ZN(n10120) );
  OR2_X1 U8894 ( .A1(n9763), .A2(n9762), .ZN(P1_U3356) );
  AOI21_X1 U8895 ( .B1(n9736), .B2(n14014), .A(n9735), .ZN(n9737) );
  NAND2_X1 U8896 ( .A1(n7215), .A2(n6756), .ZN(P1_U3557) );
  NAND2_X1 U8897 ( .A1(n14124), .A2(n14665), .ZN(n7215) );
  INV_X1 U8898 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7214) );
  NOR2_X1 U8899 ( .A1(n14454), .A2(n14455), .ZN(n14453) );
  AND2_X1 U8900 ( .A1(n7065), .A2(n7064), .ZN(n14454) );
  NOR2_X1 U8901 ( .A1(n14323), .A2(n14322), .ZN(n14331) );
  AND4_X2 U8902 ( .A1(n6760), .A2(n7550), .A3(n7552), .A4(n7553), .ZN(n6629)
         );
  NAND2_X1 U8903 ( .A1(n12892), .A2(n12711), .ZN(n6630) );
  INV_X1 U8904 ( .A(n14384), .ZN(n7358) );
  AND2_X1 U8905 ( .A1(n7475), .A2(n7476), .ZN(n6631) );
  INV_X1 U8906 ( .A(n7605), .ZN(n7642) );
  INV_X2 U8907 ( .A(n7642), .ZN(n7962) );
  AND2_X1 U8908 ( .A1(n12188), .A2(n6680), .ZN(n6632) );
  INV_X1 U8909 ( .A(n10095), .ZN(n7262) );
  XOR2_X1 U8910 ( .A(n12199), .B(n8904), .Z(n6633) );
  OR2_X1 U8911 ( .A1(n13388), .A2(n13089), .ZN(n6634) );
  AND2_X1 U8912 ( .A1(n14609), .A2(n7219), .ZN(n6635) );
  AND2_X1 U8913 ( .A1(n6720), .A2(n6919), .ZN(n6636) );
  INV_X1 U8914 ( .A(n7565), .ZN(n7002) );
  AND2_X1 U8915 ( .A1(n11918), .A2(n14334), .ZN(n6637) );
  OR2_X1 U8916 ( .A1(n14050), .A2(n14038), .ZN(n6638) );
  INV_X1 U8917 ( .A(n9940), .ZN(n7247) );
  AND2_X1 U8918 ( .A1(n10095), .A2(n9516), .ZN(n6639) );
  AND2_X1 U8919 ( .A1(n7364), .A2(n7329), .ZN(n6640) );
  NAND2_X1 U8920 ( .A1(n8632), .A2(n8631), .ZN(n13431) );
  AND2_X1 U8921 ( .A1(n7211), .A2(n7210), .ZN(n6641) );
  INV_X1 U8922 ( .A(n7274), .ZN(n7273) );
  NAND2_X1 U8923 ( .A1(n6699), .A2(n7275), .ZN(n7274) );
  AND2_X1 U8924 ( .A1(n7536), .A2(n6656), .ZN(n6642) );
  AND2_X1 U8925 ( .A1(n9011), .A2(n6631), .ZN(n6643) );
  INV_X1 U8926 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9683) );
  INV_X1 U8927 ( .A(n12090), .ZN(n6916) );
  INV_X1 U8928 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9585) );
  AND2_X1 U8929 ( .A1(n12102), .A2(n12104), .ZN(n6644) );
  NAND2_X1 U8930 ( .A1(n8833), .A2(n8832), .ZN(n13189) );
  AND2_X1 U8931 ( .A1(n6719), .A2(n6922), .ZN(n6645) );
  AND2_X1 U8932 ( .A1(n14812), .A2(n7072), .ZN(n6646) );
  NOR2_X1 U8933 ( .A1(n7534), .A2(n7004), .ZN(n6647) );
  NOR2_X1 U8934 ( .A1(n11727), .A2(n7453), .ZN(n6648) );
  AND2_X1 U8935 ( .A1(n8133), .A2(n6845), .ZN(n6649) );
  AND2_X1 U8936 ( .A1(n9218), .A2(n9219), .ZN(n12730) );
  INV_X1 U8937 ( .A(n12730), .ZN(n7461) );
  INV_X1 U8938 ( .A(n8075), .ZN(n11420) );
  INV_X1 U8939 ( .A(n12681), .ZN(n12711) );
  NAND2_X1 U8940 ( .A1(n8911), .A2(n8910), .ZN(n13377) );
  INV_X1 U8941 ( .A(n11740), .ZN(n6850) );
  INV_X1 U8942 ( .A(n12173), .ZN(n7284) );
  AND2_X1 U8943 ( .A1(n15235), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6650) );
  INV_X1 U8944 ( .A(n9099), .ZN(n7117) );
  INV_X1 U8945 ( .A(n7497), .ZN(n10586) );
  NAND2_X1 U8946 ( .A1(n8293), .A2(n6679), .ZN(n7497) );
  INV_X1 U8947 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13478) );
  OR2_X1 U8948 ( .A1(n13199), .A2(n13189), .ZN(n6651) );
  NAND2_X2 U8950 ( .A1(n8238), .A2(n8239), .ZN(n8545) );
  AND2_X1 U8951 ( .A1(n13812), .A2(n7365), .ZN(n6652) );
  AND2_X1 U8952 ( .A1(n7799), .A2(n7817), .ZN(n6653) );
  AND2_X1 U8953 ( .A1(n8152), .A2(n7463), .ZN(n8121) );
  INV_X1 U8954 ( .A(n14516), .ZN(n7352) );
  OR2_X1 U8955 ( .A1(n11918), .A2(n14334), .ZN(n6654) );
  AND2_X1 U8956 ( .A1(n10876), .A2(n9044), .ZN(n6655) );
  AND4_X1 U8957 ( .A1(n7853), .A2(n7850), .A3(n7555), .A4(n7801), .ZN(n6656)
         );
  AND2_X1 U8958 ( .A1(n6832), .A2(n6831), .ZN(n6657) );
  AND2_X1 U8959 ( .A1(n11212), .A2(n11211), .ZN(n6658) );
  NOR2_X1 U8960 ( .A1(n12107), .A2(n12105), .ZN(n6659) );
  AND2_X1 U8961 ( .A1(n8105), .A2(n9239), .ZN(n6660) );
  NOR2_X1 U8962 ( .A1(n12052), .A2(n12051), .ZN(n6661) );
  OR2_X1 U8963 ( .A1(n13248), .A2(n13092), .ZN(n6662) );
  OR2_X1 U8964 ( .A1(n12631), .A2(n9868), .ZN(n9262) );
  AND2_X1 U8965 ( .A1(n7635), .A2(n7550), .ZN(n7668) );
  AND2_X1 U8966 ( .A1(n7310), .A2(n7308), .ZN(n6663) );
  AND2_X1 U8967 ( .A1(n13896), .A2(n7206), .ZN(n6664) );
  AND2_X1 U8968 ( .A1(n13906), .A2(n7377), .ZN(n6665) );
  AND2_X1 U8969 ( .A1(n8309), .A2(n8199), .ZN(n8358) );
  INV_X1 U8970 ( .A(n11310), .ZN(n7355) );
  XOR2_X1 U8971 ( .A(n14031), .B(n10061), .Z(n10107) );
  INV_X1 U8972 ( .A(n10107), .ZN(n7325) );
  NAND2_X1 U8973 ( .A1(n13913), .A2(n14085), .ZN(n6666) );
  OAI21_X1 U8974 ( .B1(n11693), .B2(n6661), .A(n9001), .ZN(n13348) );
  NAND2_X1 U8975 ( .A1(n11999), .A2(n13109), .ZN(n6667) );
  INV_X1 U8976 ( .A(n7154), .ZN(n7153) );
  OAI21_X1 U8977 ( .B1(n13592), .B2(n12250), .A(n13590), .ZN(n7154) );
  AND2_X1 U8978 ( .A1(n9225), .A2(n7451), .ZN(n6668) );
  AND2_X1 U8979 ( .A1(n9262), .A2(n9257), .ZN(n6669) );
  XNOR2_X1 U8980 ( .A(n10727), .B(n9894), .ZN(n9890) );
  NAND2_X1 U8981 ( .A1(n9442), .A2(n9441), .ZN(n11338) );
  INV_X1 U8982 ( .A(n11338), .ZN(n7219) );
  INV_X2 U8983 ( .A(n12125), .ZN(n12137) );
  NAND2_X1 U8984 ( .A1(n8732), .A2(n8731), .ZN(n13410) );
  AND2_X1 U8985 ( .A1(n9809), .A2(n12721), .ZN(n6670) );
  OR2_X1 U8986 ( .A1(n11999), .A2(n13109), .ZN(n6671) );
  INV_X1 U8987 ( .A(n8375), .ZN(n6936) );
  OR2_X1 U8988 ( .A1(n13913), .A2(n13664), .ZN(n6672) );
  NAND2_X1 U8989 ( .A1(n7457), .A2(n8020), .ZN(n8948) );
  NAND2_X1 U8990 ( .A1(n8710), .A2(n8709), .ZN(n13415) );
  NAND3_X1 U8991 ( .A1(n7635), .A2(n6642), .A3(n6629), .ZN(n6673) );
  INV_X1 U8992 ( .A(n12192), .ZN(n13219) );
  AND2_X1 U8993 ( .A1(n9579), .A2(n9578), .ZN(n13985) );
  INV_X1 U8994 ( .A(n13985), .ZN(n14110) );
  OR2_X1 U8995 ( .A1(n11217), .A2(n11334), .ZN(n6674) );
  INV_X1 U8996 ( .A(n12021), .ZN(n7525) );
  INV_X1 U8997 ( .A(n12093), .ZN(n7524) );
  NAND2_X1 U8998 ( .A1(n6826), .A2(n12504), .ZN(n6675) );
  OR2_X1 U8999 ( .A1(n11430), .A2(n11457), .ZN(n6676) );
  OR2_X1 U9000 ( .A1(n9775), .A2(n15026), .ZN(n6677) );
  INV_X1 U9001 ( .A(n9925), .ZN(n7226) );
  INV_X1 U9002 ( .A(n10098), .ZN(n13947) );
  AND2_X1 U9003 ( .A1(n13388), .A2(n13089), .ZN(n6678) );
  NAND2_X1 U9004 ( .A1(n6974), .A2(n9322), .ZN(n14042) );
  AND3_X1 U9005 ( .A1(n8292), .A2(n8291), .A3(n8294), .ZN(n6679) );
  AND2_X1 U9006 ( .A1(n9603), .A2(n9602), .ZN(n14096) );
  INV_X1 U9007 ( .A(n14096), .ZN(n13946) );
  OR2_X1 U9008 ( .A1(n13419), .A2(n13094), .ZN(n6680) );
  AND2_X1 U9009 ( .A1(n9663), .A2(n9662), .ZN(n13813) );
  INV_X1 U9010 ( .A(n13813), .ZN(n7329) );
  AND2_X1 U9011 ( .A1(n7193), .A2(n12586), .ZN(n6681) );
  INV_X1 U9012 ( .A(n7487), .ZN(n7486) );
  NOR2_X1 U9013 ( .A1(n13217), .A2(n13090), .ZN(n7487) );
  NOR2_X1 U9014 ( .A1(n13386), .A2(n6777), .ZN(n6682) );
  INV_X1 U9015 ( .A(n6984), .ZN(n6983) );
  INV_X1 U9016 ( .A(n11998), .ZN(n6923) );
  INV_X1 U9017 ( .A(n7336), .ZN(n7335) );
  NOR2_X1 U9018 ( .A1(n14050), .A2(n13859), .ZN(n7336) );
  AND2_X1 U9019 ( .A1(n9991), .A2(n9992), .ZN(n6683) );
  INV_X1 U9020 ( .A(n9781), .ZN(n7161) );
  INV_X1 U9021 ( .A(n10021), .ZN(n7231) );
  AND2_X1 U9022 ( .A1(n9962), .A2(n9753), .ZN(n6684) );
  INV_X1 U9023 ( .A(n7167), .ZN(n7166) );
  NAND2_X1 U9024 ( .A1(n12461), .A2(n7168), .ZN(n7167) );
  INV_X1 U9025 ( .A(n7467), .ZN(n7466) );
  OAI21_X1 U9026 ( .B1(n7469), .B2(n7468), .A(n6662), .ZN(n7467) );
  AND2_X1 U9027 ( .A1(n8641), .A2(n8623), .ZN(n6685) );
  AND2_X1 U9028 ( .A1(n13189), .A2(n13088), .ZN(n6686) );
  NAND2_X1 U9029 ( .A1(n12533), .A2(n12527), .ZN(n6687) );
  AND2_X1 U9030 ( .A1(n9651), .A2(n9650), .ZN(n6688) );
  AND2_X1 U9031 ( .A1(n7461), .A2(n7901), .ZN(n6689) );
  OR2_X1 U9032 ( .A1(n9954), .A2(n9957), .ZN(n6690) );
  AND2_X1 U9033 ( .A1(n12896), .A2(n12722), .ZN(n6691) );
  AND2_X1 U9034 ( .A1(n12109), .A2(n12108), .ZN(n6692) );
  INV_X1 U9035 ( .A(n6898), .ZN(n6896) );
  NAND2_X1 U9036 ( .A1(n14057), .A2(n13873), .ZN(n6898) );
  NAND2_X1 U9037 ( .A1(n13924), .A2(n7343), .ZN(n7345) );
  NOR2_X1 U9038 ( .A1(n7524), .A2(n12092), .ZN(n6693) );
  NOR2_X1 U9039 ( .A1(n14383), .A2(n14288), .ZN(n6694) );
  INV_X1 U9040 ( .A(n7572), .ZN(n7311) );
  NOR2_X1 U9041 ( .A1(n12312), .A2(n12311), .ZN(n6695) );
  NOR2_X1 U9042 ( .A1(n9808), .A2(n12758), .ZN(n6696) );
  INV_X1 U9043 ( .A(n8999), .ZN(n6804) );
  INV_X1 U9044 ( .A(n7208), .ZN(n7207) );
  NAND2_X1 U9045 ( .A1(n13885), .A2(n7209), .ZN(n7208) );
  AND2_X1 U9046 ( .A1(n14594), .A2(n10958), .ZN(n6697) );
  AND2_X1 U9047 ( .A1(n9769), .A2(n9770), .ZN(n6698) );
  OR2_X1 U9048 ( .A1(n10075), .A2(n10074), .ZN(n6699) );
  INV_X1 U9049 ( .A(n12018), .ZN(n6920) );
  NOR2_X1 U9050 ( .A1(n14034), .A2(n13663), .ZN(n6700) );
  NAND2_X1 U9051 ( .A1(n7248), .A2(n7245), .ZN(n6701) );
  NAND2_X1 U9052 ( .A1(n7241), .A2(n7238), .ZN(n6702) );
  AND2_X1 U9053 ( .A1(n8578), .A2(n15227), .ZN(n6704) );
  INV_X1 U9054 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8233) );
  NAND2_X1 U9055 ( .A1(n9169), .A2(n9168), .ZN(n11710) );
  INV_X1 U9056 ( .A(n11710), .ZN(n7014) );
  AND2_X1 U9057 ( .A1(n12020), .A2(n7525), .ZN(n6705) );
  AND2_X1 U9058 ( .A1(n8516), .A2(n10169), .ZN(n6706) );
  AND2_X1 U9059 ( .A1(n7000), .A2(SI_0_), .ZN(n6707) );
  AND2_X1 U9060 ( .A1(n12084), .A2(n12083), .ZN(n6708) );
  INV_X1 U9061 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10173) );
  INV_X1 U9062 ( .A(n12224), .ZN(n7137) );
  AND2_X1 U9063 ( .A1(n12223), .A2(n12222), .ZN(n12224) );
  INV_X1 U9064 ( .A(n7095), .ZN(n7094) );
  NAND2_X1 U9065 ( .A1(n7099), .A2(n7774), .ZN(n7095) );
  INV_X1 U9066 ( .A(n7142), .ZN(n7141) );
  NAND2_X1 U9067 ( .A1(n7145), .A2(n7143), .ZN(n7142) );
  AND2_X1 U9068 ( .A1(n9934), .A2(n9933), .ZN(n6709) );
  NAND2_X1 U9069 ( .A1(n10108), .A2(n10076), .ZN(n6710) );
  NAND2_X1 U9070 ( .A1(n10082), .A2(n10080), .ZN(n6711) );
  AND2_X1 U9071 ( .A1(n7738), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n6712) );
  AND2_X1 U9072 ( .A1(n6858), .A2(n6654), .ZN(n6713) );
  AND2_X1 U9073 ( .A1(n13404), .A2(n13092), .ZN(n6714) );
  AND2_X1 U9074 ( .A1(n12447), .A2(n12681), .ZN(n6715) );
  OR2_X1 U9075 ( .A1(n6799), .A2(n8999), .ZN(n6716) );
  OR2_X1 U9076 ( .A1(n7328), .A2(n7325), .ZN(n6717) );
  AND2_X1 U9077 ( .A1(n7329), .A2(n7363), .ZN(n6718) );
  INV_X1 U9078 ( .A(n11872), .ZN(n7136) );
  OR2_X1 U9079 ( .A1(n12002), .A2(n12000), .ZN(n6719) );
  OR2_X1 U9080 ( .A1(n7525), .A2(n12020), .ZN(n6720) );
  AND2_X1 U9081 ( .A1(n8681), .A2(n8682), .ZN(n6721) );
  AND2_X1 U9082 ( .A1(n7328), .A2(n7325), .ZN(n6722) );
  NAND2_X1 U9083 ( .A1(n8604), .A2(n8601), .ZN(n6723) );
  INV_X1 U9084 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8127) );
  INV_X1 U9085 ( .A(n9011), .ZN(n7468) );
  OR2_X1 U9086 ( .A1(n13404), .A2(n13019), .ZN(n9011) );
  OR2_X1 U9087 ( .A1(n9073), .A2(n6678), .ZN(n6724) );
  INV_X1 U9088 ( .A(n12059), .ZN(n6907) );
  AND2_X1 U9089 ( .A1(n6855), .A2(n6654), .ZN(n6725) );
  AND2_X1 U9090 ( .A1(n7326), .A2(n7325), .ZN(n6726) );
  OR2_X1 U9091 ( .A1(n7326), .A2(n7325), .ZN(n6727) );
  AND2_X1 U9092 ( .A1(n12692), .A2(n9239), .ZN(n6728) );
  INV_X1 U9093 ( .A(n10105), .ZN(n13837) );
  XNOR2_X1 U9094 ( .A(n14042), .B(n13845), .ZN(n10105) );
  INV_X1 U9095 ( .A(n9178), .ZN(n7033) );
  INV_X1 U9096 ( .A(n6818), .ZN(n6817) );
  OAI21_X1 U9097 ( .B1(n7477), .B2(n6819), .A(n7484), .ZN(n6818) );
  INV_X1 U9098 ( .A(n9060), .ZN(n7306) );
  INV_X1 U9099 ( .A(n8473), .ZN(n7384) );
  AND2_X1 U9100 ( .A1(n8020), .A2(n8036), .ZN(n6729) );
  AND2_X1 U9101 ( .A1(n8192), .A2(n7379), .ZN(n6730) );
  AND2_X1 U9102 ( .A1(n13947), .A2(n9987), .ZN(n6731) );
  AND2_X1 U9103 ( .A1(n7047), .A2(n7048), .ZN(n6732) );
  AND2_X1 U9104 ( .A1(n6833), .A2(n9781), .ZN(n6733) );
  NAND2_X1 U9105 ( .A1(n11217), .A2(n11334), .ZN(n6734) );
  OR2_X1 U9106 ( .A1(n10000), .A2(n9998), .ZN(n6735) );
  OR2_X1 U9107 ( .A1(n9945), .A2(n9943), .ZN(n6736) );
  OR2_X1 U9108 ( .A1(n12014), .A2(n12012), .ZN(n6737) );
  OR2_X1 U9109 ( .A1(n12034), .A2(n12032), .ZN(n6738) );
  OR2_X1 U9110 ( .A1(n10011), .A2(n10009), .ZN(n6739) );
  OR2_X1 U9111 ( .A1(n10020), .A2(n7231), .ZN(n6740) );
  AND2_X1 U9112 ( .A1(n7355), .A2(n9748), .ZN(n6741) );
  INV_X1 U9113 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9319) );
  INV_X1 U9114 ( .A(n9073), .ZN(n7296) );
  INV_X1 U9115 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7282) );
  NAND2_X1 U9116 ( .A1(n9189), .A2(n8099), .ZN(n7006) );
  AND2_X1 U9117 ( .A1(n7281), .A2(n9585), .ZN(n6742) );
  INV_X1 U9118 ( .A(n13108), .ZN(n6810) );
  INV_X1 U9119 ( .A(n11528), .ZN(n11521) );
  NAND2_X1 U9120 ( .A1(n6861), .A2(n7176), .ZN(n12386) );
  NAND2_X1 U9121 ( .A1(n11881), .A2(n9790), .ZN(n12363) );
  AND2_X1 U9122 ( .A1(n14000), .A2(n7213), .ZN(n6743) );
  OR2_X1 U9123 ( .A1(n7851), .A2(n7185), .ZN(n6744) );
  INV_X1 U9124 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7103) );
  NAND2_X1 U9125 ( .A1(n13009), .A2(n8623), .ZN(n13058) );
  NAND2_X1 U9126 ( .A1(n6840), .A2(n6839), .ZN(n12434) );
  NAND2_X1 U9127 ( .A1(n6841), .A2(n7164), .ZN(n12369) );
  NAND2_X1 U9128 ( .A1(n7165), .A2(n9807), .ZN(n12460) );
  XNOR2_X1 U9129 ( .A(n14821), .B(n6810), .ZN(n11000) );
  INV_X1 U9130 ( .A(n11000), .ZN(n8988) );
  NAND2_X1 U9131 ( .A1(n9345), .A2(n9344), .ZN(n14057) );
  INV_X1 U9132 ( .A(n14057), .ZN(n7209) );
  INV_X1 U9133 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7043) );
  OR2_X1 U9134 ( .A1(n13385), .A2(n14826), .ZN(n6745) );
  NAND2_X1 U9135 ( .A1(n7172), .A2(n9812), .ZN(n12376) );
  INV_X1 U9136 ( .A(n9995), .ZN(n7240) );
  AND2_X1 U9137 ( .A1(n13415), .A2(n13093), .ZN(n6746) );
  AND4_X1 U9138 ( .A1(n8391), .A2(n8390), .A3(n8389), .A4(n8388), .ZN(n10829)
         );
  NAND2_X1 U9139 ( .A1(n7223), .A2(n9534), .ZN(n9547) );
  INV_X1 U9140 ( .A(n9012), .ZN(n13088) );
  INV_X1 U9141 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8064) );
  INV_X1 U9142 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7555) );
  INV_X1 U9143 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7889) );
  OR2_X1 U9144 ( .A1(n12278), .A2(n12277), .ZN(n6747) );
  OR2_X1 U9145 ( .A1(n7851), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n6748) );
  NOR2_X1 U9146 ( .A1(n12779), .A2(n10685), .ZN(n6749) );
  AND2_X1 U9147 ( .A1(n12745), .A2(n7901), .ZN(n6750) );
  AND2_X1 U9148 ( .A1(n10808), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n6751) );
  AND2_X1 U9149 ( .A1(n12953), .A2(n12952), .ZN(n6752) );
  OR2_X1 U9150 ( .A1(n7851), .A2(n7186), .ZN(n6753) );
  INV_X1 U9151 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7850) );
  INV_X1 U9152 ( .A(n8285), .ZN(n8457) );
  INV_X1 U9153 ( .A(n12533), .ZN(n6955) );
  XNOR2_X1 U9154 ( .A(n9711), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9879) );
  INV_X1 U9155 ( .A(n9607), .ZN(n9617) );
  AND2_X1 U9156 ( .A1(n11275), .A2(n6675), .ZN(n7174) );
  INV_X1 U9157 ( .A(n7071), .ZN(n10881) );
  INV_X1 U9158 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11285) );
  XNOR2_X1 U9159 ( .A(n11379), .B(n11401), .ZN(n14920) );
  OAI21_X1 U9160 ( .B1(n11762), .B2(n6858), .A(n6855), .ZN(n11917) );
  OAI21_X1 U9161 ( .B1(n10718), .B2(n10715), .A(n9740), .ZN(n14530) );
  NAND2_X1 U9162 ( .A1(n7320), .A2(n7322), .ZN(n14501) );
  AOI21_X1 U9163 ( .B1(n6774), .B2(n11213), .A(n6658), .ZN(n11324) );
  NAND2_X1 U9164 ( .A1(n6854), .A2(n6853), .ZN(n11927) );
  NAND2_X1 U9165 ( .A1(n9616), .A2(n9615), .ZN(n14088) );
  INV_X1 U9166 ( .A(n14088), .ZN(n7210) );
  AOI21_X1 U9167 ( .B1(n8131), .B2(P3_IR_REG_26__SCAN_IN), .A(n8130), .ZN(
        n8132) );
  NAND2_X1 U9168 ( .A1(n6836), .A2(n7159), .ZN(n11684) );
  NOR2_X1 U9169 ( .A1(n14919), .A2(n11380), .ZN(n6754) );
  AND2_X1 U9170 ( .A1(n7144), .A2(n7141), .ZN(n6755) );
  NOR2_X1 U9171 ( .A1(n9312), .A2(n9311), .ZN(n9534) );
  INV_X1 U9172 ( .A(SI_20_), .ZN(n10873) );
  INV_X1 U9173 ( .A(n12600), .ZN(n6962) );
  INV_X1 U9174 ( .A(n7946), .ZN(n7078) );
  INV_X1 U9175 ( .A(n11180), .ZN(n7323) );
  OR2_X1 U9176 ( .A1(n14665), .A2(n7214), .ZN(n6756) );
  INV_X1 U9177 ( .A(n14821), .ZN(n7072) );
  NAND2_X1 U9178 ( .A1(n8411), .A2(n8410), .ZN(n12015) );
  INV_X1 U9179 ( .A(n12015), .ZN(n7070) );
  NAND2_X1 U9180 ( .A1(n10846), .A2(n6770), .ZN(n10987) );
  INV_X1 U9181 ( .A(n10987), .ZN(n7068) );
  AND2_X1 U9182 ( .A1(n7985), .A2(n14161), .ZN(n6757) );
  NAND2_X1 U9183 ( .A1(n14157), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6758) );
  INV_X1 U9184 ( .A(n9764), .ZN(n6845) );
  AND2_X1 U9185 ( .A1(n8152), .A2(n7040), .ZN(n12927) );
  INV_X1 U9186 ( .A(n7120), .ZN(n7118) );
  NAND2_X1 U9187 ( .A1(n14144), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7120) );
  AND2_X1 U9188 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n9100), .ZN(n6759) );
  INV_X1 U9189 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6767) );
  INV_X1 U9190 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6771) );
  INV_X1 U9191 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6999) );
  INV_X1 U9192 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7049) );
  INV_X1 U9193 ( .A(n7001), .ZN(n14141) );
  NAND2_X1 U9194 ( .A1(n12976), .A2(n12975), .ZN(n12974) );
  NAND2_X1 U9195 ( .A1(n11286), .A2(n11288), .ZN(n7402) );
  NAND2_X1 U9196 ( .A1(n11194), .A2(n8490), .ZN(n11249) );
  OAI21_X1 U9197 ( .B1(n8472), .B2(n7384), .A(n11195), .ZN(n7383) );
  INV_X1 U9198 ( .A(n7383), .ZN(n7382) );
  INV_X1 U9199 ( .A(n7188), .ZN(n11375) );
  NOR2_X1 U9200 ( .A1(n11585), .A2(n15398), .ZN(n11839) );
  NAND2_X1 U9201 ( .A1(n10772), .A2(n10771), .ZN(n11374) );
  NOR2_X1 U9202 ( .A1(n14954), .A2(n11382), .ZN(n14974) );
  NOR2_X1 U9203 ( .A1(n11383), .A2(n11384), .ZN(n11515) );
  NAND2_X1 U9204 ( .A1(n6963), .A2(n6779), .ZN(P3_U3201) );
  OAI21_X1 U9205 ( .B1(n12610), .B2(n14994), .A(n6781), .ZN(n6780) );
  NAND2_X1 U9206 ( .A1(n7454), .A2(n6648), .ZN(n11726) );
  NOR2_X2 U9207 ( .A1(n8964), .A2(n12336), .ZN(n8967) );
  INV_X2 U9208 ( .A(n6761), .ZN(n12679) );
  NAND2_X1 U9209 ( .A1(n13553), .A2(n10611), .ZN(n10947) );
  NAND2_X1 U9210 ( .A1(n12266), .A2(n12265), .ZN(n13545) );
  NAND2_X1 U9211 ( .A1(n7691), .A2(n7455), .ZN(n7454) );
  XNOR2_X1 U9212 ( .A(n7570), .B(n7569), .ZN(n8074) );
  AOI22_X2 U9213 ( .A1(n13653), .A2(n13652), .B1(n12240), .B2(n12239), .ZN(
        n13580) );
  INV_X1 U9214 ( .A(n6935), .ZN(n6934) );
  NAND2_X1 U9215 ( .A1(n8724), .A2(n8723), .ZN(n8726) );
  NAND3_X1 U9216 ( .A1(n7313), .A2(n11967), .A3(n9083), .ZN(n9094) );
  NAND2_X1 U9217 ( .A1(n6766), .A2(n6752), .ZN(P2_U3186) );
  NAND2_X1 U9218 ( .A1(n12954), .A2(n12947), .ZN(n6766) );
  AOI21_X2 U9219 ( .B1(n10409), .B2(n10408), .A(n8298), .ZN(n13026) );
  INV_X1 U9220 ( .A(n8246), .ZN(n6769) );
  XNOR2_X2 U9221 ( .A(n8234), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8238) );
  NAND2_X4 U9222 ( .A1(n12214), .A2(n8917), .ZN(n8433) );
  AND2_X4 U9223 ( .A1(n8433), .A2(n10067), .ZN(n8285) );
  NAND2_X2 U9224 ( .A1(n8256), .A2(n6663), .ZN(n14791) );
  AND2_X2 U9225 ( .A1(n13114), .A2(n11972), .ZN(n8273) );
  NAND2_X1 U9226 ( .A1(n7288), .A2(n7287), .ZN(n13170) );
  NAND2_X1 U9227 ( .A1(n9047), .A2(n9046), .ZN(n11127) );
  NAND2_X1 U9228 ( .A1(n10877), .A2(n12172), .ZN(n10876) );
  NAND2_X1 U9229 ( .A1(n10929), .A2(n9045), .ZN(n11090) );
  NAND2_X1 U9230 ( .A1(n6655), .A2(n7284), .ZN(n10929) );
  NAND2_X1 U9231 ( .A1(n13218), .A2(n9074), .ZN(n7295) );
  NAND2_X1 U9232 ( .A1(n7314), .A2(n7315), .ZN(n10995) );
  XNOR2_X1 U9233 ( .A(n13111), .B(n6770), .ZN(n10845) );
  NAND2_X2 U9234 ( .A1(n8336), .A2(n8335), .ZN(n11999) );
  OR2_X1 U9235 ( .A1(n10176), .A2(n10431), .ZN(n7202) );
  AOI22_X1 U9236 ( .A1(n13509), .A2(n13510), .B1(n12319), .B2(n12318), .ZN(
        n12328) );
  OAI22_X1 U9237 ( .A1(n10703), .A2(n10348), .B1(n9363), .B2(n12284), .ZN(
        n10604) );
  AND2_X2 U9238 ( .A1(n10378), .A2(n8276), .ZN(n10409) );
  NAND2_X1 U9239 ( .A1(n10380), .A2(n10379), .ZN(n10378) );
  NAND2_X1 U9240 ( .A1(n13026), .A2(n13028), .ZN(n13027) );
  INV_X4 U9241 ( .A(n8433), .ZN(n10181) );
  NAND2_X1 U9242 ( .A1(n7381), .A2(n7382), .ZN(n11194) );
  OAI22_X1 U9243 ( .A1(n10828), .A2(n7407), .B1(n10826), .B2(n7406), .ZN(
        n11019) );
  NAND2_X1 U9244 ( .A1(n10331), .A2(n10332), .ZN(n10330) );
  NAND2_X1 U9245 ( .A1(n7402), .A2(n6778), .ZN(n11576) );
  NAND2_X1 U9246 ( .A1(n6624), .A2(n8192), .ZN(n7380) );
  AND2_X4 U9247 ( .A1(n10502), .A2(n11208), .ZN(n13359) );
  NAND2_X1 U9248 ( .A1(n11175), .A2(n11174), .ZN(n11214) );
  OAI21_X2 U9249 ( .B1(n13580), .B2(n7154), .A(n7151), .ZN(n13631) );
  AND2_X1 U9250 ( .A1(n14217), .A2(n14218), .ZN(n15523) );
  NAND3_X1 U9251 ( .A1(n7047), .A2(n7046), .A3(n7048), .ZN(n7044) );
  NOR2_X1 U9252 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n14457), .ZN(n14262) );
  NOR2_X2 U9253 ( .A1(n14225), .A2(n14226), .ZN(n14227) );
  NAND2_X1 U9254 ( .A1(n15515), .A2(n15516), .ZN(n14220) );
  OR2_X1 U9255 ( .A1(n14450), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7065) );
  NAND2_X1 U9256 ( .A1(n15520), .A2(n15521), .ZN(n14233) );
  AOI21_X1 U9257 ( .B1(n14277), .B2(n14215), .A(n14274), .ZN(n14217) );
  NOR2_X1 U9258 ( .A1(n14255), .A2(n14254), .ZN(n14450) );
  NAND2_X1 U9259 ( .A1(n13552), .A2(n13554), .ZN(n13553) );
  XNOR2_X1 U9260 ( .A(n10609), .B(n10608), .ZN(n13552) );
  NAND2_X1 U9261 ( .A1(n9676), .A2(n9683), .ZN(n7347) );
  NAND2_X1 U9262 ( .A1(n7410), .A2(n8493), .ZN(n8515) );
  NOR2_X2 U9263 ( .A1(n13156), .A2(n13161), .ZN(n13157) );
  NAND2_X1 U9264 ( .A1(n13299), .A2(n13294), .ZN(n13289) );
  NAND2_X1 U9265 ( .A1(n6934), .A2(n6936), .ZN(n6932) );
  NOR2_X2 U9266 ( .A1(n13258), .A2(n13404), .ZN(n13246) );
  OAI21_X1 U9267 ( .B1(n8355), .B2(n6936), .A(n8380), .ZN(n6935) );
  AND2_X1 U9268 ( .A1(n8325), .A2(n8303), .ZN(n8304) );
  NAND2_X1 U9269 ( .A1(n9601), .A2(n9600), .ZN(n13948) );
  INV_X1 U9270 ( .A(n7368), .ZN(n13835) );
  OAI21_X1 U9271 ( .B1(n8283), .B2(n6789), .A(n6788), .ZN(n8326) );
  NAND2_X1 U9272 ( .A1(n8326), .A2(n8325), .ZN(n8331) );
  NAND3_X1 U9273 ( .A1(n7349), .A2(n10900), .A3(n7348), .ZN(n9424) );
  AND2_X4 U9274 ( .A1(n12313), .A2(n10341), .ZN(n12321) );
  AOI22_X1 U9275 ( .A1(n10947), .A2(n10946), .B1(n10945), .B2(n10944), .ZN(
        n13537) );
  NOR2_X1 U9276 ( .A1(n10956), .A2(n10957), .ZN(n11033) );
  NAND3_X1 U9277 ( .A1(n8185), .A2(n8184), .A3(n6775), .ZN(n8202) );
  NAND2_X2 U9278 ( .A1(n12984), .A2(n6941), .ZN(n13071) );
  NAND4_X1 U9279 ( .A1(n8191), .A2(n8189), .A3(n8190), .A4(n8204), .ZN(n8213)
         );
  NAND2_X1 U9280 ( .A1(n9070), .A2(n9069), .ZN(n13239) );
  NAND2_X1 U9281 ( .A1(n7298), .A2(n7297), .ZN(n13253) );
  NAND2_X1 U9282 ( .A1(n7289), .A2(n7293), .ZN(n13185) );
  NOR2_X1 U9283 ( .A1(n8201), .A2(n8182), .ZN(n8191) );
  NAND2_X2 U9284 ( .A1(n12986), .A2(n12985), .ZN(n12984) );
  NAND2_X2 U9285 ( .A1(n13016), .A2(n8786), .ZN(n12986) );
  NAND2_X1 U9286 ( .A1(n13071), .A2(n8826), .ZN(n12949) );
  XNOR2_X2 U9287 ( .A(n12238), .B(n12239), .ZN(n13653) );
  NAND2_X1 U9288 ( .A1(n13537), .A2(n13536), .ZN(n13535) );
  NAND2_X1 U9289 ( .A1(n13613), .A2(n13612), .ZN(n13611) );
  OAI21_X2 U9290 ( .B1(n11214), .B2(n7142), .A(n7138), .ZN(n11604) );
  NOR2_X4 U9291 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7158) );
  NAND2_X1 U9292 ( .A1(n12598), .A2(n6962), .ZN(n6783) );
  INV_X1 U9293 ( .A(n12597), .ZN(n6784) );
  INV_X1 U9294 ( .A(n6787), .ZN(n6788) );
  OAI21_X1 U9295 ( .B1(n8282), .B2(n6789), .A(n8304), .ZN(n6787) );
  NAND4_X1 U9296 ( .A1(n6790), .A2(P2_DATAO_REG_1__SCAN_IN), .A3(n6887), .A4(
        n15343), .ZN(n6791) );
  NAND2_X2 U9297 ( .A1(n6793), .A2(n6794), .ZN(n8226) );
  NAND3_X1 U9298 ( .A1(n6793), .A2(n6794), .A3(P1_DATAO_REG_1__SCAN_IN), .ZN(
        n6792) );
  NAND2_X1 U9299 ( .A1(n6795), .A2(n11502), .ZN(n6796) );
  NAND2_X2 U9300 ( .A1(n6811), .A2(n8361), .ZN(n14821) );
  INV_X1 U9301 ( .A(n7465), .ZN(n6815) );
  NOR2_X1 U9302 ( .A1(n7465), .A2(n6825), .ZN(n6816) );
  OAI21_X1 U9303 ( .B1(n6818), .B2(n6815), .A(n6813), .ZN(n7480) );
  NAND2_X1 U9304 ( .A1(n7465), .A2(n7466), .ZN(n13223) );
  NAND2_X1 U9305 ( .A1(n13230), .A2(n7467), .ZN(n6824) );
  XNOR2_X1 U9306 ( .A(n6826), .B(n12504), .ZN(n11240) );
  AND2_X2 U9307 ( .A1(n7549), .A2(n7548), .ZN(n6827) );
  INV_X2 U9308 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7548) );
  NAND2_X1 U9309 ( .A1(n9836), .A2(n12399), .ZN(n12401) );
  NAND2_X1 U9310 ( .A1(n12401), .A2(n9837), .ZN(n12470) );
  NAND2_X1 U9311 ( .A1(n7174), .A2(n11239), .ZN(n6838) );
  NAND2_X1 U9312 ( .A1(n6835), .A2(n6733), .ZN(n6836) );
  NAND2_X1 U9313 ( .A1(n6838), .A2(n6837), .ZN(n11343) );
  NAND2_X1 U9314 ( .A1(n12416), .A2(n6842), .ZN(n6840) );
  NAND3_X1 U9315 ( .A1(n6846), .A2(n6848), .A3(n8133), .ZN(n11939) );
  NAND3_X1 U9316 ( .A1(n6846), .A2(n6848), .A3(n6649), .ZN(n9767) );
  NAND2_X1 U9317 ( .A1(n6725), .A2(n11762), .ZN(n6854) );
  AND2_X1 U9318 ( .A1(n7176), .A2(n6860), .ZN(n6859) );
  INV_X1 U9319 ( .A(n6864), .ZN(n8118) );
  AND2_X1 U9320 ( .A1(n6872), .A2(n6873), .ZN(n14864) );
  NAND2_X1 U9321 ( .A1(n11377), .A2(n14861), .ZN(n6873) );
  NAND2_X1 U9322 ( .A1(n14377), .A2(n6878), .ZN(n6877) );
  NAND2_X1 U9323 ( .A1(n7319), .A2(n6885), .ZN(n11109) );
  NAND2_X1 U9324 ( .A1(n8226), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6886) );
  INV_X1 U9325 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n6890) );
  OR2_X1 U9326 ( .A1(n13858), .A2(n6895), .ZN(n6891) );
  NAND2_X1 U9327 ( .A1(n6891), .A2(n6892), .ZN(n6897) );
  NAND2_X1 U9328 ( .A1(n13953), .A2(n6731), .ZN(n13938) );
  INV_X1 U9329 ( .A(n12078), .ZN(n12075) );
  NAND3_X1 U9330 ( .A1(n12074), .A2(n6906), .A3(n6905), .ZN(n6903) );
  NAND2_X1 U9331 ( .A1(n6908), .A2(n6909), .ZN(n7515) );
  NAND3_X1 U9332 ( .A1(n12101), .A2(n6910), .A3(n12100), .ZN(n6908) );
  NOR2_X1 U9333 ( .A1(n6659), .A2(n6644), .ZN(n6909) );
  INV_X1 U9334 ( .A(n12102), .ZN(n6911) );
  NAND2_X1 U9335 ( .A1(n12089), .A2(n6913), .ZN(n6912) );
  OAI21_X1 U9336 ( .B1(n6912), .B2(n6708), .A(n6914), .ZN(n7522) );
  NAND2_X1 U9337 ( .A1(n12017), .A2(n6636), .ZN(n6918) );
  OAI21_X1 U9338 ( .B1(n11997), .B2(n6924), .A(n6645), .ZN(n6926) );
  INV_X4 U9339 ( .A(n11978), .ZN(n12155) );
  NAND3_X1 U9340 ( .A1(n12201), .A2(n12161), .A3(n12131), .ZN(n11978) );
  MUX2_X1 U9341 ( .A(n13111), .B(n11983), .S(n11978), .Z(n11984) );
  OAI211_X2 U9342 ( .C1(n12125), .C2(n10127), .A(n6928), .B(n6927), .ZN(n11983) );
  INV_X1 U9343 ( .A(n12115), .ZN(n6931) );
  OAI21_X1 U9344 ( .B1(n8356), .B2(n6936), .A(n6934), .ZN(n8398) );
  NAND3_X1 U9345 ( .A1(n6933), .A2(n8397), .A3(n6932), .ZN(n8403) );
  NAND2_X1 U9346 ( .A1(n8356), .A2(n6934), .ZN(n6933) );
  NAND2_X2 U9347 ( .A1(n13010), .A2(n13011), .ZN(n13009) );
  NAND2_X1 U9348 ( .A1(n8449), .A2(n6946), .ZN(n6943) );
  NAND2_X1 U9349 ( .A1(n6943), .A2(n6944), .ZN(n8532) );
  NAND2_X1 U9350 ( .A1(n8449), .A2(n8448), .ZN(n8454) );
  OAI21_X4 U9351 ( .B1(n10807), .B2(n12125), .A(n8541), .ZN(n13452) );
  NAND3_X1 U9352 ( .A1(n7324), .A2(n6971), .A3(n6727), .ZN(n6970) );
  XNOR2_X2 U9353 ( .A(n9672), .B(n7325), .ZN(n14030) );
  NAND2_X1 U9354 ( .A1(n8576), .A2(n6979), .ZN(n6977) );
  NAND2_X1 U9355 ( .A1(n8574), .A2(n8573), .ZN(n6984) );
  NAND2_X1 U9356 ( .A1(n8680), .A2(n6986), .ZN(n6985) );
  NAND2_X1 U9357 ( .A1(n6985), .A2(n6988), .ZN(n8707) );
  NAND4_X1 U9358 ( .A1(n7433), .A2(n8787), .A3(n6997), .A4(n7430), .ZN(n6991)
         );
  NAND2_X1 U9359 ( .A1(n6992), .A2(n7433), .ZN(n6994) );
  NAND2_X1 U9360 ( .A1(n7433), .A2(n8787), .ZN(n8811) );
  NAND2_X1 U9361 ( .A1(n7572), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6998) );
  OAI21_X1 U9362 ( .B1(n7572), .B2(n6999), .A(n6998), .ZN(n8301) );
  NAND2_X2 U9363 ( .A1(n7000), .A2(P1_U3086), .ZN(n7001) );
  NAND2_X2 U9364 ( .A1(n7311), .A2(P1_U3086), .ZN(n14160) );
  MUX2_X1 U9365 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n7000), .Z(n8703) );
  MUX2_X1 U9366 ( .A(n11202), .B(n7920), .S(n7000), .Z(n8683) );
  MUX2_X1 U9367 ( .A(n10398), .B(n15235), .S(n7000), .Z(n8729) );
  MUX2_X1 U9368 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n7000), .Z(n8762) );
  MUX2_X1 U9369 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n7000), .Z(n8807) );
  MUX2_X1 U9370 ( .A(n14154), .B(n13499), .S(n7000), .Z(n8827) );
  MUX2_X1 U9371 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n7000), .Z(n8908) );
  MUX2_X1 U9372 ( .A(n14148), .B(n13490), .S(n7000), .Z(n9018) );
  MUX2_X1 U9373 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7000), .Z(n10042) );
  MUX2_X1 U9374 ( .A(n14144), .B(n13487), .S(n7000), .Z(n10040) );
  OAI21_X1 U9375 ( .B1(n12810), .B2(n7006), .A(n6647), .ZN(n7003) );
  NAND2_X1 U9376 ( .A1(n7015), .A2(n7016), .ZN(n9124) );
  NAND2_X1 U9377 ( .A1(n8947), .A2(n7019), .ZN(n7015) );
  NAND2_X1 U9378 ( .A1(n8947), .A2(n6669), .ZN(n7018) );
  NAND2_X1 U9379 ( .A1(n8947), .A2(n9257), .ZN(n8962) );
  NAND2_X1 U9380 ( .A1(n7546), .A2(n7027), .ZN(n7025) );
  NAND2_X1 U9381 ( .A1(n7025), .A2(n7026), .ZN(n12695) );
  NAND2_X1 U9382 ( .A1(n8095), .A2(n11808), .ZN(n7035) );
  NAND2_X1 U9383 ( .A1(n7030), .A2(n7031), .ZN(n8097) );
  NAND3_X1 U9384 ( .A1(n8095), .A2(n11808), .A3(n9178), .ZN(n7030) );
  OAI21_X1 U9385 ( .B1(n12692), .B2(n7038), .A(n7036), .ZN(n8106) );
  NAND2_X1 U9386 ( .A1(n12742), .A2(n7039), .ZN(n8101) );
  NAND3_X1 U9387 ( .A1(n7047), .A2(n14317), .A3(n7048), .ZN(n14316) );
  INV_X1 U9388 ( .A(n14460), .ZN(n7047) );
  NAND2_X1 U9389 ( .A1(n7060), .A2(n7063), .ZN(n14260) );
  NAND2_X1 U9390 ( .A1(n7065), .A2(n7061), .ZN(n7060) );
  NOR2_X1 U9391 ( .A1(n14451), .A2(n7062), .ZN(n7061) );
  OAI211_X2 U9392 ( .C1(n8457), .C2(n7629), .A(n7067), .B(n7066), .ZN(n11987)
         );
  NAND2_X1 U9393 ( .A1(n6646), .A2(n10973), .ZN(n7071) );
  NOR2_X2 U9394 ( .A1(n6651), .A2(n13377), .ZN(n13177) );
  NOR2_X2 U9395 ( .A1(n13226), .A2(n13393), .ZN(n13213) );
  NOR2_X2 U9396 ( .A1(n13320), .A2(n13425), .ZN(n13299) );
  NAND2_X1 U9397 ( .A1(n9080), .A2(n11640), .ZN(n13358) );
  NAND2_X1 U9398 ( .A1(n7507), .A2(n6624), .ZN(n8216) );
  INV_X1 U9399 ( .A(n7083), .ZN(n7970) );
  NAND2_X1 U9400 ( .A1(n7721), .A2(n7088), .ZN(n7085) );
  NAND2_X1 U9401 ( .A1(n7085), .A2(n7086), .ZN(n7753) );
  NAND2_X1 U9402 ( .A1(n7102), .A2(n7101), .ZN(n7828) );
  NAND2_X1 U9403 ( .A1(n7104), .A2(n7108), .ZN(n7886) );
  NAND2_X1 U9404 ( .A1(n7848), .A2(n7105), .ZN(n7104) );
  NAND2_X1 U9405 ( .A1(n7982), .A2(n14161), .ZN(n7111) );
  NAND2_X1 U9406 ( .A1(n7111), .A2(n7984), .ZN(n8000) );
  NAND2_X1 U9407 ( .A1(n7114), .A2(n7115), .ZN(n9104) );
  NAND2_X1 U9408 ( .A1(n9098), .A2(n7116), .ZN(n7114) );
  AOI21_X1 U9409 ( .B1(n9098), .B2(n9099), .A(n7118), .ZN(n9114) );
  NAND2_X1 U9410 ( .A1(n7122), .A2(n9297), .ZN(n7121) );
  OAI21_X1 U9411 ( .B1(n9273), .B2(n15058), .A(n7123), .ZN(n7122) );
  NAND2_X1 U9412 ( .A1(n9273), .A2(n9272), .ZN(n7123) );
  AND2_X2 U9413 ( .A1(n13611), .A2(n12273), .ZN(n13562) );
  NAND2_X1 U9414 ( .A1(n13545), .A2(n7542), .ZN(n13613) );
  NAND2_X2 U9415 ( .A1(n7126), .A2(n7124), .ZN(n11201) );
  NAND2_X1 U9416 ( .A1(n13570), .A2(n7130), .ZN(n7128) );
  NOR2_X1 U9417 ( .A1(n7149), .A2(n11323), .ZN(n7148) );
  NAND2_X1 U9418 ( .A1(n7158), .A2(n7548), .ZN(n7616) );
  NOR2_X1 U9419 ( .A1(n11075), .A2(n6698), .ZN(n11073) );
  NAND2_X1 U9420 ( .A1(n9771), .A2(n7162), .ZN(n11075) );
  NAND2_X1 U9421 ( .A1(n7172), .A2(n7170), .ZN(n12377) );
  NAND3_X1 U9422 ( .A1(n9819), .A2(n12711), .A3(n9820), .ZN(n12442) );
  NAND2_X1 U9423 ( .A1(n12442), .A2(n9820), .ZN(n9824) );
  NAND2_X1 U9424 ( .A1(n9819), .A2(n9820), .ZN(n12441) );
  INV_X1 U9425 ( .A(n7175), .ZN(n11238) );
  OAI21_X1 U9426 ( .B1(n7180), .B2(n7178), .A(n9792), .ZN(n7177) );
  NAND2_X2 U9427 ( .A1(n13517), .A2(n12234), .ZN(n12238) );
  NAND2_X1 U9428 ( .A1(n9703), .A2(n9702), .ZN(n9714) );
  OAI21_X1 U9429 ( .B1(n12483), .B2(n9802), .A(n9801), .ZN(n12410) );
  NAND2_X1 U9430 ( .A1(n12377), .A2(n9814), .ZN(n9818) );
  OAI22_X1 U9431 ( .A1(n11927), .A2(n9800), .B1(n12486), .B2(n9799), .ZN(
        n12483) );
  NAND2_X1 U9432 ( .A1(n12587), .A2(n12586), .ZN(n7194) );
  OR2_X1 U9433 ( .A1(n12554), .A2(n12575), .ZN(n7197) );
  NAND2_X1 U9434 ( .A1(n12584), .A2(n7196), .ZN(n7193) );
  NAND2_X1 U9435 ( .A1(n7197), .A2(n12584), .ZN(n12555) );
  OR2_X1 U9436 ( .A1(n9390), .A2(n10128), .ZN(n7203) );
  INV_X1 U9437 ( .A(n11106), .ZN(n11161) );
  NAND2_X1 U9438 ( .A1(n9919), .A2(n7228), .ZN(n7224) );
  NAND2_X1 U9439 ( .A1(n7229), .A2(n7230), .ZN(n10024) );
  NAND3_X1 U9440 ( .A1(n10019), .A2(n6740), .A3(n10018), .ZN(n7229) );
  NAND2_X1 U9441 ( .A1(n7232), .A2(n7233), .ZN(n10003) );
  NAND3_X1 U9442 ( .A1(n9997), .A2(n6735), .A3(n9996), .ZN(n7232) );
  NAND2_X1 U9443 ( .A1(n7234), .A2(n7235), .ZN(n10014) );
  NAND3_X1 U9444 ( .A1(n10008), .A2(n6739), .A3(n10007), .ZN(n7234) );
  NAND2_X1 U9445 ( .A1(n7236), .A2(n7237), .ZN(n9948) );
  NAND3_X1 U9446 ( .A1(n9942), .A2(n6736), .A3(n9941), .ZN(n7236) );
  NAND2_X1 U9447 ( .A1(n9990), .A2(n7243), .ZN(n7241) );
  NAND2_X1 U9448 ( .A1(n7241), .A2(n7239), .ZN(n9994) );
  NAND2_X1 U9449 ( .A1(n7248), .A2(n7246), .ZN(n9939) );
  NAND2_X1 U9450 ( .A1(n9955), .A2(n7251), .ZN(n7252) );
  NAND2_X1 U9451 ( .A1(n7252), .A2(n7254), .ZN(n9971) );
  INV_X1 U9452 ( .A(n7263), .ZN(n10114) );
  OAI211_X1 U9453 ( .C1(n10064), .C2(n7269), .A(n7265), .B(n7264), .ZN(n7263)
         );
  NAND2_X1 U9454 ( .A1(n10064), .A2(n7270), .ZN(n7264) );
  AND2_X1 U9455 ( .A1(n9586), .A2(n6742), .ZN(n9712) );
  AND2_X1 U9456 ( .A1(n9586), .A2(n9585), .ZN(n9703) );
  NAND2_X1 U9457 ( .A1(n9586), .A2(n7279), .ZN(n9710) );
  OAI21_X1 U9458 ( .B1(n12164), .B2(n8273), .A(n9037), .ZN(n10844) );
  NAND2_X1 U9459 ( .A1(n13218), .A2(n7290), .ZN(n7288) );
  NAND2_X1 U9460 ( .A1(n9067), .A2(n7300), .ZN(n7298) );
  NAND2_X1 U9461 ( .A1(n13345), .A2(n9060), .ZN(n7303) );
  NAND2_X1 U9462 ( .A1(n7303), .A2(n7304), .ZN(n9063) );
  XNOR2_X2 U9463 ( .A(n8214), .B(n8233), .ZN(n8917) );
  NAND3_X1 U9464 ( .A1(n8917), .A2(n12214), .A3(n14667), .ZN(n7310) );
  OAI21_X2 U9465 ( .B1(n11293), .B2(n9053), .A(n7312), .ZN(n11501) );
  NAND3_X1 U9466 ( .A1(n10583), .A2(n9041), .A3(n6667), .ZN(n7314) );
  NAND2_X1 U9467 ( .A1(n13975), .A2(n13976), .ZN(n13974) );
  NAND2_X1 U9468 ( .A1(n13842), .A2(n6726), .ZN(n7324) );
  OAI21_X1 U9469 ( .B1(n13842), .B2(n13854), .A(n7335), .ZN(n13825) );
  NAND2_X1 U9470 ( .A1(n6741), .A2(n11154), .ZN(n11307) );
  INV_X1 U9471 ( .A(n9890), .ZN(n10715) );
  NAND2_X1 U9472 ( .A1(n11907), .A2(n7337), .ZN(n13995) );
  OAI21_X1 U9473 ( .B1(n9406), .B2(n7352), .A(n7350), .ZN(n10898) );
  NAND2_X1 U9474 ( .A1(n7350), .A2(n7352), .ZN(n7348) );
  NAND2_X1 U9475 ( .A1(n9406), .A2(n7350), .ZN(n7349) );
  AOI21_X1 U9476 ( .B1(n7351), .B2(n14516), .A(n6697), .ZN(n7350) );
  NAND2_X1 U9477 ( .A1(n11306), .A2(n7354), .ZN(n7353) );
  NAND2_X1 U9478 ( .A1(n7353), .A2(n7356), .ZN(n11463) );
  NAND2_X1 U9479 ( .A1(n14052), .A2(n7364), .ZN(n7368) );
  NAND2_X1 U9480 ( .A1(n14052), .A2(n6638), .ZN(n13836) );
  NAND2_X1 U9481 ( .A1(n13834), .A2(n13845), .ZN(n7367) );
  NAND2_X1 U9482 ( .A1(n9676), .A2(n7372), .ZN(n9323) );
  OAI21_X2 U9483 ( .B1(n13973), .B2(n9584), .A(n9981), .ZN(n13952) );
  OAI21_X2 U9484 ( .B1(n13990), .B2(n9572), .A(n9573), .ZN(n13973) );
  NAND2_X1 U9485 ( .A1(n7380), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8194) );
  NAND2_X1 U9486 ( .A1(n11119), .A2(n8473), .ZN(n7381) );
  NAND3_X1 U9487 ( .A1(n7387), .A2(n7386), .A3(n8374), .ZN(n10692) );
  NAND3_X1 U9488 ( .A1(n7388), .A2(n7389), .A3(n7392), .ZN(n7386) );
  NAND3_X1 U9489 ( .A1(n7388), .A2(n13027), .A3(n7389), .ZN(n7387) );
  NAND2_X1 U9490 ( .A1(n8863), .A2(n7394), .ZN(n7393) );
  OAI211_X1 U9491 ( .C1(n8863), .C2(n7396), .A(n7399), .B(n7393), .ZN(n8933)
         );
  INV_X1 U9492 ( .A(n8862), .ZN(n7401) );
  XNOR2_X1 U9493 ( .A(n8196), .B(n12131), .ZN(n7403) );
  NAND2_X1 U9494 ( .A1(n7403), .A2(n8904), .ZN(n9077) );
  INV_X4 U9495 ( .A(n8834), .ZN(n8860) );
  NAND2_X1 U9496 ( .A1(n11019), .A2(n11020), .ZN(n8447) );
  INV_X1 U9497 ( .A(n10826), .ZN(n7408) );
  NAND3_X1 U9498 ( .A1(n8221), .A2(n8248), .A3(n8225), .ZN(n8252) );
  NAND2_X1 U9499 ( .A1(n10039), .A2(n10038), .ZN(n7423) );
  NAND2_X1 U9500 ( .A1(n8787), .A2(n8766), .ZN(n8769) );
  INV_X1 U9501 ( .A(n7433), .ZN(n7432) );
  AND2_X1 U9502 ( .A1(n7563), .A2(n7564), .ZN(n7438) );
  INV_X2 U9503 ( .A(n12505), .ZN(n7578) );
  OAI21_X2 U9504 ( .B1(n12789), .B2(n7446), .A(n7443), .ZN(n12757) );
  NAND2_X1 U9505 ( .A1(n12720), .A2(n6668), .ZN(n7448) );
  NAND2_X1 U9506 ( .A1(n7691), .A2(n7690), .ZN(n11711) );
  INV_X1 U9507 ( .A(n7690), .ZN(n7456) );
  NAND2_X1 U9508 ( .A1(n7457), .A2(n6729), .ZN(n8949) );
  AND4_X2 U9509 ( .A1(n7635), .A2(n6642), .A3(n6629), .A4(n7458), .ZN(n8068)
         );
  AND2_X1 U9510 ( .A1(n8152), .A2(n7464), .ZN(n8116) );
  NAND2_X1 U9511 ( .A1(n13264), .A2(n12977), .ZN(n7475) );
  NAND2_X1 U9512 ( .A1(n7480), .A2(n7481), .ZN(n13165) );
  INV_X1 U9513 ( .A(n7483), .ZN(n13182) );
  INV_X1 U9514 ( .A(n13186), .ZN(n7482) );
  AOI21_X1 U9515 ( .B1(n13205), .B2(n7487), .A(n7485), .ZN(n7484) );
  AND2_X1 U9516 ( .A1(n13388), .A2(n12988), .ZN(n7485) );
  NAND2_X1 U9517 ( .A1(n6624), .A2(n7506), .ZN(n8235) );
  XNOR2_X2 U9518 ( .A(n8193), .B(n8864), .ZN(n12131) );
  AND2_X2 U9519 ( .A1(n8912), .A2(n11208), .ZN(n12161) );
  NAND2_X1 U9520 ( .A1(n7509), .A2(n7510), .ZN(n12017) );
  NAND3_X1 U9521 ( .A1(n12010), .A2(n6737), .A3(n12009), .ZN(n7509) );
  NAND2_X1 U9522 ( .A1(n7511), .A2(n7512), .ZN(n12038) );
  NAND3_X1 U9523 ( .A1(n12030), .A2(n6738), .A3(n12029), .ZN(n7511) );
  NAND2_X1 U9524 ( .A1(n7515), .A2(n7516), .ZN(n12110) );
  NAND2_X1 U9525 ( .A1(n12105), .A2(n12107), .ZN(n7516) );
  OAI211_X1 U9526 ( .C1(n11986), .C2(n11984), .A(n11982), .B(n11981), .ZN(
        n7518) );
  NAND2_X1 U9527 ( .A1(n7522), .A2(n7523), .ZN(n12096) );
  XNOR2_X1 U9528 ( .A(n8937), .B(n9128), .ZN(n8939) );
  OAI21_X1 U9529 ( .B1(n8952), .B2(n15016), .A(n8951), .ZN(n8953) );
  NAND2_X1 U9530 ( .A1(n11674), .A2(n11673), .ZN(n11749) );
  NAND2_X1 U9531 ( .A1(n11604), .A2(n11605), .ZN(n11674) );
  INV_X1 U9532 ( .A(n10610), .ZN(n10608) );
  NAND2_X1 U9533 ( .A1(n9710), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9711) );
  OAI21_X1 U9534 ( .B1(n9710), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9704) );
  CLKBUF_X1 U9535 ( .A(n13552), .Z(n13555) );
  OR2_X1 U9536 ( .A1(n7675), .A2(n11429), .ZN(n7623) );
  NAND2_X1 U9537 ( .A1(n13561), .A2(n6747), .ZN(n13621) );
  NAND2_X1 U9538 ( .A1(n15038), .A2(n9136), .ZN(n15025) );
  XNOR2_X1 U9539 ( .A(n10039), .B(n10038), .ZN(n13486) );
  INV_X1 U9540 ( .A(n9712), .ZN(n9716) );
  OAI21_X1 U9541 ( .B1(n9982), .B2(n9981), .A(n9980), .ZN(n9983) );
  INV_X1 U9542 ( .A(n9363), .ZN(n10605) );
  NAND2_X2 U9543 ( .A1(n10354), .A2(n11201), .ZN(n10341) );
  OR2_X1 U9544 ( .A1(n7715), .A2(n11951), .ZN(n7580) );
  XNOR2_X1 U9545 ( .A(n11029), .B(n11028), .ZN(n10956) );
  NAND2_X1 U9546 ( .A1(n13535), .A2(n10953), .ZN(n11029) );
  CLKBUF_X1 U9547 ( .A(n13036), .Z(n13040) );
  OR2_X1 U9548 ( .A1(n9325), .A2(n14138), .ZN(n9326) );
  NAND2_X1 U9549 ( .A1(n7541), .A2(n10112), .ZN(n10113) );
  NAND2_X1 U9550 ( .A1(n13812), .A2(n9663), .ZN(n9672) );
  NAND2_X1 U9551 ( .A1(n13112), .A2(n8272), .ZN(n8263) );
  OAI21_X1 U9552 ( .B1(n6728), .B2(n8105), .A(n12664), .ZN(n12832) );
  OAI21_X1 U9553 ( .B1(n14030), .B2(n14009), .A(n9737), .ZN(n9763) );
  CLKBUF_X1 U9554 ( .A(n8657), .Z(n9032) );
  NOR2_X2 U9555 ( .A1(n11033), .A2(n11032), .ZN(n11173) );
  NAND2_X1 U9556 ( .A1(n8129), .A2(n8128), .ZN(n8130) );
  INV_X1 U9557 ( .A(n8238), .ZN(n13484) );
  AND2_X1 U9558 ( .A1(n14822), .A2(n11284), .ZN(n9091) );
  OR2_X1 U9559 ( .A1(n7568), .A2(n8127), .ZN(n7570) );
  NOR2_X1 U9560 ( .A1(n15061), .A2(n11954), .ZN(n9131) );
  AND2_X2 U9561 ( .A1(n7565), .A2(n12938), .ZN(n7605) );
  NOR2_X1 U9562 ( .A1(n13168), .A2(n13167), .ZN(n13379) );
  AND2_X1 U9563 ( .A1(n9897), .A2(n10086), .ZN(n7529) );
  NAND2_X1 U9564 ( .A1(n8913), .A2(n13354), .ZN(n13081) );
  INV_X1 U9565 ( .A(n15057), .ZN(n7577) );
  AND2_X2 U9566 ( .A1(n11066), .A2(n8172), .ZN(n15132) );
  OR2_X1 U9567 ( .A1(n12639), .A2(n12882), .ZN(n7530) );
  OR2_X1 U9568 ( .A1(n12639), .A2(n12926), .ZN(n7531) );
  NOR2_X1 U9569 ( .A1(n12622), .A2(n12926), .ZN(n8158) );
  INV_X1 U9570 ( .A(n15119), .ZN(n8156) );
  AND2_X1 U9571 ( .A1(n8924), .A2(n8906), .ZN(n13049) );
  AND2_X1 U9572 ( .A1(n7605), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7532) );
  NOR2_X1 U9573 ( .A1(n8098), .A2(n12787), .ZN(n7534) );
  INV_X1 U9574 ( .A(n12763), .ZN(n7880) );
  AND2_X1 U9575 ( .A1(n9665), .A2(n14520), .ZN(n7535) );
  NOR2_X1 U9576 ( .A1(n9879), .A2(n9719), .ZN(n10354) );
  NAND2_X1 U9577 ( .A1(n13357), .A2(n10733), .ZN(n13369) );
  INV_X1 U9578 ( .A(n12196), .ZN(n9024) );
  INV_X1 U9579 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7557) );
  INV_X1 U9580 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7559) );
  INV_X1 U9581 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7558) );
  AND2_X1 U9582 ( .A1(n6627), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7538) );
  INV_X1 U9583 ( .A(n11103), .ZN(n11107) );
  INV_X1 U9584 ( .A(n14835), .ZN(n14837) );
  AND2_X1 U9585 ( .A1(n9673), .A2(n9318), .ZN(n7539) );
  INV_X1 U9586 ( .A(n12748), .ZN(n7900) );
  AND2_X1 U9587 ( .A1(n9484), .A2(n9483), .ZN(n7540) );
  CLKBUF_X3 U9588 ( .A(n8272), .Z(n13336) );
  INV_X1 U9589 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7920) );
  XOR2_X1 U9590 ( .A(n10110), .B(n13944), .Z(n7541) );
  INV_X1 U9591 ( .A(n13991), .ZN(n9755) );
  INV_X1 U9592 ( .A(n11327), .ZN(n11177) );
  INV_X1 U9593 ( .A(n11640), .ZN(n11698) );
  INV_X1 U9594 ( .A(n15016), .ZN(n8938) );
  NOR2_X1 U9595 ( .A1(n12363), .A2(n12364), .ZN(n7544) );
  INV_X1 U9596 ( .A(n12667), .ZN(n8105) );
  NAND2_X1 U9597 ( .A1(n12691), .A2(n12690), .ZN(n12692) );
  AND2_X1 U9598 ( .A1(n12641), .A2(n15115), .ZN(n7545) );
  AND2_X1 U9599 ( .A1(n9568), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7547) );
  INV_X1 U9600 ( .A(n9363), .ZN(n10359) );
  NAND2_X1 U9601 ( .A1(n11972), .A2(n11971), .ZN(n11969) );
  AND2_X1 U9602 ( .A1(n11970), .A2(n11969), .ZN(n11975) );
  NAND2_X1 U9603 ( .A1(n11975), .A2(n11974), .ZN(n11977) );
  MUX2_X1 U9604 ( .A(n9896), .B(n9895), .S(n9894), .Z(n9897) );
  NAND2_X1 U9605 ( .A1(n12078), .A2(n12077), .ZN(n12080) );
  INV_X1 U9606 ( .A(n9719), .ZN(n9882) );
  OR2_X1 U9607 ( .A1(n8019), .A2(n8018), .ZN(n8020) );
  INV_X1 U9608 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7550) );
  INV_X1 U9609 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8208) );
  INV_X1 U9610 ( .A(n14343), .ZN(n9122) );
  INV_X1 U9611 ( .A(n9257), .ZN(n8036) );
  INV_X1 U9612 ( .A(n15028), .ZN(n9278) );
  INV_X1 U9613 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8385) );
  INV_X1 U9614 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n7788) );
  INV_X1 U9615 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n12418) );
  OR2_X1 U9616 ( .A1(n7987), .A2(n12945), .ZN(n8024) );
  INV_X1 U9617 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9100) );
  INV_X1 U9618 ( .A(n8263), .ZN(n8265) );
  NOR2_X1 U9619 ( .A1(n8733), .A2(n13053), .ZN(n8749) );
  AND2_X1 U9620 ( .A1(n8773), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8791) );
  NOR2_X1 U9621 ( .A1(n8543), .A2(n8542), .ZN(n8564) );
  NAND2_X1 U9622 ( .A1(n9023), .A2(n9022), .ZN(n9078) );
  NAND2_X1 U9623 ( .A1(n10607), .A2(n10606), .ZN(n10610) );
  INV_X1 U9624 ( .A(n10950), .ZN(n10951) );
  INV_X1 U9625 ( .A(n12229), .ZN(n9531) );
  NAND2_X1 U9626 ( .A1(n8226), .A2(n8222), .ZN(n8223) );
  INV_X1 U9627 ( .A(n9779), .ZN(n9780) );
  NOR2_X1 U9628 ( .A1(n7837), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7859) );
  OR2_X1 U9629 ( .A1(n8044), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8056) );
  NAND2_X1 U9630 ( .A1(n7939), .A2(n7938), .ZN(n7950) );
  NAND2_X1 U9631 ( .A1(n12655), .A2(n12654), .ZN(n12653) );
  INV_X1 U9632 ( .A(n11845), .ZN(n11852) );
  NAND2_X1 U9633 ( .A1(n15011), .A2(n9155), .ZN(n14996) );
  XNOR2_X1 U9634 ( .A(n8860), .B(n11983), .ZN(n8246) );
  INV_X1 U9635 ( .A(n13081), .ZN(n8914) );
  OR2_X1 U9636 ( .A1(n8688), .A2(n13044), .ZN(n8711) );
  INV_X1 U9637 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8480) );
  OR2_X1 U9638 ( .A1(n8816), .A2(n8815), .ZN(n8851) );
  OR2_X1 U9639 ( .A1(n8711), .A2(n12978), .ZN(n8733) );
  AND2_X1 U9640 ( .A1(n8564), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8583) );
  INV_X1 U9641 ( .A(n13488), .ZN(n8239) );
  AND2_X1 U9642 ( .A1(n10463), .A2(n10462), .ZN(n10570) );
  NAND2_X1 U9643 ( .A1(n8583), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8613) );
  INV_X1 U9644 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9430) );
  OR2_X1 U9645 ( .A1(n12259), .A2(n12258), .ZN(n12260) );
  NAND2_X1 U9646 ( .A1(n10600), .A2(n10599), .ZN(n10601) );
  INV_X1 U9647 ( .A(n11029), .ZN(n11030) );
  NAND2_X1 U9648 ( .A1(n10952), .A2(n10951), .ZN(n10953) );
  INV_X1 U9649 ( .A(n9347), .ZN(n9644) );
  INV_X1 U9650 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n15330) );
  NAND2_X1 U9651 ( .A1(n8603), .A2(SI_17_), .ZN(n8624) );
  INV_X4 U9652 ( .A(n7572), .ZN(n10067) );
  INV_X1 U9653 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9313) );
  NAND2_X1 U9654 ( .A1(n9780), .A2(n12503), .ZN(n9781) );
  NOR2_X1 U9655 ( .A1(n7909), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n7924) );
  AND2_X1 U9656 ( .A1(n7859), .A2(n7858), .ZN(n7874) );
  OR2_X1 U9657 ( .A1(n7745), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7767) );
  INV_X1 U9658 ( .A(n12487), .ZN(n12465) );
  INV_X1 U9659 ( .A(n8056), .ZN(n12611) );
  INV_X1 U9660 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11885) );
  INV_X1 U9661 ( .A(n9118), .ZN(n12622) );
  NAND2_X1 U9662 ( .A1(n8108), .A2(n9252), .ZN(n8947) );
  AND3_X1 U9663 ( .A1(n8008), .A2(n8007), .A3(n8006), .ZN(n12671) );
  INV_X1 U9664 ( .A(n12722), .ZN(n12700) );
  INV_X1 U9665 ( .A(n12719), .ZN(n8102) );
  INV_X1 U9666 ( .A(n12734), .ZN(n12758) );
  NOR2_X1 U9667 ( .A1(n7767), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7789) );
  OR2_X1 U9668 ( .A1(n7657), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7673) );
  OR2_X1 U9669 ( .A1(n11063), .A2(n11939), .ZN(n8164) );
  OR2_X1 U9670 ( .A1(n7987), .A2(n12942), .ZN(n8042) );
  INV_X1 U9671 ( .A(n11828), .ZN(n11834) );
  NAND3_X1 U9672 ( .A1(n10754), .A2(n10768), .A3(n10752), .ZN(n15045) );
  AND2_X1 U9673 ( .A1(n8146), .A2(n9126), .ZN(n15016) );
  NAND2_X1 U9674 ( .A1(n7886), .A2(n7885), .ZN(n7903) );
  NAND2_X1 U9675 ( .A1(n7828), .A2(n7827), .ZN(n7846) );
  INV_X1 U9676 ( .A(n12951), .ZN(n12952) );
  INV_X1 U9677 ( .A(n13377), .ZN(n8916) );
  OR2_X1 U9678 ( .A1(n8613), .A2(n8612), .ZN(n8634) );
  NOR2_X1 U9679 ( .A1(n8926), .A2(n14772), .ZN(n8924) );
  AND2_X1 U9680 ( .A1(n8851), .A2(n8817), .ZN(n13202) );
  NAND2_X1 U9681 ( .A1(n13475), .A2(n12137), .ZN(n12139) );
  NAND2_X1 U9682 ( .A1(n9015), .A2(n9014), .ZN(n9025) );
  INV_X1 U9683 ( .A(n13314), .ZN(n9064) );
  INV_X1 U9684 ( .A(n13349), .ZN(n9059) );
  INV_X1 U9685 ( .A(n13366), .ZN(n14764) );
  INV_X1 U9686 ( .A(n14826), .ZN(n14792) );
  NOR2_X1 U9687 ( .A1(n11031), .A2(n11030), .ZN(n11032) );
  NAND2_X1 U9688 ( .A1(n10603), .A2(n10709), .ZN(n10351) );
  AND2_X1 U9689 ( .A1(n9730), .A2(n9657), .ZN(n13817) );
  INV_X1 U9690 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14177) );
  INV_X1 U9691 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14184) );
  INV_X1 U9692 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n11677) );
  INV_X1 U9693 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14188) );
  NAND2_X1 U9694 ( .A1(n10357), .A2(n9717), .ZN(n10514) );
  INV_X1 U9695 ( .A(n13841), .ZN(n13854) );
  AND2_X1 U9696 ( .A1(n9540), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9554) );
  OR2_X1 U9697 ( .A1(n9510), .A2(n9509), .ZN(n9525) );
  NOR2_X1 U9698 ( .A1(n9484), .A2(n9483), .ZN(n9493) );
  OR2_X1 U9699 ( .A1(n10353), .A2(n10352), .ZN(n10513) );
  NAND2_X1 U9700 ( .A1(n10356), .A2(n10355), .ZN(n14635) );
  NAND2_X1 U9701 ( .A1(n9424), .A2(n9423), .ZN(n14500) );
  INV_X1 U9702 ( .A(n10086), .ZN(n14531) );
  INV_X1 U9703 ( .A(n14152), .ZN(n9697) );
  INV_X1 U9704 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9321) );
  AND2_X1 U9705 ( .A1(n8474), .A2(n8452), .ZN(n8453) );
  AND2_X1 U9706 ( .A1(n8375), .A2(n8354), .ZN(n8355) );
  INV_X1 U9707 ( .A(n8231), .ZN(n8228) );
  NOR2_X1 U9708 ( .A1(n9866), .A2(n15045), .ZN(n12487) );
  OR2_X1 U9709 ( .A1(n7735), .A2(n11661), .ZN(n7973) );
  NAND2_X1 U9710 ( .A1(n11047), .A2(n11204), .ZN(n12493) );
  AOI21_X1 U9711 ( .B1(n12627), .B2(n6627), .A(n8050), .ZN(n9868) );
  AND3_X1 U9712 ( .A1(n7967), .A2(n7966), .A3(n7965), .ZN(n12699) );
  INV_X1 U9713 ( .A(n12604), .ZN(n14992) );
  NAND2_X1 U9714 ( .A1(n8955), .A2(n8954), .ZN(n12636) );
  INV_X1 U9715 ( .A(n15045), .ZN(n15062) );
  NAND2_X1 U9716 ( .A1(n8114), .A2(n8165), .ZN(n14997) );
  OR2_X1 U9717 ( .A1(n14997), .A2(n15049), .ZN(n15019) );
  INV_X1 U9718 ( .A(n15071), .ZN(n12766) );
  AND2_X1 U9719 ( .A1(n8164), .A2(n8163), .ZN(n11066) );
  OR2_X1 U9720 ( .A1(n14997), .A2(n15115), .ZN(n15101) );
  AND2_X1 U9721 ( .A1(n10119), .A2(n11046), .ZN(n10749) );
  AND2_X1 U9722 ( .A1(n8081), .A2(n10752), .ZN(n15059) );
  INV_X1 U9723 ( .A(n8134), .ZN(n10399) );
  AND2_X1 U9724 ( .A1(n7637), .A2(n7636), .ZN(n11430) );
  OAI21_X1 U9725 ( .B1(n13166), .B2(n13079), .A(n8930), .ZN(n8931) );
  AND2_X1 U9726 ( .A1(n8841), .A2(n8840), .ZN(n9012) );
  AND3_X1 U9727 ( .A1(n8617), .A2(n8616), .A3(n8615), .ZN(n13061) );
  AND4_X1 U9728 ( .A1(n8508), .A2(n8507), .A3(n8506), .A4(n8505), .ZN(n9052)
         );
  OR2_X1 U9729 ( .A1(n14693), .A2(n14692), .ZN(n14694) );
  INV_X1 U9730 ( .A(n14718), .ZN(n14752) );
  AND2_X1 U9731 ( .A1(n10190), .A2(n10189), .ZN(n14729) );
  INV_X1 U9732 ( .A(n12189), .ZN(n13270) );
  INV_X1 U9733 ( .A(n12179), .ZN(n11261) );
  NAND2_X1 U9734 ( .A1(n12213), .A2(n10502), .ZN(n14826) );
  INV_X1 U9735 ( .A(n14808), .ZN(n13456) );
  OR2_X1 U9736 ( .A1(n11006), .A2(n14822), .ZN(n14808) );
  AND2_X1 U9737 ( .A1(n13496), .A2(n8884), .ZN(n14771) );
  AND2_X1 U9738 ( .A1(n8871), .A2(n8870), .ZN(n13496) );
  AND2_X1 U9739 ( .A1(n8499), .A2(n8539), .ZN(n11552) );
  INV_X1 U9740 ( .A(n13660), .ZN(n13634) );
  NAND2_X1 U9741 ( .A1(n10362), .A2(n13962), .ZN(n13658) );
  AND4_X1 U9742 ( .A1(n9640), .A2(n9639), .A3(n9638), .A4(n9637), .ZN(n13916)
         );
  AND2_X1 U9743 ( .A1(n9612), .A2(n9611), .ZN(n14103) );
  AND4_X1 U9744 ( .A1(n9545), .A2(n9544), .A3(n9543), .A4(n9542), .ZN(n14409)
         );
  INV_X1 U9745 ( .A(n14477), .ZN(n14489) );
  INV_X1 U9746 ( .A(n13930), .ZN(n13944) );
  INV_X1 U9747 ( .A(n13902), .ZN(n14548) );
  NAND2_X1 U9748 ( .A1(n9731), .A2(n13962), .ZN(n14006) );
  INV_X1 U9749 ( .A(n10513), .ZN(n10519) );
  INV_X1 U9750 ( .A(n14376), .ZN(n14533) );
  AND2_X1 U9751 ( .A1(n14602), .A2(n14601), .ZN(n14563) );
  INV_X1 U9752 ( .A(n14602), .ZN(n14536) );
  INV_X1 U9753 ( .A(n14563), .ZN(n14642) );
  INV_X1 U9754 ( .A(n14408), .ZN(n14617) );
  AND3_X1 U9755 ( .A1(n10518), .A2(n10517), .A3(n10516), .ZN(n14120) );
  NAND2_X1 U9756 ( .A1(n9685), .A2(n9697), .ZN(n10202) );
  INV_X1 U9757 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14211) );
  AND2_X1 U9758 ( .A1(n14255), .A2(n14254), .ZN(n14451) );
  OR2_X1 U9759 ( .A1(n11944), .A2(n8151), .ZN(n10119) );
  AND2_X1 U9760 ( .A1(n10784), .A2(n10783), .ZN(n14978) );
  INV_X1 U9761 ( .A(n12493), .ZN(n11768) );
  OR2_X1 U9762 ( .A1(n9303), .A2(n9302), .ZN(n9304) );
  INV_X1 U9763 ( .A(n14978), .ZN(n14952) );
  INV_X1 U9764 ( .A(n14960), .ZN(n14986) );
  OR2_X1 U9765 ( .A1(n10781), .A2(n10768), .ZN(n14994) );
  NAND2_X1 U9766 ( .A1(n15074), .A2(n15019), .ZN(n12822) );
  NAND2_X2 U9767 ( .A1(n11069), .A2(n12766), .ZN(n15074) );
  INV_X1 U9768 ( .A(n9838), .ZN(n12826) );
  NAND2_X1 U9769 ( .A1(n15132), .A2(n14345), .ZN(n12882) );
  INV_X1 U9770 ( .A(n15132), .ZN(n15130) );
  INV_X1 U9771 ( .A(n12447), .ZN(n12892) );
  NAND2_X1 U9772 ( .A1(n7823), .A2(n7822), .ZN(n12918) );
  AND2_X2 U9773 ( .A1(n8155), .A2(n10749), .ZN(n15119) );
  NOR2_X2 U9774 ( .A1(n10399), .A2(n11938), .ZN(n10637) );
  CLKBUF_X1 U9775 ( .A(n10637), .Z(n10653) );
  NAND2_X1 U9776 ( .A1(n8125), .A2(n8124), .ZN(n11740) );
  INV_X1 U9777 ( .A(n8166), .ZN(n10875) );
  INV_X1 U9778 ( .A(SI_15_), .ZN(n15227) );
  INV_X1 U9779 ( .A(n14914), .ZN(n11424) );
  INV_X1 U9780 ( .A(n8931), .ZN(n8932) );
  INV_X1 U9781 ( .A(n13049), .ZN(n13083) );
  NAND2_X1 U9782 ( .A1(n8859), .A2(n8858), .ZN(n13087) );
  INV_X1 U9783 ( .A(n12969), .ZN(n13094) );
  INV_X1 U9784 ( .A(n9052), .ZN(n13102) );
  INV_X1 U9785 ( .A(n14729), .ZN(n14745) );
  AND2_X1 U9786 ( .A1(n13313), .A2(n13312), .ZN(n13434) );
  AND2_X1 U9787 ( .A1(n10499), .A2(n13354), .ZN(n14770) );
  AND3_X1 U9788 ( .A1(n10498), .A2(n9088), .A3(n9092), .ZN(n13457) );
  INV_X1 U9789 ( .A(n13457), .ZN(n14835) );
  OR2_X1 U9790 ( .A1(n13445), .A2(n13444), .ZN(n13472) );
  NAND3_X1 U9791 ( .A1(n9093), .A2(n10498), .A3(n9092), .ZN(n14829) );
  NOR2_X1 U9792 ( .A1(n14772), .A2(n14771), .ZN(n14775) );
  INV_X1 U9793 ( .A(n14775), .ZN(n14778) );
  INV_X1 U9794 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13499) );
  INV_X1 U9795 ( .A(n13913), .ZN(n14080) );
  NAND2_X1 U9796 ( .A1(n10361), .A2(n10358), .ZN(n13660) );
  INV_X1 U9797 ( .A(n13584), .ZN(n14394) );
  INV_X1 U9798 ( .A(n14486), .ZN(n14479) );
  INV_X1 U9799 ( .A(n13792), .ZN(n14494) );
  OR2_X1 U9800 ( .A1(n9731), .A2(n13944), .ZN(n13902) );
  AND2_X1 U9801 ( .A1(n14364), .A2(n14363), .ZN(n14403) );
  INV_X2 U9802 ( .A(n14006), .ZN(n14539) );
  OR2_X1 U9803 ( .A1(n14552), .A2(n10509), .ZN(n14009) );
  AND2_X2 U9804 ( .A1(n10519), .A2(n14120), .ZN(n14665) );
  AND3_X1 U9805 ( .A1(n14419), .A2(n14418), .A3(n14417), .ZN(n14436) );
  INV_X1 U9806 ( .A(n14645), .ZN(n14643) );
  AND2_X2 U9807 ( .A1(n14121), .A2(n14120), .ZN(n14645) );
  NAND2_X1 U9808 ( .A1(n10202), .A2(n10515), .ZN(n15133) );
  INV_X1 U9809 ( .A(n9327), .ZN(n14146) );
  INV_X1 U9810 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n14161) );
  INV_X1 U9811 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10806) );
  INV_X1 U9812 ( .A(n13113), .ZN(P2_U3947) );
  INV_X1 U9813 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n7556) );
  XNOR2_X2 U9814 ( .A(n7561), .B(P3_IR_REG_29__SCAN_IN), .ZN(n7562) );
  BUF_X2 U9815 ( .A(n7562), .Z(n7567) );
  AND2_X2 U9816 ( .A1(n7565), .A2(n7562), .ZN(n7589) );
  NAND2_X1 U9817 ( .A1(n7589), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7564) );
  NAND2_X1 U9818 ( .A1(n7605), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7563) );
  INV_X1 U9819 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n7566) );
  INV_X1 U9820 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10913) );
  INV_X1 U9821 ( .A(SI_1_), .ZN(n10160) );
  OR2_X1 U9822 ( .A1(n6625), .A2(n10160), .ZN(n7576) );
  AND2_X2 U9823 ( .A1(n7585), .A2(n10067), .ZN(n7610) );
  XNOR2_X1 U9824 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7595) );
  INV_X1 U9825 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8271) );
  XNOR2_X1 U9826 ( .A(n7595), .B(n7594), .ZN(n10159) );
  NAND2_X1 U9827 ( .A1(n7610), .A2(n10159), .ZN(n7575) );
  INV_X1 U9828 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n10778) );
  NAND2_X1 U9829 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7573) );
  XNOR2_X1 U9830 ( .A(n7573), .B(n10778), .ZN(n10774) );
  OR2_X1 U9831 ( .A1(n7585), .A2(n10774), .ZN(n7574) );
  NAND2_X2 U9832 ( .A1(n7578), .A2(n7577), .ZN(n9140) );
  NAND2_X1 U9833 ( .A1(n12505), .A2(n15057), .ZN(n9138) );
  INV_X1 U9834 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11951) );
  NOR2_X1 U9835 ( .A1(n7532), .A2(n7538), .ZN(n7579) );
  AND2_X1 U9836 ( .A1(n7580), .A2(n7579), .ZN(n7582) );
  INV_X1 U9837 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10757) );
  NAND2_X2 U9838 ( .A1(n7582), .A2(n7581), .ZN(n15061) );
  INV_X1 U9839 ( .A(SI_0_), .ZN(n10132) );
  INV_X1 U9840 ( .A(n7594), .ZN(n7584) );
  INV_X1 U9841 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8222) );
  NAND2_X1 U9842 ( .A1(n8222), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7583) );
  NAND2_X1 U9843 ( .A1(n7584), .A2(n7583), .ZN(n10130) );
  NAND2_X1 U9844 ( .A1(n7610), .A2(n10130), .ZN(n7587) );
  OR2_X1 U9845 ( .A1(n7585), .A2(n10803), .ZN(n7586) );
  NAND2_X1 U9846 ( .A1(n15061), .A2(n11947), .ZN(n15064) );
  NAND2_X1 U9847 ( .A1(n9129), .A2(n15064), .ZN(n15063) );
  NAND2_X1 U9848 ( .A1(n7578), .A2(n15057), .ZN(n7588) );
  NAND2_X1 U9849 ( .A1(n15063), .A2(n7588), .ZN(n15042) );
  NAND2_X1 U9850 ( .A1(n7810), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n7593) );
  INV_X1 U9851 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10759) );
  OR2_X1 U9852 ( .A1(n7675), .A2(n10759), .ZN(n7592) );
  NAND2_X1 U9853 ( .A1(n7605), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7591) );
  NAND2_X1 U9854 ( .A1(n7595), .A2(n7594), .ZN(n7597) );
  INV_X1 U9855 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10121) );
  NAND2_X1 U9856 ( .A1(n10121), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7596) );
  NAND2_X1 U9857 ( .A1(n7597), .A2(n7596), .ZN(n7612) );
  INV_X1 U9858 ( .A(n7611), .ZN(n7598) );
  XNOR2_X1 U9859 ( .A(n7612), .B(n7598), .ZN(n10133) );
  NAND2_X1 U9860 ( .A1(n7610), .A2(n10133), .ZN(n7602) );
  INV_X1 U9861 ( .A(n10754), .ZN(n7600) );
  INV_X1 U9862 ( .A(n10773), .ZN(n7599) );
  NAND2_X1 U9863 ( .A1(n15042), .A2(n15041), .ZN(n15040) );
  INV_X1 U9864 ( .A(n15060), .ZN(n11242) );
  NAND2_X1 U9865 ( .A1(n11242), .A2(n15050), .ZN(n7603) );
  AND2_X2 U9866 ( .A1(n15040), .A2(n7603), .ZN(n15029) );
  INV_X1 U9867 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n7604) );
  NAND2_X1 U9868 ( .A1(n7810), .A2(n7604), .ZN(n7609) );
  NAND2_X1 U9869 ( .A1(n7622), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7608) );
  NAND2_X1 U9870 ( .A1(n7605), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7607) );
  INV_X1 U9871 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n14850) );
  OR2_X1 U9872 ( .A1(n7675), .A2(n14850), .ZN(n7606) );
  NAND4_X1 U9873 ( .A1(n7609), .A2(n7608), .A3(n7607), .A4(n7606), .ZN(n12504)
         );
  NAND2_X1 U9874 ( .A1(n7612), .A2(n7611), .ZN(n7614) );
  INV_X1 U9875 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10122) );
  NAND2_X1 U9876 ( .A1(n10122), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7613) );
  NAND2_X1 U9877 ( .A1(n7614), .A2(n7613), .ZN(n7628) );
  INV_X1 U9878 ( .A(n7627), .ZN(n7615) );
  XNOR2_X1 U9879 ( .A(n7628), .B(n7615), .ZN(n10135) );
  NAND2_X1 U9880 ( .A1(n7610), .A2(n10135), .ZN(n7619) );
  NAND2_X1 U9881 ( .A1(n7616), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7617) );
  XNOR2_X1 U9882 ( .A(n7617), .B(P3_IR_REG_3__SCAN_IN), .ZN(n14849) );
  OR2_X1 U9883 ( .A1(n10754), .A2(n14849), .ZN(n7618) );
  OAI211_X1 U9884 ( .C1(n7987), .C2(SI_3_), .A(n7619), .B(n7618), .ZN(n15033)
         );
  OR2_X1 U9885 ( .A1(n12504), .A2(n15033), .ZN(n9145) );
  NAND2_X1 U9886 ( .A1(n12504), .A2(n15033), .ZN(n9141) );
  INV_X1 U9887 ( .A(n15033), .ZN(n11244) );
  NAND2_X1 U9888 ( .A1(n12504), .A2(n11244), .ZN(n7620) );
  AND2_X1 U9889 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7621) );
  NOR2_X1 U9890 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7643) );
  OR2_X1 U9891 ( .A1(n7621), .A2(n7643), .ZN(n11459) );
  NAND2_X1 U9892 ( .A1(n7810), .A2(n11459), .ZN(n7625) );
  NAND2_X1 U9893 ( .A1(n6620), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7624) );
  INV_X1 U9894 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n11429) );
  NAND2_X1 U9895 ( .A1(n7628), .A2(n7627), .ZN(n7631) );
  INV_X1 U9896 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7629) );
  NAND2_X1 U9897 ( .A1(n7629), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7630) );
  NAND2_X1 U9898 ( .A1(n7631), .A2(n7630), .ZN(n7650) );
  INV_X1 U9899 ( .A(n7649), .ZN(n7632) );
  XNOR2_X1 U9900 ( .A(n7650), .B(n7632), .ZN(n10137) );
  NAND2_X1 U9901 ( .A1(n9106), .A2(n10137), .ZN(n7639) );
  NAND2_X1 U9902 ( .A1(n7633), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7634) );
  MUX2_X1 U9903 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7634), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n7637) );
  INV_X1 U9904 ( .A(n7635), .ZN(n7636) );
  OR2_X1 U9905 ( .A1(n10754), .A2(n11430), .ZN(n7638) );
  OAI211_X1 U9906 ( .C1(n7987), .C2(SI_4_), .A(n7639), .B(n7638), .ZN(n11458)
         );
  OR2_X1 U9907 ( .A1(n15026), .A2(n11458), .ZN(n9151) );
  NAND2_X1 U9908 ( .A1(n15026), .A2(n11458), .ZN(n9150) );
  NAND2_X1 U9909 ( .A1(n9151), .A2(n9150), .ZN(n11452) );
  INV_X1 U9910 ( .A(n11458), .ZN(n7640) );
  NAND2_X1 U9911 ( .A1(n15026), .A2(n7640), .ZN(n7641) );
  NAND2_X1 U9912 ( .A1(n7962), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7648) );
  NAND2_X1 U9913 ( .A1(n7643), .A2(n11344), .ZN(n7657) );
  OR2_X1 U9914 ( .A1(n7643), .A2(n11344), .ZN(n7644) );
  NAND2_X1 U9915 ( .A1(n7657), .A2(n7644), .ZN(n15021) );
  NAND2_X1 U9916 ( .A1(n7810), .A2(n15021), .ZN(n7647) );
  NAND2_X1 U9917 ( .A1(n6620), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7646) );
  INV_X1 U9918 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n14893) );
  OR2_X1 U9919 ( .A1(n7675), .A2(n14893), .ZN(n7645) );
  NAND4_X1 U9920 ( .A1(n7648), .A2(n7647), .A3(n7646), .A4(n7645), .ZN(n15002)
         );
  NAND2_X1 U9921 ( .A1(n7650), .A2(n7649), .ZN(n7652) );
  NAND2_X1 U9922 ( .A1(n10141), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7651) );
  NAND2_X1 U9923 ( .A1(n7652), .A2(n7651), .ZN(n7664) );
  INV_X1 U9924 ( .A(n7663), .ZN(n7653) );
  XNOR2_X1 U9925 ( .A(n7664), .B(n7653), .ZN(n10139) );
  NAND2_X1 U9926 ( .A1(n9106), .A2(n10139), .ZN(n7656) );
  OR2_X1 U9927 ( .A1(n7635), .A2(n8127), .ZN(n7654) );
  XNOR2_X1 U9928 ( .A(n7654), .B(P3_IR_REG_5__SCAN_IN), .ZN(n14892) );
  OR2_X1 U9929 ( .A1(n10754), .A2(n14892), .ZN(n7655) );
  OAI211_X1 U9930 ( .C1(n7735), .C2(SI_5_), .A(n7656), .B(n7655), .ZN(n15020)
         );
  OR2_X1 U9931 ( .A1(n15002), .A2(n15020), .ZN(n9155) );
  NAND2_X1 U9932 ( .A1(n15002), .A2(n15020), .ZN(n9159) );
  NAND2_X1 U9933 ( .A1(n9155), .A2(n9159), .ZN(n8091) );
  NAND2_X1 U9934 ( .A1(n7962), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7662) );
  NAND2_X1 U9935 ( .A1(n7657), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7658) );
  NAND2_X1 U9936 ( .A1(n7673), .A2(n7658), .ZN(n15007) );
  NAND2_X1 U9937 ( .A1(n7810), .A2(n15007), .ZN(n7661) );
  NAND2_X1 U9938 ( .A1(n8076), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7660) );
  INV_X1 U9939 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11396) );
  OR2_X1 U9940 ( .A1(n7675), .A2(n11396), .ZN(n7659) );
  NAND4_X1 U9941 ( .A1(n7662), .A2(n7661), .A3(n7660), .A4(n7659), .ZN(n12503)
         );
  NAND2_X1 U9942 ( .A1(n7664), .A2(n7663), .ZN(n7666) );
  NAND2_X1 U9943 ( .A1(n10147), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7665) );
  XNOR2_X1 U9944 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n7667) );
  XNOR2_X1 U9945 ( .A(n7681), .B(n7667), .ZN(n10165) );
  NAND2_X1 U9946 ( .A1(n9106), .A2(n10165), .ZN(n7672) );
  INV_X1 U9947 ( .A(SI_6_), .ZN(n15288) );
  OR2_X1 U9948 ( .A1(n7735), .A2(n15288), .ZN(n7671) );
  OR2_X1 U9949 ( .A1(n7668), .A2(n8127), .ZN(n7669) );
  XNOR2_X1 U9950 ( .A(n7669), .B(P3_IR_REG_6__SCAN_IN), .ZN(n14914) );
  OR2_X1 U9951 ( .A1(n10754), .A2(n11424), .ZN(n7670) );
  INV_X1 U9952 ( .A(n15006), .ZN(n9778) );
  NAND2_X1 U9953 ( .A1(n12503), .A2(n9778), .ZN(n11827) );
  NAND2_X1 U9954 ( .A1(n8091), .A2(n11827), .ZN(n7689) );
  NAND2_X1 U9955 ( .A1(n7962), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7679) );
  AND2_X1 U9956 ( .A1(n7673), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7674) );
  OR2_X1 U9957 ( .A1(n7674), .A2(n7693), .ZN(n11831) );
  NAND2_X1 U9958 ( .A1(n7810), .A2(n11831), .ZN(n7678) );
  NAND2_X1 U9959 ( .A1(n8076), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7677) );
  INV_X1 U9960 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11400) );
  OR2_X1 U9961 ( .A1(n7675), .A2(n11400), .ZN(n7676) );
  NAND4_X1 U9962 ( .A1(n7679), .A2(n7678), .A3(n7677), .A4(n7676), .ZN(n15001)
         );
  NAND2_X1 U9963 ( .A1(n10171), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7682) );
  XNOR2_X1 U9964 ( .A(n7700), .B(n7699), .ZN(n10155) );
  NAND2_X1 U9965 ( .A1(n9106), .A2(n10155), .ZN(n7686) );
  NAND2_X1 U9966 ( .A1(n7668), .A2(n15392), .ZN(n7704) );
  NAND2_X1 U9967 ( .A1(n7704), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7684) );
  INV_X1 U9968 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7683) );
  XNOR2_X1 U9969 ( .A(n7684), .B(n7683), .ZN(n14927) );
  INV_X1 U9970 ( .A(n14927), .ZN(n11401) );
  OR2_X1 U9971 ( .A1(n10754), .A2(n11401), .ZN(n7685) );
  OAI211_X1 U9972 ( .C1(n7735), .C2(SI_7_), .A(n7686), .B(n7685), .ZN(n15097)
         );
  NAND2_X1 U9973 ( .A1(n15001), .A2(n15097), .ZN(n9164) );
  NAND2_X1 U9974 ( .A1(n11705), .A2(n9164), .ZN(n11828) );
  NAND2_X1 U9975 ( .A1(n12503), .A2(n15006), .ZN(n9161) );
  NAND2_X1 U9976 ( .A1(n9163), .A2(n9161), .ZN(n14999) );
  INV_X1 U9977 ( .A(n15002), .ZN(n11495) );
  NAND2_X1 U9978 ( .A1(n11495), .A2(n15020), .ZN(n11825) );
  NAND2_X1 U9979 ( .A1(n14999), .A2(n11825), .ZN(n7687) );
  NAND2_X1 U9980 ( .A1(n7687), .A2(n11827), .ZN(n7688) );
  INV_X1 U9981 ( .A(n15097), .ZN(n11835) );
  NAND2_X1 U9982 ( .A1(n15001), .A2(n11835), .ZN(n7690) );
  NAND2_X1 U9983 ( .A1(n7962), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7698) );
  NOR2_X1 U9984 ( .A1(n7693), .A2(n7692), .ZN(n7694) );
  OR2_X1 U9985 ( .A1(n7713), .A2(n7694), .ZN(n11715) );
  NAND2_X1 U9986 ( .A1(n7810), .A2(n11715), .ZN(n7697) );
  NAND2_X1 U9987 ( .A1(n6620), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7696) );
  INV_X1 U9988 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11436) );
  OR2_X1 U9989 ( .A1(n7675), .A2(n11436), .ZN(n7695) );
  NAND4_X1 U9990 ( .A1(n7698), .A2(n7697), .A3(n7696), .A4(n7695), .ZN(n11730)
         );
  INV_X1 U9991 ( .A(SI_8_), .ZN(n10153) );
  NAND2_X1 U9992 ( .A1(n10180), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7701) );
  XNOR2_X1 U9993 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n7720) );
  INV_X1 U9994 ( .A(n7720), .ZN(n7703) );
  XNOR2_X1 U9995 ( .A(n7721), .B(n7703), .ZN(n10152) );
  NAND2_X1 U9996 ( .A1(n9106), .A2(n10152), .ZN(n7710) );
  INV_X1 U9997 ( .A(n7740), .ZN(n7708) );
  NAND2_X1 U9998 ( .A1(n7705), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7706) );
  MUX2_X1 U9999 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7706), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n7707) );
  NAND2_X1 U10000 ( .A1(n7708), .A2(n7707), .ZN(n14942) );
  OR2_X1 U10001 ( .A1(n10754), .A2(n14942), .ZN(n7709) );
  OAI211_X1 U10002 ( .C1(n7735), .C2(n10153), .A(n7710), .B(n7709), .ZN(n11718) );
  AND2_X1 U10003 ( .A1(n11730), .A2(n11718), .ZN(n7712) );
  INV_X1 U10004 ( .A(n11730), .ZN(n11886) );
  INV_X1 U10005 ( .A(n11718), .ZN(n15104) );
  NAND2_X1 U10006 ( .A1(n11886), .A2(n15104), .ZN(n7711) );
  NAND2_X1 U10007 ( .A1(n7962), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7719) );
  OR2_X1 U10008 ( .A1(n7713), .A2(n11885), .ZN(n7714) );
  NAND2_X1 U10009 ( .A1(n7729), .A2(n7714), .ZN(n11889) );
  NAND2_X1 U10010 ( .A1(n7810), .A2(n11889), .ZN(n7718) );
  NAND2_X1 U10011 ( .A1(n8076), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7717) );
  INV_X1 U10012 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11409) );
  OR2_X1 U10013 ( .A1(n7675), .A2(n11409), .ZN(n7716) );
  NAND4_X1 U10014 ( .A1(n7719), .A2(n7718), .A3(n7717), .A4(n7716), .ZN(n12360) );
  NAND2_X1 U10015 ( .A1(n7722), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7723) );
  XNOR2_X1 U10016 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n7736) );
  XNOR2_X1 U10017 ( .A(n7737), .B(n7736), .ZN(n10148) );
  NAND2_X1 U10018 ( .A1(n9106), .A2(n10148), .ZN(n7727) );
  OR2_X1 U10019 ( .A1(n7735), .A2(SI_9_), .ZN(n7726) );
  OR2_X1 U10020 ( .A1(n7740), .A2(n8127), .ZN(n7724) );
  INV_X1 U10021 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7739) );
  XNOR2_X1 U10022 ( .A(n7724), .B(n7739), .ZN(n14963) );
  INV_X1 U10023 ( .A(n14963), .ZN(n11410) );
  OR2_X1 U10024 ( .A1(n10754), .A2(n11410), .ZN(n7725) );
  XNOR2_X1 U10025 ( .A(n12360), .B(n11888), .ZN(n11727) );
  NAND2_X1 U10026 ( .A1(n12360), .A2(n11888), .ZN(n7728) );
  NAND2_X1 U10027 ( .A1(n11726), .A2(n7728), .ZN(n11815) );
  NAND2_X1 U10028 ( .A1(n7962), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7734) );
  NAND2_X1 U10029 ( .A1(n7729), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7730) );
  NAND2_X1 U10030 ( .A1(n7745), .A2(n7730), .ZN(n12367) );
  NAND2_X1 U10031 ( .A1(n7810), .A2(n12367), .ZN(n7733) );
  NAND2_X1 U10032 ( .A1(n8076), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n7732) );
  INV_X1 U10033 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11440) );
  OR2_X1 U10034 ( .A1(n7675), .A2(n11440), .ZN(n7731) );
  NAND4_X1 U10035 ( .A1(n7734), .A2(n7733), .A3(n7732), .A4(n7731), .ZN(n12502) );
  XNOR2_X1 U10036 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n7752) );
  XNOR2_X1 U10037 ( .A(n7753), .B(n7752), .ZN(n10157) );
  NAND2_X1 U10038 ( .A1(n9106), .A2(n10157), .ZN(n7743) );
  NAND2_X1 U10039 ( .A1(n7740), .A2(n7739), .ZN(n7758) );
  NAND2_X1 U10040 ( .A1(n7758), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7741) );
  XNOR2_X1 U10041 ( .A(n7741), .B(P3_IR_REG_10__SCAN_IN), .ZN(n11441) );
  OR2_X1 U10042 ( .A1(n10754), .A2(n11441), .ZN(n7742) );
  OAI211_X1 U10043 ( .C1(n7735), .C2(SI_10_), .A(n7743), .B(n7742), .ZN(n11819) );
  OR2_X1 U10044 ( .A1(n12502), .A2(n11819), .ZN(n9174) );
  NAND2_X1 U10045 ( .A1(n12502), .A2(n11819), .ZN(n9172) );
  NAND2_X1 U10046 ( .A1(n9174), .A2(n9172), .ZN(n11814) );
  NAND2_X1 U10047 ( .A1(n11815), .A2(n11814), .ZN(n11813) );
  INV_X1 U10048 ( .A(n11819), .ZN(n12361) );
  NAND2_X1 U10049 ( .A1(n12502), .A2(n12361), .ZN(n7744) );
  NAND2_X1 U10050 ( .A1(n11813), .A2(n7744), .ZN(n11894) );
  NAND2_X1 U10051 ( .A1(n7962), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7751) );
  NAND2_X1 U10052 ( .A1(n7745), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7746) );
  NAND2_X1 U10053 ( .A1(n7767), .A2(n7746), .ZN(n12456) );
  NAND2_X1 U10054 ( .A1(n7810), .A2(n12456), .ZN(n7750) );
  NAND2_X1 U10055 ( .A1(n6620), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7749) );
  INV_X1 U10056 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n7747) );
  OR2_X1 U10057 ( .A1(n7675), .A2(n7747), .ZN(n7748) );
  NAND4_X1 U10058 ( .A1(n7751), .A2(n7750), .A3(n7749), .A4(n7748), .ZN(n14333) );
  INV_X1 U10059 ( .A(n14333), .ZN(n12450) );
  NAND2_X1 U10060 ( .A1(n7753), .A2(n7752), .ZN(n7756) );
  NAND2_X1 U10061 ( .A1(n7754), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7755) );
  XNOR2_X1 U10062 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n7757) );
  XNOR2_X1 U10063 ( .A(n7776), .B(n7757), .ZN(n10150) );
  NAND2_X1 U10064 ( .A1(n9106), .A2(n10150), .ZN(n7762) );
  OAI21_X1 U10065 ( .B1(n7758), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7760) );
  INV_X1 U10066 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7759) );
  XNOR2_X1 U10067 ( .A(n7760), .B(n7759), .ZN(n11528) );
  OR2_X1 U10068 ( .A1(n10754), .A2(n11521), .ZN(n7761) );
  NAND2_X1 U10069 ( .A1(n12450), .A2(n12925), .ZN(n7763) );
  NAND2_X1 U10070 ( .A1(n11894), .A2(n7763), .ZN(n7766) );
  INV_X1 U10071 ( .A(n12925), .ZN(n7764) );
  NAND2_X1 U10072 ( .A1(n14333), .A2(n7764), .ZN(n7765) );
  NAND2_X1 U10073 ( .A1(n7766), .A2(n7765), .ZN(n14332) );
  AND2_X1 U10074 ( .A1(n7767), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7768) );
  OR2_X1 U10075 ( .A1(n7768), .A2(n7789), .ZN(n14336) );
  NAND2_X1 U10076 ( .A1(n7810), .A2(n14336), .ZN(n7773) );
  NAND2_X1 U10077 ( .A1(n6620), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7772) );
  NAND2_X1 U10078 ( .A1(n7962), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7771) );
  INV_X1 U10079 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n7769) );
  OR2_X1 U10080 ( .A1(n7675), .A2(n7769), .ZN(n7770) );
  NAND4_X1 U10081 ( .A1(n7773), .A2(n7772), .A3(n7771), .A4(n7770), .ZN(n12455) );
  NAND2_X1 U10082 ( .A1(n10492), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7774) );
  NAND2_X1 U10083 ( .A1(n10622), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7796) );
  NAND2_X1 U10084 ( .A1(n10625), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7777) );
  NAND2_X1 U10085 ( .A1(n7796), .A2(n7777), .ZN(n7778) );
  NAND2_X1 U10086 ( .A1(n7779), .A2(n7778), .ZN(n7780) );
  AND2_X1 U10087 ( .A1(n7797), .A2(n7780), .ZN(n10167) );
  NAND2_X1 U10088 ( .A1(n9106), .A2(n10167), .ZN(n7784) );
  NAND2_X1 U10089 ( .A1(n7800), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7781) );
  XNOR2_X1 U10090 ( .A(n7781), .B(P3_IR_REG_12__SCAN_IN), .ZN(n11594) );
  OR2_X1 U10091 ( .A1(n10754), .A2(n11586), .ZN(n7783) );
  OR2_X1 U10092 ( .A1(n7735), .A2(n10169), .ZN(n7782) );
  NAND2_X1 U10093 ( .A1(n12455), .A2(n14339), .ZN(n9185) );
  NAND2_X1 U10094 ( .A1(n9186), .A2(n9185), .ZN(n8096) );
  NAND2_X1 U10095 ( .A1(n14332), .A2(n8096), .ZN(n7787) );
  INV_X1 U10096 ( .A(n14339), .ZN(n7785) );
  NAND2_X1 U10097 ( .A1(n12455), .A2(n7785), .ZN(n7786) );
  NAND2_X1 U10098 ( .A1(n7787), .A2(n7786), .ZN(n12811) );
  NAND2_X1 U10099 ( .A1(n6620), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7795) );
  NAND2_X1 U10100 ( .A1(n7789), .A2(n7788), .ZN(n7811) );
  OR2_X1 U10101 ( .A1(n7789), .A2(n7788), .ZN(n7790) );
  NAND2_X1 U10102 ( .A1(n7811), .A2(n7790), .ZN(n12816) );
  NAND2_X1 U10103 ( .A1(n7810), .A2(n12816), .ZN(n7794) );
  NAND2_X1 U10104 ( .A1(n7962), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7793) );
  INV_X1 U10105 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n7791) );
  OR2_X1 U10106 ( .A1(n7675), .A2(n7791), .ZN(n7792) );
  NAND4_X1 U10107 ( .A1(n7795), .A2(n7794), .A3(n7793), .A4(n7792), .ZN(n14334) );
  OAI21_X1 U10108 ( .B1(n6653), .B2(P1_DATAO_REG_13__SCAN_IN), .A(n7818), .ZN(
        n10300) );
  NAND2_X1 U10109 ( .A1(n10300), .A2(n9106), .ZN(n7807) );
  NAND2_X1 U10110 ( .A1(n7803), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7802) );
  MUX2_X1 U10111 ( .A(n7802), .B(P3_IR_REG_31__SCAN_IN), .S(n7801), .Z(n7804)
         );
  NAND2_X1 U10112 ( .A1(n7804), .A2(n7830), .ZN(n11845) );
  OAI22_X1 U10113 ( .A1(n7735), .A2(SI_13_), .B1(n11852), .B2(n10754), .ZN(
        n7805) );
  INV_X1 U10114 ( .A(n7805), .ZN(n7806) );
  OR2_X1 U10115 ( .A1(n14334), .A2(n12922), .ZN(n9189) );
  NAND2_X1 U10116 ( .A1(n14334), .A2(n12922), .ZN(n9188) );
  NAND2_X1 U10117 ( .A1(n9189), .A2(n9188), .ZN(n12812) );
  NAND2_X1 U10118 ( .A1(n12811), .A2(n12812), .ZN(n7809) );
  INV_X1 U10119 ( .A(n12922), .ZN(n11924) );
  NAND2_X1 U10120 ( .A1(n14334), .A2(n11924), .ZN(n7808) );
  NAND2_X1 U10121 ( .A1(n7809), .A2(n7808), .ZN(n12799) );
  NAND2_X1 U10122 ( .A1(n7962), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7816) );
  NAND2_X1 U10123 ( .A1(n7811), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7812) );
  NAND2_X1 U10124 ( .A1(n7837), .A2(n7812), .ZN(n12804) );
  NAND2_X1 U10125 ( .A1(n7810), .A2(n12804), .ZN(n7815) );
  NAND2_X1 U10126 ( .A1(n8076), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n7814) );
  INV_X1 U10127 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12874) );
  OR2_X1 U10128 ( .A1(n7675), .A2(n12874), .ZN(n7813) );
  NAND4_X1 U10129 ( .A1(n7816), .A2(n7815), .A3(n7814), .A4(n7813), .ZN(n12486) );
  XNOR2_X1 U10130 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n7819) );
  XNOR2_X1 U10131 ( .A(n7826), .B(n7819), .ZN(n10327) );
  NAND2_X1 U10132 ( .A1(n10327), .A2(n9106), .ZN(n7823) );
  NAND2_X1 U10133 ( .A1(n7830), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7820) );
  XNOR2_X1 U10134 ( .A(n7820), .B(P3_IR_REG_14__SCAN_IN), .ZN(n11848) );
  OAI22_X1 U10135 ( .A1(n7735), .A2(SI_14_), .B1(n11848), .B2(n10754), .ZN(
        n7821) );
  INV_X1 U10136 ( .A(n7821), .ZN(n7822) );
  OR2_X1 U10137 ( .A1(n12486), .A2(n12918), .ZN(n12785) );
  NAND2_X1 U10138 ( .A1(n12918), .A2(n12486), .ZN(n9194) );
  NAND2_X1 U10139 ( .A1(n12785), .A2(n9194), .ZN(n12800) );
  NAND2_X1 U10140 ( .A1(n12799), .A2(n12800), .ZN(n7825) );
  INV_X1 U10141 ( .A(n12918), .ZN(n11934) );
  NAND2_X1 U10142 ( .A1(n11934), .A2(n12486), .ZN(n7824) );
  NAND2_X1 U10143 ( .A1(n7825), .A2(n7824), .ZN(n12789) );
  NAND2_X1 U10144 ( .A1(n10806), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7827) );
  XNOR2_X1 U10145 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n7845) );
  INV_X1 U10146 ( .A(n7845), .ZN(n7829) );
  XNOR2_X1 U10147 ( .A(n7846), .B(n7829), .ZN(n10374) );
  NAND2_X1 U10148 ( .A1(n10374), .A2(n9106), .ZN(n7836) );
  NAND2_X1 U10149 ( .A1(n7851), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7833) );
  XNOR2_X1 U10150 ( .A(n7833), .B(n7850), .ZN(n12533) );
  OAI22_X1 U10151 ( .A1(n7735), .A2(n15227), .B1(n10754), .B2(n12533), .ZN(
        n7834) );
  INV_X1 U10152 ( .A(n7834), .ZN(n7835) );
  NAND2_X1 U10153 ( .A1(n7962), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7843) );
  INV_X1 U10154 ( .A(n7859), .ZN(n7839) );
  NAND2_X1 U10155 ( .A1(n7837), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7838) );
  NAND2_X1 U10156 ( .A1(n7839), .A2(n7838), .ZN(n12793) );
  NAND2_X1 U10157 ( .A1(n7810), .A2(n12793), .ZN(n7842) );
  NAND2_X1 U10158 ( .A1(n8076), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n7841) );
  INV_X1 U10159 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n15344) );
  OR2_X1 U10160 ( .A1(n7675), .A2(n15344), .ZN(n7840) );
  NAND4_X1 U10161 ( .A1(n7843), .A2(n7842), .A3(n7841), .A4(n7840), .ZN(n12501) );
  XNOR2_X1 U10162 ( .A(n12484), .B(n12802), .ZN(n12790) );
  NAND2_X1 U10163 ( .A1(n12484), .A2(n12501), .ZN(n7844) );
  NAND2_X1 U10164 ( .A1(n7846), .A2(n7845), .ZN(n7848) );
  NAND2_X1 U10165 ( .A1(n11016), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7847) );
  XNOR2_X1 U10166 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n7866) );
  INV_X1 U10167 ( .A(n7866), .ZN(n7849) );
  XNOR2_X1 U10168 ( .A(n7867), .B(n7849), .ZN(n10455) );
  NAND2_X1 U10169 ( .A1(n10455), .A2(n9106), .ZN(n7857) );
  NAND2_X1 U10170 ( .A1(n6748), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7852) );
  MUX2_X1 U10171 ( .A(n7852), .B(P3_IR_REG_31__SCAN_IN), .S(n7853), .Z(n7854)
         );
  NAND2_X1 U10172 ( .A1(n7854), .A2(n6744), .ZN(n12556) );
  OAI22_X1 U10173 ( .A1(n7735), .A2(n10456), .B1(n10754), .B2(n12556), .ZN(
        n7855) );
  INV_X1 U10174 ( .A(n7855), .ZN(n7856) );
  NAND2_X1 U10175 ( .A1(n7962), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7864) );
  INV_X1 U10176 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n7858) );
  NOR2_X1 U10177 ( .A1(n7859), .A2(n7858), .ZN(n7860) );
  OR2_X1 U10178 ( .A1(n7874), .A2(n7860), .ZN(n12780) );
  NAND2_X1 U10179 ( .A1(n7810), .A2(n12780), .ZN(n7863) );
  NAND2_X1 U10180 ( .A1(n6620), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n7862) );
  INV_X1 U10181 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12867) );
  OR2_X1 U10182 ( .A1(n7675), .A2(n12867), .ZN(n7861) );
  NAND4_X1 U10183 ( .A1(n7864), .A2(n7863), .A3(n7862), .A4(n7861), .ZN(n10685) );
  AND2_X1 U10184 ( .A1(n12779), .A2(n10685), .ZN(n7865) );
  NAND2_X1 U10185 ( .A1(n10840), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n7868) );
  XNOR2_X1 U10186 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .ZN(n7883) );
  INV_X1 U10187 ( .A(n7883), .ZN(n7869) );
  XNOR2_X1 U10188 ( .A(n7884), .B(n7869), .ZN(n10541) );
  NAND2_X1 U10189 ( .A1(n10541), .A2(n9106), .ZN(n7873) );
  INV_X1 U10190 ( .A(SI_17_), .ZN(n10543) );
  NAND2_X1 U10191 ( .A1(n6744), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7870) );
  XNOR2_X1 U10192 ( .A(n7870), .B(n7888), .ZN(n12575) );
  OAI22_X1 U10193 ( .A1(n7735), .A2(n10543), .B1(n10754), .B2(n12575), .ZN(
        n7871) );
  INV_X1 U10194 ( .A(n7871), .ZN(n7872) );
  NAND2_X1 U10195 ( .A1(n7962), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7879) );
  OR2_X1 U10196 ( .A1(n7874), .A2(n12418), .ZN(n7875) );
  NAND2_X1 U10197 ( .A1(n7894), .A2(n7875), .ZN(n12765) );
  NAND2_X1 U10198 ( .A1(n7810), .A2(n12765), .ZN(n7878) );
  NAND2_X1 U10199 ( .A1(n8076), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n7877) );
  INV_X1 U10200 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12578) );
  OR2_X1 U10201 ( .A1(n7675), .A2(n12578), .ZN(n7876) );
  NAND4_X1 U10202 ( .A1(n7879), .A2(n7878), .A3(n7877), .A4(n7876), .ZN(n12500) );
  OR2_X1 U10203 ( .A1(n12860), .A2(n12778), .ZN(n9207) );
  NAND2_X1 U10204 ( .A1(n12860), .A2(n12778), .ZN(n9206) );
  NAND2_X1 U10205 ( .A1(n12860), .A2(n12500), .ZN(n7882) );
  INV_X1 U10206 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10869) );
  NAND2_X1 U10207 ( .A1(n10869), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7885) );
  XNOR2_X1 U10208 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .ZN(n7902) );
  INV_X1 U10209 ( .A(n7902), .ZN(n7887) );
  XNOR2_X1 U10210 ( .A(n7903), .B(n7887), .ZN(n10593) );
  NAND2_X1 U10211 ( .A1(n10593), .A2(n9106), .ZN(n7893) );
  NAND2_X1 U10212 ( .A1(n6753), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7890) );
  XNOR2_X1 U10213 ( .A(n7890), .B(n7889), .ZN(n12600) );
  OAI22_X1 U10214 ( .A1(n7735), .A2(n10595), .B1(n10754), .B2(n12600), .ZN(
        n7891) );
  INV_X1 U10215 ( .A(n7891), .ZN(n7892) );
  NAND2_X1 U10216 ( .A1(n7962), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7899) );
  NAND2_X1 U10217 ( .A1(n7894), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7895) );
  NAND2_X1 U10218 ( .A1(n7909), .A2(n7895), .ZN(n12752) );
  NAND2_X1 U10219 ( .A1(n7810), .A2(n12752), .ZN(n7898) );
  NAND2_X1 U10220 ( .A1(n8076), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n7897) );
  INV_X1 U10221 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12858) );
  OR2_X1 U10222 ( .A1(n7675), .A2(n12858), .ZN(n7896) );
  NAND4_X1 U10223 ( .A1(n7899), .A2(n7898), .A3(n7897), .A4(n7896), .ZN(n12734) );
  NAND2_X1 U10224 ( .A1(n12751), .A2(n12758), .ZN(n9213) );
  OR2_X1 U10225 ( .A1(n12751), .A2(n12734), .ZN(n7901) );
  NAND2_X1 U10226 ( .A1(n7903), .A2(n7902), .ZN(n7904) );
  INV_X1 U10227 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11228) );
  AOI22_X1 U10228 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n11226), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n11228), .ZN(n7918) );
  XNOR2_X1 U10229 ( .A(n7917), .B(n7918), .ZN(n10597) );
  NAND2_X1 U10230 ( .A1(n10597), .A2(n9106), .ZN(n7908) );
  OAI22_X1 U10231 ( .A1(n7735), .A2(SI_19_), .B1(n12595), .B2(n10754), .ZN(
        n7906) );
  INV_X1 U10232 ( .A(n7906), .ZN(n7907) );
  NAND2_X1 U10233 ( .A1(n7962), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n7914) );
  AND2_X1 U10234 ( .A1(n7909), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n7910) );
  OR2_X1 U10235 ( .A1(n7910), .A2(n7924), .ZN(n12737) );
  NAND2_X1 U10236 ( .A1(n6627), .A2(n12737), .ZN(n7913) );
  NAND2_X1 U10237 ( .A1(n6620), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n7912) );
  INV_X1 U10238 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12854) );
  OR2_X1 U10239 ( .A1(n7675), .A2(n12854), .ZN(n7911) );
  NAND4_X1 U10240 ( .A1(n7914), .A2(n7913), .A3(n7912), .A4(n7911), .ZN(n12721) );
  NAND2_X1 U10241 ( .A1(n12901), .A2(n12721), .ZN(n9219) );
  INV_X1 U10242 ( .A(n12901), .ZN(n7915) );
  NAND2_X1 U10243 ( .A1(n7915), .A2(n12721), .ZN(n7916) );
  NAND2_X1 U10244 ( .A1(n7918), .A2(n7917), .ZN(n7919) );
  XNOR2_X1 U10245 ( .A(n7933), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n10872) );
  NAND2_X1 U10246 ( .A1(n10872), .A2(n9106), .ZN(n7922) );
  NAND2_X1 U10247 ( .A1(n7962), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n7930) );
  INV_X1 U10248 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n7923) );
  NOR2_X1 U10249 ( .A1(n7924), .A2(n7923), .ZN(n7925) );
  OR2_X1 U10250 ( .A1(n7939), .A2(n7925), .ZN(n12725) );
  NAND2_X1 U10251 ( .A1(n7810), .A2(n12725), .ZN(n7929) );
  NAND2_X1 U10252 ( .A1(n6620), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n7928) );
  INV_X1 U10253 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n7926) );
  OR2_X1 U10254 ( .A1(n7675), .A2(n7926), .ZN(n7927) );
  NAND4_X1 U10255 ( .A1(n7930), .A2(n7929), .A3(n7928), .A4(n7927), .ZN(n12733) );
  XNOR2_X1 U10256 ( .A(n12848), .B(n12710), .ZN(n12719) );
  NAND2_X1 U10257 ( .A1(n12848), .A2(n12733), .ZN(n7931) );
  NAND2_X1 U10258 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n7932), .ZN(n7935) );
  INV_X1 U10259 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11282) );
  AOI22_X1 U10260 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n11285), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n11282), .ZN(n7946) );
  XNOR2_X1 U10261 ( .A(n7945), .B(n7078), .ZN(n10979) );
  NAND2_X1 U10262 ( .A1(n10979), .A2(n9106), .ZN(n7937) );
  INV_X1 U10263 ( .A(SI_21_), .ZN(n10981) );
  NAND2_X1 U10264 ( .A1(n7962), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n7944) );
  INV_X1 U10265 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n7938) );
  OR2_X1 U10266 ( .A1(n7939), .A2(n7938), .ZN(n7940) );
  NAND2_X1 U10267 ( .A1(n7950), .A2(n7940), .ZN(n12712) );
  NAND2_X1 U10268 ( .A1(n7810), .A2(n12712), .ZN(n7943) );
  NAND2_X1 U10269 ( .A1(n8076), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n7942) );
  INV_X1 U10270 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12845) );
  OR2_X1 U10271 ( .A1(n7675), .A2(n12845), .ZN(n7941) );
  NAND4_X1 U10272 ( .A1(n7944), .A2(n7943), .A3(n7942), .A4(n7941), .ZN(n12722) );
  OR2_X1 U10273 ( .A1(n12383), .A2(n12722), .ZN(n9225) );
  NAND2_X1 U10274 ( .A1(n12383), .A2(n12722), .ZN(n9224) );
  INV_X1 U10275 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10398) );
  AOI22_X1 U10276 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(
        P2_DATAO_REG_22__SCAN_IN), .B1(n10398), .B2(n15235), .ZN(n7957) );
  XNOR2_X1 U10277 ( .A(n7956), .B(n7957), .ZN(n11055) );
  NAND2_X1 U10278 ( .A1(n11055), .A2(n9106), .ZN(n7949) );
  INV_X1 U10279 ( .A(SI_22_), .ZN(n7947) );
  NAND2_X1 U10280 ( .A1(n7962), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n7955) );
  NAND2_X1 U10281 ( .A1(n7950), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n7951) );
  NAND2_X1 U10282 ( .A1(n7960), .A2(n7951), .ZN(n12701) );
  NAND2_X1 U10283 ( .A1(n6627), .A2(n12701), .ZN(n7954) );
  NAND2_X1 U10284 ( .A1(n8076), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n7953) );
  INV_X1 U10285 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12841) );
  OR2_X1 U10286 ( .A1(n7675), .A2(n12841), .ZN(n7952) );
  NAND4_X1 U10287 ( .A1(n7955), .A2(n7954), .A3(n7953), .A4(n7952), .ZN(n12681) );
  INV_X1 U10288 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11772) );
  INV_X1 U10289 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11777) );
  AOI22_X1 U10290 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(
        P1_DATAO_REG_23__SCAN_IN), .B1(n11772), .B2(n11777), .ZN(n7969) );
  XNOR2_X1 U10291 ( .A(n7970), .B(n7969), .ZN(n11203) );
  NAND2_X1 U10292 ( .A1(n11203), .A2(n9106), .ZN(n7959) );
  AND2_X1 U10293 ( .A1(n7960), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7961) );
  OR2_X1 U10294 ( .A1(n7961), .A2(n7976), .ZN(n12685) );
  NAND2_X1 U10295 ( .A1(n12685), .A2(n7810), .ZN(n7967) );
  NAND2_X1 U10296 ( .A1(n7962), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n7964) );
  INV_X1 U10297 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n15364) );
  OR2_X1 U10298 ( .A1(n7675), .A2(n15364), .ZN(n7963) );
  AND2_X1 U10299 ( .A1(n7964), .A2(n7963), .ZN(n7966) );
  NAND2_X1 U10300 ( .A1(n6620), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n7965) );
  XNOR2_X1 U10301 ( .A(n12689), .B(n12699), .ZN(n12680) );
  NAND2_X1 U10302 ( .A1(n12689), .A2(n12668), .ZN(n7968) );
  NOR2_X1 U10303 ( .A1(n7970), .A2(n7969), .ZN(n7972) );
  XNOR2_X1 U10304 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n7982), .ZN(n11659) );
  NAND2_X1 U10305 ( .A1(n11659), .A2(n9106), .ZN(n7974) );
  INV_X1 U10306 ( .A(SI_24_), .ZN(n11661) );
  INV_X1 U10307 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n7981) );
  INV_X1 U10308 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n7975) );
  NAND2_X1 U10309 ( .A1(n7976), .A2(n7975), .ZN(n8003) );
  INV_X1 U10310 ( .A(n7976), .ZN(n7977) );
  NAND2_X1 U10311 ( .A1(n7977), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n7978) );
  NAND2_X1 U10312 ( .A1(n8003), .A2(n7978), .ZN(n12673) );
  NAND2_X1 U10313 ( .A1(n12673), .A2(n6627), .ZN(n7980) );
  AOI22_X1 U10314 ( .A1(n6620), .A2(P3_REG0_REG_24__SCAN_IN), .B1(n7962), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n7979) );
  OAI211_X1 U10315 ( .C1(n7675), .C2(n7981), .A(n7980), .B(n7979), .ZN(n12682)
         );
  NAND2_X1 U10316 ( .A1(n12675), .A2(n12682), .ZN(n9240) );
  INV_X1 U10317 ( .A(n12682), .ZN(n12405) );
  NAND2_X1 U10318 ( .A1(n12831), .A2(n12405), .ZN(n9242) );
  NAND2_X1 U10319 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n7983), .ZN(n7984) );
  INV_X1 U10320 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13503) );
  NAND2_X1 U10321 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n13503), .ZN(n7985) );
  INV_X1 U10322 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14157) );
  INV_X1 U10323 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14154) );
  AOI22_X1 U10324 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n13499), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n14154), .ZN(n7986) );
  XNOR2_X1 U10325 ( .A(n8021), .B(n7986), .ZN(n11940) );
  NAND2_X1 U10326 ( .A1(n11940), .A2(n9106), .ZN(n7989) );
  INV_X1 U10327 ( .A(SI_26_), .ZN(n11941) );
  INV_X1 U10328 ( .A(n8003), .ZN(n7991) );
  INV_X1 U10329 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n7990) );
  NAND2_X1 U10330 ( .A1(n7991), .A2(n7990), .ZN(n8005) );
  NAND2_X1 U10331 ( .A1(n8005), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n7992) );
  NAND2_X1 U10332 ( .A1(n8028), .A2(n7992), .ZN(n12645) );
  NAND2_X1 U10333 ( .A1(n12645), .A2(n6627), .ZN(n7997) );
  INV_X1 U10334 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n8943) );
  NAND2_X1 U10335 ( .A1(n7962), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n7994) );
  NAND2_X1 U10336 ( .A1(n8046), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n7993) );
  OAI211_X1 U10337 ( .C1(n8943), .C2(n7715), .A(n7994), .B(n7993), .ZN(n7995)
         );
  INV_X1 U10338 ( .A(n7995), .ZN(n7996) );
  OR2_X1 U10339 ( .A1(n9838), .A2(n12656), .ZN(n8012) );
  INV_X1 U10340 ( .A(n8012), .ZN(n8011) );
  AOI22_X1 U10341 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n14157), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n13503), .ZN(n7998) );
  INV_X1 U10342 ( .A(n7998), .ZN(n7999) );
  XNOR2_X1 U10343 ( .A(n8000), .B(n7999), .ZN(n11737) );
  NAND2_X1 U10344 ( .A1(n11737), .A2(n9106), .ZN(n8002) );
  INV_X1 U10345 ( .A(SI_25_), .ZN(n11738) );
  OR2_X1 U10346 ( .A1(n7735), .A2(n11738), .ZN(n8001) );
  NAND2_X2 U10347 ( .A1(n8002), .A2(n8001), .ZN(n12396) );
  NAND2_X1 U10348 ( .A1(n8003), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8004) );
  NAND2_X1 U10349 ( .A1(n8005), .A2(n8004), .ZN(n12659) );
  NAND2_X1 U10350 ( .A1(n12659), .A2(n7810), .ZN(n8008) );
  AOI22_X1 U10351 ( .A1(n8046), .A2(P3_REG1_REG_25__SCAN_IN), .B1(n8076), .B2(
        P3_REG0_REG_25__SCAN_IN), .ZN(n8007) );
  NAND2_X1 U10352 ( .A1(n7962), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8006) );
  INV_X1 U10353 ( .A(n12671), .ZN(n12475) );
  NAND2_X1 U10354 ( .A1(n12396), .A2(n12475), .ZN(n8936) );
  NAND2_X1 U10355 ( .A1(n9838), .A2(n12656), .ZN(n8009) );
  AND2_X1 U10356 ( .A1(n8936), .A2(n8009), .ZN(n8010) );
  OR2_X2 U10357 ( .A1(n8011), .A2(n8010), .ZN(n8017) );
  INV_X1 U10358 ( .A(n8017), .ZN(n8014) );
  AND2_X1 U10359 ( .A1(n12654), .A2(n8012), .ZN(n8013) );
  AND2_X1 U10360 ( .A1(n12667), .A2(n8016), .ZN(n8015) );
  INV_X1 U10361 ( .A(n8016), .ZN(n8019) );
  NAND2_X1 U10362 ( .A1(n12831), .A2(n12682), .ZN(n8935) );
  AND2_X1 U10363 ( .A1(n8935), .A2(n8017), .ZN(n8018) );
  NOR2_X1 U10364 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n14154), .ZN(n8022) );
  OAI22_X1 U10365 ( .A1(n8022), .A2(n8021), .B1(P2_DATAO_REG_26__SCAN_IN), 
        .B2(n13499), .ZN(n8038) );
  INV_X1 U10366 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13495) );
  AOI22_X1 U10367 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n13495), .B2(n15324), .ZN(n8023) );
  XNOR2_X1 U10368 ( .A(n8038), .B(n8023), .ZN(n12943) );
  NAND2_X1 U10369 ( .A1(n12943), .A2(n9106), .ZN(n8025) );
  INV_X1 U10370 ( .A(SI_27_), .ZN(n12945) );
  INV_X1 U10371 ( .A(n8028), .ZN(n8027) );
  INV_X1 U10372 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8026) );
  NAND2_X1 U10373 ( .A1(n8027), .A2(n8026), .ZN(n8044) );
  NAND2_X1 U10374 ( .A1(n8028), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8029) );
  NAND2_X1 U10375 ( .A1(n8044), .A2(n8029), .ZN(n12637) );
  NAND2_X1 U10376 ( .A1(n12637), .A2(n7810), .ZN(n8034) );
  INV_X1 U10377 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n8956) );
  NAND2_X1 U10378 ( .A1(n7962), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8031) );
  NAND2_X1 U10379 ( .A1(n6620), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8030) );
  OAI211_X1 U10380 ( .C1(n7675), .C2(n8956), .A(n8031), .B(n8030), .ZN(n8032)
         );
  INV_X1 U10381 ( .A(n8032), .ZN(n8033) );
  NAND2_X1 U10382 ( .A1(n9842), .A2(n12477), .ZN(n8961) );
  OR2_X1 U10383 ( .A1(n9842), .A2(n12477), .ZN(n8035) );
  OR2_X1 U10384 ( .A1(n9842), .A2(n12499), .ZN(n8037) );
  NAND2_X1 U10385 ( .A1(n8949), .A2(n8037), .ZN(n8964) );
  NAND2_X1 U10386 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n13495), .ZN(n8039) );
  INV_X1 U10387 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14148) );
  AOI22_X1 U10388 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(
        P2_DATAO_REG_28__SCAN_IN), .B1(n14148), .B2(n13490), .ZN(n8040) );
  INV_X1 U10389 ( .A(n8040), .ZN(n8041) );
  XNOR2_X1 U10390 ( .A(n8052), .B(n8041), .ZN(n12940) );
  NAND2_X1 U10391 ( .A1(n12940), .A2(n9106), .ZN(n8043) );
  INV_X1 U10392 ( .A(SI_28_), .ZN(n12942) );
  NAND2_X1 U10393 ( .A1(n8044), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8045) );
  NAND2_X1 U10394 ( .A1(n8056), .A2(n8045), .ZN(n12627) );
  INV_X1 U10395 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U10396 ( .A1(n7962), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8048) );
  NAND2_X1 U10397 ( .A1(n8046), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8047) );
  OAI211_X1 U10398 ( .C1(n8049), .C2(n7715), .A(n8048), .B(n8047), .ZN(n8050)
         );
  NAND2_X1 U10399 ( .A1(n12631), .A2(n9868), .ZN(n8109) );
  INV_X1 U10400 ( .A(n9868), .ZN(n12498) );
  OR2_X2 U10401 ( .A1(n8967), .A2(n8051), .ZN(n8062) );
  NOR2_X1 U10402 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n14148), .ZN(n8053) );
  INV_X1 U10403 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13487) );
  OAI22_X1 U10404 ( .A1(n14144), .A2(n13487), .B1(P1_DATAO_REG_29__SCAN_IN), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9099) );
  XNOR2_X1 U10405 ( .A(n9098), .B(n7117), .ZN(n12936) );
  NAND2_X1 U10406 ( .A1(n12936), .A2(n9106), .ZN(n8055) );
  INV_X1 U10407 ( .A(SI_29_), .ZN(n12939) );
  NAND2_X1 U10408 ( .A1(n12611), .A2(n7810), .ZN(n9112) );
  INV_X1 U10409 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8174) );
  NAND2_X1 U10410 ( .A1(n6620), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8058) );
  NAND2_X1 U10411 ( .A1(n7962), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8057) );
  OAI211_X1 U10412 ( .C1(n8174), .C2(n7675), .A(n8058), .B(n8057), .ZN(n8059)
         );
  INV_X1 U10413 ( .A(n8059), .ZN(n8060) );
  NAND2_X1 U10414 ( .A1(n9112), .A2(n8060), .ZN(n12497) );
  XNOR2_X1 U10415 ( .A(n9118), .B(n12497), .ZN(n9291) );
  NAND2_X1 U10416 ( .A1(n8063), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8065) );
  NAND2_X1 U10417 ( .A1(n12595), .A2(n9301), .ZN(n8146) );
  NAND2_X1 U10418 ( .A1(n6673), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8066) );
  MUX2_X1 U10419 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8066), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8067) );
  INV_X1 U10420 ( .A(n8067), .ZN(n8070) );
  NOR2_X1 U10421 ( .A1(n8070), .A2(n8069), .ZN(n8166) );
  INV_X1 U10422 ( .A(n8069), .ZN(n8071) );
  NAND2_X1 U10423 ( .A1(n8071), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8073) );
  NAND2_X1 U10424 ( .A1(n8166), .A2(n11451), .ZN(n9126) );
  INV_X2 U10425 ( .A(n11420), .ZN(n11415) );
  OR2_X1 U10426 ( .A1(n6628), .A2(n11415), .ZN(n10768) );
  INV_X1 U10427 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14349) );
  NAND2_X1 U10428 ( .A1(n7962), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8078) );
  NAND2_X1 U10429 ( .A1(n6620), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8077) );
  OAI211_X1 U10430 ( .C1(n7675), .C2(n14349), .A(n8078), .B(n8077), .ZN(n8079)
         );
  INV_X1 U10431 ( .A(n8079), .ZN(n8080) );
  NAND2_X1 U10432 ( .A1(n10754), .A2(n10768), .ZN(n8081) );
  INV_X1 U10433 ( .A(P3_B_REG_SCAN_IN), .ZN(n8082) );
  OR2_X1 U10434 ( .A1(n6628), .A2(n8082), .ZN(n8083) );
  NAND2_X1 U10435 ( .A1(n15059), .A2(n8083), .ZN(n12612) );
  NOR2_X1 U10436 ( .A1(n11014), .A2(n12612), .ZN(n8084) );
  OAI21_X2 U10437 ( .B1(n8087), .B2(n15016), .A(n8086), .ZN(n12624) );
  INV_X1 U10438 ( .A(n11888), .ZN(n9786) );
  OR2_X1 U10439 ( .A1(n12360), .A2(n9786), .ZN(n11809) );
  AND2_X1 U10440 ( .A1(n11809), .A2(n9174), .ZN(n8088) );
  NAND2_X1 U10441 ( .A1(n12360), .A2(n9786), .ZN(n9173) );
  OR2_X1 U10442 ( .A1(n11730), .A2(n15104), .ZN(n9169) );
  NAND2_X1 U10443 ( .A1(n11730), .A2(n15104), .ZN(n9168) );
  AND2_X1 U10444 ( .A1(n8088), .A2(n11807), .ZN(n8095) );
  INV_X1 U10445 ( .A(n11947), .ZN(n11954) );
  NAND2_X1 U10446 ( .A1(n9131), .A2(n9138), .ZN(n9770) );
  NAND2_X1 U10447 ( .A1(n9770), .A2(n9140), .ZN(n15039) );
  INV_X1 U10448 ( .A(n15041), .ZN(n9133) );
  NAND2_X1 U10449 ( .A1(n15039), .A2(n9133), .ZN(n15038) );
  OR2_X1 U10450 ( .A1(n15060), .A2(n15050), .ZN(n9136) );
  NAND2_X1 U10451 ( .A1(n15025), .A2(n9278), .ZN(n8089) );
  NAND2_X1 U10452 ( .A1(n8089), .A2(n9145), .ZN(n11449) );
  INV_X1 U10453 ( .A(n11452), .ZN(n11450) );
  NAND2_X1 U10454 ( .A1(n11449), .A2(n11450), .ZN(n8090) );
  NAND2_X1 U10455 ( .A1(n15012), .A2(n15014), .ZN(n15011) );
  INV_X1 U10456 ( .A(n14999), .ZN(n9279) );
  NAND2_X1 U10457 ( .A1(n14996), .A2(n9279), .ZN(n8092) );
  NAND2_X1 U10458 ( .A1(n8092), .A2(n9163), .ZN(n11704) );
  AND2_X1 U10459 ( .A1(n11834), .A2(n7014), .ZN(n11706) );
  AND2_X1 U10460 ( .A1(n11706), .A2(n9173), .ZN(n8093) );
  NAND2_X1 U10461 ( .A1(n11704), .A2(n8093), .ZN(n11808) );
  INV_X1 U10462 ( .A(n9172), .ZN(n8094) );
  OR2_X1 U10463 ( .A1(n14333), .A2(n12925), .ZN(n9178) );
  NAND2_X1 U10464 ( .A1(n14333), .A2(n12925), .ZN(n9179) );
  NAND2_X1 U10465 ( .A1(n9178), .A2(n9179), .ZN(n11893) );
  INV_X1 U10466 ( .A(n11893), .ZN(n11897) );
  NAND2_X1 U10467 ( .A1(n8097), .A2(n9186), .ZN(n12810) );
  NAND2_X1 U10468 ( .A1(n12484), .A2(n12802), .ZN(n9201) );
  AND2_X1 U10469 ( .A1(n12785), .A2(n9201), .ZN(n8099) );
  INV_X1 U10470 ( .A(n9201), .ZN(n8098) );
  INV_X1 U10471 ( .A(n12790), .ZN(n12787) );
  OR2_X1 U10472 ( .A1(n12779), .A2(n12792), .ZN(n9203) );
  NAND2_X1 U10473 ( .A1(n12779), .A2(n12792), .ZN(n9202) );
  NAND2_X1 U10474 ( .A1(n12774), .A2(n12776), .ZN(n12773) );
  NAND2_X1 U10475 ( .A1(n12773), .A2(n9202), .ZN(n12764) );
  NAND2_X1 U10476 ( .A1(n12764), .A2(n12763), .ZN(n12762) );
  INV_X1 U10477 ( .A(n12744), .ZN(n8100) );
  INV_X1 U10478 ( .A(n12848), .ZN(n12727) );
  NAND2_X1 U10479 ( .A1(n12727), .A2(n12733), .ZN(n9222) );
  NAND2_X1 U10480 ( .A1(n12383), .A2(n12700), .ZN(n8103) );
  NAND2_X1 U10481 ( .A1(n12447), .A2(n12711), .ZN(n9228) );
  NAND2_X1 U10482 ( .A1(n12695), .A2(n9228), .ZN(n8104) );
  NAND2_X1 U10483 ( .A1(n8104), .A2(n9229), .ZN(n12691) );
  INV_X1 U10484 ( .A(n12680), .ZN(n12690) );
  INV_X1 U10485 ( .A(n12689), .ZN(n12838) );
  NAND2_X1 U10486 ( .A1(n12838), .A2(n12668), .ZN(n9239) );
  NAND2_X1 U10487 ( .A1(n12396), .A2(n12671), .ZN(n9246) );
  NAND2_X1 U10488 ( .A1(n8106), .A2(n9246), .ZN(n8934) );
  INV_X1 U10489 ( .A(n12656), .ZN(n8107) );
  NAND2_X1 U10490 ( .A1(n8934), .A2(n9253), .ZN(n8108) );
  NAND2_X1 U10491 ( .A1(n9838), .A2(n8107), .ZN(n9252) );
  AND2_X1 U10492 ( .A1(n8109), .A2(n8961), .ZN(n9261) );
  XNOR2_X1 U10493 ( .A(n9097), .B(n9291), .ZN(n12619) );
  NAND2_X1 U10494 ( .A1(n9301), .A2(n10875), .ZN(n8110) );
  NAND2_X1 U10495 ( .A1(n12595), .A2(n8110), .ZN(n8111) );
  NAND2_X1 U10496 ( .A1(n8111), .A2(n10980), .ZN(n8113) );
  OAI21_X1 U10497 ( .B1(n8166), .B2(n11451), .A(n11053), .ZN(n8112) );
  NAND2_X1 U10498 ( .A1(n8113), .A2(n8112), .ZN(n9859) );
  NAND2_X1 U10499 ( .A1(n9859), .A2(n15103), .ZN(n11057) );
  INV_X1 U10500 ( .A(n12595), .ZN(n12607) );
  NAND2_X1 U10501 ( .A1(n12607), .A2(n10875), .ZN(n9272) );
  OR2_X1 U10502 ( .A1(n11057), .A2(n9272), .ZN(n8114) );
  OR3_X1 U10503 ( .A1(n12595), .A2(n11053), .A3(n10875), .ZN(n8165) );
  NOR2_X1 U10504 ( .A1(n12624), .A2(n8115), .ZN(n8173) );
  INV_X1 U10505 ( .A(n8116), .ZN(n8120) );
  NAND2_X1 U10506 ( .A1(n8120), .A2(n8119), .ZN(n11662) );
  XNOR2_X1 U10507 ( .A(n11662), .B(P3_B_REG_SCAN_IN), .ZN(n8126) );
  INV_X1 U10508 ( .A(n8121), .ZN(n8125) );
  NOR2_X1 U10509 ( .A1(n8116), .A2(n8127), .ZN(n8123) );
  NOR2_X1 U10510 ( .A1(n8121), .A2(n8127), .ZN(n8131) );
  INV_X1 U10511 ( .A(n8132), .ZN(n11944) );
  OAI22_X1 U10512 ( .A1(n8134), .A2(P3_D_REG_1__SCAN_IN), .B1(n8132), .B2(
        n6850), .ZN(n11063) );
  NAND2_X1 U10513 ( .A1(n11944), .A2(n11662), .ZN(n8133) );
  INV_X1 U10514 ( .A(n8164), .ZN(n8145) );
  NOR4_X1 U10515 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_24__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n8143) );
  INV_X1 U10516 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n15265) );
  INV_X1 U10517 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10645) );
  INV_X1 U10518 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n15268) );
  INV_X1 U10519 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10641) );
  NAND4_X1 U10520 ( .A1(n15265), .A2(n10645), .A3(n15268), .A4(n10641), .ZN(
        n8140) );
  NOR4_X1 U10521 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_9__SCAN_IN), .ZN(n8138) );
  NOR4_X1 U10522 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n8137) );
  NOR4_X1 U10523 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_6__SCAN_IN), .A3(
        P3_D_REG_3__SCAN_IN), .A4(P3_D_REG_5__SCAN_IN), .ZN(n8136) );
  NOR4_X1 U10524 ( .A1(P3_D_REG_16__SCAN_IN), .A2(P3_D_REG_15__SCAN_IN), .A3(
        P3_D_REG_30__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n8135) );
  NAND4_X1 U10525 ( .A1(n8138), .A2(n8137), .A3(n8136), .A4(n8135), .ZN(n8139)
         );
  NOR4_X1 U10526 ( .A1(P3_D_REG_4__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        n8140), .A4(n8139), .ZN(n8142) );
  NOR4_X1 U10527 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_17__SCAN_IN), .A3(
        P3_D_REG_22__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n8141) );
  NAND3_X1 U10528 ( .A1(n8143), .A2(n8142), .A3(n8141), .ZN(n8144) );
  NAND2_X1 U10529 ( .A1(n10399), .A2(n8144), .ZN(n8162) );
  NAND2_X1 U10530 ( .A1(n8145), .A2(n8162), .ZN(n9858) );
  NAND2_X1 U10531 ( .A1(n8166), .A2(n10980), .ZN(n9764) );
  OR2_X1 U10532 ( .A1(n8146), .A2(n9764), .ZN(n9855) );
  OR2_X1 U10533 ( .A1(n9272), .A2(n9854), .ZN(n8147) );
  AND2_X1 U10534 ( .A1(n9855), .A2(n8147), .ZN(n8149) );
  INV_X1 U10535 ( .A(n9859), .ZN(n8148) );
  NAND3_X1 U10536 ( .A1(n11063), .A2(n11939), .A3(n8162), .ZN(n9864) );
  OAI22_X1 U10537 ( .A1(n9858), .A2(n8149), .B1(n8148), .B2(n9864), .ZN(n8155)
         );
  INV_X1 U10538 ( .A(n11662), .ZN(n8150) );
  NAND2_X1 U10539 ( .A1(n6850), .A2(n8150), .ZN(n8151) );
  INV_X1 U10540 ( .A(n8152), .ZN(n8153) );
  NAND2_X1 U10541 ( .A1(n8153), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8154) );
  OR2_X1 U10542 ( .A1(n8173), .A2(n8156), .ZN(n8161) );
  INV_X1 U10543 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8157) );
  NOR2_X1 U10544 ( .A1(n15119), .A2(n8157), .ZN(n8159) );
  NOR2_X1 U10545 ( .A1(n8159), .A2(n8158), .ZN(n8160) );
  NAND2_X1 U10546 ( .A1(n8161), .A2(n8160), .ZN(P3_U3456) );
  AND2_X1 U10547 ( .A1(n8162), .A2(n10749), .ZN(n8163) );
  NAND2_X1 U10548 ( .A1(n9272), .A2(n10752), .ZN(n11059) );
  NAND2_X1 U10549 ( .A1(n8165), .A2(n9854), .ZN(n11061) );
  NAND2_X1 U10550 ( .A1(n11059), .A2(n11061), .ZN(n8171) );
  OAI22_X1 U10551 ( .A1(n12595), .A2(n11053), .B1(n8166), .B2(n15103), .ZN(
        n8167) );
  NAND2_X1 U10552 ( .A1(n8167), .A2(n9272), .ZN(n8168) );
  NAND2_X1 U10553 ( .A1(n8168), .A2(n9854), .ZN(n8169) );
  OR2_X1 U10554 ( .A1(n11939), .A2(n8169), .ZN(n8170) );
  OAI21_X1 U10555 ( .B1(n11063), .B2(n8171), .A(n8170), .ZN(n8172) );
  OR2_X1 U10556 ( .A1(n8173), .A2(n15130), .ZN(n8178) );
  NOR2_X1 U10557 ( .A1(n15132), .A2(n8174), .ZN(n8176) );
  NOR2_X1 U10558 ( .A1(n12622), .A2(n12882), .ZN(n8175) );
  NOR2_X1 U10559 ( .A1(n8176), .A2(n8175), .ZN(n8177) );
  NAND2_X1 U10560 ( .A1(n8178), .A2(n8177), .ZN(P3_U3488) );
  NAND4_X1 U10561 ( .A1(n8199), .A2(n8181), .A3(n8180), .A4(n8179), .ZN(n8182)
         );
  INV_X2 U10562 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n15356) );
  NOR2_X4 U10563 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8218) );
  NOR2_X1 U10564 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n8188) );
  INV_X1 U10565 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8192) );
  NAND2_X1 U10566 ( .A1(n8213), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8195) );
  INV_X1 U10567 ( .A(n12203), .ZN(n8196) );
  INV_X1 U10568 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8197) );
  INV_X1 U10569 ( .A(n8202), .ZN(n8203) );
  INV_X1 U10570 ( .A(n8204), .ZN(n8205) );
  NOR2_X1 U10571 ( .A1(n8559), .A2(n8205), .ZN(n8206) );
  NAND2_X1 U10572 ( .A1(n8358), .A2(n8206), .ZN(n8629) );
  XNOR2_X1 U10573 ( .A(n8207), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8912) );
  NOR2_X1 U10574 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n8211) );
  NOR2_X1 U10575 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .ZN(n8210) );
  NOR2_X1 U10576 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .ZN(n8209) );
  NAND4_X1 U10577 ( .A1(n8211), .A2(n8210), .A3(n8209), .A4(n8208), .ZN(n8212)
         );
  OR2_X1 U10578 ( .A1(n8218), .A2(n13478), .ZN(n8219) );
  XNOR2_X1 U10579 ( .A(n8219), .B(P2_IR_REG_2__SCAN_IN), .ZN(n10242) );
  OAI21_X1 U10580 ( .B1(n8226), .B2(P1_DATAO_REG_0__SCAN_IN), .A(n8223), .ZN(
        n8224) );
  NOR2_X1 U10581 ( .A1(n8224), .A2(n10132), .ZN(n8248) );
  NAND2_X1 U10582 ( .A1(n8227), .A2(SI_2_), .ZN(n8277) );
  OAI21_X1 U10583 ( .B1(SI_2_), .B2(n8227), .A(n8277), .ZN(n8229) );
  NAND2_X1 U10584 ( .A1(n8228), .A2(n8229), .ZN(n8232) );
  INV_X1 U10585 ( .A(n8229), .ZN(n8230) );
  NAND2_X1 U10586 ( .A1(n8231), .A2(n8230), .ZN(n8278) );
  NAND2_X1 U10587 ( .A1(n8232), .A2(n8278), .ZN(n10127) );
  NAND2_X1 U10588 ( .A1(n8235), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8237) );
  AND2_X2 U10589 ( .A1(n13484), .A2(n13488), .ZN(n8313) );
  NAND2_X1 U10590 ( .A1(n8313), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8242) );
  AND2_X2 U10591 ( .A1(n8238), .A2(n13488), .ZN(n8289) );
  NAND2_X1 U10592 ( .A1(n8289), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8241) );
  NAND2_X1 U10593 ( .A1(n8288), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8240) );
  NAND2_X1 U10594 ( .A1(n13111), .A2(n8272), .ZN(n8245) );
  NAND2_X1 U10595 ( .A1(n8246), .A2(n8245), .ZN(n8276) );
  AND2_X1 U10596 ( .A1(n8247), .A2(n8276), .ZN(n10380) );
  INV_X1 U10597 ( .A(n8248), .ZN(n8249) );
  NAND2_X1 U10598 ( .A1(n8250), .A2(n8249), .ZN(n8251) );
  NAND2_X1 U10599 ( .A1(n8252), .A2(n8251), .ZN(n10129) );
  NAND2_X1 U10600 ( .A1(n8285), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8256) );
  NAND2_X1 U10601 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n13507), .ZN(n8253) );
  MUX2_X1 U10602 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8253), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8255) );
  INV_X1 U10603 ( .A(n8218), .ZN(n8254) );
  NAND2_X1 U10604 ( .A1(n8255), .A2(n8254), .ZN(n10210) );
  INV_X1 U10605 ( .A(n10210), .ZN(n14667) );
  XNOR2_X1 U10606 ( .A(n14791), .B(n8834), .ZN(n8264) );
  INV_X1 U10607 ( .A(n8264), .ZN(n8262) );
  NAND2_X1 U10608 ( .A1(n8313), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8261) );
  NAND2_X1 U10609 ( .A1(n8289), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8259) );
  INV_X1 U10610 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8257) );
  NAND4_X4 U10611 ( .A1(n8261), .A2(n8260), .A3(n8259), .A4(n8258), .ZN(n13112) );
  NAND2_X1 U10612 ( .A1(n8262), .A2(n8263), .ZN(n8275) );
  NAND2_X1 U10613 ( .A1(n8265), .A2(n8264), .ZN(n8266) );
  AND2_X1 U10614 ( .A1(n8275), .A2(n8266), .ZN(n10331) );
  NAND2_X1 U10615 ( .A1(n8313), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8270) );
  NAND2_X1 U10616 ( .A1(n8289), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8268) );
  INV_X1 U10617 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n8267) );
  XNOR2_X1 U10618 ( .A(n6707), .B(n8271), .ZN(n13508) );
  MUX2_X1 U10619 ( .A(n13507), .B(n13508), .S(n8433), .Z(n11972) );
  INV_X1 U10620 ( .A(n11972), .ZN(n11968) );
  NAND2_X1 U10621 ( .A1(n11968), .A2(n8860), .ZN(n8274) );
  AND2_X1 U10622 ( .A1(n10321), .A2(n8274), .ZN(n10332) );
  NAND2_X1 U10623 ( .A1(n10330), .A2(n8275), .ZN(n10379) );
  NAND2_X1 U10624 ( .A1(n8278), .A2(n8277), .ZN(n8283) );
  MUX2_X1 U10625 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n8226), .Z(n8280) );
  INV_X1 U10626 ( .A(n8280), .ZN(n8279) );
  INV_X1 U10627 ( .A(SI_3_), .ZN(n10134) );
  NAND2_X1 U10628 ( .A1(n8279), .A2(n10134), .ZN(n8281) );
  NAND2_X1 U10629 ( .A1(n8280), .A2(SI_3_), .ZN(n8299) );
  AND2_X1 U10630 ( .A1(n8281), .A2(n8299), .ZN(n8282) );
  OR2_X1 U10631 ( .A1(n8283), .A2(n8282), .ZN(n8284) );
  NAND2_X1 U10632 ( .A1(n8300), .A2(n8284), .ZN(n10124) );
  NAND2_X1 U10633 ( .A1(n8286), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8287) );
  XNOR2_X1 U10634 ( .A(n8287), .B(P2_IR_REG_3__SCAN_IN), .ZN(n14679) );
  XNOR2_X1 U10635 ( .A(n11987), .B(n8860), .ZN(n8295) );
  NAND2_X1 U10636 ( .A1(n8313), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8294) );
  BUF_X4 U10637 ( .A(n8288), .Z(n12126) );
  NAND2_X1 U10638 ( .A1(n12126), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8293) );
  INV_X2 U10639 ( .A(n8289), .ZN(n12130) );
  NAND2_X1 U10640 ( .A1(n9027), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8292) );
  INV_X1 U10641 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8290) );
  NAND2_X1 U10642 ( .A1(n8835), .A2(n8290), .ZN(n8291) );
  NOR2_X1 U10643 ( .A1(n10586), .A2(n13359), .ZN(n8296) );
  XNOR2_X1 U10644 ( .A(n8295), .B(n8296), .ZN(n10408) );
  INV_X1 U10645 ( .A(n8295), .ZN(n8297) );
  AND2_X1 U10646 ( .A1(n8297), .A2(n8296), .ZN(n8298) );
  NAND2_X1 U10647 ( .A1(n8301), .A2(SI_4_), .ZN(n8325) );
  INV_X1 U10648 ( .A(n8301), .ZN(n8302) );
  INV_X1 U10649 ( .A(SI_4_), .ZN(n10136) );
  NAND2_X1 U10650 ( .A1(n8302), .A2(n10136), .ZN(n8303) );
  OR2_X1 U10651 ( .A1(n8305), .A2(n8304), .ZN(n8306) );
  AND2_X1 U10652 ( .A1(n8326), .A2(n8306), .ZN(n10140) );
  NAND2_X1 U10653 ( .A1(n10140), .A2(n12137), .ZN(n8312) );
  NAND2_X1 U10654 ( .A1(n8307), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8308) );
  MUX2_X1 U10655 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8308), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8310) );
  INV_X1 U10656 ( .A(n8309), .ZN(n8333) );
  NAND2_X1 U10657 ( .A1(n8310), .A2(n8333), .ZN(n13115) );
  INV_X1 U10658 ( .A(n13115), .ZN(n13121) );
  AOI22_X1 U10659 ( .A1(n8285), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n10181), 
        .B2(n13121), .ZN(n8311) );
  XNOR2_X1 U10660 ( .A(n13031), .B(n8860), .ZN(n8319) );
  INV_X2 U10661 ( .A(n8797), .ZN(n12127) );
  NAND2_X1 U10662 ( .A1(n12127), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8318) );
  NAND2_X1 U10663 ( .A1(n12126), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8317) );
  INV_X1 U10664 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8314) );
  XNOR2_X1 U10665 ( .A(n8314), .B(P2_REG3_REG_3__SCAN_IN), .ZN(n13030) );
  NAND2_X1 U10666 ( .A1(n6619), .A2(n13030), .ZN(n8316) );
  NAND2_X1 U10667 ( .A1(n8794), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8315) );
  NAND4_X1 U10668 ( .A1(n8318), .A2(n8317), .A3(n8316), .A4(n8315), .ZN(n13110) );
  NAND2_X1 U10669 ( .A1(n13110), .A2(n8272), .ZN(n8320) );
  NAND2_X1 U10670 ( .A1(n8319), .A2(n8320), .ZN(n8324) );
  INV_X1 U10671 ( .A(n8319), .ZN(n8322) );
  INV_X1 U10672 ( .A(n8320), .ZN(n8321) );
  NAND2_X1 U10673 ( .A1(n8322), .A2(n8321), .ZN(n8323) );
  AND2_X1 U10674 ( .A1(n8324), .A2(n8323), .ZN(n13028) );
  MUX2_X1 U10675 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n10067), .Z(n8327) );
  NAND2_X1 U10676 ( .A1(n8327), .A2(SI_5_), .ZN(n8350) );
  INV_X1 U10677 ( .A(n8327), .ZN(n8328) );
  INV_X1 U10678 ( .A(SI_5_), .ZN(n10138) );
  NAND2_X1 U10679 ( .A1(n8328), .A2(n10138), .ZN(n8329) );
  OR2_X1 U10680 ( .A1(n8331), .A2(n8330), .ZN(n8332) );
  NAND2_X1 U10681 ( .A1(n8351), .A2(n8332), .ZN(n10146) );
  OR2_X1 U10682 ( .A1(n10146), .A2(n12125), .ZN(n8336) );
  NAND2_X1 U10683 ( .A1(n8333), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8334) );
  XNOR2_X1 U10684 ( .A(n8334), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10276) );
  AOI22_X1 U10685 ( .A1(n8285), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n10181), 
        .B2(n10276), .ZN(n8335) );
  XNOR2_X1 U10686 ( .A(n11999), .B(n8860), .ZN(n8344) );
  NAND2_X1 U10687 ( .A1(n9028), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8343) );
  NAND2_X1 U10688 ( .A1(n9027), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8342) );
  AND3_X1 U10689 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n8362) );
  INV_X1 U10690 ( .A(n8362), .ZN(n8364) );
  INV_X1 U10691 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8338) );
  NAND2_X1 U10692 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n8337) );
  NAND2_X1 U10693 ( .A1(n8338), .A2(n8337), .ZN(n8339) );
  AND2_X1 U10694 ( .A1(n8364), .A2(n8339), .ZN(n10974) );
  NAND2_X1 U10695 ( .A1(n6619), .A2(n10974), .ZN(n8341) );
  NAND2_X1 U10696 ( .A1(n12126), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8340) );
  NAND2_X1 U10697 ( .A1(n13109), .A2(n8272), .ZN(n8345) );
  NAND2_X1 U10698 ( .A1(n8344), .A2(n8345), .ZN(n8349) );
  INV_X1 U10699 ( .A(n8344), .ZN(n8347) );
  INV_X1 U10700 ( .A(n8345), .ZN(n8346) );
  NAND2_X1 U10701 ( .A1(n8347), .A2(n8346), .ZN(n8348) );
  AND2_X1 U10702 ( .A1(n8349), .A2(n8348), .ZN(n10628) );
  NAND2_X1 U10703 ( .A1(n8352), .A2(SI_6_), .ZN(n8375) );
  INV_X1 U10704 ( .A(n8352), .ZN(n8353) );
  NAND2_X1 U10705 ( .A1(n8353), .A2(n15288), .ZN(n8354) );
  OR2_X1 U10706 ( .A1(n8356), .A2(n8355), .ZN(n8357) );
  NAND2_X1 U10707 ( .A1(n8376), .A2(n8357), .ZN(n10172) );
  INV_X1 U10708 ( .A(n8358), .ZN(n8359) );
  NAND2_X1 U10709 ( .A1(n8359), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8360) );
  XNOR2_X1 U10710 ( .A(n8360), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10263) );
  AOI22_X1 U10711 ( .A1(n9021), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n10181), 
        .B2(n10263), .ZN(n8361) );
  XNOR2_X1 U10712 ( .A(n14821), .B(n8860), .ZN(n8370) );
  NAND2_X1 U10713 ( .A1(n8362), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8386) );
  INV_X1 U10714 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8363) );
  NAND2_X1 U10715 ( .A1(n8364), .A2(n8363), .ZN(n8365) );
  AND2_X1 U10716 ( .A1(n8386), .A2(n8365), .ZN(n10998) );
  NAND2_X1 U10717 ( .A1(n6619), .A2(n10998), .ZN(n8369) );
  NAND2_X1 U10718 ( .A1(n12127), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8368) );
  NAND2_X1 U10719 ( .A1(n9027), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8367) );
  NAND2_X1 U10720 ( .A1(n12126), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8366) );
  NAND4_X1 U10721 ( .A1(n8369), .A2(n8368), .A3(n8367), .A4(n8366), .ZN(n13108) );
  NAND2_X1 U10722 ( .A1(n13108), .A2(n13336), .ZN(n8371) );
  XNOR2_X1 U10723 ( .A(n8370), .B(n8371), .ZN(n10670) );
  INV_X1 U10724 ( .A(n8370), .ZN(n8373) );
  INV_X1 U10725 ( .A(n8371), .ZN(n8372) );
  NAND2_X1 U10726 ( .A1(n8373), .A2(n8372), .ZN(n8374) );
  MUX2_X1 U10727 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n10067), .Z(n8377) );
  NAND2_X1 U10728 ( .A1(n8377), .A2(SI_7_), .ZN(n8397) );
  INV_X1 U10729 ( .A(n8377), .ZN(n8378) );
  INV_X1 U10730 ( .A(SI_7_), .ZN(n10156) );
  NAND2_X1 U10731 ( .A1(n8378), .A2(n10156), .ZN(n8379) );
  OR2_X1 U10732 ( .A1(n10179), .A2(n12125), .ZN(n8384) );
  NAND2_X1 U10733 ( .A1(n8358), .A2(n8381), .ZN(n8405) );
  NAND2_X1 U10734 ( .A1(n8405), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8382) );
  XNOR2_X1 U10735 ( .A(n8382), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10291) );
  AOI22_X1 U10736 ( .A1(n9021), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n10181), 
        .B2(n10291), .ZN(n8383) );
  NAND2_X1 U10737 ( .A1(n8384), .A2(n8383), .ZN(n12011) );
  XNOR2_X1 U10738 ( .A(n12011), .B(n8860), .ZN(n8392) );
  NAND2_X1 U10739 ( .A1(n9028), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8391) );
  NAND2_X1 U10740 ( .A1(n12126), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8390) );
  NOR2_X1 U10741 ( .A1(n8386), .A2(n8385), .ZN(n8412) );
  INV_X1 U10742 ( .A(n8412), .ZN(n8414) );
  NAND2_X1 U10743 ( .A1(n8386), .A2(n8385), .ZN(n8387) );
  AND2_X1 U10744 ( .A1(n8414), .A2(n8387), .ZN(n14760) );
  NAND2_X1 U10745 ( .A1(n6619), .A2(n14760), .ZN(n8389) );
  NAND2_X1 U10746 ( .A1(n8794), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8388) );
  NOR2_X1 U10747 ( .A1(n10829), .A2(n13359), .ZN(n8393) );
  XNOR2_X1 U10748 ( .A(n8392), .B(n8393), .ZN(n10691) );
  NAND2_X1 U10749 ( .A1(n10692), .A2(n10691), .ZN(n8396) );
  INV_X1 U10750 ( .A(n8392), .ZN(n8394) );
  NAND2_X1 U10751 ( .A1(n8394), .A2(n8393), .ZN(n8395) );
  MUX2_X1 U10752 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n10067), .Z(n8399) );
  NAND2_X1 U10753 ( .A1(n8399), .A2(SI_8_), .ZN(n8420) );
  INV_X1 U10754 ( .A(n8399), .ZN(n8400) );
  NAND2_X1 U10755 ( .A1(n8400), .A2(n10153), .ZN(n8401) );
  NAND2_X1 U10756 ( .A1(n8403), .A2(n8402), .ZN(n8421) );
  OR2_X1 U10757 ( .A1(n8403), .A2(n8402), .ZN(n8404) );
  NAND2_X1 U10758 ( .A1(n8421), .A2(n8404), .ZN(n10303) );
  OR2_X1 U10759 ( .A1(n10303), .A2(n12125), .ZN(n8411) );
  NAND2_X1 U10760 ( .A1(n8408), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8407) );
  MUX2_X1 U10761 ( .A(n8407), .B(P2_IR_REG_31__SCAN_IN), .S(n8406), .Z(n8409)
         );
  NOR2_X1 U10762 ( .A1(n8408), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8431) );
  INV_X1 U10763 ( .A(n8431), .ZN(n8428) );
  AOI22_X1 U10764 ( .A1(n8285), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n10309), 
        .B2(n10181), .ZN(n8410) );
  XNOR2_X1 U10765 ( .A(n12015), .B(n6776), .ZN(n10826) );
  NAND2_X1 U10766 ( .A1(n12126), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8419) );
  NAND2_X1 U10767 ( .A1(n12127), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8418) );
  NAND2_X1 U10768 ( .A1(n8412), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8437) );
  INV_X1 U10769 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8413) );
  NAND2_X1 U10770 ( .A1(n8414), .A2(n8413), .ZN(n8415) );
  AND2_X1 U10771 ( .A1(n8437), .A2(n8415), .ZN(n11145) );
  NAND2_X1 U10772 ( .A1(n6619), .A2(n11145), .ZN(n8417) );
  NAND2_X1 U10773 ( .A1(n9027), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8416) );
  NAND4_X1 U10774 ( .A1(n8419), .A2(n8418), .A3(n8417), .A4(n8416), .ZN(n13106) );
  NAND2_X1 U10775 ( .A1(n13106), .A2(n13336), .ZN(n10825) );
  NAND2_X1 U10776 ( .A1(n8421), .A2(n8420), .ZN(n8426) );
  MUX2_X1 U10777 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n10067), .Z(n8422) );
  NAND2_X1 U10778 ( .A1(n8422), .A2(SI_9_), .ZN(n8448) );
  INV_X1 U10779 ( .A(n8422), .ZN(n8423) );
  INV_X1 U10780 ( .A(SI_9_), .ZN(n10149) );
  NAND2_X1 U10781 ( .A1(n8423), .A2(n10149), .ZN(n8424) );
  OR2_X1 U10782 ( .A1(n8426), .A2(n8425), .ZN(n8427) );
  NAND2_X1 U10783 ( .A1(n8449), .A2(n8427), .ZN(n10337) );
  OR2_X1 U10784 ( .A1(n10337), .A2(n12125), .ZN(n8436) );
  NAND2_X1 U10785 ( .A1(n8428), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8429) );
  MUX2_X1 U10786 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8429), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n8432) );
  NAND2_X1 U10787 ( .A1(n8431), .A2(n8430), .ZN(n8476) );
  NAND2_X1 U10788 ( .A1(n8432), .A2(n8476), .ZN(n10384) );
  INV_X1 U10789 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10338) );
  OAI22_X1 U10790 ( .A1(n10384), .A2(n8433), .B1(n8457), .B2(n10338), .ZN(
        n8434) );
  INV_X1 U10791 ( .A(n8434), .ZN(n8435) );
  XNOR2_X1 U10792 ( .A(n12019), .B(n6776), .ZN(n8443) );
  NAND2_X1 U10793 ( .A1(n12126), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8442) );
  NAND2_X1 U10794 ( .A1(n12127), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8441) );
  NAND2_X1 U10795 ( .A1(n8437), .A2(n11022), .ZN(n8438) );
  AND2_X1 U10796 ( .A1(n8461), .A2(n8438), .ZN(n11097) );
  NAND2_X1 U10797 ( .A1(n6619), .A2(n11097), .ZN(n8440) );
  NAND2_X1 U10798 ( .A1(n9027), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8439) );
  NAND4_X1 U10799 ( .A1(n8442), .A2(n8441), .A3(n8440), .A4(n8439), .ZN(n13105) );
  NAND2_X1 U10800 ( .A1(n13105), .A2(n13336), .ZN(n8444) );
  XNOR2_X1 U10801 ( .A(n8443), .B(n8444), .ZN(n11020) );
  INV_X1 U10802 ( .A(n8443), .ZN(n8445) );
  NAND2_X1 U10803 ( .A1(n8445), .A2(n8444), .ZN(n8446) );
  MUX2_X1 U10804 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n10067), .Z(n8450) );
  NAND2_X1 U10805 ( .A1(n8450), .A2(SI_10_), .ZN(n8474) );
  INV_X1 U10806 ( .A(n8450), .ZN(n8451) );
  INV_X1 U10807 ( .A(SI_10_), .ZN(n10158) );
  NAND2_X1 U10808 ( .A1(n8451), .A2(n10158), .ZN(n8452) );
  OR2_X1 U10809 ( .A1(n8454), .A2(n8453), .ZN(n8455) );
  NAND2_X1 U10810 ( .A1(n8475), .A2(n8455), .ZN(n10372) );
  OR2_X1 U10811 ( .A1(n10372), .A2(n12125), .ZN(n8459) );
  NAND2_X1 U10812 ( .A1(n8476), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8456) );
  XNOR2_X1 U10813 ( .A(n8456), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10459) );
  AOI22_X1 U10814 ( .A1(n10459), .A2(n10181), .B1(n9021), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n8458) );
  XNOR2_X1 U10815 ( .A(n12022), .B(n6776), .ZN(n8467) );
  NAND2_X1 U10816 ( .A1(n12126), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8466) );
  NAND2_X1 U10817 ( .A1(n12127), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8465) );
  INV_X1 U10818 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8460) );
  NAND2_X1 U10819 ( .A1(n8461), .A2(n8460), .ZN(n8462) );
  AND2_X1 U10820 ( .A1(n8481), .A2(n8462), .ZN(n11134) );
  NAND2_X1 U10821 ( .A1(n6619), .A2(n11134), .ZN(n8464) );
  NAND2_X1 U10822 ( .A1(n9027), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8463) );
  NAND4_X1 U10823 ( .A1(n8466), .A2(n8465), .A3(n8464), .A4(n8463), .ZN(n13104) );
  AND2_X1 U10824 ( .A1(n13104), .A2(n13336), .ZN(n8468) );
  NAND2_X1 U10825 ( .A1(n8467), .A2(n8468), .ZN(n8473) );
  INV_X1 U10826 ( .A(n8467), .ZN(n8470) );
  INV_X1 U10827 ( .A(n8468), .ZN(n8469) );
  NAND2_X1 U10828 ( .A1(n8470), .A2(n8469), .ZN(n8471) );
  NAND2_X1 U10829 ( .A1(n8473), .A2(n8471), .ZN(n11118) );
  INV_X1 U10830 ( .A(n11118), .ZN(n8472) );
  MUX2_X1 U10831 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n10067), .Z(n8491) );
  XNOR2_X1 U10832 ( .A(n8491), .B(SI_11_), .ZN(n8494) );
  NAND2_X1 U10833 ( .A1(n10490), .A2(n12137), .ZN(n8479) );
  OAI21_X1 U10834 ( .B1(n8476), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8477) );
  XNOR2_X1 U10835 ( .A(n8477), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10575) );
  AOI22_X1 U10836 ( .A1(n10575), .A2(n10181), .B1(n9021), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n8478) );
  NAND2_X1 U10837 ( .A1(n12126), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8486) );
  NAND2_X1 U10838 ( .A1(n12127), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8485) );
  INV_X1 U10839 ( .A(n8502), .ZN(n8503) );
  NAND2_X1 U10840 ( .A1(n8481), .A2(n8480), .ZN(n8482) );
  AND2_X1 U10841 ( .A1(n8503), .A2(n8482), .ZN(n11267) );
  NAND2_X1 U10842 ( .A1(n6619), .A2(n11267), .ZN(n8484) );
  NAND2_X1 U10843 ( .A1(n8794), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8483) );
  NAND4_X1 U10844 ( .A1(n8486), .A2(n8485), .A3(n8484), .A4(n8483), .ZN(n13103) );
  NAND2_X1 U10845 ( .A1(n13103), .A2(n13336), .ZN(n8487) );
  XNOR2_X1 U10846 ( .A(n8489), .B(n8487), .ZN(n11195) );
  INV_X1 U10847 ( .A(n8487), .ZN(n8488) );
  NAND2_X1 U10848 ( .A1(n8489), .A2(n8488), .ZN(n8490) );
  INV_X1 U10849 ( .A(n8491), .ZN(n8492) );
  NAND2_X1 U10850 ( .A1(n8492), .A2(n10151), .ZN(n8493) );
  MUX2_X1 U10851 ( .A(n10625), .B(n10622), .S(n10067), .Z(n8516) );
  XNOR2_X1 U10852 ( .A(n8516), .B(SI_12_), .ZN(n8514) );
  XNOR2_X1 U10853 ( .A(n8515), .B(n8514), .ZN(n10621) );
  NAND2_X1 U10854 ( .A1(n10621), .A2(n12137), .ZN(n8501) );
  NAND2_X1 U10855 ( .A1(n8358), .A2(n8496), .ZN(n8498) );
  NAND2_X1 U10856 ( .A1(n8498), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8497) );
  MUX2_X1 U10857 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8497), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8499) );
  AOI22_X1 U10858 ( .A1(n8285), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n10181), 
        .B2(n11552), .ZN(n8500) );
  XNOR2_X1 U10859 ( .A(n12035), .B(n8860), .ZN(n8509) );
  NAND2_X1 U10860 ( .A1(n12126), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8508) );
  NAND2_X1 U10861 ( .A1(n12127), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8507) );
  NAND2_X1 U10862 ( .A1(n8502), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8521) );
  INV_X1 U10863 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n15327) );
  NAND2_X1 U10864 ( .A1(n8503), .A2(n15327), .ZN(n8504) );
  AND2_X1 U10865 ( .A1(n8521), .A2(n8504), .ZN(n11299) );
  NAND2_X1 U10866 ( .A1(n6619), .A2(n11299), .ZN(n8506) );
  NAND2_X1 U10867 ( .A1(n8794), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8505) );
  OR2_X1 U10868 ( .A1(n9052), .A2(n13359), .ZN(n8510) );
  NAND2_X1 U10869 ( .A1(n8509), .A2(n8510), .ZN(n11248) );
  NAND2_X1 U10870 ( .A1(n11249), .A2(n11248), .ZN(n8513) );
  INV_X1 U10871 ( .A(n8509), .ZN(n8512) );
  INV_X1 U10872 ( .A(n8510), .ZN(n8511) );
  NAND2_X1 U10873 ( .A1(n8512), .A2(n8511), .ZN(n11247) );
  NAND2_X1 U10874 ( .A1(n8513), .A2(n11247), .ZN(n11286) );
  MUX2_X1 U10875 ( .A(n7103), .B(n10683), .S(n10067), .Z(n8533) );
  XNOR2_X1 U10876 ( .A(n8533), .B(SI_13_), .ZN(n8531) );
  XNOR2_X1 U10877 ( .A(n8532), .B(n8531), .ZN(n10681) );
  NAND2_X1 U10878 ( .A1(n10681), .A2(n12137), .ZN(n8519) );
  NAND2_X1 U10879 ( .A1(n8539), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8517) );
  XNOR2_X1 U10880 ( .A(n8517), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U10881 ( .A1(n8285), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n10181), 
        .B2(n11553), .ZN(n8518) );
  XNOR2_X1 U10882 ( .A(n12044), .B(n6776), .ZN(n8529) );
  NAND2_X1 U10883 ( .A1(n12127), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8526) );
  NAND2_X1 U10884 ( .A1(n9027), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8525) );
  INV_X1 U10885 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8520) );
  NAND2_X1 U10886 ( .A1(n8521), .A2(n8520), .ZN(n8522) );
  AND2_X1 U10887 ( .A1(n8543), .A2(n8522), .ZN(n11508) );
  NAND2_X1 U10888 ( .A1(n6619), .A2(n11508), .ZN(n8524) );
  NAND2_X1 U10889 ( .A1(n12126), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8523) );
  NAND4_X1 U10890 ( .A1(n8526), .A2(n8525), .A3(n8524), .A4(n8523), .ZN(n13101) );
  NAND2_X1 U10891 ( .A1(n13101), .A2(n13336), .ZN(n8527) );
  XNOR2_X1 U10892 ( .A(n8529), .B(n8527), .ZN(n11288) );
  INV_X1 U10893 ( .A(n8527), .ZN(n8528) );
  NAND2_X1 U10894 ( .A1(n8529), .A2(n8528), .ZN(n8530) );
  NAND2_X1 U10895 ( .A1(n8532), .A2(n8531), .ZN(n8535) );
  NAND2_X1 U10896 ( .A1(n8533), .A2(n10301), .ZN(n8534) );
  INV_X1 U10897 ( .A(SI_14_), .ZN(n10328) );
  NAND2_X1 U10898 ( .A1(n8576), .A2(n10328), .ZN(n8536) );
  NAND2_X1 U10899 ( .A1(n8556), .A2(n8536), .ZN(n8537) );
  MUX2_X1 U10900 ( .A(n10808), .B(n10806), .S(n10067), .Z(n8570) );
  OR2_X1 U10901 ( .A1(n8537), .A2(n8570), .ZN(n8557) );
  NAND2_X1 U10902 ( .A1(n8537), .A2(n8570), .ZN(n8538) );
  OAI21_X1 U10903 ( .B1(n8539), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8540) );
  XNOR2_X1 U10904 ( .A(n8540), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11554) );
  AOI22_X1 U10905 ( .A1(n10181), .A2(n11554), .B1(n9021), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n8541) );
  INV_X1 U10906 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8542) );
  INV_X1 U10907 ( .A(n8564), .ZN(n8566) );
  NAND2_X1 U10908 ( .A1(n8543), .A2(n8542), .ZN(n8544) );
  NAND2_X1 U10909 ( .A1(n8566), .A2(n8544), .ZN(n11642) );
  OR2_X1 U10910 ( .A1(n11642), .A2(n8545), .ZN(n8549) );
  NAND2_X1 U10911 ( .A1(n12127), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8548) );
  NAND2_X1 U10912 ( .A1(n8794), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U10913 ( .A1(n12126), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8546) );
  NAND4_X1 U10914 ( .A1(n8549), .A2(n8548), .A3(n8547), .A4(n8546), .ZN(n13100) );
  NAND2_X1 U10915 ( .A1(n13100), .A2(n13336), .ZN(n8551) );
  NAND2_X1 U10916 ( .A1(n8550), .A2(n8551), .ZN(n8555) );
  INV_X1 U10917 ( .A(n8550), .ZN(n8553) );
  INV_X1 U10918 ( .A(n8551), .ZN(n8552) );
  NAND2_X1 U10919 ( .A1(n8553), .A2(n8552), .ZN(n8554) );
  NAND2_X1 U10920 ( .A1(n8557), .A2(n8556), .ZN(n8558) );
  MUX2_X1 U10921 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n10067), .Z(n8577) );
  XNOR2_X1 U10922 ( .A(n8577), .B(SI_15_), .ZN(n8571) );
  XNOR2_X1 U10923 ( .A(n8558), .B(n8571), .ZN(n11015) );
  NAND2_X1 U10924 ( .A1(n11015), .A2(n12137), .ZN(n8563) );
  INV_X1 U10925 ( .A(n8559), .ZN(n8560) );
  NAND2_X1 U10926 ( .A1(n8358), .A2(n8560), .ZN(n8579) );
  NAND2_X1 U10927 ( .A1(n8579), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8561) );
  XNOR2_X1 U10928 ( .A(n8561), .B(P2_IR_REG_15__SCAN_IN), .ZN(n11559) );
  AOI22_X1 U10929 ( .A1(n8285), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n10181), 
        .B2(n11559), .ZN(n8562) );
  XNOR2_X1 U10930 ( .A(n12052), .B(n8860), .ZN(n8593) );
  INV_X1 U10931 ( .A(n8583), .ZN(n8584) );
  INV_X1 U10932 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8565) );
  NAND2_X1 U10933 ( .A1(n8566), .A2(n8565), .ZN(n8567) );
  NAND2_X1 U10934 ( .A1(n8584), .A2(n8567), .ZN(n11801) );
  AOI22_X1 U10935 ( .A1(n9028), .A2(P2_REG0_REG_15__SCAN_IN), .B1(n12126), 
        .B2(P2_REG1_REG_15__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U10936 ( .A1(n8794), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8568) );
  OAI211_X1 U10937 ( .C1(n11801), .C2(n8545), .A(n8569), .B(n8568), .ZN(n13099) );
  NAND2_X1 U10938 ( .A1(n13099), .A2(n13336), .ZN(n11799) );
  AND2_X1 U10939 ( .A1(n8593), .A2(n11799), .ZN(n8596) );
  NOR2_X1 U10940 ( .A1(n8572), .A2(SI_14_), .ZN(n8575) );
  INV_X1 U10941 ( .A(n8571), .ZN(n8574) );
  NAND2_X1 U10942 ( .A1(n8572), .A2(SI_14_), .ZN(n8573) );
  INV_X1 U10943 ( .A(n8577), .ZN(n8578) );
  MUX2_X1 U10944 ( .A(n10838), .B(n10840), .S(n10067), .Z(n8600) );
  XNOR2_X1 U10945 ( .A(n8600), .B(SI_16_), .ZN(n8598) );
  XNOR2_X1 U10946 ( .A(n8599), .B(n8598), .ZN(n10837) );
  NAND2_X1 U10947 ( .A1(n10837), .A2(n12137), .ZN(n8582) );
  NAND2_X1 U10948 ( .A1(n8608), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8580) );
  XNOR2_X1 U10949 ( .A(n8580), .B(P2_IR_REG_16__SCAN_IN), .ZN(n14727) );
  AOI22_X1 U10950 ( .A1(n8285), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n14727), 
        .B2(n10181), .ZN(n8581) );
  XNOR2_X1 U10951 ( .A(n13440), .B(n8860), .ZN(n8588) );
  INV_X1 U10952 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13356) );
  INV_X1 U10953 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n13003) );
  NAND2_X1 U10954 ( .A1(n8584), .A2(n13003), .ZN(n8585) );
  NAND2_X1 U10955 ( .A1(n8613), .A2(n8585), .ZN(n13355) );
  OR2_X1 U10956 ( .A1(n13355), .A2(n8545), .ZN(n8587) );
  AOI22_X1 U10957 ( .A1(n9028), .A2(P2_REG0_REG_16__SCAN_IN), .B1(n12126), 
        .B2(P2_REG1_REG_16__SCAN_IN), .ZN(n8586) );
  OAI211_X1 U10958 ( .C1(n12130), .C2(n13356), .A(n8587), .B(n8586), .ZN(
        n13098) );
  NAND2_X1 U10959 ( .A1(n13098), .A2(n13336), .ZN(n8589) );
  NAND2_X1 U10960 ( .A1(n8588), .A2(n8589), .ZN(n8597) );
  INV_X1 U10961 ( .A(n8588), .ZN(n8591) );
  INV_X1 U10962 ( .A(n8589), .ZN(n8590) );
  NAND2_X1 U10963 ( .A1(n8591), .A2(n8590), .ZN(n8592) );
  AND2_X1 U10964 ( .A1(n8597), .A2(n8592), .ZN(n12998) );
  INV_X1 U10965 ( .A(n8593), .ZN(n12993) );
  INV_X1 U10966 ( .A(n11799), .ZN(n12995) );
  NAND2_X1 U10967 ( .A1(n12993), .A2(n12995), .ZN(n8594) );
  AND2_X1 U10968 ( .A1(n12998), .A2(n8594), .ZN(n8595) );
  NAND2_X1 U10969 ( .A1(n12997), .A2(n8597), .ZN(n13010) );
  NAND2_X1 U10970 ( .A1(n8600), .A2(n10456), .ZN(n8601) );
  MUX2_X1 U10971 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n10067), .Z(n8603) );
  OAI21_X1 U10972 ( .B1(SI_17_), .B2(n8603), .A(n8624), .ZN(n8605) );
  NAND2_X1 U10973 ( .A1(n8606), .A2(n8605), .ZN(n8607) );
  NAND2_X1 U10974 ( .A1(n8625), .A2(n8607), .ZN(n10870) );
  OR2_X1 U10975 ( .A1(n10870), .A2(n12125), .ZN(n8611) );
  OAI21_X1 U10976 ( .B1(n8608), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8609) );
  XNOR2_X1 U10977 ( .A(n8609), .B(P2_IR_REG_17__SCAN_IN), .ZN(n14749) );
  AOI22_X1 U10978 ( .A1(n10181), .A2(n14749), .B1(n9021), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n8610) );
  XNOR2_X1 U10979 ( .A(n13437), .B(n8860), .ZN(n8618) );
  INV_X1 U10980 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8612) );
  NAND2_X1 U10981 ( .A1(n8613), .A2(n8612), .ZN(n8614) );
  AND2_X1 U10982 ( .A1(n8634), .A2(n8614), .ZN(n13339) );
  NAND2_X1 U10983 ( .A1(n13339), .A2(n6619), .ZN(n8617) );
  AOI22_X1 U10984 ( .A1(n8794), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n9028), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n8616) );
  NAND2_X1 U10985 ( .A1(n12126), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8615) );
  OR2_X1 U10986 ( .A1(n13061), .A2(n13359), .ZN(n8619) );
  NAND2_X1 U10987 ( .A1(n8618), .A2(n8619), .ZN(n8623) );
  INV_X1 U10988 ( .A(n8618), .ZN(n8621) );
  INV_X1 U10989 ( .A(n8619), .ZN(n8620) );
  NAND2_X1 U10990 ( .A1(n8621), .A2(n8620), .ZN(n8622) );
  AND2_X1 U10991 ( .A1(n8623), .A2(n8622), .ZN(n13011) );
  NAND2_X1 U10992 ( .A1(n8671), .A2(SI_18_), .ZN(n8648) );
  OR2_X1 U10993 ( .A1(n8671), .A2(SI_18_), .ZN(n8626) );
  NAND2_X1 U10994 ( .A1(n8648), .A2(n8626), .ZN(n8627) );
  MUX2_X1 U10995 ( .A(n11140), .B(n11142), .S(n10067), .Z(n8672) );
  NAND2_X1 U10996 ( .A1(n8627), .A2(n8672), .ZN(n8628) );
  NAND2_X1 U10997 ( .A1(n8629), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8630) );
  XNOR2_X1 U10998 ( .A(n8630), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13136) );
  AOI22_X1 U10999 ( .A1(n8285), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n10181), 
        .B2(n13136), .ZN(n8631) );
  XNOR2_X1 U11000 ( .A(n13431), .B(n8860), .ZN(n8642) );
  INV_X1 U11001 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8633) );
  INV_X1 U11002 ( .A(n8653), .ZN(n8655) );
  NAND2_X1 U11003 ( .A1(n8634), .A2(n8633), .ZN(n8635) );
  NAND2_X1 U11004 ( .A1(n8655), .A2(n8635), .ZN(n13318) );
  OR2_X1 U11005 ( .A1(n13318), .A2(n8545), .ZN(n8640) );
  INV_X1 U11006 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n13322) );
  NAND2_X1 U11007 ( .A1(n12126), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8637) );
  NAND2_X1 U11008 ( .A1(n9028), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8636) );
  OAI211_X1 U11009 ( .C1(n13322), .C2(n12130), .A(n8637), .B(n8636), .ZN(n8638) );
  INV_X1 U11010 ( .A(n8638), .ZN(n8639) );
  NAND2_X1 U11011 ( .A1(n8640), .A2(n8639), .ZN(n13096) );
  NAND2_X1 U11012 ( .A1(n13096), .A2(n13336), .ZN(n8643) );
  XNOR2_X1 U11013 ( .A(n8642), .B(n8643), .ZN(n13059) );
  INV_X1 U11014 ( .A(n13059), .ZN(n8641) );
  INV_X1 U11015 ( .A(n8642), .ZN(n8645) );
  INV_X1 U11016 ( .A(n8643), .ZN(n8644) );
  NAND2_X1 U11017 ( .A1(n8645), .A2(n8644), .ZN(n8646) );
  NAND2_X1 U11018 ( .A1(n8649), .A2(n8648), .ZN(n8650) );
  MUX2_X1 U11019 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n10067), .Z(n8677) );
  XNOR2_X1 U11020 ( .A(n8677), .B(SI_19_), .ZN(n8674) );
  XNOR2_X1 U11021 ( .A(n8650), .B(n8674), .ZN(n11225) );
  NAND2_X1 U11022 ( .A1(n11225), .A2(n12137), .ZN(n8652) );
  AOI22_X1 U11023 ( .A1(n8285), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10181), 
        .B2(n8912), .ZN(n8651) );
  XNOR2_X1 U11024 ( .A(n13425), .B(n8860), .ZN(n8663) );
  NAND2_X1 U11025 ( .A1(n8653), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8688) );
  INV_X1 U11026 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8654) );
  NAND2_X1 U11027 ( .A1(n8655), .A2(n8654), .ZN(n8656) );
  NAND2_X1 U11028 ( .A1(n8688), .A2(n8656), .ZN(n13305) );
  OR2_X1 U11029 ( .A1(n13305), .A2(n8545), .ZN(n8662) );
  INV_X1 U11030 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13139) );
  NAND2_X1 U11031 ( .A1(n9027), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8659) );
  NAND2_X1 U11032 ( .A1(n9028), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8658) );
  OAI211_X1 U11033 ( .C1(n9032), .C2(n13139), .A(n8659), .B(n8658), .ZN(n8660)
         );
  INV_X1 U11034 ( .A(n8660), .ZN(n8661) );
  NAND2_X1 U11035 ( .A1(n8662), .A2(n8661), .ZN(n13095) );
  NAND2_X1 U11036 ( .A1(n13095), .A2(n13336), .ZN(n8664) );
  NAND2_X1 U11037 ( .A1(n8663), .A2(n8664), .ZN(n8669) );
  INV_X1 U11038 ( .A(n8663), .ZN(n8666) );
  INV_X1 U11039 ( .A(n8664), .ZN(n8665) );
  NAND2_X1 U11040 ( .A1(n8666), .A2(n8665), .ZN(n8667) );
  NAND2_X1 U11041 ( .A1(n8669), .A2(n8667), .ZN(n12966) );
  NAND2_X1 U11042 ( .A1(n8672), .A2(n10595), .ZN(n8670) );
  NAND2_X1 U11043 ( .A1(n8671), .A2(n8670), .ZN(n8676) );
  NOR2_X1 U11044 ( .A1(n8672), .A2(n10595), .ZN(n8673) );
  NOR2_X1 U11045 ( .A1(n8674), .A2(n8673), .ZN(n8675) );
  NAND2_X1 U11046 ( .A1(n8676), .A2(n8675), .ZN(n8680) );
  INV_X1 U11047 ( .A(n8677), .ZN(n8678) );
  NAND2_X1 U11048 ( .A1(n8678), .A2(n10596), .ZN(n8679) );
  NAND2_X1 U11049 ( .A1(n8684), .A2(n8683), .ZN(n8685) );
  NAND2_X1 U11050 ( .A1(n8702), .A2(n8685), .ZN(n11207) );
  OR2_X1 U11051 ( .A1(n11207), .A2(n12125), .ZN(n8687) );
  NAND2_X1 U11052 ( .A1(n9021), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8686) );
  XNOR2_X1 U11053 ( .A(n13419), .B(n8860), .ZN(n8696) );
  INV_X1 U11054 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13044) );
  NAND2_X1 U11055 ( .A1(n8688), .A2(n13044), .ZN(n8689) );
  NAND2_X1 U11056 ( .A1(n8711), .A2(n8689), .ZN(n13290) );
  OR2_X1 U11057 ( .A1(n13290), .A2(n8545), .ZN(n8695) );
  INV_X1 U11058 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8692) );
  NAND2_X1 U11059 ( .A1(n12126), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U11060 ( .A1(n9028), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8690) );
  OAI211_X1 U11061 ( .C1(n8692), .C2(n12130), .A(n8691), .B(n8690), .ZN(n8693)
         );
  INV_X1 U11062 ( .A(n8693), .ZN(n8694) );
  NAND2_X1 U11063 ( .A1(n13094), .A2(n13336), .ZN(n8697) );
  NAND2_X1 U11064 ( .A1(n8696), .A2(n8697), .ZN(n13037) );
  NAND2_X1 U11065 ( .A1(n13036), .A2(n13037), .ZN(n8700) );
  INV_X1 U11066 ( .A(n8696), .ZN(n8699) );
  INV_X1 U11067 ( .A(n8697), .ZN(n8698) );
  NAND2_X1 U11068 ( .A1(n8699), .A2(n8698), .ZN(n13038) );
  NAND2_X1 U11069 ( .A1(n8700), .A2(n13038), .ZN(n12976) );
  NAND2_X1 U11070 ( .A1(n8703), .A2(SI_21_), .ZN(n8723) );
  INV_X1 U11071 ( .A(n8703), .ZN(n8704) );
  NAND2_X1 U11072 ( .A1(n8704), .A2(n10981), .ZN(n8705) );
  NAND2_X1 U11073 ( .A1(n8707), .A2(n8706), .ZN(n8724) );
  OR2_X1 U11074 ( .A1(n8707), .A2(n8706), .ZN(n8708) );
  NAND2_X1 U11075 ( .A1(n8724), .A2(n8708), .ZN(n11283) );
  OR2_X1 U11076 ( .A1(n11283), .A2(n12125), .ZN(n8710) );
  NAND2_X1 U11077 ( .A1(n9021), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8709) );
  XNOR2_X1 U11078 ( .A(n13415), .B(n6776), .ZN(n8721) );
  INV_X1 U11079 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12978) );
  NAND2_X1 U11080 ( .A1(n8711), .A2(n12978), .ZN(n8712) );
  AND2_X1 U11081 ( .A1(n8733), .A2(n8712), .ZN(n13276) );
  NAND2_X1 U11082 ( .A1(n13276), .A2(n6619), .ZN(n8718) );
  INV_X1 U11083 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8715) );
  NAND2_X1 U11084 ( .A1(n12126), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8714) );
  NAND2_X1 U11085 ( .A1(n8794), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8713) );
  OAI211_X1 U11086 ( .C1(n8797), .C2(n8715), .A(n8714), .B(n8713), .ZN(n8716)
         );
  INV_X1 U11087 ( .A(n8716), .ZN(n8717) );
  NAND2_X1 U11088 ( .A1(n8718), .A2(n8717), .ZN(n13093) );
  NAND2_X1 U11089 ( .A1(n13093), .A2(n13336), .ZN(n8719) );
  XNOR2_X1 U11090 ( .A(n8721), .B(n8719), .ZN(n12975) );
  INV_X1 U11091 ( .A(n8719), .ZN(n8720) );
  NAND2_X1 U11092 ( .A1(n8721), .A2(n8720), .ZN(n8722) );
  INV_X1 U11093 ( .A(n8726), .ZN(n8725) );
  NAND2_X1 U11094 ( .A1(n9625), .A2(n8729), .ZN(n8730) );
  NAND2_X1 U11095 ( .A1(n8745), .A2(n8730), .ZN(n11574) );
  NAND2_X1 U11096 ( .A1(n9021), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8731) );
  XNOR2_X1 U11097 ( .A(n13410), .B(n8860), .ZN(n8740) );
  INV_X1 U11098 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13053) );
  INV_X1 U11099 ( .A(n8749), .ZN(n8750) );
  NAND2_X1 U11100 ( .A1(n8733), .A2(n13053), .ZN(n8734) );
  NAND2_X1 U11101 ( .A1(n8750), .A2(n8734), .ZN(n13260) );
  OR2_X1 U11102 ( .A1(n13260), .A2(n8545), .ZN(n8739) );
  INV_X1 U11103 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n15218) );
  NAND2_X1 U11104 ( .A1(n9027), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8736) );
  NAND2_X1 U11105 ( .A1(n9028), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8735) );
  OAI211_X1 U11106 ( .C1(n9032), .C2(n15218), .A(n8736), .B(n8735), .ZN(n8737)
         );
  INV_X1 U11107 ( .A(n8737), .ZN(n8738) );
  NAND2_X1 U11108 ( .A1(n8739), .A2(n8738), .ZN(n12977) );
  AND2_X1 U11109 ( .A1(n12977), .A2(n13336), .ZN(n13051) );
  NAND2_X1 U11110 ( .A1(n13052), .A2(n13051), .ZN(n13050) );
  INV_X1 U11111 ( .A(n8740), .ZN(n8741) );
  NAND2_X1 U11112 ( .A1(n8742), .A2(n8741), .ZN(n8743) );
  XNOR2_X1 U11113 ( .A(n8762), .B(SI_23_), .ZN(n8746) );
  XNOR2_X1 U11114 ( .A(n8764), .B(n8746), .ZN(n11774) );
  NAND2_X1 U11115 ( .A1(n11774), .A2(n12137), .ZN(n8748) );
  NAND2_X1 U11116 ( .A1(n9021), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8747) );
  XNOR2_X1 U11117 ( .A(n13404), .B(n8860), .ZN(n8757) );
  INV_X1 U11118 ( .A(n8773), .ZN(n8774) );
  INV_X1 U11119 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n12960) );
  NAND2_X1 U11120 ( .A1(n8750), .A2(n12960), .ZN(n8751) );
  NAND2_X1 U11121 ( .A1(n8774), .A2(n8751), .ZN(n13244) );
  OR2_X1 U11122 ( .A1(n13244), .A2(n8545), .ZN(n8756) );
  INV_X1 U11123 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13247) );
  NAND2_X1 U11124 ( .A1(n12126), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8753) );
  NAND2_X1 U11125 ( .A1(n9028), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8752) );
  OAI211_X1 U11126 ( .C1(n13247), .C2(n12130), .A(n8753), .B(n8752), .ZN(n8754) );
  INV_X1 U11127 ( .A(n8754), .ZN(n8755) );
  NOR2_X1 U11128 ( .A1(n13019), .A2(n13359), .ZN(n12956) );
  NAND2_X1 U11129 ( .A1(n12957), .A2(n12956), .ZN(n12955) );
  INV_X1 U11130 ( .A(n8757), .ZN(n8758) );
  NAND2_X1 U11131 ( .A1(n8759), .A2(n8758), .ZN(n8760) );
  NAND2_X1 U11132 ( .A1(n12955), .A2(n8760), .ZN(n13018) );
  INV_X1 U11133 ( .A(n8762), .ZN(n8761) );
  NOR2_X1 U11134 ( .A1(n8761), .A2(n11206), .ZN(n8763) );
  NAND2_X1 U11135 ( .A1(n8765), .A2(n11661), .ZN(n8766) );
  INV_X1 U11136 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n13504) );
  MUX2_X1 U11137 ( .A(n13504), .B(n14161), .S(n10067), .Z(n8768) );
  NAND2_X1 U11138 ( .A1(n8769), .A2(n8768), .ZN(n8770) );
  NAND2_X1 U11139 ( .A1(n8788), .A2(n8770), .ZN(n14159) );
  OR2_X1 U11140 ( .A1(n14159), .A2(n12125), .ZN(n8772) );
  NAND2_X1 U11141 ( .A1(n9021), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8771) );
  XNOR2_X1 U11142 ( .A(n13398), .B(n6776), .ZN(n8781) );
  INV_X1 U11143 ( .A(n8791), .ZN(n8792) );
  INV_X1 U11144 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13021) );
  NAND2_X1 U11145 ( .A1(n8774), .A2(n13021), .ZN(n8775) );
  NAND2_X1 U11146 ( .A1(n13233), .A2(n6619), .ZN(n8780) );
  INV_X1 U11147 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n15285) );
  NAND2_X1 U11148 ( .A1(n8794), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U11149 ( .A1(n9028), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8776) );
  OAI211_X1 U11150 ( .C1(n9032), .C2(n15285), .A(n8777), .B(n8776), .ZN(n8778)
         );
  INV_X1 U11151 ( .A(n8778), .ZN(n8779) );
  NAND2_X1 U11152 ( .A1(n8780), .A2(n8779), .ZN(n13091) );
  AND2_X1 U11153 ( .A1(n13091), .A2(n13336), .ZN(n8782) );
  NAND2_X1 U11154 ( .A1(n8781), .A2(n8782), .ZN(n8786) );
  INV_X1 U11155 ( .A(n8781), .ZN(n8784) );
  INV_X1 U11156 ( .A(n8782), .ZN(n8783) );
  NAND2_X1 U11157 ( .A1(n8784), .A2(n8783), .ZN(n8785) );
  AND2_X1 U11158 ( .A1(n8786), .A2(n8785), .ZN(n13017) );
  NAND2_X1 U11159 ( .A1(n13018), .A2(n13017), .ZN(n13016) );
  XNOR2_X1 U11160 ( .A(n8807), .B(SI_25_), .ZN(n8810) );
  XNOR2_X1 U11161 ( .A(n8811), .B(n8810), .ZN(n13501) );
  NAND2_X1 U11162 ( .A1(n13501), .A2(n12137), .ZN(n8790) );
  NAND2_X1 U11163 ( .A1(n9021), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8789) );
  XNOR2_X1 U11164 ( .A(n13393), .B(n6776), .ZN(n8801) );
  INV_X1 U11165 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n12989) );
  NAND2_X1 U11166 ( .A1(n8792), .A2(n12989), .ZN(n8793) );
  NAND2_X1 U11167 ( .A1(n8816), .A2(n8793), .ZN(n13214) );
  OR2_X1 U11168 ( .A1(n13214), .A2(n8545), .ZN(n8800) );
  INV_X1 U11169 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n15274) );
  NAND2_X1 U11170 ( .A1(n12126), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8796) );
  NAND2_X1 U11171 ( .A1(n8794), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8795) );
  OAI211_X1 U11172 ( .C1(n8797), .C2(n15274), .A(n8796), .B(n8795), .ZN(n8798)
         );
  INV_X1 U11173 ( .A(n8798), .ZN(n8799) );
  NAND2_X1 U11174 ( .A1(n8800), .A2(n8799), .ZN(n13090) );
  AND2_X1 U11175 ( .A1(n13090), .A2(n13336), .ZN(n8802) );
  NAND2_X1 U11176 ( .A1(n8801), .A2(n8802), .ZN(n8806) );
  INV_X1 U11177 ( .A(n8801), .ZN(n8804) );
  INV_X1 U11178 ( .A(n8802), .ZN(n8803) );
  NAND2_X1 U11179 ( .A1(n8804), .A2(n8803), .ZN(n8805) );
  AND2_X1 U11180 ( .A1(n8806), .A2(n8805), .ZN(n12985) );
  INV_X1 U11181 ( .A(n8807), .ZN(n8808) );
  NAND2_X1 U11182 ( .A1(n8808), .A2(n11738), .ZN(n8809) );
  XNOR2_X1 U11183 ( .A(n8827), .B(SI_26_), .ZN(n8812) );
  XNOR2_X1 U11184 ( .A(n8829), .B(n8812), .ZN(n13497) );
  NAND2_X1 U11185 ( .A1(n13497), .A2(n12137), .ZN(n8814) );
  NAND2_X1 U11186 ( .A1(n9021), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8813) );
  XNOR2_X1 U11187 ( .A(n13388), .B(n8860), .ZN(n8825) );
  INV_X1 U11188 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8815) );
  NAND2_X1 U11189 ( .A1(n8816), .A2(n8815), .ZN(n8817) );
  NAND2_X1 U11190 ( .A1(n13202), .A2(n6619), .ZN(n8823) );
  INV_X1 U11191 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8820) );
  NAND2_X1 U11192 ( .A1(n12126), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8819) );
  NAND2_X1 U11193 ( .A1(n12127), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8818) );
  OAI211_X1 U11194 ( .C1(n8820), .C2(n12130), .A(n8819), .B(n8818), .ZN(n8821)
         );
  INV_X1 U11195 ( .A(n8821), .ZN(n8822) );
  NAND2_X1 U11196 ( .A1(n8823), .A2(n8822), .ZN(n13089) );
  NAND2_X1 U11197 ( .A1(n13089), .A2(n13336), .ZN(n8824) );
  XNOR2_X1 U11198 ( .A(n8825), .B(n8824), .ZN(n13074) );
  NAND2_X1 U11199 ( .A1(n8825), .A2(n8824), .ZN(n8826) );
  INV_X1 U11200 ( .A(n8827), .ZN(n8828) );
  XNOR2_X1 U11201 ( .A(n8908), .B(SI_27_), .ZN(n8830) );
  NAND2_X1 U11202 ( .A1(n14149), .A2(n12137), .ZN(n8833) );
  NAND2_X1 U11203 ( .A1(n9021), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8832) );
  XNOR2_X1 U11204 ( .A(n13189), .B(n6776), .ZN(n8842) );
  XNOR2_X1 U11205 ( .A(n8851), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n13188) );
  NAND2_X1 U11206 ( .A1(n13188), .A2(n6619), .ZN(n8841) );
  INV_X1 U11207 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8838) );
  NAND2_X1 U11208 ( .A1(n9028), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8837) );
  NAND2_X1 U11209 ( .A1(n12126), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8836) );
  OAI211_X1 U11210 ( .C1(n8838), .C2(n12130), .A(n8837), .B(n8836), .ZN(n8839)
         );
  INV_X1 U11211 ( .A(n8839), .ZN(n8840) );
  NOR2_X1 U11212 ( .A1(n9012), .A2(n13359), .ZN(n8843) );
  NAND2_X1 U11213 ( .A1(n8842), .A2(n8843), .ZN(n8848) );
  INV_X1 U11214 ( .A(n8842), .ZN(n8845) );
  INV_X1 U11215 ( .A(n8843), .ZN(n8844) );
  NAND2_X1 U11216 ( .A1(n8845), .A2(n8844), .ZN(n8846) );
  NAND2_X1 U11217 ( .A1(n8848), .A2(n8846), .ZN(n12948) );
  INV_X1 U11218 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8850) );
  INV_X1 U11219 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8849) );
  OAI21_X1 U11220 ( .B1(n8851), .B2(n8850), .A(n8849), .ZN(n8854) );
  INV_X1 U11221 ( .A(n8851), .ZN(n8853) );
  AND2_X1 U11222 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n8852) );
  NAND2_X1 U11223 ( .A1(n8853), .A2(n8852), .ZN(n11959) );
  NAND2_X1 U11224 ( .A1(n8854), .A2(n11959), .ZN(n13173) );
  OR2_X1 U11225 ( .A1(n13173), .A2(n8545), .ZN(n8859) );
  INV_X1 U11226 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13172) );
  NAND2_X1 U11227 ( .A1(n12126), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8856) );
  NAND2_X1 U11228 ( .A1(n12127), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8855) );
  OAI211_X1 U11229 ( .C1(n13172), .C2(n12130), .A(n8856), .B(n8855), .ZN(n8857) );
  INV_X1 U11230 ( .A(n8857), .ZN(n8858) );
  NAND2_X1 U11231 ( .A1(n13087), .A2(n13336), .ZN(n8861) );
  XNOR2_X1 U11232 ( .A(n8861), .B(n8860), .ZN(n8862) );
  NAND2_X1 U11233 ( .A1(n8865), .A2(n8864), .ZN(n8872) );
  INV_X1 U11234 ( .A(n8872), .ZN(n8867) );
  NOR2_X1 U11235 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n8866) );
  NAND2_X1 U11236 ( .A1(n8880), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8869) );
  MUX2_X1 U11237 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8869), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8871) );
  NAND2_X1 U11238 ( .A1(n8872), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8902) );
  NAND2_X1 U11239 ( .A1(n8902), .A2(n8901), .ZN(n8873) );
  NAND2_X1 U11240 ( .A1(n8873), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8875) );
  INV_X1 U11241 ( .A(n13506), .ZN(n8876) );
  NOR2_X1 U11242 ( .A1(n13496), .A2(n8876), .ZN(n14777) );
  INV_X1 U11243 ( .A(n14777), .ZN(n8886) );
  INV_X1 U11244 ( .A(n8877), .ZN(n8878) );
  NAND2_X1 U11245 ( .A1(n8878), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8879) );
  MUX2_X1 U11246 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8879), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8881) );
  INV_X1 U11247 ( .A(P2_B_REG_SCAN_IN), .ZN(n8882) );
  XOR2_X1 U11248 ( .A(n13506), .B(n8882), .Z(n8883) );
  NAND2_X1 U11249 ( .A1(n13502), .A2(n8883), .ZN(n8884) );
  INV_X1 U11250 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14776) );
  NAND2_X1 U11251 ( .A1(n14771), .A2(n14776), .ZN(n8885) );
  AND2_X1 U11252 ( .A1(n8886), .A2(n8885), .ZN(n10495) );
  INV_X1 U11253 ( .A(n13502), .ZN(n8887) );
  NOR2_X1 U11254 ( .A1(n13496), .A2(n8887), .ZN(n14780) );
  INV_X1 U11255 ( .A(n14780), .ZN(n8889) );
  INV_X1 U11256 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14779) );
  NAND2_X1 U11257 ( .A1(n14771), .A2(n14779), .ZN(n8888) );
  AND2_X1 U11258 ( .A1(n8889), .A2(n8888), .ZN(n10497) );
  NOR4_X1 U11259 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n8898) );
  INV_X1 U11260 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n14773) );
  INV_X1 U11261 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n15246) );
  INV_X1 U11262 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n14774) );
  INV_X1 U11263 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15355) );
  NAND4_X1 U11264 ( .A1(n14773), .A2(n15246), .A3(n14774), .A4(n15355), .ZN(
        n8895) );
  NOR4_X1 U11265 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n8893) );
  NOR4_X1 U11266 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n8892) );
  NOR4_X1 U11267 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8891) );
  NOR4_X1 U11268 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n8890) );
  NAND4_X1 U11269 ( .A1(n8893), .A2(n8892), .A3(n8891), .A4(n8890), .ZN(n8894)
         );
  NOR4_X1 U11270 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n8895), .A4(n8894), .ZN(n8897) );
  NOR4_X1 U11271 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8896) );
  NAND3_X1 U11272 ( .A1(n8898), .A2(n8897), .A3(n8896), .ZN(n8899) );
  NAND2_X1 U11273 ( .A1(n8899), .A2(n14771), .ZN(n9086) );
  NAND3_X1 U11274 ( .A1(n10495), .A2(n10497), .A3(n9086), .ZN(n8926) );
  NOR2_X1 U11275 ( .A1(n13506), .A2(n13502), .ZN(n8900) );
  NAND2_X1 U11276 ( .A1(n13496), .A2(n8900), .ZN(n10184) );
  AND2_X1 U11277 ( .A1(n11770), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8903) );
  INV_X1 U11278 ( .A(n14781), .ZN(n14772) );
  NAND2_X1 U11279 ( .A1(n8904), .A2(n11208), .ZN(n12213) );
  INV_X1 U11280 ( .A(n10183), .ZN(n8905) );
  AND2_X1 U11281 ( .A1(n14826), .A2(n8905), .ZN(n8906) );
  INV_X1 U11282 ( .A(n8908), .ZN(n8907) );
  NOR2_X1 U11283 ( .A1(n8907), .A2(n12945), .ZN(n8909) );
  XNOR2_X1 U11284 ( .A(n9018), .B(SI_28_), .ZN(n9016) );
  XNOR2_X1 U11285 ( .A(n9017), .B(n9016), .ZN(n13489) );
  NAND2_X1 U11286 ( .A1(n13489), .A2(n12137), .ZN(n8911) );
  NAND2_X1 U11287 ( .A1(n9021), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8910) );
  AND2_X1 U11288 ( .A1(n10502), .A2(n12163), .ZN(n10741) );
  NAND2_X1 U11289 ( .A1(n8924), .A2(n10741), .ZN(n8913) );
  INV_X1 U11290 ( .A(n13491), .ZN(n8918) );
  OR2_X1 U11291 ( .A1(n11959), .A2(n8545), .ZN(n8923) );
  INV_X1 U11292 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n11958) );
  NAND2_X1 U11293 ( .A1(n12126), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8920) );
  NAND2_X1 U11294 ( .A1(n9028), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8919) );
  OAI211_X1 U11295 ( .C1(n11958), .C2(n12130), .A(n8920), .B(n8919), .ZN(n8921) );
  INV_X1 U11296 ( .A(n8921), .ZN(n8922) );
  NAND2_X1 U11297 ( .A1(n8923), .A2(n8922), .ZN(n13086) );
  AOI22_X1 U11298 ( .A1(n13088), .A2(n13075), .B1(n13076), .B2(n13086), .ZN(
        n13166) );
  INV_X1 U11299 ( .A(n8924), .ZN(n8925) );
  INV_X1 U11300 ( .A(n13173), .ZN(n8929) );
  INV_X1 U11301 ( .A(n9091), .ZN(n9087) );
  NAND2_X1 U11302 ( .A1(n8926), .A2(n9087), .ZN(n8928) );
  NAND2_X1 U11303 ( .A1(n12213), .A2(n10183), .ZN(n9084) );
  AND3_X1 U11304 ( .A1(n10184), .A2(n11770), .A3(n9084), .ZN(n8927) );
  NAND2_X1 U11305 ( .A1(n8928), .A2(n8927), .ZN(n10322) );
  AND2_X1 U11306 ( .A1(n10322), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13077) );
  AOI22_X1 U11307 ( .A1(n8929), .A2(n13077), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n8930) );
  NAND2_X1 U11308 ( .A1(n8933), .A2(n8932), .ZN(P2_U3192) );
  XNOR2_X1 U11309 ( .A(n8934), .B(n9128), .ZN(n12644) );
  NAND2_X1 U11310 ( .A1(n12666), .A2(n12667), .ZN(n12665) );
  NAND2_X1 U11311 ( .A1(n12665), .A2(n8935), .ZN(n12655) );
  NAND2_X1 U11312 ( .A1(n12653), .A2(n8936), .ZN(n8937) );
  OAI22_X1 U11313 ( .A1(n12477), .A2(n15043), .B1(n15045), .B2(n12671), .ZN(
        n8940) );
  INV_X1 U11314 ( .A(n8940), .ZN(n8941) );
  AOI21_X1 U11315 ( .B1(n12644), .B2(n15101), .A(n12648), .ZN(n12823) );
  INV_X1 U11316 ( .A(n12926), .ZN(n8944) );
  NAND2_X1 U11317 ( .A1(n9838), .A2(n8944), .ZN(n8945) );
  NAND2_X1 U11318 ( .A1(n8946), .A2(n8945), .ZN(P3_U3453) );
  OAI21_X1 U11319 ( .B1(n8947), .B2(n9257), .A(n8962), .ZN(n12641) );
  NAND2_X1 U11320 ( .A1(n12641), .A2(n14997), .ZN(n8955) );
  INV_X1 U11321 ( .A(n8949), .ZN(n8950) );
  AOI21_X1 U11322 ( .B1(n9257), .B2(n8948), .A(n8950), .ZN(n8952) );
  AOI22_X1 U11323 ( .A1(n12498), .A2(n15059), .B1(n15062), .B2(n12656), .ZN(
        n8951) );
  MUX2_X1 U11324 ( .A(n8956), .B(n8958), .S(n15132), .Z(n8957) );
  NAND2_X1 U11325 ( .A1(n8957), .A2(n7530), .ZN(P3_U3486) );
  INV_X1 U11326 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n8959) );
  MUX2_X1 U11327 ( .A(n8959), .B(n8958), .S(n15119), .Z(n8960) );
  NAND2_X1 U11328 ( .A1(n8960), .A2(n7531), .ZN(P3_U3454) );
  INV_X1 U11329 ( .A(n12631), .ZN(n8973) );
  NAND2_X1 U11330 ( .A1(n8962), .A2(n8961), .ZN(n8963) );
  XNOR2_X1 U11331 ( .A(n8963), .B(n12336), .ZN(n12632) );
  NAND2_X1 U11332 ( .A1(n12632), .A2(n15101), .ZN(n8970) );
  NAND2_X1 U11333 ( .A1(n8964), .A2(n12336), .ZN(n8965) );
  NAND2_X1 U11334 ( .A1(n8965), .A2(n8938), .ZN(n8966) );
  OR2_X1 U11335 ( .A1(n8967), .A2(n8966), .ZN(n8969) );
  AOI22_X1 U11336 ( .A1(n12499), .A2(n15062), .B1(n12497), .B2(n15059), .ZN(
        n8968) );
  NAND2_X1 U11337 ( .A1(n8970), .A2(n12635), .ZN(n8974) );
  MUX2_X1 U11338 ( .A(n8974), .B(P3_REG1_REG_28__SCAN_IN), .S(n15130), .Z(
        n8971) );
  INV_X1 U11339 ( .A(n8971), .ZN(n8972) );
  OAI21_X1 U11340 ( .B1(n12882), .B2(n8973), .A(n8972), .ZN(P3_U3487) );
  MUX2_X1 U11341 ( .A(n8974), .B(P3_REG0_REG_28__SCAN_IN), .S(n8156), .Z(n8975) );
  INV_X1 U11342 ( .A(n8975), .ZN(n8976) );
  OAI21_X1 U11343 ( .B1(n12926), .B2(n8973), .A(n8976), .ZN(P3_U3455) );
  INV_X1 U11344 ( .A(n13425), .ZN(n13301) );
  INV_X1 U11345 ( .A(n13095), .ZN(n13041) );
  INV_X1 U11346 ( .A(n13431), .ZN(n13323) );
  XNOR2_X2 U11347 ( .A(n13112), .B(n14791), .ZN(n12164) );
  NOR2_X1 U11348 ( .A1(n13114), .A2(n11968), .ZN(n10738) );
  NAND2_X1 U11349 ( .A1(n12164), .A2(n10738), .ZN(n10737) );
  INV_X1 U11350 ( .A(n14791), .ZN(n10336) );
  OR2_X1 U11351 ( .A1(n13112), .A2(n10336), .ZN(n8977) );
  NAND2_X1 U11352 ( .A1(n10841), .A2(n12165), .ZN(n8979) );
  INV_X1 U11353 ( .A(n13111), .ZN(n10411) );
  NAND2_X1 U11354 ( .A1(n10411), .A2(n11983), .ZN(n8978) );
  NAND2_X1 U11355 ( .A1(n8979), .A2(n8978), .ZN(n10983) );
  INV_X1 U11356 ( .A(n12167), .ZN(n8980) );
  NAND2_X1 U11357 ( .A1(n10983), .A2(n8980), .ZN(n8982) );
  NAND2_X1 U11358 ( .A1(n11987), .A2(n10586), .ZN(n8981) );
  NAND2_X1 U11359 ( .A1(n8982), .A2(n8981), .ZN(n10585) );
  XNOR2_X2 U11360 ( .A(n13031), .B(n13110), .ZN(n12168) );
  NAND2_X1 U11361 ( .A1(n10585), .A2(n12168), .ZN(n8984) );
  INV_X1 U11362 ( .A(n13110), .ZN(n10410) );
  NAND2_X1 U11363 ( .A1(n13031), .A2(n10410), .ZN(n8983) );
  INV_X1 U11364 ( .A(n13109), .ZN(n8985) );
  AND2_X1 U11365 ( .A1(n11999), .A2(n8985), .ZN(n8987) );
  INV_X1 U11366 ( .A(n11999), .ZN(n14812) );
  NAND2_X1 U11367 ( .A1(n14812), .A2(n13109), .ZN(n8986) );
  NAND2_X1 U11368 ( .A1(n14821), .A2(n6810), .ZN(n8989) );
  XNOR2_X1 U11369 ( .A(n12015), .B(n13106), .ZN(n12173) );
  INV_X1 U11370 ( .A(n13106), .ZN(n10693) );
  OR2_X1 U11371 ( .A1(n12015), .A2(n10693), .ZN(n8990) );
  NAND2_X1 U11372 ( .A1(n10932), .A2(n8990), .ZN(n11092) );
  XNOR2_X1 U11373 ( .A(n12019), .B(n13105), .ZN(n12174) );
  NAND2_X1 U11374 ( .A1(n11092), .A2(n12174), .ZN(n11091) );
  INV_X1 U11375 ( .A(n13105), .ZN(n10830) );
  OR2_X1 U11376 ( .A1(n12019), .A2(n10830), .ZN(n8991) );
  XNOR2_X1 U11377 ( .A(n12022), .B(n13104), .ZN(n12176) );
  INV_X1 U11378 ( .A(n13104), .ZN(n8992) );
  OR2_X1 U11379 ( .A1(n12022), .A2(n8992), .ZN(n8993) );
  XNOR2_X1 U11380 ( .A(n12031), .B(n13103), .ZN(n12179) );
  INV_X1 U11381 ( .A(n13103), .ZN(n11251) );
  NAND2_X1 U11382 ( .A1(n12031), .A2(n11251), .ZN(n8994) );
  OR2_X1 U11383 ( .A1(n12035), .A2(n9052), .ZN(n8997) );
  NAND2_X1 U11384 ( .A1(n12035), .A2(n9052), .ZN(n8995) );
  NAND2_X1 U11385 ( .A1(n8997), .A2(n8995), .ZN(n12178) );
  INV_X1 U11386 ( .A(n12178), .ZN(n8996) );
  NAND2_X1 U11387 ( .A1(n11296), .A2(n8997), .ZN(n11503) );
  XNOR2_X1 U11388 ( .A(n12044), .B(n13101), .ZN(n12180) );
  NAND2_X1 U11389 ( .A1(n11503), .A2(n12180), .ZN(n11502) );
  INV_X1 U11390 ( .A(n13101), .ZN(n11579) );
  OR2_X1 U11391 ( .A1(n12044), .A2(n11579), .ZN(n8998) );
  INV_X1 U11392 ( .A(n13100), .ZN(n12050) );
  NAND2_X1 U11393 ( .A1(n13452), .A2(n12050), .ZN(n8999) );
  OR2_X1 U11394 ( .A1(n13452), .A2(n12050), .ZN(n9000) );
  INV_X1 U11395 ( .A(n13099), .ZN(n12051) );
  NAND2_X1 U11396 ( .A1(n12052), .A2(n12051), .ZN(n9001) );
  INV_X1 U11397 ( .A(n13440), .ZN(n13008) );
  NOR2_X1 U11398 ( .A1(n13008), .A2(n13098), .ZN(n9003) );
  INV_X1 U11399 ( .A(n13098), .ZN(n9002) );
  OR2_X1 U11400 ( .A1(n13437), .A2(n13061), .ZN(n12056) );
  INV_X1 U11401 ( .A(n12056), .ZN(n9004) );
  NAND2_X1 U11402 ( .A1(n13437), .A2(n13061), .ZN(n12055) );
  INV_X1 U11403 ( .A(n13096), .ZN(n12968) );
  NAND2_X1 U11404 ( .A1(n13419), .A2(n12969), .ZN(n13269) );
  INV_X1 U11405 ( .A(n13269), .ZN(n9007) );
  OR2_X1 U11406 ( .A1(n13419), .A2(n12969), .ZN(n12162) );
  INV_X1 U11407 ( .A(n9008), .ZN(n9010) );
  INV_X1 U11408 ( .A(n13415), .ZN(n13279) );
  INV_X1 U11409 ( .A(n13093), .ZN(n13043) );
  XNOR2_X1 U11410 ( .A(n13410), .B(n12977), .ZN(n13254) );
  INV_X1 U11411 ( .A(n13410), .ZN(n13264) );
  INV_X1 U11412 ( .A(n13404), .ZN(n13248) );
  XNOR2_X1 U11413 ( .A(n13398), .B(n13091), .ZN(n13230) );
  INV_X1 U11414 ( .A(n13091), .ZN(n12987) );
  XNOR2_X1 U11415 ( .A(n13393), .B(n13090), .ZN(n12192) );
  INV_X1 U11416 ( .A(n13393), .ZN(n13217) );
  INV_X1 U11417 ( .A(n13089), .ZN(n12988) );
  XNOR2_X1 U11418 ( .A(n13189), .B(n9012), .ZN(n13186) );
  INV_X1 U11419 ( .A(n13189), .ZN(n13385) );
  NAND2_X1 U11420 ( .A1(n13377), .A2(n13087), .ZN(n9075) );
  OR2_X1 U11421 ( .A1(n13377), .A2(n13087), .ZN(n9013) );
  NAND2_X1 U11422 ( .A1(n8916), .A2(n13087), .ZN(n9014) );
  NAND2_X1 U11423 ( .A1(n9017), .A2(n9016), .ZN(n9020) );
  NAND2_X1 U11424 ( .A1(n9018), .A2(n12942), .ZN(n9019) );
  NAND2_X1 U11425 ( .A1(n9020), .A2(n9019), .ZN(n10039) );
  XNOR2_X1 U11426 ( .A(n10040), .B(SI_29_), .ZN(n10038) );
  NAND2_X1 U11427 ( .A1(n13486), .A2(n12137), .ZN(n9023) );
  NAND2_X1 U11428 ( .A1(n9021), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n9022) );
  XNOR2_X1 U11429 ( .A(n9078), .B(n13086), .ZN(n12196) );
  XNOR2_X1 U11430 ( .A(n9025), .B(n9024), .ZN(n9036) );
  NAND2_X1 U11431 ( .A1(n8912), .A2(n12215), .ZN(n9026) );
  NAND2_X1 U11432 ( .A1(n12201), .A2(n12163), .ZN(n12206) );
  NAND2_X1 U11433 ( .A1(n13087), .A2(n13075), .ZN(n9034) );
  INV_X1 U11434 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9031) );
  NAND2_X1 U11435 ( .A1(n9027), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9030) );
  NAND2_X1 U11436 ( .A1(n9028), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9029) );
  OAI211_X1 U11437 ( .C1(n9032), .C2(n9031), .A(n9030), .B(n9029), .ZN(n13085)
         );
  INV_X1 U11438 ( .A(n12214), .ZN(n10188) );
  INV_X1 U11439 ( .A(n13076), .ZN(n13042) );
  AOI21_X1 U11440 ( .B1(n10188), .B2(P2_B_REG_SCAN_IN), .A(n13042), .ZN(n13153) );
  NAND2_X1 U11441 ( .A1(n13085), .A2(n13153), .ZN(n9033) );
  XNOR2_X1 U11442 ( .A(n12052), .B(n13099), .ZN(n12184) );
  INV_X1 U11443 ( .A(n12184), .ZN(n11692) );
  OR2_X1 U11444 ( .A1(n13112), .A2(n14791), .ZN(n9037) );
  NAND2_X1 U11445 ( .A1(n10411), .A2(n6770), .ZN(n9038) );
  NAND2_X1 U11446 ( .A1(n10986), .A2(n12167), .ZN(n9040) );
  OR2_X1 U11447 ( .A1(n7497), .A2(n11987), .ZN(n9039) );
  NAND2_X1 U11448 ( .A1(n9040), .A2(n9039), .ZN(n10583) );
  INV_X1 U11449 ( .A(n12168), .ZN(n9041) );
  OR2_X1 U11450 ( .A1(n13031), .A2(n13110), .ZN(n9042) );
  NAND2_X1 U11451 ( .A1(n10995), .A2(n11000), .ZN(n10994) );
  OR2_X1 U11452 ( .A1(n14821), .A2(n13108), .ZN(n9043) );
  NAND2_X1 U11453 ( .A1(n10994), .A2(n9043), .ZN(n10877) );
  XNOR2_X1 U11454 ( .A(n12011), .B(n10829), .ZN(n12172) );
  INV_X1 U11455 ( .A(n10829), .ZN(n13107) );
  OR2_X1 U11456 ( .A1(n12011), .A2(n13107), .ZN(n9044) );
  NAND2_X1 U11457 ( .A1(n12015), .A2(n13106), .ZN(n9045) );
  INV_X1 U11458 ( .A(n12174), .ZN(n11089) );
  NAND2_X1 U11459 ( .A1(n11090), .A2(n11089), .ZN(n9047) );
  NAND2_X1 U11460 ( .A1(n12019), .A2(n13105), .ZN(n9046) );
  INV_X1 U11461 ( .A(n12176), .ZN(n11126) );
  NAND2_X1 U11462 ( .A1(n11127), .A2(n11126), .ZN(n9049) );
  NAND2_X1 U11463 ( .A1(n12022), .A2(n13104), .ZN(n9048) );
  NAND2_X1 U11464 ( .A1(n9049), .A2(n9048), .ZN(n11257) );
  NAND2_X1 U11465 ( .A1(n11257), .A2(n11261), .ZN(n9051) );
  NAND2_X1 U11466 ( .A1(n12031), .A2(n13103), .ZN(n9050) );
  AND2_X1 U11467 ( .A1(n12035), .A2(n13102), .ZN(n9053) );
  NOR2_X1 U11468 ( .A1(n12044), .A2(n13101), .ZN(n9054) );
  NAND2_X1 U11469 ( .A1(n12044), .A2(n13101), .ZN(n9055) );
  AND2_X1 U11470 ( .A1(n13452), .A2(n13100), .ZN(n9056) );
  NAND2_X1 U11471 ( .A1(n11692), .A2(n11691), .ZN(n9058) );
  OR2_X1 U11472 ( .A1(n12052), .A2(n13099), .ZN(n9057) );
  NAND2_X1 U11473 ( .A1(n9058), .A2(n9057), .ZN(n13345) );
  XNOR2_X1 U11474 ( .A(n13440), .B(n13098), .ZN(n13349) );
  NAND2_X1 U11475 ( .A1(n13440), .A2(n13098), .ZN(n9060) );
  INV_X1 U11476 ( .A(n13061), .ZN(n13097) );
  OR2_X1 U11477 ( .A1(n13437), .A2(n13097), .ZN(n9061) );
  NAND2_X1 U11478 ( .A1(n13437), .A2(n13097), .ZN(n9062) );
  NAND2_X1 U11479 ( .A1(n9063), .A2(n9062), .ZN(n13311) );
  INV_X1 U11480 ( .A(n13311), .ZN(n9065) );
  XNOR2_X1 U11481 ( .A(n13431), .B(n13096), .ZN(n13314) );
  NAND2_X1 U11482 ( .A1(n9065), .A2(n9064), .ZN(n13313) );
  OR2_X1 U11483 ( .A1(n13431), .A2(n13096), .ZN(n9066) );
  NAND2_X1 U11484 ( .A1(n13425), .A2(n13095), .ZN(n12187) );
  OR2_X1 U11485 ( .A1(n13425), .A2(n13095), .ZN(n12188) );
  NAND2_X1 U11486 ( .A1(n13419), .A2(n13094), .ZN(n9068) );
  XNOR2_X1 U11487 ( .A(n13415), .B(n13093), .ZN(n12189) );
  INV_X1 U11488 ( .A(n13254), .ZN(n13252) );
  NAND2_X1 U11489 ( .A1(n13253), .A2(n13252), .ZN(n9070) );
  NAND2_X1 U11490 ( .A1(n13410), .A2(n12977), .ZN(n9069) );
  OR2_X1 U11491 ( .A1(n13404), .A2(n13092), .ZN(n9071) );
  NAND2_X1 U11492 ( .A1(n13398), .A2(n13091), .ZN(n9072) );
  NAND2_X1 U11493 ( .A1(n13232), .A2(n9072), .ZN(n13218) );
  OR2_X1 U11494 ( .A1(n13393), .A2(n13090), .ZN(n9074) );
  AND2_X1 U11495 ( .A1(n13393), .A2(n13090), .ZN(n9073) );
  NAND2_X1 U11496 ( .A1(n13169), .A2(n9075), .ZN(n9076) );
  XNOR2_X1 U11497 ( .A(n9076), .B(n9024), .ZN(n11964) );
  INV_X1 U11498 ( .A(n14815), .ZN(n11006) );
  INV_X1 U11499 ( .A(n9078), .ZN(n12135) );
  INV_X1 U11500 ( .A(n13388), .ZN(n13204) );
  INV_X1 U11501 ( .A(n13398), .ZN(n13235) );
  INV_X1 U11502 ( .A(n12035), .ZN(n11486) );
  INV_X1 U11503 ( .A(n12019), .ZN(n11099) );
  NOR2_X1 U11504 ( .A1(n14791), .A2(n11972), .ZN(n10846) );
  NOR2_X2 U11505 ( .A1(n13031), .A2(n10988), .ZN(n10973) );
  INV_X1 U11506 ( .A(n12011), .ZN(n14765) );
  INV_X1 U11507 ( .A(n11096), .ZN(n9079) );
  NAND2_X1 U11508 ( .A1(n11099), .A2(n9079), .ZN(n11133) );
  OR2_X1 U11509 ( .A1(n11133), .A2(n12022), .ZN(n11264) );
  NOR2_X2 U11510 ( .A1(n12031), .A2(n11264), .ZN(n11298) );
  INV_X1 U11511 ( .A(n13437), .ZN(n13342) );
  NAND2_X1 U11512 ( .A1(n13362), .A2(n13342), .ZN(n13334) );
  INV_X1 U11513 ( .A(n13419), .ZN(n13294) );
  NAND2_X1 U11514 ( .A1(n13235), .A2(n13246), .ZN(n13226) );
  NAND2_X1 U11515 ( .A1(n12135), .A2(n13177), .ZN(n13156) );
  INV_X1 U11516 ( .A(n13177), .ZN(n9081) );
  AOI21_X1 U11517 ( .B1(n9078), .B2(n9081), .A(n13336), .ZN(n9082) );
  AND2_X1 U11518 ( .A1(n13156), .A2(n9082), .ZN(n11961) );
  AOI21_X1 U11519 ( .B1(n14792), .B2(n9078), .A(n11961), .ZN(n9083) );
  AND2_X1 U11520 ( .A1(n14781), .A2(n9084), .ZN(n9085) );
  AND2_X1 U11521 ( .A1(n9086), .A2(n9085), .ZN(n10498) );
  AND2_X1 U11522 ( .A1(n10495), .A2(n9087), .ZN(n9088) );
  INV_X1 U11523 ( .A(n10497), .ZN(n9092) );
  NAND2_X1 U11524 ( .A1(n9094), .A2(n14837), .ZN(n9090) );
  NAND2_X1 U11525 ( .A1(n14835), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n9089) );
  NAND2_X1 U11526 ( .A1(n9090), .A2(n9089), .ZN(P2_U3528) );
  NOR2_X1 U11527 ( .A1(n10495), .A2(n9091), .ZN(n9093) );
  NAND2_X1 U11528 ( .A1(n9094), .A2(n6621), .ZN(n9096) );
  NAND2_X1 U11529 ( .A1(n14829), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9095) );
  NAND2_X1 U11530 ( .A1(n9096), .A2(n9095), .ZN(P2_U3496) );
  INV_X1 U11531 ( .A(n12497), .ZN(n12342) );
  OR2_X1 U11532 ( .A1(n9118), .A2(n12342), .ZN(n9265) );
  INV_X1 U11533 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13483) );
  AOI22_X1 U11534 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n13483), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9100), .ZN(n9113) );
  INV_X1 U11535 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9101) );
  INV_X1 U11536 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n15239) );
  AOI22_X1 U11537 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(n9101), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(n15239), .ZN(n9102) );
  INV_X1 U11538 ( .A(n9102), .ZN(n9103) );
  XNOR2_X1 U11539 ( .A(n9104), .B(n9103), .ZN(n12934) );
  INV_X1 U11540 ( .A(SI_31_), .ZN(n12929) );
  NOR2_X1 U11541 ( .A1(n7987), .A2(n12929), .ZN(n9105) );
  INV_X1 U11542 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n9109) );
  NAND2_X1 U11543 ( .A1(n7605), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n9108) );
  NAND2_X1 U11544 ( .A1(n6620), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n9107) );
  OAI211_X1 U11545 ( .C1(n7675), .C2(n9109), .A(n9108), .B(n9107), .ZN(n9110)
         );
  INV_X1 U11546 ( .A(n9110), .ZN(n9111) );
  NAND2_X1 U11547 ( .A1(n9112), .A2(n9111), .ZN(n12614) );
  NAND2_X1 U11548 ( .A1(n14343), .A2(n12614), .ZN(n9269) );
  XNOR2_X1 U11549 ( .A(n9114), .B(n9113), .ZN(n12351) );
  NAND2_X1 U11550 ( .A1(n9106), .A2(n12351), .ZN(n9116) );
  INV_X1 U11551 ( .A(SI_30_), .ZN(n12352) );
  OR2_X1 U11552 ( .A1(n7987), .A2(n12352), .ZN(n9115) );
  NAND2_X1 U11553 ( .A1(n9116), .A2(n9115), .ZN(n14346) );
  NAND2_X1 U11554 ( .A1(n11014), .A2(n14346), .ZN(n9117) );
  NAND2_X1 U11555 ( .A1(n9269), .A2(n9117), .ZN(n9274) );
  AND2_X1 U11556 ( .A1(n9118), .A2(n12342), .ZN(n9119) );
  NOR2_X1 U11557 ( .A1(n9274), .A2(n9119), .ZN(n9271) );
  INV_X1 U11558 ( .A(n14346), .ZN(n12618) );
  INV_X1 U11559 ( .A(n12614), .ZN(n9121) );
  NOR2_X1 U11560 ( .A1(n11014), .A2(n14346), .ZN(n9120) );
  AOI21_X1 U11561 ( .B1(n9122), .B2(n9121), .A(n9120), .ZN(n9293) );
  INV_X1 U11562 ( .A(n9293), .ZN(n9268) );
  NAND2_X1 U11563 ( .A1(n9268), .A2(n9122), .ZN(n9123) );
  NAND2_X1 U11564 ( .A1(n9124), .A2(n9123), .ZN(n9125) );
  XNOR2_X1 U11565 ( .A(n9125), .B(n12607), .ZN(n9127) );
  NOR2_X1 U11566 ( .A1(n9127), .A2(n9126), .ZN(n9299) );
  NAND2_X1 U11567 ( .A1(n9257), .A2(n9128), .ZN(n9275) );
  MUX2_X1 U11568 ( .A(n9229), .B(n9228), .S(n9854), .Z(n9236) );
  CLKBUF_X1 U11569 ( .A(n9129), .Z(n9130) );
  NAND2_X1 U11570 ( .A1(n15061), .A2(n11954), .ZN(n9276) );
  NAND2_X1 U11571 ( .A1(n9276), .A2(n10752), .ZN(n9135) );
  OAI22_X1 U11572 ( .A1(n9131), .A2(n11451), .B1(n9301), .B2(n9276), .ZN(n9132) );
  NAND2_X1 U11573 ( .A1(n9132), .A2(n9140), .ZN(n9134) );
  OAI211_X1 U11574 ( .C1(n9130), .C2(n9135), .A(n9134), .B(n9133), .ZN(n9144)
         );
  INV_X1 U11575 ( .A(n9144), .ZN(n9139) );
  NAND2_X1 U11576 ( .A1(n9145), .A2(n9136), .ZN(n9137) );
  AOI21_X1 U11577 ( .B1(n9139), .B2(n9138), .A(n9137), .ZN(n9148) );
  INV_X1 U11578 ( .A(n9140), .ZN(n9143) );
  NAND2_X1 U11579 ( .A1(n15060), .A2(n15050), .ZN(n9142) );
  OAI211_X1 U11580 ( .C1(n9144), .C2(n9143), .A(n9142), .B(n9141), .ZN(n9146)
         );
  NAND2_X1 U11581 ( .A1(n9146), .A2(n9145), .ZN(n9147) );
  MUX2_X1 U11582 ( .A(n9148), .B(n9147), .S(n10752), .Z(n9154) );
  NAND3_X1 U11583 ( .A1(n12504), .A2(n15033), .A3(n9854), .ZN(n9149) );
  NAND2_X1 U11584 ( .A1(n11450), .A2(n9149), .ZN(n9153) );
  MUX2_X1 U11585 ( .A(n9151), .B(n9150), .S(n10752), .Z(n9152) );
  OAI211_X1 U11586 ( .C1(n9154), .C2(n9153), .A(n15014), .B(n9152), .ZN(n9158)
         );
  NAND2_X1 U11587 ( .A1(n9163), .A2(n9155), .ZN(n9156) );
  NAND2_X1 U11588 ( .A1(n9156), .A2(n10752), .ZN(n9157) );
  NAND2_X1 U11589 ( .A1(n9158), .A2(n9157), .ZN(n9162) );
  AOI21_X1 U11590 ( .B1(n9161), .B2(n9159), .A(n10752), .ZN(n9160) );
  AOI21_X1 U11591 ( .B1(n9162), .B2(n9161), .A(n9160), .ZN(n9167) );
  OAI21_X1 U11592 ( .B1(n10752), .B2(n9163), .A(n11834), .ZN(n9166) );
  MUX2_X1 U11593 ( .A(n11705), .B(n9164), .S(n9854), .Z(n9165) );
  OAI211_X1 U11594 ( .C1(n9167), .C2(n9166), .A(n7014), .B(n9165), .ZN(n9171)
         );
  INV_X1 U11595 ( .A(n11814), .ZN(n11811) );
  MUX2_X1 U11596 ( .A(n9169), .B(n9168), .S(n10752), .Z(n9170) );
  NAND4_X1 U11597 ( .A1(n9171), .A2(n11727), .A3(n11811), .A4(n9170), .ZN(
        n9184) );
  OAI21_X1 U11598 ( .B1(n11814), .B2(n9173), .A(n9172), .ZN(n9176) );
  OAI21_X1 U11599 ( .B1(n11814), .B2(n11809), .A(n9174), .ZN(n9175) );
  MUX2_X1 U11600 ( .A(n9176), .B(n9175), .S(n10752), .Z(n9177) );
  NOR2_X1 U11601 ( .A1(n9177), .A2(n11893), .ZN(n9183) );
  NAND2_X1 U11602 ( .A1(n9186), .A2(n9178), .ZN(n9181) );
  NAND2_X1 U11603 ( .A1(n9185), .A2(n9179), .ZN(n9180) );
  MUX2_X1 U11604 ( .A(n9181), .B(n9180), .S(n10752), .Z(n9182) );
  AOI21_X1 U11605 ( .B1(n9184), .B2(n9183), .A(n9182), .ZN(n9192) );
  MUX2_X1 U11606 ( .A(n9186), .B(n9185), .S(n9854), .Z(n9187) );
  INV_X1 U11607 ( .A(n12812), .ZN(n12809) );
  NAND2_X1 U11608 ( .A1(n9187), .A2(n12809), .ZN(n9191) );
  MUX2_X1 U11609 ( .A(n9189), .B(n9188), .S(n10752), .Z(n9190) );
  OAI21_X1 U11610 ( .B1(n9192), .B2(n9191), .A(n9190), .ZN(n9193) );
  INV_X1 U11611 ( .A(n12800), .ZN(n9284) );
  NAND2_X1 U11612 ( .A1(n9193), .A2(n9284), .ZN(n9196) );
  MUX2_X1 U11613 ( .A(n12785), .B(n9194), .S(n10752), .Z(n9195) );
  NAND3_X1 U11614 ( .A1(n9196), .A2(n12787), .A3(n9195), .ZN(n9200) );
  OAI21_X1 U11615 ( .B1(n12802), .B2(n12484), .A(n9203), .ZN(n9197) );
  NAND2_X1 U11616 ( .A1(n9197), .A2(n9854), .ZN(n9199) );
  INV_X1 U11617 ( .A(n9202), .ZN(n9198) );
  AOI21_X1 U11618 ( .B1(n9200), .B2(n9199), .A(n9198), .ZN(n9205) );
  AOI21_X1 U11619 ( .B1(n9202), .B2(n9201), .A(n9854), .ZN(n9204) );
  OAI22_X1 U11620 ( .A1(n9205), .A2(n9204), .B1(n9203), .B2(n9854), .ZN(n9212)
         );
  INV_X1 U11621 ( .A(n9206), .ZN(n9211) );
  NAND2_X1 U11622 ( .A1(n9208), .A2(n9207), .ZN(n9209) );
  AOI21_X1 U11623 ( .B1(n9209), .B2(n9213), .A(n9854), .ZN(n9210) );
  NAND2_X1 U11624 ( .A1(n9219), .A2(n9210), .ZN(n9214) );
  AOI22_X1 U11625 ( .A1(n9212), .A2(n12763), .B1(n9211), .B2(n9214), .ZN(n9217) );
  NAND3_X1 U11626 ( .A1(n9218), .A2(n9213), .A3(n9854), .ZN(n9215) );
  NAND2_X1 U11627 ( .A1(n9215), .A2(n9214), .ZN(n9216) );
  OAI21_X1 U11628 ( .B1(n9217), .B2(n7900), .A(n9216), .ZN(n9221) );
  MUX2_X1 U11629 ( .A(n9219), .B(n9218), .S(n10752), .Z(n9220) );
  NAND3_X1 U11630 ( .A1(n9221), .A2(n8102), .A3(n9220), .ZN(n9227) );
  NAND2_X1 U11631 ( .A1(n12848), .A2(n12710), .ZN(n9223) );
  MUX2_X1 U11632 ( .A(n9223), .B(n9222), .S(n10752), .Z(n9226) );
  NAND2_X1 U11633 ( .A1(n9225), .A2(n9224), .ZN(n12708) );
  NAND3_X1 U11634 ( .A1(n9227), .A2(n9226), .A3(n12708), .ZN(n9234) );
  NAND2_X1 U11635 ( .A1(n9229), .A2(n9228), .ZN(n12697) );
  INV_X1 U11636 ( .A(n12697), .ZN(n9233) );
  NAND2_X1 U11637 ( .A1(n12722), .A2(n9854), .ZN(n9231) );
  NAND2_X1 U11638 ( .A1(n12700), .A2(n10752), .ZN(n9230) );
  MUX2_X1 U11639 ( .A(n9231), .B(n9230), .S(n12383), .Z(n9232) );
  NAND3_X1 U11640 ( .A1(n9234), .A2(n9233), .A3(n9232), .ZN(n9235) );
  NAND3_X1 U11641 ( .A1(n9236), .A2(n12690), .A3(n9235), .ZN(n9238) );
  NAND3_X1 U11642 ( .A1(n12689), .A2(n12699), .A3(n10752), .ZN(n9237) );
  AND2_X1 U11643 ( .A1(n9238), .A2(n9237), .ZN(n9245) );
  NAND2_X1 U11644 ( .A1(n9240), .A2(n9239), .ZN(n9241) );
  NAND2_X1 U11645 ( .A1(n9241), .A2(n9242), .ZN(n9243) );
  MUX2_X1 U11646 ( .A(n9243), .B(n9242), .S(n10752), .Z(n9244) );
  OAI21_X1 U11647 ( .B1(n9245), .B2(n12667), .A(n9244), .ZN(n9251) );
  NOR2_X1 U11648 ( .A1(n12396), .A2(n12671), .ZN(n9248) );
  INV_X1 U11649 ( .A(n9246), .ZN(n9247) );
  MUX2_X1 U11650 ( .A(n9248), .B(n9247), .S(n9854), .Z(n9249) );
  INV_X1 U11651 ( .A(n9249), .ZN(n9250) );
  OAI21_X1 U11652 ( .B1(n12654), .B2(n9251), .A(n9250), .ZN(n9259) );
  MUX2_X1 U11653 ( .A(n9253), .B(n9252), .S(n10752), .Z(n9254) );
  INV_X1 U11654 ( .A(n9254), .ZN(n9256) );
  NOR2_X1 U11655 ( .A1(n12477), .A2(n10752), .ZN(n9255) );
  AOI22_X1 U11656 ( .A1(n9257), .A2(n9256), .B1(n12639), .B2(n9255), .ZN(n9258) );
  OAI21_X1 U11657 ( .B1(n9275), .B2(n9259), .A(n9258), .ZN(n9260) );
  NAND2_X1 U11658 ( .A1(n9260), .A2(n12336), .ZN(n9267) );
  NAND2_X1 U11659 ( .A1(n9261), .A2(n10752), .ZN(n9263) );
  NAND2_X1 U11660 ( .A1(n9263), .A2(n9262), .ZN(n9264) );
  NAND2_X1 U11661 ( .A1(n9267), .A2(n9264), .ZN(n9266) );
  OAI211_X1 U11662 ( .C1(n9267), .C2(n10752), .A(n9266), .B(n9265), .ZN(n9270)
         );
  AOI22_X1 U11663 ( .A1(n9271), .A2(n9270), .B1(n9269), .B2(n9268), .ZN(n9273)
         );
  INV_X1 U11664 ( .A(n9272), .ZN(n9300) );
  INV_X1 U11665 ( .A(n9274), .ZN(n9294) );
  INV_X1 U11666 ( .A(n9275), .ZN(n9290) );
  INV_X1 U11667 ( .A(n9276), .ZN(n9277) );
  NOR2_X1 U11668 ( .A1(n9131), .A2(n9277), .ZN(n11950) );
  NAND4_X1 U11669 ( .A1(n11950), .A2(n15014), .A3(n7014), .A4(n11811), .ZN(
        n9282) );
  INV_X1 U11670 ( .A(n9130), .ZN(n11072) );
  NAND4_X1 U11671 ( .A1(n11834), .A2(n11450), .A3(n11072), .A4(n11897), .ZN(
        n9281) );
  NAND3_X1 U11672 ( .A1(n9279), .A2(n14337), .A3(n9278), .ZN(n9280) );
  NOR3_X1 U11673 ( .A1(n9282), .A2(n9281), .A3(n9280), .ZN(n9283) );
  AND4_X1 U11674 ( .A1(n9283), .A2(n9133), .A3(n12809), .A4(n11727), .ZN(n9285) );
  NAND4_X1 U11675 ( .A1(n9285), .A2(n12776), .A3(n9284), .A4(n12787), .ZN(
        n9286) );
  NOR4_X1 U11676 ( .A1(n7900), .A2(n7880), .A3(n7461), .A4(n9286), .ZN(n9287)
         );
  NAND3_X1 U11677 ( .A1(n9287), .A2(n8102), .A3(n12708), .ZN(n9288) );
  NOR4_X1 U11678 ( .A1(n12667), .A2(n12680), .A3(n12697), .A4(n9288), .ZN(
        n9289) );
  AND4_X1 U11679 ( .A1(n12336), .A2(n9290), .A3(n9289), .A4(n12651), .ZN(n9292) );
  NAND4_X1 U11680 ( .A1(n9294), .A2(n9293), .A3(n9292), .A4(n9291), .ZN(n9295)
         );
  XNOR2_X1 U11681 ( .A(n9295), .B(n12595), .ZN(n9296) );
  NAND2_X1 U11682 ( .A1(n9296), .A2(n6845), .ZN(n9297) );
  OR2_X1 U11683 ( .A1(n10751), .A2(P3_U3151), .ZN(n11204) );
  INV_X1 U11684 ( .A(n11204), .ZN(n9298) );
  NAND2_X1 U11685 ( .A1(n10749), .A2(n9300), .ZN(n9863) );
  NOR3_X1 U11686 ( .A1(n9863), .A2(n15045), .A3(n6628), .ZN(n9303) );
  OAI21_X1 U11687 ( .B1(n11204), .B2(n9301), .A(P3_B_REG_SCAN_IN), .ZN(n9302)
         );
  NAND2_X1 U11688 ( .A1(n9305), .A2(n9304), .ZN(P3_U3296) );
  NOR2_X1 U11689 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n9309) );
  NAND4_X1 U11690 ( .A1(n9309), .A2(n9308), .A3(n9307), .A4(n9306), .ZN(n9312)
         );
  NAND4_X1 U11691 ( .A1(n9310), .A2(n9503), .A3(n9462), .A4(n9518), .ZN(n9311)
         );
  NOR2_X1 U11692 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n9317) );
  NOR2_X1 U11693 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n9316) );
  NOR2_X1 U11694 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n9315) );
  NOR3_X1 U11695 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .A3(P1_IR_REG_25__SCAN_IN), .ZN(n9318) );
  OR2_X1 U11696 ( .A1(n6623), .A2(n15324), .ZN(n9322) );
  INV_X1 U11697 ( .A(n14042), .ZN(n13834) );
  NAND2_X1 U11698 ( .A1(n9725), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9334) );
  INV_X2 U11699 ( .A(n9552), .ZN(n10049) );
  NAND2_X1 U11700 ( .A1(n10049), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9333) );
  NAND2_X1 U11701 ( .A1(n9418), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9431) );
  NOR2_X1 U11702 ( .A1(n9431), .A2(n9430), .ZN(n9443) );
  NAND2_X1 U11703 ( .A1(n9443), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9454) );
  INV_X1 U11704 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9453) );
  INV_X1 U11705 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9483) );
  NAND2_X1 U11706 ( .A1(n9493), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9510) );
  INV_X1 U11707 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n9509) );
  INV_X1 U11708 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9524) );
  INV_X1 U11709 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9565) );
  INV_X1 U11710 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13615) );
  NAND2_X1 U11711 ( .A1(n9605), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n9628) );
  NAND2_X1 U11712 ( .A1(n9618), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9636) );
  NAND2_X1 U11713 ( .A1(n9627), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9645) );
  NAND2_X1 U11714 ( .A1(n9635), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n9347) );
  NAND2_X1 U11715 ( .A1(n9644), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9335) );
  INV_X1 U11716 ( .A(n9335), .ZN(n9346) );
  NAND2_X1 U11717 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n9346), .ZN(n9336) );
  INV_X1 U11718 ( .A(n9336), .ZN(n9329) );
  NAND2_X1 U11719 ( .A1(n9329), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9656) );
  INV_X1 U11720 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13511) );
  NAND2_X1 U11721 ( .A1(n9336), .A2(n13511), .ZN(n9330) );
  NAND2_X1 U11722 ( .A1(n9665), .A2(n13830), .ZN(n9332) );
  AND2_X2 U11723 ( .A1(n11945), .A2(n14146), .ZN(n9379) );
  NAND2_X1 U11724 ( .A1(n9379), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9331) );
  NAND4_X1 U11725 ( .A1(n9334), .A2(n9333), .A3(n9332), .A4(n9331), .ZN(n14047) );
  INV_X1 U11726 ( .A(n14047), .ZN(n13845) );
  NAND2_X1 U11727 ( .A1(n9725), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9341) );
  NAND2_X1 U11728 ( .A1(n10049), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9340) );
  INV_X1 U11729 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13643) );
  NAND2_X1 U11730 ( .A1(n13643), .A2(n9335), .ZN(n9337) );
  AND2_X1 U11731 ( .A1(n9337), .A2(n9336), .ZN(n13846) );
  NAND2_X1 U11732 ( .A1(n9665), .A2(n13846), .ZN(n9339) );
  NAND2_X1 U11733 ( .A1(n9379), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9338) );
  NAND4_X1 U11734 ( .A1(n9341), .A2(n9340), .A3(n9339), .A4(n9338), .ZN(n13859) );
  INV_X1 U11735 ( .A(n13859), .ZN(n14038) );
  NAND2_X1 U11736 ( .A1(n13497), .A2(n10071), .ZN(n9343) );
  OR2_X1 U11737 ( .A1(n6623), .A2(n14154), .ZN(n9342) );
  INV_X1 U11738 ( .A(n13851), .ZN(n14050) );
  NAND2_X1 U11739 ( .A1(n13501), .A2(n10071), .ZN(n9345) );
  OR2_X1 U11740 ( .A1(n6623), .A2(n14157), .ZN(n9344) );
  NAND2_X1 U11741 ( .A1(n9725), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9351) );
  NAND2_X1 U11742 ( .A1(n10049), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9350) );
  INV_X1 U11743 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n13572) );
  AOI21_X1 U11744 ( .B1(n13572), .B2(n9347), .A(n9346), .ZN(n13864) );
  NAND2_X1 U11745 ( .A1(n9665), .A2(n13864), .ZN(n9349) );
  NAND2_X1 U11746 ( .A1(n9379), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9348) );
  NAND4_X1 U11747 ( .A1(n9351), .A2(n9350), .A3(n9349), .A4(n9348), .ZN(n14046) );
  XNOR2_X1 U11748 ( .A(n14057), .B(n14046), .ZN(n13868) );
  INV_X1 U11749 ( .A(n13868), .ZN(n9651) );
  NAND2_X1 U11750 ( .A1(n9617), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9355) );
  NAND2_X1 U11751 ( .A1(n9379), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9354) );
  NAND2_X1 U11752 ( .A1(n9380), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9353) );
  NAND2_X1 U11753 ( .A1(n9568), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9352) );
  AND4_X2 U11754 ( .A1(n9355), .A2(n9354), .A3(n9353), .A4(n9352), .ZN(n9363)
         );
  INV_X1 U11755 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10128) );
  INV_X1 U11756 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9357) );
  NAND2_X1 U11757 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n6762), .ZN(n9356) );
  XNOR2_X1 U11758 ( .A(n9357), .B(n9356), .ZN(n10431) );
  NAND2_X1 U11759 ( .A1(n9363), .A2(n14558), .ZN(n9888) );
  NAND2_X1 U11760 ( .A1(n9617), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9361) );
  NAND2_X1 U11761 ( .A1(n9379), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9360) );
  NAND2_X1 U11762 ( .A1(n9380), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9359) );
  NAND2_X1 U11763 ( .A1(n9568), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9358) );
  AND4_X2 U11764 ( .A1(n9361), .A2(n9360), .A3(n9359), .A4(n9358), .ZN(n10706)
         );
  XNOR2_X1 U11765 ( .A(n9362), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14163) );
  MUX2_X1 U11766 ( .A(n6762), .B(n14163), .S(n10176), .Z(n14013) );
  INV_X1 U11767 ( .A(n14013), .ZN(n9877) );
  OR2_X1 U11768 ( .A1(n10706), .A2(n9877), .ZN(n10702) );
  NAND2_X1 U11769 ( .A1(n10707), .A2(n10702), .ZN(n9365) );
  NAND2_X1 U11770 ( .A1(n9363), .A2(n10703), .ZN(n9364) );
  NAND2_X1 U11771 ( .A1(n9365), .A2(n9364), .ZN(n10716) );
  NAND2_X1 U11772 ( .A1(n9568), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9369) );
  NAND2_X1 U11773 ( .A1(n9617), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9368) );
  NAND2_X1 U11774 ( .A1(n9379), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9367) );
  NAND2_X1 U11775 ( .A1(n9380), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9366) );
  NAND4_X2 U11776 ( .A1(n9369), .A2(n9368), .A3(n9367), .A4(n9366), .ZN(n9894)
         );
  NOR2_X1 U11777 ( .A1(n9370), .A2(n14138), .ZN(n9371) );
  MUX2_X1 U11778 ( .A(n14138), .B(n9371), .S(P1_IR_REG_2__SCAN_IN), .Z(n9372)
         );
  INV_X1 U11779 ( .A(n9372), .ZN(n9374) );
  INV_X1 U11780 ( .A(n9388), .ZN(n9373) );
  NAND2_X1 U11781 ( .A1(n9374), .A2(n9373), .ZN(n13690) );
  INV_X1 U11782 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10126) );
  OR2_X1 U11783 ( .A1(n6623), .A2(n10126), .ZN(n9376) );
  OR2_X1 U11784 ( .A1(n10046), .A2(n10127), .ZN(n9375) );
  OAI211_X2 U11785 ( .C1(n6772), .C2(n13690), .A(n9376), .B(n9375), .ZN(n10727) );
  NAND2_X1 U11786 ( .A1(n10716), .A2(n10715), .ZN(n9378) );
  INV_X1 U11787 ( .A(n9894), .ZN(n9739) );
  INV_X1 U11788 ( .A(n10727), .ZN(n14569) );
  NAND2_X1 U11789 ( .A1(n9739), .A2(n14569), .ZN(n9377) );
  NAND2_X1 U11790 ( .A1(n9568), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9384) );
  INV_X1 U11791 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14537) );
  NAND2_X1 U11792 ( .A1(n9665), .A2(n14537), .ZN(n9383) );
  NAND2_X1 U11793 ( .A1(n9379), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9382) );
  NAND2_X1 U11794 ( .A1(n9380), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9381) );
  NOR2_X1 U11795 ( .A1(n9388), .A2(n14138), .ZN(n9385) );
  MUX2_X1 U11796 ( .A(n14138), .B(n9385), .S(P1_IR_REG_3__SCAN_IN), .Z(n9386)
         );
  INV_X1 U11797 ( .A(n9386), .ZN(n9389) );
  INV_X1 U11798 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9387) );
  NAND2_X1 U11799 ( .A1(n9388), .A2(n9387), .ZN(n9400) );
  NAND2_X1 U11800 ( .A1(n9389), .A2(n9400), .ZN(n13705) );
  OR2_X1 U11801 ( .A1(n6772), .A2(n13705), .ZN(n9392) );
  INV_X1 U11802 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10125) );
  OR2_X1 U11803 ( .A1(n6623), .A2(n10125), .ZN(n9391) );
  XNOR2_X1 U11804 ( .A(n14583), .B(n6626), .ZN(n10086) );
  NAND2_X1 U11805 ( .A1(n14529), .A2(n14531), .ZN(n9394) );
  INV_X1 U11806 ( .A(n14583), .ZN(n10964) );
  INV_X1 U11807 ( .A(n6626), .ZN(n14576) );
  NAND2_X1 U11808 ( .A1(n10964), .A2(n14576), .ZN(n9393) );
  NAND2_X1 U11809 ( .A1(n9394), .A2(n9393), .ZN(n10891) );
  NAND2_X1 U11810 ( .A1(n10049), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9398) );
  NAND2_X1 U11811 ( .A1(n10050), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9397) );
  XNOR2_X1 U11812 ( .A(n14537), .B(P1_REG3_REG_4__SCAN_IN), .ZN(n10961) );
  NAND2_X1 U11813 ( .A1(n9665), .A2(n10961), .ZN(n9396) );
  NAND2_X1 U11814 ( .A1(n9725), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9395) );
  NAND2_X1 U11815 ( .A1(n10140), .A2(n10071), .ZN(n9403) );
  INV_X2 U11816 ( .A(n6623), .ZN(n9590) );
  NAND2_X1 U11817 ( .A1(n9400), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9399) );
  MUX2_X1 U11818 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9399), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n9401) );
  AND2_X1 U11819 ( .A1(n9401), .A2(n9536), .ZN(n10539) );
  AOI22_X1 U11820 ( .A1(n9590), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n9589), .B2(
        n10539), .ZN(n9402) );
  INV_X1 U11821 ( .A(n10959), .ZN(n14585) );
  INV_X1 U11822 ( .A(n10892), .ZN(n9404) );
  NAND2_X1 U11823 ( .A1(n10891), .A2(n9404), .ZN(n9406) );
  INV_X1 U11824 ( .A(n13671), .ZN(n11038) );
  NAND2_X1 U11825 ( .A1(n11038), .A2(n10959), .ZN(n9405) );
  AOI21_X1 U11826 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9407) );
  NOR2_X1 U11827 ( .A1(n9407), .A2(n9418), .ZN(n14520) );
  NAND2_X1 U11828 ( .A1(n10050), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9408) );
  AND2_X1 U11829 ( .A1(n9409), .A2(n9408), .ZN(n9411) );
  NAND2_X1 U11830 ( .A1(n9725), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9410) );
  OR2_X1 U11831 ( .A1(n10146), .A2(n10046), .ZN(n9414) );
  NAND2_X1 U11832 ( .A1(n9536), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9412) );
  XNOR2_X1 U11833 ( .A(n9412), .B(P1_IR_REG_5__SCAN_IN), .ZN(n13722) );
  AOI22_X1 U11834 ( .A1(n9590), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9589), .B2(
        n13722), .ZN(n9413) );
  NAND2_X1 U11835 ( .A1(n9414), .A2(n9413), .ZN(n11040) );
  INV_X1 U11836 ( .A(n11040), .ZN(n14594) );
  OR2_X1 U11837 ( .A1(n10172), .A2(n10046), .ZN(n9417) );
  NOR2_X1 U11838 ( .A1(n9536), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n9426) );
  OR2_X1 U11839 ( .A1(n9426), .A2(n14138), .ZN(n9415) );
  XNOR2_X1 U11840 ( .A(n9415), .B(P1_IR_REG_6__SCAN_IN), .ZN(n13737) );
  AOI22_X1 U11841 ( .A1(n9590), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9589), .B2(
        n13737), .ZN(n9416) );
  NAND2_X1 U11842 ( .A1(n10049), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9422) );
  NAND2_X1 U11843 ( .A1(n10050), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9421) );
  OAI21_X1 U11844 ( .B1(n9418), .B2(P1_REG3_REG_6__SCAN_IN), .A(n9431), .ZN(
        n10905) );
  INV_X1 U11845 ( .A(n10905), .ZN(n11181) );
  NAND2_X1 U11846 ( .A1(n9665), .A2(n11181), .ZN(n9420) );
  NAND2_X1 U11847 ( .A1(n9725), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9419) );
  NAND4_X1 U11848 ( .A1(n9422), .A2(n9421), .A3(n9420), .A4(n9419), .ZN(n13670) );
  XNOR2_X1 U11849 ( .A(n11180), .B(n13670), .ZN(n10897) );
  INV_X1 U11850 ( .A(n10897), .ZN(n10900) );
  OR2_X1 U11851 ( .A1(n11180), .A2(n13670), .ZN(n9423) );
  OR2_X1 U11852 ( .A1(n10179), .A2(n10046), .ZN(n9429) );
  INV_X1 U11853 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9425) );
  NAND2_X1 U11854 ( .A1(n9426), .A2(n9425), .ZN(n9439) );
  NAND2_X1 U11855 ( .A1(n9439), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9427) );
  XNOR2_X1 U11856 ( .A(n9427), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10476) );
  AOI22_X1 U11857 ( .A1(n9590), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9589), .B2(
        n10476), .ZN(n9428) );
  NAND2_X1 U11858 ( .A1(n9429), .A2(n9428), .ZN(n11217) );
  NAND2_X1 U11859 ( .A1(n9725), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9436) );
  NAND2_X1 U11860 ( .A1(n10049), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9435) );
  AND2_X1 U11861 ( .A1(n9431), .A2(n9430), .ZN(n9432) );
  NOR2_X1 U11862 ( .A1(n9443), .A2(n9432), .ZN(n14506) );
  NAND2_X1 U11863 ( .A1(n9665), .A2(n14506), .ZN(n9434) );
  NAND2_X1 U11864 ( .A1(n10050), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9433) );
  NAND4_X1 U11865 ( .A1(n9436), .A2(n9435), .A3(n9434), .A4(n9433), .ZN(n14616) );
  XNOR2_X1 U11866 ( .A(n11217), .B(n14616), .ZN(n14502) );
  INV_X1 U11867 ( .A(n14502), .ZN(n14499) );
  NAND2_X1 U11868 ( .A1(n14500), .A2(n14499), .ZN(n9438) );
  OR2_X1 U11869 ( .A1(n11217), .A2(n14616), .ZN(n9437) );
  NAND2_X1 U11870 ( .A1(n9438), .A2(n9437), .ZN(n11104) );
  OR2_X1 U11871 ( .A1(n10303), .A2(n10046), .ZN(n9442) );
  NAND2_X1 U11872 ( .A1(n9450), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9440) );
  XNOR2_X1 U11873 ( .A(n9440), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10544) );
  AOI22_X1 U11874 ( .A1(n9590), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9589), .B2(
        n10544), .ZN(n9441) );
  NAND2_X1 U11875 ( .A1(n9725), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9448) );
  NAND2_X1 U11876 ( .A1(n10049), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9447) );
  OR2_X1 U11877 ( .A1(n9443), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9444) );
  AND2_X1 U11878 ( .A1(n9454), .A2(n9444), .ZN(n11337) );
  NAND2_X1 U11879 ( .A1(n9665), .A2(n11337), .ZN(n9446) );
  NAND2_X1 U11880 ( .A1(n10050), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9445) );
  OR2_X1 U11881 ( .A1(n11338), .A2(n11607), .ZN(n9930) );
  NAND2_X1 U11882 ( .A1(n11338), .A2(n11607), .ZN(n9929) );
  NAND2_X1 U11883 ( .A1(n11104), .A2(n11107), .ZN(n9449) );
  INV_X1 U11884 ( .A(n11607), .ZN(n13669) );
  OR2_X1 U11885 ( .A1(n11338), .A2(n13669), .ZN(n9933) );
  NAND2_X1 U11886 ( .A1(n9449), .A2(n9933), .ZN(n11153) );
  OR2_X1 U11887 ( .A1(n10337), .A2(n10046), .ZN(n9452) );
  OR2_X1 U11888 ( .A1(n9477), .A2(n14138), .ZN(n9463) );
  XNOR2_X1 U11889 ( .A(n9463), .B(P1_IR_REG_9__SCAN_IN), .ZN(n13754) );
  AOI22_X1 U11890 ( .A1(n9590), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9589), .B2(
        n13754), .ZN(n9451) );
  INV_X1 U11891 ( .A(n14627), .ZN(n11162) );
  NAND2_X1 U11892 ( .A1(n10049), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9459) );
  NAND2_X1 U11893 ( .A1(n9725), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9458) );
  NAND2_X1 U11894 ( .A1(n9454), .A2(n9453), .ZN(n9455) );
  AND2_X1 U11895 ( .A1(n9468), .A2(n9455), .ZN(n11611) );
  NAND2_X1 U11896 ( .A1(n9665), .A2(n11611), .ZN(n9457) );
  NAND2_X1 U11897 ( .A1(n10050), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9456) );
  XNOR2_X1 U11898 ( .A(n11162), .B(n11678), .ZN(n10090) );
  NAND2_X1 U11899 ( .A1(n11153), .A2(n10090), .ZN(n9461) );
  NAND2_X1 U11900 ( .A1(n14627), .A2(n11678), .ZN(n9460) );
  NAND2_X1 U11901 ( .A1(n9461), .A2(n9460), .ZN(n11306) );
  OR2_X1 U11902 ( .A1(n10372), .A2(n10046), .ZN(n9467) );
  NAND2_X1 U11903 ( .A1(n9463), .A2(n9462), .ZN(n9464) );
  NAND2_X1 U11904 ( .A1(n9464), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9465) );
  XNOR2_X1 U11905 ( .A(n9465), .B(P1_IR_REG_10__SCAN_IN), .ZN(n13768) );
  AOI22_X1 U11906 ( .A1(n9590), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n13768), 
        .B2(n9589), .ZN(n9466) );
  NAND2_X1 U11907 ( .A1(n10049), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9473) );
  NAND2_X1 U11908 ( .A1(n10050), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n9472) );
  NAND2_X1 U11909 ( .A1(n9468), .A2(n11677), .ZN(n9469) );
  AND2_X1 U11910 ( .A1(n9484), .A2(n9469), .ZN(n11680) );
  NAND2_X1 U11911 ( .A1(n9665), .A2(n11680), .ZN(n9471) );
  NAND2_X1 U11912 ( .A1(n9725), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9470) );
  NAND4_X1 U11913 ( .A1(n9473), .A2(n9472), .A3(n9471), .A4(n9470), .ZN(n13668) );
  INV_X1 U11914 ( .A(n13668), .ZN(n11608) );
  OR2_X1 U11915 ( .A1(n14636), .A2(n11608), .ZN(n9749) );
  NAND2_X1 U11916 ( .A1(n14636), .A2(n11608), .ZN(n9474) );
  NAND2_X1 U11917 ( .A1(n9749), .A2(n9474), .ZN(n11310) );
  OR2_X1 U11918 ( .A1(n14636), .A2(n13668), .ZN(n9475) );
  NAND2_X1 U11919 ( .A1(n10490), .A2(n10071), .ZN(n9482) );
  NOR2_X1 U11920 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n9476) );
  NAND2_X1 U11921 ( .A1(n9477), .A2(n9476), .ZN(n9489) );
  NAND2_X1 U11922 ( .A1(n9489), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9479) );
  INV_X1 U11923 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9478) );
  XNOR2_X1 U11924 ( .A(n9479), .B(n9478), .ZN(n10660) );
  OAI22_X1 U11925 ( .A1(n6623), .A2(n10494), .B1(n10660), .B2(n6772), .ZN(
        n9480) );
  INV_X1 U11926 ( .A(n9480), .ZN(n9481) );
  NAND2_X1 U11927 ( .A1(n10049), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9488) );
  NOR2_X1 U11928 ( .A1(n9493), .A2(n7540), .ZN(n14381) );
  NAND2_X1 U11929 ( .A1(n9665), .A2(n14381), .ZN(n9487) );
  NAND2_X1 U11930 ( .A1(n10050), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9486) );
  NAND2_X1 U11931 ( .A1(n9725), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9485) );
  NAND4_X1 U11932 ( .A1(n9488), .A2(n9487), .A3(n9486), .A4(n9485), .ZN(n14288) );
  XNOR2_X1 U11933 ( .A(n14383), .B(n11792), .ZN(n14384) );
  NAND2_X1 U11934 ( .A1(n10621), .A2(n10071), .ZN(n9492) );
  OR2_X1 U11935 ( .A1(n9489), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9490) );
  NAND2_X1 U11936 ( .A1(n9490), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9504) );
  XNOR2_X1 U11937 ( .A(n9504), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10815) );
  AOI22_X1 U11938 ( .A1(n9589), .A2(n10815), .B1(n9590), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n9491) );
  NAND2_X1 U11939 ( .A1(n9725), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9498) );
  NAND2_X1 U11940 ( .A1(n10049), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9497) );
  OR2_X1 U11941 ( .A1(n9493), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9494) );
  AND2_X1 U11942 ( .A1(n9494), .A2(n9510), .ZN(n11789) );
  NAND2_X1 U11943 ( .A1(n9665), .A2(n11789), .ZN(n9496) );
  NAND2_X1 U11944 ( .A1(n10050), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9495) );
  NAND4_X1 U11945 ( .A1(n9498), .A2(n9497), .A3(n9496), .A4(n9495), .ZN(n13667) );
  INV_X1 U11946 ( .A(n13667), .ZN(n9499) );
  OR2_X1 U11947 ( .A1(n14290), .A2(n9499), .ZN(n9751) );
  NAND2_X1 U11948 ( .A1(n14290), .A2(n9499), .ZN(n9500) );
  NAND2_X1 U11949 ( .A1(n9751), .A2(n9500), .ZN(n10092) );
  NAND2_X1 U11950 ( .A1(n11463), .A2(n10092), .ZN(n9502) );
  OR2_X1 U11951 ( .A1(n14290), .A2(n13667), .ZN(n9501) );
  NAND2_X1 U11952 ( .A1(n9502), .A2(n9501), .ZN(n14308) );
  NAND2_X1 U11953 ( .A1(n10681), .A2(n10071), .ZN(n9508) );
  NAND2_X1 U11954 ( .A1(n9504), .A2(n9503), .ZN(n9505) );
  NAND2_X1 U11955 ( .A1(n9505), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9519) );
  XNOR2_X1 U11956 ( .A(n9519), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10857) );
  NOR2_X1 U11957 ( .A1(n6623), .A2(n10683), .ZN(n9506) );
  AOI21_X1 U11958 ( .B1(n10857), .B2(n9589), .A(n9506), .ZN(n9507) );
  NAND2_X1 U11959 ( .A1(n10049), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9515) );
  NAND2_X1 U11960 ( .A1(n10050), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9514) );
  NAND2_X1 U11961 ( .A1(n9510), .A2(n9509), .ZN(n9511) );
  AND2_X1 U11962 ( .A1(n9525), .A2(n9511), .ZN(n14306) );
  NAND2_X1 U11963 ( .A1(n9665), .A2(n14306), .ZN(n9513) );
  NAND2_X1 U11964 ( .A1(n9725), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9512) );
  NAND4_X1 U11965 ( .A1(n9515), .A2(n9514), .A3(n9513), .A4(n9512), .ZN(n14289) );
  XNOR2_X1 U11966 ( .A(n14310), .B(n14289), .ZN(n14302) );
  INV_X1 U11967 ( .A(n14302), .ZN(n14307) );
  OR2_X1 U11968 ( .A1(n14310), .A2(n14289), .ZN(n9516) );
  OR2_X1 U11969 ( .A1(n10807), .A2(n10046), .ZN(n9523) );
  NAND2_X1 U11970 ( .A1(n9519), .A2(n9518), .ZN(n9520) );
  NAND2_X1 U11971 ( .A1(n9520), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9521) );
  XNOR2_X1 U11972 ( .A(n9521), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11350) );
  AOI22_X1 U11973 ( .A1(n11350), .A2(n9589), .B1(n9590), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9522) );
  NAND2_X1 U11974 ( .A1(n10049), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9530) );
  NAND2_X1 U11975 ( .A1(n9725), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9529) );
  AND2_X1 U11976 ( .A1(n9525), .A2(n9524), .ZN(n9526) );
  NOR2_X1 U11977 ( .A1(n9540), .A2(n9526), .ZN(n13523) );
  NAND2_X1 U11978 ( .A1(n9665), .A2(n13523), .ZN(n9528) );
  NAND2_X1 U11979 ( .A1(n10050), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9527) );
  NAND2_X1 U11980 ( .A1(n14414), .A2(n12229), .ZN(n9958) );
  NAND2_X1 U11981 ( .A1(n9959), .A2(n9958), .ZN(n10095) );
  NAND2_X1 U11982 ( .A1(n14414), .A2(n9531), .ZN(n9533) );
  NAND2_X1 U11983 ( .A1(n11015), .A2(n10071), .ZN(n9539) );
  INV_X1 U11984 ( .A(n9534), .ZN(n9535) );
  OAI21_X1 U11985 ( .B1(n9536), .B2(n9535), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9537) );
  XNOR2_X1 U11986 ( .A(n9537), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11364) );
  AOI22_X1 U11987 ( .A1(n9590), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9589), 
        .B2(n11364), .ZN(n9538) );
  NOR2_X1 U11988 ( .A1(n9540), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9541) );
  NOR2_X1 U11989 ( .A1(n9554), .A2(n9541), .ZN(n14365) );
  NAND2_X1 U11990 ( .A1(n14365), .A2(n9665), .ZN(n9545) );
  NAND2_X1 U11991 ( .A1(n9725), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9544) );
  NAND2_X1 U11992 ( .A1(n10049), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n9543) );
  NAND2_X1 U11993 ( .A1(n10050), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n9542) );
  NAND2_X1 U11994 ( .A1(n14366), .A2(n14409), .ZN(n9963) );
  NAND2_X1 U11995 ( .A1(n14370), .A2(n14369), .ZN(n14368) );
  INV_X1 U11996 ( .A(n14409), .ZN(n14393) );
  OR2_X1 U11997 ( .A1(n14366), .A2(n14393), .ZN(n9546) );
  NAND2_X1 U11998 ( .A1(n14368), .A2(n9546), .ZN(n11903) );
  NAND2_X1 U11999 ( .A1(n10837), .A2(n10071), .ZN(n9551) );
  NAND2_X1 U12000 ( .A1(n9547), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9548) );
  MUX2_X1 U12001 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9548), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n9549) );
  INV_X1 U12002 ( .A(n9575), .ZN(n9561) );
  AND2_X1 U12003 ( .A1(n9549), .A2(n9561), .ZN(n11360) );
  AOI22_X1 U12004 ( .A1(n9590), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9589), 
        .B2(n11360), .ZN(n9550) );
  INV_X1 U12005 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9553) );
  INV_X1 U12006 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11623) );
  OAI22_X1 U12007 ( .A1(n10053), .A2(n9553), .B1(n9552), .B2(n11623), .ZN(
        n9558) );
  OR2_X1 U12008 ( .A1(n9554), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9555) );
  NAND2_X1 U12009 ( .A1(n9566), .A2(n9555), .ZN(n11909) );
  INV_X1 U12010 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9556) );
  OAI22_X1 U12011 ( .A1(n11909), .A2(n9607), .B1(n9729), .B2(n9556), .ZN(n9557) );
  INV_X1 U12012 ( .A(n13666), .ZN(n13993) );
  XNOR2_X1 U12013 ( .A(n12244), .B(n13993), .ZN(n11904) );
  NAND2_X1 U12014 ( .A1(n11903), .A2(n11904), .ZN(n9560) );
  OR2_X1 U12015 ( .A1(n12244), .A2(n13666), .ZN(n9559) );
  OR2_X1 U12016 ( .A1(n10870), .A2(n10046), .ZN(n9564) );
  NAND2_X1 U12017 ( .A1(n9561), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9562) );
  XNOR2_X1 U12018 ( .A(n9562), .B(P1_IR_REG_17__SCAN_IN), .ZN(n13778) );
  AOI22_X1 U12019 ( .A1(n9590), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9589), 
        .B2(n13778), .ZN(n9563) );
  NAND2_X1 U12020 ( .A1(n9566), .A2(n9565), .ZN(n9567) );
  AND2_X1 U12021 ( .A1(n9580), .A2(n9567), .ZN(n14001) );
  NAND2_X1 U12022 ( .A1(n14001), .A2(n9665), .ZN(n9571) );
  AOI22_X1 U12023 ( .A1(n9725), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n10049), 
        .B2(P1_REG2_REG_17__SCAN_IN), .ZN(n9570) );
  NAND2_X1 U12024 ( .A1(n10050), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9569) );
  NOR2_X1 U12025 ( .A1(n14116), .A2(n14394), .ZN(n9572) );
  NAND2_X1 U12026 ( .A1(n14116), .A2(n14394), .ZN(n9573) );
  OR2_X1 U12027 ( .A1(n11141), .A2(n10046), .ZN(n9579) );
  INV_X1 U12028 ( .A(n9586), .ZN(n9576) );
  NAND2_X1 U12029 ( .A1(n9576), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9577) );
  XNOR2_X1 U12030 ( .A(n9577), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13787) );
  AOI22_X1 U12031 ( .A1(n9590), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9589), 
        .B2(n13787), .ZN(n9578) );
  AND2_X1 U12032 ( .A1(n9580), .A2(n15330), .ZN(n9581) );
  OR2_X1 U12033 ( .A1(n9581), .A2(n9593), .ZN(n13636) );
  AOI22_X1 U12034 ( .A1(n10049), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10050), 
        .B2(P1_REG0_REG_18__SCAN_IN), .ZN(n9583) );
  NAND2_X1 U12035 ( .A1(n9725), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9582) );
  OAI211_X1 U12036 ( .C1(n13636), .C2(n9607), .A(n9583), .B(n9582), .ZN(n13959) );
  NAND2_X1 U12037 ( .A1(n14110), .A2(n13959), .ZN(n9984) );
  INV_X1 U12038 ( .A(n9984), .ZN(n9584) );
  OR2_X1 U12039 ( .A1(n14110), .A2(n13959), .ZN(n9981) );
  NAND2_X1 U12040 ( .A1(n11225), .A2(n10071), .ZN(n9592) );
  INV_X1 U12041 ( .A(n9703), .ZN(n9587) );
  NAND2_X1 U12042 ( .A1(n9587), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9588) );
  AOI22_X1 U12043 ( .A1(n9590), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n13944), 
        .B2(n9589), .ZN(n9591) );
  OR2_X1 U12044 ( .A1(n9593), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9594) );
  NAND2_X1 U12045 ( .A1(n9604), .A2(n9594), .ZN(n13961) );
  OR2_X1 U12046 ( .A1(n13961), .A2(n9607), .ZN(n9599) );
  INV_X1 U12047 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13784) );
  NAND2_X1 U12048 ( .A1(n10050), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U12049 ( .A1(n10049), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n9595) );
  OAI211_X1 U12050 ( .C1(n10053), .C2(n13784), .A(n9596), .B(n9595), .ZN(n9597) );
  INV_X1 U12051 ( .A(n9597), .ZN(n9598) );
  NAND2_X1 U12052 ( .A1(n9599), .A2(n9598), .ZN(n13665) );
  INV_X1 U12053 ( .A(n13954), .ZN(n10101) );
  NAND2_X1 U12054 ( .A1(n13952), .A2(n10101), .ZN(n9601) );
  OR2_X1 U12055 ( .A1(n14106), .A2(n13665), .ZN(n9600) );
  INV_X1 U12056 ( .A(n13948), .ZN(n9613) );
  OR2_X1 U12057 ( .A1(n11207), .A2(n10046), .ZN(n9603) );
  OR2_X1 U12058 ( .A1(n6623), .A2(n11202), .ZN(n9602) );
  NAND2_X1 U12059 ( .A1(n9604), .A2(n13615), .ZN(n9606) );
  INV_X1 U12060 ( .A(n9605), .ZN(n9619) );
  NAND2_X1 U12061 ( .A1(n9606), .A2(n9619), .ZN(n13943) );
  OR2_X1 U12062 ( .A1(n13943), .A2(n9607), .ZN(n9612) );
  INV_X1 U12063 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n15390) );
  NAND2_X1 U12064 ( .A1(n9725), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n9609) );
  NAND2_X1 U12065 ( .A1(n10049), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9608) );
  OAI211_X1 U12066 ( .C1(n15390), .C2(n9729), .A(n9609), .B(n9608), .ZN(n9610)
         );
  INV_X1 U12067 ( .A(n9610), .ZN(n9611) );
  XNOR2_X1 U12068 ( .A(n13946), .B(n14103), .ZN(n10098) );
  NAND2_X2 U12069 ( .A1(n9613), .A2(n10098), .ZN(n14093) );
  OR2_X1 U12070 ( .A1(n14096), .A2(n14103), .ZN(n9614) );
  OR2_X1 U12071 ( .A1(n11283), .A2(n10046), .ZN(n9616) );
  OR2_X1 U12072 ( .A1(n6623), .A2(n11282), .ZN(n9615) );
  NAND2_X1 U12073 ( .A1(n9725), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n9623) );
  NAND2_X1 U12074 ( .A1(n10049), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9622) );
  INV_X1 U12075 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13565) );
  AOI21_X1 U12076 ( .B1(n13565), .B2(n9619), .A(n9618), .ZN(n13929) );
  NAND2_X1 U12077 ( .A1(n9665), .A2(n13929), .ZN(n9621) );
  NAND2_X1 U12078 ( .A1(n9379), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9620) );
  NAND4_X1 U12079 ( .A1(n9623), .A2(n9622), .A3(n9621), .A4(n9620), .ZN(n14076) );
  INV_X1 U12080 ( .A(n14076), .ZN(n13624) );
  XNOR2_X1 U12081 ( .A(n14088), .B(n13624), .ZN(n10100) );
  OR2_X1 U12082 ( .A1(n14088), .A2(n14076), .ZN(n9624) );
  OR2_X1 U12083 ( .A1(n9625), .A2(n7572), .ZN(n9626) );
  XNOR2_X1 U12084 ( .A(n9626), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14162) );
  NAND2_X1 U12085 ( .A1(n9725), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n9632) );
  NAND2_X1 U12086 ( .A1(n10049), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9631) );
  INV_X1 U12087 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13626) );
  AOI21_X1 U12088 ( .B1(n13626), .B2(n9628), .A(n9627), .ZN(n13625) );
  NAND2_X1 U12089 ( .A1(n9665), .A2(n13625), .ZN(n9630) );
  NAND2_X1 U12090 ( .A1(n9379), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9629) );
  NAND4_X1 U12091 ( .A1(n9632), .A2(n9631), .A3(n9630), .A4(n9629), .ZN(n13664) );
  XNOR2_X1 U12092 ( .A(n14080), .B(n13664), .ZN(n13906) );
  NAND2_X1 U12093 ( .A1(n11774), .A2(n10071), .ZN(n9634) );
  OR2_X1 U12094 ( .A1(n6623), .A2(n11777), .ZN(n9633) );
  NAND2_X1 U12095 ( .A1(n9725), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9640) );
  NAND2_X1 U12096 ( .A1(n10049), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9639) );
  INV_X1 U12097 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13530) );
  AOI21_X1 U12098 ( .B1(n13530), .B2(n9636), .A(n9635), .ZN(n13898) );
  NAND2_X1 U12099 ( .A1(n9665), .A2(n13898), .ZN(n9638) );
  NAND2_X1 U12100 ( .A1(n9379), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9637) );
  XNOR2_X1 U12101 ( .A(n13899), .B(n13916), .ZN(n13892) );
  NAND2_X1 U12102 ( .A1(n13893), .A2(n13892), .ZN(n13895) );
  OR2_X1 U12103 ( .A1(n14071), .A2(n13916), .ZN(n9641) );
  OR2_X1 U12104 ( .A1(n6623), .A2(n14161), .ZN(n9642) );
  NAND2_X1 U12105 ( .A1(n10049), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9649) );
  NAND2_X1 U12106 ( .A1(n9379), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9648) );
  INV_X1 U12107 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13605) );
  AOI21_X1 U12108 ( .B1(n13605), .B2(n9645), .A(n9644), .ZN(n13882) );
  NAND2_X1 U12109 ( .A1(n9665), .A2(n13882), .ZN(n9647) );
  NAND2_X1 U12110 ( .A1(n9725), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9646) );
  NAND4_X1 U12111 ( .A1(n9649), .A2(n9648), .A3(n9647), .A4(n9646), .ZN(n13860) );
  XNOR2_X1 U12112 ( .A(n14066), .B(n13860), .ZN(n13871) );
  INV_X1 U12113 ( .A(n13860), .ZN(n13574) );
  NAND2_X1 U12114 ( .A1(n13885), .A2(n13574), .ZN(n9650) );
  NAND2_X1 U12115 ( .A1(n14057), .A2(n14046), .ZN(n9652) );
  NAND2_X1 U12116 ( .A1(n14060), .A2(n9652), .ZN(n13855) );
  XNOR2_X1 U12117 ( .A(n13851), .B(n13859), .ZN(n13841) );
  NAND2_X1 U12118 ( .A1(n13855), .A2(n13854), .ZN(n14052) );
  NAND2_X1 U12119 ( .A1(n13489), .A2(n10071), .ZN(n9654) );
  OR2_X1 U12120 ( .A1(n6623), .A2(n14148), .ZN(n9653) );
  NAND2_X1 U12121 ( .A1(n9725), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9661) );
  NAND2_X1 U12122 ( .A1(n10049), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9660) );
  INV_X1 U12123 ( .A(n9656), .ZN(n9655) );
  NAND2_X1 U12124 ( .A1(n9655), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9730) );
  INV_X1 U12125 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n12329) );
  NAND2_X1 U12126 ( .A1(n9656), .A2(n12329), .ZN(n9657) );
  NAND2_X1 U12127 ( .A1(n9665), .A2(n13817), .ZN(n9659) );
  NAND2_X1 U12128 ( .A1(n9379), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9658) );
  NAND4_X1 U12129 ( .A1(n9661), .A2(n9660), .A3(n9659), .A4(n9658), .ZN(n13663) );
  NAND2_X1 U12130 ( .A1(n13821), .A2(n13663), .ZN(n9663) );
  OR2_X1 U12131 ( .A1(n13821), .A2(n13663), .ZN(n9662) );
  NAND2_X1 U12132 ( .A1(n9725), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9669) );
  NAND2_X1 U12133 ( .A1(n10049), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9668) );
  INV_X1 U12134 ( .A(n9730), .ZN(n9664) );
  NAND2_X1 U12135 ( .A1(n9665), .A2(n9664), .ZN(n9667) );
  NAND2_X1 U12136 ( .A1(n10050), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n9666) );
  NAND4_X1 U12137 ( .A1(n9669), .A2(n9668), .A3(n9667), .A4(n9666), .ZN(n14031) );
  NAND2_X1 U12138 ( .A1(n13486), .A2(n10071), .ZN(n9671) );
  OR2_X1 U12139 ( .A1(n6623), .A2(n14144), .ZN(n9670) );
  INV_X1 U12140 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9674) );
  NAND2_X1 U12141 ( .A1(n9678), .A2(n9674), .ZN(n9679) );
  NAND2_X1 U12142 ( .A1(n9679), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9675) );
  MUX2_X1 U12143 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9675), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9677) );
  INV_X1 U12144 ( .A(n9676), .ZN(n9682) );
  NAND2_X1 U12145 ( .A1(n14155), .A2(P1_B_REG_SCAN_IN), .ZN(n9681) );
  MUX2_X1 U12146 ( .A(P1_B_REG_SCAN_IN), .B(n9681), .S(n14158), .Z(n9685) );
  NAND2_X1 U12147 ( .A1(n9682), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9684) );
  NOR4_X1 U12148 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n9694) );
  NOR4_X1 U12149 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n9693) );
  INV_X1 U12150 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n15300) );
  INV_X1 U12151 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n14553) );
  INV_X1 U12152 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15286) );
  INV_X1 U12153 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n14554) );
  NAND4_X1 U12154 ( .A1(n15300), .A2(n14553), .A3(n15286), .A4(n14554), .ZN(
        n9691) );
  NOR4_X1 U12155 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9689) );
  NOR4_X1 U12156 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n9688) );
  NOR4_X1 U12157 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9687) );
  NOR4_X1 U12158 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9686) );
  NAND4_X1 U12159 ( .A1(n9689), .A2(n9688), .A3(n9687), .A4(n9686), .ZN(n9690)
         );
  NOR4_X1 U12160 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9691), .A4(n9690), .ZN(n9692) );
  AND3_X1 U12161 ( .A1(n9694), .A2(n9693), .A3(n9692), .ZN(n9695) );
  NOR2_X1 U12162 ( .A1(n10202), .A2(n9695), .ZN(n10352) );
  INV_X1 U12163 ( .A(n10352), .ZN(n9698) );
  INV_X1 U12164 ( .A(n14158), .ZN(n9696) );
  OAI22_X1 U12165 ( .A1(n10202), .A2(P1_D_REG_0__SCAN_IN), .B1(n9697), .B2(
        n9696), .ZN(n10353) );
  AND2_X1 U12166 ( .A1(n9698), .A2(n10353), .ZN(n14121) );
  INV_X1 U12167 ( .A(n10202), .ZN(n9699) );
  INV_X1 U12168 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10164) );
  NAND2_X1 U12169 ( .A1(n9699), .A2(n10164), .ZN(n9701) );
  NAND2_X1 U12170 ( .A1(n14155), .A2(n14152), .ZN(n9700) );
  NAND2_X1 U12171 ( .A1(n9701), .A2(n9700), .ZN(n10518) );
  INV_X1 U12172 ( .A(n10366), .ZN(n9708) );
  NOR2_X1 U12173 ( .A1(n14158), .A2(n14152), .ZN(n9705) );
  NAND2_X2 U12174 ( .A1(n9705), .A2(n9706), .ZN(n10344) );
  INV_X1 U12175 ( .A(n10515), .ZN(n9709) );
  NOR2_X1 U12176 ( .A1(n10518), .A2(n9709), .ZN(n10162) );
  XNOR2_X2 U12177 ( .A(n9713), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9719) );
  NAND2_X1 U12178 ( .A1(n9879), .A2(n9719), .ZN(n10175) );
  NAND2_X1 U12179 ( .A1(n9714), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9715) );
  NAND2_X1 U12180 ( .A1(n11201), .A2(n13930), .ZN(n9717) );
  NAND3_X1 U12181 ( .A1(n14121), .A2(n10162), .A3(n10514), .ZN(n9731) );
  INV_X1 U12182 ( .A(n10516), .ZN(n9718) );
  NAND2_X1 U12183 ( .A1(n9880), .A2(n10342), .ZN(n11327) );
  OAI21_X1 U12184 ( .B1(n9880), .B2(n10342), .A(n12323), .ZN(n10509) );
  INV_X1 U12185 ( .A(n14290), .ZN(n11467) );
  OR2_X1 U12186 ( .A1(n10723), .A2(n10727), .ZN(n14543) );
  NAND2_X1 U12187 ( .A1(n14544), .A2(n10959), .ZN(n14523) );
  OR2_X1 U12188 ( .A1(n14523), .A2(n11040), .ZN(n14524) );
  INV_X1 U12189 ( .A(n11217), .ZN(n14609) );
  OR2_X1 U12190 ( .A1(n14636), .A2(n11312), .ZN(n11311) );
  NOR2_X2 U12191 ( .A1(n13821), .A2(n13827), .ZN(n13815) );
  NAND2_X1 U12192 ( .A1(n10061), .A2(n13815), .ZN(n13806) );
  OAI21_X1 U12193 ( .B1(n10061), .B2(n13815), .A(n13806), .ZN(n14026) );
  INV_X1 U12194 ( .A(n14026), .ZN(n9736) );
  NOR2_X1 U12195 ( .A1(n13902), .A2(n10341), .ZN(n14014) );
  INV_X1 U12196 ( .A(n11201), .ZN(n9759) );
  NAND2_X1 U12197 ( .A1(n9882), .A2(n9759), .ZN(n10111) );
  NOR2_X1 U12198 ( .A1(n9879), .A2(n10111), .ZN(n10360) );
  INV_X1 U12199 ( .A(n10360), .ZN(n10355) );
  NAND2_X1 U12200 ( .A1(n10357), .A2(n9721), .ZN(n14408) );
  INV_X1 U12201 ( .A(P1_B_REG_SCAN_IN), .ZN(n9723) );
  NOR2_X1 U12202 ( .A1(n14150), .A2(n9723), .ZN(n9724) );
  NOR2_X1 U12203 ( .A1(n14408), .A2(n9724), .ZN(n13802) );
  INV_X1 U12204 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9728) );
  NAND2_X1 U12205 ( .A1(n10049), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9727) );
  NAND2_X1 U12206 ( .A1(n9725), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n9726) );
  OAI211_X1 U12207 ( .C1(n9729), .C2(n9728), .A(n9727), .B(n9726), .ZN(n13662)
         );
  NAND2_X1 U12208 ( .A1(n13802), .A2(n13662), .ZN(n14025) );
  OAI22_X1 U12209 ( .A1(n9731), .A2(n14025), .B1(n9730), .B2(n13962), .ZN(
        n9733) );
  INV_X1 U12210 ( .A(n9721), .ZN(n10523) );
  OR2_X1 U12211 ( .A1(n14552), .A2(n14410), .ZN(n13849) );
  INV_X1 U12212 ( .A(n13663), .ZN(n14039) );
  NOR2_X1 U12213 ( .A1(n13849), .A2(n14039), .ZN(n9732) );
  AOI211_X1 U12214 ( .C1(n14539), .C2(P1_REG2_REG_29__SCAN_IN), .A(n9733), .B(
        n9732), .ZN(n9734) );
  OAI21_X1 U12215 ( .B1(n10061), .B2(n14541), .A(n9734), .ZN(n9735) );
  NAND2_X1 U12216 ( .A1(n9888), .A2(n9884), .ZN(n9738) );
  NAND2_X1 U12217 ( .A1(n9738), .A2(n9889), .ZN(n10718) );
  NAND2_X1 U12218 ( .A1(n9739), .A2(n10727), .ZN(n9740) );
  NAND2_X1 U12219 ( .A1(n10964), .A2(n6626), .ZN(n9741) );
  NAND2_X1 U12220 ( .A1(n9742), .A2(n9741), .ZN(n10888) );
  NAND2_X1 U12221 ( .A1(n10888), .A2(n10892), .ZN(n9744) );
  NAND2_X1 U12222 ( .A1(n14585), .A2(n11038), .ZN(n9743) );
  NAND2_X1 U12223 ( .A1(n9744), .A2(n9743), .ZN(n14515) );
  NAND2_X1 U12224 ( .A1(n14515), .A2(n7352), .ZN(n9746) );
  NAND2_X1 U12225 ( .A1(n11040), .A2(n10958), .ZN(n9745) );
  NAND2_X1 U12226 ( .A1(n9746), .A2(n9745), .ZN(n10899) );
  INV_X1 U12227 ( .A(n13670), .ZN(n11039) );
  AND2_X1 U12228 ( .A1(n11180), .A2(n11039), .ZN(n9747) );
  INV_X1 U12229 ( .A(n14616), .ZN(n11334) );
  INV_X1 U12230 ( .A(n10090), .ZN(n11155) );
  NAND2_X1 U12231 ( .A1(n11156), .A2(n11155), .ZN(n11154) );
  INV_X1 U12232 ( .A(n11678), .ZN(n14633) );
  OR2_X1 U12233 ( .A1(n14627), .A2(n14633), .ZN(n9748) );
  NAND2_X1 U12234 ( .A1(n14378), .A2(n7358), .ZN(n14377) );
  OR2_X1 U12235 ( .A1(n14383), .A2(n11792), .ZN(n9750) );
  INV_X1 U12236 ( .A(n14289), .ZN(n14411) );
  OR2_X1 U12237 ( .A1(n14310), .A2(n14411), .ZN(n9752) );
  NAND2_X1 U12238 ( .A1(n14301), .A2(n9752), .ZN(n11650) );
  NAND2_X1 U12239 ( .A1(n11650), .A2(n7262), .ZN(n11649) );
  NAND2_X1 U12240 ( .A1(n11649), .A2(n9959), .ZN(n14362) );
  INV_X1 U12241 ( .A(n11904), .ZN(n9753) );
  NAND2_X1 U12242 ( .A1(n12244), .A2(n13993), .ZN(n9754) );
  XNOR2_X1 U12243 ( .A(n14116), .B(n13584), .ZN(n13991) );
  OR2_X1 U12244 ( .A1(n14116), .A2(n13584), .ZN(n9969) );
  NAND2_X1 U12245 ( .A1(n13995), .A2(n9969), .ZN(n13975) );
  INV_X1 U12246 ( .A(n13959), .ZN(n14102) );
  XNOR2_X1 U12247 ( .A(n14110), .B(n14102), .ZN(n13972) );
  INV_X1 U12248 ( .A(n13972), .ZN(n13976) );
  NAND2_X1 U12249 ( .A1(n13985), .A2(n13959), .ZN(n9756) );
  INV_X1 U12250 ( .A(n13665), .ZN(n9986) );
  NAND2_X1 U12251 ( .A1(n14106), .A2(n9986), .ZN(n9987) );
  INV_X1 U12252 ( .A(n14103), .ZN(n13933) );
  NAND2_X1 U12253 ( .A1(n14096), .A2(n13933), .ZN(n9757) );
  NAND2_X1 U12254 ( .A1(n13938), .A2(n9757), .ZN(n13926) );
  OR2_X1 U12255 ( .A1(n14088), .A2(n13624), .ZN(n9758) );
  INV_X1 U12256 ( .A(n13664), .ZN(n14085) );
  INV_X1 U12257 ( .A(n13916), .ZN(n14077) );
  INV_X1 U12258 ( .A(n13871), .ZN(n13876) );
  INV_X1 U12259 ( .A(n14046), .ZN(n13873) );
  INV_X1 U12260 ( .A(n13821), .ZN(n14034) );
  NAND2_X1 U12261 ( .A1(n9879), .A2(n13944), .ZN(n9761) );
  NAND2_X1 U12262 ( .A1(n9719), .A2(n9759), .ZN(n9760) );
  NOR2_X1 U12263 ( .A1(n14029), .A2(n14539), .ZN(n9762) );
  NAND2_X1 U12264 ( .A1(n12595), .A2(n10980), .ZN(n9765) );
  NAND2_X1 U12265 ( .A1(n9765), .A2(n10875), .ZN(n9766) );
  NAND2_X2 U12266 ( .A1(n9767), .A2(n9766), .ZN(n9774) );
  NAND2_X1 U12267 ( .A1(n15064), .A2(n12335), .ZN(n9769) );
  XOR2_X1 U12268 ( .A(n9774), .B(n15057), .Z(n9768) );
  INV_X1 U12269 ( .A(n9771), .ZN(n9772) );
  XNOR2_X1 U12270 ( .A(n9773), .B(n15060), .ZN(n11045) );
  OAI22_X1 U12271 ( .A1(n11044), .A2(n11045), .B1(n15060), .B2(n9773), .ZN(
        n11239) );
  XNOR2_X1 U12272 ( .A(n11458), .B(n9774), .ZN(n9775) );
  XOR2_X1 U12273 ( .A(n15026), .B(n9775), .Z(n11275) );
  XNOR2_X1 U12274 ( .A(n15020), .B(n9774), .ZN(n9776) );
  XNOR2_X1 U12275 ( .A(n11495), .B(n9776), .ZN(n11342) );
  INV_X1 U12276 ( .A(n9776), .ZN(n9777) );
  XNOR2_X1 U12277 ( .A(n9778), .B(n9774), .ZN(n9779) );
  INV_X1 U12278 ( .A(n12503), .ZN(n15018) );
  XNOR2_X1 U12279 ( .A(n9779), .B(n12503), .ZN(n11493) );
  XNOR2_X1 U12280 ( .A(n11828), .B(n12335), .ZN(n11685) );
  INV_X1 U12281 ( .A(n15001), .ZN(n11763) );
  XNOR2_X1 U12282 ( .A(n11718), .B(n9774), .ZN(n9783) );
  XNOR2_X1 U12283 ( .A(n9783), .B(n11730), .ZN(n11761) );
  INV_X1 U12284 ( .A(n9783), .ZN(n9784) );
  NAND2_X1 U12285 ( .A1(n9784), .A2(n11730), .ZN(n9785) );
  XNOR2_X1 U12286 ( .A(n9786), .B(n9774), .ZN(n9787) );
  XNOR2_X1 U12287 ( .A(n9787), .B(n12360), .ZN(n11884) );
  INV_X1 U12288 ( .A(n9787), .ZN(n9789) );
  INV_X1 U12289 ( .A(n12360), .ZN(n9788) );
  NAND2_X1 U12290 ( .A1(n9789), .A2(n9788), .ZN(n9790) );
  XNOR2_X1 U12291 ( .A(n11819), .B(n9774), .ZN(n9791) );
  XNOR2_X1 U12292 ( .A(n9791), .B(n12502), .ZN(n12364) );
  NAND2_X1 U12293 ( .A1(n9791), .A2(n12502), .ZN(n9792) );
  XNOR2_X1 U12294 ( .A(n12335), .B(n12925), .ZN(n9793) );
  XNOR2_X1 U12295 ( .A(n14339), .B(n9774), .ZN(n12388) );
  NAND2_X1 U12296 ( .A1(n12388), .A2(n12455), .ZN(n9795) );
  OAI21_X1 U12297 ( .B1(n12450), .B2(n9793), .A(n9795), .ZN(n9798) );
  INV_X1 U12298 ( .A(n9793), .ZN(n12387) );
  NOR2_X1 U12299 ( .A1(n12387), .A2(n14333), .ZN(n9796) );
  INV_X1 U12300 ( .A(n12455), .ZN(n12814) );
  INV_X1 U12301 ( .A(n12388), .ZN(n9794) );
  AOI22_X1 U12302 ( .A1(n9796), .A2(n9795), .B1(n12814), .B2(n9794), .ZN(n9797) );
  XNOR2_X1 U12303 ( .A(n12922), .B(n9774), .ZN(n11918) );
  XNOR2_X1 U12304 ( .A(n12918), .B(n12335), .ZN(n11928) );
  INV_X1 U12305 ( .A(n12486), .ZN(n12815) );
  NOR2_X1 U12306 ( .A1(n11928), .A2(n12815), .ZN(n9800) );
  INV_X1 U12307 ( .A(n11928), .ZN(n9799) );
  XOR2_X1 U12308 ( .A(n9774), .B(n12484), .Z(n12481) );
  NOR2_X1 U12309 ( .A1(n12481), .A2(n12501), .ZN(n9802) );
  NAND2_X1 U12310 ( .A1(n12481), .A2(n12501), .ZN(n9801) );
  XNOR2_X1 U12311 ( .A(n12779), .B(n9774), .ZN(n9803) );
  XNOR2_X1 U12312 ( .A(n9803), .B(n10685), .ZN(n12409) );
  NAND2_X1 U12313 ( .A1(n12410), .A2(n12409), .ZN(n9805) );
  OR2_X1 U12314 ( .A1(n9803), .A2(n12792), .ZN(n9804) );
  NAND2_X1 U12315 ( .A1(n9805), .A2(n9804), .ZN(n12416) );
  XNOR2_X1 U12316 ( .A(n12860), .B(n9774), .ZN(n9806) );
  XNOR2_X1 U12317 ( .A(n9806), .B(n12500), .ZN(n12417) );
  XNOR2_X1 U12318 ( .A(n12751), .B(n9774), .ZN(n9808) );
  XNOR2_X1 U12319 ( .A(n9808), .B(n12734), .ZN(n12461) );
  XNOR2_X1 U12320 ( .A(n12901), .B(n9774), .ZN(n9809) );
  XNOR2_X1 U12321 ( .A(n12848), .B(n9774), .ZN(n9810) );
  INV_X1 U12322 ( .A(n9810), .ZN(n9811) );
  NAND2_X1 U12323 ( .A1(n9811), .A2(n12733), .ZN(n9812) );
  XNOR2_X1 U12324 ( .A(n12383), .B(n9774), .ZN(n9813) );
  NAND2_X1 U12325 ( .A1(n9813), .A2(n12700), .ZN(n9814) );
  OAI21_X1 U12326 ( .B1(n9813), .B2(n12700), .A(n9814), .ZN(n12379) );
  INV_X1 U12327 ( .A(n9818), .ZN(n9816) );
  XNOR2_X1 U12328 ( .A(n12447), .B(n9774), .ZN(n9817) );
  INV_X1 U12329 ( .A(n9817), .ZN(n9815) );
  NAND2_X1 U12330 ( .A1(n9816), .A2(n9815), .ZN(n9819) );
  NAND2_X1 U12331 ( .A1(n9818), .A2(n9817), .ZN(n9820) );
  INV_X1 U12332 ( .A(n9824), .ZN(n9822) );
  XNOR2_X1 U12333 ( .A(n12689), .B(n9774), .ZN(n9823) );
  INV_X1 U12334 ( .A(n9823), .ZN(n9821) );
  NAND2_X1 U12335 ( .A1(n9822), .A2(n9821), .ZN(n9825) );
  NAND2_X1 U12336 ( .A1(n9824), .A2(n9823), .ZN(n12424) );
  NAND2_X1 U12337 ( .A1(n9825), .A2(n12424), .ZN(n12354) );
  XNOR2_X1 U12338 ( .A(n12675), .B(n12335), .ZN(n9826) );
  NAND2_X1 U12339 ( .A1(n9826), .A2(n12405), .ZN(n12398) );
  INV_X1 U12340 ( .A(n9826), .ZN(n9827) );
  NAND2_X1 U12341 ( .A1(n9827), .A2(n12682), .ZN(n9828) );
  OR2_X1 U12342 ( .A1(n12668), .A2(n9830), .ZN(n9829) );
  NOR2_X1 U12343 ( .A1(n12354), .A2(n9829), .ZN(n9832) );
  NOR2_X1 U12344 ( .A1(n9830), .A2(n12424), .ZN(n9831) );
  NOR2_X1 U12345 ( .A1(n9832), .A2(n9831), .ZN(n12397) );
  NAND2_X1 U12346 ( .A1(n12397), .A2(n12398), .ZN(n9836) );
  XNOR2_X1 U12347 ( .A(n12396), .B(n9774), .ZN(n9833) );
  NAND2_X1 U12348 ( .A1(n9833), .A2(n12671), .ZN(n9837) );
  INV_X1 U12349 ( .A(n9833), .ZN(n9834) );
  NAND2_X1 U12350 ( .A1(n9834), .A2(n12475), .ZN(n9835) );
  XNOR2_X1 U12351 ( .A(n9838), .B(n12335), .ZN(n9839) );
  NOR2_X1 U12352 ( .A1(n9839), .A2(n12656), .ZN(n9840) );
  AOI21_X1 U12353 ( .B1(n9839), .B2(n12656), .A(n9840), .ZN(n12472) );
  INV_X1 U12354 ( .A(n9840), .ZN(n9841) );
  INV_X1 U12355 ( .A(n9846), .ZN(n9844) );
  XNOR2_X1 U12356 ( .A(n9842), .B(n12335), .ZN(n12343) );
  NOR2_X1 U12357 ( .A1(n12343), .A2(n12499), .ZN(n12338) );
  AOI21_X1 U12358 ( .B1(n12343), .B2(n12499), .A(n12338), .ZN(n9845) );
  INV_X1 U12359 ( .A(n9845), .ZN(n9843) );
  NAND2_X1 U12360 ( .A1(n9844), .A2(n9843), .ZN(n9847) );
  NAND2_X1 U12361 ( .A1(n9847), .A2(n12349), .ZN(n9849) );
  OAI22_X1 U12362 ( .A1(n9858), .A2(n11057), .B1(n9855), .B2(n9864), .ZN(n9848) );
  NAND2_X1 U12363 ( .A1(n9849), .A2(n12473), .ZN(n9873) );
  INV_X1 U12364 ( .A(n9858), .ZN(n9851) );
  AND2_X1 U12365 ( .A1(n10749), .A2(n14345), .ZN(n9850) );
  NAND2_X1 U12366 ( .A1(n9851), .A2(n9850), .ZN(n9853) );
  NOR2_X1 U12367 ( .A1(n9863), .A2(n9854), .ZN(n9862) );
  INV_X1 U12368 ( .A(n9864), .ZN(n9856) );
  OAI211_X1 U12369 ( .C1(n9856), .C2(n9855), .A(n11059), .B(n10119), .ZN(n9857) );
  AOI21_X1 U12370 ( .B1(n9859), .B2(n9858), .A(n9857), .ZN(n9860) );
  NOR2_X1 U12371 ( .A1(n9860), .A2(P3_U3151), .ZN(n9861) );
  AOI21_X1 U12372 ( .B1(n9862), .B2(n9864), .A(n9861), .ZN(n11047) );
  OR2_X1 U12373 ( .A1(n9864), .A2(n9863), .ZN(n9866) );
  INV_X1 U12374 ( .A(n9866), .ZN(n9865) );
  AOI22_X1 U12375 ( .A1(n12656), .A2(n12487), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n9867) );
  OAI21_X1 U12376 ( .B1(n9868), .B2(n12490), .A(n9867), .ZN(n9869) );
  AOI21_X1 U12377 ( .B1(n12637), .B2(n12493), .A(n9869), .ZN(n9870) );
  INV_X1 U12378 ( .A(n9871), .ZN(n9872) );
  NAND2_X1 U12379 ( .A1(n9873), .A2(n9872), .ZN(P3_U3154) );
  INV_X1 U12380 ( .A(n9879), .ZN(n10511) );
  NAND2_X1 U12381 ( .A1(n10511), .A2(n11201), .ZN(n9874) );
  NAND2_X1 U12382 ( .A1(n10175), .A2(n9874), .ZN(n9875) );
  OR2_X1 U12383 ( .A1(n10342), .A2(n13930), .ZN(n10717) );
  AND2_X1 U12384 ( .A1(n9875), .A2(n10717), .ZN(n10080) );
  INV_X1 U12385 ( .A(n10080), .ZN(n9876) );
  NAND2_X1 U12386 ( .A1(n9876), .A2(n10111), .ZN(n10081) );
  INV_X1 U12387 ( .A(n10081), .ZN(n10085) );
  NAND2_X1 U12388 ( .A1(n10709), .A2(n9877), .ZN(n9878) );
  NAND2_X1 U12389 ( .A1(n9884), .A2(n9878), .ZN(n14010) );
  OAI21_X2 U12390 ( .B1(n9883), .B2(n11201), .A(n10058), .ZN(n9904) );
  XNOR2_X1 U12391 ( .A(n9884), .B(n9899), .ZN(n9885) );
  OAI21_X1 U12392 ( .B1(n14010), .B2(n10342), .A(n9885), .ZN(n9887) );
  MUX2_X1 U12393 ( .A(n9888), .B(n9889), .S(n9899), .Z(n9886) );
  NAND2_X1 U12394 ( .A1(n9887), .A2(n9886), .ZN(n9893) );
  MUX2_X1 U12395 ( .A(n9889), .B(n9888), .S(n9899), .Z(n9891) );
  NAND2_X1 U12396 ( .A1(n9893), .A2(n9892), .ZN(n9898) );
  NAND2_X1 U12397 ( .A1(n9904), .A2(n10727), .ZN(n9896) );
  NAND2_X1 U12398 ( .A1(n9899), .A2(n14569), .ZN(n9895) );
  NAND2_X1 U12399 ( .A1(n9898), .A2(n7529), .ZN(n9903) );
  NAND2_X1 U12400 ( .A1(n10056), .A2(n14583), .ZN(n9901) );
  NAND2_X1 U12401 ( .A1(n9899), .A2(n10964), .ZN(n9900) );
  MUX2_X1 U12402 ( .A(n9901), .B(n9900), .S(n6626), .Z(n9902) );
  NAND2_X1 U12403 ( .A1(n9903), .A2(n9902), .ZN(n9907) );
  MUX2_X1 U12404 ( .A(n10959), .B(n11038), .S(n9899), .Z(n9906) );
  MUX2_X1 U12405 ( .A(n13671), .B(n14585), .S(n9899), .Z(n9905) );
  OAI21_X1 U12406 ( .B1(n9907), .B2(n9906), .A(n9905), .ZN(n9909) );
  NAND2_X1 U12407 ( .A1(n9907), .A2(n9906), .ZN(n9908) );
  NAND2_X1 U12408 ( .A1(n9909), .A2(n9908), .ZN(n9912) );
  MUX2_X1 U12409 ( .A(n14584), .B(n11040), .S(n9899), .Z(n9913) );
  NAND2_X1 U12410 ( .A1(n9912), .A2(n9913), .ZN(n9911) );
  MUX2_X1 U12411 ( .A(n11040), .B(n14584), .S(n9899), .Z(n9910) );
  NAND2_X1 U12412 ( .A1(n9911), .A2(n9910), .ZN(n9917) );
  INV_X1 U12413 ( .A(n9912), .ZN(n9915) );
  INV_X1 U12414 ( .A(n9913), .ZN(n9914) );
  NAND2_X1 U12415 ( .A1(n9915), .A2(n9914), .ZN(n9916) );
  NAND2_X1 U12416 ( .A1(n9917), .A2(n9916), .ZN(n9919) );
  MUX2_X1 U12417 ( .A(n11180), .B(n13670), .S(n9899), .Z(n9920) );
  MUX2_X1 U12418 ( .A(n11180), .B(n13670), .S(n10056), .Z(n9918) );
  INV_X1 U12419 ( .A(n9920), .ZN(n9921) );
  MUX2_X1 U12420 ( .A(n14616), .B(n11217), .S(n9899), .Z(n9925) );
  MUX2_X1 U12421 ( .A(n14616), .B(n11217), .S(n10056), .Z(n9922) );
  NAND2_X1 U12422 ( .A1(n9923), .A2(n9922), .ZN(n9928) );
  INV_X1 U12423 ( .A(n9924), .ZN(n9926) );
  NAND2_X1 U12424 ( .A1(n9926), .A2(n7226), .ZN(n9927) );
  NAND2_X1 U12425 ( .A1(n9928), .A2(n9927), .ZN(n9932) );
  MUX2_X1 U12426 ( .A(n9930), .B(n9929), .S(n9899), .Z(n9931) );
  NAND2_X1 U12427 ( .A1(n9932), .A2(n9931), .ZN(n9935) );
  MUX2_X1 U12428 ( .A(n11607), .B(n7219), .S(n9899), .Z(n9934) );
  MUX2_X1 U12429 ( .A(n11678), .B(n14627), .S(n9899), .Z(n9937) );
  MUX2_X1 U12430 ( .A(n14633), .B(n11162), .S(n10056), .Z(n9936) );
  MUX2_X1 U12431 ( .A(n13668), .B(n14636), .S(n10056), .Z(n9940) );
  MUX2_X1 U12432 ( .A(n13668), .B(n14636), .S(n9899), .Z(n9938) );
  NAND2_X1 U12433 ( .A1(n9939), .A2(n9938), .ZN(n9942) );
  NAND2_X1 U12434 ( .A1(n6701), .A2(n7247), .ZN(n9941) );
  MUX2_X1 U12435 ( .A(n14288), .B(n14383), .S(n9899), .Z(n9944) );
  MUX2_X1 U12436 ( .A(n14288), .B(n14383), .S(n10056), .Z(n9943) );
  INV_X1 U12437 ( .A(n9944), .ZN(n9945) );
  MUX2_X1 U12438 ( .A(n13667), .B(n14290), .S(n10056), .Z(n9949) );
  NAND2_X1 U12439 ( .A1(n9948), .A2(n9949), .ZN(n9947) );
  MUX2_X1 U12440 ( .A(n13667), .B(n14290), .S(n9899), .Z(n9946) );
  NAND2_X1 U12441 ( .A1(n9947), .A2(n9946), .ZN(n9953) );
  INV_X1 U12442 ( .A(n9948), .ZN(n9951) );
  INV_X1 U12443 ( .A(n9949), .ZN(n9950) );
  NAND2_X1 U12444 ( .A1(n9951), .A2(n9950), .ZN(n9952) );
  NAND2_X1 U12445 ( .A1(n9953), .A2(n9952), .ZN(n9955) );
  MUX2_X1 U12446 ( .A(n14289), .B(n14310), .S(n9899), .Z(n9956) );
  MUX2_X1 U12447 ( .A(n14289), .B(n14310), .S(n10056), .Z(n9954) );
  INV_X1 U12448 ( .A(n9956), .ZN(n9957) );
  NAND2_X1 U12449 ( .A1(n9963), .A2(n9958), .ZN(n9961) );
  NAND2_X1 U12450 ( .A1(n9962), .A2(n9959), .ZN(n9960) );
  MUX2_X1 U12451 ( .A(n9961), .B(n9960), .S(n9899), .Z(n9965) );
  MUX2_X1 U12452 ( .A(n9963), .B(n9962), .S(n10056), .Z(n9964) );
  INV_X1 U12453 ( .A(n12244), .ZN(n14397) );
  MUX2_X1 U12454 ( .A(n13993), .B(n14397), .S(n9899), .Z(n9975) );
  NAND2_X1 U12455 ( .A1(n12244), .A2(n10056), .ZN(n9968) );
  NAND2_X1 U12456 ( .A1(n14116), .A2(n13584), .ZN(n9967) );
  NAND2_X1 U12457 ( .A1(n9899), .A2(n13666), .ZN(n9966) );
  NAND4_X1 U12458 ( .A1(n9969), .A2(n9968), .A3(n9967), .A4(n9966), .ZN(n9976)
         );
  OAI21_X1 U12459 ( .B1(n13991), .B2(n9975), .A(n9976), .ZN(n9970) );
  NAND2_X1 U12460 ( .A1(n9971), .A2(n9970), .ZN(n9979) );
  AND2_X1 U12461 ( .A1(n14394), .A2(n10056), .ZN(n9973) );
  OAI21_X1 U12462 ( .B1(n14394), .B2(n10056), .A(n14116), .ZN(n9972) );
  OAI21_X1 U12463 ( .B1(n9973), .B2(n14116), .A(n9972), .ZN(n9974) );
  OAI21_X1 U12464 ( .B1(n9976), .B2(n9975), .A(n9974), .ZN(n9977) );
  INV_X1 U12465 ( .A(n9977), .ZN(n9978) );
  NAND2_X1 U12466 ( .A1(n9979), .A2(n9978), .ZN(n9982) );
  INV_X1 U12467 ( .A(n9982), .ZN(n9985) );
  MUX2_X1 U12468 ( .A(n14102), .B(n13985), .S(n10056), .Z(n9980) );
  OAI211_X1 U12469 ( .C1(n9985), .C2(n9984), .A(n9983), .B(n13954), .ZN(n9990)
         );
  OR2_X1 U12470 ( .A1(n14106), .A2(n9986), .ZN(n9988) );
  MUX2_X1 U12471 ( .A(n9988), .B(n9987), .S(n10056), .Z(n9989) );
  MUX2_X1 U12472 ( .A(n14103), .B(n14096), .S(n9899), .Z(n9992) );
  MUX2_X1 U12473 ( .A(n13933), .B(n13946), .S(n10056), .Z(n9991) );
  MUX2_X1 U12474 ( .A(n14076), .B(n14088), .S(n10056), .Z(n9995) );
  MUX2_X1 U12475 ( .A(n14076), .B(n14088), .S(n9899), .Z(n9993) );
  NAND2_X1 U12476 ( .A1(n9994), .A2(n9993), .ZN(n9997) );
  NAND2_X1 U12477 ( .A1(n6702), .A2(n7240), .ZN(n9996) );
  MUX2_X1 U12478 ( .A(n13664), .B(n13913), .S(n9899), .Z(n9999) );
  MUX2_X1 U12479 ( .A(n13664), .B(n13913), .S(n10056), .Z(n9998) );
  INV_X1 U12480 ( .A(n9999), .ZN(n10000) );
  MUX2_X1 U12481 ( .A(n13916), .B(n14071), .S(n9899), .Z(n10004) );
  NAND2_X1 U12482 ( .A1(n10003), .A2(n10004), .ZN(n10002) );
  MUX2_X1 U12483 ( .A(n13916), .B(n14071), .S(n10056), .Z(n10001) );
  NAND2_X1 U12484 ( .A1(n10002), .A2(n10001), .ZN(n10008) );
  INV_X1 U12485 ( .A(n10003), .ZN(n10006) );
  INV_X1 U12486 ( .A(n10004), .ZN(n10005) );
  NAND2_X1 U12487 ( .A1(n10006), .A2(n10005), .ZN(n10007) );
  MUX2_X1 U12488 ( .A(n14066), .B(n13860), .S(n9904), .Z(n10010) );
  MUX2_X1 U12489 ( .A(n14066), .B(n13860), .S(n9899), .Z(n10009) );
  INV_X1 U12490 ( .A(n10010), .ZN(n10011) );
  MUX2_X1 U12491 ( .A(n14046), .B(n14057), .S(n9904), .Z(n10015) );
  NAND2_X1 U12492 ( .A1(n10014), .A2(n10015), .ZN(n10013) );
  MUX2_X1 U12493 ( .A(n14046), .B(n14057), .S(n9899), .Z(n10012) );
  NAND2_X1 U12494 ( .A1(n10013), .A2(n10012), .ZN(n10019) );
  INV_X1 U12495 ( .A(n10014), .ZN(n10017) );
  INV_X1 U12496 ( .A(n10015), .ZN(n10016) );
  NAND2_X1 U12497 ( .A1(n10017), .A2(n10016), .ZN(n10018) );
  MUX2_X1 U12498 ( .A(n13859), .B(n13851), .S(n9899), .Z(n10021) );
  MUX2_X1 U12499 ( .A(n13851), .B(n13859), .S(n9899), .Z(n10020) );
  MUX2_X1 U12500 ( .A(n14047), .B(n14042), .S(n9904), .Z(n10025) );
  NAND2_X1 U12501 ( .A1(n10024), .A2(n10025), .ZN(n10023) );
  MUX2_X1 U12502 ( .A(n14047), .B(n14042), .S(n9899), .Z(n10022) );
  NAND2_X1 U12503 ( .A1(n10023), .A2(n10022), .ZN(n10029) );
  INV_X1 U12504 ( .A(n10024), .ZN(n10027) );
  INV_X1 U12505 ( .A(n10025), .ZN(n10026) );
  NAND2_X1 U12506 ( .A1(n10027), .A2(n10026), .ZN(n10028) );
  NAND2_X1 U12507 ( .A1(n10029), .A2(n10028), .ZN(n10032) );
  MUX2_X1 U12508 ( .A(n13663), .B(n13821), .S(n9899), .Z(n10033) );
  NAND2_X1 U12509 ( .A1(n10032), .A2(n10033), .ZN(n10031) );
  MUX2_X1 U12510 ( .A(n13663), .B(n13821), .S(n9904), .Z(n10030) );
  NAND2_X1 U12511 ( .A1(n10031), .A2(n10030), .ZN(n10037) );
  INV_X1 U12512 ( .A(n10032), .ZN(n10035) );
  INV_X1 U12513 ( .A(n10033), .ZN(n10034) );
  NAND2_X1 U12514 ( .A1(n10035), .A2(n10034), .ZN(n10036) );
  NAND2_X1 U12515 ( .A1(n10037), .A2(n10036), .ZN(n10064) );
  MUX2_X1 U12516 ( .A(n14031), .B(n14028), .S(n9904), .Z(n10063) );
  NAND2_X1 U12517 ( .A1(n10040), .A2(n12939), .ZN(n10041) );
  NAND2_X1 U12518 ( .A1(n10042), .A2(SI_30_), .ZN(n10065) );
  OAI21_X1 U12519 ( .B1(n10042), .B2(SI_30_), .A(n10065), .ZN(n10043) );
  NAND2_X1 U12520 ( .A1(n10044), .A2(n10043), .ZN(n10045) );
  OR2_X1 U12521 ( .A1(n6623), .A2(n9100), .ZN(n10047) );
  INV_X1 U12522 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n15333) );
  NAND2_X1 U12523 ( .A1(n10049), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n10052) );
  NAND2_X1 U12524 ( .A1(n10050), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n10051) );
  OAI211_X1 U12525 ( .C1(n10053), .C2(n15333), .A(n10052), .B(n10051), .ZN(
        n13801) );
  OAI21_X1 U12526 ( .B1(n13801), .B2(n11201), .A(n13662), .ZN(n10054) );
  INV_X1 U12527 ( .A(n10054), .ZN(n10055) );
  MUX2_X1 U12528 ( .A(n13808), .B(n10055), .S(n9899), .Z(n10075) );
  NAND2_X1 U12529 ( .A1(n10056), .A2(n13801), .ZN(n10059) );
  INV_X1 U12530 ( .A(n13662), .ZN(n10057) );
  AOI21_X1 U12531 ( .B1(n10059), .B2(n10058), .A(n10057), .ZN(n10060) );
  AOI21_X1 U12532 ( .B1(n13808), .B2(n9899), .A(n10060), .ZN(n10074) );
  INV_X1 U12533 ( .A(n14031), .ZN(n13816) );
  MUX2_X1 U12534 ( .A(n13816), .B(n10061), .S(n9899), .Z(n10062) );
  MUX2_X1 U12535 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7311), .Z(n10068) );
  XNOR2_X1 U12536 ( .A(n10068), .B(SI_31_), .ZN(n10069) );
  NAND2_X1 U12537 ( .A1(n13475), .A2(n10071), .ZN(n10073) );
  OR2_X1 U12538 ( .A1(n6623), .A2(n15239), .ZN(n10072) );
  XNOR2_X1 U12539 ( .A(n14019), .B(n13801), .ZN(n10108) );
  NAND2_X1 U12540 ( .A1(n10075), .A2(n10074), .ZN(n10076) );
  NAND2_X1 U12541 ( .A1(n9899), .A2(n13801), .ZN(n10079) );
  INV_X1 U12542 ( .A(n13801), .ZN(n10077) );
  NAND2_X1 U12543 ( .A1(n9904), .A2(n10077), .ZN(n10078) );
  MUX2_X1 U12544 ( .A(n10079), .B(n10078), .S(n14019), .Z(n10082) );
  AND2_X1 U12545 ( .A1(n10366), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10174) );
  XOR2_X1 U12546 ( .A(n13662), .B(n13808), .Z(n10106) );
  NOR2_X1 U12547 ( .A1(n10707), .A2(n14010), .ZN(n10087) );
  NAND4_X1 U12548 ( .A1(n10087), .A2(n10892), .A3(n10086), .A4(n9890), .ZN(
        n10088) );
  NOR2_X1 U12549 ( .A1(n10088), .A2(n14516), .ZN(n10089) );
  NAND4_X1 U12550 ( .A1(n11103), .A2(n10089), .A3(n14502), .A4(n10897), .ZN(
        n10091) );
  OR3_X1 U12551 ( .A1(n11310), .A2(n10091), .A3(n10090), .ZN(n10093) );
  OR3_X1 U12552 ( .A1(n10093), .A2(n10092), .A3(n14384), .ZN(n10094) );
  NOR2_X1 U12553 ( .A1(n10095), .A2(n10094), .ZN(n10096) );
  NAND4_X1 U12554 ( .A1(n14367), .A2(n9755), .A3(n10096), .A4(n14302), .ZN(
        n10097) );
  OR4_X1 U12555 ( .A1(n10098), .A2(n13972), .A3(n11904), .A4(n10097), .ZN(
        n10099) );
  OR4_X1 U12556 ( .A1(n13906), .A2(n10101), .A3(n10100), .A4(n10099), .ZN(
        n10102) );
  NOR2_X1 U12557 ( .A1(n13892), .A2(n10102), .ZN(n10103) );
  NAND4_X1 U12558 ( .A1(n13841), .A2(n10103), .A3(n13868), .A4(n13871), .ZN(
        n10104) );
  NOR4_X1 U12559 ( .A1(n10106), .A2(n10105), .A3(n13813), .A4(n10104), .ZN(
        n10109) );
  NAND3_X1 U12560 ( .A1(n10109), .A2(n10108), .A3(n10107), .ZN(n10110) );
  INV_X1 U12561 ( .A(n10111), .ZN(n10112) );
  NAND2_X1 U12562 ( .A1(n10114), .A2(n10113), .ZN(n10117) );
  INV_X1 U12563 ( .A(n10174), .ZN(n11775) );
  INV_X1 U12564 ( .A(n14150), .ZN(n14466) );
  NAND4_X1 U12565 ( .A1(n14634), .A2(n10515), .A3(n14466), .A4(n10514), .ZN(
        n10115) );
  OAI211_X1 U12566 ( .C1(n9879), .C2(n11775), .A(n10115), .B(P1_B_REG_SCAN_IN), 
        .ZN(n10116) );
  NAND2_X1 U12567 ( .A1(n10117), .A2(n10116), .ZN(P1_U3242) );
  INV_X1 U12568 ( .A(n10184), .ZN(n10118) );
  NAND2_X1 U12569 ( .A1(n10118), .A2(n11770), .ZN(n10182) );
  NOR2_X4 U12570 ( .A1(n10119), .A2(n11938), .ZN(P3_U3897) );
  NOR2_X4 U12571 ( .A1(n10366), .A2(n10120), .ZN(P1_U4016) );
  AND2_X1 U12572 ( .A1(n7572), .A2(P2_U3088), .ZN(n13492) );
  INV_X2 U12573 ( .A(n13492), .ZN(n13505) );
  AND2_X1 U12574 ( .A1(n10067), .A2(P2_U3088), .ZN(n13481) );
  INV_X2 U12575 ( .A(n13481), .ZN(n13498) );
  OAI222_X1 U12576 ( .A1(n13505), .A2(n10129), .B1(n13498), .B2(n10121), .C1(
        P2_U3088), .C2(n10210), .ZN(P2_U3326) );
  INV_X1 U12577 ( .A(n10242), .ZN(n10220) );
  OAI222_X1 U12578 ( .A1(n13498), .A2(n10122), .B1(n13505), .B2(n10127), .C1(
        n10220), .C2(P2_U3088), .ZN(P2_U3325) );
  AOI22_X1 U12579 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n13481), .B1(n14679), 
        .B2(P2_STATE_REG_SCAN_IN), .ZN(n10123) );
  OAI21_X1 U12580 ( .B1(n10124), .B2(n13505), .A(n10123), .ZN(P2_U3324) );
  OAI222_X1 U12581 ( .A1(n7001), .A2(n10125), .B1(n14160), .B2(n10124), .C1(
        n13705), .C2(P1_U3086), .ZN(P1_U3352) );
  INV_X1 U12582 ( .A(n14160), .ZN(n11773) );
  OAI222_X1 U12583 ( .A1(P1_U3086), .A2(n13690), .B1(n14160), .B2(n10127), 
        .C1(n10126), .C2(n7001), .ZN(P1_U3353) );
  OAI222_X1 U12584 ( .A1(P1_U3086), .A2(n10431), .B1(n14160), .B2(n10129), 
        .C1(n10128), .C2(n7001), .ZN(P1_U3354) );
  AND2_X1 U12585 ( .A1(n10067), .A2(P3_U3151), .ZN(n12933) );
  INV_X1 U12586 ( .A(n10130), .ZN(n10131) );
  INV_X1 U12587 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10803) );
  OAI222_X1 U12588 ( .A1(n12944), .A2(n10132), .B1(n11943), .B2(n10131), .C1(
        P3_U3151), .C2(n10803), .ZN(P3_U3295) );
  INV_X1 U12589 ( .A(SI_2_), .ZN(n15232) );
  OAI222_X1 U12590 ( .A1(n7599), .A2(P3_U3151), .B1(n11943), .B2(n10133), .C1(
        n15232), .C2(n12944), .ZN(P3_U3293) );
  INV_X1 U12591 ( .A(n14849), .ZN(n11426) );
  OAI222_X1 U12592 ( .A1(n11426), .A2(P3_U3151), .B1(n11943), .B2(n10135), 
        .C1(n10134), .C2(n12944), .ZN(P3_U3292) );
  INV_X1 U12593 ( .A(n11430), .ZN(n14875) );
  OAI222_X1 U12594 ( .A1(n14875), .A2(P3_U3151), .B1(n11943), .B2(n10137), 
        .C1(n10136), .C2(n12944), .ZN(P3_U3291) );
  OAI222_X1 U12595 ( .A1(n11431), .A2(P3_U3151), .B1(n11943), .B2(n10139), 
        .C1(n10138), .C2(n12944), .ZN(P3_U3290) );
  INV_X1 U12596 ( .A(n10140), .ZN(n10143) );
  OAI222_X1 U12597 ( .A1(n13498), .A2(n10141), .B1(n13505), .B2(n10143), .C1(
        n13115), .C2(P2_U3088), .ZN(P2_U3323) );
  INV_X1 U12598 ( .A(n10539), .ZN(n10142) );
  OAI222_X1 U12599 ( .A1(n7001), .A2(n6999), .B1(n14160), .B2(n10143), .C1(
        n10142), .C2(P1_U3086), .ZN(P1_U3351) );
  INV_X1 U12600 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10145) );
  INV_X1 U12601 ( .A(n13722), .ZN(n10144) );
  OAI222_X1 U12602 ( .A1(n7001), .A2(n10145), .B1(n14160), .B2(n10146), .C1(
        n10144), .C2(P1_U3086), .ZN(P1_U3350) );
  INV_X1 U12603 ( .A(n10276), .ZN(n10283) );
  OAI222_X1 U12604 ( .A1(n13498), .A2(n10147), .B1(n13505), .B2(n10146), .C1(
        n10283), .C2(P2_U3088), .ZN(P2_U3322) );
  OAI222_X1 U12605 ( .A1(P3_U3151), .A2(n14963), .B1(n12944), .B2(n10149), 
        .C1(n11943), .C2(n10148), .ZN(P3_U3286) );
  OAI222_X1 U12606 ( .A1(P3_U3151), .A2(n11528), .B1(n12944), .B2(n10151), 
        .C1(n11943), .C2(n10150), .ZN(P3_U3284) );
  INV_X1 U12607 ( .A(n10152), .ZN(n10154) );
  OAI222_X1 U12608 ( .A1(n11943), .A2(n10154), .B1(n12944), .B2(n10153), .C1(
        P3_U3151), .C2(n14942), .ZN(P3_U3287) );
  OAI222_X1 U12609 ( .A1(P3_U3151), .A2(n14927), .B1(n12944), .B2(n10156), 
        .C1(n11943), .C2(n10155), .ZN(P3_U3288) );
  INV_X1 U12610 ( .A(n11441), .ZN(n14981) );
  OAI222_X1 U12611 ( .A1(P3_U3151), .A2(n14981), .B1(n12944), .B2(n10158), 
        .C1(n11943), .C2(n10157), .ZN(P3_U3285) );
  INV_X1 U12612 ( .A(n10159), .ZN(n10161) );
  OAI222_X1 U12613 ( .A1(n11943), .A2(n10161), .B1(n12944), .B2(n10160), .C1(
        P3_U3151), .C2(n10774), .ZN(P3_U3294) );
  INV_X1 U12614 ( .A(n10162), .ZN(n10163) );
  OAI21_X1 U12615 ( .B1(n10515), .B2(n10164), .A(n10163), .ZN(P1_U3446) );
  INV_X1 U12616 ( .A(n10165), .ZN(n10166) );
  OAI222_X1 U12617 ( .A1(P3_U3151), .A2(n11424), .B1(n11943), .B2(n10166), 
        .C1(n15288), .C2(n12944), .ZN(P3_U3289) );
  INV_X1 U12618 ( .A(n10167), .ZN(n10168) );
  OAI222_X1 U12619 ( .A1(n12944), .A2(n10169), .B1(n11943), .B2(n10168), .C1(
        n11586), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U12620 ( .A(n13737), .ZN(n10170) );
  OAI222_X1 U12621 ( .A1(n7001), .A2(n10171), .B1(n14160), .B2(n10172), .C1(
        n10170), .C2(P1_U3086), .ZN(P1_U3349) );
  INV_X1 U12622 ( .A(n10263), .ZN(n10269) );
  OAI222_X1 U12623 ( .A1(n13498), .A2(n10173), .B1(n13505), .B2(n10172), .C1(
        n10269), .C2(P2_U3088), .ZN(P2_U3321) );
  OR2_X1 U12624 ( .A1(n10515), .A2(n10174), .ZN(n10424) );
  OR2_X1 U12625 ( .A1(n10175), .A2(n10366), .ZN(n10177) );
  NAND2_X1 U12626 ( .A1(n10177), .A2(n6772), .ZN(n10423) );
  AND2_X1 U12627 ( .A1(n10424), .A2(n10423), .ZN(n14468) );
  NOR2_X1 U12628 ( .A1(n14468), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12629 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10178) );
  INV_X1 U12630 ( .A(n10291), .ZN(n10299) );
  OAI222_X1 U12631 ( .A1(n13498), .A2(n10178), .B1(n13505), .B2(n10179), .C1(
        n10299), .C2(P2_U3088), .ZN(P2_U3320) );
  INV_X1 U12632 ( .A(n10476), .ZN(n10489) );
  OAI222_X1 U12633 ( .A1(n7001), .A2(n10180), .B1(n14160), .B2(n10179), .C1(
        n10489), .C2(P1_U3086), .ZN(P1_U3348) );
  NAND2_X1 U12634 ( .A1(n10182), .A2(n10181), .ZN(n10186) );
  NAND3_X1 U12635 ( .A1(n10184), .A2(n10183), .A3(n11770), .ZN(n10185) );
  NAND2_X1 U12636 ( .A1(n10186), .A2(n10185), .ZN(n10199) );
  NOR2_X1 U12637 ( .A1(n10199), .A2(P2_U3088), .ZN(n10194) );
  NOR2_X1 U12638 ( .A1(n13491), .A2(n10188), .ZN(n10187) );
  NAND2_X1 U12639 ( .A1(n10194), .A2(n10187), .ZN(n14718) );
  INV_X1 U12640 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10192) );
  INV_X1 U12641 ( .A(n10199), .ZN(n10190) );
  NAND2_X1 U12642 ( .A1(n10188), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13493) );
  NOR2_X1 U12643 ( .A1(n13493), .A2(n13491), .ZN(n10189) );
  NAND2_X1 U12644 ( .A1(n14729), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10191) );
  OAI21_X1 U12645 ( .B1(n14718), .B2(n10192), .A(n10191), .ZN(n10197) );
  INV_X1 U12646 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10193) );
  NAND2_X1 U12647 ( .A1(n14729), .A2(n10193), .ZN(n10195) );
  NAND2_X1 U12648 ( .A1(n10194), .A2(n13491), .ZN(n14722) );
  OAI211_X1 U12649 ( .C1(n14718), .C2(P2_REG1_REG_0__SCAN_IN), .A(n10195), .B(
        n14722), .ZN(n10196) );
  MUX2_X1 U12650 ( .A(n10197), .B(n10196), .S(n13507), .Z(n10198) );
  INV_X1 U12651 ( .A(n10198), .ZN(n10201) );
  AND2_X1 U12652 ( .A1(n10199), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14726) );
  AOI22_X1 U12653 ( .A1(n14726), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n10200) );
  NAND2_X1 U12654 ( .A1(n10201), .A2(n10200), .ZN(P2_U3214) );
  INV_X1 U12655 ( .A(n15133), .ZN(n14555) );
  NAND3_X1 U12656 ( .A1(n14158), .A2(P1_STATE_REG_SCAN_IN), .A3(n14152), .ZN(
        n10203) );
  OAI22_X1 U12657 ( .A1(n14555), .A2(P1_D_REG_0__SCAN_IN), .B1(n10366), .B2(
        n10203), .ZN(n10204) );
  INV_X1 U12658 ( .A(n10204), .ZN(P1_U3445) );
  NAND2_X1 U12659 ( .A1(n14667), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10206) );
  INV_X1 U12660 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10743) );
  NAND2_X1 U12661 ( .A1(n10210), .A2(n10743), .ZN(n10205) );
  AND2_X1 U12662 ( .A1(n10206), .A2(n10205), .ZN(n14673) );
  AND2_X1 U12663 ( .A1(n13507), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n14672) );
  NAND2_X1 U12664 ( .A1(n14673), .A2(n14672), .ZN(n14671) );
  NAND2_X1 U12665 ( .A1(n14671), .A2(n10206), .ZN(n10241) );
  INV_X1 U12666 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10207) );
  XNOR2_X1 U12667 ( .A(n10242), .B(n10207), .ZN(n10240) );
  XNOR2_X1 U12668 ( .A(n10241), .B(n10240), .ZN(n10208) );
  OAI22_X1 U12669 ( .A1(n14745), .A2(n10208), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6767), .ZN(n10209) );
  AOI21_X1 U12670 ( .B1(n14726), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n10209), .ZN(
        n10219) );
  INV_X1 U12671 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10211) );
  MUX2_X1 U12672 ( .A(n10211), .B(P2_REG1_REG_1__SCAN_IN), .S(n10210), .Z(
        n14669) );
  AND2_X1 U12673 ( .A1(n13507), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n14670) );
  NAND2_X1 U12674 ( .A1(n14669), .A2(n14670), .ZN(n14668) );
  NAND2_X1 U12675 ( .A1(n14667), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10216) );
  NAND2_X1 U12676 ( .A1(n14668), .A2(n10216), .ZN(n10214) );
  INV_X1 U12677 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10212) );
  MUX2_X1 U12678 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10212), .S(n10242), .Z(
        n10213) );
  NAND2_X1 U12679 ( .A1(n10214), .A2(n10213), .ZN(n10222) );
  MUX2_X1 U12680 ( .A(n10212), .B(P2_REG1_REG_2__SCAN_IN), .S(n10242), .Z(
        n10215) );
  NAND3_X1 U12681 ( .A1(n14668), .A2(n10216), .A3(n10215), .ZN(n10217) );
  NAND3_X1 U12682 ( .A1(n14752), .A2(n10222), .A3(n10217), .ZN(n10218) );
  OAI211_X1 U12683 ( .C1(n14722), .C2(n10220), .A(n10219), .B(n10218), .ZN(
        P2_U3216) );
  NAND2_X1 U12684 ( .A1(n10242), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10221) );
  NAND2_X1 U12685 ( .A1(n10222), .A2(n10221), .ZN(n14682) );
  INV_X1 U12686 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10223) );
  MUX2_X1 U12687 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10223), .S(n14679), .Z(
        n14681) );
  NAND2_X1 U12688 ( .A1(n14682), .A2(n14681), .ZN(n14680) );
  NAND2_X1 U12689 ( .A1(n14679), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n13116) );
  NAND2_X1 U12690 ( .A1(n14680), .A2(n13116), .ZN(n10226) );
  INV_X1 U12691 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10224) );
  MUX2_X1 U12692 ( .A(n10224), .B(P2_REG1_REG_4__SCAN_IN), .S(n13115), .Z(
        n10225) );
  NAND2_X1 U12693 ( .A1(n10226), .A2(n10225), .ZN(n13119) );
  NAND2_X1 U12694 ( .A1(n13121), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10278) );
  NAND2_X1 U12695 ( .A1(n13119), .A2(n10278), .ZN(n10229) );
  INV_X1 U12696 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10227) );
  MUX2_X1 U12697 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10227), .S(n10276), .Z(
        n10228) );
  NAND2_X1 U12698 ( .A1(n10229), .A2(n10228), .ZN(n10280) );
  NAND2_X1 U12699 ( .A1(n10276), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10265) );
  NAND2_X1 U12700 ( .A1(n10280), .A2(n10265), .ZN(n10232) );
  INV_X1 U12701 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10230) );
  MUX2_X1 U12702 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10230), .S(n10263), .Z(
        n10231) );
  NAND2_X1 U12703 ( .A1(n10232), .A2(n10231), .ZN(n10294) );
  NAND2_X1 U12704 ( .A1(n10263), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10293) );
  NAND2_X1 U12705 ( .A1(n10294), .A2(n10293), .ZN(n10235) );
  INV_X1 U12706 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10233) );
  MUX2_X1 U12707 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10233), .S(n10291), .Z(
        n10234) );
  NAND2_X1 U12708 ( .A1(n10235), .A2(n10234), .ZN(n10296) );
  NAND2_X1 U12709 ( .A1(n10291), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10237) );
  INV_X1 U12710 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10938) );
  MUX2_X1 U12711 ( .A(n10938), .B(P2_REG1_REG_8__SCAN_IN), .S(n10309), .Z(
        n10236) );
  AOI21_X1 U12712 ( .B1(n10296), .B2(n10237), .A(n10236), .ZN(n10305) );
  NAND3_X1 U12713 ( .A1(n10296), .A2(n10237), .A3(n10236), .ZN(n10238) );
  NAND2_X1 U12714 ( .A1(n14752), .A2(n10238), .ZN(n10256) );
  INV_X1 U12715 ( .A(n14722), .ZN(n14750) );
  INV_X1 U12716 ( .A(n14726), .ZN(n14741) );
  INV_X1 U12717 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10239) );
  NAND2_X1 U12718 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n10832) );
  OAI21_X1 U12719 ( .B1(n14741), .B2(n10239), .A(n10832), .ZN(n10254) );
  NAND2_X1 U12720 ( .A1(n10241), .A2(n10240), .ZN(n10244) );
  NAND2_X1 U12721 ( .A1(n10242), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10243) );
  NAND2_X1 U12722 ( .A1(n10244), .A2(n10243), .ZN(n14685) );
  INV_X1 U12723 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10245) );
  MUX2_X1 U12724 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10245), .S(n14679), .Z(
        n14684) );
  NAND2_X1 U12725 ( .A1(n14685), .A2(n14684), .ZN(n14683) );
  NAND2_X1 U12726 ( .A1(n14679), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n13124) );
  INV_X1 U12727 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10246) );
  MUX2_X1 U12728 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10246), .S(n13115), .Z(
        n13123) );
  AOI21_X1 U12729 ( .B1(n14683), .B2(n13124), .A(n13123), .ZN(n13122) );
  NOR2_X1 U12730 ( .A1(n13115), .A2(n10246), .ZN(n10272) );
  INV_X1 U12731 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10972) );
  MUX2_X1 U12732 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10972), .S(n10276), .Z(
        n10271) );
  OAI21_X1 U12733 ( .B1(n13122), .B2(n10272), .A(n10271), .ZN(n10270) );
  NAND2_X1 U12734 ( .A1(n10276), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10259) );
  INV_X1 U12735 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10247) );
  MUX2_X1 U12736 ( .A(n10247), .B(P2_REG2_REG_6__SCAN_IN), .S(n10263), .Z(
        n10258) );
  AOI21_X1 U12737 ( .B1(n10270), .B2(n10259), .A(n10258), .ZN(n10287) );
  NOR2_X1 U12738 ( .A1(n10269), .A2(n10247), .ZN(n10286) );
  INV_X1 U12739 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10248) );
  MUX2_X1 U12740 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10248), .S(n10291), .Z(
        n10285) );
  OAI21_X1 U12741 ( .B1(n10287), .B2(n10286), .A(n10285), .ZN(n10284) );
  NAND2_X1 U12742 ( .A1(n10291), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10251) );
  INV_X1 U12743 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10249) );
  MUX2_X1 U12744 ( .A(n10249), .B(P2_REG2_REG_8__SCAN_IN), .S(n10309), .Z(
        n10250) );
  AOI21_X1 U12745 ( .B1(n10284), .B2(n10251), .A(n10250), .ZN(n10308) );
  AND3_X1 U12746 ( .A1(n10284), .A2(n10251), .A3(n10250), .ZN(n10252) );
  NOR3_X1 U12747 ( .A1(n14745), .A2(n10308), .A3(n10252), .ZN(n10253) );
  AOI211_X1 U12748 ( .C1(n14750), .C2(n10309), .A(n10254), .B(n10253), .ZN(
        n10255) );
  OAI21_X1 U12749 ( .B1(n10305), .B2(n10256), .A(n10255), .ZN(P2_U3222) );
  AOI22_X1 U12750 ( .A1(n10544), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n14141), .ZN(n10257) );
  OAI21_X1 U12751 ( .B1(n10303), .B2(n14160), .A(n10257), .ZN(P1_U3347) );
  NAND2_X1 U12752 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10675) );
  INV_X1 U12753 ( .A(n10675), .ZN(n10262) );
  AND3_X1 U12754 ( .A1(n10270), .A2(n10259), .A3(n10258), .ZN(n10260) );
  NOR3_X1 U12755 ( .A1(n14745), .A2(n10287), .A3(n10260), .ZN(n10261) );
  AOI211_X1 U12756 ( .C1(n14726), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n10262), .B(
        n10261), .ZN(n10268) );
  MUX2_X1 U12757 ( .A(n10230), .B(P2_REG1_REG_6__SCAN_IN), .S(n10263), .Z(
        n10264) );
  NAND3_X1 U12758 ( .A1(n10280), .A2(n10265), .A3(n10264), .ZN(n10266) );
  NAND3_X1 U12759 ( .A1(n14752), .A2(n10294), .A3(n10266), .ZN(n10267) );
  OAI211_X1 U12760 ( .C1(n14722), .C2(n10269), .A(n10268), .B(n10267), .ZN(
        P2_U3220) );
  AND2_X1 U12761 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10634) );
  INV_X1 U12762 ( .A(n10270), .ZN(n10274) );
  NOR3_X1 U12763 ( .A1(n13122), .A2(n10272), .A3(n10271), .ZN(n10273) );
  NOR3_X1 U12764 ( .A1(n14745), .A2(n10274), .A3(n10273), .ZN(n10275) );
  AOI211_X1 U12765 ( .C1(n14726), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n10634), .B(
        n10275), .ZN(n10282) );
  MUX2_X1 U12766 ( .A(n10227), .B(P2_REG1_REG_5__SCAN_IN), .S(n10276), .Z(
        n10277) );
  NAND3_X1 U12767 ( .A1(n13119), .A2(n10278), .A3(n10277), .ZN(n10279) );
  NAND3_X1 U12768 ( .A1(n14752), .A2(n10280), .A3(n10279), .ZN(n10281) );
  OAI211_X1 U12769 ( .C1(n14722), .C2(n10283), .A(n10282), .B(n10281), .ZN(
        P2_U3219) );
  AND2_X1 U12770 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10694) );
  INV_X1 U12771 ( .A(n10284), .ZN(n10289) );
  NOR3_X1 U12772 ( .A1(n10287), .A2(n10286), .A3(n10285), .ZN(n10288) );
  NOR3_X1 U12773 ( .A1(n14745), .A2(n10289), .A3(n10288), .ZN(n10290) );
  AOI211_X1 U12774 ( .C1(n14726), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n10694), .B(
        n10290), .ZN(n10298) );
  MUX2_X1 U12775 ( .A(n10233), .B(P2_REG1_REG_7__SCAN_IN), .S(n10291), .Z(
        n10292) );
  NAND3_X1 U12776 ( .A1(n10294), .A2(n10293), .A3(n10292), .ZN(n10295) );
  NAND3_X1 U12777 ( .A1(n14752), .A2(n10296), .A3(n10295), .ZN(n10297) );
  OAI211_X1 U12778 ( .C1(n14722), .C2(n10299), .A(n10298), .B(n10297), .ZN(
        P2_U3221) );
  OAI222_X1 U12779 ( .A1(P3_U3151), .A2(n11845), .B1(n12944), .B2(n10301), 
        .C1(n11943), .C2(n10300), .ZN(P3_U3282) );
  INV_X1 U12780 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10304) );
  INV_X1 U12781 ( .A(n10309), .ZN(n10302) );
  OAI222_X1 U12782 ( .A1(n13498), .A2(n10304), .B1(n13505), .B2(n10303), .C1(
        n10302), .C2(P2_U3088), .ZN(P2_U3319) );
  AOI21_X1 U12783 ( .B1(n10309), .B2(P2_REG1_REG_8__SCAN_IN), .A(n10305), .ZN(
        n10307) );
  INV_X1 U12784 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n11190) );
  MUX2_X1 U12785 ( .A(n11190), .B(P2_REG1_REG_9__SCAN_IN), .S(n10384), .Z(
        n10306) );
  NAND2_X1 U12786 ( .A1(n10307), .A2(n10306), .ZN(n10389) );
  OAI21_X1 U12787 ( .B1(n10307), .B2(n10306), .A(n10389), .ZN(n10318) );
  AOI21_X1 U12788 ( .B1(n10309), .B2(P2_REG2_REG_8__SCAN_IN), .A(n10308), .ZN(
        n10312) );
  INV_X1 U12789 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10310) );
  MUX2_X1 U12790 ( .A(n10310), .B(P2_REG2_REG_9__SCAN_IN), .S(n10384), .Z(
        n10311) );
  NAND2_X1 U12791 ( .A1(n10312), .A2(n10311), .ZN(n10385) );
  OAI21_X1 U12792 ( .B1(n10312), .B2(n10311), .A(n10385), .ZN(n10313) );
  NAND2_X1 U12793 ( .A1(n10313), .A2(n14729), .ZN(n10316) );
  AND2_X1 U12794 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10314) );
  AOI21_X1 U12795 ( .B1(n14726), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n10314), .ZN(
        n10315) );
  OAI211_X1 U12796 ( .C1(n14722), .C2(n10384), .A(n10316), .B(n10315), .ZN(
        n10317) );
  AOI21_X1 U12797 ( .B1(n14752), .B2(n10318), .A(n10317), .ZN(n10319) );
  INV_X1 U12798 ( .A(n10319), .ZN(P2_U3223) );
  AOI22_X1 U12799 ( .A1(n13754), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n14141), .ZN(n10320) );
  OAI21_X1 U12800 ( .B1(n10337), .B2(n14160), .A(n10320), .ZN(P1_U3346) );
  AOI21_X1 U12801 ( .B1(n13049), .B2(n10321), .A(n13081), .ZN(n10326) );
  OR2_X1 U12802 ( .A1(n10322), .A2(P2_U3088), .ZN(n10377) );
  NAND2_X1 U12803 ( .A1(n13112), .A2(n13076), .ZN(n10503) );
  NAND4_X1 U12804 ( .A1(n13049), .A2(n13336), .A3(n13114), .A4(n10734), .ZN(
        n10323) );
  OAI21_X1 U12805 ( .B1(n13079), .B2(n10503), .A(n10323), .ZN(n10324) );
  AOI21_X1 U12806 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n10377), .A(n10324), .ZN(
        n10325) );
  OAI21_X1 U12807 ( .B1(n10326), .B2(n11968), .A(n10325), .ZN(P2_U3204) );
  INV_X1 U12808 ( .A(n11848), .ZN(n11864) );
  OAI222_X1 U12809 ( .A1(P3_U3151), .A2(n11864), .B1(n12944), .B2(n10328), 
        .C1(n11943), .C2(n10327), .ZN(P3_U3281) );
  INV_X1 U12810 ( .A(n13114), .ZN(n10329) );
  OAI22_X1 U12811 ( .A1(n10329), .A2(n13060), .B1(n10411), .B2(n13042), .ZN(
        n10739) );
  AOI22_X1 U12812 ( .A1(n13065), .A2(n10739), .B1(n10377), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n10335) );
  OAI21_X1 U12813 ( .B1(n10332), .B2(n10331), .A(n10330), .ZN(n10333) );
  NAND2_X1 U12814 ( .A1(n13049), .A2(n10333), .ZN(n10334) );
  OAI211_X1 U12815 ( .C1(n8914), .C2(n10336), .A(n10335), .B(n10334), .ZN(
        P2_U3194) );
  OAI222_X1 U12816 ( .A1(n13498), .A2(n10338), .B1(n13505), .B2(n10337), .C1(
        n10384), .C2(P2_U3088), .ZN(P2_U3318) );
  NAND2_X1 U12817 ( .A1(n11938), .A2(P3_D_REG_1__SCAN_IN), .ZN(n10339) );
  OAI21_X1 U12818 ( .B1(n11063), .B2(n11938), .A(n10339), .ZN(P3_U3377) );
  AOI22_X1 U12819 ( .A1(n13768), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n14141), .ZN(n10340) );
  OAI21_X1 U12820 ( .B1(n10372), .B2(n14160), .A(n10340), .ZN(P1_U3345) );
  INV_X1 U12821 ( .A(n10344), .ZN(n10365) );
  AND2_X1 U12822 ( .A1(n10347), .A2(n10346), .ZN(n10599) );
  AND2_X1 U12823 ( .A1(n10351), .A2(n10350), .ZN(n10598) );
  XNOR2_X1 U12824 ( .A(n10598), .B(n10599), .ZN(n10522) );
  NOR2_X1 U12825 ( .A1(n10513), .A2(n10518), .ZN(n10363) );
  AND2_X1 U12826 ( .A1(n10363), .A2(n10515), .ZN(n10361) );
  NAND2_X1 U12827 ( .A1(n10354), .A2(n13944), .ZN(n10356) );
  NOR2_X1 U12828 ( .A1(n14635), .A2(n10357), .ZN(n10358) );
  NAND2_X1 U12829 ( .A1(n10361), .A2(n10514), .ZN(n13656) );
  INV_X1 U12830 ( .A(n13647), .ZN(n13595) );
  NAND2_X1 U12831 ( .A1(n10361), .A2(n10360), .ZN(n10362) );
  AOI22_X1 U12832 ( .A1(n13595), .A2(n10359), .B1(n14013), .B2(n13658), .ZN(
        n10371) );
  INV_X1 U12833 ( .A(n10363), .ZN(n10364) );
  NAND2_X1 U12834 ( .A1(n10364), .A2(n10516), .ZN(n10369) );
  NOR2_X1 U12835 ( .A1(n10366), .A2(n10365), .ZN(n10367) );
  AND2_X1 U12836 ( .A1(n10514), .A2(n10367), .ZN(n10368) );
  NAND2_X1 U12837 ( .A1(n10369), .A2(n10368), .ZN(n10960) );
  OR2_X1 U12838 ( .A1(n10960), .A2(P1_U3086), .ZN(n13557) );
  NAND2_X1 U12839 ( .A1(n13557), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n10370) );
  OAI211_X1 U12840 ( .C1(n10522), .C2(n13660), .A(n10371), .B(n10370), .ZN(
        P1_U3232) );
  INV_X1 U12841 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10373) );
  INV_X1 U12842 ( .A(n10459), .ZN(n10467) );
  OAI222_X1 U12843 ( .A1(n13498), .A2(n10373), .B1(n13505), .B2(n10372), .C1(
        n10467), .C2(P2_U3088), .ZN(P2_U3317) );
  INV_X1 U12844 ( .A(n10374), .ZN(n10375) );
  OAI222_X1 U12845 ( .A1(n12944), .A2(n15227), .B1(n11943), .B2(n10375), .C1(
        n12533), .C2(P3_U3151), .ZN(P3_U3280) );
  INV_X1 U12846 ( .A(n13112), .ZN(n10376) );
  OAI22_X1 U12847 ( .A1(n10376), .A2(n13060), .B1(n10586), .B2(n13042), .ZN(
        n10842) );
  AOI22_X1 U12848 ( .A1(n13065), .A2(n10842), .B1(n10377), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n10383) );
  OAI21_X1 U12849 ( .B1(n10380), .B2(n10379), .A(n10378), .ZN(n10381) );
  NAND2_X1 U12850 ( .A1(n13049), .A2(n10381), .ZN(n10382) );
  OAI211_X1 U12851 ( .C1(n8914), .C2(n6770), .A(n10383), .B(n10382), .ZN(
        P2_U3209) );
  INV_X1 U12852 ( .A(n10384), .ZN(n10390) );
  OAI21_X1 U12853 ( .B1(n10390), .B2(P2_REG2_REG_9__SCAN_IN), .A(n10385), .ZN(
        n10388) );
  INV_X1 U12854 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10386) );
  MUX2_X1 U12855 ( .A(n10386), .B(P2_REG2_REG_10__SCAN_IN), .S(n10459), .Z(
        n10387) );
  NOR2_X1 U12856 ( .A1(n10388), .A2(n10387), .ZN(n10458) );
  AOI211_X1 U12857 ( .C1(n10388), .C2(n10387), .A(n14745), .B(n10458), .ZN(
        n10396) );
  OAI21_X1 U12858 ( .B1(n10390), .B2(P2_REG1_REG_9__SCAN_IN), .A(n10389), .ZN(
        n10392) );
  INV_X1 U12859 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n11234) );
  MUX2_X1 U12860 ( .A(n11234), .B(P2_REG1_REG_10__SCAN_IN), .S(n10459), .Z(
        n10391) );
  NOR2_X1 U12861 ( .A1(n10392), .A2(n10391), .ZN(n10473) );
  AOI211_X1 U12862 ( .C1(n10392), .C2(n10391), .A(n14718), .B(n10473), .ZN(
        n10395) );
  NAND2_X1 U12863 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n11122)
         );
  NAND2_X1 U12864 ( .A1(n14726), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n10393) );
  OAI211_X1 U12865 ( .C1(n14722), .C2(n10467), .A(n11122), .B(n10393), .ZN(
        n10394) );
  OR3_X1 U12866 ( .A1(n10396), .A2(n10395), .A3(n10394), .ZN(P2_U3224) );
  NAND2_X1 U12867 ( .A1(n12977), .A2(P2_U3947), .ZN(n10397) );
  OAI21_X1 U12868 ( .B1(P2_U3947), .B2(n10398), .A(n10397), .ZN(P2_U3553) );
  INV_X1 U12869 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10400) );
  NOR2_X1 U12870 ( .A1(n10637), .A2(n10400), .ZN(P3_U3250) );
  INV_X1 U12871 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n15334) );
  NOR2_X1 U12872 ( .A1(n10637), .A2(n15334), .ZN(P3_U3254) );
  INV_X1 U12873 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10401) );
  NOR2_X1 U12874 ( .A1(n10637), .A2(n10401), .ZN(P3_U3246) );
  INV_X1 U12875 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n15417) );
  NOR2_X1 U12876 ( .A1(n10637), .A2(n15417), .ZN(P3_U3252) );
  INV_X1 U12877 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10402) );
  NOR2_X1 U12878 ( .A1(n10637), .A2(n10402), .ZN(P3_U3248) );
  INV_X1 U12879 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10403) );
  NOR2_X1 U12880 ( .A1(n10637), .A2(n10403), .ZN(P3_U3247) );
  INV_X1 U12881 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n15377) );
  NOR2_X1 U12882 ( .A1(n10637), .A2(n15377), .ZN(P3_U3253) );
  INV_X1 U12883 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10404) );
  NOR2_X1 U12884 ( .A1(n10637), .A2(n10404), .ZN(P3_U3251) );
  INV_X1 U12885 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10405) );
  NOR2_X1 U12886 ( .A1(n10637), .A2(n10405), .ZN(P3_U3243) );
  INV_X1 U12887 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10406) );
  NOR2_X1 U12888 ( .A1(n10637), .A2(n10406), .ZN(P3_U3249) );
  INV_X1 U12889 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10407) );
  NOR2_X1 U12890 ( .A1(n10637), .A2(n10407), .ZN(P3_U3242) );
  INV_X1 U12891 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n15340) );
  NOR2_X1 U12892 ( .A1(n10637), .A2(n15340), .ZN(P3_U3241) );
  XNOR2_X1 U12893 ( .A(n10409), .B(n10408), .ZN(n10414) );
  OAI22_X1 U12894 ( .A1(n10411), .A2(n13060), .B1(n10410), .B2(n13042), .ZN(
        n10984) );
  AOI22_X1 U12895 ( .A1(n13065), .A2(n10984), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10413) );
  AOI22_X1 U12896 ( .A1(n13081), .A2(n11987), .B1(n13077), .B2(n8290), .ZN(
        n10412) );
  OAI211_X1 U12897 ( .C1(n10414), .C2(n13083), .A(n10413), .B(n10412), .ZN(
        P2_U3190) );
  MUX2_X1 U12898 ( .A(n14658), .B(P1_REG1_REG_8__SCAN_IN), .S(n10544), .Z(
        n10422) );
  INV_X1 U12899 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n14656) );
  INV_X1 U12900 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10415) );
  MUX2_X1 U12901 ( .A(n10415), .B(P1_REG1_REG_2__SCAN_IN), .S(n13690), .Z(
        n10418) );
  INV_X1 U12902 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10416) );
  MUX2_X1 U12903 ( .A(n10416), .B(P1_REG1_REG_1__SCAN_IN), .S(n10431), .Z(
        n13678) );
  AND2_X1 U12904 ( .A1(n6762), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n13679) );
  NAND2_X1 U12905 ( .A1(n13678), .A2(n13679), .ZN(n13677) );
  INV_X1 U12906 ( .A(n10431), .ZN(n13676) );
  NAND2_X1 U12907 ( .A1(n13676), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10417) );
  NAND2_X1 U12908 ( .A1(n13677), .A2(n10417), .ZN(n13686) );
  NAND2_X1 U12909 ( .A1(n10418), .A2(n13686), .ZN(n13707) );
  OR2_X1 U12910 ( .A1(n13690), .A2(n10415), .ZN(n13706) );
  NAND2_X1 U12911 ( .A1(n13707), .A2(n13706), .ZN(n10420) );
  MUX2_X1 U12912 ( .A(n14648), .B(P1_REG1_REG_3__SCAN_IN), .S(n13705), .Z(
        n10419) );
  NAND2_X1 U12913 ( .A1(n10420), .A2(n10419), .ZN(n13710) );
  INV_X1 U12914 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n14648) );
  OR2_X1 U12915 ( .A1(n13705), .A2(n14648), .ZN(n10528) );
  INV_X1 U12916 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n14650) );
  MUX2_X1 U12917 ( .A(n14650), .B(P1_REG1_REG_4__SCAN_IN), .S(n10539), .Z(
        n10527) );
  AOI21_X1 U12918 ( .B1(n13710), .B2(n10528), .A(n10527), .ZN(n10526) );
  AOI21_X1 U12919 ( .B1(n10539), .B2(P1_REG1_REG_4__SCAN_IN), .A(n10526), .ZN(
        n13719) );
  INV_X1 U12920 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n14652) );
  MUX2_X1 U12921 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n14652), .S(n13722), .Z(
        n13720) );
  NAND2_X1 U12922 ( .A1(n13719), .A2(n13720), .ZN(n13718) );
  OAI21_X1 U12923 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n13722), .A(n13718), .ZN(
        n13733) );
  INV_X1 U12924 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14654) );
  MUX2_X1 U12925 ( .A(n14654), .B(P1_REG1_REG_6__SCAN_IN), .S(n13737), .Z(
        n13732) );
  NOR2_X1 U12926 ( .A1(n13733), .A2(n13732), .ZN(n13731) );
  AOI21_X1 U12927 ( .B1(n13737), .B2(P1_REG1_REG_6__SCAN_IN), .A(n13731), .ZN(
        n10482) );
  MUX2_X1 U12928 ( .A(n14656), .B(P1_REG1_REG_7__SCAN_IN), .S(n10476), .Z(
        n10481) );
  OR2_X1 U12929 ( .A1(n10482), .A2(n10481), .ZN(n10483) );
  OAI21_X1 U12930 ( .B1(n14656), .B2(n10489), .A(n10483), .ZN(n10421) );
  NOR2_X1 U12931 ( .A1(n10421), .A2(n10422), .ZN(n13749) );
  AOI21_X1 U12932 ( .B1(n10422), .B2(n10421), .A(n13749), .ZN(n10454) );
  INV_X1 U12933 ( .A(n10423), .ZN(n10425) );
  NAND2_X1 U12934 ( .A1(n10425), .A2(n10424), .ZN(n14470) );
  NOR2_X2 U12935 ( .A1(n14470), .A2(n14466), .ZN(n14486) );
  INV_X1 U12936 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10426) );
  NOR2_X1 U12937 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10426), .ZN(n11336) );
  NOR2_X1 U12938 ( .A1(n14470), .A2(n10523), .ZN(n13792) );
  INV_X1 U12939 ( .A(n10544), .ZN(n10427) );
  NOR2_X1 U12940 ( .A1(n14494), .A2(n10427), .ZN(n10428) );
  AOI211_X1 U12941 ( .C1(n14468), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n11336), .B(
        n10428), .ZN(n10453) );
  INV_X1 U12942 ( .A(n14470), .ZN(n10430) );
  NOR2_X1 U12943 ( .A1(n9721), .A2(n14150), .ZN(n10429) );
  NAND2_X1 U12944 ( .A1(n10430), .A2(n10429), .ZN(n14477) );
  INV_X1 U12945 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10722) );
  MUX2_X1 U12946 ( .A(n10722), .B(P1_REG2_REG_2__SCAN_IN), .S(n13690), .Z(
        n13685) );
  INV_X1 U12947 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10432) );
  MUX2_X1 U12948 ( .A(n10432), .B(P1_REG2_REG_1__SCAN_IN), .S(n10431), .Z(
        n13674) );
  AND2_X1 U12949 ( .A1(n6762), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n13675) );
  NAND2_X1 U12950 ( .A1(n13674), .A2(n13675), .ZN(n13673) );
  NAND2_X1 U12951 ( .A1(n13676), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10433) );
  NAND2_X1 U12952 ( .A1(n13673), .A2(n10433), .ZN(n13684) );
  NAND2_X1 U12953 ( .A1(n13685), .A2(n13684), .ZN(n13700) );
  OR2_X1 U12954 ( .A1(n13690), .A2(n10722), .ZN(n13699) );
  NAND2_X1 U12955 ( .A1(n13700), .A2(n13699), .ZN(n10436) );
  INV_X1 U12956 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10434) );
  MUX2_X1 U12957 ( .A(n10434), .B(P1_REG2_REG_3__SCAN_IN), .S(n13705), .Z(
        n10435) );
  NAND2_X1 U12958 ( .A1(n10436), .A2(n10435), .ZN(n13703) );
  OR2_X1 U12959 ( .A1(n13705), .A2(n10434), .ZN(n10533) );
  NAND2_X1 U12960 ( .A1(n13703), .A2(n10533), .ZN(n10438) );
  INV_X1 U12961 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10531) );
  MUX2_X1 U12962 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10531), .S(n10539), .Z(
        n10437) );
  NAND2_X1 U12963 ( .A1(n10438), .A2(n10437), .ZN(n13726) );
  NAND2_X1 U12964 ( .A1(n10539), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n13725) );
  NAND2_X1 U12965 ( .A1(n13726), .A2(n13725), .ZN(n10440) );
  INV_X1 U12966 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n13723) );
  MUX2_X1 U12967 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n13723), .S(n13722), .Z(
        n10439) );
  NAND2_X1 U12968 ( .A1(n10440), .A2(n10439), .ZN(n13740) );
  NAND2_X1 U12969 ( .A1(n13722), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n13739) );
  NAND2_X1 U12970 ( .A1(n13740), .A2(n13739), .ZN(n10442) );
  INV_X1 U12971 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10904) );
  MUX2_X1 U12972 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10904), .S(n13737), .Z(
        n10441) );
  NAND2_X1 U12973 ( .A1(n10442), .A2(n10441), .ZN(n13742) );
  NAND2_X1 U12974 ( .A1(n13737), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10478) );
  NAND2_X1 U12975 ( .A1(n13742), .A2(n10478), .ZN(n10445) );
  INV_X1 U12976 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10443) );
  MUX2_X1 U12977 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10443), .S(n10476), .Z(
        n10444) );
  NAND2_X1 U12978 ( .A1(n10445), .A2(n10444), .ZN(n10480) );
  NAND2_X1 U12979 ( .A1(n10476), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10450) );
  NAND2_X1 U12980 ( .A1(n10480), .A2(n10450), .ZN(n10448) );
  INV_X1 U12981 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10446) );
  MUX2_X1 U12982 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10446), .S(n10544), .Z(
        n10447) );
  NAND2_X1 U12983 ( .A1(n10448), .A2(n10447), .ZN(n13757) );
  MUX2_X1 U12984 ( .A(n10446), .B(P1_REG2_REG_8__SCAN_IN), .S(n10544), .Z(
        n10449) );
  NAND3_X1 U12985 ( .A1(n10480), .A2(n10450), .A3(n10449), .ZN(n10451) );
  NAND3_X1 U12986 ( .A1(n14489), .A2(n13757), .A3(n10451), .ZN(n10452) );
  OAI211_X1 U12987 ( .C1(n10454), .C2(n14479), .A(n10453), .B(n10452), .ZN(
        P1_U3251) );
  INV_X1 U12988 ( .A(n10455), .ZN(n10457) );
  OAI222_X1 U12989 ( .A1(P3_U3151), .A2(n12556), .B1(n11943), .B2(n10457), 
        .C1(n10456), .C2(n12944), .ZN(P3_U3279) );
  AOI21_X1 U12990 ( .B1(n10459), .B2(P2_REG2_REG_10__SCAN_IN), .A(n10458), 
        .ZN(n10463) );
  INV_X1 U12991 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10460) );
  MUX2_X1 U12992 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10460), .S(n10575), .Z(
        n10462) );
  INV_X1 U12993 ( .A(n10570), .ZN(n10461) );
  OAI21_X1 U12994 ( .B1(n10463), .B2(n10462), .A(n10461), .ZN(n10466) );
  INV_X1 U12995 ( .A(n10575), .ZN(n10491) );
  NAND2_X1 U12996 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11197)
         );
  NAND2_X1 U12997 ( .A1(n14726), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n10464) );
  OAI211_X1 U12998 ( .C1(n14722), .C2(n10491), .A(n11197), .B(n10464), .ZN(
        n10465) );
  AOI21_X1 U12999 ( .B1(n10466), .B2(n14729), .A(n10465), .ZN(n10475) );
  NOR2_X1 U13000 ( .A1(n10467), .A2(n11234), .ZN(n10471) );
  INV_X1 U13001 ( .A(n10471), .ZN(n10469) );
  INV_X1 U13002 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11480) );
  MUX2_X1 U13003 ( .A(n11480), .B(P2_REG1_REG_11__SCAN_IN), .S(n10575), .Z(
        n10468) );
  NAND2_X1 U13004 ( .A1(n10469), .A2(n10468), .ZN(n10472) );
  MUX2_X1 U13005 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n11480), .S(n10575), .Z(
        n10470) );
  OAI21_X1 U13006 ( .B1(n10473), .B2(n10471), .A(n10470), .ZN(n10578) );
  OAI211_X1 U13007 ( .C1(n10473), .C2(n10472), .A(n10578), .B(n14752), .ZN(
        n10474) );
  NAND2_X1 U13008 ( .A1(n10475), .A2(n10474), .ZN(P2_U3225) );
  MUX2_X1 U13009 ( .A(n10443), .B(P1_REG2_REG_7__SCAN_IN), .S(n10476), .Z(
        n10477) );
  NAND3_X1 U13010 ( .A1(n13742), .A2(n10478), .A3(n10477), .ZN(n10479) );
  NAND3_X1 U13011 ( .A1(n14489), .A2(n10480), .A3(n10479), .ZN(n10488) );
  NAND2_X1 U13012 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11220) );
  AOI21_X1 U13013 ( .B1(n10482), .B2(n10481), .A(n14479), .ZN(n10484) );
  NAND2_X1 U13014 ( .A1(n10484), .A2(n10483), .ZN(n10485) );
  NAND2_X1 U13015 ( .A1(n11220), .A2(n10485), .ZN(n10486) );
  AOI21_X1 U13016 ( .B1(n14468), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n10486), .ZN(
        n10487) );
  OAI211_X1 U13017 ( .C1(n14494), .C2(n10489), .A(n10488), .B(n10487), .ZN(
        P1_U3250) );
  INV_X1 U13018 ( .A(n10490), .ZN(n10493) );
  OAI222_X1 U13019 ( .A1(n13498), .A2(n10492), .B1(n13505), .B2(n10493), .C1(
        P2_U3088), .C2(n10491), .ZN(P2_U3316) );
  OAI222_X1 U13020 ( .A1(n7001), .A2(n10494), .B1(n14160), .B2(n10493), .C1(
        P1_U3086), .C2(n10660), .ZN(P1_U3344) );
  INV_X1 U13021 ( .A(n10495), .ZN(n10496) );
  NAND3_X1 U13022 ( .A1(n10498), .A2(n10497), .A3(n10496), .ZN(n10499) );
  NAND2_X1 U13023 ( .A1(n12161), .A2(n12201), .ZN(n10732) );
  INV_X1 U13024 ( .A(n10732), .ZN(n10500) );
  NAND2_X1 U13025 ( .A1(n13357), .A2(n10500), .ZN(n10993) );
  OR2_X1 U13026 ( .A1(n13114), .A2(n11972), .ZN(n10501) );
  NAND2_X1 U13027 ( .A1(n10734), .A2(n10501), .ZN(n14785) );
  NAND2_X1 U13028 ( .A1(n11972), .A2(n10502), .ZN(n14782) );
  AOI21_X1 U13029 ( .B1(n13332), .B2(n14815), .A(n14785), .ZN(n10505) );
  INV_X1 U13030 ( .A(n10503), .ZN(n10504) );
  NOR2_X1 U13031 ( .A1(n10505), .A2(n10504), .ZN(n14783) );
  OAI21_X1 U13032 ( .B1(n12161), .B2(n14782), .A(n14783), .ZN(n10506) );
  INV_X1 U13033 ( .A(n13354), .ZN(n14759) );
  AOI22_X1 U13034 ( .A1(n13357), .A2(n10506), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n14759), .ZN(n10508) );
  NAND2_X1 U13035 ( .A1(n14761), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10507) );
  OAI211_X1 U13036 ( .C1(n10993), .C2(n14785), .A(n10508), .B(n10507), .ZN(
        P2_U3265) );
  OR2_X1 U13037 ( .A1(n10509), .A2(n13944), .ZN(n14602) );
  AND2_X1 U13038 ( .A1(n11201), .A2(n13944), .ZN(n10510) );
  NAND2_X1 U13039 ( .A1(n10511), .A2(n10510), .ZN(n14601) );
  NAND2_X1 U13040 ( .A1(n14563), .A2(n14533), .ZN(n10512) );
  AOI222_X1 U13041 ( .A1(n14010), .A2(n10512), .B1(n10354), .B2(n14013), .C1(
        n10359), .C2(n14617), .ZN(n14557) );
  AND2_X1 U13042 ( .A1(n10515), .A2(n10514), .ZN(n10517) );
  NAND2_X1 U13043 ( .A1(n14662), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10520) );
  OAI21_X1 U13044 ( .B1(n14557), .B2(n14662), .A(n10520), .ZN(P1_U3528) );
  INV_X1 U13045 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10521) );
  AOI21_X1 U13046 ( .B1(n14466), .B2(n10521), .A(n9721), .ZN(n14465) );
  MUX2_X1 U13047 ( .A(n13675), .B(n10522), .S(n14150), .Z(n10524) );
  NAND2_X1 U13048 ( .A1(n10524), .A2(n10523), .ZN(n10525) );
  OAI211_X1 U13049 ( .C1(n6762), .C2(n14465), .A(n10525), .B(P1_U4016), .ZN(
        n13698) );
  INV_X1 U13050 ( .A(n10526), .ZN(n10530) );
  NAND3_X1 U13051 ( .A1(n13710), .A2(n10528), .A3(n10527), .ZN(n10529) );
  AND3_X1 U13052 ( .A1(n14486), .A2(n10530), .A3(n10529), .ZN(n10538) );
  INV_X1 U13053 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10536) );
  INV_X1 U13054 ( .A(n14468), .ZN(n14498) );
  MUX2_X1 U13055 ( .A(n10531), .B(P1_REG2_REG_4__SCAN_IN), .S(n10539), .Z(
        n10532) );
  NAND3_X1 U13056 ( .A1(n13703), .A2(n10533), .A3(n10532), .ZN(n10534) );
  NAND3_X1 U13057 ( .A1(n14489), .A2(n13726), .A3(n10534), .ZN(n10535) );
  NAND2_X1 U13058 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n10963) );
  OAI211_X1 U13059 ( .C1(n10536), .C2(n14498), .A(n10535), .B(n10963), .ZN(
        n10537) );
  AOI211_X1 U13060 ( .C1(n13792), .C2(n10539), .A(n10538), .B(n10537), .ZN(
        n10540) );
  NAND2_X1 U13061 ( .A1(n13698), .A2(n10540), .ZN(P1_U3247) );
  INV_X1 U13062 ( .A(n10541), .ZN(n10542) );
  OAI222_X1 U13063 ( .A1(P3_U3151), .A2(n12575), .B1(n12944), .B2(n10543), 
        .C1(n11943), .C2(n10542), .ZN(P3_U3278) );
  NOR2_X1 U13064 ( .A1(n10544), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n13747) );
  INV_X1 U13065 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n14660) );
  MUX2_X1 U13066 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n14660), .S(n13754), .Z(
        n13748) );
  OAI21_X1 U13067 ( .B1(n13749), .B2(n13747), .A(n13748), .ZN(n13746) );
  OAI21_X1 U13068 ( .B1(n13754), .B2(P1_REG1_REG_9__SCAN_IN), .A(n13746), .ZN(
        n13764) );
  INV_X1 U13069 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14663) );
  MUX2_X1 U13070 ( .A(n14663), .B(P1_REG1_REG_10__SCAN_IN), .S(n13768), .Z(
        n13763) );
  NOR2_X1 U13071 ( .A1(n13764), .A2(n13763), .ZN(n13762) );
  AOI21_X1 U13072 ( .B1(n13768), .B2(P1_REG1_REG_10__SCAN_IN), .A(n13762), 
        .ZN(n10561) );
  INV_X1 U13073 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n14431) );
  NOR3_X1 U13074 ( .A1(n10561), .A2(n14431), .A3(n14479), .ZN(n10552) );
  NAND2_X1 U13075 ( .A1(n10544), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n13756) );
  NAND2_X1 U13076 ( .A1(n13757), .A2(n13756), .ZN(n10547) );
  INV_X1 U13077 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10545) );
  MUX2_X1 U13078 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10545), .S(n13754), .Z(
        n10546) );
  NAND2_X1 U13079 ( .A1(n10547), .A2(n10546), .ZN(n13772) );
  NAND2_X1 U13080 ( .A1(n13754), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n13771) );
  NAND2_X1 U13081 ( .A1(n13772), .A2(n13771), .ZN(n10549) );
  MUX2_X1 U13082 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n13769), .S(n13768), .Z(
        n10548) );
  NAND2_X1 U13083 ( .A1(n10549), .A2(n10548), .ZN(n13774) );
  NAND2_X1 U13084 ( .A1(n13768), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10550) );
  NAND2_X1 U13085 ( .A1(n13774), .A2(n10550), .ZN(n10556) );
  NOR3_X1 U13086 ( .A1(n10556), .A2(n14477), .A3(P1_REG2_REG_11__SCAN_IN), 
        .ZN(n10551) );
  NOR3_X1 U13087 ( .A1(n10552), .A2(n13792), .A3(n10551), .ZN(n10565) );
  AOI21_X1 U13088 ( .B1(n10660), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10556), 
        .ZN(n10553) );
  NOR2_X1 U13089 ( .A1(n10553), .A2(n14477), .ZN(n10558) );
  INV_X1 U13090 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10554) );
  MUX2_X1 U13091 ( .A(n10554), .B(P1_REG2_REG_11__SCAN_IN), .S(n10660), .Z(
        n10555) );
  NAND2_X1 U13092 ( .A1(n10556), .A2(n10555), .ZN(n10659) );
  NAND2_X1 U13093 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n11756)
         );
  OAI21_X1 U13094 ( .B1(n14498), .B2(n14188), .A(n11756), .ZN(n10557) );
  AOI21_X1 U13095 ( .B1(n10558), .B2(n10659), .A(n10557), .ZN(n10564) );
  INV_X1 U13096 ( .A(n10660), .ZN(n10559) );
  NOR3_X1 U13097 ( .A1(n10561), .A2(P1_REG1_REG_11__SCAN_IN), .A3(n10559), 
        .ZN(n10562) );
  MUX2_X1 U13098 ( .A(n14431), .B(P1_REG1_REG_11__SCAN_IN), .S(n10660), .Z(
        n10560) );
  AND2_X1 U13099 ( .A1(n10561), .A2(n10560), .ZN(n10654) );
  OAI21_X1 U13100 ( .B1(n10562), .B2(n10654), .A(n14486), .ZN(n10563) );
  OAI211_X1 U13101 ( .C1(n10565), .C2(n10660), .A(n10564), .B(n10563), .ZN(
        P1_U3254) );
  INV_X1 U13102 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14448) );
  NAND2_X1 U13103 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n10566)
         );
  OAI21_X1 U13104 ( .B1(n14741), .B2(n14448), .A(n10566), .ZN(n10573) );
  NOR2_X1 U13105 ( .A1(n10575), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10568) );
  INV_X1 U13106 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10567) );
  MUX2_X1 U13107 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n10567), .S(n11552), .Z(
        n10569) );
  OAI21_X1 U13108 ( .B1(n10570), .B2(n10568), .A(n10569), .ZN(n11542) );
  OR3_X1 U13109 ( .A1(n10570), .A2(n10569), .A3(n10568), .ZN(n10571) );
  AOI21_X1 U13110 ( .B1(n11542), .B2(n10571), .A(n14745), .ZN(n10572) );
  AOI211_X1 U13111 ( .C1(n14750), .C2(n11552), .A(n10573), .B(n10572), .ZN(
        n10582) );
  INV_X1 U13112 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10574) );
  XNOR2_X1 U13113 ( .A(n11552), .B(n10574), .ZN(n10576) );
  NAND2_X1 U13114 ( .A1(n10575), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10577) );
  NAND3_X1 U13115 ( .A1(n10578), .A2(n10576), .A3(n10577), .ZN(n11551) );
  INV_X1 U13116 ( .A(n11551), .ZN(n10580) );
  AOI21_X1 U13117 ( .B1(n10578), .B2(n10577), .A(n10576), .ZN(n10579) );
  OAI21_X1 U13118 ( .B1(n10580), .B2(n10579), .A(n14752), .ZN(n10581) );
  NAND2_X1 U13119 ( .A1(n10582), .A2(n10581), .ZN(P2_U3226) );
  INV_X1 U13120 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10592) );
  CLKBUF_X1 U13121 ( .A(n10583), .Z(n10584) );
  XNOR2_X1 U13122 ( .A(n10584), .B(n12168), .ZN(n11088) );
  AOI211_X1 U13123 ( .C1(n13031), .C2(n10988), .A(n13336), .B(n10973), .ZN(
        n11084) );
  AOI21_X1 U13124 ( .B1(n14792), .B2(n13031), .A(n11084), .ZN(n10590) );
  XNOR2_X1 U13125 ( .A(n10585), .B(n12168), .ZN(n10589) );
  OR2_X1 U13126 ( .A1(n10586), .A2(n13060), .ZN(n10588) );
  NAND2_X1 U13127 ( .A1(n13109), .A2(n13076), .ZN(n10587) );
  NAND2_X1 U13128 ( .A1(n10588), .A2(n10587), .ZN(n13032) );
  AOI21_X1 U13129 ( .B1(n10589), .B2(n13350), .A(n13032), .ZN(n11085) );
  OAI211_X1 U13130 ( .C1(n13456), .C2(n11088), .A(n10590), .B(n11085), .ZN(
        n10689) );
  NAND2_X1 U13131 ( .A1(n10689), .A2(n6621), .ZN(n10591) );
  OAI21_X1 U13132 ( .B1(n6621), .B2(n10592), .A(n10591), .ZN(P2_U3442) );
  INV_X1 U13133 ( .A(n10593), .ZN(n10594) );
  OAI222_X1 U13134 ( .A1(P3_U3151), .A2(n12600), .B1(n12944), .B2(n10595), 
        .C1(n11943), .C2(n10594), .ZN(P3_U3277) );
  OAI222_X1 U13135 ( .A1(n11943), .A2(n10597), .B1(n12944), .B2(n10596), .C1(
        P3_U3151), .C2(n12607), .ZN(P3_U3276) );
  INV_X1 U13136 ( .A(n13658), .ZN(n13640) );
  NAND2_X1 U13137 ( .A1(n10598), .A2(n11327), .ZN(n10602) );
  INV_X1 U13138 ( .A(n10598), .ZN(n10600) );
  NAND2_X1 U13139 ( .A1(n10602), .A2(n10601), .ZN(n13554) );
  XNOR2_X1 U13140 ( .A(n10604), .B(n11327), .ZN(n10609) );
  NAND2_X1 U13141 ( .A1(n10603), .A2(n14558), .ZN(n10607) );
  NAND2_X1 U13142 ( .A1(n10605), .A2(n12321), .ZN(n10606) );
  OR2_X1 U13143 ( .A1(n10610), .A2(n10609), .ZN(n10611) );
  NAND2_X1 U13144 ( .A1(n9894), .A2(n10603), .ZN(n10614) );
  NAND2_X1 U13145 ( .A1(n10727), .A2(n12313), .ZN(n10613) );
  NAND2_X1 U13146 ( .A1(n10614), .A2(n10613), .ZN(n10615) );
  XNOR2_X1 U13147 ( .A(n10615), .B(n11327), .ZN(n10943) );
  AOI22_X1 U13148 ( .A1(n12321), .A2(n9894), .B1(n10603), .B2(n10727), .ZN(
        n10944) );
  XNOR2_X1 U13149 ( .A(n10943), .B(n10944), .ZN(n10946) );
  XNOR2_X1 U13150 ( .A(n10947), .B(n10946), .ZN(n10616) );
  NAND2_X1 U13151 ( .A1(n10616), .A2(n13634), .ZN(n10620) );
  INV_X1 U13152 ( .A(n13656), .ZN(n13540) );
  OR2_X1 U13153 ( .A1(n9363), .A2(n14410), .ZN(n10618) );
  NAND2_X1 U13154 ( .A1(n14583), .A2(n14617), .ZN(n10617) );
  NAND2_X1 U13155 ( .A1(n10618), .A2(n10617), .ZN(n10721) );
  AOI22_X1 U13156 ( .A1(n13540), .A2(n10721), .B1(n13557), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n10619) );
  OAI211_X1 U13157 ( .C1(n14569), .C2(n13640), .A(n10620), .B(n10619), .ZN(
        P1_U3237) );
  INV_X1 U13158 ( .A(n10621), .ZN(n10624) );
  INV_X1 U13159 ( .A(n10815), .ZN(n10657) );
  OAI222_X1 U13160 ( .A1(n7001), .A2(n10622), .B1(n14160), .B2(n10624), .C1(
        n10657), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U13161 ( .A(n11552), .ZN(n10623) );
  OAI222_X1 U13162 ( .A1(n13498), .A2(n10625), .B1(n13505), .B2(n10624), .C1(
        n10623), .C2(P2_U3088), .ZN(P2_U3315) );
  OAI21_X1 U13163 ( .B1(n10628), .B2(n10627), .A(n10626), .ZN(n10629) );
  NAND2_X1 U13164 ( .A1(n10629), .A2(n13049), .ZN(n10636) );
  NAND2_X1 U13165 ( .A1(n13108), .A2(n13076), .ZN(n10631) );
  NAND2_X1 U13166 ( .A1(n13110), .A2(n13075), .ZN(n10630) );
  NAND2_X1 U13167 ( .A1(n10631), .A2(n10630), .ZN(n10970) );
  INV_X1 U13168 ( .A(n13077), .ZN(n13067) );
  INV_X1 U13169 ( .A(n10974), .ZN(n10632) );
  NOR2_X1 U13170 ( .A1(n13067), .A2(n10632), .ZN(n10633) );
  AOI211_X1 U13171 ( .C1(n13065), .C2(n10970), .A(n10634), .B(n10633), .ZN(
        n10635) );
  OAI211_X1 U13172 ( .C1(n14812), .C2(n8914), .A(n10636), .B(n10635), .ZN(
        P2_U3199) );
  NOR2_X1 U13173 ( .A1(n10653), .A2(n15265), .ZN(P3_U3255) );
  INV_X1 U13174 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10638) );
  NOR2_X1 U13175 ( .A1(n10653), .A2(n10638), .ZN(P3_U3256) );
  INV_X1 U13176 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10639) );
  NOR2_X1 U13177 ( .A1(n10653), .A2(n10639), .ZN(P3_U3236) );
  INV_X1 U13178 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10640) );
  NOR2_X1 U13179 ( .A1(n10653), .A2(n10640), .ZN(P3_U3235) );
  NOR2_X1 U13180 ( .A1(n10653), .A2(n10641), .ZN(P3_U3263) );
  NOR2_X1 U13181 ( .A1(n10653), .A2(n15268), .ZN(P3_U3234) );
  INV_X1 U13182 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10642) );
  NOR2_X1 U13183 ( .A1(n10653), .A2(n10642), .ZN(P3_U3238) );
  INV_X1 U13184 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10643) );
  NOR2_X1 U13185 ( .A1(n10653), .A2(n10643), .ZN(P3_U3245) );
  INV_X1 U13186 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10644) );
  NOR2_X1 U13187 ( .A1(n10653), .A2(n10644), .ZN(P3_U3244) );
  NOR2_X1 U13188 ( .A1(n10653), .A2(n10645), .ZN(P3_U3258) );
  INV_X1 U13189 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10646) );
  NOR2_X1 U13190 ( .A1(n10653), .A2(n10646), .ZN(P3_U3237) );
  INV_X1 U13191 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10647) );
  NOR2_X1 U13192 ( .A1(n10653), .A2(n10647), .ZN(P3_U3261) );
  INV_X1 U13193 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10648) );
  NOR2_X1 U13194 ( .A1(n10653), .A2(n10648), .ZN(P3_U3260) );
  INV_X1 U13195 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10649) );
  NOR2_X1 U13196 ( .A1(n10653), .A2(n10649), .ZN(P3_U3240) );
  INV_X1 U13197 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n15341) );
  NOR2_X1 U13198 ( .A1(n10653), .A2(n15341), .ZN(P3_U3239) );
  INV_X1 U13199 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10650) );
  NOR2_X1 U13200 ( .A1(n10653), .A2(n10650), .ZN(P3_U3262) );
  INV_X1 U13201 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10651) );
  NOR2_X1 U13202 ( .A1(n10653), .A2(n10651), .ZN(P3_U3257) );
  INV_X1 U13203 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10652) );
  NOR2_X1 U13204 ( .A1(n10653), .A2(n10652), .ZN(P3_U3259) );
  AOI21_X1 U13205 ( .B1(n14431), .B2(n10660), .A(n10654), .ZN(n10656) );
  INV_X1 U13206 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14299) );
  AOI22_X1 U13207 ( .A1(n10815), .A2(n14299), .B1(P1_REG1_REG_12__SCAN_IN), 
        .B2(n10657), .ZN(n10655) );
  NOR2_X1 U13208 ( .A1(n10656), .A2(n10655), .ZN(n10817) );
  AOI21_X1 U13209 ( .B1(n10656), .B2(n10655), .A(n10817), .ZN(n10669) );
  INV_X1 U13210 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U13211 ( .A1(n10815), .A2(n10658), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n10657), .ZN(n10662) );
  OAI21_X1 U13212 ( .B1(n10660), .B2(n10554), .A(n10659), .ZN(n10661) );
  NOR2_X1 U13213 ( .A1(n10662), .A2(n10661), .ZN(n10809) );
  AOI21_X1 U13214 ( .B1(n10662), .B2(n10661), .A(n10809), .ZN(n10666) );
  INV_X1 U13215 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n11790) );
  NOR2_X1 U13216 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11790), .ZN(n10663) );
  AOI21_X1 U13217 ( .B1(n14468), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n10663), 
        .ZN(n10665) );
  NAND2_X1 U13218 ( .A1(n13792), .A2(n10815), .ZN(n10664) );
  OAI211_X1 U13219 ( .C1(n10666), .C2(n14477), .A(n10665), .B(n10664), .ZN(
        n10667) );
  INV_X1 U13220 ( .A(n10667), .ZN(n10668) );
  OAI21_X1 U13221 ( .B1(n10669), .B2(n14479), .A(n10668), .ZN(P1_U3255) );
  XNOR2_X1 U13222 ( .A(n10671), .B(n10670), .ZN(n10679) );
  INV_X1 U13223 ( .A(n10998), .ZN(n10676) );
  OR2_X1 U13224 ( .A1(n10829), .A2(n13042), .ZN(n10673) );
  NAND2_X1 U13225 ( .A1(n13109), .A2(n13075), .ZN(n10672) );
  NAND2_X1 U13226 ( .A1(n10673), .A2(n10672), .ZN(n11004) );
  NAND2_X1 U13227 ( .A1(n13065), .A2(n11004), .ZN(n10674) );
  OAI211_X1 U13228 ( .C1(n13067), .C2(n10676), .A(n10675), .B(n10674), .ZN(
        n10677) );
  AOI21_X1 U13229 ( .B1(n14821), .B2(n13081), .A(n10677), .ZN(n10678) );
  OAI21_X1 U13230 ( .B1(n10679), .B2(n13083), .A(n10678), .ZN(P2_U3211) );
  INV_X1 U13231 ( .A(P3_DATAO_REG_8__SCAN_IN), .ZN(n15220) );
  NAND2_X1 U13232 ( .A1(n11730), .A2(P3_U3897), .ZN(n10680) );
  OAI21_X1 U13233 ( .B1(P3_U3897), .B2(n15220), .A(n10680), .ZN(P3_U3499) );
  INV_X1 U13234 ( .A(n10681), .ZN(n10682) );
  INV_X1 U13235 ( .A(n11553), .ZN(n14689) );
  OAI222_X1 U13236 ( .A1(n13498), .A2(n7103), .B1(n13505), .B2(n10682), .C1(
        n14689), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U13237 ( .A(n10857), .ZN(n10854) );
  OAI222_X1 U13238 ( .A1(n7001), .A2(n10683), .B1(n14160), .B2(n10682), .C1(
        n10854), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U13239 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n15283) );
  NAND2_X1 U13240 ( .A1(n12486), .A2(P3_U3897), .ZN(n10684) );
  OAI21_X1 U13241 ( .B1(P3_U3897), .B2(n15283), .A(n10684), .ZN(P3_U3505) );
  INV_X1 U13242 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n15411) );
  NAND2_X1 U13243 ( .A1(n10685), .A2(P3_U3897), .ZN(n10686) );
  OAI21_X1 U13244 ( .B1(P3_U3897), .B2(n15411), .A(n10686), .ZN(P3_U3507) );
  INV_X1 U13245 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n15217) );
  NAND2_X1 U13246 ( .A1(n12360), .A2(P3_U3897), .ZN(n10687) );
  OAI21_X1 U13247 ( .B1(P3_U3897), .B2(n15217), .A(n10687), .ZN(P3_U3500) );
  INV_X1 U13248 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n15399) );
  NAND2_X1 U13249 ( .A1(n12455), .A2(P3_U3897), .ZN(n10688) );
  OAI21_X1 U13250 ( .B1(P3_U3897), .B2(n15399), .A(n10688), .ZN(P3_U3503) );
  NAND2_X1 U13251 ( .A1(n10689), .A2(n14837), .ZN(n10690) );
  OAI21_X1 U13252 ( .B1(n14837), .B2(n10224), .A(n10690), .ZN(P2_U3503) );
  XNOR2_X1 U13253 ( .A(n10692), .B(n10691), .ZN(n10699) );
  INV_X1 U13254 ( .A(n14760), .ZN(n10696) );
  OAI22_X1 U13255 ( .A1(n6810), .A2(n13060), .B1(n10693), .B2(n13042), .ZN(
        n10879) );
  AOI21_X1 U13256 ( .B1(n13065), .B2(n10879), .A(n10694), .ZN(n10695) );
  OAI21_X1 U13257 ( .B1(n10696), .B2(n13067), .A(n10695), .ZN(n10697) );
  AOI21_X1 U13258 ( .B1(n12011), .B2(n13081), .A(n10697), .ZN(n10698) );
  OAI21_X1 U13259 ( .B1(n10699), .B2(n13083), .A(n10698), .ZN(P2_U3185) );
  NAND2_X1 U13260 ( .A1(n14558), .A2(n14013), .ZN(n10700) );
  AND2_X1 U13261 ( .A1(n10723), .A2(n10700), .ZN(n14560) );
  INV_X1 U13262 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10701) );
  OAI22_X1 U13263 ( .A1(n14006), .A2(n10432), .B1(n10701), .B2(n13962), .ZN(
        n10705) );
  XOR2_X1 U13264 ( .A(n10702), .B(n10707), .Z(n14564) );
  OAI22_X1 U13265 ( .A1(n14564), .A2(n14009), .B1(n14541), .B2(n10703), .ZN(
        n10704) );
  AOI211_X1 U13266 ( .C1(n14014), .C2(n14560), .A(n10705), .B(n10704), .ZN(
        n10714) );
  OR2_X1 U13267 ( .A1(n14539), .A2(n14408), .ZN(n13966) );
  INV_X1 U13268 ( .A(n13966), .ZN(n14012) );
  OAI21_X1 U13269 ( .B1(n10707), .B2(n10706), .A(n14376), .ZN(n10712) );
  INV_X1 U13270 ( .A(n14560), .ZN(n10708) );
  XNOR2_X1 U13271 ( .A(n10359), .B(n10708), .ZN(n10710) );
  AOI21_X1 U13272 ( .B1(n10710), .B2(n14376), .A(n10709), .ZN(n10711) );
  AOI21_X1 U13273 ( .B1(n14410), .B2(n10712), .A(n10711), .ZN(n14565) );
  AOI22_X1 U13274 ( .A1(n14012), .A2(n9894), .B1(n14565), .B2(n14006), .ZN(
        n10713) );
  NAND2_X1 U13275 ( .A1(n10714), .A2(n10713), .ZN(P1_U3292) );
  XNOR2_X1 U13276 ( .A(n10716), .B(n10715), .ZN(n14573) );
  INV_X1 U13277 ( .A(n14573), .ZN(n10730) );
  NOR2_X1 U13278 ( .A1(n14539), .A2(n10717), .ZN(n14549) );
  INV_X1 U13279 ( .A(n14549), .ZN(n13986) );
  XNOR2_X1 U13280 ( .A(n9890), .B(n10718), .ZN(n10719) );
  NOR2_X1 U13281 ( .A1(n10719), .A2(n14533), .ZN(n10720) );
  AOI211_X1 U13282 ( .C1(n14536), .C2(n14573), .A(n10721), .B(n10720), .ZN(
        n14570) );
  MUX2_X1 U13283 ( .A(n10722), .B(n14570), .S(n14006), .Z(n10729) );
  INV_X1 U13284 ( .A(n10723), .ZN(n10724) );
  OAI211_X1 U13285 ( .C1(n10724), .C2(n14569), .A(n14559), .B(n14543), .ZN(
        n14568) );
  INV_X1 U13286 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10725) );
  OAI22_X1 U13287 ( .A1(n13902), .A2(n14568), .B1(n10725), .B2(n13962), .ZN(
        n10726) );
  AOI21_X1 U13288 ( .B1(n14382), .B2(n10727), .A(n10726), .ZN(n10728) );
  OAI211_X1 U13289 ( .C1(n10730), .C2(n13986), .A(n10729), .B(n10728), .ZN(
        P1_U3291) );
  INV_X1 U13290 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n15423) );
  NAND2_X1 U13291 ( .A1(n12682), .A2(P3_U3897), .ZN(n10731) );
  OAI21_X1 U13292 ( .B1(P3_U3897), .B2(n15423), .A(n10731), .ZN(P3_U3515) );
  NAND2_X1 U13293 ( .A1(n10732), .A2(n14815), .ZN(n10733) );
  XNOR2_X1 U13294 ( .A(n12164), .B(n10734), .ZN(n14794) );
  NAND2_X1 U13295 ( .A1(n14791), .A2(n11972), .ZN(n10735) );
  NAND2_X1 U13296 ( .A1(n10735), .A2(n13359), .ZN(n10736) );
  NOR2_X1 U13297 ( .A1(n10846), .A2(n10736), .ZN(n14790) );
  OAI21_X1 U13298 ( .B1(n10738), .B2(n12164), .A(n10737), .ZN(n10740) );
  AOI21_X1 U13299 ( .B1(n10740), .B2(n13350), .A(n10739), .ZN(n14788) );
  NOR2_X1 U13300 ( .A1(n14788), .A2(n14761), .ZN(n10747) );
  INV_X1 U13301 ( .A(n10741), .ZN(n10742) );
  NOR2_X2 U13302 ( .A1(n14761), .A2(n10742), .ZN(n13366) );
  NAND2_X1 U13303 ( .A1(n13366), .A2(n14791), .ZN(n10745) );
  AOI22_X1 U13304 ( .A1(n14761), .A2(P2_REG2_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(n14759), .ZN(n10744) );
  NAND2_X1 U13305 ( .A1(n10745), .A2(n10744), .ZN(n10746) );
  AOI211_X1 U13306 ( .C1(n14790), .C2(n13338), .A(n10747), .B(n10746), .ZN(
        n10748) );
  OAI21_X1 U13307 ( .B1(n13369), .B2(n14794), .A(n10748), .ZN(P2_U3264) );
  INV_X1 U13308 ( .A(n10749), .ZN(n10750) );
  NAND2_X1 U13309 ( .A1(n10750), .A2(n11204), .ZN(n10784) );
  NAND2_X1 U13310 ( .A1(n10752), .A2(n10751), .ZN(n10753) );
  NAND2_X1 U13311 ( .A1(n10784), .A2(n10782), .ZN(n10781) );
  MUX2_X1 U13312 ( .A(n12506), .B(n10781), .S(n6628), .Z(n14982) );
  INV_X1 U13313 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10755) );
  MUX2_X1 U13314 ( .A(n10755), .B(n10913), .S(n8075), .Z(n10756) );
  INV_X1 U13315 ( .A(n10774), .ZN(n10927) );
  NAND2_X1 U13316 ( .A1(n10756), .A2(n10927), .ZN(n10758) );
  OAI21_X1 U13317 ( .B1(n10756), .B2(n10927), .A(n10758), .ZN(n10922) );
  INV_X1 U13318 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11068) );
  MUX2_X1 U13319 ( .A(n11068), .B(n10757), .S(n11415), .Z(n10791) );
  NAND2_X1 U13320 ( .A1(n10791), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10923) );
  INV_X1 U13321 ( .A(n10758), .ZN(n10765) );
  INV_X1 U13322 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10760) );
  MUX2_X1 U13323 ( .A(n10760), .B(n10759), .S(n11415), .Z(n10761) );
  NAND2_X1 U13324 ( .A1(n10761), .A2(n10773), .ZN(n14843) );
  INV_X1 U13325 ( .A(n10761), .ZN(n10762) );
  NAND2_X1 U13326 ( .A1(n10762), .A2(n7599), .ZN(n10763) );
  AND2_X1 U13327 ( .A1(n14843), .A2(n10763), .ZN(n10764) );
  OAI21_X1 U13328 ( .B1(n10921), .B2(n10765), .A(n10764), .ZN(n14844) );
  INV_X1 U13329 ( .A(n14844), .ZN(n10767) );
  NOR3_X1 U13330 ( .A1(n10921), .A2(n10765), .A3(n10764), .ZN(n10766) );
  AND2_X1 U13331 ( .A1(P3_U3897), .A2(n6628), .ZN(n14960) );
  OAI21_X1 U13332 ( .B1(n10767), .B2(n10766), .A(n14960), .ZN(n10790) );
  INV_X1 U13333 ( .A(n14994), .ZN(n14872) );
  MUX2_X1 U13334 ( .A(n10760), .B(P3_REG2_REG_2__SCAN_IN), .S(n10773), .Z(
        n10772) );
  NAND2_X1 U13335 ( .A1(n10803), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10797) );
  INV_X1 U13336 ( .A(n10797), .ZN(n10769) );
  OR3_X1 U13337 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        n11068), .ZN(n10770) );
  OAI21_X1 U13338 ( .B1(n10774), .B2(n10769), .A(n10770), .ZN(n10909) );
  NAND2_X1 U13339 ( .A1(n10911), .A2(n10770), .ZN(n10771) );
  OAI21_X1 U13340 ( .B1(n10772), .B2(n10771), .A(n11374), .ZN(n10788) );
  MUX2_X1 U13341 ( .A(P3_REG1_REG_2__SCAN_IN), .B(n10759), .S(n10773), .Z(
        n10780) );
  NAND2_X1 U13342 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10803), .ZN(n10796) );
  INV_X1 U13343 ( .A(n10796), .ZN(n10777) );
  OR2_X1 U13344 ( .A1(n10774), .A2(n10777), .ZN(n10776) );
  OR2_X1 U13345 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10796), .ZN(n10775) );
  NAND2_X1 U13346 ( .A1(n10776), .A2(n10775), .ZN(n10914) );
  NOR2_X1 U13347 ( .A1(n10914), .A2(n10913), .ZN(n10912) );
  AOI21_X1 U13348 ( .B1(n10780), .B2(n10779), .A(n11425), .ZN(n10786) );
  OR2_X1 U13349 ( .A1(n10781), .A2(n11420), .ZN(n12604) );
  INV_X1 U13350 ( .A(n10782), .ZN(n10783) );
  AOI22_X1 U13351 ( .A1(n14978), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10785) );
  OAI21_X1 U13352 ( .B1(n10786), .B2(n12604), .A(n10785), .ZN(n10787) );
  AOI21_X1 U13353 ( .B1(n14872), .B2(n10788), .A(n10787), .ZN(n10789) );
  OAI211_X1 U13354 ( .C1(n14982), .C2(n7599), .A(n10790), .B(n10789), .ZN(
        P3_U3184) );
  INV_X1 U13355 ( .A(n10923), .ZN(n10801) );
  NAND3_X1 U13356 ( .A1(n14994), .A2(n12604), .A3(n14986), .ZN(n10800) );
  INV_X1 U13357 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10795) );
  NAND2_X1 U13358 ( .A1(n14978), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n10794) );
  INV_X1 U13359 ( .A(n10791), .ZN(n10792) );
  NAND3_X1 U13360 ( .A1(n14960), .A2(n10792), .A3(n10803), .ZN(n10793) );
  OAI211_X1 U13361 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n10795), .A(n10794), .B(
        n10793), .ZN(n10799) );
  OAI22_X1 U13362 ( .A1(n10797), .A2(n14994), .B1(n12604), .B2(n10796), .ZN(
        n10798) );
  AOI211_X1 U13363 ( .C1(n10801), .C2(n10800), .A(n10799), .B(n10798), .ZN(
        n10802) );
  OAI21_X1 U13364 ( .B1(n10803), .B2(n14982), .A(n10802), .ZN(P3_U3182) );
  INV_X1 U13365 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n10805) );
  NAND2_X1 U13366 ( .A1(n12475), .A2(P3_U3897), .ZN(n10804) );
  OAI21_X1 U13367 ( .B1(P3_U3897), .B2(n10805), .A(n10804), .ZN(P3_U3516) );
  INV_X1 U13368 ( .A(n11350), .ZN(n11363) );
  OAI222_X1 U13369 ( .A1(n7001), .A2(n10806), .B1(n14160), .B2(n10807), .C1(
        n11363), .C2(P1_U3086), .ZN(P1_U3341) );
  INV_X1 U13370 ( .A(n11554), .ZN(n14706) );
  OAI222_X1 U13371 ( .A1(n13498), .A2(n10808), .B1(n13505), .B2(n10807), .C1(
        n14706), .C2(P2_U3088), .ZN(P2_U3313) );
  NOR2_X1 U13372 ( .A1(n10815), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10810) );
  NOR2_X1 U13373 ( .A1(n10810), .A2(n10809), .ZN(n10814) );
  INV_X1 U13374 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10811) );
  MUX2_X1 U13375 ( .A(n10811), .B(P1_REG2_REG_13__SCAN_IN), .S(n10857), .Z(
        n10812) );
  INV_X1 U13376 ( .A(n10812), .ZN(n10813) );
  NAND2_X1 U13377 ( .A1(n10813), .A2(n10814), .ZN(n10858) );
  OAI211_X1 U13378 ( .C1(n10814), .C2(n10813), .A(n14489), .B(n10858), .ZN(
        n10824) );
  NAND2_X1 U13379 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n11876)
         );
  NOR2_X1 U13380 ( .A1(n10815), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10816) );
  NOR2_X1 U13381 ( .A1(n10817), .A2(n10816), .ZN(n10820) );
  INV_X1 U13382 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10818) );
  MUX2_X1 U13383 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10818), .S(n10857), .Z(
        n10819) );
  NAND2_X1 U13384 ( .A1(n10820), .A2(n10819), .ZN(n10853) );
  OAI211_X1 U13385 ( .C1(n10820), .C2(n10819), .A(n14486), .B(n10853), .ZN(
        n10821) );
  NAND2_X1 U13386 ( .A1(n11876), .A2(n10821), .ZN(n10822) );
  AOI21_X1 U13387 ( .B1(n14468), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10822), 
        .ZN(n10823) );
  OAI211_X1 U13388 ( .C1(n14494), .C2(n10854), .A(n10824), .B(n10823), .ZN(
        P1_U3256) );
  XNOR2_X1 U13389 ( .A(n10826), .B(n10825), .ZN(n10827) );
  XNOR2_X1 U13390 ( .A(n10828), .B(n10827), .ZN(n10836) );
  INV_X1 U13391 ( .A(n11145), .ZN(n10833) );
  OAI22_X1 U13392 ( .A1(n10830), .A2(n13042), .B1(n10829), .B2(n13060), .ZN(
        n10931) );
  NAND2_X1 U13393 ( .A1(n13065), .A2(n10931), .ZN(n10831) );
  OAI211_X1 U13394 ( .C1(n13067), .C2(n10833), .A(n10832), .B(n10831), .ZN(
        n10834) );
  AOI21_X1 U13395 ( .B1(n12015), .B2(n13081), .A(n10834), .ZN(n10835) );
  OAI21_X1 U13396 ( .B1(n10836), .B2(n13083), .A(n10835), .ZN(P2_U3193) );
  INV_X1 U13397 ( .A(n10837), .ZN(n10839) );
  INV_X1 U13398 ( .A(n14727), .ZN(n11562) );
  OAI222_X1 U13399 ( .A1(n13498), .A2(n10838), .B1(n13505), .B2(n10839), .C1(
        n11562), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U13400 ( .A(n11360), .ZN(n11630) );
  OAI222_X1 U13401 ( .A1(n7001), .A2(n10840), .B1(n14160), .B2(n10839), .C1(
        n11630), .C2(P1_U3086), .ZN(P1_U3339) );
  XNOR2_X1 U13402 ( .A(n10841), .B(n12165), .ZN(n10843) );
  AOI21_X1 U13403 ( .B1(n10843), .B2(n13350), .A(n10842), .ZN(n14799) );
  INV_X1 U13404 ( .A(n13369), .ZN(n11149) );
  XNOR2_X1 U13405 ( .A(n10845), .B(n10844), .ZN(n14802) );
  OAI211_X1 U13406 ( .C1(n10846), .C2(n6770), .A(n10987), .B(n13359), .ZN(
        n14798) );
  INV_X1 U13407 ( .A(n14798), .ZN(n10847) );
  NAND2_X1 U13408 ( .A1(n13338), .A2(n10847), .ZN(n10850) );
  NAND2_X1 U13409 ( .A1(n13366), .A2(n11983), .ZN(n10849) );
  AOI22_X1 U13410 ( .A1(n14761), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n14759), .ZN(n10848) );
  NAND3_X1 U13411 ( .A1(n10850), .A2(n10849), .A3(n10848), .ZN(n10851) );
  AOI21_X1 U13412 ( .B1(n11149), .B2(n14802), .A(n10851), .ZN(n10852) );
  OAI21_X1 U13413 ( .B1(n14770), .B2(n14799), .A(n10852), .ZN(P2_U3263) );
  INV_X1 U13414 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14420) );
  AOI22_X1 U13415 ( .A1(n11350), .A2(n14420), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n11363), .ZN(n10856) );
  OAI21_X1 U13416 ( .B1(n10854), .B2(n10818), .A(n10853), .ZN(n10855) );
  NOR2_X1 U13417 ( .A1(n10856), .A2(n10855), .ZN(n11362) );
  AOI21_X1 U13418 ( .B1(n10856), .B2(n10855), .A(n11362), .ZN(n10868) );
  NAND2_X1 U13419 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n10857), .ZN(n10859) );
  NAND2_X1 U13420 ( .A1(n10859), .A2(n10858), .ZN(n10863) );
  INV_X1 U13421 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10860) );
  MUX2_X1 U13422 ( .A(n10860), .B(P1_REG2_REG_14__SCAN_IN), .S(n11350), .Z(
        n10861) );
  INV_X1 U13423 ( .A(n10861), .ZN(n10862) );
  NAND2_X1 U13424 ( .A1(n10862), .A2(n10863), .ZN(n11351) );
  OAI211_X1 U13425 ( .C1(n10863), .C2(n10862), .A(n14489), .B(n11351), .ZN(
        n10865) );
  AND2_X1 U13426 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n13522) );
  AOI21_X1 U13427 ( .B1(n14468), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n13522), 
        .ZN(n10864) );
  OAI211_X1 U13428 ( .C1(n14494), .C2(n11363), .A(n10865), .B(n10864), .ZN(
        n10866) );
  INV_X1 U13429 ( .A(n10866), .ZN(n10867) );
  OAI21_X1 U13430 ( .B1(n10868), .B2(n14479), .A(n10867), .ZN(P1_U3257) );
  INV_X1 U13431 ( .A(n13778), .ZN(n11636) );
  OAI222_X1 U13432 ( .A1(n7001), .A2(n10869), .B1(n14160), .B2(n10870), .C1(
        n11636), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U13433 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10871) );
  INV_X1 U13434 ( .A(n14749), .ZN(n11563) );
  OAI222_X1 U13435 ( .A1(n13498), .A2(n10871), .B1(n13505), .B2(n10870), .C1(
        n11563), .C2(P2_U3088), .ZN(P2_U3310) );
  INV_X1 U13436 ( .A(n10872), .ZN(n10874) );
  OAI222_X1 U13437 ( .A1(P3_U3151), .A2(n10875), .B1(n11943), .B2(n10874), 
        .C1(n10873), .C2(n12944), .ZN(P3_U3275) );
  INV_X1 U13438 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15418) );
  OAI21_X1 U13439 ( .B1(n10877), .B2(n12172), .A(n10876), .ZN(n14767) );
  INV_X1 U13440 ( .A(n14767), .ZN(n10884) );
  XOR2_X1 U13441 ( .A(n10878), .B(n12172), .Z(n10880) );
  AOI21_X1 U13442 ( .B1(n10880), .B2(n13350), .A(n10879), .ZN(n14769) );
  INV_X1 U13443 ( .A(n10934), .ZN(n10882) );
  AOI211_X1 U13444 ( .C1(n12011), .C2(n7071), .A(n13336), .B(n10882), .ZN(
        n14758) );
  AOI21_X1 U13445 ( .B1(n14792), .B2(n12011), .A(n14758), .ZN(n10883) );
  OAI211_X1 U13446 ( .C1(n13456), .C2(n10884), .A(n14769), .B(n10883), .ZN(
        n10886) );
  NAND2_X1 U13447 ( .A1(n10886), .A2(n6621), .ZN(n10885) );
  OAI21_X1 U13448 ( .B1(n6621), .B2(n15418), .A(n10885), .ZN(P2_U3451) );
  NAND2_X1 U13449 ( .A1(n10886), .A2(n13457), .ZN(n10887) );
  OAI21_X1 U13450 ( .B1(n14837), .B2(n10233), .A(n10887), .ZN(P2_U3506) );
  OAI211_X1 U13451 ( .C1(n14544), .C2(n10959), .A(n14559), .B(n14523), .ZN(
        n14587) );
  XNOR2_X1 U13452 ( .A(n10892), .B(n10888), .ZN(n10889) );
  NAND2_X1 U13453 ( .A1(n10889), .A2(n14376), .ZN(n14589) );
  OAI21_X1 U13454 ( .B1(n13944), .B2(n14587), .A(n14589), .ZN(n10890) );
  MUX2_X1 U13455 ( .A(n10890), .B(P1_REG2_REG_4__SCAN_IN), .S(n14539), .Z(
        n10896) );
  XNOR2_X1 U13456 ( .A(n10892), .B(n10891), .ZN(n14582) );
  AOI22_X1 U13457 ( .A1(n14382), .A2(n14585), .B1(n10961), .B2(n14538), .ZN(
        n10894) );
  INV_X1 U13458 ( .A(n13849), .ZN(n13960) );
  AOI22_X1 U13459 ( .A1(n13960), .A2(n14583), .B1(n14012), .B2(n14584), .ZN(
        n10893) );
  OAI211_X1 U13460 ( .C1(n14582), .C2(n14009), .A(n10894), .B(n10893), .ZN(
        n10895) );
  OR2_X1 U13461 ( .A1(n10896), .A2(n10895), .ZN(P1_U3289) );
  XNOR2_X1 U13462 ( .A(n10898), .B(n10897), .ZN(n14600) );
  XNOR2_X1 U13463 ( .A(n10899), .B(n10900), .ZN(n10902) );
  OAI22_X1 U13464 ( .A1(n11334), .A2(n14408), .B1(n10958), .B2(n14410), .ZN(
        n11179) );
  INV_X1 U13465 ( .A(n11179), .ZN(n10901) );
  OAI21_X1 U13466 ( .B1(n10902), .B2(n14533), .A(n10901), .ZN(n14605) );
  INV_X1 U13467 ( .A(n14605), .ZN(n10903) );
  MUX2_X1 U13468 ( .A(n10904), .B(n10903), .S(n14006), .Z(n10908) );
  AOI211_X1 U13469 ( .C1(n11180), .C2(n14524), .A(n10341), .B(n14510), .ZN(
        n14603) );
  OAI22_X1 U13470 ( .A1(n14541), .A2(n7323), .B1(n10905), .B2(n13962), .ZN(
        n10906) );
  AOI21_X1 U13471 ( .B1(n14603), .B2(n14548), .A(n10906), .ZN(n10907) );
  OAI211_X1 U13472 ( .C1(n14009), .C2(n14600), .A(n10908), .B(n10907), .ZN(
        P1_U3287) );
  INV_X1 U13473 ( .A(n14982), .ZN(n14915) );
  NAND2_X1 U13474 ( .A1(n10909), .A2(n10755), .ZN(n10910) );
  AND2_X1 U13475 ( .A1(n10911), .A2(n10910), .ZN(n10920) );
  INV_X1 U13476 ( .A(n10912), .ZN(n10916) );
  NAND2_X1 U13477 ( .A1(n10914), .A2(n10913), .ZN(n10915) );
  NAND2_X1 U13478 ( .A1(n10916), .A2(n10915), .ZN(n10917) );
  NAND2_X1 U13479 ( .A1(n14992), .A2(n10917), .ZN(n10919) );
  AOI22_X1 U13480 ( .A1(n14978), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10918) );
  OAI211_X1 U13481 ( .C1(n10920), .C2(n14994), .A(n10919), .B(n10918), .ZN(
        n10926) );
  AOI21_X1 U13482 ( .B1(n10923), .B2(n10922), .A(n10921), .ZN(n10924) );
  NOR2_X1 U13483 ( .A1(n10924), .A2(n14986), .ZN(n10925) );
  AOI211_X1 U13484 ( .C1(n14915), .C2(n10927), .A(n10926), .B(n10925), .ZN(
        n10928) );
  INV_X1 U13485 ( .A(n10928), .ZN(P3_U3183) );
  OAI21_X1 U13486 ( .B1(n6655), .B2(n7284), .A(n10929), .ZN(n11143) );
  AOI21_X1 U13487 ( .B1(n10930), .B2(n7284), .A(n13332), .ZN(n10933) );
  AOI21_X1 U13488 ( .B1(n10933), .B2(n10932), .A(n10931), .ZN(n11152) );
  NAND2_X1 U13489 ( .A1(n12015), .A2(n10934), .ZN(n10935) );
  AND3_X1 U13490 ( .A1(n11096), .A2(n13359), .A3(n10935), .ZN(n11144) );
  AOI21_X1 U13491 ( .B1(n14792), .B2(n12015), .A(n11144), .ZN(n10936) );
  OAI211_X1 U13492 ( .C1(n11143), .C2(n13456), .A(n11152), .B(n10936), .ZN(
        n10939) );
  NAND2_X1 U13493 ( .A1(n10939), .A2(n13457), .ZN(n10937) );
  OAI21_X1 U13494 ( .B1(n14837), .B2(n10938), .A(n10937), .ZN(P2_U3507) );
  INV_X1 U13495 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10941) );
  NAND2_X1 U13496 ( .A1(n10939), .A2(n6621), .ZN(n10940) );
  OAI21_X1 U13497 ( .B1(n6621), .B2(n10941), .A(n10940), .ZN(P2_U3454) );
  OAI22_X1 U13498 ( .A1(n11038), .A2(n10612), .B1(n10959), .B2(n10348), .ZN(
        n10942) );
  XOR2_X1 U13499 ( .A(n12323), .B(n10942), .Z(n10957) );
  INV_X1 U13500 ( .A(n10943), .ZN(n10945) );
  AOI22_X1 U13501 ( .A1(n12321), .A2(n14583), .B1(n10603), .B2(n6626), .ZN(
        n10950) );
  AOI22_X1 U13502 ( .A1(n14583), .A2(n10603), .B1(n12320), .B2(n13538), .ZN(
        n10948) );
  XNOR2_X1 U13503 ( .A(n10948), .B(n11327), .ZN(n10949) );
  XOR2_X1 U13504 ( .A(n10950), .B(n10949), .Z(n13536) );
  INV_X1 U13505 ( .A(n10949), .ZN(n10952) );
  INV_X1 U13506 ( .A(n12321), .ZN(n10954) );
  OR2_X1 U13507 ( .A1(n11038), .A2(n10954), .ZN(n10955) );
  OAI21_X1 U13508 ( .B1(n10959), .B2(n10612), .A(n10955), .ZN(n11028) );
  AOI211_X1 U13509 ( .C1(n10957), .C2(n10956), .A(n13660), .B(n11033), .ZN(
        n10967) );
  OAI22_X1 U13510 ( .A1(n13640), .A2(n10959), .B1(n13647), .B2(n10958), .ZN(
        n10966) );
  INV_X1 U13511 ( .A(n13645), .ZN(n13654) );
  NAND2_X1 U13512 ( .A1(n13654), .A2(n10961), .ZN(n10962) );
  OAI211_X1 U13513 ( .C1(n13646), .C2(n10964), .A(n10963), .B(n10962), .ZN(
        n10965) );
  OR3_X1 U13514 ( .A1(n10967), .A2(n10966), .A3(n10965), .ZN(P1_U3230) );
  XNOR2_X1 U13515 ( .A(n11999), .B(n13109), .ZN(n12169) );
  XNOR2_X1 U13516 ( .A(n10968), .B(n12169), .ZN(n14816) );
  XNOR2_X1 U13517 ( .A(n10969), .B(n12169), .ZN(n10971) );
  AOI21_X1 U13518 ( .B1(n10971), .B2(n13350), .A(n10970), .ZN(n14818) );
  MUX2_X1 U13519 ( .A(n10972), .B(n14818), .S(n13357), .Z(n10978) );
  INV_X1 U13520 ( .A(n13338), .ZN(n13363) );
  OAI211_X1 U13521 ( .C1(n14812), .C2(n10973), .A(n13359), .B(n10996), .ZN(
        n14811) );
  AOI22_X1 U13522 ( .A1(n13366), .A2(n11999), .B1(n14759), .B2(n10974), .ZN(
        n10975) );
  OAI21_X1 U13523 ( .B1(n13363), .B2(n14811), .A(n10975), .ZN(n10976) );
  INV_X1 U13524 ( .A(n10976), .ZN(n10977) );
  OAI211_X1 U13525 ( .C1(n13369), .C2(n14816), .A(n10978), .B(n10977), .ZN(
        P2_U3260) );
  INV_X1 U13526 ( .A(n10979), .ZN(n10982) );
  OAI222_X1 U13527 ( .A1(n11943), .A2(n10982), .B1(n12944), .B2(n10981), .C1(
        P3_U3151), .C2(n10980), .ZN(P3_U3274) );
  XNOR2_X1 U13528 ( .A(n10983), .B(n8980), .ZN(n10985) );
  AOI21_X1 U13529 ( .B1(n10985), .B2(n13350), .A(n10984), .ZN(n14805) );
  XNOR2_X1 U13530 ( .A(n12167), .B(n10986), .ZN(n14809) );
  OAI211_X1 U13531 ( .C1(n7068), .C2(n7498), .A(n13359), .B(n10988), .ZN(
        n14804) );
  OAI22_X1 U13532 ( .A1(n13357), .A2(n10245), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n13354), .ZN(n10989) );
  AOI21_X1 U13533 ( .B1(n13366), .B2(n11987), .A(n10989), .ZN(n10990) );
  OAI21_X1 U13534 ( .B1(n13363), .B2(n14804), .A(n10990), .ZN(n10991) );
  AOI21_X1 U13535 ( .B1(n11149), .B2(n14809), .A(n10991), .ZN(n10992) );
  OAI21_X1 U13536 ( .B1(n14770), .B2(n14805), .A(n10992), .ZN(P2_U3262) );
  INV_X1 U13537 ( .A(n10993), .ZN(n11011) );
  OAI21_X1 U13538 ( .B1(n10995), .B2(n11000), .A(n10994), .ZN(n14823) );
  NAND2_X1 U13539 ( .A1(n14821), .A2(n10996), .ZN(n10997) );
  NAND3_X1 U13540 ( .A1(n7071), .A2(n13359), .A3(n10997), .ZN(n14824) );
  AOI22_X1 U13541 ( .A1(n13366), .A2(n14821), .B1(n14759), .B2(n10998), .ZN(
        n10999) );
  OAI21_X1 U13542 ( .B1(n13363), .B2(n14824), .A(n10999), .ZN(n11010) );
  NAND2_X1 U13543 ( .A1(n11001), .A2(n11000), .ZN(n11002) );
  NAND2_X1 U13544 ( .A1(n11003), .A2(n11002), .ZN(n11005) );
  AOI21_X1 U13545 ( .B1(n11005), .B2(n13350), .A(n11004), .ZN(n11008) );
  NAND2_X1 U13546 ( .A1(n14823), .A2(n11006), .ZN(n11007) );
  NAND2_X1 U13547 ( .A1(n11008), .A2(n11007), .ZN(n14827) );
  MUX2_X1 U13548 ( .A(n14827), .B(P2_REG2_REG_6__SCAN_IN), .S(n14761), .Z(
        n11009) );
  AOI211_X1 U13549 ( .C1(n11011), .C2(n14823), .A(n11010), .B(n11009), .ZN(
        n11012) );
  INV_X1 U13550 ( .A(n11012), .ZN(P2_U3259) );
  NAND2_X1 U13551 ( .A1(n12506), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n11013) );
  OAI21_X1 U13552 ( .B1(n11014), .B2(n12506), .A(n11013), .ZN(P3_U3521) );
  INV_X1 U13553 ( .A(n11015), .ZN(n11017) );
  INV_X1 U13554 ( .A(n11364), .ZN(n14480) );
  OAI222_X1 U13555 ( .A1(n7001), .A2(n11016), .B1(n14160), .B2(n11017), .C1(
        P1_U3086), .C2(n14480), .ZN(P1_U3340) );
  INV_X1 U13556 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11018) );
  INV_X1 U13557 ( .A(n11559), .ZN(n14721) );
  OAI222_X1 U13558 ( .A1(n13498), .A2(n11018), .B1(n13505), .B2(n11017), .C1(
        P2_U3088), .C2(n14721), .ZN(P2_U3312) );
  XOR2_X1 U13559 ( .A(n11021), .B(n11020), .Z(n11026) );
  AOI22_X1 U13560 ( .A1(n13075), .A2(n13106), .B1(n13104), .B2(n13076), .ZN(
        n11093) );
  OAI22_X1 U13561 ( .A1(n13079), .A2(n11093), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11022), .ZN(n11024) );
  NOR2_X1 U13562 ( .A1(n11099), .A2(n8914), .ZN(n11023) );
  AOI211_X1 U13563 ( .C1(n13077), .C2(n11097), .A(n11024), .B(n11023), .ZN(
        n11025) );
  OAI21_X1 U13564 ( .B1(n11026), .B2(n13083), .A(n11025), .ZN(P2_U3203) );
  INV_X1 U13565 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n15424) );
  NAND2_X1 U13566 ( .A1(n12614), .A2(P3_U3897), .ZN(n11027) );
  OAI21_X1 U13567 ( .B1(P3_U3897), .B2(n15424), .A(n11027), .ZN(P3_U3522) );
  INV_X1 U13568 ( .A(n11028), .ZN(n11031) );
  AOI22_X1 U13569 ( .A1(n11040), .A2(n12320), .B1(n12322), .B2(n14584), .ZN(
        n11034) );
  XOR2_X1 U13570 ( .A(n12323), .B(n11034), .Z(n11168) );
  NAND2_X1 U13571 ( .A1(n11040), .A2(n12322), .ZN(n11036) );
  NAND2_X1 U13572 ( .A1(n12321), .A2(n14584), .ZN(n11035) );
  NAND2_X1 U13573 ( .A1(n11036), .A2(n11035), .ZN(n11172) );
  XNOR2_X1 U13574 ( .A(n11168), .B(n11172), .ZN(n11037) );
  XNOR2_X1 U13575 ( .A(n11173), .B(n11037), .ZN(n11043) );
  OAI22_X1 U13576 ( .A1(n11039), .A2(n14408), .B1(n11038), .B2(n14410), .ZN(
        n14519) );
  AOI22_X1 U13577 ( .A1(n13540), .A2(n14519), .B1(P1_REG3_REG_5__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11042) );
  AOI22_X1 U13578 ( .A1(n14520), .A2(n13654), .B1(n13658), .B2(n11040), .ZN(
        n11041) );
  OAI211_X1 U13579 ( .C1(n11043), .C2(n13660), .A(n11042), .B(n11041), .ZN(
        P1_U3227) );
  XOR2_X1 U13580 ( .A(n11045), .B(n11044), .Z(n11051) );
  NAND2_X1 U13581 ( .A1(n11047), .A2(n11046), .ZN(n11946) );
  NOR2_X1 U13582 ( .A1(n12465), .A2(n7578), .ZN(n11049) );
  INV_X1 U13583 ( .A(n12504), .ZN(n15044) );
  OAI22_X1 U13584 ( .A1(n12485), .A2(n15050), .B1(n15044), .B2(n12490), .ZN(
        n11048) );
  AOI211_X1 U13585 ( .C1(n11946), .C2(P3_REG3_REG_2__SCAN_IN), .A(n11049), .B(
        n11048), .ZN(n11050) );
  OAI21_X1 U13586 ( .B1(n11051), .B2(n12495), .A(n11050), .ZN(P3_U3177) );
  NOR2_X1 U13587 ( .A1(n12944), .A2(SI_22_), .ZN(n11052) );
  AOI21_X1 U13588 ( .B1(n11053), .B2(P3_STATE_REG_SCAN_IN), .A(n11052), .ZN(
        n11054) );
  OAI21_X1 U13589 ( .B1(n11055), .B2(n11943), .A(n11054), .ZN(n11056) );
  INV_X1 U13590 ( .A(n11056), .ZN(P3_U3273) );
  AOI21_X1 U13591 ( .B1(n15016), .B2(n11057), .A(n11950), .ZN(n11058) );
  AOI21_X1 U13592 ( .B1(n15059), .B2(n12505), .A(n11058), .ZN(n11957) );
  INV_X1 U13593 ( .A(n11059), .ZN(n11060) );
  OAI21_X1 U13594 ( .B1(n11939), .B2(n11060), .A(n11061), .ZN(n11065) );
  INV_X1 U13595 ( .A(n11061), .ZN(n11062) );
  NAND2_X1 U13596 ( .A1(n11063), .A2(n11062), .ZN(n11064) );
  AND2_X1 U13597 ( .A1(n11065), .A2(n11064), .ZN(n11067) );
  MUX2_X1 U13598 ( .A(n11068), .B(n11957), .S(n15074), .Z(n11071) );
  INV_X1 U13599 ( .A(n12818), .ZN(n12770) );
  AOI22_X1 U13600 ( .A1(n12770), .A2(n11947), .B1(n15071), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n11070) );
  NAND2_X1 U13601 ( .A1(n11071), .A2(n11070), .ZN(P3_U3233) );
  INV_X1 U13602 ( .A(n15064), .ZN(n11076) );
  NOR3_X1 U13603 ( .A1(n11072), .A2(n9131), .A3(n12335), .ZN(n11074) );
  AOI211_X1 U13604 ( .C1(n11076), .C2(n11075), .A(n11074), .B(n11073), .ZN(
        n11080) );
  OAI22_X1 U13605 ( .A1(n12485), .A2(n15057), .B1(n11242), .B2(n12490), .ZN(
        n11077) );
  AOI21_X1 U13606 ( .B1(n12487), .B2(n15061), .A(n11077), .ZN(n11079) );
  NAND2_X1 U13607 ( .A1(n11946), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n11078) );
  OAI211_X1 U13608 ( .C1(n11080), .C2(n12495), .A(n11079), .B(n11078), .ZN(
        P3_U3162) );
  INV_X1 U13609 ( .A(n13031), .ZN(n11082) );
  INV_X1 U13610 ( .A(n13030), .ZN(n11081) );
  OAI22_X1 U13611 ( .A1(n14764), .A2(n11082), .B1(n13354), .B2(n11081), .ZN(
        n11083) );
  AOI21_X1 U13612 ( .B1(n14757), .B2(n11084), .A(n11083), .ZN(n11087) );
  MUX2_X1 U13613 ( .A(n10246), .B(n11085), .S(n13357), .Z(n11086) );
  OAI211_X1 U13614 ( .C1(n13369), .C2(n11088), .A(n11087), .B(n11086), .ZN(
        P2_U3261) );
  XNOR2_X1 U13615 ( .A(n11090), .B(n11089), .ZN(n11188) );
  OAI211_X1 U13616 ( .C1(n11092), .C2(n12174), .A(n11091), .B(n13350), .ZN(
        n11094) );
  NAND2_X1 U13617 ( .A1(n11094), .A2(n11093), .ZN(n11185) );
  NAND2_X1 U13618 ( .A1(n11185), .A2(n13357), .ZN(n11102) );
  INV_X1 U13619 ( .A(n11133), .ZN(n11095) );
  AOI211_X1 U13620 ( .C1(n12019), .C2(n11096), .A(n13336), .B(n11095), .ZN(
        n11186) );
  AOI22_X1 U13621 ( .A1(n14761), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n11097), 
        .B2(n14759), .ZN(n11098) );
  OAI21_X1 U13622 ( .B1(n11099), .B2(n14764), .A(n11098), .ZN(n11100) );
  AOI21_X1 U13623 ( .B1(n11186), .B2(n14757), .A(n11100), .ZN(n11101) );
  OAI211_X1 U13624 ( .C1(n13369), .C2(n11188), .A(n11102), .B(n11101), .ZN(
        P2_U3256) );
  XNOR2_X1 U13625 ( .A(n11104), .B(n11103), .ZN(n14615) );
  NAND2_X1 U13626 ( .A1(n14509), .A2(n11338), .ZN(n11105) );
  NAND3_X1 U13627 ( .A1(n11106), .A2(n14559), .A3(n11105), .ZN(n14619) );
  AOI21_X1 U13628 ( .B1(n11108), .B2(n11107), .A(n14533), .ZN(n11110) );
  NAND2_X1 U13629 ( .A1(n11110), .A2(n11109), .ZN(n14620) );
  OAI21_X1 U13630 ( .B1(n13944), .B2(n14619), .A(n14620), .ZN(n11111) );
  MUX2_X1 U13631 ( .A(n11111), .B(P1_REG2_REG_8__SCAN_IN), .S(n14539), .Z(
        n11112) );
  INV_X1 U13632 ( .A(n11112), .ZN(n11117) );
  NOR2_X1 U13633 ( .A1(n13966), .A2(n11678), .ZN(n11115) );
  INV_X1 U13634 ( .A(n11337), .ZN(n11113) );
  OAI22_X1 U13635 ( .A1(n13849), .A2(n11334), .B1(n11113), .B2(n13962), .ZN(
        n11114) );
  AOI211_X1 U13636 ( .C1(n14382), .C2(n11338), .A(n11115), .B(n11114), .ZN(
        n11116) );
  OAI211_X1 U13637 ( .C1(n14615), .C2(n14009), .A(n11117), .B(n11116), .ZN(
        P1_U3285) );
  INV_X1 U13638 ( .A(n12022), .ZN(n11136) );
  AOI21_X1 U13639 ( .B1(n11119), .B2(n11118), .A(n13083), .ZN(n11121) );
  NAND2_X1 U13640 ( .A1(n11121), .A2(n11120), .ZN(n11125) );
  AOI22_X1 U13641 ( .A1(n13076), .A2(n13103), .B1(n13105), .B2(n13075), .ZN(
        n11130) );
  OAI21_X1 U13642 ( .B1(n13079), .B2(n11130), .A(n11122), .ZN(n11123) );
  AOI21_X1 U13643 ( .B1(n11134), .B2(n13077), .A(n11123), .ZN(n11124) );
  OAI211_X1 U13644 ( .C1(n11136), .C2(n8914), .A(n11125), .B(n11124), .ZN(
        P2_U3189) );
  XNOR2_X1 U13645 ( .A(n11127), .B(n11126), .ZN(n11232) );
  OAI211_X1 U13646 ( .C1(n11129), .C2(n12176), .A(n11128), .B(n13350), .ZN(
        n11131) );
  NAND2_X1 U13647 ( .A1(n11131), .A2(n11130), .ZN(n11229) );
  NAND2_X1 U13648 ( .A1(n11229), .A2(n13357), .ZN(n11139) );
  INV_X1 U13649 ( .A(n11264), .ZN(n11132) );
  AOI211_X1 U13650 ( .C1(n12022), .C2(n11133), .A(n13336), .B(n11132), .ZN(
        n11230) );
  AOI22_X1 U13651 ( .A1(n14761), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11134), 
        .B2(n14759), .ZN(n11135) );
  OAI21_X1 U13652 ( .B1(n11136), .B2(n14764), .A(n11135), .ZN(n11137) );
  AOI21_X1 U13653 ( .B1(n11230), .B2(n14757), .A(n11137), .ZN(n11138) );
  OAI211_X1 U13654 ( .C1(n13369), .C2(n11232), .A(n11139), .B(n11138), .ZN(
        P2_U3255) );
  INV_X1 U13655 ( .A(n13136), .ZN(n11570) );
  OAI222_X1 U13656 ( .A1(n13498), .A2(n11140), .B1(n13505), .B2(n11141), .C1(
        n11570), .C2(P2_U3088), .ZN(P2_U3309) );
  INV_X1 U13657 ( .A(n13787), .ZN(n14493) );
  OAI222_X1 U13658 ( .A1(n7001), .A2(n11142), .B1(n14160), .B2(n11141), .C1(
        n14493), .C2(P1_U3086), .ZN(P1_U3337) );
  INV_X1 U13659 ( .A(n11143), .ZN(n11150) );
  NAND2_X1 U13660 ( .A1(n11144), .A2(n14757), .ZN(n11147) );
  AOI22_X1 U13661 ( .A1(n14761), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n11145), 
        .B2(n14759), .ZN(n11146) );
  OAI211_X1 U13662 ( .C1(n7070), .C2(n14764), .A(n11147), .B(n11146), .ZN(
        n11148) );
  AOI21_X1 U13663 ( .B1(n11150), .B2(n11149), .A(n11148), .ZN(n11151) );
  OAI21_X1 U13664 ( .B1(n14770), .B2(n11152), .A(n11151), .ZN(P2_U3257) );
  XNOR2_X1 U13665 ( .A(n11153), .B(n11155), .ZN(n11160) );
  OAI21_X1 U13666 ( .B1(n11156), .B2(n11155), .A(n11154), .ZN(n11158) );
  OAI22_X1 U13667 ( .A1(n11608), .A2(n14408), .B1(n11607), .B2(n14410), .ZN(
        n11157) );
  AOI21_X1 U13668 ( .B1(n11158), .B2(n14376), .A(n11157), .ZN(n11159) );
  OAI21_X1 U13669 ( .B1(n14602), .B2(n11160), .A(n11159), .ZN(n14628) );
  INV_X1 U13670 ( .A(n14628), .ZN(n11167) );
  INV_X1 U13671 ( .A(n11160), .ZN(n14630) );
  OAI211_X1 U13672 ( .C1(n14627), .C2(n11161), .A(n14559), .B(n11312), .ZN(
        n14625) );
  AOI22_X1 U13673 ( .A1(n14539), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n11611), 
        .B2(n14538), .ZN(n11164) );
  NAND2_X1 U13674 ( .A1(n11162), .A2(n14382), .ZN(n11163) );
  OAI211_X1 U13675 ( .C1(n14625), .C2(n13902), .A(n11164), .B(n11163), .ZN(
        n11165) );
  AOI21_X1 U13676 ( .B1(n14630), .B2(n14549), .A(n11165), .ZN(n11166) );
  OAI21_X1 U13677 ( .B1(n11167), .B2(n14539), .A(n11166), .ZN(P1_U3284) );
  INV_X1 U13678 ( .A(n11172), .ZN(n11170) );
  INV_X1 U13679 ( .A(n11168), .ZN(n11169) );
  AOI21_X1 U13680 ( .B1(n11173), .B2(n11170), .A(n11169), .ZN(n11171) );
  INV_X1 U13681 ( .A(n11171), .ZN(n11175) );
  AND2_X1 U13682 ( .A1(n12321), .A2(n13670), .ZN(n11176) );
  AOI21_X1 U13683 ( .B1(n11180), .B2(n12322), .A(n11176), .ZN(n11210) );
  AOI22_X1 U13684 ( .A1(n11180), .A2(n12320), .B1(n12322), .B2(n13670), .ZN(
        n11178) );
  INV_X2 U13685 ( .A(n11177), .ZN(n12323) );
  XNOR2_X1 U13686 ( .A(n11178), .B(n12323), .ZN(n11209) );
  XOR2_X1 U13687 ( .A(n11210), .B(n11209), .Z(n11213) );
  XNOR2_X1 U13688 ( .A(n6774), .B(n11213), .ZN(n11184) );
  AND2_X1 U13689 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n13736) );
  AOI21_X1 U13690 ( .B1(n13540), .B2(n11179), .A(n13736), .ZN(n11183) );
  AOI22_X1 U13691 ( .A1(n11181), .A2(n13654), .B1(n13658), .B2(n11180), .ZN(
        n11182) );
  OAI211_X1 U13692 ( .C1(n11184), .C2(n13660), .A(n11183), .B(n11182), .ZN(
        P1_U3239) );
  AOI211_X1 U13693 ( .C1(n14792), .C2(n12019), .A(n11186), .B(n11185), .ZN(
        n11187) );
  OAI21_X1 U13694 ( .B1(n13456), .B2(n11188), .A(n11187), .ZN(n11191) );
  NAND2_X1 U13695 ( .A1(n11191), .A2(n13457), .ZN(n11189) );
  OAI21_X1 U13696 ( .B1(n13457), .B2(n11190), .A(n11189), .ZN(P2_U3508) );
  INV_X1 U13697 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11193) );
  NAND2_X1 U13698 ( .A1(n11191), .A2(n6621), .ZN(n11192) );
  OAI21_X1 U13699 ( .B1(n6621), .B2(n11193), .A(n11192), .ZN(P2_U3457) );
  INV_X1 U13700 ( .A(n12031), .ZN(n11270) );
  OAI211_X1 U13701 ( .C1(n11196), .C2(n11195), .A(n11194), .B(n13049), .ZN(
        n11200) );
  AOI22_X1 U13702 ( .A1(n13102), .A2(n13076), .B1(n13075), .B2(n13104), .ZN(
        n11262) );
  OAI21_X1 U13703 ( .B1(n13079), .B2(n11262), .A(n11197), .ZN(n11198) );
  AOI21_X1 U13704 ( .B1(n11267), .B2(n13077), .A(n11198), .ZN(n11199) );
  OAI211_X1 U13705 ( .C1(n11270), .C2(n8914), .A(n11200), .B(n11199), .ZN(
        P2_U3208) );
  OAI222_X1 U13706 ( .A1(n7001), .A2(n11202), .B1(n14160), .B2(n11207), .C1(
        n11201), .C2(P1_U3086), .ZN(P1_U3335) );
  NAND2_X1 U13707 ( .A1(n11203), .A2(n12933), .ZN(n11205) );
  OAI211_X1 U13708 ( .C1(n11206), .C2(n12944), .A(n11205), .B(n11204), .ZN(
        P3_U3272) );
  OAI222_X1 U13709 ( .A1(n13498), .A2(n7920), .B1(P2_U3088), .B2(n11208), .C1(
        n13505), .C2(n11207), .ZN(P2_U3307) );
  INV_X1 U13710 ( .A(n11209), .ZN(n11212) );
  INV_X1 U13711 ( .A(n11210), .ZN(n11211) );
  AOI22_X1 U13712 ( .A1(n11217), .A2(n12320), .B1(n12322), .B2(n14616), .ZN(
        n11215) );
  XNOR2_X1 U13713 ( .A(n11215), .B(n12323), .ZN(n11321) );
  AND2_X1 U13714 ( .A1(n12321), .A2(n14616), .ZN(n11216) );
  AOI21_X1 U13715 ( .B1(n11217), .B2(n12322), .A(n11216), .ZN(n11322) );
  XNOR2_X1 U13716 ( .A(n11321), .B(n11322), .ZN(n11323) );
  XNOR2_X1 U13717 ( .A(n11324), .B(n11323), .ZN(n11224) );
  OR2_X1 U13718 ( .A1(n11607), .A2(n14408), .ZN(n11219) );
  NAND2_X1 U13719 ( .A1(n13670), .A2(n14634), .ZN(n11218) );
  AND2_X1 U13720 ( .A1(n11219), .A2(n11218), .ZN(n14503) );
  OAI21_X1 U13721 ( .B1(n13656), .B2(n14503), .A(n11220), .ZN(n11222) );
  NOR2_X1 U13722 ( .A1(n13640), .A2(n14609), .ZN(n11221) );
  AOI211_X1 U13723 ( .C1(n13654), .C2(n14506), .A(n11222), .B(n11221), .ZN(
        n11223) );
  OAI21_X1 U13724 ( .B1(n11224), .B2(n13660), .A(n11223), .ZN(P1_U3213) );
  INV_X1 U13725 ( .A(n11225), .ZN(n11227) );
  OAI222_X1 U13726 ( .A1(n13498), .A2(n11226), .B1(n13505), .B2(n11227), .C1(
        n8904), .C2(P2_U3088), .ZN(P2_U3308) );
  OAI222_X1 U13727 ( .A1(n7001), .A2(n11228), .B1(n14160), .B2(n11227), .C1(
        P1_U3086), .C2(n13930), .ZN(P1_U3336) );
  AOI211_X1 U13728 ( .C1(n14792), .C2(n12022), .A(n11230), .B(n11229), .ZN(
        n11231) );
  OAI21_X1 U13729 ( .B1(n13456), .B2(n11232), .A(n11231), .ZN(n11235) );
  NAND2_X1 U13730 ( .A1(n11235), .A2(n13457), .ZN(n11233) );
  OAI21_X1 U13731 ( .B1(n13457), .B2(n11234), .A(n11233), .ZN(P2_U3509) );
  INV_X1 U13732 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n11237) );
  NAND2_X1 U13733 ( .A1(n11235), .A2(n6621), .ZN(n11236) );
  OAI21_X1 U13734 ( .B1(n6621), .B2(n11237), .A(n11236), .ZN(P2_U3460) );
  AOI211_X1 U13735 ( .C1(n11240), .C2(n11239), .A(n12495), .B(n11238), .ZN(
        n11241) );
  INV_X1 U13736 ( .A(n11241), .ZN(n11246) );
  NOR2_X1 U13737 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7604), .ZN(n14840) );
  INV_X1 U13738 ( .A(n15026), .ZN(n15017) );
  OAI22_X1 U13739 ( .A1(n12465), .A2(n11242), .B1(n15017), .B2(n12490), .ZN(
        n11243) );
  AOI211_X1 U13740 ( .C1(n11244), .C2(n12467), .A(n14840), .B(n11243), .ZN(
        n11245) );
  OAI211_X1 U13741 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n11768), .A(n11246), .B(
        n11245), .ZN(P3_U3158) );
  NAND2_X1 U13742 ( .A1(n11248), .A2(n11247), .ZN(n11250) );
  XOR2_X1 U13743 ( .A(n11250), .B(n11249), .Z(n11256) );
  INV_X1 U13744 ( .A(n11299), .ZN(n11253) );
  OAI22_X1 U13745 ( .A1(n11251), .A2(n13060), .B1(n11579), .B2(n13042), .ZN(
        n11295) );
  AOI22_X1 U13746 ( .A1(n13065), .A2(n11295), .B1(P2_REG3_REG_12__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11252) );
  OAI21_X1 U13747 ( .B1(n11253), .B2(n13067), .A(n11252), .ZN(n11254) );
  AOI21_X1 U13748 ( .B1(n12035), .B2(n13081), .A(n11254), .ZN(n11255) );
  OAI21_X1 U13749 ( .B1(n11256), .B2(n13083), .A(n11255), .ZN(P2_U3196) );
  XNOR2_X1 U13750 ( .A(n11257), .B(n11261), .ZN(n11478) );
  INV_X1 U13751 ( .A(n11258), .ZN(n11259) );
  AOI21_X1 U13752 ( .B1(n11261), .B2(n11260), .A(n11259), .ZN(n11263) );
  OAI21_X1 U13753 ( .B1(n11263), .B2(n13332), .A(n11262), .ZN(n11475) );
  NAND2_X1 U13754 ( .A1(n12031), .A2(n11264), .ZN(n11265) );
  NAND2_X1 U13755 ( .A1(n11265), .A2(n13359), .ZN(n11266) );
  NOR2_X1 U13756 ( .A1(n11298), .A2(n11266), .ZN(n11476) );
  NAND2_X1 U13757 ( .A1(n11476), .A2(n14757), .ZN(n11269) );
  AOI22_X1 U13758 ( .A1(n14761), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11267), 
        .B2(n14759), .ZN(n11268) );
  OAI211_X1 U13759 ( .C1(n11270), .C2(n14764), .A(n11269), .B(n11268), .ZN(
        n11271) );
  AOI21_X1 U13760 ( .B1(n11475), .B2(n13357), .A(n11271), .ZN(n11272) );
  OAI21_X1 U13761 ( .B1(n13369), .B2(n11478), .A(n11272), .ZN(P2_U3254) );
  INV_X1 U13762 ( .A(n11459), .ZN(n11281) );
  OAI21_X1 U13763 ( .B1(n11275), .B2(n11274), .A(n11273), .ZN(n11276) );
  NAND2_X1 U13764 ( .A1(n11276), .A2(n12473), .ZN(n11280) );
  NAND2_X1 U13765 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n14877) );
  INV_X1 U13766 ( .A(n14877), .ZN(n11278) );
  OAI22_X1 U13767 ( .A1(n12485), .A2(n11458), .B1(n12465), .B2(n15044), .ZN(
        n11277) );
  AOI211_X1 U13768 ( .C1(n12462), .C2(n15002), .A(n11278), .B(n11277), .ZN(
        n11279) );
  OAI211_X1 U13769 ( .C1(n11281), .C2(n11768), .A(n11280), .B(n11279), .ZN(
        P3_U3170) );
  OAI222_X1 U13770 ( .A1(n7001), .A2(n11282), .B1(n14160), .B2(n11283), .C1(
        n9882), .C2(P1_U3086), .ZN(P1_U3334) );
  OAI222_X1 U13771 ( .A1(n13498), .A2(n11285), .B1(P2_U3088), .B2(n11284), 
        .C1(n13505), .C2(n11283), .ZN(P2_U3306) );
  XNOR2_X1 U13772 ( .A(n11287), .B(n11288), .ZN(n11292) );
  AND2_X1 U13773 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n14691) );
  AOI22_X1 U13774 ( .A1(n13102), .A2(n13075), .B1(n13076), .B2(n13100), .ZN(
        n11504) );
  NOR2_X1 U13775 ( .A1(n13079), .A2(n11504), .ZN(n11289) );
  AOI211_X1 U13776 ( .C1(n13077), .C2(n11508), .A(n14691), .B(n11289), .ZN(
        n11291) );
  NAND2_X1 U13777 ( .A1(n12044), .A2(n13081), .ZN(n11290) );
  OAI211_X1 U13778 ( .C1(n11292), .C2(n13083), .A(n11291), .B(n11290), .ZN(
        P2_U3206) );
  XOR2_X1 U13779 ( .A(n11293), .B(n12178), .Z(n11488) );
  INV_X1 U13780 ( .A(n11488), .ZN(n11305) );
  AOI21_X1 U13781 ( .B1(n11294), .B2(n12178), .A(n13332), .ZN(n11297) );
  AOI21_X1 U13782 ( .B1(n11297), .B2(n11296), .A(n11295), .ZN(n11485) );
  INV_X1 U13783 ( .A(n11485), .ZN(n11303) );
  OAI211_X1 U13784 ( .C1(n11486), .C2(n11298), .A(n13359), .B(n11506), .ZN(
        n11484) );
  AOI22_X1 U13785 ( .A1(n14761), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11299), 
        .B2(n14759), .ZN(n11301) );
  NAND2_X1 U13786 ( .A1(n12035), .A2(n13366), .ZN(n11300) );
  OAI211_X1 U13787 ( .C1(n11484), .C2(n13363), .A(n11301), .B(n11300), .ZN(
        n11302) );
  AOI21_X1 U13788 ( .B1(n11303), .B2(n13357), .A(n11302), .ZN(n11304) );
  OAI21_X1 U13789 ( .B1(n13369), .B2(n11305), .A(n11304), .ZN(P2_U3253) );
  XNOR2_X1 U13790 ( .A(n11306), .B(n11310), .ZN(n14641) );
  INV_X1 U13791 ( .A(n14641), .ZN(n11320) );
  INV_X1 U13792 ( .A(n11307), .ZN(n11308) );
  AOI211_X1 U13793 ( .C1(n11310), .C2(n11309), .A(n14533), .B(n11308), .ZN(
        n14639) );
  INV_X1 U13794 ( .A(n11311), .ZN(n14388) );
  AOI211_X1 U13795 ( .C1(n14636), .C2(n11312), .A(n10341), .B(n14388), .ZN(
        n11313) );
  AOI21_X1 U13796 ( .B1(n14617), .B2(n14288), .A(n11313), .ZN(n14638) );
  NOR2_X1 U13797 ( .A1(n13849), .A2(n11678), .ZN(n11316) );
  INV_X1 U13798 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n13769) );
  INV_X1 U13799 ( .A(n11680), .ZN(n11314) );
  OAI22_X1 U13800 ( .A1(n14006), .A2(n13769), .B1(n11314), .B2(n13962), .ZN(
        n11315) );
  AOI211_X1 U13801 ( .C1(n14636), .C2(n14382), .A(n11316), .B(n11315), .ZN(
        n11317) );
  OAI21_X1 U13802 ( .B1(n14638), .B2(n13902), .A(n11317), .ZN(n11318) );
  AOI21_X1 U13803 ( .B1(n14639), .B2(n14006), .A(n11318), .ZN(n11319) );
  OAI21_X1 U13804 ( .B1(n11320), .B2(n14009), .A(n11319), .ZN(P1_U3283) );
  NAND2_X1 U13805 ( .A1(n11338), .A2(n12320), .ZN(n11326) );
  OR2_X1 U13806 ( .A1(n11607), .A2(n10612), .ZN(n11325) );
  NAND2_X1 U13807 ( .A1(n11326), .A2(n11325), .ZN(n11328) );
  XNOR2_X1 U13808 ( .A(n11328), .B(n11177), .ZN(n11331) );
  NOR2_X1 U13809 ( .A1(n11607), .A2(n10954), .ZN(n11329) );
  AOI21_X1 U13810 ( .B1(n11338), .B2(n12322), .A(n11329), .ZN(n11330) );
  NAND2_X1 U13811 ( .A1(n11331), .A2(n11330), .ZN(n11603) );
  OAI21_X1 U13812 ( .B1(n11331), .B2(n11330), .A(n11603), .ZN(n11332) );
  AOI21_X1 U13813 ( .B1(n11333), .B2(n11332), .A(n6755), .ZN(n11341) );
  OAI22_X1 U13814 ( .A1(n11678), .A2(n13647), .B1(n13646), .B2(n11334), .ZN(
        n11335) );
  AOI211_X1 U13815 ( .C1(n13654), .C2(n11337), .A(n11336), .B(n11335), .ZN(
        n11340) );
  NAND2_X1 U13816 ( .A1(n11338), .A2(n13658), .ZN(n11339) );
  OAI211_X1 U13817 ( .C1(n11341), .C2(n13660), .A(n11340), .B(n11339), .ZN(
        P1_U3221) );
  XOR2_X1 U13818 ( .A(n11343), .B(n11342), .Z(n11349) );
  INV_X1 U13819 ( .A(n15020), .ZN(n11346) );
  NOR2_X1 U13820 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11344), .ZN(n14882) );
  OAI22_X1 U13821 ( .A1(n12465), .A2(n15017), .B1(n15018), .B2(n12490), .ZN(
        n11345) );
  AOI211_X1 U13822 ( .C1(n11346), .C2(n12467), .A(n14882), .B(n11345), .ZN(
        n11348) );
  NAND2_X1 U13823 ( .A1(n12493), .A2(n15021), .ZN(n11347) );
  OAI211_X1 U13824 ( .C1(n11349), .C2(n12495), .A(n11348), .B(n11347), .ZN(
        P3_U3167) );
  NAND2_X1 U13825 ( .A1(n11350), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11352) );
  NAND2_X1 U13826 ( .A1(n11352), .A2(n11351), .ZN(n11353) );
  NOR2_X1 U13827 ( .A1(n11364), .A2(n11353), .ZN(n11354) );
  XOR2_X1 U13828 ( .A(n14480), .B(n11353), .Z(n14475) );
  NOR2_X1 U13829 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14475), .ZN(n14474) );
  NOR2_X1 U13830 ( .A1(n11354), .A2(n14474), .ZN(n11358) );
  NAND2_X1 U13831 ( .A1(n11360), .A2(n11623), .ZN(n11355) );
  OAI21_X1 U13832 ( .B1(n11360), .B2(n11623), .A(n11355), .ZN(n11357) );
  NAND2_X1 U13833 ( .A1(n11630), .A2(n11623), .ZN(n11356) );
  OAI211_X1 U13834 ( .C1(n11630), .C2(n11623), .A(n11358), .B(n11356), .ZN(
        n11622) );
  OAI211_X1 U13835 ( .C1(n11358), .C2(n11357), .A(n11622), .B(n14489), .ZN(
        n11372) );
  NAND2_X1 U13836 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13583)
         );
  NAND2_X1 U13837 ( .A1(n11360), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11359) );
  OAI21_X1 U13838 ( .B1(n11360), .B2(P1_REG1_REG_16__SCAN_IN), .A(n11359), 
        .ZN(n11361) );
  INV_X1 U13839 ( .A(n11361), .ZN(n11368) );
  AOI21_X1 U13840 ( .B1(n11363), .B2(n14420), .A(n11362), .ZN(n11365) );
  NOR2_X1 U13841 ( .A1(n11364), .A2(n11365), .ZN(n11366) );
  XOR2_X1 U13842 ( .A(n14480), .B(n11365), .Z(n14473) );
  NOR2_X1 U13843 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14473), .ZN(n14472) );
  NOR2_X1 U13844 ( .A1(n11366), .A2(n14472), .ZN(n11367) );
  NAND2_X1 U13845 ( .A1(n11367), .A2(n11368), .ZN(n11629) );
  OAI211_X1 U13846 ( .C1(n11368), .C2(n11367), .A(n14486), .B(n11629), .ZN(
        n11369) );
  NAND2_X1 U13847 ( .A1(n13583), .A2(n11369), .ZN(n11370) );
  AOI21_X1 U13848 ( .B1(n14468), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11370), 
        .ZN(n11371) );
  OAI211_X1 U13849 ( .C1(n14494), .C2(n11630), .A(n11372), .B(n11371), .ZN(
        P1_U3259) );
  INV_X1 U13850 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11384) );
  INV_X1 U13851 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11457) );
  NAND2_X1 U13852 ( .A1(n7599), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n11373) );
  NAND2_X1 U13853 ( .A1(n11375), .A2(n14849), .ZN(n11376) );
  INV_X1 U13854 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n15036) );
  INV_X1 U13855 ( .A(n14862), .ZN(n11377) );
  MUX2_X1 U13856 ( .A(n11457), .B(P3_REG2_REG_4__SCAN_IN), .S(n11430), .Z(
        n14861) );
  XNOR2_X1 U13857 ( .A(n11378), .B(n11431), .ZN(n14881) );
  INV_X1 U13858 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15023) );
  NOR2_X1 U13859 ( .A1(n14881), .A2(n15023), .ZN(n14880) );
  AOI21_X1 U13860 ( .B1(n11431), .B2(n11378), .A(n14880), .ZN(n14901) );
  INV_X1 U13861 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n15009) );
  AOI22_X1 U13862 ( .A1(n14914), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n15009), 
        .B2(n11424), .ZN(n14900) );
  NOR2_X1 U13863 ( .A1(n14901), .A2(n14900), .ZN(n14899) );
  NOR2_X1 U13864 ( .A1(n11401), .A2(n11379), .ZN(n11380) );
  INV_X1 U13865 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n14921) );
  INV_X1 U13866 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11716) );
  MUX2_X1 U13867 ( .A(n11716), .B(P3_REG2_REG_8__SCAN_IN), .S(n14942), .Z(
        n14940) );
  NOR2_X1 U13868 ( .A1(n11410), .A2(n11381), .ZN(n11382) );
  INV_X1 U13869 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n14956) );
  XNOR2_X1 U13870 ( .A(n11410), .B(n11381), .ZN(n14955) );
  NOR2_X1 U13871 ( .A1(n14956), .A2(n14955), .ZN(n14954) );
  INV_X1 U13872 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11821) );
  MUX2_X1 U13873 ( .A(P3_REG2_REG_10__SCAN_IN), .B(n11821), .S(n11441), .Z(
        n14973) );
  AOI21_X1 U13874 ( .B1(n11384), .B2(n11383), .A(n11515), .ZN(n11448) );
  MUX2_X1 U13875 ( .A(n15036), .B(n14850), .S(n11415), .Z(n11385) );
  NAND2_X1 U13876 ( .A1(n11385), .A2(n14849), .ZN(n11388) );
  INV_X1 U13877 ( .A(n11385), .ZN(n11386) );
  NAND2_X1 U13878 ( .A1(n11386), .A2(n11426), .ZN(n11387) );
  NAND2_X1 U13879 ( .A1(n11388), .A2(n11387), .ZN(n14842) );
  AOI21_X1 U13880 ( .B1(n14844), .B2(n14843), .A(n14842), .ZN(n14858) );
  INV_X1 U13881 ( .A(n11388), .ZN(n14857) );
  MUX2_X1 U13882 ( .A(n11457), .B(n11429), .S(n11415), .Z(n11389) );
  NAND2_X1 U13883 ( .A1(n11389), .A2(n11430), .ZN(n14886) );
  INV_X1 U13884 ( .A(n11389), .ZN(n11390) );
  NAND2_X1 U13885 ( .A1(n11390), .A2(n14875), .ZN(n11391) );
  AND2_X1 U13886 ( .A1(n14886), .A2(n11391), .ZN(n14856) );
  OAI21_X1 U13887 ( .B1(n14858), .B2(n14857), .A(n14856), .ZN(n14887) );
  MUX2_X1 U13888 ( .A(n15023), .B(n14893), .S(n11415), .Z(n11392) );
  NAND2_X1 U13889 ( .A1(n11392), .A2(n14892), .ZN(n11395) );
  INV_X1 U13890 ( .A(n11392), .ZN(n11393) );
  NAND2_X1 U13891 ( .A1(n11393), .A2(n11431), .ZN(n11394) );
  NAND2_X1 U13892 ( .A1(n11395), .A2(n11394), .ZN(n14885) );
  INV_X1 U13893 ( .A(n11395), .ZN(n14909) );
  MUX2_X1 U13894 ( .A(n15009), .B(n11396), .S(n11415), .Z(n11397) );
  NAND2_X1 U13895 ( .A1(n11397), .A2(n14914), .ZN(n14923) );
  INV_X1 U13896 ( .A(n11397), .ZN(n11398) );
  NAND2_X1 U13897 ( .A1(n11398), .A2(n11424), .ZN(n11399) );
  AND2_X1 U13898 ( .A1(n14923), .A2(n11399), .ZN(n14908) );
  OAI21_X1 U13899 ( .B1(n14910), .B2(n14909), .A(n14908), .ZN(n14924) );
  MUX2_X1 U13900 ( .A(n14921), .B(n11400), .S(n11415), .Z(n11402) );
  NAND2_X1 U13901 ( .A1(n11402), .A2(n11401), .ZN(n11405) );
  INV_X1 U13902 ( .A(n11402), .ZN(n11403) );
  NAND2_X1 U13903 ( .A1(n11403), .A2(n14927), .ZN(n11404) );
  NAND2_X1 U13904 ( .A1(n11405), .A2(n11404), .ZN(n14922) );
  AOI21_X1 U13905 ( .B1(n14924), .B2(n14923), .A(n14922), .ZN(n14945) );
  INV_X1 U13906 ( .A(n11405), .ZN(n14944) );
  MUX2_X1 U13907 ( .A(n11716), .B(n11436), .S(n11415), .Z(n11406) );
  INV_X1 U13908 ( .A(n14942), .ZN(n11437) );
  NAND2_X1 U13909 ( .A1(n11406), .A2(n11437), .ZN(n14958) );
  INV_X1 U13910 ( .A(n11406), .ZN(n11407) );
  NAND2_X1 U13911 ( .A1(n11407), .A2(n14942), .ZN(n11408) );
  AND2_X1 U13912 ( .A1(n14958), .A2(n11408), .ZN(n14943) );
  OAI21_X1 U13913 ( .B1(n14945), .B2(n14944), .A(n14943), .ZN(n14959) );
  MUX2_X1 U13914 ( .A(n14956), .B(n11409), .S(n11415), .Z(n11411) );
  NAND2_X1 U13915 ( .A1(n11411), .A2(n11410), .ZN(n11414) );
  INV_X1 U13916 ( .A(n11411), .ZN(n11412) );
  NAND2_X1 U13917 ( .A1(n11412), .A2(n14963), .ZN(n11413) );
  NAND2_X1 U13918 ( .A1(n11414), .A2(n11413), .ZN(n14957) );
  INV_X1 U13919 ( .A(n11414), .ZN(n14984) );
  MUX2_X1 U13920 ( .A(n11821), .B(n11440), .S(n11415), .Z(n11416) );
  NAND2_X1 U13921 ( .A1(n11416), .A2(n11441), .ZN(n11419) );
  INV_X1 U13922 ( .A(n11416), .ZN(n11417) );
  NAND2_X1 U13923 ( .A1(n11417), .A2(n14981), .ZN(n11418) );
  AND2_X1 U13924 ( .A1(n11419), .A2(n11418), .ZN(n14983) );
  OAI21_X1 U13925 ( .B1(n14985), .B2(n14984), .A(n14983), .ZN(n14988) );
  NAND2_X1 U13926 ( .A1(n14988), .A2(n11419), .ZN(n11422) );
  MUX2_X1 U13927 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n11415), .Z(n11520) );
  XNOR2_X1 U13928 ( .A(n11520), .B(n11521), .ZN(n11421) );
  NAND2_X1 U13929 ( .A1(n11422), .A2(n11421), .ZN(n11524) );
  OAI21_X1 U13930 ( .B1(n11422), .B2(n11421), .A(n11524), .ZN(n11423) );
  NAND2_X1 U13931 ( .A1(n11423), .A2(n14960), .ZN(n11447) );
  AOI22_X1 U13932 ( .A1(n14914), .A2(n11396), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n11424), .ZN(n14903) );
  XNOR2_X1 U13933 ( .A(n11427), .B(n11426), .ZN(n14851) );
  OAI22_X1 U13934 ( .A1(n11428), .A2(n14849), .B1(n14850), .B2(n14851), .ZN(
        n14868) );
  MUX2_X1 U13935 ( .A(n11429), .B(P3_REG1_REG_4__SCAN_IN), .S(n11430), .Z(
        n14869) );
  NAND2_X1 U13936 ( .A1(n14868), .A2(n14869), .ZN(n14867) );
  OAI21_X1 U13937 ( .B1(n11430), .B2(n11429), .A(n14867), .ZN(n11432) );
  XNOR2_X1 U13938 ( .A(n11432), .B(n11431), .ZN(n14894) );
  INV_X1 U13939 ( .A(n11432), .ZN(n11433) );
  OAI22_X1 U13940 ( .A1(n14894), .A2(n14893), .B1(n14892), .B2(n11433), .ZN(
        n14904) );
  NAND2_X1 U13941 ( .A1(n14903), .A2(n14904), .ZN(n14902) );
  NAND2_X1 U13942 ( .A1(n14927), .A2(n11434), .ZN(n11435) );
  MUX2_X1 U13943 ( .A(P3_REG1_REG_8__SCAN_IN), .B(n11436), .S(n14942), .Z(
        n14937) );
  NAND2_X1 U13944 ( .A1(n14938), .A2(n14937), .ZN(n14936) );
  NAND2_X1 U13945 ( .A1(n14963), .A2(n11438), .ZN(n11439) );
  MUX2_X1 U13946 ( .A(n11440), .B(P3_REG1_REG_10__SCAN_IN), .S(n11441), .Z(
        n14976) );
  NAND2_X1 U13947 ( .A1(n14977), .A2(n14976), .ZN(n14975) );
  OAI21_X1 U13948 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n11442), .A(n11529), 
        .ZN(n11445) );
  INV_X1 U13949 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n15211) );
  NOR2_X1 U13950 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15211), .ZN(n12454) );
  AOI21_X1 U13951 ( .B1(n14978), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n12454), 
        .ZN(n11443) );
  OAI21_X1 U13952 ( .B1(n14982), .B2(n11528), .A(n11443), .ZN(n11444) );
  AOI21_X1 U13953 ( .B1(n11445), .B2(n14992), .A(n11444), .ZN(n11446) );
  OAI211_X1 U13954 ( .C1(n11448), .C2(n14994), .A(n11447), .B(n11446), .ZN(
        P3_U3193) );
  XNOR2_X1 U13955 ( .A(n11450), .B(n11449), .ZN(n15089) );
  INV_X1 U13956 ( .A(n15089), .ZN(n11462) );
  AND2_X1 U13957 ( .A1(n15058), .A2(n11451), .ZN(n15049) );
  AND2_X1 U13958 ( .A1(n15074), .A2(n15049), .ZN(n15072) );
  INV_X1 U13959 ( .A(n15072), .ZN(n11721) );
  XNOR2_X1 U13960 ( .A(n11453), .B(n11452), .ZN(n11455) );
  AOI22_X1 U13961 ( .A1(n15062), .A2(n12504), .B1(n15002), .B2(n15059), .ZN(
        n11454) );
  OAI21_X1 U13962 ( .B1(n11455), .B2(n15016), .A(n11454), .ZN(n11456) );
  AOI21_X1 U13963 ( .B1(n15089), .B2(n14997), .A(n11456), .ZN(n15086) );
  MUX2_X1 U13964 ( .A(n11457), .B(n15086), .S(n15074), .Z(n11461) );
  NOR2_X1 U13965 ( .A1(n11458), .A2(n15103), .ZN(n15088) );
  AOI22_X1 U13966 ( .A1(n15034), .A2(n15088), .B1(n15071), .B2(n11459), .ZN(
        n11460) );
  OAI211_X1 U13967 ( .C1(n11462), .C2(n11721), .A(n11461), .B(n11460), .ZN(
        P3_U3229) );
  XNOR2_X1 U13968 ( .A(n11463), .B(n11465), .ZN(n14287) );
  OAI211_X1 U13969 ( .C1(n11466), .C2(n11465), .A(n11464), .B(n14376), .ZN(
        n14294) );
  INV_X1 U13970 ( .A(n14294), .ZN(n11473) );
  OAI211_X1 U13971 ( .C1(n11467), .C2(n14386), .A(n14559), .B(n14309), .ZN(
        n14292) );
  OR2_X1 U13972 ( .A1(n13966), .A2(n14411), .ZN(n11469) );
  AOI22_X1 U13973 ( .A1(n14539), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n11789), 
        .B2(n14538), .ZN(n11468) );
  OAI211_X1 U13974 ( .C1(n11792), .C2(n13849), .A(n11469), .B(n11468), .ZN(
        n11470) );
  AOI21_X1 U13975 ( .B1(n14290), .B2(n14382), .A(n11470), .ZN(n11471) );
  OAI21_X1 U13976 ( .B1(n14292), .B2(n13902), .A(n11471), .ZN(n11472) );
  AOI21_X1 U13977 ( .B1(n11473), .B2(n14006), .A(n11472), .ZN(n11474) );
  OAI21_X1 U13978 ( .B1(n14009), .B2(n14287), .A(n11474), .ZN(P1_U3281) );
  AOI211_X1 U13979 ( .C1(n14792), .C2(n12031), .A(n11476), .B(n11475), .ZN(
        n11477) );
  OAI21_X1 U13980 ( .B1(n13456), .B2(n11478), .A(n11477), .ZN(n11481) );
  NAND2_X1 U13981 ( .A1(n11481), .A2(n14837), .ZN(n11479) );
  OAI21_X1 U13982 ( .B1(n13457), .B2(n11480), .A(n11479), .ZN(P2_U3510) );
  INV_X1 U13983 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11483) );
  NAND2_X1 U13984 ( .A1(n11481), .A2(n6621), .ZN(n11482) );
  OAI21_X1 U13985 ( .B1(n6621), .B2(n11483), .A(n11482), .ZN(P2_U3463) );
  OAI211_X1 U13986 ( .C1(n11486), .C2(n14826), .A(n11485), .B(n11484), .ZN(
        n11487) );
  AOI21_X1 U13987 ( .B1(n11488), .B2(n14808), .A(n11487), .ZN(n11491) );
  NAND2_X1 U13988 ( .A1(n14835), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n11489) );
  OAI21_X1 U13989 ( .B1(n11491), .B2(n14835), .A(n11489), .ZN(P2_U3511) );
  NAND2_X1 U13990 ( .A1(n14829), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n11490) );
  OAI21_X1 U13991 ( .B1(n11491), .B2(n14829), .A(n11490), .ZN(P2_U3466) );
  INV_X1 U13992 ( .A(n15007), .ZN(n11500) );
  OAI211_X1 U13993 ( .C1(n11494), .C2(n11493), .A(n11492), .B(n12473), .ZN(
        n11499) );
  NAND2_X1 U13994 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n14916) );
  INV_X1 U13995 ( .A(n14916), .ZN(n11497) );
  OAI22_X1 U13996 ( .A1(n12485), .A2(n15006), .B1(n12465), .B2(n11495), .ZN(
        n11496) );
  AOI211_X1 U13997 ( .C1(n12462), .C2(n15001), .A(n11497), .B(n11496), .ZN(
        n11498) );
  OAI211_X1 U13998 ( .C1(n11500), .C2(n11768), .A(n11499), .B(n11498), .ZN(
        P3_U3179) );
  XOR2_X1 U13999 ( .A(n12180), .B(n11501), .Z(n11618) );
  INV_X1 U14000 ( .A(n11618), .ZN(n11513) );
  OAI211_X1 U14001 ( .C1(n11503), .C2(n12180), .A(n11502), .B(n13350), .ZN(
        n11505) );
  NAND2_X1 U14002 ( .A1(n11505), .A2(n11504), .ZN(n11616) );
  AOI21_X1 U14003 ( .B1(n11506), .B2(n12044), .A(n13336), .ZN(n11507) );
  NAND2_X1 U14004 ( .A1(n11507), .A2(n11641), .ZN(n11614) );
  AOI22_X1 U14005 ( .A1(n14761), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11508), 
        .B2(n14759), .ZN(n11510) );
  NAND2_X1 U14006 ( .A1(n12044), .A2(n13366), .ZN(n11509) );
  OAI211_X1 U14007 ( .C1(n11614), .C2(n13363), .A(n11510), .B(n11509), .ZN(
        n11511) );
  AOI21_X1 U14008 ( .B1(n11616), .B2(n13357), .A(n11511), .ZN(n11512) );
  OAI21_X1 U14009 ( .B1(n13369), .B2(n11513), .A(n11512), .ZN(P2_U3252) );
  NOR2_X1 U14010 ( .A1(n11521), .A2(n11514), .ZN(n11516) );
  INV_X1 U14011 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11517) );
  AOI22_X1 U14012 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n11594), .B1(n11586), 
        .B2(n11517), .ZN(n11518) );
  AOI21_X1 U14013 ( .B1(n11519), .B2(n11518), .A(n11584), .ZN(n11539) );
  INV_X1 U14014 ( .A(n11520), .ZN(n11522) );
  NAND2_X1 U14015 ( .A1(n11522), .A2(n11521), .ZN(n11523) );
  AND2_X1 U14016 ( .A1(n11524), .A2(n11523), .ZN(n11526) );
  MUX2_X1 U14017 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n11415), .Z(n11587) );
  XNOR2_X1 U14018 ( .A(n11587), .B(n11594), .ZN(n11525) );
  NAND3_X1 U14019 ( .A1(n11524), .A2(n11523), .A3(n11525), .ZN(n11590) );
  OAI211_X1 U14020 ( .C1(n11526), .C2(n11525), .A(n14960), .B(n11590), .ZN(
        n11538) );
  AOI22_X1 U14021 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n11586), .B1(n11594), 
        .B2(n7769), .ZN(n11532) );
  NAND2_X1 U14022 ( .A1(n11528), .A2(n11527), .ZN(n11530) );
  NAND2_X1 U14023 ( .A1(n11532), .A2(n11531), .ZN(n11593) );
  OAI21_X1 U14024 ( .B1(n11532), .B2(n11531), .A(n11593), .ZN(n11536) );
  INV_X1 U14025 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11533) );
  NOR2_X1 U14026 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11533), .ZN(n12392) );
  AOI21_X1 U14027 ( .B1(n14978), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12392), 
        .ZN(n11534) );
  OAI21_X1 U14028 ( .B1(n14982), .B2(n11586), .A(n11534), .ZN(n11535) );
  AOI21_X1 U14029 ( .B1(n11536), .B2(n14992), .A(n11535), .ZN(n11537) );
  OAI211_X1 U14030 ( .C1(n11539), .C2(n14994), .A(n11538), .B(n11537), .ZN(
        P3_U3194) );
  NAND2_X1 U14031 ( .A1(n14749), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11549) );
  INV_X1 U14032 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11540) );
  AOI22_X1 U14033 ( .A1(n14749), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n11540), 
        .B2(n11563), .ZN(n14744) );
  NAND2_X1 U14034 ( .A1(n14727), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11548) );
  INV_X1 U14035 ( .A(n11548), .ZN(n11541) );
  AOI21_X1 U14036 ( .B1(n13356), .B2(n11562), .A(n11541), .ZN(n14730) );
  INV_X1 U14037 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11543) );
  OAI21_X1 U14038 ( .B1(n11552), .B2(P2_REG2_REG_12__SCAN_IN), .A(n11542), 
        .ZN(n14693) );
  MUX2_X1 U14039 ( .A(n11543), .B(P2_REG2_REG_13__SCAN_IN), .S(n11553), .Z(
        n14692) );
  OAI21_X1 U14040 ( .B1(n11543), .B2(n14689), .A(n14694), .ZN(n11544) );
  NAND2_X1 U14041 ( .A1(n11554), .A2(n11544), .ZN(n11545) );
  XNOR2_X1 U14042 ( .A(n11544), .B(n14706), .ZN(n14710) );
  NAND2_X1 U14043 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n14710), .ZN(n14709) );
  NAND2_X1 U14044 ( .A1(n11545), .A2(n14709), .ZN(n11546) );
  NAND2_X1 U14045 ( .A1(n11559), .A2(n11546), .ZN(n11547) );
  XOR2_X1 U14046 ( .A(n11559), .B(n11546), .Z(n14714) );
  NAND2_X1 U14047 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14714), .ZN(n14713) );
  NAND2_X1 U14048 ( .A1(n11547), .A2(n14713), .ZN(n14731) );
  NAND2_X1 U14049 ( .A1(n14730), .A2(n14731), .ZN(n14728) );
  NAND2_X1 U14050 ( .A1(n11548), .A2(n14728), .ZN(n14743) );
  NAND2_X1 U14051 ( .A1(n14744), .A2(n14743), .ZN(n14742) );
  NAND2_X1 U14052 ( .A1(n11549), .A2(n14742), .ZN(n13131) );
  XOR2_X1 U14053 ( .A(n11570), .B(n13131), .Z(n11550) );
  NOR2_X1 U14054 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n11550), .ZN(n13133) );
  AOI21_X1 U14055 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n11550), .A(n13133), 
        .ZN(n11573) );
  INV_X1 U14056 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11564) );
  XNOR2_X1 U14057 ( .A(n11563), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14754) );
  INV_X1 U14058 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n11561) );
  XNOR2_X1 U14059 ( .A(n11562), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14733) );
  INV_X1 U14060 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11556) );
  OAI21_X1 U14061 ( .B1(n11552), .B2(P2_REG1_REG_12__SCAN_IN), .A(n11551), 
        .ZN(n14697) );
  XNOR2_X1 U14062 ( .A(n11553), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n14698) );
  NOR2_X1 U14063 ( .A1(n14697), .A2(n14698), .ZN(n14696) );
  AOI21_X1 U14064 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n11553), .A(n14696), 
        .ZN(n14703) );
  XNOR2_X1 U14065 ( .A(n11554), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n14704) );
  OR2_X1 U14066 ( .A1(n14703), .A2(n14704), .ZN(n11555) );
  OAI21_X1 U14067 ( .B1(n11556), .B2(n14706), .A(n11555), .ZN(n11557) );
  NAND2_X1 U14068 ( .A1(n11559), .A2(n11557), .ZN(n11560) );
  INV_X1 U14069 ( .A(n11557), .ZN(n11558) );
  XNOR2_X1 U14070 ( .A(n11559), .B(n11558), .ZN(n14716) );
  NAND2_X1 U14071 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n14716), .ZN(n14715) );
  NAND2_X1 U14072 ( .A1(n11560), .A2(n14715), .ZN(n14734) );
  NAND2_X1 U14073 ( .A1(n14733), .A2(n14734), .ZN(n14732) );
  OAI21_X1 U14074 ( .B1(n11562), .B2(n11561), .A(n14732), .ZN(n14753) );
  NAND2_X1 U14075 ( .A1(n14754), .A2(n14753), .ZN(n14751) );
  OAI21_X1 U14076 ( .B1(n11564), .B2(n11563), .A(n14751), .ZN(n13135) );
  INV_X1 U14077 ( .A(n13135), .ZN(n11565) );
  XNOR2_X1 U14078 ( .A(n13136), .B(n11565), .ZN(n11566) );
  NAND2_X1 U14079 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n11566), .ZN(n13138) );
  OAI21_X1 U14080 ( .B1(n11566), .B2(P2_REG1_REG_18__SCAN_IN), .A(n13138), 
        .ZN(n11567) );
  OR2_X1 U14081 ( .A1(n14718), .A2(n11567), .ZN(n11569) );
  AND2_X1 U14082 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13064) );
  AOI21_X1 U14083 ( .B1(n14726), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n13064), 
        .ZN(n11568) );
  OAI211_X1 U14084 ( .C1(n14722), .C2(n11570), .A(n11569), .B(n11568), .ZN(
        n11571) );
  INV_X1 U14085 ( .A(n11571), .ZN(n11572) );
  OAI21_X1 U14086 ( .B1(n11573), .B2(n14745), .A(n11572), .ZN(P2_U3232) );
  OAI222_X1 U14087 ( .A1(n13498), .A2(n15235), .B1(P2_U3088), .B2(n12131), 
        .C1(n13505), .C2(n11574), .ZN(P2_U3305) );
  INV_X1 U14088 ( .A(n11576), .ZN(n11577) );
  AOI21_X1 U14089 ( .B1(n11578), .B2(n11575), .A(n11577), .ZN(n11583) );
  NAND2_X1 U14090 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14705)
         );
  OAI22_X1 U14091 ( .A1(n12051), .A2(n13042), .B1(n11579), .B2(n13060), .ZN(
        n11638) );
  NAND2_X1 U14092 ( .A1(n13065), .A2(n11638), .ZN(n11580) );
  OAI211_X1 U14093 ( .C1(n13067), .C2(n11642), .A(n14705), .B(n11580), .ZN(
        n11581) );
  AOI21_X1 U14094 ( .B1(n13452), .B2(n13081), .A(n11581), .ZN(n11582) );
  OAI21_X1 U14095 ( .B1(n11583), .B2(n13083), .A(n11582), .ZN(P2_U3187) );
  INV_X1 U14096 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n15398) );
  AOI21_X1 U14097 ( .B1(n15398), .B2(n11585), .A(n11839), .ZN(n11601) );
  NAND2_X1 U14098 ( .A1(n11587), .A2(n11586), .ZN(n11589) );
  MUX2_X1 U14099 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n11415), .Z(n11851) );
  XNOR2_X1 U14100 ( .A(n11851), .B(n11852), .ZN(n11588) );
  NAND3_X1 U14101 ( .A1(n11590), .A2(n11589), .A3(n11588), .ZN(n11858) );
  INV_X1 U14102 ( .A(n11858), .ZN(n11592) );
  AOI21_X1 U14103 ( .B1(n11590), .B2(n11589), .A(n11588), .ZN(n11591) );
  OAI21_X1 U14104 ( .B1(n11592), .B2(n11591), .A(n14960), .ZN(n11600) );
  OAI21_X1 U14105 ( .B1(n11594), .B2(n7769), .A(n11593), .ZN(n11844) );
  XNOR2_X1 U14106 ( .A(n11844), .B(n11852), .ZN(n11595) );
  NAND2_X1 U14107 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n11595), .ZN(n11846) );
  OAI21_X1 U14108 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n11595), .A(n11846), 
        .ZN(n11598) );
  NOR2_X1 U14109 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7788), .ZN(n11920) );
  AOI21_X1 U14110 ( .B1(n14978), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n11920), 
        .ZN(n11596) );
  OAI21_X1 U14111 ( .B1(n14982), .B2(n11845), .A(n11596), .ZN(n11597) );
  AOI21_X1 U14112 ( .B1(n11598), .B2(n14992), .A(n11597), .ZN(n11599) );
  OAI211_X1 U14113 ( .C1(n11601), .C2(n14994), .A(n11600), .B(n11599), .ZN(
        P3_U3195) );
  OAI22_X1 U14114 ( .A1(n14627), .A2(n10612), .B1(n11678), .B2(n10954), .ZN(
        n11664) );
  OAI22_X1 U14115 ( .A1(n14627), .A2(n10348), .B1(n11678), .B2(n10612), .ZN(
        n11602) );
  XNOR2_X1 U14116 ( .A(n11602), .B(n12323), .ZN(n11663) );
  XOR2_X1 U14117 ( .A(n11664), .B(n11663), .Z(n11605) );
  OAI21_X1 U14118 ( .B1(n11605), .B2(n11604), .A(n11667), .ZN(n11606) );
  NAND2_X1 U14119 ( .A1(n11606), .A2(n13634), .ZN(n11613) );
  NAND2_X1 U14120 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n13752) );
  INV_X1 U14121 ( .A(n13752), .ZN(n11610) );
  OAI22_X1 U14122 ( .A1(n11608), .A2(n13647), .B1(n13646), .B2(n11607), .ZN(
        n11609) );
  AOI211_X1 U14123 ( .C1(n11611), .C2(n13654), .A(n11610), .B(n11609), .ZN(
        n11612) );
  OAI211_X1 U14124 ( .C1(n14627), .C2(n13640), .A(n11613), .B(n11612), .ZN(
        P1_U3231) );
  INV_X1 U14125 ( .A(n12044), .ZN(n11615) );
  OAI21_X1 U14126 ( .B1(n11615), .B2(n14826), .A(n11614), .ZN(n11617) );
  AOI211_X1 U14127 ( .C1(n11618), .C2(n14808), .A(n11617), .B(n11616), .ZN(
        n11621) );
  NAND2_X1 U14128 ( .A1(n14829), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n11619) );
  OAI21_X1 U14129 ( .B1(n11621), .B2(n14829), .A(n11619), .ZN(P2_U3469) );
  NAND2_X1 U14130 ( .A1(n14835), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11620) );
  OAI21_X1 U14131 ( .B1(n11621), .B2(n14835), .A(n11620), .ZN(P2_U3512) );
  OAI21_X1 U14132 ( .B1(n11630), .B2(n11623), .A(n11622), .ZN(n11627) );
  INV_X1 U14133 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11625) );
  NAND2_X1 U14134 ( .A1(n13778), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n13786) );
  INV_X1 U14135 ( .A(n13786), .ZN(n11624) );
  AOI21_X1 U14136 ( .B1(n11625), .B2(n11636), .A(n11624), .ZN(n11626) );
  NAND2_X1 U14137 ( .A1(n11626), .A2(n11627), .ZN(n13785) );
  OAI211_X1 U14138 ( .C1(n11627), .C2(n11626), .A(n14489), .B(n13785), .ZN(
        n11635) );
  NAND2_X1 U14139 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13597)
         );
  INV_X1 U14140 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n11628) );
  XNOR2_X1 U14141 ( .A(n13778), .B(n11628), .ZN(n13779) );
  OAI21_X1 U14142 ( .B1(n9553), .B2(n11630), .A(n11629), .ZN(n13780) );
  XOR2_X1 U14143 ( .A(n13779), .B(n13780), .Z(n11631) );
  NAND2_X1 U14144 ( .A1(n14486), .A2(n11631), .ZN(n11632) );
  NAND2_X1 U14145 ( .A1(n13597), .A2(n11632), .ZN(n11633) );
  AOI21_X1 U14146 ( .B1(n14468), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n11633), 
        .ZN(n11634) );
  OAI211_X1 U14147 ( .C1(n14494), .C2(n11636), .A(n11635), .B(n11634), .ZN(
        P1_U3260) );
  XNOR2_X1 U14148 ( .A(n13452), .B(n13100), .ZN(n12182) );
  XOR2_X1 U14149 ( .A(n11637), .B(n12182), .Z(n11639) );
  AOI21_X1 U14150 ( .B1(n11639), .B2(n13350), .A(n11638), .ZN(n13454) );
  AOI211_X1 U14151 ( .C1(n13452), .C2(n11641), .A(n13336), .B(n11640), .ZN(
        n13451) );
  INV_X1 U14152 ( .A(n13452), .ZN(n12049) );
  INV_X1 U14153 ( .A(n11642), .ZN(n11643) );
  AOI22_X1 U14154 ( .A1(n14761), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11643), 
        .B2(n14759), .ZN(n11644) );
  OAI21_X1 U14155 ( .B1(n12049), .B2(n14764), .A(n11644), .ZN(n11647) );
  XOR2_X1 U14156 ( .A(n12182), .B(n11645), .Z(n13455) );
  NOR2_X1 U14157 ( .A1(n13455), .A2(n13369), .ZN(n11646) );
  AOI211_X1 U14158 ( .C1(n13451), .C2(n14757), .A(n11647), .B(n11646), .ZN(
        n11648) );
  OAI21_X1 U14159 ( .B1(n14770), .B2(n13454), .A(n11648), .ZN(P2_U3251) );
  OAI211_X1 U14160 ( .C1(n11650), .C2(n7262), .A(n11649), .B(n14376), .ZN(
        n14418) );
  INV_X1 U14161 ( .A(n11651), .ZN(n14372) );
  AOI211_X1 U14162 ( .C1(n14414), .C2(n14311), .A(n10341), .B(n14372), .ZN(
        n14412) );
  AOI22_X1 U14163 ( .A1(n14539), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n13523), 
        .B2(n14538), .ZN(n11652) );
  OAI21_X1 U14164 ( .B1(n13966), .B2(n14409), .A(n11652), .ZN(n11653) );
  AOI21_X1 U14165 ( .B1(n13960), .B2(n14289), .A(n11653), .ZN(n11654) );
  OAI21_X1 U14166 ( .B1(n9532), .B2(n14541), .A(n11654), .ZN(n11655) );
  AOI21_X1 U14167 ( .B1(n14412), .B2(n14548), .A(n11655), .ZN(n11658) );
  NAND2_X1 U14168 ( .A1(n11656), .A2(n7262), .ZN(n14415) );
  NAND3_X1 U14169 ( .A1(n14416), .A2(n14415), .A3(n14390), .ZN(n11657) );
  OAI211_X1 U14170 ( .C1(n14418), .C2(n14552), .A(n11658), .B(n11657), .ZN(
        P1_U3279) );
  INV_X1 U14171 ( .A(n11659), .ZN(n11660) );
  OAI222_X1 U14172 ( .A1(P3_U3151), .A2(n11662), .B1(n12944), .B2(n11661), 
        .C1(n11943), .C2(n11660), .ZN(P3_U3271) );
  INV_X1 U14173 ( .A(n14636), .ZN(n11683) );
  INV_X1 U14174 ( .A(n11663), .ZN(n11666) );
  INV_X1 U14175 ( .A(n11664), .ZN(n11665) );
  NAND2_X1 U14176 ( .A1(n11666), .A2(n11665), .ZN(n11672) );
  AND2_X1 U14177 ( .A1(n11667), .A2(n11672), .ZN(n11676) );
  NAND2_X1 U14178 ( .A1(n14636), .A2(n12320), .ZN(n11669) );
  NAND2_X1 U14179 ( .A1(n13668), .A2(n12322), .ZN(n11668) );
  NAND2_X1 U14180 ( .A1(n11669), .A2(n11668), .ZN(n11670) );
  XNOR2_X1 U14181 ( .A(n11670), .B(n12323), .ZN(n11747) );
  AND2_X1 U14182 ( .A1(n12321), .A2(n13668), .ZN(n11671) );
  AOI21_X1 U14183 ( .B1(n14636), .B2(n12322), .A(n11671), .ZN(n11745) );
  XNOR2_X1 U14184 ( .A(n11747), .B(n11745), .ZN(n11675) );
  AND2_X1 U14185 ( .A1(n11675), .A2(n11672), .ZN(n11673) );
  OAI211_X1 U14186 ( .C1(n11676), .C2(n11675), .A(n13634), .B(n11753), .ZN(
        n11682) );
  NOR2_X1 U14187 ( .A1(n11677), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13767) );
  OAI22_X1 U14188 ( .A1(n11792), .A2(n13647), .B1(n13646), .B2(n11678), .ZN(
        n11679) );
  AOI211_X1 U14189 ( .C1(n13654), .C2(n11680), .A(n13767), .B(n11679), .ZN(
        n11681) );
  OAI211_X1 U14190 ( .C1(n11683), .C2(n13640), .A(n11682), .B(n11681), .ZN(
        P1_U3217) );
  INV_X1 U14191 ( .A(n11831), .ZN(n11690) );
  OAI211_X1 U14192 ( .C1(n11686), .C2(n11685), .A(n11684), .B(n12473), .ZN(
        n11689) );
  AND2_X1 U14193 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n14929) );
  OAI22_X1 U14194 ( .A1(n12465), .A2(n15018), .B1(n11886), .B2(n12490), .ZN(
        n11687) );
  AOI211_X1 U14195 ( .C1(n11835), .C2(n12467), .A(n14929), .B(n11687), .ZN(
        n11688) );
  OAI211_X1 U14196 ( .C1(n11690), .C2(n11768), .A(n11689), .B(n11688), .ZN(
        P3_U3153) );
  XNOR2_X1 U14197 ( .A(n11691), .B(n12184), .ZN(n13446) );
  XNOR2_X1 U14198 ( .A(n11693), .B(n11692), .ZN(n11694) );
  NAND2_X1 U14199 ( .A1(n11694), .A2(n13350), .ZN(n11696) );
  AND2_X1 U14200 ( .A1(n13100), .A2(n13075), .ZN(n11695) );
  AOI21_X1 U14201 ( .B1(n13098), .B2(n13076), .A(n11695), .ZN(n11802) );
  NAND2_X1 U14202 ( .A1(n11696), .A2(n11802), .ZN(n13450) );
  NAND2_X1 U14203 ( .A1(n13450), .A2(n13357), .ZN(n11703) );
  INV_X1 U14204 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n11697) );
  OAI22_X1 U14205 ( .A1(n13357), .A2(n11697), .B1(n11801), .B2(n13354), .ZN(
        n11701) );
  AOI21_X1 U14206 ( .B1(n12052), .B2(n11698), .A(n13336), .ZN(n11699) );
  NAND2_X1 U14207 ( .A1(n11699), .A2(n13358), .ZN(n13447) );
  NOR2_X1 U14208 ( .A1(n13447), .A2(n13363), .ZN(n11700) );
  AOI211_X1 U14209 ( .C1(n13366), .C2(n12052), .A(n11701), .B(n11700), .ZN(
        n11702) );
  OAI211_X1 U14210 ( .C1(n13369), .C2(n13446), .A(n11703), .B(n11702), .ZN(
        P2_U3250) );
  NAND2_X1 U14211 ( .A1(n11704), .A2(n11834), .ZN(n11833) );
  NAND2_X1 U14212 ( .A1(n11833), .A2(n11705), .ZN(n11709) );
  NAND2_X1 U14213 ( .A1(n11704), .A2(n11706), .ZN(n11724) );
  AND2_X1 U14214 ( .A1(n11724), .A2(n11707), .ZN(n11708) );
  OAI21_X1 U14215 ( .B1(n11709), .B2(n7014), .A(n11708), .ZN(n15107) );
  INV_X1 U14216 ( .A(n15107), .ZN(n11722) );
  XNOR2_X1 U14217 ( .A(n11711), .B(n11710), .ZN(n11714) );
  NAND2_X1 U14218 ( .A1(n15107), .A2(n14997), .ZN(n11713) );
  AOI22_X1 U14219 ( .A1(n15059), .A2(n12360), .B1(n15001), .B2(n15062), .ZN(
        n11712) );
  OAI211_X1 U14220 ( .C1(n15016), .C2(n11714), .A(n11713), .B(n11712), .ZN(
        n15105) );
  NAND2_X1 U14221 ( .A1(n15105), .A2(n15074), .ZN(n11720) );
  INV_X1 U14222 ( .A(n11715), .ZN(n11769) );
  OAI22_X1 U14223 ( .A1(n15074), .A2(n11716), .B1(n11769), .B2(n12766), .ZN(
        n11717) );
  AOI21_X1 U14224 ( .B1(n12770), .B2(n11718), .A(n11717), .ZN(n11719) );
  OAI211_X1 U14225 ( .C1(n11722), .C2(n11721), .A(n11720), .B(n11719), .ZN(
        P3_U3225) );
  NAND2_X1 U14226 ( .A1(n11724), .A2(n11723), .ZN(n11725) );
  XNOR2_X1 U14227 ( .A(n11725), .B(n11727), .ZN(n15110) );
  NAND2_X1 U14228 ( .A1(n11728), .A2(n11727), .ZN(n11729) );
  NAND3_X1 U14229 ( .A1(n11726), .A2(n8938), .A3(n11729), .ZN(n11732) );
  AOI22_X1 U14230 ( .A1(n15062), .A2(n11730), .B1(n12502), .B2(n15059), .ZN(
        n11731) );
  NAND2_X1 U14231 ( .A1(n11732), .A2(n11731), .ZN(n11733) );
  AOI21_X1 U14232 ( .B1(n15110), .B2(n14997), .A(n11733), .ZN(n15112) );
  AND2_X1 U14233 ( .A1(n11888), .A2(n14345), .ZN(n15109) );
  AOI22_X1 U14234 ( .A1(n15034), .A2(n15109), .B1(n15071), .B2(n11889), .ZN(
        n11734) );
  OAI21_X1 U14235 ( .B1(n14956), .B2(n15074), .A(n11734), .ZN(n11735) );
  AOI21_X1 U14236 ( .B1(n15110), .B2(n15072), .A(n11735), .ZN(n11736) );
  OAI21_X1 U14237 ( .B1(n15112), .B2(n15056), .A(n11736), .ZN(P3_U3224) );
  INV_X1 U14238 ( .A(n11737), .ZN(n11739) );
  OAI222_X1 U14239 ( .A1(P3_U3151), .A2(n11740), .B1(n11943), .B2(n11739), 
        .C1(n11738), .C2(n12944), .ZN(P3_U3270) );
  INV_X1 U14240 ( .A(n14383), .ZN(n14428) );
  NAND2_X1 U14241 ( .A1(n14383), .A2(n12320), .ZN(n11742) );
  NAND2_X1 U14242 ( .A1(n14288), .A2(n12322), .ZN(n11741) );
  NAND2_X1 U14243 ( .A1(n11742), .A2(n11741), .ZN(n11743) );
  XNOR2_X1 U14244 ( .A(n11743), .B(n12323), .ZN(n11782) );
  AND2_X1 U14245 ( .A1(n12321), .A2(n14288), .ZN(n11744) );
  AOI21_X1 U14246 ( .B1(n14383), .B2(n12322), .A(n11744), .ZN(n11783) );
  XNOR2_X1 U14247 ( .A(n11782), .B(n11783), .ZN(n11751) );
  INV_X1 U14248 ( .A(n11745), .ZN(n11746) );
  NAND2_X1 U14249 ( .A1(n11747), .A2(n11746), .ZN(n11752) );
  AND2_X1 U14250 ( .A1(n11751), .A2(n11752), .ZN(n11748) );
  NAND2_X1 U14251 ( .A1(n11749), .A2(n11748), .ZN(n11786) );
  INV_X1 U14252 ( .A(n11750), .ZN(n11755) );
  AOI21_X1 U14253 ( .B1(n11753), .B2(n11752), .A(n11751), .ZN(n11754) );
  OAI21_X1 U14254 ( .B1(n11755), .B2(n11754), .A(n13634), .ZN(n11759) );
  AOI22_X1 U14255 ( .A1(n14617), .A2(n13667), .B1(n13668), .B2(n14634), .ZN(
        n14379) );
  OAI21_X1 U14256 ( .B1(n13656), .B2(n14379), .A(n11756), .ZN(n11757) );
  AOI21_X1 U14257 ( .B1(n14381), .B2(n13654), .A(n11757), .ZN(n11758) );
  OAI211_X1 U14258 ( .C1(n14428), .C2(n13640), .A(n11759), .B(n11758), .ZN(
        P1_U3236) );
  OAI211_X1 U14259 ( .C1(n11762), .C2(n11761), .A(n11760), .B(n12473), .ZN(
        n11767) );
  NAND2_X1 U14260 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n14950) );
  INV_X1 U14261 ( .A(n14950), .ZN(n11765) );
  OAI22_X1 U14262 ( .A1(n12485), .A2(n15104), .B1(n12465), .B2(n11763), .ZN(
        n11764) );
  AOI211_X1 U14263 ( .C1(n12462), .C2(n12360), .A(n11765), .B(n11764), .ZN(
        n11766) );
  OAI211_X1 U14264 ( .C1(n11769), .C2(n11768), .A(n11767), .B(n11766), .ZN(
        P3_U3161) );
  NAND2_X1 U14265 ( .A1(n11774), .A2(n13492), .ZN(n11771) );
  OR2_X1 U14266 ( .A1(n11770), .A2(P2_U3088), .ZN(n12218) );
  OAI211_X1 U14267 ( .C1(n11772), .C2(n13498), .A(n11771), .B(n12218), .ZN(
        P2_U3304) );
  NAND2_X1 U14268 ( .A1(n11774), .A2(n11773), .ZN(n11776) );
  OAI211_X1 U14269 ( .C1(n11777), .C2(n7001), .A(n11776), .B(n11775), .ZN(
        P1_U3332) );
  NAND2_X1 U14270 ( .A1(n14290), .A2(n12320), .ZN(n11779) );
  NAND2_X1 U14271 ( .A1(n13667), .A2(n12322), .ZN(n11778) );
  NAND2_X1 U14272 ( .A1(n11779), .A2(n11778), .ZN(n11780) );
  XNOR2_X1 U14273 ( .A(n11780), .B(n12323), .ZN(n11869) );
  AND2_X1 U14274 ( .A1(n12321), .A2(n13667), .ZN(n11781) );
  AOI21_X1 U14275 ( .B1(n14290), .B2(n12322), .A(n11781), .ZN(n11870) );
  XNOR2_X1 U14276 ( .A(n11869), .B(n11870), .ZN(n11787) );
  INV_X1 U14277 ( .A(n11782), .ZN(n11784) );
  NAND2_X1 U14278 ( .A1(n11784), .A2(n11783), .ZN(n11788) );
  NAND2_X1 U14279 ( .A1(n11873), .A2(n13634), .ZN(n11797) );
  AOI21_X1 U14280 ( .B1(n11750), .B2(n11788), .A(n11787), .ZN(n11796) );
  INV_X1 U14281 ( .A(n11789), .ZN(n11791) );
  OAI22_X1 U14282 ( .A1(n13645), .A2(n11791), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11790), .ZN(n11794) );
  OAI22_X1 U14283 ( .A1(n14411), .A2(n13647), .B1(n13646), .B2(n11792), .ZN(
        n11793) );
  AOI211_X1 U14284 ( .C1(n14290), .C2(n13658), .A(n11794), .B(n11793), .ZN(
        n11795) );
  OAI21_X1 U14285 ( .B1(n11797), .B2(n11796), .A(n11795), .ZN(P1_U3224) );
  XNOR2_X1 U14286 ( .A(n11798), .B(n12993), .ZN(n12996) );
  XNOR2_X1 U14287 ( .A(n12996), .B(n11799), .ZN(n11800) );
  NAND2_X1 U14288 ( .A1(n11800), .A2(n13049), .ZN(n11806) );
  INV_X1 U14289 ( .A(n11801), .ZN(n11804) );
  AND2_X1 U14290 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n14724) );
  NOR2_X1 U14291 ( .A1(n13079), .A2(n11802), .ZN(n11803) );
  AOI211_X1 U14292 ( .C1(n13077), .C2(n11804), .A(n14724), .B(n11803), .ZN(
        n11805) );
  OAI211_X1 U14293 ( .C1(n9080), .C2(n8914), .A(n11806), .B(n11805), .ZN(
        P2_U3213) );
  AND2_X1 U14294 ( .A1(n11808), .A2(n11807), .ZN(n11810) );
  NAND2_X1 U14295 ( .A1(n11810), .A2(n11809), .ZN(n11812) );
  XNOR2_X1 U14296 ( .A(n11812), .B(n11811), .ZN(n15116) );
  OAI211_X1 U14297 ( .C1(n11815), .C2(n11814), .A(n11813), .B(n8938), .ZN(
        n11817) );
  AOI22_X1 U14298 ( .A1(n15062), .A2(n12360), .B1(n14333), .B2(n15059), .ZN(
        n11816) );
  NAND2_X1 U14299 ( .A1(n11817), .A2(n11816), .ZN(n11818) );
  AOI21_X1 U14300 ( .B1(n15116), .B2(n14997), .A(n11818), .ZN(n15118) );
  NOR2_X1 U14301 ( .A1(n11819), .A2(n15103), .ZN(n15114) );
  AOI22_X1 U14302 ( .A1(n15034), .A2(n15114), .B1(n15071), .B2(n12367), .ZN(
        n11820) );
  OAI21_X1 U14303 ( .B1(n11821), .B2(n15074), .A(n11820), .ZN(n11822) );
  AOI21_X1 U14304 ( .B1(n15116), .B2(n15072), .A(n11822), .ZN(n11823) );
  OAI21_X1 U14305 ( .B1(n15118), .B2(n15056), .A(n11823), .ZN(P3_U3223) );
  NOR2_X1 U14306 ( .A1(n11824), .A2(n15014), .ZN(n15013) );
  INV_X1 U14307 ( .A(n11825), .ZN(n11826) );
  NOR2_X1 U14308 ( .A1(n15013), .A2(n11826), .ZN(n15000) );
  NAND2_X1 U14309 ( .A1(n15000), .A2(n14999), .ZN(n14998) );
  NAND2_X1 U14310 ( .A1(n14998), .A2(n11827), .ZN(n11829) );
  XNOR2_X1 U14311 ( .A(n11829), .B(n11828), .ZN(n11830) );
  OAI222_X1 U14312 ( .A1(n15043), .A2(n11886), .B1(n15045), .B2(n15018), .C1(
        n11830), .C2(n15016), .ZN(n15098) );
  AOI21_X1 U14313 ( .B1(n15071), .B2(n11831), .A(n15098), .ZN(n11832) );
  MUX2_X1 U14314 ( .A(n14921), .B(n11832), .S(n15074), .Z(n11837) );
  OAI21_X1 U14315 ( .B1(n11704), .B2(n11834), .A(n11833), .ZN(n15100) );
  AOI22_X1 U14316 ( .A1(n15100), .A2(n14340), .B1(n11835), .B2(n12770), .ZN(
        n11836) );
  NAND2_X1 U14317 ( .A1(n11837), .A2(n11836), .ZN(P3_U3226) );
  NOR2_X1 U14318 ( .A1(n11852), .A2(n11838), .ZN(n11840) );
  NAND2_X1 U14319 ( .A1(n11864), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12516) );
  INV_X1 U14320 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n11841) );
  NAND2_X1 U14321 ( .A1(n11848), .A2(n11841), .ZN(n11842) );
  NAND2_X1 U14322 ( .A1(n12516), .A2(n11842), .ZN(n11854) );
  AOI21_X1 U14323 ( .B1(n11843), .B2(n11854), .A(n12507), .ZN(n11868) );
  NAND2_X1 U14324 ( .A1(n11845), .A2(n11844), .ZN(n11847) );
  NAND2_X1 U14325 ( .A1(n11847), .A2(n11846), .ZN(n11850) );
  NAND2_X1 U14326 ( .A1(n11864), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12515) );
  NAND2_X1 U14327 ( .A1(n11848), .A2(n12874), .ZN(n11849) );
  AND2_X1 U14328 ( .A1(n12515), .A2(n11849), .ZN(n11855) );
  NAND2_X1 U14329 ( .A1(n11855), .A2(n11850), .ZN(n12511) );
  OAI21_X1 U14330 ( .B1(n11850), .B2(n11855), .A(n12511), .ZN(n11866) );
  INV_X1 U14331 ( .A(n11851), .ZN(n11853) );
  NAND2_X1 U14332 ( .A1(n11853), .A2(n11852), .ZN(n11857) );
  AND2_X1 U14333 ( .A1(n11858), .A2(n11857), .ZN(n11860) );
  INV_X1 U14334 ( .A(n11854), .ZN(n11856) );
  MUX2_X1 U14335 ( .A(n11856), .B(n11855), .S(n11415), .Z(n11859) );
  NAND3_X1 U14336 ( .A1(n11858), .A2(n11859), .A3(n11857), .ZN(n12518) );
  OAI211_X1 U14337 ( .C1(n11860), .C2(n11859), .A(n14960), .B(n12518), .ZN(
        n11863) );
  INV_X1 U14338 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n11861) );
  NOR2_X1 U14339 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11861), .ZN(n11930) );
  AOI21_X1 U14340 ( .B1(n14978), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n11930), 
        .ZN(n11862) );
  OAI211_X1 U14341 ( .C1(n14982), .C2(n11864), .A(n11863), .B(n11862), .ZN(
        n11865) );
  AOI21_X1 U14342 ( .B1(n14992), .B2(n11866), .A(n11865), .ZN(n11867) );
  OAI21_X1 U14343 ( .B1(n11868), .B2(n14994), .A(n11867), .ZN(P3_U3196) );
  INV_X1 U14344 ( .A(n11870), .ZN(n11871) );
  NAND2_X1 U14345 ( .A1(n11869), .A2(n11871), .ZN(n11872) );
  AND2_X1 U14346 ( .A1(n12321), .A2(n14289), .ZN(n11874) );
  AOI21_X1 U14347 ( .B1(n14310), .B2(n12322), .A(n11874), .ZN(n12221) );
  AOI22_X1 U14348 ( .A1(n14310), .A2(n12320), .B1(n12322), .B2(n14289), .ZN(
        n11875) );
  XNOR2_X1 U14349 ( .A(n11875), .B(n12323), .ZN(n12220) );
  XOR2_X1 U14350 ( .A(n12221), .B(n12220), .Z(n12225) );
  XNOR2_X1 U14351 ( .A(n12226), .B(n12225), .ZN(n11880) );
  AOI22_X1 U14352 ( .A1(n9531), .A2(n14617), .B1(n14634), .B2(n13667), .ZN(
        n14304) );
  NAND2_X1 U14353 ( .A1(n13654), .A2(n14306), .ZN(n11877) );
  OAI211_X1 U14354 ( .C1(n14304), .C2(n13656), .A(n11877), .B(n11876), .ZN(
        n11878) );
  AOI21_X1 U14355 ( .B1(n14310), .B2(n13658), .A(n11878), .ZN(n11879) );
  OAI21_X1 U14356 ( .B1(n11880), .B2(n13660), .A(n11879), .ZN(P1_U3234) );
  INV_X1 U14357 ( .A(n11881), .ZN(n11882) );
  AOI21_X1 U14358 ( .B1(n11884), .B2(n11883), .A(n11882), .ZN(n11892) );
  NOR2_X1 U14359 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11885), .ZN(n14965) );
  INV_X1 U14360 ( .A(n12502), .ZN(n12452) );
  OAI22_X1 U14361 ( .A1(n12465), .A2(n11886), .B1(n12452), .B2(n12490), .ZN(
        n11887) );
  AOI211_X1 U14362 ( .C1(n11888), .C2(n12467), .A(n14965), .B(n11887), .ZN(
        n11891) );
  NAND2_X1 U14363 ( .A1(n12493), .A2(n11889), .ZN(n11890) );
  OAI211_X1 U14364 ( .C1(n11892), .C2(n12495), .A(n11891), .B(n11890), .ZN(
        P3_U3171) );
  XNOR2_X1 U14365 ( .A(n11894), .B(n11893), .ZN(n11895) );
  OAI222_X1 U14366 ( .A1(n15043), .A2(n12814), .B1(n15045), .B2(n12452), .C1(
        n11895), .C2(n15016), .ZN(n12879) );
  INV_X1 U14367 ( .A(n12879), .ZN(n11902) );
  OAI21_X1 U14368 ( .B1(n11898), .B2(n11897), .A(n11896), .ZN(n12880) );
  AOI22_X1 U14369 ( .A1(n15056), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n15071), 
        .B2(n12456), .ZN(n11899) );
  OAI21_X1 U14370 ( .B1(n12818), .B2(n12925), .A(n11899), .ZN(n11900) );
  AOI21_X1 U14371 ( .B1(n12880), .B2(n14340), .A(n11900), .ZN(n11901) );
  OAI21_X1 U14372 ( .B1(n11902), .B2(n15056), .A(n11901), .ZN(P3_U3222) );
  XNOR2_X1 U14373 ( .A(n11903), .B(n11904), .ZN(n14400) );
  INV_X1 U14374 ( .A(n14400), .ZN(n11916) );
  NAND2_X1 U14375 ( .A1(n11905), .A2(n11904), .ZN(n11906) );
  AOI21_X1 U14376 ( .B1(n11907), .B2(n11906), .A(n14533), .ZN(n14398) );
  AOI21_X1 U14377 ( .B1(n14371), .B2(n12244), .A(n10341), .ZN(n11908) );
  NAND2_X1 U14378 ( .A1(n11908), .A2(n13997), .ZN(n14396) );
  OR2_X1 U14379 ( .A1(n13966), .A2(n13584), .ZN(n11911) );
  INV_X1 U14380 ( .A(n11909), .ZN(n13587) );
  AOI22_X1 U14381 ( .A1(n14539), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n13587), 
        .B2(n14538), .ZN(n11910) );
  OAI211_X1 U14382 ( .C1(n14409), .C2(n13849), .A(n11911), .B(n11910), .ZN(
        n11912) );
  AOI21_X1 U14383 ( .B1(n12244), .B2(n14382), .A(n11912), .ZN(n11913) );
  OAI21_X1 U14384 ( .B1(n14396), .B2(n13902), .A(n11913), .ZN(n11914) );
  AOI21_X1 U14385 ( .B1(n14398), .B2(n14006), .A(n11914), .ZN(n11915) );
  OAI21_X1 U14386 ( .B1(n14009), .B2(n11916), .A(n11915), .ZN(P1_U3277) );
  XNOR2_X1 U14387 ( .A(n11918), .B(n14334), .ZN(n11919) );
  XNOR2_X1 U14388 ( .A(n11917), .B(n11919), .ZN(n11926) );
  NAND2_X1 U14389 ( .A1(n12493), .A2(n12816), .ZN(n11922) );
  AOI21_X1 U14390 ( .B1(n12462), .B2(n12486), .A(n11920), .ZN(n11921) );
  OAI211_X1 U14391 ( .C1(n12814), .C2(n12465), .A(n11922), .B(n11921), .ZN(
        n11923) );
  AOI21_X1 U14392 ( .B1(n11924), .B2(n12467), .A(n11923), .ZN(n11925) );
  OAI21_X1 U14393 ( .B1(n11926), .B2(n12495), .A(n11925), .ZN(P3_U3174) );
  XNOR2_X1 U14394 ( .A(n11928), .B(n12486), .ZN(n11929) );
  XNOR2_X1 U14395 ( .A(n11927), .B(n11929), .ZN(n11936) );
  INV_X1 U14396 ( .A(n14334), .ZN(n12803) );
  NAND2_X1 U14397 ( .A1(n12493), .A2(n12804), .ZN(n11932) );
  AOI21_X1 U14398 ( .B1(n12462), .B2(n12501), .A(n11930), .ZN(n11931) );
  OAI211_X1 U14399 ( .C1(n12803), .C2(n12465), .A(n11932), .B(n11931), .ZN(
        n11933) );
  AOI21_X1 U14400 ( .B1(n11934), .B2(n12467), .A(n11933), .ZN(n11935) );
  OAI21_X1 U14401 ( .B1(n11936), .B2(n12495), .A(n11935), .ZN(P3_U3155) );
  NAND2_X1 U14402 ( .A1(n11938), .A2(P3_D_REG_0__SCAN_IN), .ZN(n11937) );
  OAI21_X1 U14403 ( .B1(n11939), .B2(n11938), .A(n11937), .ZN(P3_U3376) );
  INV_X1 U14404 ( .A(n11940), .ZN(n11942) );
  OAI222_X1 U14405 ( .A1(n11944), .A2(P3_U3151), .B1(n11943), .B2(n11942), 
        .C1(n11941), .C2(n12944), .ZN(P3_U3269) );
  OAI222_X1 U14406 ( .A1(n11945), .A2(P1_U3086), .B1(n14160), .B2(n13485), 
        .C1(n9100), .C2(n7001), .ZN(P1_U3325) );
  NAND2_X1 U14407 ( .A1(n11946), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U14408 ( .A1(n12467), .A2(n11947), .B1(n12462), .B2(n12505), .ZN(
        n11948) );
  OAI211_X1 U14409 ( .C1(n11950), .C2(n12495), .A(n11949), .B(n11948), .ZN(
        P3_U3172) );
  OAI22_X1 U14410 ( .A1(n12926), .A2(n11954), .B1(n15119), .B2(n11951), .ZN(
        n11952) );
  INV_X1 U14411 ( .A(n11952), .ZN(n11953) );
  OAI21_X1 U14412 ( .B1(n11957), .B2(n8156), .A(n11953), .ZN(P3_U3390) );
  OAI22_X1 U14413 ( .A1(n12882), .A2(n11954), .B1(n15132), .B2(n10757), .ZN(
        n11955) );
  INV_X1 U14414 ( .A(n11955), .ZN(n11956) );
  OAI21_X1 U14415 ( .B1(n11957), .B2(n15130), .A(n11956), .ZN(P3_U3459) );
  OAI22_X1 U14416 ( .A1(n11959), .A2(n13354), .B1(n11958), .B2(n13357), .ZN(
        n11960) );
  AOI21_X1 U14417 ( .B1(n9078), .B2(n13366), .A(n11960), .ZN(n11963) );
  NAND2_X1 U14418 ( .A1(n11961), .A2(n13338), .ZN(n11962) );
  OAI211_X1 U14419 ( .C1(n11964), .C2(n13369), .A(n11963), .B(n11962), .ZN(
        n11965) );
  INV_X1 U14420 ( .A(n11965), .ZN(n11966) );
  OAI21_X1 U14421 ( .B1(n11967), .B2(n14761), .A(n11966), .ZN(P2_U3236) );
  NAND3_X1 U14422 ( .A1(n13114), .A2(n12155), .A3(n11968), .ZN(n11970) );
  AOI21_X1 U14423 ( .B1(n8912), .B2(n12131), .A(n12203), .ZN(n11971) );
  AOI21_X1 U14424 ( .B1(n6622), .B2(n11972), .A(n11971), .ZN(n11973) );
  OR2_X1 U14425 ( .A1(n13114), .A2(n11973), .ZN(n11974) );
  MUX2_X1 U14426 ( .A(n13112), .B(n14791), .S(n6622), .Z(n11976) );
  OR2_X1 U14427 ( .A1(n11977), .A2(n11976), .ZN(n11982) );
  NAND2_X1 U14428 ( .A1(n11977), .A2(n11976), .ZN(n11980) );
  MUX2_X1 U14429 ( .A(n14791), .B(n13112), .S(n6622), .Z(n11979) );
  NAND2_X1 U14430 ( .A1(n11980), .A2(n11979), .ZN(n11981) );
  MUX2_X1 U14431 ( .A(n11983), .B(n13111), .S(n6622), .Z(n11985) );
  INV_X1 U14432 ( .A(n11985), .ZN(n11986) );
  MUX2_X1 U14433 ( .A(n7497), .B(n11987), .S(n6622), .Z(n11991) );
  NAND2_X1 U14434 ( .A1(n11990), .A2(n11991), .ZN(n11989) );
  MUX2_X1 U14435 ( .A(n7497), .B(n11987), .S(n12155), .Z(n11988) );
  NAND2_X1 U14436 ( .A1(n11989), .A2(n11988), .ZN(n11995) );
  INV_X1 U14437 ( .A(n11990), .ZN(n11993) );
  INV_X1 U14438 ( .A(n11991), .ZN(n11992) );
  NAND2_X1 U14439 ( .A1(n11993), .A2(n11992), .ZN(n11994) );
  NAND2_X1 U14440 ( .A1(n11995), .A2(n11994), .ZN(n11997) );
  MUX2_X1 U14441 ( .A(n13031), .B(n13110), .S(n6622), .Z(n11998) );
  MUX2_X1 U14442 ( .A(n13031), .B(n13110), .S(n12155), .Z(n11996) );
  MUX2_X1 U14443 ( .A(n11999), .B(n13109), .S(n12155), .Z(n12001) );
  MUX2_X1 U14444 ( .A(n13109), .B(n11999), .S(n12155), .Z(n12000) );
  INV_X1 U14445 ( .A(n12001), .ZN(n12002) );
  MUX2_X1 U14446 ( .A(n14821), .B(n13108), .S(n6622), .Z(n12006) );
  NAND2_X1 U14447 ( .A1(n12005), .A2(n12006), .ZN(n12004) );
  MUX2_X1 U14448 ( .A(n14821), .B(n13108), .S(n12155), .Z(n12003) );
  NAND2_X1 U14449 ( .A1(n12004), .A2(n12003), .ZN(n12010) );
  INV_X1 U14450 ( .A(n12005), .ZN(n12008) );
  INV_X1 U14451 ( .A(n12006), .ZN(n12007) );
  NAND2_X1 U14452 ( .A1(n12008), .A2(n12007), .ZN(n12009) );
  MUX2_X1 U14453 ( .A(n13107), .B(n12011), .S(n6622), .Z(n12013) );
  MUX2_X1 U14454 ( .A(n13107), .B(n12011), .S(n12155), .Z(n12012) );
  INV_X1 U14455 ( .A(n12013), .ZN(n12014) );
  MUX2_X1 U14456 ( .A(n13106), .B(n12015), .S(n12155), .Z(n12018) );
  MUX2_X1 U14457 ( .A(n13106), .B(n12015), .S(n6622), .Z(n12016) );
  MUX2_X1 U14458 ( .A(n13105), .B(n12019), .S(n6622), .Z(n12021) );
  MUX2_X1 U14459 ( .A(n13105), .B(n12019), .S(n12155), .Z(n12020) );
  MUX2_X1 U14460 ( .A(n13104), .B(n12022), .S(n12155), .Z(n12026) );
  NAND2_X1 U14461 ( .A1(n12025), .A2(n12026), .ZN(n12024) );
  MUX2_X1 U14462 ( .A(n13104), .B(n12022), .S(n6622), .Z(n12023) );
  NAND2_X1 U14463 ( .A1(n12024), .A2(n12023), .ZN(n12030) );
  INV_X1 U14464 ( .A(n12025), .ZN(n12028) );
  INV_X1 U14465 ( .A(n12026), .ZN(n12027) );
  NAND2_X1 U14466 ( .A1(n12028), .A2(n12027), .ZN(n12029) );
  MUX2_X1 U14467 ( .A(n13103), .B(n12031), .S(n6622), .Z(n12033) );
  MUX2_X1 U14468 ( .A(n13103), .B(n12031), .S(n12155), .Z(n12032) );
  INV_X1 U14469 ( .A(n12033), .ZN(n12034) );
  MUX2_X1 U14470 ( .A(n13102), .B(n12035), .S(n12155), .Z(n12039) );
  NAND2_X1 U14471 ( .A1(n12038), .A2(n12039), .ZN(n12037) );
  MUX2_X1 U14472 ( .A(n13102), .B(n12035), .S(n6622), .Z(n12036) );
  NAND2_X1 U14473 ( .A1(n12037), .A2(n12036), .ZN(n12043) );
  INV_X1 U14474 ( .A(n12038), .ZN(n12041) );
  INV_X1 U14475 ( .A(n12039), .ZN(n12040) );
  NAND2_X1 U14476 ( .A1(n12041), .A2(n12040), .ZN(n12042) );
  NAND2_X1 U14477 ( .A1(n12043), .A2(n12042), .ZN(n12046) );
  MUX2_X1 U14478 ( .A(n13101), .B(n12044), .S(n6622), .Z(n12047) );
  MUX2_X1 U14479 ( .A(n13101), .B(n12044), .S(n12155), .Z(n12045) );
  INV_X1 U14480 ( .A(n12047), .ZN(n12048) );
  MUX2_X1 U14481 ( .A(n12050), .B(n12049), .S(n12155), .Z(n12059) );
  MUX2_X1 U14482 ( .A(n12051), .B(n9080), .S(n6622), .Z(n12065) );
  MUX2_X1 U14483 ( .A(n13099), .B(n12052), .S(n12155), .Z(n12064) );
  XNOR2_X1 U14484 ( .A(n13437), .B(n13061), .ZN(n13327) );
  INV_X1 U14485 ( .A(n13327), .ZN(n13329) );
  MUX2_X1 U14486 ( .A(n13098), .B(n13440), .S(n12155), .Z(n12063) );
  NAND2_X1 U14487 ( .A1(n13329), .A2(n12063), .ZN(n12057) );
  NAND2_X1 U14488 ( .A1(n13440), .A2(n6622), .ZN(n12054) );
  NAND2_X1 U14489 ( .A1(n13098), .A2(n12155), .ZN(n12053) );
  NAND4_X1 U14490 ( .A1(n12056), .A2(n12055), .A3(n12054), .A4(n12053), .ZN(
        n12071) );
  NAND2_X1 U14491 ( .A1(n12057), .A2(n12071), .ZN(n12066) );
  OAI21_X1 U14492 ( .B1(n12065), .B2(n12064), .A(n12066), .ZN(n12058) );
  MUX2_X1 U14493 ( .A(n13100), .B(n13452), .S(n6622), .Z(n12061) );
  NAND2_X1 U14494 ( .A1(n12062), .A2(n12061), .ZN(n12074) );
  INV_X1 U14495 ( .A(n12063), .ZN(n12072) );
  NAND3_X1 U14496 ( .A1(n12066), .A2(n12065), .A3(n12064), .ZN(n12070) );
  AND2_X1 U14497 ( .A1(n13097), .A2(n6622), .ZN(n12068) );
  OAI21_X1 U14498 ( .B1(n13097), .B2(n6622), .A(n13437), .ZN(n12067) );
  OAI21_X1 U14499 ( .B1(n12068), .B2(n13437), .A(n12067), .ZN(n12069) );
  OAI211_X1 U14500 ( .C1(n12072), .C2(n12071), .A(n12070), .B(n12069), .ZN(
        n12073) );
  MUX2_X1 U14501 ( .A(n12968), .B(n13323), .S(n12155), .Z(n12076) );
  NAND2_X1 U14502 ( .A1(n12075), .A2(n12076), .ZN(n12082) );
  INV_X1 U14503 ( .A(n12076), .ZN(n12077) );
  MUX2_X1 U14504 ( .A(n13096), .B(n13431), .S(n6622), .Z(n12079) );
  NAND2_X1 U14505 ( .A1(n12080), .A2(n12079), .ZN(n12081) );
  NAND2_X1 U14506 ( .A1(n12082), .A2(n12081), .ZN(n12085) );
  MUX2_X1 U14507 ( .A(n13095), .B(n13425), .S(n6622), .Z(n12086) );
  NAND2_X1 U14508 ( .A1(n12085), .A2(n12086), .ZN(n12084) );
  MUX2_X1 U14509 ( .A(n13095), .B(n13425), .S(n12155), .Z(n12083) );
  INV_X1 U14510 ( .A(n12085), .ZN(n12088) );
  INV_X1 U14511 ( .A(n12086), .ZN(n12087) );
  NAND2_X1 U14512 ( .A1(n12088), .A2(n12087), .ZN(n12089) );
  MUX2_X1 U14513 ( .A(n13094), .B(n13419), .S(n12155), .Z(n12091) );
  MUX2_X1 U14514 ( .A(n13094), .B(n13419), .S(n6622), .Z(n12090) );
  MUX2_X1 U14515 ( .A(n13093), .B(n13415), .S(n6622), .Z(n12093) );
  MUX2_X1 U14516 ( .A(n13093), .B(n13415), .S(n12155), .Z(n12092) );
  MUX2_X1 U14517 ( .A(n12977), .B(n13410), .S(n12155), .Z(n12097) );
  NAND2_X1 U14518 ( .A1(n12096), .A2(n12097), .ZN(n12095) );
  MUX2_X1 U14519 ( .A(n12977), .B(n13410), .S(n6622), .Z(n12094) );
  NAND2_X1 U14520 ( .A1(n12095), .A2(n12094), .ZN(n12101) );
  INV_X1 U14521 ( .A(n12096), .ZN(n12099) );
  INV_X1 U14522 ( .A(n12097), .ZN(n12098) );
  NAND2_X1 U14523 ( .A1(n12099), .A2(n12098), .ZN(n12100) );
  MUX2_X1 U14524 ( .A(n13092), .B(n13404), .S(n6622), .Z(n12103) );
  MUX2_X1 U14525 ( .A(n13092), .B(n13404), .S(n12155), .Z(n12102) );
  INV_X1 U14526 ( .A(n12103), .ZN(n12104) );
  MUX2_X1 U14527 ( .A(n13398), .B(n13091), .S(n6622), .Z(n12106) );
  MUX2_X1 U14528 ( .A(n13398), .B(n13091), .S(n12155), .Z(n12105) );
  INV_X1 U14529 ( .A(n12106), .ZN(n12107) );
  MUX2_X1 U14530 ( .A(n13090), .B(n13393), .S(n6622), .Z(n12111) );
  NAND2_X1 U14531 ( .A1(n12110), .A2(n12111), .ZN(n12109) );
  MUX2_X1 U14532 ( .A(n13090), .B(n13393), .S(n12155), .Z(n12108) );
  INV_X1 U14533 ( .A(n12110), .ZN(n12113) );
  INV_X1 U14534 ( .A(n12111), .ZN(n12112) );
  NAND2_X1 U14535 ( .A1(n12113), .A2(n12112), .ZN(n12114) );
  MUX2_X1 U14536 ( .A(n13089), .B(n13388), .S(n12155), .Z(n12116) );
  MUX2_X1 U14537 ( .A(n13388), .B(n13089), .S(n12155), .Z(n12115) );
  MUX2_X1 U14538 ( .A(n13088), .B(n13189), .S(n6622), .Z(n12120) );
  INV_X1 U14539 ( .A(n13087), .ZN(n12117) );
  MUX2_X1 U14540 ( .A(n12117), .B(n8916), .S(n12155), .Z(n12144) );
  MUX2_X1 U14541 ( .A(n13087), .B(n13377), .S(n6622), .Z(n12143) );
  OAI22_X1 U14542 ( .A1(n12121), .A2(n12120), .B1(n12144), .B2(n12143), .ZN(
        n12123) );
  MUX2_X1 U14543 ( .A(n13088), .B(n13189), .S(n12155), .Z(n12118) );
  INV_X1 U14544 ( .A(n12118), .ZN(n12119) );
  AOI21_X1 U14545 ( .B1(n12121), .B2(n12120), .A(n12119), .ZN(n12122) );
  NOR2_X1 U14546 ( .A1(n12123), .A2(n12122), .ZN(n12142) );
  NAND2_X1 U14547 ( .A1(n8285), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12124) );
  MUX2_X1 U14548 ( .A(n13085), .B(n13161), .S(n6622), .Z(n12151) );
  INV_X1 U14549 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n13151) );
  NAND2_X1 U14550 ( .A1(n12126), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n12129) );
  NAND2_X1 U14551 ( .A1(n12127), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n12128) );
  OAI211_X1 U14552 ( .C1(n12130), .C2(n13151), .A(n12129), .B(n12128), .ZN(
        n13152) );
  NAND2_X1 U14553 ( .A1(n13152), .A2(n6622), .ZN(n12156) );
  INV_X1 U14554 ( .A(n12161), .ZN(n12132) );
  OR2_X1 U14555 ( .A1(n12132), .A2(n12131), .ZN(n12205) );
  NAND4_X1 U14556 ( .A1(n12156), .A2(n12201), .A3(n12205), .A4(n12213), .ZN(
        n12133) );
  AND2_X1 U14557 ( .A1(n12133), .A2(n13085), .ZN(n12134) );
  AOI21_X1 U14558 ( .B1(n13161), .B2(n12155), .A(n12134), .ZN(n12150) );
  INV_X1 U14559 ( .A(n13086), .ZN(n12136) );
  MUX2_X1 U14560 ( .A(n13086), .B(n9078), .S(n6622), .Z(n12145) );
  OAI22_X1 U14561 ( .A1(n12151), .A2(n12150), .B1(n12146), .B2(n12145), .ZN(
        n12141) );
  NAND2_X1 U14562 ( .A1(n9021), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n12138) );
  NAND2_X1 U14563 ( .A1(n13370), .A2(n13152), .ZN(n12140) );
  NAND2_X1 U14564 ( .A1(n12141), .A2(n12197), .ZN(n12149) );
  NAND2_X1 U14565 ( .A1(n12142), .A2(n12149), .ZN(n12154) );
  AOI22_X1 U14566 ( .A1(n12146), .A2(n12145), .B1(n12144), .B2(n12143), .ZN(
        n12147) );
  NAND2_X1 U14567 ( .A1(n12197), .A2(n12147), .ZN(n12148) );
  NAND2_X1 U14568 ( .A1(n12149), .A2(n12148), .ZN(n12153) );
  NAND2_X1 U14569 ( .A1(n12151), .A2(n12150), .ZN(n12152) );
  NAND3_X1 U14570 ( .A1(n12154), .A2(n12153), .A3(n12152), .ZN(n12160) );
  NAND2_X1 U14571 ( .A1(n13370), .A2(n12155), .ZN(n12157) );
  NAND3_X1 U14572 ( .A1(n12158), .A2(n12157), .A3(n12156), .ZN(n12159) );
  XOR2_X1 U14573 ( .A(n13085), .B(n13161), .Z(n12195) );
  XNOR2_X1 U14574 ( .A(n13404), .B(n13019), .ZN(n13241) );
  NAND2_X1 U14575 ( .A1(n12162), .A2(n13269), .ZN(n13268) );
  NAND4_X1 U14576 ( .A1(n12165), .A2(n12164), .A3(n14785), .A4(n12163), .ZN(
        n12166) );
  NOR2_X1 U14577 ( .A1(n12167), .A2(n12166), .ZN(n12170) );
  NAND4_X1 U14578 ( .A1(n8988), .A2(n12170), .A3(n12169), .A4(n12168), .ZN(
        n12171) );
  NOR2_X1 U14579 ( .A1(n12172), .A2(n12171), .ZN(n12175) );
  NAND4_X1 U14580 ( .A1(n12176), .A2(n12175), .A3(n12174), .A4(n12173), .ZN(
        n12177) );
  NOR2_X1 U14581 ( .A1(n12178), .A2(n12177), .ZN(n12181) );
  NAND4_X1 U14582 ( .A1(n12182), .A2(n12181), .A3(n12180), .A4(n12179), .ZN(
        n12183) );
  NOR2_X1 U14583 ( .A1(n13327), .A2(n12183), .ZN(n12185) );
  NAND4_X1 U14584 ( .A1(n13314), .A2(n12185), .A3(n12184), .A4(n13349), .ZN(
        n12186) );
  NOR2_X1 U14585 ( .A1(n13268), .A2(n12186), .ZN(n12190) );
  NAND2_X1 U14586 ( .A1(n12188), .A2(n12187), .ZN(n13302) );
  NAND4_X1 U14587 ( .A1(n13254), .A2(n12190), .A3(n12189), .A4(n13302), .ZN(
        n12191) );
  NOR2_X1 U14588 ( .A1(n13241), .A2(n12191), .ZN(n12193) );
  NAND4_X1 U14589 ( .A1(n13205), .A2(n12193), .A3(n12192), .A4(n13230), .ZN(
        n12194) );
  NAND3_X1 U14590 ( .A1(n12198), .A2(n12197), .A3(n12196), .ZN(n12199) );
  INV_X1 U14591 ( .A(n12200), .ZN(n12212) );
  NAND2_X1 U14592 ( .A1(n8904), .A2(n12201), .ZN(n12202) );
  OAI211_X1 U14593 ( .C1(n12215), .C2(n12203), .A(n12213), .B(n12202), .ZN(
        n12204) );
  INV_X1 U14594 ( .A(n12204), .ZN(n12209) );
  OAI21_X1 U14595 ( .B1(n12206), .B2(n8904), .A(n12205), .ZN(n12207) );
  NAND2_X1 U14596 ( .A1(n12210), .A2(n12207), .ZN(n12208) );
  OAI21_X1 U14597 ( .B1(n12210), .B2(n12209), .A(n12208), .ZN(n12211) );
  NOR2_X1 U14598 ( .A1(n12212), .A2(n12211), .ZN(n12219) );
  NOR4_X1 U14599 ( .A1(n14772), .A2(n12214), .A3(n12213), .A4(n13060), .ZN(
        n12217) );
  OAI21_X1 U14600 ( .B1(n12218), .B2(n12215), .A(P2_B_REG_SCAN_IN), .ZN(n12216) );
  OAI22_X1 U14601 ( .A1(n12219), .A2(n12218), .B1(n12217), .B2(n12216), .ZN(
        P2_U3328) );
  INV_X1 U14602 ( .A(n12220), .ZN(n12223) );
  INV_X1 U14603 ( .A(n12221), .ZN(n12222) );
  NOR2_X1 U14604 ( .A1(n12229), .A2(n10612), .ZN(n12227) );
  AOI21_X1 U14605 ( .B1(n14414), .B2(n12320), .A(n12227), .ZN(n12228) );
  XNOR2_X1 U14606 ( .A(n12228), .B(n12323), .ZN(n12232) );
  NOR2_X1 U14607 ( .A1(n12229), .A2(n10954), .ZN(n12230) );
  AOI21_X1 U14608 ( .B1(n14414), .B2(n12322), .A(n12230), .ZN(n12231) );
  NAND2_X1 U14609 ( .A1(n12232), .A2(n12231), .ZN(n12234) );
  OAI21_X1 U14610 ( .B1(n12232), .B2(n12231), .A(n12234), .ZN(n12233) );
  INV_X1 U14611 ( .A(n12233), .ZN(n13519) );
  NAND2_X1 U14612 ( .A1(n14366), .A2(n12320), .ZN(n12236) );
  OR2_X1 U14613 ( .A1(n14409), .A2(n10612), .ZN(n12235) );
  NAND2_X1 U14614 ( .A1(n12236), .A2(n12235), .ZN(n12237) );
  XNOR2_X1 U14615 ( .A(n12237), .B(n12323), .ZN(n12239) );
  INV_X1 U14616 ( .A(n14366), .ZN(n14402) );
  OAI22_X1 U14617 ( .A1(n14402), .A2(n10612), .B1(n14409), .B2(n10954), .ZN(
        n13652) );
  INV_X1 U14618 ( .A(n12238), .ZN(n12240) );
  NAND2_X1 U14619 ( .A1(n12244), .A2(n12320), .ZN(n12242) );
  NAND2_X1 U14620 ( .A1(n13666), .A2(n12322), .ZN(n12241) );
  NAND2_X1 U14621 ( .A1(n12242), .A2(n12241), .ZN(n12243) );
  XNOR2_X1 U14622 ( .A(n12243), .B(n12323), .ZN(n12248) );
  NAND2_X1 U14623 ( .A1(n12244), .A2(n12322), .ZN(n12246) );
  NAND2_X1 U14624 ( .A1(n12321), .A2(n13666), .ZN(n12245) );
  NAND2_X1 U14625 ( .A1(n12246), .A2(n12245), .ZN(n12247) );
  NOR2_X1 U14626 ( .A1(n12248), .A2(n12247), .ZN(n12249) );
  AOI21_X1 U14627 ( .B1(n12248), .B2(n12247), .A(n12249), .ZN(n13581) );
  INV_X1 U14628 ( .A(n12249), .ZN(n12250) );
  NAND2_X1 U14629 ( .A1(n14116), .A2(n12320), .ZN(n12252) );
  OR2_X1 U14630 ( .A1(n13584), .A2(n10612), .ZN(n12251) );
  NAND2_X1 U14631 ( .A1(n12252), .A2(n12251), .ZN(n12253) );
  XNOR2_X1 U14632 ( .A(n12253), .B(n11177), .ZN(n12256) );
  NOR2_X1 U14633 ( .A1(n13584), .A2(n10954), .ZN(n12254) );
  AOI21_X1 U14634 ( .B1(n14116), .B2(n12322), .A(n12254), .ZN(n12255) );
  NOR2_X1 U14635 ( .A1(n12256), .A2(n12255), .ZN(n13592) );
  NAND2_X1 U14636 ( .A1(n12256), .A2(n12255), .ZN(n13590) );
  OAI22_X1 U14637 ( .A1(n13985), .A2(n10612), .B1(n14102), .B2(n10954), .ZN(
        n12258) );
  OAI22_X1 U14638 ( .A1(n13985), .A2(n10348), .B1(n14102), .B2(n10612), .ZN(
        n12257) );
  XNOR2_X1 U14639 ( .A(n12257), .B(n12323), .ZN(n12259) );
  XOR2_X1 U14640 ( .A(n12258), .B(n12259), .Z(n13633) );
  NAND2_X1 U14641 ( .A1(n13631), .A2(n12260), .ZN(n13547) );
  INV_X1 U14642 ( .A(n13547), .ZN(n12266) );
  AND2_X1 U14643 ( .A1(n13665), .A2(n12321), .ZN(n12261) );
  AOI21_X1 U14644 ( .B1(n14106), .B2(n12322), .A(n12261), .ZN(n12268) );
  NAND2_X1 U14645 ( .A1(n14106), .A2(n12320), .ZN(n12263) );
  NAND2_X1 U14646 ( .A1(n13665), .A2(n12322), .ZN(n12262) );
  NAND2_X1 U14647 ( .A1(n12263), .A2(n12262), .ZN(n12264) );
  XNOR2_X1 U14648 ( .A(n12264), .B(n12323), .ZN(n12267) );
  XOR2_X1 U14649 ( .A(n12268), .B(n12267), .Z(n13548) );
  INV_X1 U14650 ( .A(n13548), .ZN(n12265) );
  INV_X1 U14651 ( .A(n12267), .ZN(n12269) );
  OAI22_X1 U14652 ( .A1(n14096), .A2(n10612), .B1(n14103), .B2(n10954), .ZN(
        n12271) );
  OAI22_X1 U14653 ( .A1(n14096), .A2(n10348), .B1(n14103), .B2(n10612), .ZN(
        n12270) );
  XNOR2_X1 U14654 ( .A(n12270), .B(n12323), .ZN(n12272) );
  XOR2_X1 U14655 ( .A(n12271), .B(n12272), .Z(n13612) );
  NAND2_X1 U14656 ( .A1(n12272), .A2(n12271), .ZN(n12273) );
  AOI22_X1 U14657 ( .A1(n14088), .A2(n12322), .B1(n12321), .B2(n14076), .ZN(
        n12276) );
  AOI22_X1 U14658 ( .A1(n14088), .A2(n12320), .B1(n12322), .B2(n14076), .ZN(
        n12274) );
  XNOR2_X1 U14659 ( .A(n12274), .B(n12323), .ZN(n12275) );
  XOR2_X1 U14660 ( .A(n12276), .B(n12275), .Z(n13563) );
  INV_X1 U14661 ( .A(n12275), .ZN(n12278) );
  INV_X1 U14662 ( .A(n12276), .ZN(n12277) );
  AND2_X1 U14663 ( .A1(n12321), .A2(n13664), .ZN(n12279) );
  AOI21_X1 U14664 ( .B1(n13913), .B2(n12322), .A(n12279), .ZN(n12281) );
  AOI22_X1 U14665 ( .A1(n13913), .A2(n12320), .B1(n12322), .B2(n13664), .ZN(
        n12280) );
  XNOR2_X1 U14666 ( .A(n12280), .B(n12323), .ZN(n12282) );
  XOR2_X1 U14667 ( .A(n12281), .B(n12282), .Z(n13622) );
  NAND2_X1 U14668 ( .A1(n13621), .A2(n13622), .ZN(n13620) );
  NAND2_X1 U14669 ( .A1(n12282), .A2(n12281), .ZN(n12283) );
  NAND2_X1 U14670 ( .A1(n13620), .A2(n12283), .ZN(n13526) );
  OAI22_X1 U14671 ( .A1(n14071), .A2(n10612), .B1(n13916), .B2(n10954), .ZN(
        n12287) );
  OAI22_X1 U14672 ( .A1(n14071), .A2(n10348), .B1(n13916), .B2(n10612), .ZN(
        n12285) );
  XNOR2_X1 U14673 ( .A(n12285), .B(n12323), .ZN(n12286) );
  XOR2_X1 U14674 ( .A(n12287), .B(n12286), .Z(n13527) );
  NAND2_X1 U14675 ( .A1(n13526), .A2(n13527), .ZN(n12291) );
  INV_X1 U14676 ( .A(n12286), .ZN(n12289) );
  INV_X1 U14677 ( .A(n12287), .ZN(n12288) );
  NAND2_X1 U14678 ( .A1(n12289), .A2(n12288), .ZN(n12290) );
  NAND2_X1 U14679 ( .A1(n12291), .A2(n12290), .ZN(n13603) );
  NAND2_X1 U14680 ( .A1(n14066), .A2(n12320), .ZN(n12293) );
  NAND2_X1 U14681 ( .A1(n13860), .A2(n12322), .ZN(n12292) );
  NAND2_X1 U14682 ( .A1(n12293), .A2(n12292), .ZN(n12294) );
  XNOR2_X1 U14683 ( .A(n12294), .B(n12323), .ZN(n12295) );
  AOI22_X1 U14684 ( .A1(n14066), .A2(n12322), .B1(n12321), .B2(n13860), .ZN(
        n12296) );
  XNOR2_X1 U14685 ( .A(n12295), .B(n12296), .ZN(n13604) );
  NAND2_X1 U14686 ( .A1(n13603), .A2(n13604), .ZN(n12299) );
  INV_X1 U14687 ( .A(n12295), .ZN(n12297) );
  NAND2_X1 U14688 ( .A1(n12297), .A2(n12296), .ZN(n12298) );
  NAND2_X1 U14689 ( .A1(n14057), .A2(n12320), .ZN(n12301) );
  NAND2_X1 U14690 ( .A1(n14046), .A2(n12322), .ZN(n12300) );
  NAND2_X1 U14691 ( .A1(n12301), .A2(n12300), .ZN(n12302) );
  XNOR2_X1 U14692 ( .A(n12302), .B(n12323), .ZN(n12303) );
  AOI22_X1 U14693 ( .A1(n14057), .A2(n12322), .B1(n12321), .B2(n14046), .ZN(
        n12304) );
  XNOR2_X1 U14694 ( .A(n12303), .B(n12304), .ZN(n13571) );
  INV_X1 U14695 ( .A(n12303), .ZN(n12305) );
  NAND2_X1 U14696 ( .A1(n12305), .A2(n12304), .ZN(n12306) );
  NAND2_X1 U14697 ( .A1(n13851), .A2(n12320), .ZN(n12308) );
  NAND2_X1 U14698 ( .A1(n13859), .A2(n12322), .ZN(n12307) );
  NAND2_X1 U14699 ( .A1(n12308), .A2(n12307), .ZN(n12309) );
  XNOR2_X1 U14700 ( .A(n12309), .B(n12323), .ZN(n12312) );
  AOI22_X1 U14701 ( .A1(n13851), .A2(n12322), .B1(n12321), .B2(n13859), .ZN(
        n12310) );
  XNOR2_X1 U14702 ( .A(n12312), .B(n12310), .ZN(n13642) );
  INV_X1 U14703 ( .A(n12310), .ZN(n12311) );
  NAND2_X1 U14704 ( .A1(n14042), .A2(n12320), .ZN(n12315) );
  NAND2_X1 U14705 ( .A1(n14047), .A2(n12322), .ZN(n12314) );
  NAND2_X1 U14706 ( .A1(n12315), .A2(n12314), .ZN(n12316) );
  XNOR2_X1 U14707 ( .A(n12316), .B(n12323), .ZN(n12317) );
  AOI22_X1 U14708 ( .A1(n14042), .A2(n12322), .B1(n12321), .B2(n14047), .ZN(
        n12318) );
  XNOR2_X1 U14709 ( .A(n12317), .B(n12318), .ZN(n13510) );
  INV_X1 U14710 ( .A(n12317), .ZN(n12319) );
  AOI22_X1 U14711 ( .A1(n13821), .A2(n12313), .B1(n12322), .B2(n13663), .ZN(
        n12326) );
  AOI22_X1 U14712 ( .A1(n13821), .A2(n12322), .B1(n12321), .B2(n13663), .ZN(
        n12324) );
  XNOR2_X1 U14713 ( .A(n12324), .B(n12323), .ZN(n12325) );
  XOR2_X1 U14714 ( .A(n12326), .B(n12325), .Z(n12327) );
  XNOR2_X1 U14715 ( .A(n12328), .B(n12327), .ZN(n12334) );
  INV_X1 U14716 ( .A(n13817), .ZN(n12330) );
  OAI22_X1 U14717 ( .A1(n13645), .A2(n12330), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12329), .ZN(n12332) );
  OAI22_X1 U14718 ( .A1(n13816), .A2(n13647), .B1(n13646), .B2(n13845), .ZN(
        n12331) );
  AOI211_X1 U14719 ( .C1(n13821), .C2(n13658), .A(n12332), .B(n12331), .ZN(
        n12333) );
  OAI21_X1 U14720 ( .B1(n12334), .B2(n13660), .A(n12333), .ZN(P1_U3220) );
  XNOR2_X1 U14721 ( .A(n12336), .B(n12335), .ZN(n12344) );
  INV_X1 U14722 ( .A(n12344), .ZN(n12337) );
  NAND2_X1 U14723 ( .A1(n12337), .A2(n12473), .ZN(n12350) );
  INV_X1 U14724 ( .A(n12338), .ZN(n12339) );
  NAND4_X1 U14725 ( .A1(n12349), .A2(n12473), .A3(n12339), .A4(n12344), .ZN(
        n12348) );
  AOI22_X1 U14726 ( .A1(n12499), .A2(n12487), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12341) );
  NAND2_X1 U14727 ( .A1(n12493), .A2(n12627), .ZN(n12340) );
  OAI211_X1 U14728 ( .C1(n12342), .C2(n12490), .A(n12341), .B(n12340), .ZN(
        n12346) );
  NOR4_X1 U14729 ( .A1(n12344), .A2(n12343), .A3(n12495), .A4(n12499), .ZN(
        n12345) );
  AOI211_X1 U14730 ( .C1(n12631), .C2(n12467), .A(n12346), .B(n12345), .ZN(
        n12347) );
  OAI211_X1 U14731 ( .C1(n12350), .C2(n12349), .A(n12348), .B(n12347), .ZN(
        P3_U3160) );
  INV_X1 U14732 ( .A(n12351), .ZN(n12353) );
  OAI222_X1 U14733 ( .A1(P3_U3151), .A2(n7002), .B1(n11943), .B2(n12353), .C1(
        n12352), .C2(n12944), .ZN(P3_U3265) );
  NOR2_X1 U14734 ( .A1(n12354), .A2(n12668), .ZN(n12427) );
  AOI21_X1 U14735 ( .B1(n12668), .B2(n12354), .A(n12427), .ZN(n12359) );
  NAND2_X1 U14736 ( .A1(n12493), .A2(n12685), .ZN(n12356) );
  AOI22_X1 U14737 ( .A1(n12682), .A2(n12462), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12355) );
  OAI211_X1 U14738 ( .C1(n12711), .C2(n12465), .A(n12356), .B(n12355), .ZN(
        n12357) );
  AOI21_X1 U14739 ( .B1(n12689), .B2(n12467), .A(n12357), .ZN(n12358) );
  OAI21_X1 U14740 ( .B1(n12359), .B2(n12495), .A(n12358), .ZN(P3_U3156) );
  AOI22_X1 U14741 ( .A1(n12467), .A2(n12361), .B1(n12487), .B2(n12360), .ZN(
        n12362) );
  NAND2_X1 U14742 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n14980)
         );
  OAI211_X1 U14743 ( .C1(n12450), .C2(n12490), .A(n12362), .B(n14980), .ZN(
        n12366) );
  AOI211_X1 U14744 ( .C1(n12364), .C2(n12363), .A(n12495), .B(n7544), .ZN(
        n12365) );
  AOI211_X1 U14745 ( .C1(n12367), .C2(n12493), .A(n12366), .B(n12365), .ZN(
        n12368) );
  INV_X1 U14746 ( .A(n12368), .ZN(P3_U3157) );
  XNOR2_X1 U14747 ( .A(n12369), .B(n12370), .ZN(n12375) );
  NAND2_X1 U14748 ( .A1(n12487), .A2(n12734), .ZN(n12371) );
  NAND2_X1 U14749 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12606)
         );
  OAI211_X1 U14750 ( .C1(n12710), .C2(n12490), .A(n12371), .B(n12606), .ZN(
        n12373) );
  NOR2_X1 U14751 ( .A1(n12901), .A2(n12485), .ZN(n12372) );
  AOI211_X1 U14752 ( .C1(n12737), .C2(n12493), .A(n12373), .B(n12372), .ZN(
        n12374) );
  OAI21_X1 U14753 ( .B1(n12375), .B2(n12495), .A(n12374), .ZN(P3_U3159) );
  INV_X1 U14754 ( .A(n12377), .ZN(n12378) );
  AOI21_X1 U14755 ( .B1(n12379), .B2(n12376), .A(n12378), .ZN(n12385) );
  NAND2_X1 U14756 ( .A1(n12493), .A2(n12712), .ZN(n12381) );
  AOI22_X1 U14757 ( .A1(n12462), .A2(n12681), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12380) );
  OAI211_X1 U14758 ( .C1(n12710), .C2(n12465), .A(n12381), .B(n12380), .ZN(
        n12382) );
  AOI21_X1 U14759 ( .B1(n12383), .B2(n12467), .A(n12382), .ZN(n12384) );
  OAI21_X1 U14760 ( .B1(n12385), .B2(n12495), .A(n12384), .ZN(P3_U3163) );
  XNOR2_X1 U14761 ( .A(n12386), .B(n12387), .ZN(n12451) );
  OAI22_X1 U14762 ( .A1(n12451), .A2(n14333), .B1(n12386), .B2(n12387), .ZN(
        n12390) );
  XNOR2_X1 U14763 ( .A(n12388), .B(n12455), .ZN(n12389) );
  XNOR2_X1 U14764 ( .A(n12390), .B(n12389), .ZN(n12395) );
  OAI22_X1 U14765 ( .A1(n12485), .A2(n14339), .B1(n12465), .B2(n12450), .ZN(
        n12391) );
  AOI211_X1 U14766 ( .C1(n12462), .C2(n14334), .A(n12392), .B(n12391), .ZN(
        n12394) );
  NAND2_X1 U14767 ( .A1(n12493), .A2(n14336), .ZN(n12393) );
  OAI211_X1 U14768 ( .C1(n12395), .C2(n12495), .A(n12394), .B(n12393), .ZN(
        P3_U3164) );
  INV_X1 U14769 ( .A(n12398), .ZN(n12400) );
  NOR3_X1 U14770 ( .A1(n12428), .A2(n12400), .A3(n12399), .ZN(n12403) );
  INV_X1 U14771 ( .A(n12401), .ZN(n12402) );
  OAI21_X1 U14772 ( .B1(n12403), .B2(n12402), .A(n12473), .ZN(n12408) );
  AOI22_X1 U14773 ( .A1(n12656), .A2(n12462), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12404) );
  OAI21_X1 U14774 ( .B1(n12405), .B2(n12465), .A(n12404), .ZN(n12406) );
  AOI21_X1 U14775 ( .B1(n12493), .B2(n12659), .A(n12406), .ZN(n12407) );
  OAI211_X1 U14776 ( .C1(n12886), .C2(n12485), .A(n12408), .B(n12407), .ZN(
        P3_U3165) );
  XNOR2_X1 U14777 ( .A(n12410), .B(n12409), .ZN(n12415) );
  NAND2_X1 U14778 ( .A1(n12487), .A2(n12501), .ZN(n12411) );
  NAND2_X1 U14779 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12536)
         );
  OAI211_X1 U14780 ( .C1(n12778), .C2(n12490), .A(n12411), .B(n12536), .ZN(
        n12412) );
  AOI21_X1 U14781 ( .B1(n12493), .B2(n12780), .A(n12412), .ZN(n12414) );
  NAND2_X1 U14782 ( .A1(n12779), .A2(n12467), .ZN(n12413) );
  OAI211_X1 U14783 ( .C1(n12415), .C2(n12495), .A(n12414), .B(n12413), .ZN(
        P3_U3166) );
  XNOR2_X1 U14784 ( .A(n12416), .B(n12417), .ZN(n12423) );
  NAND2_X1 U14785 ( .A1(n12493), .A2(n12765), .ZN(n12420) );
  NOR2_X1 U14786 ( .A1(n12418), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12559) );
  AOI21_X1 U14787 ( .B1(n12462), .B2(n12734), .A(n12559), .ZN(n12419) );
  OAI211_X1 U14788 ( .C1(n12792), .C2(n12465), .A(n12420), .B(n12419), .ZN(
        n12421) );
  AOI21_X1 U14789 ( .B1(n12860), .B2(n12467), .A(n12421), .ZN(n12422) );
  OAI21_X1 U14790 ( .B1(n12423), .B2(n12495), .A(n12422), .ZN(P3_U3168) );
  INV_X1 U14791 ( .A(n12424), .ZN(n12426) );
  NOR3_X1 U14792 ( .A1(n12427), .A2(n12426), .A3(n12425), .ZN(n12429) );
  OAI21_X1 U14793 ( .B1(n12429), .B2(n12428), .A(n12473), .ZN(n12433) );
  AOI22_X1 U14794 ( .A1(n12668), .A2(n12487), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12430) );
  OAI21_X1 U14795 ( .B1(n12671), .B2(n12490), .A(n12430), .ZN(n12431) );
  AOI21_X1 U14796 ( .B1(n12493), .B2(n12673), .A(n12431), .ZN(n12432) );
  OAI211_X1 U14797 ( .C1(n12675), .C2(n12485), .A(n12433), .B(n12432), .ZN(
        P3_U3169) );
  XNOR2_X1 U14798 ( .A(n12434), .B(n12435), .ZN(n12440) );
  INV_X1 U14799 ( .A(n12721), .ZN(n12750) );
  NAND2_X1 U14800 ( .A1(n12493), .A2(n12725), .ZN(n12437) );
  AOI22_X1 U14801 ( .A1(n12462), .A2(n12722), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12436) );
  OAI211_X1 U14802 ( .C1(n12750), .C2(n12465), .A(n12437), .B(n12436), .ZN(
        n12438) );
  AOI21_X1 U14803 ( .B1(n12848), .B2(n12467), .A(n12438), .ZN(n12439) );
  OAI21_X1 U14804 ( .B1(n12440), .B2(n12495), .A(n12439), .ZN(P3_U3173) );
  INV_X1 U14805 ( .A(n12442), .ZN(n12443) );
  AOI21_X1 U14806 ( .B1(n12681), .B2(n12441), .A(n12443), .ZN(n12449) );
  NAND2_X1 U14807 ( .A1(n12493), .A2(n12701), .ZN(n12445) );
  AOI22_X1 U14808 ( .A1(n12668), .A2(n12462), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12444) );
  OAI211_X1 U14809 ( .C1(n12700), .C2(n12465), .A(n12445), .B(n12444), .ZN(
        n12446) );
  AOI21_X1 U14810 ( .B1(n12447), .B2(n12467), .A(n12446), .ZN(n12448) );
  OAI21_X1 U14811 ( .B1(n12449), .B2(n12495), .A(n12448), .ZN(P3_U3175) );
  XNOR2_X1 U14812 ( .A(n12451), .B(n12450), .ZN(n12459) );
  OAI22_X1 U14813 ( .A1(n12485), .A2(n12925), .B1(n12465), .B2(n12452), .ZN(
        n12453) );
  AOI211_X1 U14814 ( .C1(n12462), .C2(n12455), .A(n12454), .B(n12453), .ZN(
        n12458) );
  NAND2_X1 U14815 ( .A1(n12493), .A2(n12456), .ZN(n12457) );
  OAI211_X1 U14816 ( .C1(n12459), .C2(n12495), .A(n12458), .B(n12457), .ZN(
        P3_U3176) );
  XNOR2_X1 U14817 ( .A(n12460), .B(n12461), .ZN(n12469) );
  NAND2_X1 U14818 ( .A1(n12493), .A2(n12752), .ZN(n12464) );
  INV_X1 U14819 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n15378) );
  NOR2_X1 U14820 ( .A1(n15378), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12580) );
  AOI21_X1 U14821 ( .B1(n12462), .B2(n12721), .A(n12580), .ZN(n12463) );
  OAI211_X1 U14822 ( .C1(n12778), .C2(n12465), .A(n12464), .B(n12463), .ZN(
        n12466) );
  AOI21_X1 U14823 ( .B1(n12751), .B2(n12467), .A(n12466), .ZN(n12468) );
  OAI21_X1 U14824 ( .B1(n12469), .B2(n12495), .A(n12468), .ZN(P3_U3178) );
  OAI21_X1 U14825 ( .B1(n12472), .B2(n12470), .A(n12471), .ZN(n12474) );
  NAND2_X1 U14826 ( .A1(n12474), .A2(n12473), .ZN(n12480) );
  AOI22_X1 U14827 ( .A1(n12475), .A2(n12487), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12476) );
  OAI21_X1 U14828 ( .B1(n12477), .B2(n12490), .A(n12476), .ZN(n12478) );
  AOI21_X1 U14829 ( .B1(n12645), .B2(n12493), .A(n12478), .ZN(n12479) );
  OAI211_X1 U14830 ( .C1(n12826), .C2(n12485), .A(n12480), .B(n12479), .ZN(
        P3_U3180) );
  XNOR2_X1 U14831 ( .A(n12481), .B(n12501), .ZN(n12482) );
  XNOR2_X1 U14832 ( .A(n12483), .B(n12482), .ZN(n12496) );
  INV_X1 U14833 ( .A(n12484), .ZN(n12914) );
  NOR2_X1 U14834 ( .A1(n12914), .A2(n12485), .ZN(n12492) );
  NAND2_X1 U14835 ( .A1(n12487), .A2(n12486), .ZN(n12489) );
  NAND2_X1 U14836 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12513)
         );
  OAI211_X1 U14837 ( .C1(n12792), .C2(n12490), .A(n12489), .B(n12513), .ZN(
        n12491) );
  AOI211_X1 U14838 ( .C1(n12493), .C2(n12793), .A(n12492), .B(n12491), .ZN(
        n12494) );
  OAI21_X1 U14839 ( .B1(n12496), .B2(n12495), .A(n12494), .ZN(P3_U3181) );
  MUX2_X1 U14840 ( .A(n12497), .B(P3_DATAO_REG_29__SCAN_IN), .S(n12506), .Z(
        P3_U3520) );
  MUX2_X1 U14841 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12498), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14842 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12499), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14843 ( .A(n12656), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12506), .Z(
        P3_U3517) );
  MUX2_X1 U14844 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12668), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14845 ( .A(n12681), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12506), .Z(
        P3_U3513) );
  MUX2_X1 U14846 ( .A(n12722), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12506), .Z(
        P3_U3512) );
  MUX2_X1 U14847 ( .A(n12733), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12506), .Z(
        P3_U3511) );
  MUX2_X1 U14848 ( .A(n12721), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12506), .Z(
        P3_U3510) );
  MUX2_X1 U14849 ( .A(n12734), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12506), .Z(
        P3_U3509) );
  MUX2_X1 U14850 ( .A(n12500), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12506), .Z(
        P3_U3508) );
  MUX2_X1 U14851 ( .A(n12501), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12506), .Z(
        P3_U3506) );
  MUX2_X1 U14852 ( .A(n14334), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12506), .Z(
        P3_U3504) );
  MUX2_X1 U14853 ( .A(n14333), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12506), .Z(
        P3_U3502) );
  MUX2_X1 U14854 ( .A(n12502), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12506), .Z(
        P3_U3501) );
  MUX2_X1 U14855 ( .A(n15001), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12506), .Z(
        P3_U3498) );
  MUX2_X1 U14856 ( .A(n12503), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12506), .Z(
        P3_U3497) );
  MUX2_X1 U14857 ( .A(n15002), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12506), .Z(
        P3_U3496) );
  MUX2_X1 U14858 ( .A(n15026), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12506), .Z(
        P3_U3495) );
  MUX2_X1 U14859 ( .A(n12504), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12506), .Z(
        P3_U3494) );
  MUX2_X1 U14860 ( .A(n15060), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12506), .Z(
        P3_U3493) );
  MUX2_X1 U14861 ( .A(n12505), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12506), .Z(
        P3_U3492) );
  MUX2_X1 U14862 ( .A(n15061), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12506), .Z(
        P3_U3491) );
  INV_X1 U14863 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12510) );
  NAND2_X1 U14864 ( .A1(n12516), .A2(n12508), .ZN(n12527) );
  AOI21_X1 U14865 ( .B1(n12510), .B2(n12509), .A(n12528), .ZN(n12526) );
  NAND2_X1 U14866 ( .A1(n12515), .A2(n12511), .ZN(n12532) );
  OAI21_X1 U14867 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12512), .A(n12534), 
        .ZN(n12524) );
  INV_X1 U14868 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14196) );
  NAND2_X1 U14869 ( .A1(n14915), .A2(n6955), .ZN(n12514) );
  OAI211_X1 U14870 ( .C1(n14196), .C2(n14952), .A(n12514), .B(n12513), .ZN(
        n12523) );
  MUX2_X1 U14871 ( .A(n12516), .B(n12515), .S(n11415), .Z(n12517) );
  NAND2_X1 U14872 ( .A1(n12518), .A2(n12517), .ZN(n12540) );
  XNOR2_X1 U14873 ( .A(n12540), .B(n12533), .ZN(n12520) );
  MUX2_X1 U14874 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n11415), .Z(n12519) );
  NOR2_X1 U14875 ( .A1(n12520), .A2(n12519), .ZN(n12541) );
  AOI21_X1 U14876 ( .B1(n12520), .B2(n12519), .A(n12541), .ZN(n12521) );
  NOR2_X1 U14877 ( .A1(n12521), .A2(n14986), .ZN(n12522) );
  AOI211_X1 U14878 ( .C1(n14992), .C2(n12524), .A(n12523), .B(n12522), .ZN(
        n12525) );
  OAI21_X1 U14879 ( .B1(n12526), .B2(n14994), .A(n12525), .ZN(P3_U3197) );
  INV_X1 U14880 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12543) );
  MUX2_X1 U14881 ( .A(n12543), .B(P3_REG2_REG_16__SCAN_IN), .S(n12556), .Z(
        n12530) );
  INV_X1 U14882 ( .A(n12553), .ZN(n12529) );
  AOI21_X1 U14883 ( .B1(n12531), .B2(n12530), .A(n12529), .ZN(n12551) );
  NAND2_X1 U14884 ( .A1(n12533), .A2(n12532), .ZN(n12535) );
  XOR2_X1 U14885 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n12556), .Z(n12557) );
  XNOR2_X1 U14886 ( .A(n12558), .B(n12557), .ZN(n12539) );
  NOR2_X1 U14887 ( .A1(n14982), .A2(n12556), .ZN(n12538) );
  INV_X1 U14888 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14264) );
  OAI21_X1 U14889 ( .B1(n14952), .B2(n14264), .A(n12536), .ZN(n12537) );
  AOI211_X1 U14890 ( .C1(n12539), .C2(n14992), .A(n12538), .B(n12537), .ZN(
        n12550) );
  INV_X1 U14891 ( .A(n12540), .ZN(n12542) );
  AOI21_X1 U14892 ( .B1(n12542), .B2(n6955), .A(n12541), .ZN(n12563) );
  MUX2_X1 U14893 ( .A(n12543), .B(n12867), .S(n11415), .Z(n12545) );
  INV_X1 U14894 ( .A(n12556), .ZN(n12544) );
  NOR2_X1 U14895 ( .A1(n12545), .A2(n12544), .ZN(n12562) );
  INV_X1 U14896 ( .A(n12562), .ZN(n12546) );
  NAND2_X1 U14897 ( .A1(n12545), .A2(n12544), .ZN(n12561) );
  NAND2_X1 U14898 ( .A1(n12546), .A2(n12561), .ZN(n12547) );
  XNOR2_X1 U14899 ( .A(n12563), .B(n12547), .ZN(n12548) );
  NAND2_X1 U14900 ( .A1(n12548), .A2(n14960), .ZN(n12549) );
  OAI211_X1 U14901 ( .C1(n12551), .C2(n14994), .A(n12550), .B(n12549), .ZN(
        P3_U3198) );
  INV_X1 U14902 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12768) );
  NAND2_X1 U14903 ( .A1(n12556), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12552) );
  NAND2_X1 U14904 ( .A1(n12553), .A2(n12552), .ZN(n12554) );
  NAND2_X1 U14905 ( .A1(n12554), .A2(n12575), .ZN(n12584) );
  AOI21_X1 U14906 ( .B1(n12768), .B2(n12555), .A(n12588), .ZN(n12570) );
  XOR2_X1 U14907 ( .A(n12575), .B(n12576), .Z(n12579) );
  XOR2_X1 U14908 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12579), .Z(n12568) );
  AOI21_X1 U14909 ( .B1(n14978), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n12559), 
        .ZN(n12560) );
  OAI21_X1 U14910 ( .B1(n14982), .B2(n12575), .A(n12560), .ZN(n12567) );
  MUX2_X1 U14911 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n11415), .Z(n12572) );
  XNOR2_X1 U14912 ( .A(n12572), .B(n12575), .ZN(n12565) );
  NOR2_X1 U14913 ( .A1(n12564), .A2(n12565), .ZN(n12571) );
  AOI211_X1 U14914 ( .C1(n12565), .C2(n12564), .A(n14986), .B(n12571), .ZN(
        n12566) );
  AOI211_X1 U14915 ( .C1(n14992), .C2(n12568), .A(n12567), .B(n12566), .ZN(
        n12569) );
  OAI21_X1 U14916 ( .B1(n12570), .B2(n14994), .A(n12569), .ZN(P3_U3199) );
  MUX2_X1 U14917 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n11415), .Z(n12574) );
  AOI21_X1 U14918 ( .B1(n12572), .B2(n12575), .A(n12571), .ZN(n12598) );
  XOR2_X1 U14919 ( .A(n12600), .B(n12598), .Z(n12573) );
  NOR2_X1 U14920 ( .A1(n12573), .A2(n12574), .ZN(n12597) );
  AOI21_X1 U14921 ( .B1(n12574), .B2(n12573), .A(n12597), .ZN(n12592) );
  INV_X1 U14922 ( .A(n12575), .ZN(n12577) );
  OAI22_X1 U14923 ( .A1(n12579), .A2(n12578), .B1(n12577), .B2(n12576), .ZN(
        n12602) );
  XOR2_X1 U14924 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n12600), .Z(n12601) );
  XNOR2_X1 U14925 ( .A(n12602), .B(n12601), .ZN(n12583) );
  AOI21_X1 U14926 ( .B1(n14978), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n12580), 
        .ZN(n12581) );
  OAI21_X1 U14927 ( .B1(n14982), .B2(n12600), .A(n12581), .ZN(n12582) );
  AOI21_X1 U14928 ( .B1(n12583), .B2(n14992), .A(n12582), .ZN(n12591) );
  INV_X1 U14929 ( .A(n12584), .ZN(n12587) );
  NAND2_X1 U14930 ( .A1(n12600), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12593) );
  OR2_X1 U14931 ( .A1(n12600), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12585) );
  AND2_X1 U14932 ( .A1(n12593), .A2(n12585), .ZN(n12586) );
  NOR3_X1 U14933 ( .A1(n12588), .A2(n12587), .A3(n12586), .ZN(n12589) );
  OAI21_X1 U14934 ( .B1(n6681), .B2(n12589), .A(n14872), .ZN(n12590) );
  OAI211_X1 U14935 ( .C1(n12592), .C2(n14986), .A(n12591), .B(n12590), .ZN(
        P3_U3200) );
  XNOR2_X1 U14936 ( .A(n12595), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12596) );
  XOR2_X1 U14937 ( .A(n12596), .B(n12594), .Z(n12610) );
  XNOR2_X1 U14938 ( .A(n12595), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12603) );
  MUX2_X1 U14939 ( .A(n12596), .B(n12603), .S(n11415), .Z(n12599) );
  NAND2_X1 U14940 ( .A1(n14978), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12605) );
  OAI211_X1 U14941 ( .C1(n14982), .C2(n12607), .A(n12606), .B(n12605), .ZN(
        n12608) );
  NAND2_X1 U14942 ( .A1(n12611), .A2(n15071), .ZN(n12621) );
  INV_X1 U14943 ( .A(n12612), .ZN(n12613) );
  NAND2_X1 U14944 ( .A1(n12614), .A2(n12613), .ZN(n14348) );
  AOI21_X1 U14945 ( .B1(n12621), .B2(n14348), .A(n15056), .ZN(n12616) );
  AOI21_X1 U14946 ( .B1(n15056), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12616), 
        .ZN(n12615) );
  OAI21_X1 U14947 ( .B1(n14343), .B2(n12818), .A(n12615), .ZN(P3_U3202) );
  AOI21_X1 U14948 ( .B1(n15056), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12616), 
        .ZN(n12617) );
  OAI21_X1 U14949 ( .B1(n12818), .B2(n12618), .A(n12617), .ZN(P3_U3203) );
  INV_X1 U14950 ( .A(n12619), .ZN(n12626) );
  NAND2_X1 U14951 ( .A1(n15056), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n12620) );
  OAI211_X1 U14952 ( .C1(n12622), .C2(n12818), .A(n12621), .B(n12620), .ZN(
        n12623) );
  AOI21_X1 U14953 ( .B1(n12624), .B2(n15074), .A(n12623), .ZN(n12625) );
  OAI21_X1 U14954 ( .B1(n12626), .B2(n12822), .A(n12625), .ZN(P3_U3204) );
  INV_X1 U14955 ( .A(n12627), .ZN(n12629) );
  INV_X1 U14956 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12628) );
  OAI22_X1 U14957 ( .A1(n12629), .A2(n12766), .B1(n15074), .B2(n12628), .ZN(
        n12630) );
  AOI21_X1 U14958 ( .B1(n12631), .B2(n12770), .A(n12630), .ZN(n12634) );
  NAND2_X1 U14959 ( .A1(n12632), .A2(n14340), .ZN(n12633) );
  OAI211_X1 U14960 ( .C1(n12635), .C2(n15056), .A(n12634), .B(n12633), .ZN(
        P3_U3205) );
  INV_X1 U14961 ( .A(n12636), .ZN(n12643) );
  AOI22_X1 U14962 ( .A1(n12637), .A2(n15071), .B1(n15056), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12638) );
  OAI21_X1 U14963 ( .B1(n12639), .B2(n12818), .A(n12638), .ZN(n12640) );
  AOI21_X1 U14964 ( .B1(n12641), .B2(n15072), .A(n12640), .ZN(n12642) );
  OAI21_X1 U14965 ( .B1(n12643), .B2(n15056), .A(n12642), .ZN(P3_U3206) );
  INV_X1 U14966 ( .A(n12644), .ZN(n12650) );
  AOI22_X1 U14967 ( .A1(n15071), .A2(n12645), .B1(n15056), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12646) );
  OAI21_X1 U14968 ( .B1(n12826), .B2(n12818), .A(n12646), .ZN(n12647) );
  AOI21_X1 U14969 ( .B1(n12648), .B2(n15074), .A(n12647), .ZN(n12649) );
  OAI21_X1 U14970 ( .B1(n12822), .B2(n12650), .A(n12649), .ZN(P3_U3207) );
  XNOR2_X1 U14971 ( .A(n12652), .B(n12651), .ZN(n12828) );
  INV_X1 U14972 ( .A(n12828), .ZN(n12663) );
  OAI211_X1 U14973 ( .C1(n12655), .C2(n12654), .A(n12653), .B(n8938), .ZN(
        n12658) );
  AOI22_X1 U14974 ( .A1(n12656), .A2(n15059), .B1(n15062), .B2(n12682), .ZN(
        n12657) );
  NAND2_X1 U14975 ( .A1(n12658), .A2(n12657), .ZN(n12827) );
  AOI22_X1 U14976 ( .A1(n15056), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n15071), 
        .B2(n12659), .ZN(n12660) );
  OAI21_X1 U14977 ( .B1(n12886), .B2(n12818), .A(n12660), .ZN(n12661) );
  AOI21_X1 U14978 ( .B1(n12827), .B2(n15074), .A(n12661), .ZN(n12662) );
  OAI21_X1 U14979 ( .B1(n12663), .B2(n12822), .A(n12662), .ZN(P3_U3208) );
  OAI211_X1 U14980 ( .C1(n12667), .C2(n12666), .A(n12665), .B(n8938), .ZN(
        n12670) );
  NAND2_X1 U14981 ( .A1(n12668), .A2(n15062), .ZN(n12669) );
  OAI211_X1 U14982 ( .C1(n12671), .C2(n15043), .A(n12670), .B(n12669), .ZN(
        n12672) );
  AOI21_X1 U14983 ( .B1(n12832), .B2(n14997), .A(n12672), .ZN(n12834) );
  AOI22_X1 U14984 ( .A1(n15056), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15071), 
        .B2(n12673), .ZN(n12674) );
  OAI21_X1 U14985 ( .B1(n12675), .B2(n12818), .A(n12674), .ZN(n12676) );
  AOI21_X1 U14986 ( .B1(n12832), .B2(n15072), .A(n12676), .ZN(n12677) );
  OAI21_X1 U14987 ( .B1(n12834), .B2(n15056), .A(n12677), .ZN(P3_U3209) );
  OAI211_X1 U14988 ( .C1(n12680), .C2(n12679), .A(n12678), .B(n8938), .ZN(
        n12684) );
  AOI22_X1 U14989 ( .A1(n12682), .A2(n15059), .B1(n15062), .B2(n12681), .ZN(
        n12683) );
  AND2_X1 U14990 ( .A1(n12684), .A2(n12683), .ZN(n12837) );
  INV_X1 U14991 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12687) );
  INV_X1 U14992 ( .A(n12685), .ZN(n12686) );
  OAI22_X1 U14993 ( .A1(n15074), .A2(n12687), .B1(n12686), .B2(n12766), .ZN(
        n12688) );
  AOI21_X1 U14994 ( .B1(n12689), .B2(n12770), .A(n12688), .ZN(n12694) );
  OR2_X1 U14995 ( .A1(n12691), .A2(n12690), .ZN(n12835) );
  NAND3_X1 U14996 ( .A1(n12835), .A2(n12692), .A3(n14340), .ZN(n12693) );
  OAI211_X1 U14997 ( .C1(n12837), .C2(n15056), .A(n12694), .B(n12693), .ZN(
        P3_U3210) );
  XNOR2_X1 U14998 ( .A(n12695), .B(n12697), .ZN(n12840) );
  INV_X1 U14999 ( .A(n12840), .ZN(n12705) );
  XNOR2_X1 U15000 ( .A(n12696), .B(n12697), .ZN(n12698) );
  OAI222_X1 U15001 ( .A1(n15045), .A2(n12700), .B1(n15043), .B2(n12699), .C1(
        n12698), .C2(n15016), .ZN(n12839) );
  AOI22_X1 U15002 ( .A1(n15056), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15071), 
        .B2(n12701), .ZN(n12702) );
  OAI21_X1 U15003 ( .B1(n12892), .B2(n12818), .A(n12702), .ZN(n12703) );
  AOI21_X1 U15004 ( .B1(n12839), .B2(n15074), .A(n12703), .ZN(n12704) );
  OAI21_X1 U15005 ( .B1(n12705), .B2(n12822), .A(n12704), .ZN(P3_U3211) );
  XOR2_X1 U15006 ( .A(n12708), .B(n12706), .Z(n12844) );
  INV_X1 U15007 ( .A(n12844), .ZN(n12716) );
  XOR2_X1 U15008 ( .A(n12708), .B(n12707), .Z(n12709) );
  OAI222_X1 U15009 ( .A1(n15043), .A2(n12711), .B1(n15045), .B2(n12710), .C1(
        n15016), .C2(n12709), .ZN(n12843) );
  AOI22_X1 U15010 ( .A1(n15056), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15071), 
        .B2(n12712), .ZN(n12713) );
  OAI21_X1 U15011 ( .B1(n12896), .B2(n12818), .A(n12713), .ZN(n12714) );
  AOI21_X1 U15012 ( .B1(n12843), .B2(n15074), .A(n12714), .ZN(n12715) );
  OAI21_X1 U15013 ( .B1(n12822), .B2(n12716), .A(n12715), .ZN(P3_U3212) );
  OAI21_X1 U15014 ( .B1(n7546), .B2(n8102), .A(n12717), .ZN(n12851) );
  OAI211_X1 U15015 ( .C1(n12720), .C2(n12719), .A(n12718), .B(n8938), .ZN(
        n12724) );
  AOI22_X1 U15016 ( .A1(n15059), .A2(n12722), .B1(n12721), .B2(n15062), .ZN(
        n12723) );
  NAND2_X1 U15017 ( .A1(n12724), .A2(n12723), .ZN(n12847) );
  AOI22_X1 U15018 ( .A1(n15056), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15071), 
        .B2(n12725), .ZN(n12726) );
  OAI21_X1 U15019 ( .B1(n12727), .B2(n12818), .A(n12726), .ZN(n12728) );
  AOI21_X1 U15020 ( .B1(n12847), .B2(n15074), .A(n12728), .ZN(n12729) );
  OAI21_X1 U15021 ( .B1(n12851), .B2(n12822), .A(n12729), .ZN(P3_U3213) );
  XOR2_X1 U15022 ( .A(n12731), .B(n12730), .Z(n12853) );
  INV_X1 U15023 ( .A(n12853), .ZN(n12741) );
  OAI211_X1 U15024 ( .C1(n6750), .C2(n7461), .A(n8938), .B(n12732), .ZN(n12736) );
  AOI22_X1 U15025 ( .A1(n15062), .A2(n12734), .B1(n12733), .B2(n15059), .ZN(
        n12735) );
  NAND2_X1 U15026 ( .A1(n12736), .A2(n12735), .ZN(n12852) );
  AOI22_X1 U15027 ( .A1(n15056), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15071), 
        .B2(n12737), .ZN(n12738) );
  OAI21_X1 U15028 ( .B1(n12901), .B2(n12818), .A(n12738), .ZN(n12739) );
  AOI21_X1 U15029 ( .B1(n12852), .B2(n15074), .A(n12739), .ZN(n12740) );
  OAI21_X1 U15030 ( .B1(n12741), .B2(n12822), .A(n12740), .ZN(P3_U3214) );
  INV_X1 U15031 ( .A(n12742), .ZN(n12743) );
  AOI21_X1 U15032 ( .B1(n7900), .B2(n12744), .A(n12743), .ZN(n12857) );
  INV_X1 U15033 ( .A(n12857), .ZN(n12756) );
  INV_X1 U15034 ( .A(n12745), .ZN(n12746) );
  AOI21_X1 U15035 ( .B1(n12748), .B2(n12747), .A(n12746), .ZN(n12749) );
  OAI222_X1 U15036 ( .A1(n15043), .A2(n12750), .B1(n15045), .B2(n12778), .C1(
        n15016), .C2(n12749), .ZN(n12856) );
  INV_X1 U15037 ( .A(n12751), .ZN(n12905) );
  AOI22_X1 U15038 ( .A1(n15056), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15071), 
        .B2(n12752), .ZN(n12753) );
  OAI21_X1 U15039 ( .B1(n12905), .B2(n12818), .A(n12753), .ZN(n12754) );
  AOI21_X1 U15040 ( .B1(n12856), .B2(n15074), .A(n12754), .ZN(n12755) );
  OAI21_X1 U15041 ( .B1(n12822), .B2(n12756), .A(n12755), .ZN(P3_U3215) );
  AOI21_X1 U15042 ( .B1(n12757), .B2(n12763), .A(n15016), .ZN(n12761) );
  OAI22_X1 U15043 ( .A1(n12792), .A2(n15045), .B1(n12758), .B2(n15043), .ZN(
        n12759) );
  AOI21_X1 U15044 ( .B1(n12761), .B2(n12760), .A(n12759), .ZN(n12862) );
  OAI21_X1 U15045 ( .B1(n12764), .B2(n12763), .A(n12762), .ZN(n12861) );
  NAND2_X1 U15046 ( .A1(n12861), .A2(n14340), .ZN(n12772) );
  INV_X1 U15047 ( .A(n12765), .ZN(n12767) );
  OAI22_X1 U15048 ( .A1(n15074), .A2(n12768), .B1(n12767), .B2(n12766), .ZN(
        n12769) );
  AOI21_X1 U15049 ( .B1(n12860), .B2(n12770), .A(n12769), .ZN(n12771) );
  OAI211_X1 U15050 ( .C1(n15056), .C2(n12862), .A(n12772), .B(n12771), .ZN(
        P3_U3216) );
  OAI21_X1 U15051 ( .B1(n12774), .B2(n12776), .A(n12773), .ZN(n12866) );
  INV_X1 U15052 ( .A(n12866), .ZN(n12784) );
  XOR2_X1 U15053 ( .A(n12776), .B(n12775), .Z(n12777) );
  OAI222_X1 U15054 ( .A1(n15043), .A2(n12778), .B1(n15045), .B2(n12802), .C1(
        n12777), .C2(n15016), .ZN(n12865) );
  INV_X1 U15055 ( .A(n12779), .ZN(n12910) );
  AOI22_X1 U15056 ( .A1(n15056), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15071), 
        .B2(n12780), .ZN(n12781) );
  OAI21_X1 U15057 ( .B1(n12910), .B2(n12818), .A(n12781), .ZN(n12782) );
  AOI21_X1 U15058 ( .B1(n12865), .B2(n15074), .A(n12782), .ZN(n12783) );
  OAI21_X1 U15059 ( .B1(n12784), .B2(n12822), .A(n12783), .ZN(P3_U3217) );
  NAND2_X1 U15060 ( .A1(n12786), .A2(n12785), .ZN(n12788) );
  XNOR2_X1 U15061 ( .A(n12788), .B(n12787), .ZN(n12870) );
  INV_X1 U15062 ( .A(n12870), .ZN(n12797) );
  XNOR2_X1 U15063 ( .A(n12789), .B(n12790), .ZN(n12791) );
  OAI222_X1 U15064 ( .A1(n15043), .A2(n12792), .B1(n15045), .B2(n12815), .C1(
        n15016), .C2(n12791), .ZN(n12869) );
  AOI22_X1 U15065 ( .A1(n15056), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15071), 
        .B2(n12793), .ZN(n12794) );
  OAI21_X1 U15066 ( .B1(n12914), .B2(n12818), .A(n12794), .ZN(n12795) );
  AOI21_X1 U15067 ( .B1(n12869), .B2(n15074), .A(n12795), .ZN(n12796) );
  OAI21_X1 U15068 ( .B1(n12797), .B2(n12822), .A(n12796), .ZN(P3_U3218) );
  XNOR2_X1 U15069 ( .A(n12798), .B(n12800), .ZN(n12873) );
  INV_X1 U15070 ( .A(n12873), .ZN(n12808) );
  XNOR2_X1 U15071 ( .A(n12799), .B(n12800), .ZN(n12801) );
  OAI222_X1 U15072 ( .A1(n15045), .A2(n12803), .B1(n15043), .B2(n12802), .C1(
        n12801), .C2(n15016), .ZN(n12872) );
  AOI22_X1 U15073 ( .A1(n15056), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15071), 
        .B2(n12804), .ZN(n12805) );
  OAI21_X1 U15074 ( .B1(n12818), .B2(n12918), .A(n12805), .ZN(n12806) );
  AOI21_X1 U15075 ( .B1(n12872), .B2(n15074), .A(n12806), .ZN(n12807) );
  OAI21_X1 U15076 ( .B1(n12808), .B2(n12822), .A(n12807), .ZN(P3_U3219) );
  XNOR2_X1 U15077 ( .A(n12810), .B(n12809), .ZN(n12877) );
  INV_X1 U15078 ( .A(n12877), .ZN(n12821) );
  XNOR2_X1 U15079 ( .A(n12811), .B(n12812), .ZN(n12813) );
  OAI222_X1 U15080 ( .A1(n15043), .A2(n12815), .B1(n15045), .B2(n12814), .C1(
        n12813), .C2(n15016), .ZN(n12876) );
  AOI22_X1 U15081 ( .A1(n15056), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n15071), 
        .B2(n12816), .ZN(n12817) );
  OAI21_X1 U15082 ( .B1(n12818), .B2(n12922), .A(n12817), .ZN(n12819) );
  AOI21_X1 U15083 ( .B1(n12876), .B2(n15074), .A(n12819), .ZN(n12820) );
  OAI21_X1 U15084 ( .B1(n12822), .B2(n12821), .A(n12820), .ZN(P3_U3220) );
  INV_X1 U15085 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12824) );
  OAI21_X1 U15086 ( .B1(n12826), .B2(n12882), .A(n12825), .ZN(P3_U3485) );
  INV_X1 U15087 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12829) );
  AOI21_X1 U15088 ( .B1(n12828), .B2(n15101), .A(n12827), .ZN(n12883) );
  MUX2_X1 U15089 ( .A(n12829), .B(n12883), .S(n15132), .Z(n12830) );
  OAI21_X1 U15090 ( .B1(n12886), .B2(n12882), .A(n12830), .ZN(P3_U3484) );
  AOI22_X1 U15091 ( .A1(n12832), .A2(n15115), .B1(n14345), .B2(n12831), .ZN(
        n12833) );
  NAND2_X1 U15092 ( .A1(n12834), .A2(n12833), .ZN(n12887) );
  MUX2_X1 U15093 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n12887), .S(n15132), .Z(
        P3_U3483) );
  NAND3_X1 U15094 ( .A1(n12835), .A2(n12692), .A3(n15101), .ZN(n12836) );
  OAI211_X1 U15095 ( .C1(n12838), .C2(n15103), .A(n12837), .B(n12836), .ZN(
        n12888) );
  MUX2_X1 U15096 ( .A(n12888), .B(P3_REG1_REG_23__SCAN_IN), .S(n15130), .Z(
        P3_U3482) );
  AOI21_X1 U15097 ( .B1(n15101), .B2(n12840), .A(n12839), .ZN(n12889) );
  MUX2_X1 U15098 ( .A(n12841), .B(n12889), .S(n15132), .Z(n12842) );
  OAI21_X1 U15099 ( .B1(n12892), .B2(n12882), .A(n12842), .ZN(P3_U3481) );
  AOI21_X1 U15100 ( .B1(n12844), .B2(n15101), .A(n12843), .ZN(n12893) );
  MUX2_X1 U15101 ( .A(n12845), .B(n12893), .S(n15132), .Z(n12846) );
  OAI21_X1 U15102 ( .B1(n12896), .B2(n12882), .A(n12846), .ZN(P3_U3480) );
  INV_X1 U15103 ( .A(n15101), .ZN(n12850) );
  AOI21_X1 U15104 ( .B1(n14345), .B2(n12848), .A(n12847), .ZN(n12849) );
  OAI21_X1 U15105 ( .B1(n12851), .B2(n12850), .A(n12849), .ZN(n12897) );
  MUX2_X1 U15106 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n12897), .S(n15132), .Z(
        P3_U3479) );
  AOI21_X1 U15107 ( .B1(n12853), .B2(n15101), .A(n12852), .ZN(n12898) );
  MUX2_X1 U15108 ( .A(n12854), .B(n12898), .S(n15132), .Z(n12855) );
  OAI21_X1 U15109 ( .B1(n12882), .B2(n12901), .A(n12855), .ZN(P3_U3478) );
  AOI21_X1 U15110 ( .B1(n12857), .B2(n15101), .A(n12856), .ZN(n12902) );
  MUX2_X1 U15111 ( .A(n12858), .B(n12902), .S(n15132), .Z(n12859) );
  OAI21_X1 U15112 ( .B1(n12905), .B2(n12882), .A(n12859), .ZN(P3_U3477) );
  INV_X1 U15113 ( .A(n12860), .ZN(n12864) );
  NAND2_X1 U15114 ( .A1(n12861), .A2(n15101), .ZN(n12863) );
  OAI211_X1 U15115 ( .C1(n12864), .C2(n15103), .A(n12863), .B(n12862), .ZN(
        n12906) );
  MUX2_X1 U15116 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12906), .S(n15132), .Z(
        P3_U3476) );
  AOI21_X1 U15117 ( .B1(n15101), .B2(n12866), .A(n12865), .ZN(n12907) );
  MUX2_X1 U15118 ( .A(n12867), .B(n12907), .S(n15132), .Z(n12868) );
  OAI21_X1 U15119 ( .B1(n12910), .B2(n12882), .A(n12868), .ZN(P3_U3475) );
  AOI21_X1 U15120 ( .B1(n15101), .B2(n12870), .A(n12869), .ZN(n12911) );
  MUX2_X1 U15121 ( .A(n15344), .B(n12911), .S(n15132), .Z(n12871) );
  OAI21_X1 U15122 ( .B1(n12914), .B2(n12882), .A(n12871), .ZN(P3_U3474) );
  AOI21_X1 U15123 ( .B1(n15101), .B2(n12873), .A(n12872), .ZN(n12915) );
  MUX2_X1 U15124 ( .A(n12874), .B(n12915), .S(n15132), .Z(n12875) );
  OAI21_X1 U15125 ( .B1(n12882), .B2(n12918), .A(n12875), .ZN(P3_U3473) );
  AOI21_X1 U15126 ( .B1(n12877), .B2(n15101), .A(n12876), .ZN(n12919) );
  MUX2_X1 U15127 ( .A(n7791), .B(n12919), .S(n15132), .Z(n12878) );
  OAI21_X1 U15128 ( .B1(n12882), .B2(n12922), .A(n12878), .ZN(P3_U3472) );
  AOI21_X1 U15129 ( .B1(n15101), .B2(n12880), .A(n12879), .ZN(n12923) );
  MUX2_X1 U15130 ( .A(n7747), .B(n12923), .S(n15132), .Z(n12881) );
  OAI21_X1 U15131 ( .B1(n12882), .B2(n12925), .A(n12881), .ZN(P3_U3470) );
  INV_X1 U15132 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12884) );
  MUX2_X1 U15133 ( .A(n12884), .B(n12883), .S(n15119), .Z(n12885) );
  OAI21_X1 U15134 ( .B1(n12886), .B2(n12926), .A(n12885), .ZN(P3_U3452) );
  MUX2_X1 U15135 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n12887), .S(n15119), .Z(
        P3_U3451) );
  MUX2_X1 U15136 ( .A(n12888), .B(P3_REG0_REG_23__SCAN_IN), .S(n8156), .Z(
        P3_U3450) );
  INV_X1 U15137 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12890) );
  MUX2_X1 U15138 ( .A(n12890), .B(n12889), .S(n15119), .Z(n12891) );
  OAI21_X1 U15139 ( .B1(n12892), .B2(n12926), .A(n12891), .ZN(P3_U3449) );
  INV_X1 U15140 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12894) );
  MUX2_X1 U15141 ( .A(n12894), .B(n12893), .S(n15119), .Z(n12895) );
  OAI21_X1 U15142 ( .B1(n12896), .B2(n12926), .A(n12895), .ZN(P3_U3448) );
  MUX2_X1 U15143 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n12897), .S(n15119), .Z(
        P3_U3447) );
  INV_X1 U15144 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12899) );
  MUX2_X1 U15145 ( .A(n12899), .B(n12898), .S(n15119), .Z(n12900) );
  OAI21_X1 U15146 ( .B1(n12926), .B2(n12901), .A(n12900), .ZN(P3_U3446) );
  INV_X1 U15147 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12903) );
  MUX2_X1 U15148 ( .A(n12903), .B(n12902), .S(n15119), .Z(n12904) );
  OAI21_X1 U15149 ( .B1(n12905), .B2(n12926), .A(n12904), .ZN(P3_U3444) );
  MUX2_X1 U15150 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n12906), .S(n15119), .Z(
        P3_U3441) );
  INV_X1 U15151 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12908) );
  MUX2_X1 U15152 ( .A(n12908), .B(n12907), .S(n15119), .Z(n12909) );
  OAI21_X1 U15153 ( .B1(n12910), .B2(n12926), .A(n12909), .ZN(P3_U3438) );
  INV_X1 U15154 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12912) );
  MUX2_X1 U15155 ( .A(n12912), .B(n12911), .S(n15119), .Z(n12913) );
  OAI21_X1 U15156 ( .B1(n12914), .B2(n12926), .A(n12913), .ZN(P3_U3435) );
  INV_X1 U15157 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12916) );
  MUX2_X1 U15158 ( .A(n12916), .B(n12915), .S(n15119), .Z(n12917) );
  OAI21_X1 U15159 ( .B1(n12926), .B2(n12918), .A(n12917), .ZN(P3_U3432) );
  INV_X1 U15160 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n12920) );
  MUX2_X1 U15161 ( .A(n12920), .B(n12919), .S(n15119), .Z(n12921) );
  OAI21_X1 U15162 ( .B1(n12926), .B2(n12922), .A(n12921), .ZN(P3_U3429) );
  INV_X1 U15163 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n15209) );
  MUX2_X1 U15164 ( .A(n15209), .B(n12923), .S(n15119), .Z(n12924) );
  OAI21_X1 U15165 ( .B1(n12926), .B2(n12925), .A(n12924), .ZN(P3_U3423) );
  INV_X1 U15166 ( .A(n12927), .ZN(n12931) );
  INV_X1 U15167 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n12928) );
  NAND3_X1 U15168 ( .A1(n12928), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n12930) );
  OAI22_X1 U15169 ( .A1(n12931), .A2(n12930), .B1(n12929), .B2(n12944), .ZN(
        n12932) );
  AOI21_X1 U15170 ( .B1(n12934), .B2(n12933), .A(n12932), .ZN(n12935) );
  INV_X1 U15171 ( .A(n12935), .ZN(P3_U3264) );
  INV_X1 U15172 ( .A(n12936), .ZN(n12937) );
  OAI222_X1 U15173 ( .A1(n12944), .A2(n12939), .B1(P3_U3151), .B2(n12938), 
        .C1(n11943), .C2(n12937), .ZN(P3_U3266) );
  INV_X1 U15174 ( .A(n12940), .ZN(n12941) );
  OAI222_X1 U15175 ( .A1(n12944), .A2(n12942), .B1(P3_U3151), .B2(n6628), .C1(
        n11943), .C2(n12941), .ZN(P3_U3267) );
  INV_X1 U15176 ( .A(n12943), .ZN(n12946) );
  OAI222_X1 U15177 ( .A1(P3_U3151), .A2(n11415), .B1(n11943), .B2(n12946), 
        .C1(n12945), .C2(n12944), .ZN(P3_U3268) );
  AOI21_X1 U15178 ( .B1(n12949), .B2(n12948), .A(n13083), .ZN(n12954) );
  NAND2_X1 U15179 ( .A1(n13189), .A2(n13081), .ZN(n12953) );
  AOI22_X1 U15180 ( .A1(n13087), .A2(n13076), .B1(n13075), .B2(n13089), .ZN(
        n13183) );
  AOI22_X1 U15181 ( .A1(n13188), .A2(n13077), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12950) );
  OAI21_X1 U15182 ( .B1(n13183), .B2(n13079), .A(n12950), .ZN(n12951) );
  OAI211_X1 U15183 ( .C1(n12957), .C2(n12956), .A(n12955), .B(n13049), .ZN(
        n12963) );
  NAND2_X1 U15184 ( .A1(n13091), .A2(n13076), .ZN(n12959) );
  NAND2_X1 U15185 ( .A1(n12977), .A2(n13075), .ZN(n12958) );
  NAND2_X1 U15186 ( .A1(n12959), .A2(n12958), .ZN(n13403) );
  OAI22_X1 U15187 ( .A1(n13244), .A2(n13067), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12960), .ZN(n12961) );
  AOI21_X1 U15188 ( .B1(n13403), .B2(n13065), .A(n12961), .ZN(n12962) );
  OAI211_X1 U15189 ( .C1(n13248), .C2(n8914), .A(n12963), .B(n12962), .ZN(
        P2_U3188) );
  INV_X1 U15190 ( .A(n12964), .ZN(n12965) );
  AOI21_X1 U15191 ( .B1(n12967), .B2(n12966), .A(n12965), .ZN(n12973) );
  OAI22_X1 U15192 ( .A1(n12969), .A2(n13042), .B1(n12968), .B2(n13060), .ZN(
        n13424) );
  NAND2_X1 U15193 ( .A1(n13424), .A2(n13065), .ZN(n12970) );
  NAND2_X1 U15194 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13147)
         );
  OAI211_X1 U15195 ( .C1(n13067), .C2(n13305), .A(n12970), .B(n13147), .ZN(
        n12971) );
  AOI21_X1 U15196 ( .B1(n13425), .B2(n13081), .A(n12971), .ZN(n12972) );
  OAI21_X1 U15197 ( .B1(n12973), .B2(n13083), .A(n12972), .ZN(P2_U3191) );
  OAI211_X1 U15198 ( .C1(n12976), .C2(n12975), .A(n12974), .B(n13049), .ZN(
        n12983) );
  AOI22_X1 U15199 ( .A1(n12977), .A2(n13076), .B1(n13075), .B2(n13094), .ZN(
        n13272) );
  INV_X1 U15200 ( .A(n13272), .ZN(n12981) );
  INV_X1 U15201 ( .A(n13276), .ZN(n12979) );
  OAI22_X1 U15202 ( .A1(n13067), .A2(n12979), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12978), .ZN(n12980) );
  AOI21_X1 U15203 ( .B1(n12981), .B2(n13065), .A(n12980), .ZN(n12982) );
  OAI211_X1 U15204 ( .C1(n13279), .C2(n8914), .A(n12983), .B(n12982), .ZN(
        P2_U3195) );
  OAI211_X1 U15205 ( .C1(n12986), .C2(n12985), .A(n12984), .B(n13049), .ZN(
        n12992) );
  OAI22_X1 U15206 ( .A1(n12988), .A2(n13042), .B1(n12987), .B2(n13060), .ZN(
        n13211) );
  OAI22_X1 U15207 ( .A1(n13214), .A2(n13067), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12989), .ZN(n12990) );
  AOI21_X1 U15208 ( .B1(n13211), .B2(n13065), .A(n12990), .ZN(n12991) );
  OAI211_X1 U15209 ( .C1(n13217), .C2(n8914), .A(n12992), .B(n12991), .ZN(
        P2_U3197) );
  INV_X1 U15210 ( .A(n11798), .ZN(n12994) );
  AOI22_X1 U15211 ( .A1(n12996), .A2(n12995), .B1(n12994), .B2(n12993), .ZN(
        n12999) );
  OAI21_X1 U15212 ( .B1(n12999), .B2(n12998), .A(n12997), .ZN(n13000) );
  NAND2_X1 U15213 ( .A1(n13000), .A2(n13049), .ZN(n13007) );
  INV_X1 U15214 ( .A(n13355), .ZN(n13005) );
  OR2_X1 U15215 ( .A1(n13061), .A2(n13042), .ZN(n13002) );
  NAND2_X1 U15216 ( .A1(n13099), .A2(n13075), .ZN(n13001) );
  AND2_X1 U15217 ( .A1(n13002), .A2(n13001), .ZN(n13352) );
  OAI22_X1 U15218 ( .A1(n13079), .A2(n13352), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13003), .ZN(n13004) );
  AOI21_X1 U15219 ( .B1(n13005), .B2(n13077), .A(n13004), .ZN(n13006) );
  OAI211_X1 U15220 ( .C1(n13008), .C2(n8914), .A(n13007), .B(n13006), .ZN(
        P2_U3198) );
  OAI21_X1 U15221 ( .B1(n13011), .B2(n13010), .A(n13009), .ZN(n13012) );
  NAND2_X1 U15222 ( .A1(n13012), .A2(n13049), .ZN(n13015) );
  AOI22_X1 U15223 ( .A1(n13096), .A2(n13076), .B1(n13075), .B2(n13098), .ZN(
        n13331) );
  NAND2_X1 U15224 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n14739)
         );
  OAI21_X1 U15225 ( .B1(n13331), .B2(n13079), .A(n14739), .ZN(n13013) );
  AOI21_X1 U15226 ( .B1(n13339), .B2(n13077), .A(n13013), .ZN(n13014) );
  OAI211_X1 U15227 ( .C1(n13342), .C2(n8914), .A(n13015), .B(n13014), .ZN(
        P2_U3200) );
  OAI211_X1 U15228 ( .C1(n13018), .C2(n13017), .A(n13016), .B(n13049), .ZN(
        n13025) );
  INV_X1 U15229 ( .A(n13090), .ZN(n13020) );
  OAI22_X1 U15230 ( .A1(n13020), .A2(n13042), .B1(n13019), .B2(n13060), .ZN(
        n13224) );
  INV_X1 U15231 ( .A(n13233), .ZN(n13022) );
  OAI22_X1 U15232 ( .A1(n13022), .A2(n13067), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13021), .ZN(n13023) );
  AOI21_X1 U15233 ( .B1(n13224), .B2(n13065), .A(n13023), .ZN(n13024) );
  OAI211_X1 U15234 ( .C1(n13235), .C2(n8914), .A(n13025), .B(n13024), .ZN(
        P2_U3201) );
  OAI21_X1 U15235 ( .B1(n13026), .B2(n13028), .A(n13027), .ZN(n13029) );
  NAND2_X1 U15236 ( .A1(n13029), .A2(n13049), .ZN(n13035) );
  AOI22_X1 U15237 ( .A1(n13081), .A2(n13031), .B1(n13077), .B2(n13030), .ZN(
        n13034) );
  NAND2_X1 U15238 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n13129) );
  NAND2_X1 U15239 ( .A1(n13065), .A2(n13032), .ZN(n13033) );
  NAND4_X1 U15240 ( .A1(n13035), .A2(n13034), .A3(n13129), .A4(n13033), .ZN(
        P2_U3202) );
  NAND2_X1 U15241 ( .A1(n13038), .A2(n13037), .ZN(n13039) );
  XOR2_X1 U15242 ( .A(n13040), .B(n13039), .Z(n13048) );
  OAI22_X1 U15243 ( .A1(n13043), .A2(n13042), .B1(n13041), .B2(n13060), .ZN(
        n13286) );
  OAI22_X1 U15244 ( .A1(n13067), .A2(n13290), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13044), .ZN(n13046) );
  NOR2_X1 U15245 ( .A1(n13294), .A2(n8914), .ZN(n13045) );
  AOI211_X1 U15246 ( .C1(n13065), .C2(n13286), .A(n13046), .B(n13045), .ZN(
        n13047) );
  OAI21_X1 U15247 ( .B1(n13048), .B2(n13083), .A(n13047), .ZN(P2_U3205) );
  OAI211_X1 U15248 ( .C1(n13052), .C2(n13051), .A(n13050), .B(n13049), .ZN(
        n13057) );
  AOI22_X1 U15249 ( .A1(n13092), .A2(n13076), .B1(n13075), .B2(n13093), .ZN(
        n13256) );
  INV_X1 U15250 ( .A(n13256), .ZN(n13055) );
  OAI22_X1 U15251 ( .A1(n13260), .A2(n13067), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13053), .ZN(n13054) );
  AOI21_X1 U15252 ( .B1(n13055), .B2(n13065), .A(n13054), .ZN(n13056) );
  OAI211_X1 U15253 ( .C1(n13264), .C2(n8914), .A(n13057), .B(n13056), .ZN(
        P2_U3207) );
  XNOR2_X1 U15254 ( .A(n13058), .B(n13059), .ZN(n13070) );
  NAND2_X1 U15255 ( .A1(n13095), .A2(n13076), .ZN(n13063) );
  OR2_X1 U15256 ( .A1(n13061), .A2(n13060), .ZN(n13062) );
  NAND2_X1 U15257 ( .A1(n13063), .A2(n13062), .ZN(n13430) );
  AOI21_X1 U15258 ( .B1(n13065), .B2(n13430), .A(n13064), .ZN(n13066) );
  OAI21_X1 U15259 ( .B1(n13318), .B2(n13067), .A(n13066), .ZN(n13068) );
  AOI21_X1 U15260 ( .B1(n13431), .B2(n13081), .A(n13068), .ZN(n13069) );
  OAI21_X1 U15261 ( .B1(n13070), .B2(n13083), .A(n13069), .ZN(P2_U3210) );
  INV_X1 U15262 ( .A(n13071), .ZN(n13072) );
  AOI21_X1 U15263 ( .B1(n13074), .B2(n13073), .A(n13072), .ZN(n13084) );
  AOI22_X1 U15264 ( .A1(n13088), .A2(n13076), .B1(n13075), .B2(n13090), .ZN(
        n13196) );
  AOI22_X1 U15265 ( .A1(n13202), .A2(n13077), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13078) );
  OAI21_X1 U15266 ( .B1(n13196), .B2(n13079), .A(n13078), .ZN(n13080) );
  AOI21_X1 U15267 ( .B1(n13388), .B2(n13081), .A(n13080), .ZN(n13082) );
  OAI21_X1 U15268 ( .B1(n13084), .B2(n13083), .A(n13082), .ZN(P2_U3212) );
  MUX2_X1 U15269 ( .A(n13152), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13113), .Z(
        P2_U3562) );
  MUX2_X1 U15270 ( .A(n13085), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13113), .Z(
        P2_U3561) );
  MUX2_X1 U15271 ( .A(n13086), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13113), .Z(
        P2_U3560) );
  MUX2_X1 U15272 ( .A(n13087), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13113), .Z(
        P2_U3559) );
  MUX2_X1 U15273 ( .A(n13088), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13113), .Z(
        P2_U3558) );
  MUX2_X1 U15274 ( .A(n13089), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13113), .Z(
        P2_U3557) );
  MUX2_X1 U15275 ( .A(n13090), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13113), .Z(
        P2_U3556) );
  MUX2_X1 U15276 ( .A(n13091), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13113), .Z(
        P2_U3555) );
  MUX2_X1 U15277 ( .A(n13092), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13113), .Z(
        P2_U3554) );
  MUX2_X1 U15278 ( .A(n13093), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13113), .Z(
        P2_U3552) );
  MUX2_X1 U15279 ( .A(n13094), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13113), .Z(
        P2_U3551) );
  MUX2_X1 U15280 ( .A(n13095), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13113), .Z(
        P2_U3550) );
  MUX2_X1 U15281 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13096), .S(P2_U3947), .Z(
        P2_U3549) );
  MUX2_X1 U15282 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13097), .S(P2_U3947), .Z(
        P2_U3548) );
  MUX2_X1 U15283 ( .A(n13098), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13113), .Z(
        P2_U3547) );
  MUX2_X1 U15284 ( .A(n13099), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13113), .Z(
        P2_U3546) );
  MUX2_X1 U15285 ( .A(n13100), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13113), .Z(
        P2_U3545) );
  MUX2_X1 U15286 ( .A(n13101), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13113), .Z(
        P2_U3544) );
  MUX2_X1 U15287 ( .A(n13102), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13113), .Z(
        P2_U3543) );
  MUX2_X1 U15288 ( .A(n13103), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13113), .Z(
        P2_U3542) );
  MUX2_X1 U15289 ( .A(n13104), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13113), .Z(
        P2_U3541) );
  MUX2_X1 U15290 ( .A(n13105), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13113), .Z(
        P2_U3540) );
  MUX2_X1 U15291 ( .A(n13106), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13113), .Z(
        P2_U3539) );
  MUX2_X1 U15292 ( .A(n13107), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13113), .Z(
        P2_U3538) );
  MUX2_X1 U15293 ( .A(n13108), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13113), .Z(
        P2_U3537) );
  MUX2_X1 U15294 ( .A(n13109), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13113), .Z(
        P2_U3536) );
  MUX2_X1 U15295 ( .A(n13110), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13113), .Z(
        P2_U3535) );
  MUX2_X1 U15296 ( .A(n7497), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13113), .Z(
        P2_U3534) );
  MUX2_X1 U15297 ( .A(n13111), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13113), .Z(
        P2_U3533) );
  MUX2_X1 U15298 ( .A(n13112), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13113), .Z(
        P2_U3532) );
  MUX2_X1 U15299 ( .A(n13114), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13113), .Z(
        P2_U3531) );
  MUX2_X1 U15300 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10224), .S(n13115), .Z(
        n13117) );
  NAND3_X1 U15301 ( .A1(n13117), .A2(n14680), .A3(n13116), .ZN(n13118) );
  AND3_X1 U15302 ( .A1(n14752), .A2(n13119), .A3(n13118), .ZN(n13120) );
  AOI21_X1 U15303 ( .B1(n14750), .B2(n13121), .A(n13120), .ZN(n13130) );
  NAND2_X1 U15304 ( .A1(n14726), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n13128) );
  INV_X1 U15305 ( .A(n13122), .ZN(n13126) );
  NAND3_X1 U15306 ( .A1(n14683), .A2(n13124), .A3(n13123), .ZN(n13125) );
  NAND3_X1 U15307 ( .A1(n14729), .A2(n13126), .A3(n13125), .ZN(n13127) );
  NAND4_X1 U15308 ( .A1(n13130), .A2(n13129), .A3(n13128), .A4(n13127), .ZN(
        P2_U3218) );
  INV_X1 U15309 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n13149) );
  NOR2_X1 U15310 ( .A1(n13136), .A2(n13131), .ZN(n13132) );
  NOR2_X1 U15311 ( .A1(n13133), .A2(n13132), .ZN(n13134) );
  XOR2_X1 U15312 ( .A(n13134), .B(P2_REG2_REG_19__SCAN_IN), .Z(n13144) );
  INV_X1 U15313 ( .A(n13144), .ZN(n13142) );
  NAND2_X1 U15314 ( .A1(n13136), .A2(n13135), .ZN(n13137) );
  NAND2_X1 U15315 ( .A1(n13138), .A2(n13137), .ZN(n13140) );
  XNOR2_X1 U15316 ( .A(n13140), .B(n13139), .ZN(n13143) );
  OAI21_X1 U15317 ( .B1(n13143), .B2(n14718), .A(n14722), .ZN(n13141) );
  AOI21_X1 U15318 ( .B1(n13142), .B2(n14729), .A(n13141), .ZN(n13146) );
  AOI22_X1 U15319 ( .A1(n13144), .A2(n14729), .B1(n14752), .B2(n13143), .ZN(
        n13145) );
  MUX2_X1 U15320 ( .A(n13146), .B(n13145), .S(n8904), .Z(n13148) );
  OAI211_X1 U15321 ( .C1(n13149), .C2(n14741), .A(n13148), .B(n13147), .ZN(
        P2_U3233) );
  XNOR2_X1 U15322 ( .A(n13157), .B(n13370), .ZN(n13150) );
  NAND2_X1 U15323 ( .A1(n13150), .A2(n13359), .ZN(n13371) );
  NOR2_X1 U15324 ( .A1(n13357), .A2(n13151), .ZN(n13154) );
  NAND2_X1 U15325 ( .A1(n13153), .A2(n13152), .ZN(n13373) );
  NOR2_X1 U15326 ( .A1(n14761), .A2(n13373), .ZN(n13160) );
  AOI211_X1 U15327 ( .C1(n13370), .C2(n13366), .A(n13154), .B(n13160), .ZN(
        n13155) );
  OAI21_X1 U15328 ( .B1(n13371), .B2(n13363), .A(n13155), .ZN(P2_U3234) );
  INV_X1 U15329 ( .A(n13161), .ZN(n13375) );
  INV_X1 U15330 ( .A(n13156), .ZN(n13159) );
  INV_X1 U15331 ( .A(n13157), .ZN(n13158) );
  OAI211_X1 U15332 ( .C1(n13375), .C2(n13159), .A(n13158), .B(n13359), .ZN(
        n13374) );
  AOI21_X1 U15333 ( .B1(n14761), .B2(P2_REG2_REG_30__SCAN_IN), .A(n13160), 
        .ZN(n13163) );
  NAND2_X1 U15334 ( .A1(n13161), .A2(n13366), .ZN(n13162) );
  OAI211_X1 U15335 ( .C1(n13374), .C2(n13363), .A(n13163), .B(n13162), .ZN(
        P2_U3235) );
  AOI211_X1 U15336 ( .C1(n13171), .C2(n13165), .A(n13332), .B(n13164), .ZN(
        n13168) );
  INV_X1 U15337 ( .A(n13166), .ZN(n13167) );
  OAI21_X1 U15338 ( .B1(n13171), .B2(n13170), .A(n13169), .ZN(n13380) );
  OAI22_X1 U15339 ( .A1(n13173), .A2(n13354), .B1(n13172), .B2(n13357), .ZN(
        n13174) );
  AOI21_X1 U15340 ( .B1(n13377), .B2(n13366), .A(n13174), .ZN(n13179) );
  NAND2_X1 U15341 ( .A1(n13377), .A2(n6651), .ZN(n13175) );
  NAND2_X1 U15342 ( .A1(n13175), .A2(n13359), .ZN(n13176) );
  NOR2_X1 U15343 ( .A1(n13177), .A2(n13176), .ZN(n13376) );
  NAND2_X1 U15344 ( .A1(n13376), .A2(n13338), .ZN(n13178) );
  OAI211_X1 U15345 ( .C1(n13380), .C2(n13369), .A(n13179), .B(n13178), .ZN(
        n13180) );
  INV_X1 U15346 ( .A(n13180), .ZN(n13181) );
  OAI21_X1 U15347 ( .B1(n13379), .B2(n14761), .A(n13181), .ZN(P2_U3237) );
  XOR2_X1 U15348 ( .A(n13182), .B(n13186), .Z(n13184) );
  OAI21_X1 U15349 ( .B1(n13184), .B2(n13332), .A(n13183), .ZN(n13386) );
  OR2_X1 U15350 ( .A1(n13186), .A2(n13185), .ZN(n13382) );
  AND3_X1 U15351 ( .A1(n13381), .A2(n13382), .A3(n11149), .ZN(n13193) );
  AOI21_X1 U15352 ( .B1(n13189), .B2(n13199), .A(n13336), .ZN(n13187) );
  NAND2_X1 U15353 ( .A1(n13187), .A2(n6651), .ZN(n13383) );
  AOI22_X1 U15354 ( .A1(n13188), .A2(n14759), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14761), .ZN(n13191) );
  NAND2_X1 U15355 ( .A1(n13189), .A2(n13366), .ZN(n13190) );
  OAI211_X1 U15356 ( .C1(n13383), .C2(n13363), .A(n13191), .B(n13190), .ZN(
        n13192) );
  AOI211_X1 U15357 ( .C1(n13386), .C2(n13357), .A(n13193), .B(n13192), .ZN(
        n13194) );
  INV_X1 U15358 ( .A(n13194), .ZN(P2_U3238) );
  XNOR2_X1 U15359 ( .A(n13195), .B(n13205), .ZN(n13198) );
  INV_X1 U15360 ( .A(n13196), .ZN(n13197) );
  AOI21_X1 U15361 ( .B1(n13198), .B2(n13350), .A(n13197), .ZN(n13390) );
  INV_X1 U15362 ( .A(n13213), .ZN(n13201) );
  INV_X1 U15363 ( .A(n13199), .ZN(n13200) );
  AOI211_X1 U15364 ( .C1(n13388), .C2(n13201), .A(n13336), .B(n13200), .ZN(
        n13387) );
  AOI22_X1 U15365 ( .A1(n13202), .A2(n14759), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14761), .ZN(n13203) );
  OAI21_X1 U15366 ( .B1(n13204), .B2(n14764), .A(n13203), .ZN(n13208) );
  XNOR2_X1 U15367 ( .A(n13206), .B(n13205), .ZN(n13391) );
  NOR2_X1 U15368 ( .A1(n13391), .A2(n13369), .ZN(n13207) );
  OAI21_X1 U15369 ( .B1(n13390), .B2(n14761), .A(n13209), .ZN(P2_U3239) );
  XNOR2_X1 U15370 ( .A(n13210), .B(n13219), .ZN(n13212) );
  AOI21_X1 U15371 ( .B1(n13212), .B2(n13350), .A(n13211), .ZN(n13395) );
  AOI211_X1 U15372 ( .C1(n13393), .C2(n13226), .A(n13336), .B(n13213), .ZN(
        n13392) );
  INV_X1 U15373 ( .A(n13214), .ZN(n13215) );
  AOI22_X1 U15374 ( .A1(n13215), .A2(n14759), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n14761), .ZN(n13216) );
  OAI21_X1 U15375 ( .B1(n13217), .B2(n14764), .A(n13216), .ZN(n13221) );
  XNOR2_X1 U15376 ( .A(n13219), .B(n13218), .ZN(n13396) );
  NOR2_X1 U15377 ( .A1(n13396), .A2(n13369), .ZN(n13220) );
  AOI211_X1 U15378 ( .C1(n13392), .C2(n14757), .A(n13221), .B(n13220), .ZN(
        n13222) );
  OAI21_X1 U15379 ( .B1(n13395), .B2(n14761), .A(n13222), .ZN(P2_U3240) );
  XNOR2_X1 U15380 ( .A(n13223), .B(n13230), .ZN(n13225) );
  AOI21_X1 U15381 ( .B1(n13225), .B2(n13350), .A(n13224), .ZN(n13400) );
  INV_X1 U15382 ( .A(n13246), .ZN(n13228) );
  INV_X1 U15383 ( .A(n13226), .ZN(n13227) );
  AOI211_X1 U15384 ( .C1(n13398), .C2(n13228), .A(n13336), .B(n13227), .ZN(
        n13397) );
  NAND2_X1 U15385 ( .A1(n13230), .A2(n13229), .ZN(n13231) );
  NAND2_X1 U15386 ( .A1(n13232), .A2(n13231), .ZN(n13401) );
  NOR2_X1 U15387 ( .A1(n13401), .A2(n13369), .ZN(n13237) );
  AOI22_X1 U15388 ( .A1(n13233), .A2(n14759), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n14761), .ZN(n13234) );
  OAI21_X1 U15389 ( .B1(n13235), .B2(n14764), .A(n13234), .ZN(n13236) );
  AOI211_X1 U15390 ( .C1(n13397), .C2(n13338), .A(n13237), .B(n13236), .ZN(
        n13238) );
  OAI21_X1 U15391 ( .B1(n13400), .B2(n14761), .A(n13238), .ZN(P2_U3241) );
  XNOR2_X1 U15392 ( .A(n13239), .B(n13241), .ZN(n13407) );
  XOR2_X1 U15393 ( .A(n13241), .B(n13240), .Z(n13242) );
  NAND2_X1 U15394 ( .A1(n13242), .A2(n13350), .ZN(n13406) );
  INV_X1 U15395 ( .A(n13403), .ZN(n13243) );
  OAI211_X1 U15396 ( .C1(n13354), .C2(n13244), .A(n13406), .B(n13243), .ZN(
        n13245) );
  NAND2_X1 U15397 ( .A1(n13245), .A2(n13357), .ZN(n13251) );
  AOI211_X1 U15398 ( .C1(n13404), .C2(n13258), .A(n13336), .B(n13246), .ZN(
        n13402) );
  OAI22_X1 U15399 ( .A1(n13248), .A2(n14764), .B1(n13357), .B2(n13247), .ZN(
        n13249) );
  AOI21_X1 U15400 ( .B1(n13402), .B2(n14757), .A(n13249), .ZN(n13250) );
  OAI211_X1 U15401 ( .C1(n13407), .C2(n13369), .A(n13251), .B(n13250), .ZN(
        P2_U3242) );
  XNOR2_X1 U15402 ( .A(n13253), .B(n13252), .ZN(n13412) );
  XNOR2_X1 U15403 ( .A(n13255), .B(n13254), .ZN(n13257) );
  OAI21_X1 U15404 ( .B1(n13257), .B2(n13332), .A(n13256), .ZN(n13408) );
  INV_X1 U15405 ( .A(n13258), .ZN(n13259) );
  AOI211_X1 U15406 ( .C1(n13410), .C2(n13274), .A(n13336), .B(n13259), .ZN(
        n13409) );
  NAND2_X1 U15407 ( .A1(n13409), .A2(n14757), .ZN(n13263) );
  INV_X1 U15408 ( .A(n13260), .ZN(n13261) );
  AOI22_X1 U15409 ( .A1(n13261), .A2(n14759), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n14761), .ZN(n13262) );
  OAI211_X1 U15410 ( .C1(n13264), .C2(n14764), .A(n13263), .B(n13262), .ZN(
        n13265) );
  AOI21_X1 U15411 ( .B1(n13408), .B2(n13357), .A(n13265), .ZN(n13266) );
  OAI21_X1 U15412 ( .B1(n13412), .B2(n13369), .A(n13266), .ZN(P2_U3243) );
  XNOR2_X1 U15413 ( .A(n13267), .B(n13270), .ZN(n13417) );
  NAND2_X1 U15414 ( .A1(n13284), .A2(n13285), .ZN(n13283) );
  NAND2_X1 U15415 ( .A1(n13283), .A2(n13269), .ZN(n13271) );
  XNOR2_X1 U15416 ( .A(n13271), .B(n13270), .ZN(n13273) );
  OAI21_X1 U15417 ( .B1(n13273), .B2(n13332), .A(n13272), .ZN(n13413) );
  AOI21_X1 U15418 ( .B1(n13289), .B2(n13415), .A(n13336), .ZN(n13275) );
  AND2_X1 U15419 ( .A1(n13275), .A2(n13274), .ZN(n13414) );
  NAND2_X1 U15420 ( .A1(n13414), .A2(n14757), .ZN(n13278) );
  AOI22_X1 U15421 ( .A1(n13276), .A2(n14759), .B1(n14761), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n13277) );
  OAI211_X1 U15422 ( .C1(n13279), .C2(n14764), .A(n13278), .B(n13277), .ZN(
        n13280) );
  AOI21_X1 U15423 ( .B1(n13413), .B2(n13357), .A(n13280), .ZN(n13281) );
  OAI21_X1 U15424 ( .B1(n13417), .B2(n13369), .A(n13281), .ZN(P2_U3244) );
  XNOR2_X1 U15425 ( .A(n13282), .B(n13285), .ZN(n13422) );
  OAI21_X1 U15426 ( .B1(n13285), .B2(n13284), .A(n13283), .ZN(n13287) );
  AOI21_X1 U15427 ( .B1(n13287), .B2(n13350), .A(n13286), .ZN(n13421) );
  INV_X1 U15428 ( .A(n13421), .ZN(n13296) );
  OR2_X1 U15429 ( .A1(n13299), .A2(n13294), .ZN(n13288) );
  AND3_X1 U15430 ( .A1(n13289), .A2(n13359), .A3(n13288), .ZN(n13418) );
  NAND2_X1 U15431 ( .A1(n13418), .A2(n13338), .ZN(n13293) );
  INV_X1 U15432 ( .A(n13290), .ZN(n13291) );
  AOI22_X1 U15433 ( .A1(P2_REG2_REG_20__SCAN_IN), .A2(n14761), .B1(n13291), 
        .B2(n14759), .ZN(n13292) );
  OAI211_X1 U15434 ( .C1(n13294), .C2(n14764), .A(n13293), .B(n13292), .ZN(
        n13295) );
  AOI21_X1 U15435 ( .B1(n13296), .B2(n13357), .A(n13295), .ZN(n13297) );
  OAI21_X1 U15436 ( .B1(n13422), .B2(n13369), .A(n13297), .ZN(P2_U3245) );
  XNOR2_X1 U15437 ( .A(n13298), .B(n13302), .ZN(n13428) );
  AOI211_X1 U15438 ( .C1(n13425), .C2(n13320), .A(n13336), .B(n13299), .ZN(
        n13423) );
  INV_X1 U15439 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13300) );
  OAI22_X1 U15440 ( .A1(n13301), .A2(n14764), .B1(n13357), .B2(n13300), .ZN(
        n13309) );
  XNOR2_X1 U15441 ( .A(n13303), .B(n13302), .ZN(n13304) );
  NAND2_X1 U15442 ( .A1(n13304), .A2(n13350), .ZN(n13427) );
  INV_X1 U15443 ( .A(n13305), .ZN(n13306) );
  AOI21_X1 U15444 ( .B1(n13306), .B2(n14759), .A(n13424), .ZN(n13307) );
  AOI21_X1 U15445 ( .B1(n13427), .B2(n13307), .A(n14761), .ZN(n13308) );
  AOI211_X1 U15446 ( .C1(n13423), .C2(n14757), .A(n13309), .B(n13308), .ZN(
        n13310) );
  OAI21_X1 U15447 ( .B1(n13369), .B2(n13428), .A(n13310), .ZN(P2_U3246) );
  NAND2_X1 U15448 ( .A1(n13311), .A2(n13314), .ZN(n13312) );
  XNOR2_X1 U15449 ( .A(n13315), .B(n13314), .ZN(n13316) );
  NAND2_X1 U15450 ( .A1(n13316), .A2(n13350), .ZN(n13432) );
  INV_X1 U15451 ( .A(n13430), .ZN(n13317) );
  OAI211_X1 U15452 ( .C1(n13354), .C2(n13318), .A(n13432), .B(n13317), .ZN(
        n13319) );
  NAND2_X1 U15453 ( .A1(n13319), .A2(n13357), .ZN(n13326) );
  INV_X1 U15454 ( .A(n13320), .ZN(n13321) );
  AOI211_X1 U15455 ( .C1(n13431), .C2(n13334), .A(n13336), .B(n13321), .ZN(
        n13429) );
  OAI22_X1 U15456 ( .A1(n13323), .A2(n14764), .B1(n13357), .B2(n13322), .ZN(
        n13324) );
  AOI21_X1 U15457 ( .B1(n13429), .B2(n14757), .A(n13324), .ZN(n13325) );
  OAI211_X1 U15458 ( .C1(n13434), .C2(n13369), .A(n13326), .B(n13325), .ZN(
        P2_U3247) );
  XNOR2_X1 U15459 ( .A(n13328), .B(n13327), .ZN(n13439) );
  XNOR2_X1 U15460 ( .A(n13330), .B(n13329), .ZN(n13333) );
  OAI21_X1 U15461 ( .B1(n13333), .B2(n13332), .A(n13331), .ZN(n13435) );
  INV_X1 U15462 ( .A(n13362), .ZN(n13337) );
  INV_X1 U15463 ( .A(n13334), .ZN(n13335) );
  AOI211_X1 U15464 ( .C1(n13437), .C2(n13337), .A(n13336), .B(n13335), .ZN(
        n13436) );
  NAND2_X1 U15465 ( .A1(n13436), .A2(n13338), .ZN(n13341) );
  AOI22_X1 U15466 ( .A1(n14761), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13339), 
        .B2(n14759), .ZN(n13340) );
  OAI211_X1 U15467 ( .C1(n13342), .C2(n14764), .A(n13341), .B(n13340), .ZN(
        n13343) );
  AOI21_X1 U15468 ( .B1(n13357), .B2(n13435), .A(n13343), .ZN(n13344) );
  OAI21_X1 U15469 ( .B1(n13439), .B2(n13369), .A(n13344), .ZN(P2_U3248) );
  NAND2_X1 U15470 ( .A1(n13345), .A2(n13349), .ZN(n13346) );
  NAND2_X1 U15471 ( .A1(n13347), .A2(n13346), .ZN(n13443) );
  XNOR2_X1 U15472 ( .A(n13348), .B(n13349), .ZN(n13351) );
  NAND2_X1 U15473 ( .A1(n13351), .A2(n13350), .ZN(n13353) );
  NAND2_X1 U15474 ( .A1(n13353), .A2(n13352), .ZN(n13445) );
  NAND2_X1 U15475 ( .A1(n13445), .A2(n13357), .ZN(n13368) );
  OAI22_X1 U15476 ( .A1(n13357), .A2(n13356), .B1(n13355), .B2(n13354), .ZN(
        n13365) );
  NAND2_X1 U15477 ( .A1(n13358), .A2(n13440), .ZN(n13360) );
  NAND2_X1 U15478 ( .A1(n13360), .A2(n13359), .ZN(n13361) );
  OR2_X1 U15479 ( .A1(n13362), .A2(n13361), .ZN(n13442) );
  NOR2_X1 U15480 ( .A1(n13442), .A2(n13363), .ZN(n13364) );
  AOI211_X1 U15481 ( .C1(n13366), .C2(n13440), .A(n13365), .B(n13364), .ZN(
        n13367) );
  OAI211_X1 U15482 ( .C1(n13369), .C2(n13443), .A(n13368), .B(n13367), .ZN(
        P2_U3249) );
  INV_X1 U15483 ( .A(n13370), .ZN(n13372) );
  OAI211_X1 U15484 ( .C1(n13372), .C2(n14826), .A(n13371), .B(n13373), .ZN(
        n13458) );
  MUX2_X1 U15485 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13458), .S(n13457), .Z(
        P2_U3530) );
  OAI211_X1 U15486 ( .C1(n13375), .C2(n14826), .A(n13374), .B(n13373), .ZN(
        n13459) );
  MUX2_X1 U15487 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13459), .S(n14837), .Z(
        P2_U3529) );
  AOI21_X1 U15488 ( .B1(n14792), .B2(n13377), .A(n13376), .ZN(n13378) );
  OAI211_X1 U15489 ( .C1(n13456), .C2(n13380), .A(n13379), .B(n13378), .ZN(
        n13460) );
  MUX2_X1 U15490 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13460), .S(n14837), .Z(
        P2_U3527) );
  NAND3_X1 U15491 ( .A1(n13382), .A2(n14808), .A3(n13381), .ZN(n13384) );
  MUX2_X1 U15492 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13461), .S(n14837), .Z(
        P2_U3526) );
  AOI21_X1 U15493 ( .B1(n14792), .B2(n13388), .A(n13387), .ZN(n13389) );
  OAI211_X1 U15494 ( .C1(n13456), .C2(n13391), .A(n13390), .B(n13389), .ZN(
        n13462) );
  MUX2_X1 U15495 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13462), .S(n14837), .Z(
        P2_U3525) );
  AOI21_X1 U15496 ( .B1(n14792), .B2(n13393), .A(n13392), .ZN(n13394) );
  OAI211_X1 U15497 ( .C1(n13456), .C2(n13396), .A(n13395), .B(n13394), .ZN(
        n13463) );
  MUX2_X1 U15498 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13463), .S(n14837), .Z(
        P2_U3524) );
  AOI21_X1 U15499 ( .B1(n14792), .B2(n13398), .A(n13397), .ZN(n13399) );
  OAI211_X1 U15500 ( .C1(n13456), .C2(n13401), .A(n13400), .B(n13399), .ZN(
        n13464) );
  MUX2_X1 U15501 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13464), .S(n14837), .Z(
        P2_U3523) );
  AOI211_X1 U15502 ( .C1(n14792), .C2(n13404), .A(n13403), .B(n13402), .ZN(
        n13405) );
  OAI211_X1 U15503 ( .C1(n13456), .C2(n13407), .A(n13406), .B(n13405), .ZN(
        n13465) );
  MUX2_X1 U15504 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13465), .S(n13457), .Z(
        P2_U3522) );
  AOI211_X1 U15505 ( .C1(n14792), .C2(n13410), .A(n13409), .B(n13408), .ZN(
        n13411) );
  OAI21_X1 U15506 ( .B1(n13456), .B2(n13412), .A(n13411), .ZN(n13466) );
  MUX2_X1 U15507 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13466), .S(n13457), .Z(
        P2_U3521) );
  AOI211_X1 U15508 ( .C1(n14792), .C2(n13415), .A(n13414), .B(n13413), .ZN(
        n13416) );
  OAI21_X1 U15509 ( .B1(n13456), .B2(n13417), .A(n13416), .ZN(n13467) );
  MUX2_X1 U15510 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13467), .S(n13457), .Z(
        P2_U3520) );
  AOI21_X1 U15511 ( .B1(n14792), .B2(n13419), .A(n13418), .ZN(n13420) );
  OAI211_X1 U15512 ( .C1(n13456), .C2(n13422), .A(n13421), .B(n13420), .ZN(
        n13468) );
  MUX2_X1 U15513 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13468), .S(n13457), .Z(
        P2_U3519) );
  AOI211_X1 U15514 ( .C1(n14792), .C2(n13425), .A(n13424), .B(n13423), .ZN(
        n13426) );
  OAI211_X1 U15515 ( .C1(n13456), .C2(n13428), .A(n13427), .B(n13426), .ZN(
        n13469) );
  MUX2_X1 U15516 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13469), .S(n13457), .Z(
        P2_U3518) );
  AOI211_X1 U15517 ( .C1(n14792), .C2(n13431), .A(n13430), .B(n13429), .ZN(
        n13433) );
  OAI211_X1 U15518 ( .C1(n13456), .C2(n13434), .A(n13433), .B(n13432), .ZN(
        n13470) );
  MUX2_X1 U15519 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13470), .S(n13457), .Z(
        P2_U3517) );
  AOI211_X1 U15520 ( .C1(n14792), .C2(n13437), .A(n13436), .B(n13435), .ZN(
        n13438) );
  OAI21_X1 U15521 ( .B1(n13456), .B2(n13439), .A(n13438), .ZN(n13471) );
  MUX2_X1 U15522 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13471), .S(n13457), .Z(
        P2_U3516) );
  NAND2_X1 U15523 ( .A1(n13440), .A2(n14792), .ZN(n13441) );
  OAI211_X1 U15524 ( .C1(n13443), .C2(n13456), .A(n13442), .B(n13441), .ZN(
        n13444) );
  MUX2_X1 U15525 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13472), .S(n13457), .Z(
        P2_U3515) );
  NOR2_X1 U15526 ( .A1(n13446), .A2(n13456), .ZN(n13449) );
  OAI21_X1 U15527 ( .B1(n9080), .B2(n14826), .A(n13447), .ZN(n13448) );
  OR3_X1 U15528 ( .A1(n13450), .A2(n13449), .A3(n13448), .ZN(n13473) );
  MUX2_X1 U15529 ( .A(n13473), .B(P2_REG1_REG_15__SCAN_IN), .S(n14835), .Z(
        P2_U3514) );
  AOI21_X1 U15530 ( .B1(n14792), .B2(n13452), .A(n13451), .ZN(n13453) );
  OAI211_X1 U15531 ( .C1(n13456), .C2(n13455), .A(n13454), .B(n13453), .ZN(
        n13474) );
  MUX2_X1 U15532 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13474), .S(n13457), .Z(
        P2_U3513) );
  MUX2_X1 U15533 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13458), .S(n6621), .Z(
        P2_U3498) );
  MUX2_X1 U15534 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13459), .S(n6621), .Z(
        P2_U3497) );
  MUX2_X1 U15535 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13460), .S(n6621), .Z(
        P2_U3495) );
  MUX2_X1 U15536 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13461), .S(n6621), .Z(
        P2_U3494) );
  MUX2_X1 U15537 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13462), .S(n6621), .Z(
        P2_U3493) );
  MUX2_X1 U15538 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13463), .S(n6621), .Z(
        P2_U3492) );
  MUX2_X1 U15539 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13464), .S(n6621), .Z(
        P2_U3491) );
  MUX2_X1 U15540 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13465), .S(n6621), .Z(
        P2_U3490) );
  MUX2_X1 U15541 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13466), .S(n6621), .Z(
        P2_U3489) );
  MUX2_X1 U15542 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13467), .S(n6621), .Z(
        P2_U3488) );
  MUX2_X1 U15543 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13468), .S(n6621), .Z(
        P2_U3487) );
  MUX2_X1 U15544 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13469), .S(n6621), .Z(
        P2_U3486) );
  MUX2_X1 U15545 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13470), .S(n6621), .Z(
        P2_U3484) );
  MUX2_X1 U15546 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13471), .S(n6621), .Z(
        P2_U3481) );
  MUX2_X1 U15547 ( .A(n13472), .B(P2_REG0_REG_16__SCAN_IN), .S(n14829), .Z(
        P2_U3478) );
  MUX2_X1 U15548 ( .A(n13473), .B(P2_REG0_REG_15__SCAN_IN), .S(n14829), .Z(
        P2_U3475) );
  MUX2_X1 U15549 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13474), .S(n6621), .Z(
        P2_U3472) );
  INV_X1 U15550 ( .A(n13475), .ZN(n14143) );
  INV_X1 U15551 ( .A(n13477), .ZN(n13479) );
  NOR4_X1 U15552 ( .A1(n13479), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13478), .A4(
        P2_U3088), .ZN(n13480) );
  AOI21_X1 U15553 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n13481), .A(n13480), 
        .ZN(n13482) );
  OAI21_X1 U15554 ( .B1(n14143), .B2(n13505), .A(n13482), .ZN(P2_U3296) );
  OAI222_X1 U15555 ( .A1(n13505), .A2(n13485), .B1(P2_U3088), .B2(n13484), 
        .C1(n13483), .C2(n13498), .ZN(P2_U3297) );
  INV_X1 U15556 ( .A(n13486), .ZN(n14145) );
  OAI222_X1 U15557 ( .A1(n13505), .A2(n14145), .B1(P2_U3088), .B2(n13488), 
        .C1(n13487), .C2(n13498), .ZN(P2_U3298) );
  INV_X1 U15558 ( .A(n13489), .ZN(n14147) );
  OAI222_X1 U15559 ( .A1(n13505), .A2(n14147), .B1(P2_U3088), .B2(n13491), 
        .C1(n13490), .C2(n13498), .ZN(P2_U3299) );
  NAND2_X1 U15560 ( .A1(n14149), .A2(n13492), .ZN(n13494) );
  OAI211_X1 U15561 ( .C1(n13498), .C2(n13495), .A(n13494), .B(n13493), .ZN(
        P2_U3300) );
  INV_X1 U15562 ( .A(n13496), .ZN(n13500) );
  INV_X1 U15563 ( .A(n13497), .ZN(n14153) );
  OAI222_X1 U15564 ( .A1(P2_U3088), .A2(n13500), .B1(n13505), .B2(n14153), 
        .C1(n13499), .C2(n13498), .ZN(P2_U3301) );
  INV_X1 U15565 ( .A(n13501), .ZN(n14156) );
  OAI222_X1 U15566 ( .A1(n13498), .A2(n13503), .B1(n13505), .B2(n14156), .C1(
        P2_U3088), .C2(n13502), .ZN(P2_U3302) );
  OAI222_X1 U15567 ( .A1(P2_U3088), .A2(n13506), .B1(n13505), .B2(n14159), 
        .C1(n13504), .C2(n13498), .ZN(P2_U3303) );
  MUX2_X1 U15568 ( .A(n13508), .B(n13507), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3327) );
  XOR2_X1 U15569 ( .A(n13510), .B(n13509), .Z(n13516) );
  INV_X1 U15570 ( .A(n13830), .ZN(n13512) );
  OAI22_X1 U15571 ( .A1(n13645), .A2(n13512), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13511), .ZN(n13514) );
  OAI22_X1 U15572 ( .A1(n14039), .A2(n13647), .B1(n13646), .B2(n14038), .ZN(
        n13513) );
  AOI211_X1 U15573 ( .C1(n14042), .C2(n13658), .A(n13514), .B(n13513), .ZN(
        n13515) );
  OAI21_X1 U15574 ( .B1(n13516), .B2(n13660), .A(n13515), .ZN(P1_U3214) );
  OAI21_X1 U15575 ( .B1(n13519), .B2(n13518), .A(n13517), .ZN(n13520) );
  NAND2_X1 U15576 ( .A1(n13520), .A2(n13634), .ZN(n13525) );
  OAI22_X1 U15577 ( .A1(n14411), .A2(n13646), .B1(n13647), .B2(n14409), .ZN(
        n13521) );
  AOI211_X1 U15578 ( .C1(n13523), .C2(n13654), .A(n13522), .B(n13521), .ZN(
        n13524) );
  OAI211_X1 U15579 ( .C1(n9532), .C2(n13640), .A(n13525), .B(n13524), .ZN(
        P1_U3215) );
  XOR2_X1 U15580 ( .A(n13527), .B(n13526), .Z(n13534) );
  NAND2_X1 U15581 ( .A1(n13664), .A2(n14634), .ZN(n13529) );
  NAND2_X1 U15582 ( .A1(n13860), .A2(n14617), .ZN(n13528) );
  AND2_X1 U15583 ( .A1(n13529), .A2(n13528), .ZN(n13889) );
  OAI22_X1 U15584 ( .A1(n13656), .A2(n13889), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13530), .ZN(n13531) );
  AOI21_X1 U15585 ( .B1(n13898), .B2(n13654), .A(n13531), .ZN(n13533) );
  NAND2_X1 U15586 ( .A1(n13899), .A2(n13658), .ZN(n13532) );
  OAI211_X1 U15587 ( .C1(n13534), .C2(n13660), .A(n13533), .B(n13532), .ZN(
        P1_U3216) );
  OAI211_X1 U15588 ( .C1(n13537), .C2(n13536), .A(n13535), .B(n13634), .ZN(
        n13543) );
  AOI22_X1 U15589 ( .A1(n13671), .A2(n14617), .B1(n14634), .B2(n9894), .ZN(
        n14532) );
  INV_X1 U15590 ( .A(n14532), .ZN(n13539) );
  AOI22_X1 U15591 ( .A1(n13540), .A2(n13539), .B1(n13658), .B2(n6626), .ZN(
        n13542) );
  MUX2_X1 U15592 ( .A(P1_STATE_REG_SCAN_IN), .B(n13645), .S(n14537), .Z(n13541) );
  NAND3_X1 U15593 ( .A1(n13543), .A2(n13542), .A3(n13541), .ZN(P1_U3218) );
  INV_X1 U15594 ( .A(n13646), .ZN(n13596) );
  AOI22_X1 U15595 ( .A1(n13596), .A2(n13959), .B1(n13595), .B2(n13933), .ZN(
        n13544) );
  NAND2_X1 U15596 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13798)
         );
  OAI211_X1 U15597 ( .C1(n13645), .C2(n13961), .A(n13544), .B(n13798), .ZN(
        n13550) );
  INV_X1 U15598 ( .A(n13545), .ZN(n13546) );
  AOI211_X1 U15599 ( .C1(n13548), .C2(n13547), .A(n13660), .B(n13546), .ZN(
        n13549) );
  AOI211_X1 U15600 ( .C1(n14106), .C2(n13658), .A(n13550), .B(n13549), .ZN(
        n13551) );
  INV_X1 U15601 ( .A(n13551), .ZN(P1_U3219) );
  OAI21_X1 U15602 ( .B1(n13555), .B2(n13554), .A(n13553), .ZN(n13556) );
  NAND2_X1 U15603 ( .A1(n13556), .A2(n13634), .ZN(n13560) );
  AOI22_X1 U15604 ( .A1(n13658), .A2(n14558), .B1(n13557), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n13559) );
  AOI22_X1 U15605 ( .A1(n13595), .A2(n9894), .B1(n13596), .B2(n10709), .ZN(
        n13558) );
  NAND3_X1 U15606 ( .A1(n13560), .A2(n13559), .A3(n13558), .ZN(P1_U3222) );
  OAI21_X1 U15607 ( .B1(n13563), .B2(n13562), .A(n13561), .ZN(n13564) );
  NAND2_X1 U15608 ( .A1(n13564), .A2(n13634), .ZN(n13569) );
  NOR2_X1 U15609 ( .A1(n13565), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13567) );
  OAI22_X1 U15610 ( .A1(n14103), .A2(n13646), .B1(n13647), .B2(n14085), .ZN(
        n13566) );
  AOI211_X1 U15611 ( .C1(n13654), .C2(n13929), .A(n13567), .B(n13566), .ZN(
        n13568) );
  OAI211_X1 U15612 ( .C1(n7210), .C2(n13640), .A(n13569), .B(n13568), .ZN(
        P1_U3223) );
  XOR2_X1 U15613 ( .A(n13571), .B(n13570), .Z(n13578) );
  INV_X1 U15614 ( .A(n13864), .ZN(n13573) );
  OAI22_X1 U15615 ( .A1(n13645), .A2(n13573), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13572), .ZN(n13576) );
  OAI22_X1 U15616 ( .A1(n14038), .A2(n13647), .B1(n13646), .B2(n13574), .ZN(
        n13575) );
  AOI211_X1 U15617 ( .C1(n14057), .C2(n13658), .A(n13576), .B(n13575), .ZN(
        n13577) );
  OAI21_X1 U15618 ( .B1(n13578), .B2(n13660), .A(n13577), .ZN(P1_U3225) );
  OAI21_X1 U15619 ( .B1(n13581), .B2(n13580), .A(n13579), .ZN(n13582) );
  NAND2_X1 U15620 ( .A1(n13582), .A2(n13634), .ZN(n13589) );
  INV_X1 U15621 ( .A(n13583), .ZN(n13586) );
  OAI22_X1 U15622 ( .A1(n13584), .A2(n13647), .B1(n13646), .B2(n14409), .ZN(
        n13585) );
  AOI211_X1 U15623 ( .C1(n13654), .C2(n13587), .A(n13586), .B(n13585), .ZN(
        n13588) );
  OAI211_X1 U15624 ( .C1(n14397), .C2(n13640), .A(n13589), .B(n13588), .ZN(
        P1_U3226) );
  INV_X1 U15625 ( .A(n13590), .ZN(n13591) );
  NOR2_X1 U15626 ( .A1(n13592), .A2(n13591), .ZN(n13593) );
  XNOR2_X1 U15627 ( .A(n13594), .B(n13593), .ZN(n13602) );
  INV_X1 U15628 ( .A(n14001), .ZN(n13599) );
  AOI22_X1 U15629 ( .A1(n13596), .A2(n13666), .B1(n13595), .B2(n13959), .ZN(
        n13598) );
  OAI211_X1 U15630 ( .C1(n13645), .C2(n13599), .A(n13598), .B(n13597), .ZN(
        n13600) );
  AOI21_X1 U15631 ( .B1(n14116), .B2(n13658), .A(n13600), .ZN(n13601) );
  OAI21_X1 U15632 ( .B1(n13602), .B2(n13660), .A(n13601), .ZN(P1_U3228) );
  XOR2_X1 U15633 ( .A(n13604), .B(n13603), .Z(n13610) );
  INV_X1 U15634 ( .A(n13882), .ZN(n13606) );
  OAI22_X1 U15635 ( .A1(n13645), .A2(n13606), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13605), .ZN(n13608) );
  OAI22_X1 U15636 ( .A1(n13873), .A2(n13647), .B1(n13646), .B2(n13916), .ZN(
        n13607) );
  AOI211_X1 U15637 ( .C1(n14066), .C2(n13658), .A(n13608), .B(n13607), .ZN(
        n13609) );
  OAI21_X1 U15638 ( .B1(n13610), .B2(n13660), .A(n13609), .ZN(P1_U3229) );
  OAI211_X1 U15639 ( .C1(n13613), .C2(n13612), .A(n13611), .B(n13634), .ZN(
        n13619) );
  INV_X1 U15640 ( .A(n13943), .ZN(n13617) );
  AND2_X1 U15641 ( .A1(n14076), .A2(n14617), .ZN(n13614) );
  AOI21_X1 U15642 ( .B1(n13665), .B2(n14634), .A(n13614), .ZN(n13940) );
  OAI22_X1 U15643 ( .A1(n13656), .A2(n13940), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13615), .ZN(n13616) );
  AOI21_X1 U15644 ( .B1(n13617), .B2(n13654), .A(n13616), .ZN(n13618) );
  OAI211_X1 U15645 ( .C1(n14096), .C2(n13640), .A(n13619), .B(n13618), .ZN(
        P1_U3233) );
  OAI21_X1 U15646 ( .B1(n13622), .B2(n13621), .A(n13620), .ZN(n13623) );
  NAND2_X1 U15647 ( .A1(n13623), .A2(n13634), .ZN(n13630) );
  OAI22_X1 U15648 ( .A1(n13916), .A2(n13647), .B1(n13646), .B2(n13624), .ZN(
        n13628) );
  INV_X1 U15649 ( .A(n13625), .ZN(n13911) );
  OAI22_X1 U15650 ( .A1(n13645), .A2(n13911), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13626), .ZN(n13627) );
  NOR2_X1 U15651 ( .A1(n13628), .A2(n13627), .ZN(n13629) );
  OAI211_X1 U15652 ( .C1(n13640), .C2(n14080), .A(n13630), .B(n13629), .ZN(
        P1_U3235) );
  OAI21_X1 U15653 ( .B1(n13633), .B2(n13632), .A(n13631), .ZN(n13635) );
  NAND2_X1 U15654 ( .A1(n13635), .A2(n13634), .ZN(n13639) );
  INV_X1 U15655 ( .A(n13636), .ZN(n13983) );
  AOI22_X1 U15656 ( .A1(n13665), .A2(n14617), .B1(n14634), .B2(n14394), .ZN(
        n13977) );
  NAND2_X1 U15657 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14496)
         );
  OAI21_X1 U15658 ( .B1(n13656), .B2(n13977), .A(n14496), .ZN(n13637) );
  AOI21_X1 U15659 ( .B1(n13983), .B2(n13654), .A(n13637), .ZN(n13638) );
  OAI211_X1 U15660 ( .C1(n13985), .C2(n13640), .A(n13639), .B(n13638), .ZN(
        P1_U3238) );
  XOR2_X1 U15661 ( .A(n13642), .B(n13641), .Z(n13651) );
  INV_X1 U15662 ( .A(n13846), .ZN(n13644) );
  OAI22_X1 U15663 ( .A1(n13645), .A2(n13644), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13643), .ZN(n13649) );
  OAI22_X1 U15664 ( .A1(n13845), .A2(n13647), .B1(n13646), .B2(n13873), .ZN(
        n13648) );
  AOI211_X1 U15665 ( .C1(n13851), .C2(n13658), .A(n13649), .B(n13648), .ZN(
        n13650) );
  OAI21_X1 U15666 ( .B1(n13651), .B2(n13660), .A(n13650), .ZN(P1_U3240) );
  XNOR2_X1 U15667 ( .A(n13653), .B(n13652), .ZN(n13661) );
  AOI22_X1 U15668 ( .A1(n9531), .A2(n14634), .B1(n14617), .B2(n13666), .ZN(
        n14363) );
  NAND2_X1 U15669 ( .A1(n13654), .A2(n14365), .ZN(n13655) );
  NAND2_X1 U15670 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14482)
         );
  OAI211_X1 U15671 ( .C1(n14363), .C2(n13656), .A(n13655), .B(n14482), .ZN(
        n13657) );
  AOI21_X1 U15672 ( .B1(n14366), .B2(n13658), .A(n13657), .ZN(n13659) );
  OAI21_X1 U15673 ( .B1(n13661), .B2(n13660), .A(n13659), .ZN(P1_U3241) );
  MUX2_X1 U15674 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13801), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15675 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13662), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15676 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14031), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15677 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13663), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15678 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14047), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15679 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13859), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15680 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14046), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15681 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13860), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15682 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14077), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15683 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13664), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15684 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14076), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15685 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13933), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15686 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13665), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15687 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13959), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15688 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14394), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15689 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13666), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15690 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14393), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15691 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9531), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15692 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14289), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15693 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13667), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15694 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14288), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15695 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13668), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U15696 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14633), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15697 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13669), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U15698 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14616), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15699 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13670), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15700 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14584), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15701 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13671), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15702 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14583), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U15703 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9894), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15704 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n10359), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15705 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n10709), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U15706 ( .C1(n13675), .C2(n13674), .A(n14489), .B(n13673), .ZN(
        n13683) );
  AOI22_X1 U15707 ( .A1(n14468), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n13682) );
  NAND2_X1 U15708 ( .A1(n13792), .A2(n13676), .ZN(n13681) );
  OAI211_X1 U15709 ( .C1(n13679), .C2(n13678), .A(n14486), .B(n13677), .ZN(
        n13680) );
  NAND4_X1 U15710 ( .A1(n13683), .A2(n13682), .A3(n13681), .A4(n13680), .ZN(
        P1_U3244) );
  AOI22_X1 U15711 ( .A1(n14468), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n13697) );
  OAI21_X1 U15712 ( .B1(n13685), .B2(n13684), .A(n13700), .ZN(n13694) );
  MUX2_X1 U15713 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10415), .S(n13690), .Z(
        n13688) );
  INV_X1 U15714 ( .A(n13686), .ZN(n13687) );
  NAND2_X1 U15715 ( .A1(n13688), .A2(n13687), .ZN(n13689) );
  NAND3_X1 U15716 ( .A1(n14486), .A2(n13707), .A3(n13689), .ZN(n13693) );
  INV_X1 U15717 ( .A(n13690), .ZN(n13691) );
  NAND2_X1 U15718 ( .A1(n13792), .A2(n13691), .ZN(n13692) );
  OAI211_X1 U15719 ( .C1(n14477), .C2(n13694), .A(n13693), .B(n13692), .ZN(
        n13695) );
  INV_X1 U15720 ( .A(n13695), .ZN(n13696) );
  NAND3_X1 U15721 ( .A1(n13698), .A2(n13697), .A3(n13696), .ZN(P1_U3245) );
  MUX2_X1 U15722 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10434), .S(n13705), .Z(
        n13701) );
  NAND3_X1 U15723 ( .A1(n13701), .A2(n13700), .A3(n13699), .ZN(n13702) );
  NAND3_X1 U15724 ( .A1(n14489), .A2(n13703), .A3(n13702), .ZN(n13714) );
  AOI22_X1 U15725 ( .A1(n14468), .A2(P1_ADDR_REG_3__SCAN_IN), .B1(
        P1_REG3_REG_3__SCAN_IN), .B2(P1_U3086), .ZN(n13713) );
  INV_X1 U15726 ( .A(n13705), .ZN(n13704) );
  NAND2_X1 U15727 ( .A1(n13792), .A2(n13704), .ZN(n13712) );
  MUX2_X1 U15728 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n14648), .S(n13705), .Z(
        n13708) );
  NAND3_X1 U15729 ( .A1(n13708), .A2(n13707), .A3(n13706), .ZN(n13709) );
  NAND3_X1 U15730 ( .A1(n14486), .A2(n13710), .A3(n13709), .ZN(n13711) );
  NAND4_X1 U15731 ( .A1(n13714), .A2(n13713), .A3(n13712), .A4(n13711), .ZN(
        P1_U3246) );
  INV_X1 U15732 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n13716) );
  NAND2_X1 U15733 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n13715) );
  OAI21_X1 U15734 ( .B1(n14498), .B2(n13716), .A(n13715), .ZN(n13717) );
  AOI21_X1 U15735 ( .B1(n13722), .B2(n13792), .A(n13717), .ZN(n13730) );
  OAI21_X1 U15736 ( .B1(n13720), .B2(n13719), .A(n13718), .ZN(n13721) );
  NAND2_X1 U15737 ( .A1(n14486), .A2(n13721), .ZN(n13729) );
  MUX2_X1 U15738 ( .A(n13723), .B(P1_REG2_REG_5__SCAN_IN), .S(n13722), .Z(
        n13724) );
  NAND3_X1 U15739 ( .A1(n13726), .A2(n13725), .A3(n13724), .ZN(n13727) );
  NAND3_X1 U15740 ( .A1(n14489), .A2(n13740), .A3(n13727), .ZN(n13728) );
  NAND3_X1 U15741 ( .A1(n13730), .A2(n13729), .A3(n13728), .ZN(P1_U3248) );
  AOI211_X1 U15742 ( .C1(n13733), .C2(n13732), .A(n13731), .B(n14479), .ZN(
        n13734) );
  INV_X1 U15743 ( .A(n13734), .ZN(n13745) );
  NOR2_X1 U15744 ( .A1(n14498), .A2(n14177), .ZN(n13735) );
  AOI211_X1 U15745 ( .C1(n13792), .C2(n13737), .A(n13736), .B(n13735), .ZN(
        n13744) );
  MUX2_X1 U15746 ( .A(n10904), .B(P1_REG2_REG_6__SCAN_IN), .S(n13737), .Z(
        n13738) );
  NAND3_X1 U15747 ( .A1(n13740), .A2(n13739), .A3(n13738), .ZN(n13741) );
  NAND3_X1 U15748 ( .A1(n14489), .A2(n13742), .A3(n13741), .ZN(n13743) );
  NAND3_X1 U15749 ( .A1(n13745), .A2(n13744), .A3(n13743), .ZN(P1_U3249) );
  INV_X1 U15750 ( .A(n13746), .ZN(n13751) );
  NOR3_X1 U15751 ( .A1(n13749), .A2(n13748), .A3(n13747), .ZN(n13750) );
  OAI21_X1 U15752 ( .B1(n13751), .B2(n13750), .A(n14486), .ZN(n13761) );
  OAI21_X1 U15753 ( .B1(n14498), .B2(n14184), .A(n13752), .ZN(n13753) );
  AOI21_X1 U15754 ( .B1(n13754), .B2(n13792), .A(n13753), .ZN(n13760) );
  MUX2_X1 U15755 ( .A(n10545), .B(P1_REG2_REG_9__SCAN_IN), .S(n13754), .Z(
        n13755) );
  NAND3_X1 U15756 ( .A1(n13757), .A2(n13756), .A3(n13755), .ZN(n13758) );
  NAND3_X1 U15757 ( .A1(n14489), .A2(n13772), .A3(n13758), .ZN(n13759) );
  NAND3_X1 U15758 ( .A1(n13761), .A2(n13760), .A3(n13759), .ZN(P1_U3252) );
  AOI211_X1 U15759 ( .C1(n13764), .C2(n13763), .A(n14479), .B(n13762), .ZN(
        n13765) );
  INV_X1 U15760 ( .A(n13765), .ZN(n13777) );
  INV_X1 U15761 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14186) );
  NOR2_X1 U15762 ( .A1(n14498), .A2(n14186), .ZN(n13766) );
  AOI211_X1 U15763 ( .C1(n13792), .C2(n13768), .A(n13767), .B(n13766), .ZN(
        n13776) );
  MUX2_X1 U15764 ( .A(n13769), .B(P1_REG2_REG_10__SCAN_IN), .S(n13768), .Z(
        n13770) );
  NAND3_X1 U15765 ( .A1(n13772), .A2(n13771), .A3(n13770), .ZN(n13773) );
  NAND3_X1 U15766 ( .A1(n14489), .A2(n13774), .A3(n13773), .ZN(n13775) );
  NAND3_X1 U15767 ( .A1(n13777), .A2(n13776), .A3(n13775), .ZN(P1_U3253) );
  AOI22_X1 U15768 ( .A1(n13780), .A2(n13779), .B1(n13778), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n13781) );
  OR2_X1 U15769 ( .A1(n13781), .A2(n14493), .ZN(n13782) );
  XNOR2_X1 U15770 ( .A(n13781), .B(n13787), .ZN(n14487) );
  NAND2_X1 U15771 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n14487), .ZN(n14485) );
  NAND2_X1 U15772 ( .A1(n13782), .A2(n14485), .ZN(n13783) );
  XNOR2_X1 U15773 ( .A(n13784), .B(n13783), .ZN(n13795) );
  INV_X1 U15774 ( .A(n13795), .ZN(n13793) );
  NAND2_X1 U15775 ( .A1(n13786), .A2(n13785), .ZN(n13788) );
  XOR2_X1 U15776 ( .A(n13787), .B(n13788), .Z(n14490) );
  NAND2_X1 U15777 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14490), .ZN(n14488) );
  NAND2_X1 U15778 ( .A1(n13788), .A2(n13787), .ZN(n13789) );
  NAND2_X1 U15779 ( .A1(n14488), .A2(n13789), .ZN(n13790) );
  XOR2_X1 U15780 ( .A(n13790), .B(P1_REG2_REG_19__SCAN_IN), .Z(n13794) );
  NOR2_X1 U15781 ( .A1(n13794), .A2(n14477), .ZN(n13791) );
  AOI211_X1 U15782 ( .C1(n13793), .C2(n14486), .A(n13792), .B(n13791), .ZN(
        n13797) );
  AOI22_X1 U15783 ( .A1(n13795), .A2(n14486), .B1(n14489), .B2(n13794), .ZN(
        n13796) );
  MUX2_X1 U15784 ( .A(n13797), .B(n13796), .S(n13930), .Z(n13799) );
  OAI211_X1 U15785 ( .C1(n6890), .C2(n14498), .A(n13799), .B(n13798), .ZN(
        P1_U3262) );
  NOR2_X1 U15786 ( .A1(n13806), .A2(n13808), .ZN(n13800) );
  XOR2_X1 U15787 ( .A(n13800), .B(n14019), .Z(n14021) );
  INV_X1 U15788 ( .A(n14014), .ZN(n13805) );
  NAND2_X1 U15789 ( .A1(n13802), .A2(n13801), .ZN(n14022) );
  NOR2_X1 U15790 ( .A1(n14539), .A2(n14022), .ZN(n13810) );
  AOI21_X1 U15791 ( .B1(n14539), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13810), 
        .ZN(n13804) );
  NAND2_X1 U15792 ( .A1(n14019), .A2(n14382), .ZN(n13803) );
  OAI211_X1 U15793 ( .C1(n14021), .C2(n13805), .A(n13804), .B(n13803), .ZN(
        P1_U3263) );
  XOR2_X1 U15794 ( .A(n13808), .B(n13806), .Z(n13807) );
  NAND2_X1 U15795 ( .A1(n13807), .A2(n14559), .ZN(n14023) );
  INV_X1 U15796 ( .A(n13808), .ZN(n14024) );
  NOR2_X1 U15797 ( .A1(n14024), .A2(n14541), .ZN(n13809) );
  AOI211_X1 U15798 ( .C1(n14539), .C2(P1_REG2_REG_30__SCAN_IN), .A(n13810), 
        .B(n13809), .ZN(n13811) );
  OAI21_X1 U15799 ( .B1(n13902), .B2(n14023), .A(n13811), .ZN(P1_U3264) );
  NAND2_X1 U15800 ( .A1(n14006), .A2(n14376), .ZN(n13956) );
  AND2_X1 U15801 ( .A1(n13821), .A2(n13827), .ZN(n13814) );
  OR3_X1 U15802 ( .A1(n13815), .A2(n13814), .A3(n10341), .ZN(n14033) );
  OR2_X1 U15803 ( .A1(n13966), .A2(n13816), .ZN(n13819) );
  AOI22_X1 U15804 ( .A1(n14539), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n13817), 
        .B2(n14538), .ZN(n13818) );
  OAI211_X1 U15805 ( .C1(n13845), .C2(n13849), .A(n13819), .B(n13818), .ZN(
        n13820) );
  AOI21_X1 U15806 ( .B1(n13821), .B2(n14382), .A(n13820), .ZN(n13822) );
  OAI21_X1 U15807 ( .B1(n14033), .B2(n13902), .A(n13822), .ZN(n13823) );
  AOI21_X1 U15808 ( .B1(n6652), .B2(n14390), .A(n13823), .ZN(n13824) );
  OAI21_X1 U15809 ( .B1(n14037), .B2(n13956), .A(n13824), .ZN(P1_U3265) );
  XNOR2_X1 U15810 ( .A(n13825), .B(n13837), .ZN(n13826) );
  NAND2_X1 U15811 ( .A1(n13826), .A2(n14376), .ZN(n14044) );
  INV_X1 U15812 ( .A(n6664), .ZN(n13829) );
  INV_X1 U15813 ( .A(n13827), .ZN(n13828) );
  AOI211_X1 U15814 ( .C1(n14042), .C2(n13829), .A(n10341), .B(n13828), .ZN(
        n14040) );
  AOI22_X1 U15815 ( .A1(n14539), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13830), 
        .B2(n14538), .ZN(n13831) );
  OAI21_X1 U15816 ( .B1(n13966), .B2(n14039), .A(n13831), .ZN(n13832) );
  AOI21_X1 U15817 ( .B1(n13960), .B2(n13859), .A(n13832), .ZN(n13833) );
  OAI21_X1 U15818 ( .B1(n13834), .B2(n14541), .A(n13833), .ZN(n13839) );
  AOI21_X1 U15819 ( .B1(n13837), .B2(n13836), .A(n13835), .ZN(n14045) );
  NOR2_X1 U15820 ( .A1(n14045), .A2(n14009), .ZN(n13838) );
  AOI211_X1 U15821 ( .C1(n14040), .C2(n14548), .A(n13839), .B(n13838), .ZN(
        n13840) );
  OAI21_X1 U15822 ( .B1(n14539), .B2(n14044), .A(n13840), .ZN(P1_U3266) );
  XNOR2_X1 U15823 ( .A(n13842), .B(n13841), .ZN(n14056) );
  NAND2_X1 U15824 ( .A1(n13851), .A2(n13863), .ZN(n13843) );
  NAND2_X1 U15825 ( .A1(n13843), .A2(n14559), .ZN(n13844) );
  OR2_X1 U15826 ( .A1(n6664), .A2(n13844), .ZN(n14049) );
  OR2_X1 U15827 ( .A1(n13966), .A2(n13845), .ZN(n13848) );
  AOI22_X1 U15828 ( .A1(n14539), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n13846), 
        .B2(n14538), .ZN(n13847) );
  OAI211_X1 U15829 ( .C1(n13873), .C2(n13849), .A(n13848), .B(n13847), .ZN(
        n13850) );
  AOI21_X1 U15830 ( .B1(n13851), .B2(n14382), .A(n13850), .ZN(n13852) );
  OAI21_X1 U15831 ( .B1(n14049), .B2(n13902), .A(n13852), .ZN(n13853) );
  INV_X1 U15832 ( .A(n13853), .ZN(n13857) );
  OR2_X1 U15833 ( .A1(n13855), .A2(n13854), .ZN(n14053) );
  NAND3_X1 U15834 ( .A1(n14053), .A2(n14390), .A3(n14052), .ZN(n13856) );
  OAI211_X1 U15835 ( .C1(n14056), .C2(n13956), .A(n13857), .B(n13856), .ZN(
        P1_U3267) );
  XNOR2_X1 U15836 ( .A(n13868), .B(n13858), .ZN(n13861) );
  AOI222_X1 U15837 ( .A1(n14376), .A2(n13861), .B1(n13860), .B2(n14634), .C1(
        n13859), .C2(n14617), .ZN(n14063) );
  NAND2_X1 U15838 ( .A1(n14057), .A2(n13879), .ZN(n13862) );
  AND2_X1 U15839 ( .A1(n13863), .A2(n13862), .ZN(n14058) );
  AOI22_X1 U15840 ( .A1(n14539), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n13864), 
        .B2(n14538), .ZN(n13865) );
  OAI21_X1 U15841 ( .B1(n7209), .B2(n14541), .A(n13865), .ZN(n13866) );
  AOI21_X1 U15842 ( .B1(n14014), .B2(n14058), .A(n13866), .ZN(n13870) );
  NAND2_X1 U15843 ( .A1(n13868), .A2(n13867), .ZN(n14059) );
  NAND3_X1 U15844 ( .A1(n14060), .A2(n14390), .A3(n14059), .ZN(n13869) );
  OAI211_X1 U15845 ( .C1(n14063), .C2(n14552), .A(n13870), .B(n13869), .ZN(
        P1_U3268) );
  XNOR2_X1 U15846 ( .A(n13872), .B(n13871), .ZN(n14064) );
  OAI22_X1 U15847 ( .A1(n13873), .A2(n14408), .B1(n13916), .B2(n14410), .ZN(
        n13878) );
  AOI211_X1 U15848 ( .C1(n13876), .C2(n13875), .A(n14533), .B(n13874), .ZN(
        n13877) );
  AOI211_X1 U15849 ( .C1(n14536), .C2(n14064), .A(n13878), .B(n13877), .ZN(
        n14068) );
  INV_X1 U15850 ( .A(n13896), .ZN(n13881) );
  INV_X1 U15851 ( .A(n13879), .ZN(n13880) );
  AOI211_X1 U15852 ( .C1(n14066), .C2(n13881), .A(n10341), .B(n13880), .ZN(
        n14065) );
  NAND2_X1 U15853 ( .A1(n14065), .A2(n14548), .ZN(n13884) );
  AOI22_X1 U15854 ( .A1(n14539), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n13882), 
        .B2(n14538), .ZN(n13883) );
  OAI211_X1 U15855 ( .C1(n13885), .C2(n14541), .A(n13884), .B(n13883), .ZN(
        n13886) );
  AOI21_X1 U15856 ( .B1(n14549), .B2(n14064), .A(n13886), .ZN(n13887) );
  OAI21_X1 U15857 ( .B1(n14068), .B2(n14539), .A(n13887), .ZN(P1_U3269) );
  XNOR2_X1 U15858 ( .A(n13888), .B(n13892), .ZN(n13891) );
  INV_X1 U15859 ( .A(n13889), .ZN(n13890) );
  AOI21_X1 U15860 ( .B1(n13891), .B2(n14376), .A(n13890), .ZN(n14075) );
  OR2_X1 U15861 ( .A1(n13893), .A2(n13892), .ZN(n13894) );
  AND2_X1 U15862 ( .A1(n13895), .A2(n13894), .ZN(n14073) );
  NOR2_X1 U15863 ( .A1(n14071), .A2(n13910), .ZN(n13897) );
  OR3_X1 U15864 ( .A1(n13897), .A2(n13896), .A3(n10341), .ZN(n14070) );
  AOI22_X1 U15865 ( .A1(n14539), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n13898), 
        .B2(n14538), .ZN(n13901) );
  NAND2_X1 U15866 ( .A1(n13899), .A2(n14382), .ZN(n13900) );
  OAI211_X1 U15867 ( .C1(n14070), .C2(n13902), .A(n13901), .B(n13900), .ZN(
        n13903) );
  AOI21_X1 U15868 ( .B1(n14073), .B2(n14390), .A(n13903), .ZN(n13904) );
  OAI21_X1 U15869 ( .B1(n14075), .B2(n14539), .A(n13904), .ZN(P1_U3270) );
  XNOR2_X1 U15870 ( .A(n13905), .B(n13906), .ZN(n14083) );
  INV_X1 U15871 ( .A(n14083), .ZN(n13920) );
  NAND2_X1 U15872 ( .A1(n13907), .A2(n13906), .ZN(n13908) );
  AOI21_X1 U15873 ( .B1(n7345), .B2(n13908), .A(n14533), .ZN(n14081) );
  AND2_X1 U15874 ( .A1(n13913), .A2(n13927), .ZN(n13909) );
  OR3_X1 U15875 ( .A1(n13910), .A2(n13909), .A3(n10341), .ZN(n14079) );
  OAI22_X1 U15876 ( .A1(n14079), .A2(n13944), .B1(n13962), .B2(n13911), .ZN(
        n13912) );
  OR2_X1 U15877 ( .A1(n14081), .A2(n13912), .ZN(n13918) );
  NAND2_X1 U15878 ( .A1(n13913), .A2(n14382), .ZN(n13915) );
  AOI22_X1 U15879 ( .A1(n13960), .A2(n14076), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n14539), .ZN(n13914) );
  OAI211_X1 U15880 ( .C1(n13916), .C2(n13966), .A(n13915), .B(n13914), .ZN(
        n13917) );
  AOI21_X1 U15881 ( .B1(n13918), .B2(n14006), .A(n13917), .ZN(n13919) );
  OAI21_X1 U15882 ( .B1(n13920), .B2(n14009), .A(n13919), .ZN(P1_U3271) );
  INV_X1 U15883 ( .A(n13921), .ZN(n13922) );
  AOI21_X1 U15884 ( .B1(n13925), .B2(n13923), .A(n13922), .ZN(n14091) );
  OAI211_X1 U15885 ( .C1(n13926), .C2(n13925), .A(n14376), .B(n13924), .ZN(
        n14089) );
  AOI21_X1 U15886 ( .B1(n13942), .B2(n14088), .A(n10341), .ZN(n13928) );
  AND2_X1 U15887 ( .A1(n13928), .A2(n13927), .ZN(n14086) );
  AOI22_X1 U15888 ( .A1(n14086), .A2(n13930), .B1(n14538), .B2(n13929), .ZN(
        n13931) );
  AOI21_X1 U15889 ( .B1(n14089), .B2(n13931), .A(n14539), .ZN(n13932) );
  INV_X1 U15890 ( .A(n13932), .ZN(n13937) );
  AOI22_X1 U15891 ( .A1(n13960), .A2(n13933), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n14539), .ZN(n13934) );
  OAI21_X1 U15892 ( .B1(n14085), .B2(n13966), .A(n13934), .ZN(n13935) );
  AOI21_X1 U15893 ( .B1(n14088), .B2(n14382), .A(n13935), .ZN(n13936) );
  OAI211_X1 U15894 ( .C1(n14091), .C2(n14009), .A(n13937), .B(n13936), .ZN(
        P1_U3272) );
  OAI211_X1 U15895 ( .C1(n13939), .C2(n13947), .A(n13938), .B(n14376), .ZN(
        n13941) );
  NAND2_X1 U15896 ( .A1(n13941), .A2(n13940), .ZN(n14098) );
  OAI211_X1 U15897 ( .C1(n6743), .C2(n14096), .A(n14559), .B(n13942), .ZN(
        n14094) );
  OAI22_X1 U15898 ( .A1(n14094), .A2(n13944), .B1(n13962), .B2(n13943), .ZN(
        n13945) );
  OAI21_X1 U15899 ( .B1(n14098), .B2(n13945), .A(n14006), .ZN(n13951) );
  AOI22_X1 U15900 ( .A1(n13946), .A2(n14382), .B1(P1_REG2_REG_20__SCAN_IN), 
        .B2(n14539), .ZN(n13950) );
  NAND2_X1 U15901 ( .A1(n13948), .A2(n13947), .ZN(n14092) );
  NAND3_X1 U15902 ( .A1(n14093), .A2(n14092), .A3(n14390), .ZN(n13949) );
  NAND3_X1 U15903 ( .A1(n13951), .A2(n13950), .A3(n13949), .ZN(P1_U3273) );
  XNOR2_X1 U15904 ( .A(n13952), .B(n13954), .ZN(n14109) );
  OAI21_X1 U15905 ( .B1(n13955), .B2(n13954), .A(n13953), .ZN(n14101) );
  INV_X1 U15906 ( .A(n13956), .ZN(n14011) );
  NAND2_X1 U15907 ( .A1(n14106), .A2(n13980), .ZN(n13957) );
  NAND2_X1 U15908 ( .A1(n13957), .A2(n14559), .ZN(n13958) );
  NOR2_X1 U15909 ( .A1(n6743), .A2(n13958), .ZN(n14104) );
  NAND2_X1 U15910 ( .A1(n14104), .A2(n14548), .ZN(n13969) );
  NAND2_X1 U15911 ( .A1(n13960), .A2(n13959), .ZN(n13965) );
  NOR2_X1 U15912 ( .A1(n13962), .A2(n13961), .ZN(n13963) );
  AOI21_X1 U15913 ( .B1(n14539), .B2(P1_REG2_REG_19__SCAN_IN), .A(n13963), 
        .ZN(n13964) );
  OAI211_X1 U15914 ( .C1(n14103), .C2(n13966), .A(n13965), .B(n13964), .ZN(
        n13967) );
  AOI21_X1 U15915 ( .B1(n14106), .B2(n14382), .A(n13967), .ZN(n13968) );
  NAND2_X1 U15916 ( .A1(n13969), .A2(n13968), .ZN(n13970) );
  AOI21_X1 U15917 ( .B1(n14101), .B2(n14011), .A(n13970), .ZN(n13971) );
  OAI21_X1 U15918 ( .B1(n14009), .B2(n14109), .A(n13971), .ZN(P1_U3274) );
  XNOR2_X1 U15919 ( .A(n13973), .B(n13972), .ZN(n14114) );
  OAI211_X1 U15920 ( .C1(n13976), .C2(n13975), .A(n13974), .B(n14376), .ZN(
        n13978) );
  OAI211_X1 U15921 ( .C1(n14114), .C2(n14602), .A(n13978), .B(n13977), .ZN(
        n13979) );
  INV_X1 U15922 ( .A(n13979), .ZN(n14113) );
  INV_X1 U15923 ( .A(n14000), .ZN(n13982) );
  INV_X1 U15924 ( .A(n13980), .ZN(n13981) );
  AOI21_X1 U15925 ( .B1(n14110), .B2(n13982), .A(n13981), .ZN(n14111) );
  AOI22_X1 U15926 ( .A1(n14539), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n13983), 
        .B2(n14538), .ZN(n13984) );
  OAI21_X1 U15927 ( .B1(n13985), .B2(n14541), .A(n13984), .ZN(n13988) );
  NOR2_X1 U15928 ( .A1(n14114), .A2(n13986), .ZN(n13987) );
  AOI211_X1 U15929 ( .C1(n14111), .C2(n14014), .A(n13988), .B(n13987), .ZN(
        n13989) );
  OAI21_X1 U15930 ( .B1(n14113), .B2(n14539), .A(n13989), .ZN(P1_U3275) );
  XNOR2_X1 U15931 ( .A(n13990), .B(n9755), .ZN(n14119) );
  AOI21_X1 U15932 ( .B1(n13992), .B2(n13991), .A(n14533), .ZN(n13996) );
  OAI22_X1 U15933 ( .A1(n14102), .A2(n14408), .B1(n13993), .B2(n14410), .ZN(
        n13994) );
  AOI21_X1 U15934 ( .B1(n13996), .B2(n13995), .A(n13994), .ZN(n14118) );
  INV_X1 U15935 ( .A(n14118), .ZN(n14007) );
  INV_X1 U15936 ( .A(n14116), .ZN(n14004) );
  NAND2_X1 U15937 ( .A1(n13997), .A2(n14116), .ZN(n13998) );
  NAND2_X1 U15938 ( .A1(n13998), .A2(n14559), .ZN(n13999) );
  NOR2_X1 U15939 ( .A1(n14000), .A2(n13999), .ZN(n14115) );
  NAND2_X1 U15940 ( .A1(n14115), .A2(n14548), .ZN(n14003) );
  AOI22_X1 U15941 ( .A1(n14539), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n14001), 
        .B2(n14538), .ZN(n14002) );
  OAI211_X1 U15942 ( .C1(n14004), .C2(n14541), .A(n14003), .B(n14002), .ZN(
        n14005) );
  AOI21_X1 U15943 ( .B1(n14007), .B2(n14006), .A(n14005), .ZN(n14008) );
  OAI21_X1 U15944 ( .B1(n14009), .B2(n14119), .A(n14008), .ZN(P1_U3276) );
  OAI21_X1 U15945 ( .B1(n14011), .B2(n14390), .A(n14010), .ZN(n14018) );
  AOI22_X1 U15946 ( .A1(n14552), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n14538), .ZN(n14017) );
  NAND2_X1 U15947 ( .A1(n14012), .A2(n10359), .ZN(n14016) );
  OAI21_X1 U15948 ( .B1(n14382), .B2(n14014), .A(n14013), .ZN(n14015) );
  NAND4_X1 U15949 ( .A1(n14018), .A2(n14017), .A3(n14016), .A4(n14015), .ZN(
        P1_U3293) );
  NAND2_X1 U15950 ( .A1(n14019), .A2(n14635), .ZN(n14020) );
  OAI211_X1 U15951 ( .C1(n14021), .C2(n10341), .A(n14020), .B(n14022), .ZN(
        n14122) );
  MUX2_X1 U15952 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14122), .S(n14665), .Z(
        P1_U3559) );
  OAI211_X1 U15953 ( .C1(n14626), .C2(n14024), .A(n14023), .B(n14022), .ZN(
        n14123) );
  MUX2_X1 U15954 ( .A(n14123), .B(P1_REG1_REG_30__SCAN_IN), .S(n14662), .Z(
        P1_U3558) );
  OAI21_X1 U15955 ( .B1(n14039), .B2(n14410), .A(n14025), .ZN(n14027) );
  AOI22_X1 U15956 ( .A1(n14617), .A2(n14031), .B1(n14047), .B2(n14634), .ZN(
        n14032) );
  OAI211_X1 U15957 ( .C1(n14034), .C2(n14626), .A(n14033), .B(n14032), .ZN(
        n14035) );
  OAI21_X1 U15958 ( .B1(n14037), .B2(n14533), .A(n14036), .ZN(n14125) );
  MUX2_X1 U15959 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14125), .S(n14665), .Z(
        P1_U3556) );
  OAI22_X1 U15960 ( .A1(n14039), .A2(n14408), .B1(n14038), .B2(n14410), .ZN(
        n14041) );
  AOI211_X1 U15961 ( .C1(n14042), .C2(n14635), .A(n14041), .B(n14040), .ZN(
        n14043) );
  OAI211_X1 U15962 ( .C1(n14563), .C2(n14045), .A(n14044), .B(n14043), .ZN(
        n14126) );
  MUX2_X1 U15963 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14126), .S(n14665), .Z(
        P1_U3555) );
  AOI22_X1 U15964 ( .A1(n14617), .A2(n14047), .B1(n14046), .B2(n14634), .ZN(
        n14048) );
  OAI211_X1 U15965 ( .C1(n14050), .C2(n14626), .A(n14049), .B(n14048), .ZN(
        n14051) );
  INV_X1 U15966 ( .A(n14051), .ZN(n14055) );
  NAND3_X1 U15967 ( .A1(n14053), .A2(n14642), .A3(n14052), .ZN(n14054) );
  OAI211_X1 U15968 ( .C1(n14056), .C2(n14533), .A(n14055), .B(n14054), .ZN(
        n14127) );
  MUX2_X1 U15969 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14127), .S(n14665), .Z(
        P1_U3554) );
  AOI22_X1 U15970 ( .A1(n14058), .A2(n14559), .B1(n14057), .B2(n14635), .ZN(
        n14062) );
  NAND3_X1 U15971 ( .A1(n14060), .A2(n14642), .A3(n14059), .ZN(n14061) );
  NAND3_X1 U15972 ( .A1(n14063), .A2(n14062), .A3(n14061), .ZN(n14128) );
  MUX2_X1 U15973 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14128), .S(n14665), .Z(
        P1_U3553) );
  INV_X1 U15974 ( .A(n14064), .ZN(n14069) );
  AOI21_X1 U15975 ( .B1(n14066), .B2(n14635), .A(n14065), .ZN(n14067) );
  OAI211_X1 U15976 ( .C1(n14069), .C2(n14601), .A(n14068), .B(n14067), .ZN(
        n14129) );
  MUX2_X1 U15977 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14129), .S(n14665), .Z(
        P1_U3552) );
  OAI21_X1 U15978 ( .B1(n14071), .B2(n14626), .A(n14070), .ZN(n14072) );
  AOI21_X1 U15979 ( .B1(n14073), .B2(n14642), .A(n14072), .ZN(n14074) );
  NAND2_X1 U15980 ( .A1(n14075), .A2(n14074), .ZN(n14130) );
  MUX2_X1 U15981 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14130), .S(n14665), .Z(
        P1_U3551) );
  AOI22_X1 U15982 ( .A1(n14077), .A2(n14617), .B1(n14634), .B2(n14076), .ZN(
        n14078) );
  OAI211_X1 U15983 ( .C1(n14626), .C2(n14080), .A(n14079), .B(n14078), .ZN(
        n14082) );
  AOI211_X1 U15984 ( .C1(n14642), .C2(n14083), .A(n14082), .B(n14081), .ZN(
        n14084) );
  INV_X1 U15985 ( .A(n14084), .ZN(n14131) );
  MUX2_X1 U15986 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14131), .S(n14665), .Z(
        P1_U3550) );
  OAI22_X1 U15987 ( .A1(n14103), .A2(n14410), .B1(n14085), .B2(n14408), .ZN(
        n14087) );
  AOI211_X1 U15988 ( .C1(n14088), .C2(n14635), .A(n14087), .B(n14086), .ZN(
        n14090) );
  OAI211_X1 U15989 ( .C1(n14091), .C2(n14563), .A(n14090), .B(n14089), .ZN(
        n14132) );
  MUX2_X1 U15990 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14132), .S(n14665), .Z(
        P1_U3549) );
  INV_X1 U15991 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n14099) );
  NAND3_X1 U15992 ( .A1(n14093), .A2(n14642), .A3(n14092), .ZN(n14095) );
  OAI211_X1 U15993 ( .C1(n14096), .C2(n14626), .A(n14095), .B(n14094), .ZN(
        n14097) );
  NOR2_X1 U15994 ( .A1(n14098), .A2(n14097), .ZN(n14133) );
  MUX2_X1 U15995 ( .A(n14099), .B(n14133), .S(n14665), .Z(n14100) );
  INV_X1 U15996 ( .A(n14100), .ZN(P1_U3548) );
  NAND2_X1 U15997 ( .A1(n14101), .A2(n14376), .ZN(n14108) );
  OAI22_X1 U15998 ( .A1(n14103), .A2(n14408), .B1(n14102), .B2(n14410), .ZN(
        n14105) );
  AOI211_X1 U15999 ( .C1(n14106), .C2(n14635), .A(n14105), .B(n14104), .ZN(
        n14107) );
  OAI211_X1 U16000 ( .C1(n14563), .C2(n14109), .A(n14108), .B(n14107), .ZN(
        n14135) );
  MUX2_X1 U16001 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14135), .S(n14665), .Z(
        P1_U3547) );
  AOI22_X1 U16002 ( .A1(n14111), .A2(n14559), .B1(n14110), .B2(n14635), .ZN(
        n14112) );
  OAI211_X1 U16003 ( .C1(n14114), .C2(n14601), .A(n14113), .B(n14112), .ZN(
        n14136) );
  MUX2_X1 U16004 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14136), .S(n14665), .Z(
        P1_U3546) );
  AOI21_X1 U16005 ( .B1(n14116), .B2(n14635), .A(n14115), .ZN(n14117) );
  OAI211_X1 U16006 ( .C1(n14563), .C2(n14119), .A(n14118), .B(n14117), .ZN(
        n14137) );
  MUX2_X1 U16007 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14137), .S(n14665), .Z(
        P1_U3545) );
  MUX2_X1 U16008 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14122), .S(n14645), .Z(
        P1_U3527) );
  MUX2_X1 U16009 ( .A(n14123), .B(P1_REG0_REG_30__SCAN_IN), .S(n14643), .Z(
        P1_U3526) );
  MUX2_X1 U16010 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14124), .S(n14645), .Z(
        P1_U3525) );
  MUX2_X1 U16011 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14125), .S(n14645), .Z(
        P1_U3524) );
  MUX2_X1 U16012 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14126), .S(n14645), .Z(
        P1_U3523) );
  MUX2_X1 U16013 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14127), .S(n14645), .Z(
        P1_U3522) );
  MUX2_X1 U16014 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14128), .S(n14645), .Z(
        P1_U3521) );
  MUX2_X1 U16015 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14129), .S(n14645), .Z(
        P1_U3520) );
  MUX2_X1 U16016 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14130), .S(n14645), .Z(
        P1_U3519) );
  MUX2_X1 U16017 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14131), .S(n14645), .Z(
        P1_U3518) );
  MUX2_X1 U16018 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14132), .S(n14645), .Z(
        P1_U3517) );
  MUX2_X1 U16019 ( .A(n15390), .B(n14133), .S(n14645), .Z(n14134) );
  INV_X1 U16020 ( .A(n14134), .ZN(P1_U3516) );
  MUX2_X1 U16021 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14135), .S(n14645), .Z(
        P1_U3515) );
  MUX2_X1 U16022 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14136), .S(n14645), .Z(
        P1_U3513) );
  MUX2_X1 U16023 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14137), .S(n14645), .Z(
        P1_U3510) );
  NOR4_X1 U16024 ( .A1(n14139), .A2(P1_IR_REG_30__SCAN_IN), .A3(n14138), .A4(
        P1_U3086), .ZN(n14140) );
  AOI21_X1 U16025 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n14141), .A(n14140), 
        .ZN(n14142) );
  OAI21_X1 U16026 ( .B1(n14143), .B2(n14160), .A(n14142), .ZN(P1_U3324) );
  OAI222_X1 U16027 ( .A1(n14146), .A2(P1_U3086), .B1(n14160), .B2(n14145), 
        .C1(n14144), .C2(n7001), .ZN(P1_U3326) );
  OAI222_X1 U16028 ( .A1(n7001), .A2(n14148), .B1(n14160), .B2(n14147), .C1(
        n9721), .C2(P1_U3086), .ZN(P1_U3327) );
  INV_X1 U16029 ( .A(n14149), .ZN(n14151) );
  OAI222_X1 U16030 ( .A1(n7001), .A2(n15324), .B1(n14160), .B2(n14151), .C1(
        P1_U3086), .C2(n14150), .ZN(P1_U3328) );
  OAI222_X1 U16031 ( .A1(n7001), .A2(n14154), .B1(n14160), .B2(n14153), .C1(
        n14152), .C2(P1_U3086), .ZN(P1_U3329) );
  OAI222_X1 U16032 ( .A1(n7001), .A2(n14157), .B1(n14160), .B2(n14156), .C1(
        P1_U3086), .C2(n14155), .ZN(P1_U3330) );
  OAI222_X1 U16033 ( .A1(n7001), .A2(n14161), .B1(n14160), .B2(n14159), .C1(
        n14158), .C2(P1_U3086), .ZN(P1_U3331) );
  MUX2_X1 U16034 ( .A(n9879), .B(n14162), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16035 ( .A(n14163), .B(n6762), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  INV_X1 U16036 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14463) );
  NAND2_X1 U16037 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14264), .ZN(n14265) );
  OAI21_X1 U16038 ( .B1(n14264), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n14265), 
        .ZN(n14198) );
  INV_X1 U16039 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14484) );
  NOR2_X1 U16040 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14484), .ZN(n14197) );
  INV_X1 U16041 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14164) );
  NOR2_X1 U16042 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n14164), .ZN(n14195) );
  INV_X1 U16043 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14193) );
  INV_X1 U16044 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14191) );
  INV_X1 U16045 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14165) );
  XOR2_X1 U16046 ( .A(n14165), .B(n14188), .Z(n14200) );
  INV_X1 U16047 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14953) );
  XNOR2_X1 U16048 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n14203) );
  INV_X1 U16049 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n15267) );
  XNOR2_X1 U16050 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n14209) );
  NAND2_X1 U16051 ( .A1(n14210), .A2(n14209), .ZN(n14166) );
  NAND2_X1 U16052 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14167), .ZN(n14170) );
  NAND2_X1 U16053 ( .A1(n14216), .A2(n14168), .ZN(n14169) );
  NAND2_X1 U16054 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14171), .ZN(n14172) );
  NAND2_X1 U16055 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14173), .ZN(n14175) );
  INV_X1 U16056 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14918) );
  NAND2_X1 U16057 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n14918), .ZN(n14176) );
  INV_X1 U16058 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n14178) );
  NAND2_X1 U16059 ( .A1(n14179), .A2(n14178), .ZN(n14181) );
  XNOR2_X1 U16060 ( .A(n14179), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n14231) );
  NAND2_X1 U16061 ( .A1(n14231), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14180) );
  NAND2_X1 U16062 ( .A1(n14181), .A2(n14180), .ZN(n14204) );
  XNOR2_X1 U16063 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n14239) );
  XNOR2_X1 U16064 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(P3_ADDR_REG_10__SCAN_IN), 
        .ZN(n14201) );
  NAND2_X1 U16065 ( .A1(n14202), .A2(n14201), .ZN(n14185) );
  INV_X1 U16066 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14189) );
  XOR2_X1 U16067 ( .A(n14189), .B(n14191), .Z(n14248) );
  AND2_X1 U16068 ( .A1(n14193), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14192) );
  INV_X1 U16069 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14194) );
  OAI22_X1 U16070 ( .A1(n14195), .A2(n14256), .B1(P3_ADDR_REG_14__SCAN_IN), 
        .B2(n14194), .ZN(n14258) );
  OAI22_X1 U16071 ( .A1(n14197), .A2(n14258), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n14196), .ZN(n14266) );
  XOR2_X1 U16072 ( .A(n14198), .B(n14266), .Z(n14461) );
  INV_X1 U16073 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n15237) );
  XNOR2_X1 U16074 ( .A(n14200), .B(n14199), .ZN(n14443) );
  XOR2_X1 U16075 ( .A(n14202), .B(n14201), .Z(n14284) );
  XOR2_X1 U16076 ( .A(n14204), .B(n14203), .Z(n14236) );
  XNOR2_X1 U16077 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n14205), .ZN(n14206) );
  NAND2_X1 U16078 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14206), .ZN(n14221) );
  INV_X1 U16079 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n15225) );
  XNOR2_X1 U16080 ( .A(n14206), .B(n15225), .ZN(n15516) );
  INV_X1 U16081 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14277) );
  XNOR2_X1 U16082 ( .A(n14208), .B(n14207), .ZN(n14275) );
  XNOR2_X1 U16083 ( .A(n14210), .B(n14209), .ZN(n14212) );
  NAND2_X1 U16084 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14212), .ZN(n14214) );
  AOI21_X1 U16085 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14211), .A(n14210), .ZN(
        n15519) );
  INV_X1 U16086 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15518) );
  NOR2_X1 U16087 ( .A1(n15519), .A2(n15518), .ZN(n15526) );
  NAND2_X1 U16088 ( .A1(n14275), .A2(n14276), .ZN(n14215) );
  NOR2_X1 U16089 ( .A1(n14275), .A2(n14276), .ZN(n14274) );
  XOR2_X1 U16090 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14216), .Z(n14218) );
  NOR2_X1 U16091 ( .A1(n14217), .A2(n14218), .ZN(n15522) );
  NOR2_X1 U16092 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(n15523), .ZN(n14219) );
  NAND2_X1 U16093 ( .A1(n14221), .A2(n14220), .ZN(n14224) );
  XNOR2_X1 U16094 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n14222), .ZN(n14223) );
  NOR2_X1 U16095 ( .A1(n14224), .A2(n14223), .ZN(n14226) );
  XNOR2_X1 U16096 ( .A(n14224), .B(n14223), .ZN(n15517) );
  NOR2_X1 U16097 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n15517), .ZN(n14225) );
  NAND2_X1 U16098 ( .A1(n14227), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14230) );
  XNOR2_X1 U16099 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n14229) );
  XNOR2_X1 U16100 ( .A(n14229), .B(n14228), .ZN(n14279) );
  NAND2_X1 U16101 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14232), .ZN(n14234) );
  XOR2_X1 U16102 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14231), .Z(n15521) );
  NAND2_X1 U16103 ( .A1(n14234), .A2(n14233), .ZN(n14235) );
  NOR2_X1 U16104 ( .A1(n14236), .A2(n14235), .ZN(n14238) );
  XNOR2_X1 U16105 ( .A(n14236), .B(n14235), .ZN(n14281) );
  NOR2_X1 U16106 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n14281), .ZN(n14237) );
  XNOR2_X1 U16107 ( .A(n14240), .B(n14239), .ZN(n14242) );
  NAND2_X1 U16108 ( .A1(n14241), .A2(n14242), .ZN(n14243) );
  NOR2_X1 U16109 ( .A1(n14284), .A2(n14285), .ZN(n14245) );
  INV_X1 U16110 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14244) );
  NAND2_X1 U16111 ( .A1(n14284), .A2(n14285), .ZN(n14283) );
  NOR2_X1 U16112 ( .A1(n14443), .A2(n14442), .ZN(n14247) );
  INV_X1 U16113 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14246) );
  NAND2_X1 U16114 ( .A1(n14443), .A2(n14442), .ZN(n14441) );
  XNOR2_X1 U16115 ( .A(n14249), .B(n14248), .ZN(n14447) );
  NAND2_X1 U16116 ( .A1(n14446), .A2(n14447), .ZN(n14250) );
  NOR2_X1 U16117 ( .A1(n14446), .A2(n14447), .ZN(n14445) );
  AOI21_X1 U16118 ( .B1(n14448), .B2(n14250), .A(n14445), .ZN(n14251) );
  INV_X1 U16119 ( .A(n14251), .ZN(n14255) );
  XOR2_X1 U16120 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n14252) );
  XOR2_X1 U16121 ( .A(n14253), .B(n14252), .Z(n14254) );
  XNOR2_X1 U16122 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n14257) );
  XNOR2_X1 U16123 ( .A(n14257), .B(n14256), .ZN(n14455) );
  XNOR2_X1 U16124 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n14259) );
  XOR2_X1 U16125 ( .A(n14259), .B(n14258), .Z(n14261) );
  NOR2_X1 U16126 ( .A1(n14260), .A2(n14261), .ZN(n14458) );
  NOR2_X2 U16127 ( .A1(n14458), .A2(n14262), .ZN(n14462) );
  NAND2_X1 U16128 ( .A1(n14461), .A2(n14462), .ZN(n14263) );
  NOR2_X1 U16129 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14264), .ZN(n14267) );
  OAI21_X1 U16130 ( .B1(n14267), .B2(n14266), .A(n14265), .ZN(n14268) );
  XOR2_X1 U16131 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14268), .Z(n14269) );
  XNOR2_X1 U16132 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14269), .ZN(n14317) );
  INV_X1 U16133 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14740) );
  NOR2_X1 U16134 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14268), .ZN(n14271) );
  AND2_X1 U16135 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14269), .ZN(n14270) );
  NOR2_X1 U16136 ( .A1(n14271), .A2(n14270), .ZN(n14325) );
  XOR2_X1 U16137 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n14324) );
  XNOR2_X1 U16138 ( .A(n14325), .B(n14324), .ZN(n14320) );
  XNOR2_X1 U16139 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14319), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16140 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14272) );
  OAI21_X1 U16141 ( .B1(P1_WR_REG_SCAN_IN), .B2(P2_WR_REG_SCAN_IN), .A(n14272), 
        .ZN(U28) );
  AOI21_X1 U16142 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14273) );
  OAI21_X1 U16143 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14273), 
        .ZN(U29) );
  AOI21_X1 U16144 ( .B1(n14276), .B2(n14275), .A(n14274), .ZN(n14278) );
  XNOR2_X1 U16145 ( .A(n14278), .B(n14277), .ZN(SUB_1596_U61) );
  XOR2_X1 U16146 ( .A(n14280), .B(n14279), .Z(SUB_1596_U57) );
  XNOR2_X1 U16147 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14281), .ZN(SUB_1596_U55)
         );
  XOR2_X1 U16148 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14282), .Z(SUB_1596_U54) );
  OAI21_X1 U16149 ( .B1(n14285), .B2(n14284), .A(n14283), .ZN(n14286) );
  XNOR2_X1 U16150 ( .A(n14286), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  INV_X1 U16151 ( .A(n14287), .ZN(n14297) );
  NOR2_X1 U16152 ( .A1(n14287), .A2(n14601), .ZN(n14296) );
  AOI22_X1 U16153 ( .A1(n14617), .A2(n14289), .B1(n14288), .B2(n14634), .ZN(
        n14293) );
  NAND2_X1 U16154 ( .A1(n14290), .A2(n14635), .ZN(n14291) );
  NAND4_X1 U16155 ( .A1(n14294), .A2(n14293), .A3(n14292), .A4(n14291), .ZN(
        n14295) );
  AOI211_X1 U16156 ( .C1(n14536), .C2(n14297), .A(n14296), .B(n14295), .ZN(
        n14300) );
  INV_X1 U16157 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14298) );
  AOI22_X1 U16158 ( .A1(n14645), .A2(n14300), .B1(n14298), .B2(n14643), .ZN(
        P1_U3495) );
  AOI22_X1 U16159 ( .A1(n14665), .A2(n14300), .B1(n14299), .B2(n14662), .ZN(
        P1_U3540) );
  OAI211_X1 U16160 ( .C1(n14303), .C2(n14302), .A(n14301), .B(n14376), .ZN(
        n14305) );
  AND2_X1 U16161 ( .A1(n14305), .A2(n14304), .ZN(n14422) );
  AOI222_X1 U16162 ( .A1(n14310), .A2(n14382), .B1(n14306), .B2(n14538), .C1(
        P1_REG2_REG_13__SCAN_IN), .C2(n14539), .ZN(n14315) );
  XNOR2_X1 U16163 ( .A(n14308), .B(n14307), .ZN(n14425) );
  INV_X1 U16164 ( .A(n14309), .ZN(n14312) );
  INV_X1 U16165 ( .A(n14310), .ZN(n14423) );
  OAI211_X1 U16166 ( .C1(n14312), .C2(n14423), .A(n14559), .B(n14311), .ZN(
        n14421) );
  INV_X1 U16167 ( .A(n14421), .ZN(n14313) );
  AOI22_X1 U16168 ( .A1(n14425), .A2(n14390), .B1(n14548), .B2(n14313), .ZN(
        n14314) );
  OAI211_X1 U16169 ( .C1(n14552), .C2(n14422), .A(n14315), .B(n14314), .ZN(
        P1_U3280) );
  OAI21_X1 U16170 ( .B1(n14317), .B2(n6732), .A(n14316), .ZN(n14318) );
  XNOR2_X1 U16171 ( .A(n14318), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  NOR2_X1 U16172 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n14319), .ZN(n14323) );
  NOR2_X1 U16173 ( .A1(n14321), .A2(n14320), .ZN(n14322) );
  INV_X1 U16174 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15248) );
  NOR2_X1 U16175 ( .A1(n14325), .A2(n14324), .ZN(n14326) );
  AOI21_X1 U16176 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n15248), .A(n14326), 
        .ZN(n14329) );
  XNOR2_X1 U16177 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14327) );
  XOR2_X1 U16178 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(n14327), .Z(n14328) );
  XNOR2_X1 U16179 ( .A(n14329), .B(n14328), .ZN(n14330) );
  XNOR2_X1 U16180 ( .A(n14331), .B(n14330), .ZN(SUB_1596_U4) );
  XNOR2_X1 U16181 ( .A(n14332), .B(n14337), .ZN(n14335) );
  AOI222_X1 U16182 ( .A1(n8938), .A2(n14335), .B1(n14334), .B2(n15059), .C1(
        n14333), .C2(n15062), .ZN(n14350) );
  AOI22_X1 U16183 ( .A1(n15071), .A2(n14336), .B1(n15056), .B2(
        P3_REG2_REG_12__SCAN_IN), .ZN(n14342) );
  XNOR2_X1 U16184 ( .A(n14338), .B(n14337), .ZN(n14353) );
  NOR2_X1 U16185 ( .A1(n14339), .A2(n15103), .ZN(n14352) );
  AOI22_X1 U16186 ( .A1(n14353), .A2(n14340), .B1(n15034), .B2(n14352), .ZN(
        n14341) );
  OAI211_X1 U16187 ( .C1(n15056), .C2(n14350), .A(n14342), .B(n14341), .ZN(
        P3_U3221) );
  OR2_X1 U16188 ( .A1(n14343), .A2(n15103), .ZN(n14344) );
  AOI22_X1 U16189 ( .A1(n15132), .A2(n14354), .B1(n9109), .B2(n15130), .ZN(
        P3_U3490) );
  NAND2_X1 U16190 ( .A1(n14346), .A2(n14345), .ZN(n14347) );
  AOI22_X1 U16191 ( .A1(n15132), .A2(n14356), .B1(n14349), .B2(n15130), .ZN(
        P3_U3489) );
  INV_X1 U16192 ( .A(n14350), .ZN(n14351) );
  AOI211_X1 U16193 ( .C1(n14353), .C2(n15101), .A(n14352), .B(n14351), .ZN(
        n14359) );
  AOI22_X1 U16194 ( .A1(n15132), .A2(n14359), .B1(n7769), .B2(n15130), .ZN(
        P3_U3471) );
  INV_X1 U16195 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14355) );
  AOI22_X1 U16196 ( .A1(n8156), .A2(n14355), .B1(n14354), .B2(n15119), .ZN(
        P3_U3458) );
  INV_X1 U16197 ( .A(n14356), .ZN(n14357) );
  OAI22_X1 U16198 ( .A1(n15119), .A2(P3_REG0_REG_30__SCAN_IN), .B1(n14357), 
        .B2(n8156), .ZN(n14358) );
  INV_X1 U16199 ( .A(n14358), .ZN(P3_U3457) );
  INV_X1 U16200 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14360) );
  AOI22_X1 U16201 ( .A1(n8156), .A2(n14360), .B1(n14359), .B2(n15119), .ZN(
        P3_U3426) );
  OAI211_X1 U16202 ( .C1(n14362), .C2(n14367), .A(n14361), .B(n14376), .ZN(
        n14364) );
  AOI222_X1 U16203 ( .A1(n14366), .A2(n14382), .B1(n14365), .B2(n14538), .C1(
        P1_REG2_REG_15__SCAN_IN), .C2(n14539), .ZN(n14375) );
  INV_X1 U16204 ( .A(n14367), .ZN(n14369) );
  OAI21_X1 U16205 ( .B1(n14370), .B2(n14369), .A(n14368), .ZN(n14406) );
  OAI211_X1 U16206 ( .C1(n14402), .C2(n14372), .A(n14559), .B(n14371), .ZN(
        n14401) );
  INV_X1 U16207 ( .A(n14401), .ZN(n14373) );
  AOI22_X1 U16208 ( .A1(n14406), .A2(n14390), .B1(n14548), .B2(n14373), .ZN(
        n14374) );
  OAI211_X1 U16209 ( .C1(n14552), .C2(n14403), .A(n14375), .B(n14374), .ZN(
        P1_U3278) );
  OAI211_X1 U16210 ( .C1(n14378), .C2(n7358), .A(n14377), .B(n14376), .ZN(
        n14380) );
  AND2_X1 U16211 ( .A1(n14380), .A2(n14379), .ZN(n14427) );
  AOI222_X1 U16212 ( .A1(n14383), .A2(n14382), .B1(n14381), .B2(n14538), .C1(
        P1_REG2_REG_11__SCAN_IN), .C2(n14539), .ZN(n14392) );
  XNOR2_X1 U16213 ( .A(n14385), .B(n14384), .ZN(n14430) );
  INV_X1 U16214 ( .A(n14386), .ZN(n14387) );
  OAI211_X1 U16215 ( .C1(n14428), .C2(n14388), .A(n14387), .B(n14559), .ZN(
        n14426) );
  INV_X1 U16216 ( .A(n14426), .ZN(n14389) );
  AOI22_X1 U16217 ( .A1(n14430), .A2(n14390), .B1(n14548), .B2(n14389), .ZN(
        n14391) );
  OAI211_X1 U16218 ( .C1(n14552), .C2(n14427), .A(n14392), .B(n14391), .ZN(
        P1_U3282) );
  AOI22_X1 U16219 ( .A1(n14394), .A2(n14617), .B1(n14634), .B2(n14393), .ZN(
        n14395) );
  OAI211_X1 U16220 ( .C1(n14397), .C2(n14626), .A(n14396), .B(n14395), .ZN(
        n14399) );
  AOI211_X1 U16221 ( .C1(n14400), .C2(n14642), .A(n14399), .B(n14398), .ZN(
        n14432) );
  AOI22_X1 U16222 ( .A1(n14665), .A2(n14432), .B1(n9553), .B2(n14662), .ZN(
        P1_U3544) );
  OAI21_X1 U16223 ( .B1(n14402), .B2(n14626), .A(n14401), .ZN(n14405) );
  INV_X1 U16224 ( .A(n14403), .ZN(n14404) );
  AOI211_X1 U16225 ( .C1(n14642), .C2(n14406), .A(n14405), .B(n14404), .ZN(
        n14434) );
  INV_X1 U16226 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14407) );
  AOI22_X1 U16227 ( .A1(n14665), .A2(n14434), .B1(n14407), .B2(n14662), .ZN(
        P1_U3543) );
  OAI22_X1 U16228 ( .A1(n14411), .A2(n14410), .B1(n14409), .B2(n14408), .ZN(
        n14413) );
  AOI211_X1 U16229 ( .C1(n14414), .C2(n14635), .A(n14413), .B(n14412), .ZN(
        n14419) );
  NAND3_X1 U16230 ( .A1(n14416), .A2(n14415), .A3(n14642), .ZN(n14417) );
  AOI22_X1 U16231 ( .A1(n14665), .A2(n14436), .B1(n14420), .B2(n14662), .ZN(
        P1_U3542) );
  OAI211_X1 U16232 ( .C1(n14423), .C2(n14626), .A(n14422), .B(n14421), .ZN(
        n14424) );
  AOI21_X1 U16233 ( .B1(n14425), .B2(n14642), .A(n14424), .ZN(n14438) );
  AOI22_X1 U16234 ( .A1(n14665), .A2(n14438), .B1(n10818), .B2(n14662), .ZN(
        P1_U3541) );
  OAI211_X1 U16235 ( .C1(n14428), .C2(n14626), .A(n14427), .B(n14426), .ZN(
        n14429) );
  AOI21_X1 U16236 ( .B1(n14430), .B2(n14642), .A(n14429), .ZN(n14440) );
  AOI22_X1 U16237 ( .A1(n14665), .A2(n14440), .B1(n14431), .B2(n14662), .ZN(
        P1_U3539) );
  AOI22_X1 U16238 ( .A1(n14645), .A2(n14432), .B1(n9556), .B2(n14643), .ZN(
        P1_U3507) );
  INV_X1 U16239 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14433) );
  AOI22_X1 U16240 ( .A1(n14645), .A2(n14434), .B1(n14433), .B2(n14643), .ZN(
        P1_U3504) );
  INV_X1 U16241 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14435) );
  AOI22_X1 U16242 ( .A1(n14645), .A2(n14436), .B1(n14435), .B2(n14643), .ZN(
        P1_U3501) );
  INV_X1 U16243 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14437) );
  AOI22_X1 U16244 ( .A1(n14645), .A2(n14438), .B1(n14437), .B2(n14643), .ZN(
        P1_U3498) );
  INV_X1 U16245 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14439) );
  AOI22_X1 U16246 ( .A1(n14645), .A2(n14440), .B1(n14439), .B2(n14643), .ZN(
        P1_U3492) );
  OAI21_X1 U16247 ( .B1(n14443), .B2(n14442), .A(n14441), .ZN(n14444) );
  XNOR2_X1 U16248 ( .A(n14444), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  AOI21_X1 U16249 ( .B1(n14447), .B2(n14446), .A(n14445), .ZN(n14449) );
  XNOR2_X1 U16250 ( .A(n14449), .B(n14448), .ZN(SUB_1596_U68) );
  NOR2_X1 U16251 ( .A1(n14451), .A2(n14450), .ZN(n14452) );
  XOR2_X1 U16252 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n14452), .Z(SUB_1596_U67)
         );
  AOI21_X1 U16253 ( .B1(n14455), .B2(n14454), .A(n14453), .ZN(n14456) );
  XNOR2_X1 U16254 ( .A(n14456), .B(n15237), .ZN(SUB_1596_U66) );
  NOR2_X1 U16255 ( .A1(n14458), .A2(n14457), .ZN(n14459) );
  XOR2_X1 U16256 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14459), .Z(SUB_1596_U65)
         );
  AOI21_X1 U16257 ( .B1(n14462), .B2(n14461), .A(n14460), .ZN(n14464) );
  XNOR2_X1 U16258 ( .A(n14464), .B(n14463), .ZN(SUB_1596_U64) );
  OAI21_X1 U16259 ( .B1(n14466), .B2(P1_REG1_REG_0__SCAN_IN), .A(n14465), .ZN(
        n14467) );
  XOR2_X1 U16260 ( .A(n6762), .B(n14467), .Z(n14471) );
  AOI22_X1 U16261 ( .A1(n14468), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14469) );
  OAI21_X1 U16262 ( .B1(n14471), .B2(n14470), .A(n14469), .ZN(P1_U3243) );
  AOI21_X1 U16263 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n14473), .A(n14472), 
        .ZN(n14478) );
  AOI21_X1 U16264 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14475), .A(n14474), 
        .ZN(n14476) );
  OAI222_X1 U16265 ( .A1(n14494), .A2(n14480), .B1(n14479), .B2(n14478), .C1(
        n14477), .C2(n14476), .ZN(n14481) );
  INV_X1 U16266 ( .A(n14481), .ZN(n14483) );
  OAI211_X1 U16267 ( .C1(n14484), .C2(n14498), .A(n14483), .B(n14482), .ZN(
        P1_U3258) );
  OAI211_X1 U16268 ( .C1(n14487), .C2(P1_REG1_REG_18__SCAN_IN), .A(n14486), 
        .B(n14485), .ZN(n14492) );
  OAI211_X1 U16269 ( .C1(n14490), .C2(P1_REG2_REG_18__SCAN_IN), .A(n14489), 
        .B(n14488), .ZN(n14491) );
  OAI211_X1 U16270 ( .C1(n14494), .C2(n14493), .A(n14492), .B(n14491), .ZN(
        n14495) );
  INV_X1 U16271 ( .A(n14495), .ZN(n14497) );
  OAI211_X1 U16272 ( .C1(n15248), .C2(n14498), .A(n14497), .B(n14496), .ZN(
        P1_U3261) );
  XNOR2_X1 U16273 ( .A(n14500), .B(n14499), .ZN(n14613) );
  XNOR2_X1 U16274 ( .A(n14501), .B(n14502), .ZN(n14504) );
  OAI21_X1 U16275 ( .B1(n14504), .B2(n14533), .A(n14503), .ZN(n14505) );
  AOI21_X1 U16276 ( .B1(n14536), .B2(n14613), .A(n14505), .ZN(n14610) );
  AOI22_X1 U16277 ( .A1(n14539), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n14506), 
        .B2(n14538), .ZN(n14507) );
  OAI21_X1 U16278 ( .B1(n14541), .B2(n14609), .A(n14507), .ZN(n14508) );
  INV_X1 U16279 ( .A(n14508), .ZN(n14513) );
  OAI211_X1 U16280 ( .C1(n14510), .C2(n14609), .A(n14559), .B(n14509), .ZN(
        n14608) );
  INV_X1 U16281 ( .A(n14608), .ZN(n14511) );
  AOI22_X1 U16282 ( .A1(n14613), .A2(n14549), .B1(n14548), .B2(n14511), .ZN(
        n14512) );
  OAI211_X1 U16283 ( .C1(n14552), .C2(n14610), .A(n14513), .B(n14512), .ZN(
        P1_U3286) );
  XNOR2_X1 U16284 ( .A(n14516), .B(n14514), .ZN(n14598) );
  XNOR2_X1 U16285 ( .A(n14516), .B(n14515), .ZN(n14517) );
  NOR2_X1 U16286 ( .A1(n14517), .A2(n14533), .ZN(n14518) );
  AOI211_X1 U16287 ( .C1(n14536), .C2(n14598), .A(n14519), .B(n14518), .ZN(
        n14595) );
  AOI22_X1 U16288 ( .A1(n14539), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n14520), 
        .B2(n14538), .ZN(n14521) );
  OAI21_X1 U16289 ( .B1(n14541), .B2(n14594), .A(n14521), .ZN(n14522) );
  INV_X1 U16290 ( .A(n14522), .ZN(n14528) );
  INV_X1 U16291 ( .A(n14523), .ZN(n14525) );
  OAI211_X1 U16292 ( .C1(n14525), .C2(n14594), .A(n14559), .B(n14524), .ZN(
        n14593) );
  INV_X1 U16293 ( .A(n14593), .ZN(n14526) );
  AOI22_X1 U16294 ( .A1(n14598), .A2(n14549), .B1(n14548), .B2(n14526), .ZN(
        n14527) );
  OAI211_X1 U16295 ( .C1(n14552), .C2(n14595), .A(n14528), .B(n14527), .ZN(
        P1_U3288) );
  XNOR2_X1 U16296 ( .A(n14529), .B(n14531), .ZN(n14580) );
  XNOR2_X1 U16297 ( .A(n14530), .B(n14531), .ZN(n14534) );
  OAI21_X1 U16298 ( .B1(n14534), .B2(n14533), .A(n14532), .ZN(n14535) );
  AOI21_X1 U16299 ( .B1(n14536), .B2(n14580), .A(n14535), .ZN(n14577) );
  AOI22_X1 U16300 ( .A1(n14539), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n14538), 
        .B2(n14537), .ZN(n14540) );
  OAI21_X1 U16301 ( .B1(n14541), .B2(n14576), .A(n14540), .ZN(n14542) );
  INV_X1 U16302 ( .A(n14542), .ZN(n14551) );
  INV_X1 U16303 ( .A(n14543), .ZN(n14546) );
  INV_X1 U16304 ( .A(n14544), .ZN(n14545) );
  OAI211_X1 U16305 ( .C1(n14576), .C2(n14546), .A(n14545), .B(n14559), .ZN(
        n14575) );
  INV_X1 U16306 ( .A(n14575), .ZN(n14547) );
  AOI22_X1 U16307 ( .A1(n14580), .A2(n14549), .B1(n14548), .B2(n14547), .ZN(
        n14550) );
  OAI211_X1 U16308 ( .C1(n14552), .C2(n14577), .A(n14551), .B(n14550), .ZN(
        P1_U3290) );
  AND2_X1 U16309 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15133), .ZN(P1_U3294) );
  AND2_X1 U16310 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15133), .ZN(P1_U3295) );
  AND2_X1 U16311 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15133), .ZN(P1_U3296) );
  AND2_X1 U16312 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15133), .ZN(P1_U3297) );
  AND2_X1 U16313 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15133), .ZN(P1_U3298) );
  NOR2_X1 U16314 ( .A1(n14555), .A2(n14553), .ZN(P1_U3299) );
  INV_X1 U16315 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n15240) );
  NOR2_X1 U16316 ( .A1(n14555), .A2(n15240), .ZN(P1_U3300) );
  NOR2_X1 U16317 ( .A1(n14555), .A2(n15286), .ZN(P1_U3301) );
  AND2_X1 U16318 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15133), .ZN(P1_U3303) );
  AND2_X1 U16319 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15133), .ZN(P1_U3304) );
  AND2_X1 U16320 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15133), .ZN(P1_U3305) );
  AND2_X1 U16321 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15133), .ZN(P1_U3306) );
  AND2_X1 U16322 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15133), .ZN(P1_U3307) );
  AND2_X1 U16323 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15133), .ZN(P1_U3308) );
  INV_X1 U16324 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n15328) );
  NOR2_X1 U16325 ( .A1(n14555), .A2(n15328), .ZN(P1_U3309) );
  AND2_X1 U16326 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15133), .ZN(P1_U3310) );
  INV_X1 U16327 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n15374) );
  NOR2_X1 U16328 ( .A1(n14555), .A2(n15374), .ZN(P1_U3311) );
  AND2_X1 U16329 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15133), .ZN(P1_U3312) );
  AND2_X1 U16330 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15133), .ZN(P1_U3313) );
  AND2_X1 U16331 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15133), .ZN(P1_U3314) );
  AND2_X1 U16332 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15133), .ZN(P1_U3315) );
  AND2_X1 U16333 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15133), .ZN(P1_U3316) );
  AND2_X1 U16334 ( .A1(n15133), .A2(P1_D_REG_8__SCAN_IN), .ZN(P1_U3317) );
  INV_X1 U16335 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15407) );
  NOR2_X1 U16336 ( .A1(n14555), .A2(n15407), .ZN(P1_U3318) );
  NOR2_X1 U16337 ( .A1(n14555), .A2(n14554), .ZN(P1_U3319) );
  AND2_X1 U16338 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15133), .ZN(P1_U3320) );
  INV_X1 U16339 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15420) );
  NOR2_X1 U16340 ( .A1(n14555), .A2(n15420), .ZN(P1_U3321) );
  AND2_X1 U16341 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15133), .ZN(P1_U3322) );
  INV_X1 U16342 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n15405) );
  NOR2_X1 U16343 ( .A1(n14555), .A2(n15405), .ZN(P1_U3323) );
  INV_X1 U16344 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n14556) );
  AOI22_X1 U16345 ( .A1(n14645), .A2(n14557), .B1(n14556), .B2(n14643), .ZN(
        P1_U3459) );
  AOI22_X1 U16346 ( .A1(n14617), .A2(n9894), .B1(n14635), .B2(n14558), .ZN(
        n14562) );
  NAND2_X1 U16347 ( .A1(n14560), .A2(n14559), .ZN(n14561) );
  OAI211_X1 U16348 ( .C1(n14564), .C2(n14563), .A(n14562), .B(n14561), .ZN(
        n14566) );
  NOR2_X1 U16349 ( .A1(n14566), .A2(n14565), .ZN(n14646) );
  INV_X1 U16350 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14567) );
  AOI22_X1 U16351 ( .A1(n14645), .A2(n14646), .B1(n14567), .B2(n14643), .ZN(
        P1_U3462) );
  INV_X1 U16352 ( .A(n14601), .ZN(n14631) );
  OAI21_X1 U16353 ( .B1(n14569), .B2(n14626), .A(n14568), .ZN(n14572) );
  INV_X1 U16354 ( .A(n14570), .ZN(n14571) );
  AOI211_X1 U16355 ( .C1(n14631), .C2(n14573), .A(n14572), .B(n14571), .ZN(
        n14647) );
  INV_X1 U16356 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14574) );
  AOI22_X1 U16357 ( .A1(n14645), .A2(n14647), .B1(n14574), .B2(n14643), .ZN(
        P1_U3465) );
  OAI21_X1 U16358 ( .B1(n14576), .B2(n14626), .A(n14575), .ZN(n14579) );
  INV_X1 U16359 ( .A(n14577), .ZN(n14578) );
  AOI211_X1 U16360 ( .C1(n14631), .C2(n14580), .A(n14579), .B(n14578), .ZN(
        n14649) );
  INV_X1 U16361 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n14581) );
  AOI22_X1 U16362 ( .A1(n14645), .A2(n14649), .B1(n14581), .B2(n14643), .ZN(
        P1_U3468) );
  INV_X1 U16363 ( .A(n14582), .ZN(n14591) );
  AOI22_X1 U16364 ( .A1(n14617), .A2(n14584), .B1(n14583), .B2(n14634), .ZN(
        n14588) );
  NAND2_X1 U16365 ( .A1(n14585), .A2(n14635), .ZN(n14586) );
  NAND4_X1 U16366 ( .A1(n14589), .A2(n14588), .A3(n14587), .A4(n14586), .ZN(
        n14590) );
  AOI21_X1 U16367 ( .B1(n14591), .B2(n14642), .A(n14590), .ZN(n14651) );
  INV_X1 U16368 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14592) );
  AOI22_X1 U16369 ( .A1(n14645), .A2(n14651), .B1(n14592), .B2(n14643), .ZN(
        P1_U3471) );
  OAI21_X1 U16370 ( .B1(n14594), .B2(n14626), .A(n14593), .ZN(n14597) );
  INV_X1 U16371 ( .A(n14595), .ZN(n14596) );
  AOI211_X1 U16372 ( .C1(n14631), .C2(n14598), .A(n14597), .B(n14596), .ZN(
        n14653) );
  INV_X1 U16373 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14599) );
  AOI22_X1 U16374 ( .A1(n14645), .A2(n14653), .B1(n14599), .B2(n14643), .ZN(
        P1_U3474) );
  AOI21_X1 U16375 ( .B1(n14602), .B2(n14601), .A(n14600), .ZN(n14606) );
  NOR2_X1 U16376 ( .A1(n7323), .A2(n14626), .ZN(n14604) );
  NOR4_X1 U16377 ( .A1(n14606), .A2(n14605), .A3(n14604), .A4(n14603), .ZN(
        n14655) );
  INV_X1 U16378 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14607) );
  AOI22_X1 U16379 ( .A1(n14645), .A2(n14655), .B1(n14607), .B2(n14643), .ZN(
        P1_U3477) );
  OAI21_X1 U16380 ( .B1(n14609), .B2(n14626), .A(n14608), .ZN(n14612) );
  INV_X1 U16381 ( .A(n14610), .ZN(n14611) );
  AOI211_X1 U16382 ( .C1(n14631), .C2(n14613), .A(n14612), .B(n14611), .ZN(
        n14657) );
  INV_X1 U16383 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14614) );
  AOI22_X1 U16384 ( .A1(n14645), .A2(n14657), .B1(n14614), .B2(n14643), .ZN(
        P1_U3480) );
  INV_X1 U16385 ( .A(n14615), .ZN(n14623) );
  AOI22_X1 U16386 ( .A1(n14633), .A2(n14617), .B1(n14634), .B2(n14616), .ZN(
        n14618) );
  OAI211_X1 U16387 ( .C1(n7219), .C2(n14626), .A(n14619), .B(n14618), .ZN(
        n14622) );
  INV_X1 U16388 ( .A(n14620), .ZN(n14621) );
  AOI211_X1 U16389 ( .C1(n14642), .C2(n14623), .A(n14622), .B(n14621), .ZN(
        n14659) );
  INV_X1 U16390 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14624) );
  AOI22_X1 U16391 ( .A1(n14645), .A2(n14659), .B1(n14624), .B2(n14643), .ZN(
        P1_U3483) );
  OAI21_X1 U16392 ( .B1(n14627), .B2(n14626), .A(n14625), .ZN(n14629) );
  AOI211_X1 U16393 ( .C1(n14631), .C2(n14630), .A(n14629), .B(n14628), .ZN(
        n14661) );
  INV_X1 U16394 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14632) );
  AOI22_X1 U16395 ( .A1(n14645), .A2(n14661), .B1(n14632), .B2(n14643), .ZN(
        P1_U3486) );
  AOI22_X1 U16396 ( .A1(n14636), .A2(n14635), .B1(n14634), .B2(n14633), .ZN(
        n14637) );
  NAND2_X1 U16397 ( .A1(n14638), .A2(n14637), .ZN(n14640) );
  AOI211_X1 U16398 ( .C1(n14642), .C2(n14641), .A(n14640), .B(n14639), .ZN(
        n14664) );
  INV_X1 U16399 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14644) );
  AOI22_X1 U16400 ( .A1(n14645), .A2(n14664), .B1(n14644), .B2(n14643), .ZN(
        P1_U3489) );
  AOI22_X1 U16401 ( .A1(n14665), .A2(n14646), .B1(n10416), .B2(n14662), .ZN(
        P1_U3529) );
  AOI22_X1 U16402 ( .A1(n14665), .A2(n14647), .B1(n10415), .B2(n14662), .ZN(
        P1_U3530) );
  AOI22_X1 U16403 ( .A1(n14665), .A2(n14649), .B1(n14648), .B2(n14662), .ZN(
        P1_U3531) );
  AOI22_X1 U16404 ( .A1(n14665), .A2(n14651), .B1(n14650), .B2(n14662), .ZN(
        P1_U3532) );
  AOI22_X1 U16405 ( .A1(n14665), .A2(n14653), .B1(n14652), .B2(n14662), .ZN(
        P1_U3533) );
  AOI22_X1 U16406 ( .A1(n14665), .A2(n14655), .B1(n14654), .B2(n14662), .ZN(
        P1_U3534) );
  AOI22_X1 U16407 ( .A1(n14665), .A2(n14657), .B1(n14656), .B2(n14662), .ZN(
        P1_U3535) );
  INV_X1 U16408 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n14658) );
  AOI22_X1 U16409 ( .A1(n14665), .A2(n14659), .B1(n14658), .B2(n14662), .ZN(
        P1_U3536) );
  AOI22_X1 U16410 ( .A1(n14665), .A2(n14661), .B1(n14660), .B2(n14662), .ZN(
        P1_U3537) );
  AOI22_X1 U16411 ( .A1(n14665), .A2(n14664), .B1(n14663), .B2(n14662), .ZN(
        P1_U3538) );
  NOR2_X1 U16412 ( .A1(n14726), .A2(P2_U3947), .ZN(P2_U3087) );
  OAI22_X1 U16413 ( .A1(n14741), .A2(n6771), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8257), .ZN(n14666) );
  AOI21_X1 U16414 ( .B1(n14667), .B2(n14750), .A(n14666), .ZN(n14676) );
  OAI211_X1 U16415 ( .C1(n14670), .C2(n14669), .A(n14752), .B(n14668), .ZN(
        n14675) );
  OAI211_X1 U16416 ( .C1(n14673), .C2(n14672), .A(n14729), .B(n14671), .ZN(
        n14674) );
  NAND3_X1 U16417 ( .A1(n14676), .A2(n14675), .A3(n14674), .ZN(P2_U3215) );
  INV_X1 U16418 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n14677) );
  OAI22_X1 U16419 ( .A1(n14741), .A2(n14677), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8290), .ZN(n14678) );
  AOI21_X1 U16420 ( .B1(n14679), .B2(n14750), .A(n14678), .ZN(n14688) );
  OAI211_X1 U16421 ( .C1(n14682), .C2(n14681), .A(n14752), .B(n14680), .ZN(
        n14687) );
  OAI211_X1 U16422 ( .C1(n14685), .C2(n14684), .A(n14729), .B(n14683), .ZN(
        n14686) );
  NAND3_X1 U16423 ( .A1(n14688), .A2(n14687), .A3(n14686), .ZN(P2_U3217) );
  NOR2_X1 U16424 ( .A1(n14722), .A2(n14689), .ZN(n14690) );
  AOI211_X1 U16425 ( .C1(n14726), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n14691), 
        .B(n14690), .ZN(n14702) );
  AOI21_X1 U16426 ( .B1(n14693), .B2(n14692), .A(n14745), .ZN(n14695) );
  NAND2_X1 U16427 ( .A1(n14695), .A2(n14694), .ZN(n14701) );
  AOI211_X1 U16428 ( .C1(n14698), .C2(n14697), .A(n14718), .B(n14696), .ZN(
        n14699) );
  INV_X1 U16429 ( .A(n14699), .ZN(n14700) );
  NAND3_X1 U16430 ( .A1(n14702), .A2(n14701), .A3(n14700), .ZN(P2_U3227) );
  XOR2_X1 U16431 ( .A(n14704), .B(n14703), .Z(n14708) );
  OAI21_X1 U16432 ( .B1(n14722), .B2(n14706), .A(n14705), .ZN(n14707) );
  AOI21_X1 U16433 ( .B1(n14708), .B2(n14752), .A(n14707), .ZN(n14712) );
  OAI211_X1 U16434 ( .C1(n14710), .C2(P2_REG2_REG_14__SCAN_IN), .A(n14729), 
        .B(n14709), .ZN(n14711) );
  OAI211_X1 U16435 ( .C1(n14741), .C2(n15237), .A(n14712), .B(n14711), .ZN(
        P2_U3228) );
  OAI211_X1 U16436 ( .C1(n14714), .C2(P2_REG2_REG_15__SCAN_IN), .A(n14729), 
        .B(n14713), .ZN(n14720) );
  OAI21_X1 U16437 ( .B1(n14716), .B2(P2_REG1_REG_15__SCAN_IN), .A(n14715), 
        .ZN(n14717) );
  OR2_X1 U16438 ( .A1(n14718), .A2(n14717), .ZN(n14719) );
  OAI211_X1 U16439 ( .C1(n14722), .C2(n14721), .A(n14720), .B(n14719), .ZN(
        n14723) );
  AOI211_X1 U16440 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n14726), .A(n14724), 
        .B(n14723), .ZN(n14725) );
  INV_X1 U16441 ( .A(n14725), .ZN(P2_U3229) );
  AOI22_X1 U16442 ( .A1(n14726), .A2(P2_ADDR_REG_16__SCAN_IN), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(P2_U3088), .ZN(n14738) );
  NAND2_X1 U16443 ( .A1(n14750), .A2(n14727), .ZN(n14737) );
  OAI211_X1 U16444 ( .C1(n14731), .C2(n14730), .A(n14729), .B(n14728), .ZN(
        n14736) );
  OAI211_X1 U16445 ( .C1(n14734), .C2(n14733), .A(n14752), .B(n14732), .ZN(
        n14735) );
  NAND4_X1 U16446 ( .A1(n14738), .A2(n14737), .A3(n14736), .A4(n14735), .ZN(
        P2_U3230) );
  OAI21_X1 U16447 ( .B1(n14741), .B2(n14740), .A(n14739), .ZN(n14748) );
  OAI21_X1 U16448 ( .B1(n14744), .B2(n14743), .A(n14742), .ZN(n14746) );
  NOR2_X1 U16449 ( .A1(n14746), .A2(n14745), .ZN(n14747) );
  AOI211_X1 U16450 ( .C1(n14750), .C2(n14749), .A(n14748), .B(n14747), .ZN(
        n14756) );
  OAI211_X1 U16451 ( .C1(n14754), .C2(n14753), .A(n14752), .B(n14751), .ZN(
        n14755) );
  NAND2_X1 U16452 ( .A1(n14756), .A2(n14755), .ZN(P2_U3231) );
  NAND2_X1 U16453 ( .A1(n14758), .A2(n14757), .ZN(n14763) );
  AOI22_X1 U16454 ( .A1(n14761), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n14760), 
        .B2(n14759), .ZN(n14762) );
  OAI211_X1 U16455 ( .C1(n14765), .C2(n14764), .A(n14763), .B(n14762), .ZN(
        n14766) );
  AOI21_X1 U16456 ( .B1(n11149), .B2(n14767), .A(n14766), .ZN(n14768) );
  OAI21_X1 U16457 ( .B1(n14770), .B2(n14769), .A(n14768), .ZN(P2_U3258) );
  AND2_X1 U16458 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14778), .ZN(P2_U3266) );
  AND2_X1 U16459 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14778), .ZN(P2_U3267) );
  AND2_X1 U16460 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14778), .ZN(P2_U3268) );
  AND2_X1 U16461 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14778), .ZN(P2_U3269) );
  AND2_X1 U16462 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14778), .ZN(P2_U3270) );
  NOR2_X1 U16463 ( .A1(n14775), .A2(n15246), .ZN(P2_U3271) );
  AND2_X1 U16464 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14778), .ZN(P2_U3272) );
  AND2_X1 U16465 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14778), .ZN(P2_U3273) );
  AND2_X1 U16466 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14778), .ZN(P2_U3274) );
  AND2_X1 U16467 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14778), .ZN(P2_U3275) );
  AND2_X1 U16468 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14778), .ZN(P2_U3276) );
  NOR2_X1 U16469 ( .A1(n14775), .A2(n15355), .ZN(P2_U3277) );
  INV_X1 U16470 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15362) );
  NOR2_X1 U16471 ( .A1(n14775), .A2(n15362), .ZN(P2_U3278) );
  AND2_X1 U16472 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14778), .ZN(P2_U3279) );
  AND2_X1 U16473 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14778), .ZN(P2_U3280) );
  AND2_X1 U16474 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14778), .ZN(P2_U3281) );
  INV_X1 U16475 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15421) );
  NOR2_X1 U16476 ( .A1(n14775), .A2(n15421), .ZN(P2_U3282) );
  AND2_X1 U16477 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14778), .ZN(P2_U3283) );
  AND2_X1 U16478 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14778), .ZN(P2_U3284) );
  AND2_X1 U16479 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14778), .ZN(P2_U3285) );
  AND2_X1 U16480 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14778), .ZN(P2_U3286) );
  AND2_X1 U16481 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14778), .ZN(P2_U3287) );
  AND2_X1 U16482 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14778), .ZN(P2_U3288) );
  NOR2_X1 U16483 ( .A1(n14775), .A2(n14773), .ZN(P2_U3289) );
  AND2_X1 U16484 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14778), .ZN(P2_U3290) );
  AND2_X1 U16485 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14778), .ZN(P2_U3291) );
  AND2_X1 U16486 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14778), .ZN(P2_U3292) );
  AND2_X1 U16487 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14778), .ZN(P2_U3293) );
  AND2_X1 U16488 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14778), .ZN(P2_U3294) );
  NOR2_X1 U16489 ( .A1(n14775), .A2(n14774), .ZN(P2_U3295) );
  AOI22_X1 U16490 ( .A1(n14781), .A2(n14777), .B1(n14776), .B2(n14778), .ZN(
        P2_U3416) );
  AOI22_X1 U16491 ( .A1(n14781), .A2(n14780), .B1(n14779), .B2(n14778), .ZN(
        P2_U3417) );
  INV_X1 U16492 ( .A(n14822), .ZN(n14784) );
  OAI211_X1 U16493 ( .C1(n14785), .C2(n14784), .A(n14783), .B(n14782), .ZN(
        n14786) );
  INV_X1 U16494 ( .A(n14786), .ZN(n14830) );
  INV_X1 U16495 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14787) );
  AOI22_X1 U16496 ( .A1(n6621), .A2(n14830), .B1(n14787), .B2(n14829), .ZN(
        P2_U3430) );
  INV_X1 U16497 ( .A(n14794), .ZN(n14796) );
  INV_X1 U16498 ( .A(n14788), .ZN(n14789) );
  AOI211_X1 U16499 ( .C1(n14792), .C2(n14791), .A(n14790), .B(n14789), .ZN(
        n14793) );
  OAI21_X1 U16500 ( .B1(n14815), .B2(n14794), .A(n14793), .ZN(n14795) );
  AOI21_X1 U16501 ( .B1(n14822), .B2(n14796), .A(n14795), .ZN(n14831) );
  INV_X1 U16502 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n14797) );
  AOI22_X1 U16503 ( .A1(n6621), .A2(n14831), .B1(n14797), .B2(n14829), .ZN(
        P2_U3433) );
  OAI21_X1 U16504 ( .B1(n6770), .B2(n14826), .A(n14798), .ZN(n14801) );
  INV_X1 U16505 ( .A(n14799), .ZN(n14800) );
  AOI211_X1 U16506 ( .C1(n14802), .C2(n14808), .A(n14801), .B(n14800), .ZN(
        n14832) );
  INV_X1 U16507 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n14803) );
  AOI22_X1 U16508 ( .A1(n6621), .A2(n14832), .B1(n14803), .B2(n14829), .ZN(
        P2_U3436) );
  OAI21_X1 U16509 ( .B1(n7498), .B2(n14826), .A(n14804), .ZN(n14807) );
  INV_X1 U16510 ( .A(n14805), .ZN(n14806) );
  AOI211_X1 U16511 ( .C1(n14809), .C2(n14808), .A(n14807), .B(n14806), .ZN(
        n14833) );
  INV_X1 U16512 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14810) );
  AOI22_X1 U16513 ( .A1(n6621), .A2(n14833), .B1(n14810), .B2(n14829), .ZN(
        P2_U3439) );
  INV_X1 U16514 ( .A(n14816), .ZN(n14814) );
  OAI21_X1 U16515 ( .B1(n14812), .B2(n14826), .A(n14811), .ZN(n14813) );
  AOI21_X1 U16516 ( .B1(n14814), .B2(n14822), .A(n14813), .ZN(n14819) );
  OR2_X1 U16517 ( .A1(n14816), .A2(n14815), .ZN(n14817) );
  AND3_X1 U16518 ( .A1(n14819), .A2(n14818), .A3(n14817), .ZN(n14834) );
  INV_X1 U16519 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14820) );
  AOI22_X1 U16520 ( .A1(n6621), .A2(n14834), .B1(n14820), .B2(n14829), .ZN(
        P2_U3445) );
  NAND2_X1 U16521 ( .A1(n14823), .A2(n14822), .ZN(n14825) );
  OAI211_X1 U16522 ( .C1(n7072), .C2(n14826), .A(n14825), .B(n14824), .ZN(
        n14828) );
  NOR2_X1 U16523 ( .A1(n14828), .A2(n14827), .ZN(n14836) );
  INV_X1 U16524 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n15397) );
  AOI22_X1 U16525 ( .A1(n6621), .A2(n14836), .B1(n15397), .B2(n14829), .ZN(
        P2_U3448) );
  AOI22_X1 U16526 ( .A1(n14837), .A2(n14830), .B1(n10192), .B2(n14835), .ZN(
        P2_U3499) );
  AOI22_X1 U16527 ( .A1(n14837), .A2(n14831), .B1(n10211), .B2(n14835), .ZN(
        P2_U3500) );
  AOI22_X1 U16528 ( .A1(n14837), .A2(n14832), .B1(n10212), .B2(n14835), .ZN(
        P2_U3501) );
  AOI22_X1 U16529 ( .A1(n14837), .A2(n14833), .B1(n10223), .B2(n14835), .ZN(
        P2_U3502) );
  AOI22_X1 U16530 ( .A1(n14837), .A2(n14834), .B1(n10227), .B2(n14835), .ZN(
        P2_U3504) );
  AOI22_X1 U16531 ( .A1(n14837), .A2(n14836), .B1(n10230), .B2(n14835), .ZN(
        P2_U3505) );
  NOR2_X1 U16532 ( .A1(P3_U3897), .A2(n14978), .ZN(P3_U3150) );
  AND2_X1 U16533 ( .A1(n14838), .A2(n15036), .ZN(n14839) );
  NOR2_X1 U16534 ( .A1(n14866), .A2(n14839), .ZN(n14855) );
  INV_X1 U16535 ( .A(n14840), .ZN(n14841) );
  OAI21_X1 U16536 ( .B1(n14952), .B2(n7049), .A(n14841), .ZN(n14848) );
  INV_X1 U16537 ( .A(n14858), .ZN(n14846) );
  NAND3_X1 U16538 ( .A1(n14844), .A2(n14843), .A3(n14842), .ZN(n14845) );
  AOI21_X1 U16539 ( .B1(n14846), .B2(n14845), .A(n14986), .ZN(n14847) );
  AOI211_X1 U16540 ( .C1(n14915), .C2(n14849), .A(n14848), .B(n14847), .ZN(
        n14854) );
  XNOR2_X1 U16541 ( .A(n14851), .B(n14850), .ZN(n14852) );
  NAND2_X1 U16542 ( .A1(n14992), .A2(n14852), .ZN(n14853) );
  OAI211_X1 U16543 ( .C1(n14855), .C2(n14994), .A(n14854), .B(n14853), .ZN(
        P3_U3185) );
  INV_X1 U16544 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14879) );
  INV_X1 U16545 ( .A(n14887), .ZN(n14860) );
  NOR3_X1 U16546 ( .A1(n14858), .A2(n14857), .A3(n14856), .ZN(n14859) );
  OAI21_X1 U16547 ( .B1(n14860), .B2(n14859), .A(n14960), .ZN(n14874) );
  INV_X1 U16548 ( .A(n14861), .ZN(n14863) );
  NAND2_X1 U16549 ( .A1(n14863), .A2(n14862), .ZN(n14865) );
  OAI21_X1 U16550 ( .B1(n14866), .B2(n14865), .A(n14864), .ZN(n14871) );
  OAI21_X1 U16551 ( .B1(n14869), .B2(n14868), .A(n14867), .ZN(n14870) );
  AOI22_X1 U16552 ( .A1(n14872), .A2(n14871), .B1(n14992), .B2(n14870), .ZN(
        n14873) );
  OAI211_X1 U16553 ( .C1(n14982), .C2(n14875), .A(n14874), .B(n14873), .ZN(
        n14876) );
  INV_X1 U16554 ( .A(n14876), .ZN(n14878) );
  OAI211_X1 U16555 ( .C1(n14879), .C2(n14952), .A(n14878), .B(n14877), .ZN(
        P3_U3186) );
  AOI21_X1 U16556 ( .B1(n15023), .B2(n14881), .A(n14880), .ZN(n14898) );
  INV_X1 U16557 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n14884) );
  INV_X1 U16558 ( .A(n14882), .ZN(n14883) );
  OAI21_X1 U16559 ( .B1(n14952), .B2(n14884), .A(n14883), .ZN(n14891) );
  INV_X1 U16560 ( .A(n14910), .ZN(n14889) );
  NAND3_X1 U16561 ( .A1(n14887), .A2(n14886), .A3(n14885), .ZN(n14888) );
  AOI21_X1 U16562 ( .B1(n14889), .B2(n14888), .A(n14986), .ZN(n14890) );
  AOI211_X1 U16563 ( .C1(n14915), .C2(n14892), .A(n14891), .B(n14890), .ZN(
        n14897) );
  XNOR2_X1 U16564 ( .A(n14894), .B(n14893), .ZN(n14895) );
  NAND2_X1 U16565 ( .A1(n14992), .A2(n14895), .ZN(n14896) );
  OAI211_X1 U16566 ( .C1(n14898), .C2(n14994), .A(n14897), .B(n14896), .ZN(
        P3_U3187) );
  AOI21_X1 U16567 ( .B1(n14901), .B2(n14900), .A(n14899), .ZN(n14907) );
  OAI21_X1 U16568 ( .B1(n14904), .B2(n14903), .A(n14902), .ZN(n14905) );
  NAND2_X1 U16569 ( .A1(n14992), .A2(n14905), .ZN(n14906) );
  OAI21_X1 U16570 ( .B1(n14907), .B2(n14994), .A(n14906), .ZN(n14913) );
  OR3_X1 U16571 ( .A1(n14910), .A2(n14909), .A3(n14908), .ZN(n14911) );
  AOI21_X1 U16572 ( .B1(n14924), .B2(n14911), .A(n14986), .ZN(n14912) );
  AOI211_X1 U16573 ( .C1(n14915), .C2(n14914), .A(n14913), .B(n14912), .ZN(
        n14917) );
  OAI211_X1 U16574 ( .C1(n14918), .C2(n14952), .A(n14917), .B(n14916), .ZN(
        P3_U3188) );
  AOI21_X1 U16575 ( .B1(n14921), .B2(n14920), .A(n14919), .ZN(n14935) );
  AND3_X1 U16576 ( .A1(n14924), .A2(n14923), .A3(n14922), .ZN(n14925) );
  OAI21_X1 U16577 ( .B1(n14945), .B2(n14925), .A(n14960), .ZN(n14926) );
  OAI21_X1 U16578 ( .B1(n14982), .B2(n14927), .A(n14926), .ZN(n14928) );
  AOI211_X1 U16579 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n14978), .A(n14929), .B(
        n14928), .ZN(n14934) );
  OAI21_X1 U16580 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n14931), .A(n14930), .ZN(
        n14932) );
  NAND2_X1 U16581 ( .A1(n14992), .A2(n14932), .ZN(n14933) );
  OAI211_X1 U16582 ( .C1(n14935), .C2(n14994), .A(n14934), .B(n14933), .ZN(
        P3_U3189) );
  OAI21_X1 U16583 ( .B1(n14938), .B2(n14937), .A(n14936), .ZN(n14949) );
  AOI21_X1 U16584 ( .B1(n6754), .B2(n14940), .A(n14939), .ZN(n14941) );
  OAI22_X1 U16585 ( .A1(n14982), .A2(n14942), .B1(n14941), .B2(n14994), .ZN(
        n14948) );
  OR3_X1 U16586 ( .A1(n14945), .A2(n14944), .A3(n14943), .ZN(n14946) );
  AOI21_X1 U16587 ( .B1(n14959), .B2(n14946), .A(n14986), .ZN(n14947) );
  AOI211_X1 U16588 ( .C1(n14992), .C2(n14949), .A(n14948), .B(n14947), .ZN(
        n14951) );
  OAI211_X1 U16589 ( .C1(n14953), .C2(n14952), .A(n14951), .B(n14950), .ZN(
        P3_U3190) );
  AOI21_X1 U16590 ( .B1(n14956), .B2(n14955), .A(n14954), .ZN(n14971) );
  AND3_X1 U16591 ( .A1(n14959), .A2(n14958), .A3(n14957), .ZN(n14961) );
  OAI21_X1 U16592 ( .B1(n14985), .B2(n14961), .A(n14960), .ZN(n14962) );
  OAI21_X1 U16593 ( .B1(n14982), .B2(n14963), .A(n14962), .ZN(n14964) );
  AOI211_X1 U16594 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n14978), .A(n14965), .B(
        n14964), .ZN(n14970) );
  OAI21_X1 U16595 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n14967), .A(n14966), .ZN(
        n14968) );
  NAND2_X1 U16596 ( .A1(n14968), .A2(n14992), .ZN(n14969) );
  OAI211_X1 U16597 ( .C1(n14971), .C2(n14994), .A(n14970), .B(n14969), .ZN(
        P3_U3191) );
  AOI21_X1 U16598 ( .B1(n14974), .B2(n14973), .A(n14972), .ZN(n14995) );
  OAI21_X1 U16599 ( .B1(n14977), .B2(n14976), .A(n14975), .ZN(n14991) );
  NAND2_X1 U16600 ( .A1(n14978), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n14979) );
  OAI211_X1 U16601 ( .C1(n14982), .C2(n14981), .A(n14980), .B(n14979), .ZN(
        n14990) );
  OR3_X1 U16602 ( .A1(n14985), .A2(n14984), .A3(n14983), .ZN(n14987) );
  AOI21_X1 U16603 ( .B1(n14988), .B2(n14987), .A(n14986), .ZN(n14989) );
  AOI211_X1 U16604 ( .C1(n14992), .C2(n14991), .A(n14990), .B(n14989), .ZN(
        n14993) );
  OAI21_X1 U16605 ( .B1(n14995), .B2(n14994), .A(n14993), .ZN(P3_U3192) );
  XNOR2_X1 U16606 ( .A(n14996), .B(n14999), .ZN(n15005) );
  INV_X1 U16607 ( .A(n15005), .ZN(n15095) );
  INV_X1 U16608 ( .A(n14997), .ZN(n15068) );
  OAI211_X1 U16609 ( .C1(n15000), .C2(n14999), .A(n14998), .B(n8938), .ZN(
        n15004) );
  AOI22_X1 U16610 ( .A1(n15062), .A2(n15002), .B1(n15001), .B2(n15059), .ZN(
        n15003) );
  OAI211_X1 U16611 ( .C1(n15068), .C2(n15005), .A(n15004), .B(n15003), .ZN(
        n15093) );
  AOI21_X1 U16612 ( .B1(n15049), .B2(n15095), .A(n15093), .ZN(n15010) );
  NOR2_X1 U16613 ( .A1(n15006), .A2(n15103), .ZN(n15094) );
  AOI22_X1 U16614 ( .A1(n15034), .A2(n15094), .B1(n15071), .B2(n15007), .ZN(
        n15008) );
  OAI221_X1 U16615 ( .B1(n15056), .B2(n15010), .C1(n15074), .C2(n15009), .A(
        n15008), .ZN(P3_U3227) );
  OAI21_X1 U16616 ( .B1(n15012), .B2(n15014), .A(n15011), .ZN(n15092) );
  AOI21_X1 U16617 ( .B1(n15014), .B2(n11824), .A(n15013), .ZN(n15015) );
  OAI222_X1 U16618 ( .A1(n15043), .A2(n15018), .B1(n15045), .B2(n15017), .C1(
        n15016), .C2(n15015), .ZN(n15090) );
  AOI21_X1 U16619 ( .B1(n15019), .B2(n15092), .A(n15090), .ZN(n15024) );
  NOR2_X1 U16620 ( .A1(n15020), .A2(n15103), .ZN(n15091) );
  AOI22_X1 U16621 ( .A1(n15034), .A2(n15091), .B1(n15071), .B2(n15021), .ZN(
        n15022) );
  OAI221_X1 U16622 ( .B1(n15056), .B2(n15024), .C1(n15074), .C2(n15023), .A(
        n15022), .ZN(P3_U3228) );
  XNOR2_X1 U16623 ( .A(n15028), .B(n15025), .ZN(n15032) );
  INV_X1 U16624 ( .A(n15032), .ZN(n15084) );
  AOI22_X1 U16625 ( .A1(n15062), .A2(n15060), .B1(n15026), .B2(n15059), .ZN(
        n15031) );
  OAI211_X1 U16626 ( .C1(n15029), .C2(n15028), .A(n15027), .B(n8938), .ZN(
        n15030) );
  OAI211_X1 U16627 ( .C1(n15032), .C2(n15068), .A(n15031), .B(n15030), .ZN(
        n15082) );
  AOI21_X1 U16628 ( .B1(n15049), .B2(n15084), .A(n15082), .ZN(n15037) );
  NOR2_X1 U16629 ( .A1(n15033), .A2(n15103), .ZN(n15083) );
  AOI22_X1 U16630 ( .A1(n15034), .A2(n15083), .B1(n15071), .B2(n7604), .ZN(
        n15035) );
  OAI221_X1 U16631 ( .B1(n15056), .B2(n15037), .C1(n15074), .C2(n15036), .A(
        n15035), .ZN(P3_U3230) );
  OAI21_X1 U16632 ( .B1(n15039), .B2(n9133), .A(n15038), .ZN(n15081) );
  INV_X1 U16633 ( .A(n15081), .ZN(n15053) );
  OAI21_X1 U16634 ( .B1(n15042), .B2(n15041), .A(n15040), .ZN(n15047) );
  OAI22_X1 U16635 ( .A1(n7578), .A2(n15045), .B1(n15044), .B2(n15043), .ZN(
        n15046) );
  AOI21_X1 U16636 ( .B1(n15047), .B2(n8938), .A(n15046), .ZN(n15048) );
  OAI21_X1 U16637 ( .B1(n15053), .B2(n15068), .A(n15048), .ZN(n15079) );
  INV_X1 U16638 ( .A(n15049), .ZN(n15052) );
  NOR2_X1 U16639 ( .A1(n15050), .A2(n15103), .ZN(n15080) );
  INV_X1 U16640 ( .A(n15080), .ZN(n15051) );
  OAI22_X1 U16641 ( .A1(n15053), .A2(n15052), .B1(n15058), .B2(n15051), .ZN(
        n15054) );
  AOI211_X1 U16642 ( .C1(n15071), .C2(P3_REG3_REG_2__SCAN_IN), .A(n15079), .B(
        n15054), .ZN(n15055) );
  AOI22_X1 U16643 ( .A1(n15056), .A2(n10760), .B1(n15055), .B2(n15074), .ZN(
        P3_U3231) );
  NOR2_X1 U16644 ( .A1(n15057), .A2(n15103), .ZN(n15077) );
  INV_X1 U16645 ( .A(n15058), .ZN(n15069) );
  XNOR2_X1 U16646 ( .A(n9131), .B(n9130), .ZN(n15070) );
  AOI22_X1 U16647 ( .A1(n15062), .A2(n15061), .B1(n15060), .B2(n15059), .ZN(
        n15067) );
  OAI21_X1 U16648 ( .B1(n9130), .B2(n15064), .A(n15063), .ZN(n15065) );
  NAND2_X1 U16649 ( .A1(n15065), .A2(n8938), .ZN(n15066) );
  OAI211_X1 U16650 ( .C1(n15070), .C2(n15068), .A(n15067), .B(n15066), .ZN(
        n15076) );
  AOI21_X1 U16651 ( .B1(n15077), .B2(n15069), .A(n15076), .ZN(n15075) );
  INV_X1 U16652 ( .A(n15070), .ZN(n15078) );
  AOI22_X1 U16653 ( .A1(n15078), .A2(n15072), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15071), .ZN(n15073) );
  OAI221_X1 U16654 ( .B1(n15056), .B2(n15075), .C1(n15074), .C2(n10755), .A(
        n15073), .ZN(P3_U3232) );
  AOI211_X1 U16655 ( .C1(n15115), .C2(n15078), .A(n15077), .B(n15076), .ZN(
        n15121) );
  AOI22_X1 U16656 ( .A1(n8156), .A2(n7566), .B1(n15121), .B2(n15119), .ZN(
        P3_U3393) );
  INV_X1 U16657 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15296) );
  AOI211_X1 U16658 ( .C1(n15115), .C2(n15081), .A(n15080), .B(n15079), .ZN(
        n15122) );
  AOI22_X1 U16659 ( .A1(n8156), .A2(n15296), .B1(n15122), .B2(n15119), .ZN(
        P3_U3396) );
  INV_X1 U16660 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15085) );
  AOI211_X1 U16661 ( .C1(n15084), .C2(n15115), .A(n15083), .B(n15082), .ZN(
        n15123) );
  AOI22_X1 U16662 ( .A1(n8156), .A2(n15085), .B1(n15123), .B2(n15119), .ZN(
        P3_U3399) );
  INV_X1 U16663 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15381) );
  INV_X1 U16664 ( .A(n15086), .ZN(n15087) );
  AOI211_X1 U16665 ( .C1(n15089), .C2(n15115), .A(n15088), .B(n15087), .ZN(
        n15124) );
  AOI22_X1 U16666 ( .A1(n8156), .A2(n15381), .B1(n15124), .B2(n15119), .ZN(
        P3_U3402) );
  INV_X1 U16667 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15375) );
  AOI211_X1 U16668 ( .C1(n15101), .C2(n15092), .A(n15091), .B(n15090), .ZN(
        n15125) );
  AOI22_X1 U16669 ( .A1(n8156), .A2(n15375), .B1(n15125), .B2(n15119), .ZN(
        P3_U3405) );
  INV_X1 U16670 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15096) );
  AOI211_X1 U16671 ( .C1(n15095), .C2(n15115), .A(n15094), .B(n15093), .ZN(
        n15126) );
  AOI22_X1 U16672 ( .A1(n8156), .A2(n15096), .B1(n15126), .B2(n15119), .ZN(
        P3_U3408) );
  INV_X1 U16673 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15102) );
  NOR2_X1 U16674 ( .A1(n15097), .A2(n15103), .ZN(n15099) );
  AOI211_X1 U16675 ( .C1(n15101), .C2(n15100), .A(n15099), .B(n15098), .ZN(
        n15127) );
  AOI22_X1 U16676 ( .A1(n8156), .A2(n15102), .B1(n15127), .B2(n15119), .ZN(
        P3_U3411) );
  INV_X1 U16677 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15108) );
  NOR2_X1 U16678 ( .A1(n15104), .A2(n15103), .ZN(n15106) );
  AOI211_X1 U16679 ( .C1(n15115), .C2(n15107), .A(n15106), .B(n15105), .ZN(
        n15128) );
  AOI22_X1 U16680 ( .A1(n8156), .A2(n15108), .B1(n15128), .B2(n15119), .ZN(
        P3_U3414) );
  INV_X1 U16681 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15113) );
  AOI21_X1 U16682 ( .B1(n15110), .B2(n15115), .A(n15109), .ZN(n15111) );
  AND2_X1 U16683 ( .A1(n15112), .A2(n15111), .ZN(n15129) );
  AOI22_X1 U16684 ( .A1(n8156), .A2(n15113), .B1(n15129), .B2(n15119), .ZN(
        P3_U3417) );
  INV_X1 U16685 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15120) );
  AOI21_X1 U16686 ( .B1(n15116), .B2(n15115), .A(n15114), .ZN(n15117) );
  AND2_X1 U16687 ( .A1(n15118), .A2(n15117), .ZN(n15131) );
  AOI22_X1 U16688 ( .A1(n8156), .A2(n15120), .B1(n15131), .B2(n15119), .ZN(
        P3_U3420) );
  AOI22_X1 U16689 ( .A1(n15132), .A2(n15121), .B1(n10913), .B2(n15130), .ZN(
        P3_U3460) );
  AOI22_X1 U16690 ( .A1(n15132), .A2(n15122), .B1(n10759), .B2(n15130), .ZN(
        P3_U3461) );
  AOI22_X1 U16691 ( .A1(n15132), .A2(n15123), .B1(n14850), .B2(n15130), .ZN(
        P3_U3462) );
  AOI22_X1 U16692 ( .A1(n15132), .A2(n15124), .B1(n11429), .B2(n15130), .ZN(
        P3_U3463) );
  AOI22_X1 U16693 ( .A1(n15132), .A2(n15125), .B1(n14893), .B2(n15130), .ZN(
        P3_U3464) );
  AOI22_X1 U16694 ( .A1(n15132), .A2(n15126), .B1(n11396), .B2(n15130), .ZN(
        P3_U3465) );
  AOI22_X1 U16695 ( .A1(n15132), .A2(n15127), .B1(n11400), .B2(n15130), .ZN(
        P3_U3466) );
  AOI22_X1 U16696 ( .A1(n15132), .A2(n15128), .B1(n11436), .B2(n15130), .ZN(
        P3_U3467) );
  AOI22_X1 U16697 ( .A1(n15132), .A2(n15129), .B1(n11409), .B2(n15130), .ZN(
        P3_U3468) );
  AOI22_X1 U16698 ( .A1(n15132), .A2(n15131), .B1(n11440), .B2(n15130), .ZN(
        P3_U3469) );
  NAND2_X1 U16699 ( .A1(n15133), .A2(P1_D_REG_23__SCAN_IN), .ZN(n15514) );
  AOI22_X1 U16700 ( .A1(P1_D_REG_16__SCAN_IN), .A2(keyinput190), .B1(
        P3_REG3_REG_15__SCAN_IN), .B2(keyinput155), .ZN(n15134) );
  OAI221_X1 U16701 ( .B1(P1_D_REG_16__SCAN_IN), .B2(keyinput190), .C1(
        P3_REG3_REG_15__SCAN_IN), .C2(keyinput155), .A(n15134), .ZN(n15141) );
  AOI22_X1 U16702 ( .A1(P2_REG0_REG_7__SCAN_IN), .A2(keyinput252), .B1(
        P3_ADDR_REG_19__SCAN_IN), .B2(keyinput207), .ZN(n15135) );
  OAI221_X1 U16703 ( .B1(P2_REG0_REG_7__SCAN_IN), .B2(keyinput252), .C1(
        P3_ADDR_REG_19__SCAN_IN), .C2(keyinput207), .A(n15135), .ZN(n15140) );
  AOI22_X1 U16704 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(keyinput152), .B1(
        P3_D_REG_12__SCAN_IN), .B2(keyinput129), .ZN(n15136) );
  OAI221_X1 U16705 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(keyinput152), .C1(
        P3_D_REG_12__SCAN_IN), .C2(keyinput129), .A(n15136), .ZN(n15139) );
  AOI22_X1 U16706 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(keyinput202), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(keyinput158), .ZN(n15137) );
  OAI221_X1 U16707 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(keyinput202), .C1(
        P1_ADDR_REG_10__SCAN_IN), .C2(keyinput158), .A(n15137), .ZN(n15138) );
  NOR4_X1 U16708 ( .A1(n15141), .A2(n15140), .A3(n15139), .A4(n15138), .ZN(
        n15169) );
  AOI22_X1 U16709 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(keyinput171), .B1(
        P2_REG2_REG_1__SCAN_IN), .B2(keyinput144), .ZN(n15142) );
  OAI221_X1 U16710 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(keyinput171), .C1(
        P2_REG2_REG_1__SCAN_IN), .C2(keyinput144), .A(n15142), .ZN(n15149) );
  AOI22_X1 U16711 ( .A1(P2_D_REG_19__SCAN_IN), .A2(keyinput164), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(keyinput142), .ZN(n15143) );
  OAI221_X1 U16712 ( .B1(P2_D_REG_19__SCAN_IN), .B2(keyinput164), .C1(
        P2_DATAO_REG_2__SCAN_IN), .C2(keyinput142), .A(n15143), .ZN(n15148) );
  AOI22_X1 U16713 ( .A1(P2_REG2_REG_25__SCAN_IN), .A2(keyinput180), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(keyinput136), .ZN(n15144) );
  OAI221_X1 U16714 ( .B1(P2_REG2_REG_25__SCAN_IN), .B2(keyinput180), .C1(
        P2_DATAO_REG_25__SCAN_IN), .C2(keyinput136), .A(n15144), .ZN(n15147)
         );
  AOI22_X1 U16715 ( .A1(P1_D_REG_14__SCAN_IN), .A2(keyinput245), .B1(
        P2_IR_REG_5__SCAN_IN), .B2(keyinput221), .ZN(n15145) );
  OAI221_X1 U16716 ( .B1(P1_D_REG_14__SCAN_IN), .B2(keyinput245), .C1(
        P2_IR_REG_5__SCAN_IN), .C2(keyinput221), .A(n15145), .ZN(n15146) );
  NOR4_X1 U16717 ( .A1(n15149), .A2(n15148), .A3(n15147), .A4(n15146), .ZN(
        n15168) );
  AOI22_X1 U16718 ( .A1(P2_D_REG_2__SCAN_IN), .A2(keyinput206), .B1(
        P3_REG1_REG_18__SCAN_IN), .B2(keyinput232), .ZN(n15150) );
  OAI221_X1 U16719 ( .B1(P2_D_REG_2__SCAN_IN), .B2(keyinput206), .C1(
        P3_REG1_REG_18__SCAN_IN), .C2(keyinput232), .A(n15150), .ZN(n15157) );
  AOI22_X1 U16720 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput176), .B1(
        P3_REG1_REG_30__SCAN_IN), .B2(keyinput137), .ZN(n15151) );
  OAI221_X1 U16721 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput176), .C1(
        P3_REG1_REG_30__SCAN_IN), .C2(keyinput137), .A(n15151), .ZN(n15156) );
  AOI22_X1 U16722 ( .A1(P2_REG1_REG_30__SCAN_IN), .A2(keyinput216), .B1(
        P2_REG2_REG_2__SCAN_IN), .B2(keyinput241), .ZN(n15152) );
  OAI221_X1 U16723 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(keyinput216), .C1(
        P2_REG2_REG_2__SCAN_IN), .C2(keyinput241), .A(n15152), .ZN(n15155) );
  AOI22_X1 U16724 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(keyinput218), .B1(
        P1_REG0_REG_30__SCAN_IN), .B2(keyinput185), .ZN(n15153) );
  OAI221_X1 U16725 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(keyinput218), .C1(
        P1_REG0_REG_30__SCAN_IN), .C2(keyinput185), .A(n15153), .ZN(n15154) );
  NOR4_X1 U16726 ( .A1(n15157), .A2(n15156), .A3(n15155), .A4(n15154), .ZN(
        n15167) );
  AOI22_X1 U16727 ( .A1(P2_D_REG_15__SCAN_IN), .A2(keyinput244), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(keyinput191), .ZN(n15158) );
  OAI221_X1 U16728 ( .B1(P2_D_REG_15__SCAN_IN), .B2(keyinput244), .C1(
        P2_DATAO_REG_14__SCAN_IN), .C2(keyinput191), .A(n15158), .ZN(n15165)
         );
  AOI22_X1 U16729 ( .A1(P1_D_REG_26__SCAN_IN), .A2(keyinput146), .B1(
        P2_D_REG_20__SCAN_IN), .B2(keyinput224), .ZN(n15159) );
  OAI221_X1 U16730 ( .B1(P1_D_REG_26__SCAN_IN), .B2(keyinput146), .C1(
        P2_D_REG_20__SCAN_IN), .C2(keyinput224), .A(n15159), .ZN(n15164) );
  AOI22_X1 U16731 ( .A1(P3_REG0_REG_5__SCAN_IN), .A2(keyinput149), .B1(SI_17_), 
        .B2(keyinput173), .ZN(n15160) );
  OAI221_X1 U16732 ( .B1(P3_REG0_REG_5__SCAN_IN), .B2(keyinput149), .C1(SI_17_), .C2(keyinput173), .A(n15160), .ZN(n15163) );
  AOI22_X1 U16733 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(keyinput133), .B1(
        P3_REG2_REG_13__SCAN_IN), .B2(keyinput228), .ZN(n15161) );
  OAI221_X1 U16734 ( .B1(P2_IR_REG_10__SCAN_IN), .B2(keyinput133), .C1(
        P3_REG2_REG_13__SCAN_IN), .C2(keyinput228), .A(n15161), .ZN(n15162) );
  NOR4_X1 U16735 ( .A1(n15165), .A2(n15164), .A3(n15163), .A4(n15162), .ZN(
        n15166) );
  NAND4_X1 U16736 ( .A1(n15169), .A2(n15168), .A3(n15167), .A4(n15166), .ZN(
        n15314) );
  AOI22_X1 U16737 ( .A1(P1_D_REG_6__SCAN_IN), .A2(keyinput251), .B1(
        P3_D_REG_11__SCAN_IN), .B2(keyinput165), .ZN(n15170) );
  OAI221_X1 U16738 ( .B1(P1_D_REG_6__SCAN_IN), .B2(keyinput251), .C1(
        P3_D_REG_11__SCAN_IN), .C2(keyinput165), .A(n15170), .ZN(n15177) );
  AOI22_X1 U16739 ( .A1(P3_D_REG_2__SCAN_IN), .A2(keyinput179), .B1(
        P3_REG3_REG_5__SCAN_IN), .B2(keyinput255), .ZN(n15171) );
  OAI221_X1 U16740 ( .B1(P3_D_REG_2__SCAN_IN), .B2(keyinput179), .C1(
        P3_REG3_REG_5__SCAN_IN), .C2(keyinput255), .A(n15171), .ZN(n15176) );
  AOI22_X1 U16741 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(keyinput237), .B1(
        P2_REG1_REG_7__SCAN_IN), .B2(keyinput169), .ZN(n15172) );
  OAI221_X1 U16742 ( .B1(P1_IR_REG_21__SCAN_IN), .B2(keyinput237), .C1(
        P2_REG1_REG_7__SCAN_IN), .C2(keyinput169), .A(n15172), .ZN(n15175) );
  AOI22_X1 U16743 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput150), .B1(
        P3_D_REG_7__SCAN_IN), .B2(keyinput189), .ZN(n15173) );
  OAI221_X1 U16744 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput150), .C1(
        P3_D_REG_7__SCAN_IN), .C2(keyinput189), .A(n15173), .ZN(n15174) );
  NOR4_X1 U16745 ( .A1(n15177), .A2(n15176), .A3(n15175), .A4(n15174), .ZN(
        n15205) );
  AOI22_X1 U16746 ( .A1(P1_REG0_REG_19__SCAN_IN), .A2(keyinput223), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(keyinput242), .ZN(n15178) );
  OAI221_X1 U16747 ( .B1(P1_REG0_REG_19__SCAN_IN), .B2(keyinput223), .C1(
        P2_DATAO_REG_1__SCAN_IN), .C2(keyinput242), .A(n15178), .ZN(n15185) );
  AOI22_X1 U16748 ( .A1(P2_D_REG_8__SCAN_IN), .A2(keyinput174), .B1(
        P3_REG3_REG_9__SCAN_IN), .B2(keyinput187), .ZN(n15179) );
  OAI221_X1 U16749 ( .B1(P2_D_REG_8__SCAN_IN), .B2(keyinput174), .C1(
        P3_REG3_REG_9__SCAN_IN), .C2(keyinput187), .A(n15179), .ZN(n15184) );
  AOI22_X1 U16750 ( .A1(P1_REG1_REG_19__SCAN_IN), .A2(keyinput148), .B1(
        P3_REG0_REG_8__SCAN_IN), .B2(keyinput203), .ZN(n15180) );
  OAI221_X1 U16751 ( .B1(P1_REG1_REG_19__SCAN_IN), .B2(keyinput148), .C1(
        P3_REG0_REG_8__SCAN_IN), .C2(keyinput203), .A(n15180), .ZN(n15183) );
  AOI22_X1 U16752 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput205), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput157), .ZN(n15181) );
  OAI221_X1 U16753 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput205), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput157), .A(n15181), .ZN(n15182) );
  NOR4_X1 U16754 ( .A1(n15185), .A2(n15184), .A3(n15183), .A4(n15182), .ZN(
        n15204) );
  AOI22_X1 U16755 ( .A1(P2_REG1_REG_25__SCAN_IN), .A2(keyinput247), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(keyinput227), .ZN(n15186) );
  OAI221_X1 U16756 ( .B1(P2_REG1_REG_25__SCAN_IN), .B2(keyinput247), .C1(
        P1_DATAO_REG_28__SCAN_IN), .C2(keyinput227), .A(n15186), .ZN(n15193)
         );
  AOI22_X1 U16757 ( .A1(P1_D_REG_8__SCAN_IN), .A2(keyinput234), .B1(
        P3_REG0_REG_4__SCAN_IN), .B2(keyinput162), .ZN(n15187) );
  OAI221_X1 U16758 ( .B1(P1_D_REG_8__SCAN_IN), .B2(keyinput234), .C1(
        P3_REG0_REG_4__SCAN_IN), .C2(keyinput162), .A(n15187), .ZN(n15192) );
  AOI22_X1 U16759 ( .A1(P3_DATAO_REG_25__SCAN_IN), .A2(keyinput168), .B1(
        P1_REG2_REG_14__SCAN_IN), .B2(keyinput128), .ZN(n15188) );
  OAI221_X1 U16760 ( .B1(P3_DATAO_REG_25__SCAN_IN), .B2(keyinput168), .C1(
        P1_REG2_REG_14__SCAN_IN), .C2(keyinput128), .A(n15188), .ZN(n15191) );
  AOI22_X1 U16761 ( .A1(P1_REG0_REG_20__SCAN_IN), .A2(keyinput167), .B1(
        P1_IR_REG_29__SCAN_IN), .B2(keyinput163), .ZN(n15189) );
  OAI221_X1 U16762 ( .B1(P1_REG0_REG_20__SCAN_IN), .B2(keyinput167), .C1(
        P1_IR_REG_29__SCAN_IN), .C2(keyinput163), .A(n15189), .ZN(n15190) );
  NOR4_X1 U16763 ( .A1(n15193), .A2(n15192), .A3(n15191), .A4(n15190), .ZN(
        n15203) );
  AOI22_X1 U16764 ( .A1(P1_REG2_REG_24__SCAN_IN), .A2(keyinput194), .B1(
        P3_D_REG_1__SCAN_IN), .B2(keyinput236), .ZN(n15194) );
  OAI221_X1 U16765 ( .B1(P1_REG2_REG_24__SCAN_IN), .B2(keyinput194), .C1(
        P3_D_REG_1__SCAN_IN), .C2(keyinput236), .A(n15194), .ZN(n15201) );
  AOI22_X1 U16766 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(keyinput220), .B1(
        P3_REG3_REG_16__SCAN_IN), .B2(keyinput222), .ZN(n15195) );
  OAI221_X1 U16767 ( .B1(P2_IR_REG_8__SCAN_IN), .B2(keyinput220), .C1(
        P3_REG3_REG_16__SCAN_IN), .C2(keyinput222), .A(n15195), .ZN(n15200) );
  AOI22_X1 U16768 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput208), .B1(
        P3_REG1_REG_27__SCAN_IN), .B2(keyinput219), .ZN(n15196) );
  OAI221_X1 U16769 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput208), .C1(
        P3_REG1_REG_27__SCAN_IN), .C2(keyinput219), .A(n15196), .ZN(n15199) );
  AOI22_X1 U16770 ( .A1(P1_REG1_REG_23__SCAN_IN), .A2(keyinput140), .B1(
        P1_D_REG_7__SCAN_IN), .B2(keyinput239), .ZN(n15197) );
  OAI221_X1 U16771 ( .B1(P1_REG1_REG_23__SCAN_IN), .B2(keyinput140), .C1(
        P1_D_REG_7__SCAN_IN), .C2(keyinput239), .A(n15197), .ZN(n15198) );
  NOR4_X1 U16772 ( .A1(n15201), .A2(n15200), .A3(n15199), .A4(n15198), .ZN(
        n15202) );
  NAND4_X1 U16773 ( .A1(n15205), .A2(n15204), .A3(n15203), .A4(n15202), .ZN(
        n15313) );
  INV_X1 U16774 ( .A(P1_WR_REG_SCAN_IN), .ZN(n15404) );
  AOI22_X1 U16775 ( .A1(keyinput230), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n15404), .B2(keyinput212), .ZN(n15206) );
  OAI221_X1 U16776 ( .B1(keyinput230), .B2(P1_REG2_REG_26__SCAN_IN), .C1(
        n15404), .C2(keyinput212), .A(n15206), .ZN(n15215) );
  AOI22_X1 U16777 ( .A1(n15330), .A2(keyinput253), .B1(keyinput188), .B2(
        n15333), .ZN(n15207) );
  OAI221_X1 U16778 ( .B1(n15330), .B2(keyinput253), .C1(n15333), .C2(
        keyinput188), .A(n15207), .ZN(n15214) );
  AOI22_X1 U16779 ( .A1(n15209), .A2(keyinput151), .B1(keyinput135), .B2(
        n14893), .ZN(n15208) );
  OAI221_X1 U16780 ( .B1(n15209), .B2(keyinput151), .C1(n14893), .C2(
        keyinput135), .A(n15208), .ZN(n15213) );
  AOI22_X1 U16781 ( .A1(n15211), .A2(keyinput214), .B1(keyinput138), .B2(
        n10818), .ZN(n15210) );
  OAI221_X1 U16782 ( .B1(n15211), .B2(keyinput214), .C1(n10818), .C2(
        keyinput138), .A(n15210), .ZN(n15212) );
  NOR4_X1 U16783 ( .A1(n15215), .A2(n15214), .A3(n15213), .A4(n15212), .ZN(
        n15259) );
  AOI22_X1 U16784 ( .A1(n15218), .A2(keyinput145), .B1(keyinput182), .B2(
        n15217), .ZN(n15216) );
  OAI221_X1 U16785 ( .B1(n15218), .B2(keyinput145), .C1(n15217), .C2(
        keyinput182), .A(n15216), .ZN(n15223) );
  XNOR2_X1 U16786 ( .A(n15219), .B(keyinput229), .ZN(n15222) );
  XNOR2_X1 U16787 ( .A(n15220), .B(keyinput147), .ZN(n15221) );
  OR3_X1 U16788 ( .A1(n15223), .A2(n15222), .A3(n15221), .ZN(n15230) );
  AOI22_X1 U16789 ( .A1(n15397), .A2(keyinput250), .B1(keyinput238), .B2(
        n15225), .ZN(n15224) );
  OAI221_X1 U16790 ( .B1(n15397), .B2(keyinput250), .C1(n15225), .C2(
        keyinput238), .A(n15224), .ZN(n15229) );
  AOI22_X1 U16791 ( .A1(n15227), .A2(keyinput153), .B1(keyinput193), .B2(
        n15420), .ZN(n15226) );
  OAI221_X1 U16792 ( .B1(n15227), .B2(keyinput153), .C1(n15420), .C2(
        keyinput193), .A(n15226), .ZN(n15228) );
  NOR3_X1 U16793 ( .A1(n15230), .A2(n15229), .A3(n15228), .ZN(n15258) );
  INV_X1 U16794 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n15233) );
  AOI22_X1 U16795 ( .A1(n15233), .A2(keyinput134), .B1(keyinput198), .B2(
        n15232), .ZN(n15231) );
  OAI221_X1 U16796 ( .B1(n15233), .B2(keyinput134), .C1(n15232), .C2(
        keyinput198), .A(n15231), .ZN(n15244) );
  INV_X1 U16797 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n15353) );
  AOI22_X1 U16798 ( .A1(n15353), .A2(keyinput141), .B1(n15235), .B2(
        keyinput130), .ZN(n15234) );
  OAI221_X1 U16799 ( .B1(n15353), .B2(keyinput141), .C1(n15235), .C2(
        keyinput130), .A(n15234), .ZN(n15243) );
  AOI22_X1 U16800 ( .A1(n13172), .A2(keyinput254), .B1(keyinput181), .B2(
        n15237), .ZN(n15236) );
  OAI221_X1 U16801 ( .B1(n13172), .B2(keyinput254), .C1(n15237), .C2(
        keyinput181), .A(n15236), .ZN(n15242) );
  AOI22_X1 U16802 ( .A1(n15240), .A2(keyinput177), .B1(n15239), .B2(
        keyinput196), .ZN(n15238) );
  OAI221_X1 U16803 ( .B1(n15240), .B2(keyinput177), .C1(n15239), .C2(
        keyinput196), .A(n15238), .ZN(n15241) );
  NOR4_X1 U16804 ( .A1(n15244), .A2(n15243), .A3(n15242), .A4(n15241), .ZN(
        n15257) );
  AOI22_X1 U16805 ( .A1(n15424), .A2(keyinput249), .B1(n15246), .B2(
        keyinput201), .ZN(n15245) );
  OAI221_X1 U16806 ( .B1(n15424), .B2(keyinput249), .C1(n15246), .C2(
        keyinput201), .A(n15245), .ZN(n15255) );
  AOI22_X1 U16807 ( .A1(n15248), .A2(keyinput197), .B1(n15324), .B2(
        keyinput235), .ZN(n15247) );
  OAI221_X1 U16808 ( .B1(n15248), .B2(keyinput197), .C1(n15324), .C2(
        keyinput235), .A(n15247), .ZN(n15254) );
  INV_X1 U16809 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n15365) );
  XOR2_X1 U16810 ( .A(n15365), .B(keyinput132), .Z(n15251) );
  XNOR2_X1 U16811 ( .A(P3_IR_REG_12__SCAN_IN), .B(keyinput186), .ZN(n15250) );
  XNOR2_X1 U16812 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput211), .ZN(n15249)
         );
  NAND3_X1 U16813 ( .A1(n15251), .A2(n15250), .A3(n15249), .ZN(n15253) );
  XNOR2_X1 U16814 ( .A(n15340), .B(keyinput246), .ZN(n15252) );
  NOR4_X1 U16815 ( .A1(n15255), .A2(n15254), .A3(n15253), .A4(n15252), .ZN(
        n15256) );
  NAND4_X1 U16816 ( .A1(n15259), .A2(n15258), .A3(n15257), .A4(n15256), .ZN(
        n15312) );
  AOI22_X1 U16817 ( .A1(n15399), .A2(keyinput172), .B1(n8654), .B2(keyinput192), .ZN(n15260) );
  OAI221_X1 U16818 ( .B1(n15399), .B2(keyinput172), .C1(n8654), .C2(
        keyinput192), .A(n15260), .ZN(n15263) );
  XOR2_X1 U16819 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput156), .Z(n15262) );
  XNOR2_X1 U16820 ( .A(n15405), .B(keyinput161), .ZN(n15261) );
  OR3_X1 U16821 ( .A1(n15263), .A2(n15262), .A3(n15261), .ZN(n15271) );
  AOI22_X1 U16822 ( .A1(n15265), .A2(keyinput183), .B1(n7788), .B2(keyinput143), .ZN(n15264) );
  OAI221_X1 U16823 ( .B1(n15265), .B2(keyinput183), .C1(n7788), .C2(
        keyinput143), .A(n15264), .ZN(n15270) );
  AOI22_X1 U16824 ( .A1(n15268), .A2(keyinput184), .B1(keyinput215), .B2(
        n15267), .ZN(n15266) );
  OAI221_X1 U16825 ( .B1(n15268), .B2(keyinput184), .C1(n15267), .C2(
        keyinput215), .A(n15266), .ZN(n15269) );
  NOR3_X1 U16826 ( .A1(n15271), .A2(n15270), .A3(n15269), .ZN(n15310) );
  AOI22_X1 U16827 ( .A1(n12928), .A2(keyinput159), .B1(keyinput200), .B2(
        n15423), .ZN(n15272) );
  OAI221_X1 U16828 ( .B1(n12928), .B2(keyinput159), .C1(n15423), .C2(
        keyinput200), .A(n15272), .ZN(n15281) );
  AOI22_X1 U16829 ( .A1(n15341), .A2(keyinput175), .B1(keyinput217), .B2(
        n15274), .ZN(n15273) );
  OAI221_X1 U16830 ( .B1(n15341), .B2(keyinput175), .C1(n15274), .C2(
        keyinput217), .A(n15273), .ZN(n15280) );
  XNOR2_X1 U16831 ( .A(P3_REG3_REG_18__SCAN_IN), .B(keyinput160), .ZN(n15278)
         );
  XNOR2_X1 U16832 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput210), .ZN(n15277)
         );
  XNOR2_X1 U16833 ( .A(P1_REG3_REG_1__SCAN_IN), .B(keyinput195), .ZN(n15276)
         );
  XNOR2_X1 U16834 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(keyinput131), .ZN(n15275)
         );
  NAND4_X1 U16835 ( .A1(n15278), .A2(n15277), .A3(n15276), .A4(n15275), .ZN(
        n15279) );
  NOR3_X1 U16836 ( .A1(n15281), .A2(n15280), .A3(n15279), .ZN(n15309) );
  INV_X1 U16837 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n15361) );
  AOI22_X1 U16838 ( .A1(n15361), .A2(keyinput213), .B1(keyinput204), .B2(
        n15283), .ZN(n15282) );
  OAI221_X1 U16839 ( .B1(n15361), .B2(keyinput213), .C1(n15283), .C2(
        keyinput204), .A(n15282), .ZN(n15294) );
  AOI22_X1 U16840 ( .A1(n15286), .A2(keyinput225), .B1(n15285), .B2(
        keyinput166), .ZN(n15284) );
  OAI221_X1 U16841 ( .B1(n15286), .B2(keyinput225), .C1(n15285), .C2(
        keyinput166), .A(n15284), .ZN(n15293) );
  AOI22_X1 U16842 ( .A1(n15411), .A2(keyinput243), .B1(n15288), .B2(
        keyinput139), .ZN(n15287) );
  OAI221_X1 U16843 ( .B1(n15411), .B2(keyinput243), .C1(n15288), .C2(
        keyinput139), .A(n15287), .ZN(n15292) );
  XNOR2_X1 U16844 ( .A(P3_IR_REG_6__SCAN_IN), .B(keyinput226), .ZN(n15290) );
  XNOR2_X1 U16845 ( .A(P2_REG0_REG_21__SCAN_IN), .B(keyinput248), .ZN(n15289)
         );
  NAND2_X1 U16846 ( .A1(n15290), .A2(n15289), .ZN(n15291) );
  NOR4_X1 U16847 ( .A1(n15294), .A2(n15293), .A3(n15292), .A4(n15291), .ZN(
        n15308) );
  AOI22_X1 U16848 ( .A1(n15296), .A2(keyinput170), .B1(keyinput199), .B2(
        n10248), .ZN(n15295) );
  OAI221_X1 U16849 ( .B1(n15296), .B2(keyinput170), .C1(n10248), .C2(
        keyinput199), .A(n15295), .ZN(n15306) );
  INV_X1 U16850 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n15298) );
  AOI22_X1 U16851 ( .A1(n15364), .A2(keyinput231), .B1(keyinput209), .B2(
        n15298), .ZN(n15297) );
  OAI221_X1 U16852 ( .B1(n15364), .B2(keyinput231), .C1(n15298), .C2(
        keyinput209), .A(n15297), .ZN(n15305) );
  AOI22_X1 U16853 ( .A1(n15417), .A2(keyinput178), .B1(keyinput233), .B2(
        n15300), .ZN(n15299) );
  OAI221_X1 U16854 ( .B1(n15417), .B2(keyinput178), .C1(n15300), .C2(
        keyinput233), .A(n15299), .ZN(n15304) );
  INV_X1 U16855 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n15302) );
  AOI22_X1 U16856 ( .A1(n15302), .A2(keyinput240), .B1(n15344), .B2(
        keyinput154), .ZN(n15301) );
  OAI221_X1 U16857 ( .B1(n15302), .B2(keyinput240), .C1(n15344), .C2(
        keyinput154), .A(n15301), .ZN(n15303) );
  NOR4_X1 U16858 ( .A1(n15306), .A2(n15305), .A3(n15304), .A4(n15303), .ZN(
        n15307) );
  NAND4_X1 U16859 ( .A1(n15310), .A2(n15309), .A3(n15308), .A4(n15307), .ZN(
        n15311) );
  NOR4_X1 U16860 ( .A1(n15314), .A2(n15313), .A3(n15312), .A4(n15311), .ZN(
        n15512) );
  AOI22_X1 U16861 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput48), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput29), .ZN(n15315) );
  OAI221_X1 U16862 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput48), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput29), .A(n15315), .ZN(n15322) );
  AOI22_X1 U16863 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(keyinput99), .B1(
        P3_D_REG_2__SCAN_IN), .B2(keyinput51), .ZN(n15316) );
  OAI221_X1 U16864 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(keyinput99), .C1(
        P3_D_REG_2__SCAN_IN), .C2(keyinput51), .A(n15316), .ZN(n15321) );
  AOI22_X1 U16865 ( .A1(P3_DATAO_REG_8__SCAN_IN), .A2(keyinput19), .B1(
        P2_REG2_REG_1__SCAN_IN), .B2(keyinput16), .ZN(n15317) );
  OAI221_X1 U16866 ( .B1(P3_DATAO_REG_8__SCAN_IN), .B2(keyinput19), .C1(
        P2_REG2_REG_1__SCAN_IN), .C2(keyinput16), .A(n15317), .ZN(n15320) );
  AOI22_X1 U16867 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(keyinput92), .B1(
        P3_REG3_REG_9__SCAN_IN), .B2(keyinput59), .ZN(n15318) );
  OAI221_X1 U16868 ( .B1(P2_IR_REG_8__SCAN_IN), .B2(keyinput92), .C1(
        P3_REG3_REG_9__SCAN_IN), .C2(keyinput59), .A(n15318), .ZN(n15319) );
  NOR4_X1 U16869 ( .A1(n15322), .A2(n15321), .A3(n15320), .A4(n15319), .ZN(
        n15372) );
  INV_X1 U16870 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n15325) );
  AOI22_X1 U16871 ( .A1(n15325), .A2(keyinput66), .B1(n15324), .B2(keyinput107), .ZN(n15323) );
  OAI221_X1 U16872 ( .B1(n15325), .B2(keyinput66), .C1(n15324), .C2(
        keyinput107), .A(n15323), .ZN(n15338) );
  AOI22_X1 U16873 ( .A1(n15328), .A2(keyinput62), .B1(n15327), .B2(keyinput22), 
        .ZN(n15326) );
  OAI221_X1 U16874 ( .B1(n15328), .B2(keyinput62), .C1(n15327), .C2(keyinput22), .A(n15326), .ZN(n15337) );
  INV_X1 U16875 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n15331) );
  AOI22_X1 U16876 ( .A1(n15331), .A2(keyinput108), .B1(keyinput125), .B2(
        n15330), .ZN(n15329) );
  OAI221_X1 U16877 ( .B1(n15331), .B2(keyinput108), .C1(n15330), .C2(
        keyinput125), .A(n15329), .ZN(n15336) );
  AOI22_X1 U16878 ( .A1(n15334), .A2(keyinput37), .B1(keyinput60), .B2(n15333), 
        .ZN(n15332) );
  OAI221_X1 U16879 ( .B1(n15334), .B2(keyinput37), .C1(n15333), .C2(keyinput60), .A(n15332), .ZN(n15335) );
  NOR4_X1 U16880 ( .A1(n15338), .A2(n15337), .A3(n15336), .A4(n15335), .ZN(
        n15371) );
  AOI22_X1 U16881 ( .A1(n15341), .A2(keyinput47), .B1(keyinput118), .B2(n15340), .ZN(n15339) );
  OAI221_X1 U16882 ( .B1(n15341), .B2(keyinput47), .C1(n15340), .C2(
        keyinput118), .A(n15339), .ZN(n15351) );
  AOI22_X1 U16883 ( .A1(n15344), .A2(keyinput26), .B1(n15343), .B2(keyinput79), 
        .ZN(n15342) );
  OAI221_X1 U16884 ( .B1(n15344), .B2(keyinput26), .C1(n15343), .C2(keyinput79), .A(n15342), .ZN(n15350) );
  XNOR2_X1 U16885 ( .A(P1_REG1_REG_23__SCAN_IN), .B(keyinput12), .ZN(n15348)
         );
  XNOR2_X1 U16886 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput83), .ZN(n15347) );
  XNOR2_X1 U16887 ( .A(P2_IR_REG_15__SCAN_IN), .B(keyinput101), .ZN(n15346) );
  XNOR2_X1 U16888 ( .A(P1_REG1_REG_19__SCAN_IN), .B(keyinput20), .ZN(n15345)
         );
  NAND4_X1 U16889 ( .A1(n15348), .A2(n15347), .A3(n15346), .A4(n15345), .ZN(
        n15349) );
  NOR3_X1 U16890 ( .A1(n15351), .A2(n15350), .A3(n15349), .ZN(n15370) );
  INV_X1 U16891 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n15354) );
  AOI22_X1 U16892 ( .A1(n15354), .A2(keyinput102), .B1(keyinput13), .B2(n15353), .ZN(n15352) );
  OAI221_X1 U16893 ( .B1(n15354), .B2(keyinput102), .C1(n15353), .C2(
        keyinput13), .A(n15352), .ZN(n15359) );
  XNOR2_X1 U16894 ( .A(n15355), .B(keyinput96), .ZN(n15358) );
  XNOR2_X1 U16895 ( .A(n15356), .B(keyinput5), .ZN(n15357) );
  OR3_X1 U16896 ( .A1(n15359), .A2(n15358), .A3(n15357), .ZN(n15368) );
  AOI22_X1 U16897 ( .A1(n15362), .A2(keyinput36), .B1(n15361), .B2(keyinput85), 
        .ZN(n15360) );
  OAI221_X1 U16898 ( .B1(n15362), .B2(keyinput36), .C1(n15361), .C2(keyinput85), .A(n15360), .ZN(n15367) );
  AOI22_X1 U16899 ( .A1(n15365), .A2(keyinput4), .B1(n15364), .B2(keyinput103), 
        .ZN(n15363) );
  OAI221_X1 U16900 ( .B1(n15365), .B2(keyinput4), .C1(n15364), .C2(keyinput103), .A(n15363), .ZN(n15366) );
  NOR3_X1 U16901 ( .A1(n15368), .A2(n15367), .A3(n15366), .ZN(n15369) );
  NAND4_X1 U16902 ( .A1(n15372), .A2(n15371), .A3(n15370), .A4(n15369), .ZN(
        n15511) );
  AOI22_X1 U16903 ( .A1(n15375), .A2(keyinput21), .B1(keyinput117), .B2(n15374), .ZN(n15373) );
  OAI221_X1 U16904 ( .B1(n15375), .B2(keyinput21), .C1(n15374), .C2(
        keyinput117), .A(n15373), .ZN(n15387) );
  AOI22_X1 U16905 ( .A1(n15378), .A2(keyinput32), .B1(keyinput1), .B2(n15377), 
        .ZN(n15376) );
  OAI221_X1 U16906 ( .B1(n15378), .B2(keyinput32), .C1(n15377), .C2(keyinput1), 
        .A(n15376), .ZN(n15386) );
  INV_X1 U16907 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n15380) );
  AOI22_X1 U16908 ( .A1(n15380), .A2(keyinput119), .B1(n8654), .B2(keyinput64), 
        .ZN(n15379) );
  OAI221_X1 U16909 ( .B1(n15380), .B2(keyinput119), .C1(n8654), .C2(keyinput64), .A(n15379), .ZN(n15385) );
  XOR2_X1 U16910 ( .A(n15381), .B(keyinput34), .Z(n15383) );
  XNOR2_X1 U16911 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput77), .ZN(n15382) );
  NAND2_X1 U16912 ( .A1(n15383), .A2(n15382), .ZN(n15384) );
  NOR4_X1 U16913 ( .A1(n15387), .A2(n15386), .A3(n15385), .A4(n15384), .ZN(
        n15434) );
  AOI22_X1 U16914 ( .A1(n11716), .A2(keyinput24), .B1(keyinput74), .B2(n14677), 
        .ZN(n15388) );
  OAI221_X1 U16915 ( .B1(n11716), .B2(keyinput24), .C1(n14677), .C2(keyinput74), .A(n15388), .ZN(n15395) );
  INV_X1 U16916 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n15391) );
  AOI22_X1 U16917 ( .A1(n15391), .A2(keyinput27), .B1(keyinput39), .B2(n15390), 
        .ZN(n15389) );
  OAI221_X1 U16918 ( .B1(n15391), .B2(keyinput27), .C1(n15390), .C2(keyinput39), .A(n15389), .ZN(n15394) );
  XNOR2_X1 U16919 ( .A(n15392), .B(keyinput98), .ZN(n15393) );
  OR3_X1 U16920 ( .A1(n15395), .A2(n15394), .A3(n15393), .ZN(n15402) );
  AOI22_X1 U16921 ( .A1(n15398), .A2(keyinput100), .B1(keyinput122), .B2(
        n15397), .ZN(n15396) );
  OAI221_X1 U16922 ( .B1(n15398), .B2(keyinput100), .C1(n15397), .C2(
        keyinput122), .A(n15396), .ZN(n15401) );
  XNOR2_X1 U16923 ( .A(n15399), .B(keyinput44), .ZN(n15400) );
  NOR3_X1 U16924 ( .A1(n15402), .A2(n15401), .A3(n15400), .ZN(n15433) );
  AOI22_X1 U16925 ( .A1(n15405), .A2(keyinput33), .B1(keyinput84), .B2(n15404), 
        .ZN(n15403) );
  OAI221_X1 U16926 ( .B1(n15405), .B2(keyinput33), .C1(n15404), .C2(keyinput84), .A(n15403), .ZN(n15415) );
  AOI22_X1 U16927 ( .A1(n7788), .A2(keyinput15), .B1(keyinput111), .B2(n15407), 
        .ZN(n15406) );
  OAI221_X1 U16928 ( .B1(n7788), .B2(keyinput15), .C1(n15407), .C2(keyinput111), .A(n15406), .ZN(n15414) );
  XNOR2_X1 U16929 ( .A(P3_IR_REG_12__SCAN_IN), .B(keyinput58), .ZN(n15410) );
  XNOR2_X1 U16930 ( .A(P2_REG1_REG_22__SCAN_IN), .B(keyinput17), .ZN(n15409)
         );
  XNOR2_X1 U16931 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput14), .ZN(n15408)
         );
  NAND3_X1 U16932 ( .A1(n15410), .A2(n15409), .A3(n15408), .ZN(n15413) );
  XNOR2_X1 U16933 ( .A(n15411), .B(keyinput115), .ZN(n15412) );
  NOR4_X1 U16934 ( .A1(n15415), .A2(n15414), .A3(n15413), .A4(n15412), .ZN(
        n15432) );
  AOI22_X1 U16935 ( .A1(n15418), .A2(keyinput124), .B1(n15417), .B2(keyinput50), .ZN(n15416) );
  OAI221_X1 U16936 ( .B1(n15418), .B2(keyinput124), .C1(n15417), .C2(
        keyinput50), .A(n15416), .ZN(n15430) );
  AOI22_X1 U16937 ( .A1(n15421), .A2(keyinput116), .B1(keyinput65), .B2(n15420), .ZN(n15419) );
  OAI221_X1 U16938 ( .B1(n15421), .B2(keyinput116), .C1(n15420), .C2(
        keyinput65), .A(n15419), .ZN(n15429) );
  AOI22_X1 U16939 ( .A1(n15424), .A2(keyinput121), .B1(n15423), .B2(keyinput72), .ZN(n15422) );
  OAI221_X1 U16940 ( .B1(n15424), .B2(keyinput121), .C1(n15423), .C2(
        keyinput72), .A(n15422), .ZN(n15428) );
  XNOR2_X1 U16941 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput82), .ZN(n15426)
         );
  XNOR2_X1 U16942 ( .A(P1_REG0_REG_19__SCAN_IN), .B(keyinput95), .ZN(n15425)
         );
  NAND2_X1 U16943 ( .A1(n15426), .A2(n15425), .ZN(n15427) );
  NOR4_X1 U16944 ( .A1(n15430), .A2(n15429), .A3(n15428), .A4(n15427), .ZN(
        n15431) );
  NAND4_X1 U16945 ( .A1(n15434), .A2(n15433), .A3(n15432), .A4(n15431), .ZN(
        n15510) );
  OAI22_X1 U16946 ( .A1(P3_REG3_REG_16__SCAN_IN), .A2(keyinput94), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(keyinput8), .ZN(n15435) );
  AOI221_X1 U16947 ( .B1(P3_REG3_REG_16__SCAN_IN), .B2(keyinput94), .C1(
        keyinput8), .C2(P2_DATAO_REG_25__SCAN_IN), .A(n15435), .ZN(n15442) );
  OAI22_X1 U16948 ( .A1(P3_REG1_REG_27__SCAN_IN), .A2(keyinput91), .B1(
        keyinput123), .B2(P1_D_REG_6__SCAN_IN), .ZN(n15436) );
  AOI221_X1 U16949 ( .B1(P3_REG1_REG_27__SCAN_IN), .B2(keyinput91), .C1(
        P1_D_REG_6__SCAN_IN), .C2(keyinput123), .A(n15436), .ZN(n15441) );
  OAI22_X1 U16950 ( .A1(P3_D_REG_31__SCAN_IN), .A2(keyinput56), .B1(
        keyinput105), .B2(P1_D_REG_23__SCAN_IN), .ZN(n15437) );
  AOI221_X1 U16951 ( .B1(P3_D_REG_31__SCAN_IN), .B2(keyinput56), .C1(
        P1_D_REG_23__SCAN_IN), .C2(keyinput105), .A(n15437), .ZN(n15440) );
  OAI22_X1 U16952 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(keyinput43), .B1(
        keyinput87), .B2(P3_ADDR_REG_1__SCAN_IN), .ZN(n15438) );
  AOI221_X1 U16953 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(keyinput43), .C1(
        P3_ADDR_REG_1__SCAN_IN), .C2(keyinput87), .A(n15438), .ZN(n15439) );
  NAND4_X1 U16954 ( .A1(n15442), .A2(n15441), .A3(n15440), .A4(n15439), .ZN(
        n15470) );
  OAI22_X1 U16955 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(keyinput127), .B1(
        P2_D_REG_2__SCAN_IN), .B2(keyinput78), .ZN(n15443) );
  AOI221_X1 U16956 ( .B1(P3_REG3_REG_5__SCAN_IN), .B2(keyinput127), .C1(
        keyinput78), .C2(P2_D_REG_2__SCAN_IN), .A(n15443), .ZN(n15450) );
  OAI22_X1 U16957 ( .A1(P1_D_REG_24__SCAN_IN), .A2(keyinput97), .B1(
        P1_REG2_REG_14__SCAN_IN), .B2(keyinput0), .ZN(n15444) );
  AOI221_X1 U16958 ( .B1(P1_D_REG_24__SCAN_IN), .B2(keyinput97), .C1(keyinput0), .C2(P1_REG2_REG_14__SCAN_IN), .A(n15444), .ZN(n15449) );
  OAI22_X1 U16959 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(keyinput114), .B1(
        P2_REG1_REG_13__SCAN_IN), .B2(keyinput112), .ZN(n15445) );
  AOI221_X1 U16960 ( .B1(P2_DATAO_REG_1__SCAN_IN), .B2(keyinput114), .C1(
        keyinput112), .C2(P2_REG1_REG_13__SCAN_IN), .A(n15445), .ZN(n15448) );
  OAI22_X1 U16961 ( .A1(P3_REG1_REG_30__SCAN_IN), .A2(keyinput9), .B1(
        keyinput90), .B2(P1_ADDR_REG_17__SCAN_IN), .ZN(n15446) );
  AOI221_X1 U16962 ( .B1(P3_REG1_REG_30__SCAN_IN), .B2(keyinput9), .C1(
        P1_ADDR_REG_17__SCAN_IN), .C2(keyinput90), .A(n15446), .ZN(n15447) );
  NAND4_X1 U16963 ( .A1(n15450), .A2(n15449), .A3(n15448), .A4(n15447), .ZN(
        n15469) );
  OAI22_X1 U16964 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(keyinput104), .B1(
        keyinput93), .B2(P2_IR_REG_5__SCAN_IN), .ZN(n15451) );
  AOI221_X1 U16965 ( .B1(P3_REG1_REG_18__SCAN_IN), .B2(keyinput104), .C1(
        P2_IR_REG_5__SCAN_IN), .C2(keyinput93), .A(n15451), .ZN(n15458) );
  OAI22_X1 U16966 ( .A1(P2_REG2_REG_28__SCAN_IN), .A2(keyinput126), .B1(
        P1_D_REG_25__SCAN_IN), .B2(keyinput49), .ZN(n15452) );
  AOI221_X1 U16967 ( .B1(P2_REG2_REG_28__SCAN_IN), .B2(keyinput126), .C1(
        keyinput49), .C2(P1_D_REG_25__SCAN_IN), .A(n15452), .ZN(n15457) );
  OAI22_X1 U16968 ( .A1(P3_REG0_REG_11__SCAN_IN), .A2(keyinput23), .B1(
        keyinput57), .B2(P1_REG0_REG_30__SCAN_IN), .ZN(n15453) );
  AOI221_X1 U16969 ( .B1(P3_REG0_REG_11__SCAN_IN), .B2(keyinput23), .C1(
        P1_REG0_REG_30__SCAN_IN), .C2(keyinput57), .A(n15453), .ZN(n15456) );
  OAI22_X1 U16970 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(keyinput35), .B1(
        keyinput53), .B2(P2_ADDR_REG_14__SCAN_IN), .ZN(n15454) );
  AOI221_X1 U16971 ( .B1(P1_IR_REG_29__SCAN_IN), .B2(keyinput35), .C1(
        P2_ADDR_REG_14__SCAN_IN), .C2(keyinput53), .A(n15454), .ZN(n15455) );
  NAND4_X1 U16972 ( .A1(n15458), .A2(n15457), .A3(n15456), .A4(n15455), .ZN(
        n15468) );
  OAI22_X1 U16973 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(keyinput86), .B1(
        P3_DATAO_REG_14__SCAN_IN), .B2(keyinput76), .ZN(n15459) );
  AOI221_X1 U16974 ( .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput86), .C1(
        keyinput76), .C2(P3_DATAO_REG_14__SCAN_IN), .A(n15459), .ZN(n15466) );
  OAI22_X1 U16975 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(keyinput63), .B1(
        P1_D_REG_8__SCAN_IN), .B2(keyinput106), .ZN(n15460) );
  AOI221_X1 U16976 ( .B1(P2_DATAO_REG_14__SCAN_IN), .B2(keyinput63), .C1(
        keyinput106), .C2(P1_D_REG_8__SCAN_IN), .A(n15460), .ZN(n15465) );
  OAI22_X1 U16977 ( .A1(P3_REG0_REG_8__SCAN_IN), .A2(keyinput75), .B1(
        P3_DATAO_REG_9__SCAN_IN), .B2(keyinput54), .ZN(n15461) );
  AOI221_X1 U16978 ( .B1(P3_REG0_REG_8__SCAN_IN), .B2(keyinput75), .C1(
        keyinput54), .C2(P3_DATAO_REG_9__SCAN_IN), .A(n15461), .ZN(n15464) );
  OAI22_X1 U16979 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(keyinput28), .B1(
        keyinput110), .B2(P2_ADDR_REG_4__SCAN_IN), .ZN(n15462) );
  AOI221_X1 U16980 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(keyinput28), .C1(
        P2_ADDR_REG_4__SCAN_IN), .C2(keyinput110), .A(n15462), .ZN(n15463) );
  NAND4_X1 U16981 ( .A1(n15466), .A2(n15465), .A3(n15464), .A4(n15463), .ZN(
        n15467) );
  NOR4_X1 U16982 ( .A1(n15470), .A2(n15469), .A3(n15468), .A4(n15467), .ZN(
        n15508) );
  OAI22_X1 U16983 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput68), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(keyinput30), .ZN(n15471) );
  AOI221_X1 U16984 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput68), .C1(
        keyinput30), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n15471), .ZN(n15478) );
  OAI22_X1 U16985 ( .A1(SI_15_), .A2(keyinput25), .B1(P1_REG1_REG_13__SCAN_IN), 
        .B2(keyinput10), .ZN(n15472) );
  AOI221_X1 U16986 ( .B1(SI_15_), .B2(keyinput25), .C1(keyinput10), .C2(
        P1_REG1_REG_13__SCAN_IN), .A(n15472), .ZN(n15477) );
  OAI22_X1 U16987 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(keyinput2), .B1(
        P2_REG2_REG_2__SCAN_IN), .B2(keyinput113), .ZN(n15473) );
  AOI221_X1 U16988 ( .B1(P1_DATAO_REG_22__SCAN_IN), .B2(keyinput2), .C1(
        keyinput113), .C2(P2_REG2_REG_2__SCAN_IN), .A(n15473), .ZN(n15476) );
  OAI22_X1 U16989 ( .A1(SI_6_), .A2(keyinput11), .B1(keyinput67), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n15474) );
  AOI221_X1 U16990 ( .B1(SI_6_), .B2(keyinput11), .C1(P1_REG3_REG_1__SCAN_IN), 
        .C2(keyinput67), .A(n15474), .ZN(n15475) );
  NAND4_X1 U16991 ( .A1(n15478), .A2(n15477), .A3(n15476), .A4(n15475), .ZN(
        n15506) );
  OAI22_X1 U16992 ( .A1(P3_D_REG_10__SCAN_IN), .A2(keyinput55), .B1(
        P3_REG0_REG_23__SCAN_IN), .B2(keyinput6), .ZN(n15479) );
  AOI221_X1 U16993 ( .B1(P3_D_REG_10__SCAN_IN), .B2(keyinput55), .C1(keyinput6), .C2(P3_REG0_REG_23__SCAN_IN), .A(n15479), .ZN(n15486) );
  OAI22_X1 U16994 ( .A1(SI_2_), .A2(keyinput70), .B1(keyinput41), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n15480) );
  AOI221_X1 U16995 ( .B1(SI_2_), .B2(keyinput70), .C1(P2_REG1_REG_7__SCAN_IN), 
        .C2(keyinput41), .A(n15480), .ZN(n15485) );
  OAI22_X1 U16996 ( .A1(P3_IR_REG_30__SCAN_IN), .A2(keyinput31), .B1(
        keyinput42), .B2(P3_REG0_REG_2__SCAN_IN), .ZN(n15481) );
  AOI221_X1 U16997 ( .B1(P3_IR_REG_30__SCAN_IN), .B2(keyinput31), .C1(
        P3_REG0_REG_2__SCAN_IN), .C2(keyinput42), .A(n15481), .ZN(n15484) );
  OAI22_X1 U16998 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(keyinput109), .B1(
        P1_ADDR_REG_18__SCAN_IN), .B2(keyinput69), .ZN(n15482) );
  AOI221_X1 U16999 ( .B1(P1_IR_REG_21__SCAN_IN), .B2(keyinput109), .C1(
        keyinput69), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n15482), .ZN(n15483) );
  NAND4_X1 U17000 ( .A1(n15486), .A2(n15485), .A3(n15484), .A4(n15483), .ZN(
        n15505) );
  OAI22_X1 U17001 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(keyinput3), .B1(
        keyinput45), .B2(SI_17_), .ZN(n15487) );
  AOI221_X1 U17002 ( .B1(P1_DATAO_REG_25__SCAN_IN), .B2(keyinput3), .C1(SI_17_), .C2(keyinput45), .A(n15487), .ZN(n15494) );
  OAI22_X1 U17003 ( .A1(P2_D_REG_26__SCAN_IN), .A2(keyinput73), .B1(keyinput88), .B2(P2_REG1_REG_30__SCAN_IN), .ZN(n15488) );
  AOI221_X1 U17004 ( .B1(P2_D_REG_26__SCAN_IN), .B2(keyinput73), .C1(
        P2_REG1_REG_30__SCAN_IN), .C2(keyinput88), .A(n15488), .ZN(n15493) );
  OAI22_X1 U17005 ( .A1(P3_D_REG_7__SCAN_IN), .A2(keyinput61), .B1(
        P1_IR_REG_5__SCAN_IN), .B2(keyinput80), .ZN(n15489) );
  AOI221_X1 U17006 ( .B1(P3_D_REG_7__SCAN_IN), .B2(keyinput61), .C1(keyinput80), .C2(P1_IR_REG_5__SCAN_IN), .A(n15489), .ZN(n15492) );
  OAI22_X1 U17007 ( .A1(P2_REG1_REG_24__SCAN_IN), .A2(keyinput38), .B1(
        keyinput18), .B2(P1_D_REG_26__SCAN_IN), .ZN(n15490) );
  AOI221_X1 U17008 ( .B1(P2_REG1_REG_24__SCAN_IN), .B2(keyinput38), .C1(
        P1_D_REG_26__SCAN_IN), .C2(keyinput18), .A(n15490), .ZN(n15491) );
  NAND4_X1 U17009 ( .A1(n15494), .A2(n15493), .A3(n15492), .A4(n15491), .ZN(
        n15504) );
  OAI22_X1 U17010 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(keyinput7), .B1(
        P2_REG0_REG_25__SCAN_IN), .B2(keyinput89), .ZN(n15495) );
  AOI221_X1 U17011 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(keyinput7), .C1(
        keyinput89), .C2(P2_REG0_REG_25__SCAN_IN), .A(n15495), .ZN(n15502) );
  OAI22_X1 U17012 ( .A1(P2_REG2_REG_25__SCAN_IN), .A2(keyinput52), .B1(
        P3_DATAO_REG_25__SCAN_IN), .B2(keyinput40), .ZN(n15496) );
  AOI221_X1 U17013 ( .B1(P2_REG2_REG_25__SCAN_IN), .B2(keyinput52), .C1(
        keyinput40), .C2(P3_DATAO_REG_25__SCAN_IN), .A(n15496), .ZN(n15501) );
  OAI22_X1 U17014 ( .A1(P2_D_REG_8__SCAN_IN), .A2(keyinput46), .B1(
        P1_REG0_REG_17__SCAN_IN), .B2(keyinput81), .ZN(n15497) );
  AOI221_X1 U17015 ( .B1(P2_D_REG_8__SCAN_IN), .B2(keyinput46), .C1(keyinput81), .C2(P1_REG0_REG_17__SCAN_IN), .A(n15497), .ZN(n15500) );
  OAI22_X1 U17016 ( .A1(P2_REG0_REG_21__SCAN_IN), .A2(keyinput120), .B1(
        P2_REG2_REG_7__SCAN_IN), .B2(keyinput71), .ZN(n15498) );
  AOI221_X1 U17017 ( .B1(P2_REG0_REG_21__SCAN_IN), .B2(keyinput120), .C1(
        keyinput71), .C2(P2_REG2_REG_7__SCAN_IN), .A(n15498), .ZN(n15499) );
  NAND4_X1 U17018 ( .A1(n15502), .A2(n15501), .A3(n15500), .A4(n15499), .ZN(
        n15503) );
  NOR4_X1 U17019 ( .A1(n15506), .A2(n15505), .A3(n15504), .A4(n15503), .ZN(
        n15507) );
  NAND2_X1 U17020 ( .A1(n15508), .A2(n15507), .ZN(n15509) );
  NOR4_X1 U17021 ( .A1(n15512), .A2(n15511), .A3(n15510), .A4(n15509), .ZN(
        n15513) );
  XNOR2_X1 U17022 ( .A(n15514), .B(n15513), .ZN(P1_U3302) );
  XOR2_X1 U17023 ( .A(n15516), .B(n15515), .Z(SUB_1596_U59) );
  XNOR2_X1 U17024 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n15517), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U17025 ( .B1(n15519), .B2(n15518), .A(n15526), .ZN(SUB_1596_U53) );
  XOR2_X1 U17026 ( .A(n15521), .B(n15520), .Z(SUB_1596_U56) );
  NOR2_X1 U17027 ( .A1(n15523), .A2(n15522), .ZN(n15524) );
  XNOR2_X1 U17028 ( .A(n15524), .B(n14677), .ZN(SUB_1596_U60) );
  XOR2_X1 U17029 ( .A(n15526), .B(n15525), .Z(SUB_1596_U5) );
  CLKBUF_X1 U7368 ( .A(n9904), .Z(n10056) );
  CLKBUF_X3 U7385 ( .A(n7585), .Z(n10754) );
  INV_X2 U7399 ( .A(n10603), .ZN(n10612) );
  AOI21_X1 U7432 ( .B1(n13885), .B2(n13860), .A(n13874), .ZN(n13858) );
  CLKBUF_X1 U7454 ( .A(n10176), .Z(n6772) );
  CLKBUF_X1 U7457 ( .A(n13538), .Z(n6626) );
  CLKBUF_X1 U7462 ( .A(n7572), .Z(n7000) );
  CLKBUF_X1 U8949 ( .A(n8074), .Z(n6628) );
endmodule

