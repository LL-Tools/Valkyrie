

module b14_C_gen_AntiSAT_k_256_4 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091;

  OR2_X1 U2469 ( .A1(n3093), .A2(n3092), .ZN(n3655) );
  OR2_X1 U2470 ( .A1(n4217), .A2(n4145), .ZN(n4196) );
  NAND2_X1 U2471 ( .A1(n2276), .A2(n3562), .ZN(n3574) );
  CLKBUF_X2 U2472 ( .A(n2513), .Z(n2735) );
  OAI21_X1 U2473 ( .B1(n2227), .B2(n2346), .A(n2345), .ZN(n3256) );
  INV_X1 U2474 ( .A(n2955), .ZN(n2877) );
  AND2_X1 U2475 ( .A1(n2856), .A2(n2816), .ZN(n2488) );
  INV_X4 U2476 ( .A(n2242), .ZN(n2955) );
  OAI21_X1 U2477 ( .B1(n3422), .B2(n3908), .A(n3902), .ZN(n3535) );
  OAI21_X1 U2478 ( .B1(n3303), .B2(n3892), .A(n3909), .ZN(n3334) );
  INV_X1 U2479 ( .A(n3030), .ZN(n3038) );
  INV_X1 U2480 ( .A(n2542), .ZN(n2502) );
  NAND2_X1 U2481 ( .A1(n2808), .A2(n3880), .ZN(n2866) );
  NAND2_X1 U2482 ( .A1(n3093), .A2(n3816), .ZN(n4299) );
  CLKBUF_X3 U2483 ( .A(n2551), .Z(n2227) );
  AND2_X1 U2484 ( .A1(n3473), .A2(n3477), .ZN(n3471) );
  XNOR2_X1 U2485 ( .A(n2505), .B(IR_REG_1__SCAN_IN), .ZN(n2347) );
  NOR2_X1 U2486 ( .A1(n2519), .A2(n2518), .ZN(n4494) );
  INV_X4 U2487 ( .A(n2498), .ZN(n2625) );
  XNOR2_X2 U2488 ( .A(n2783), .B(n2782), .ZN(n2808) );
  OAI21_X1 U2489 ( .B1(n2861), .B2(n2860), .A(n4646), .ZN(n2862) );
  INV_X1 U2490 ( .A(n3655), .ZN(n3095) );
  OAI21_X1 U2491 ( .B1(n3660), .B2(n3661), .A(n3662), .ZN(n2978) );
  OAI22_X1 U2492 ( .A1(n2849), .A2(n2283), .B1(n2285), .B2(n3837), .ZN(n4104)
         );
  OR2_X1 U2493 ( .A1(n4260), .A2(n4143), .ZN(n4217) );
  AND2_X1 U2494 ( .A1(n2865), .A2(n3119), .ZN(n2242) );
  NAND2_X2 U2495 ( .A1(n3119), .A2(n2866), .ZN(n3040) );
  NAND2_X1 U2496 ( .A1(n2824), .A2(n3881), .ZN(n3350) );
  NAND3_X1 U2497 ( .A1(n2252), .A2(n2229), .A3(n2236), .ZN(n3881) );
  INV_X1 U2498 ( .A(n3311), .ZN(n2888) );
  NAND2_X2 U2499 ( .A1(n2499), .A2(n2477), .ZN(n2544) );
  XNOR2_X1 U2500 ( .A(n2474), .B(IR_REG_29__SCAN_IN), .ZN(n4484) );
  INV_X1 U2501 ( .A(n2243), .ZN(n2282) );
  AND2_X1 U2502 ( .A1(n2469), .A2(n2471), .ZN(n2339) );
  AND4_X1 U2503 ( .A1(n2468), .A2(n2467), .A3(n2466), .A4(n2484), .ZN(n2469)
         );
  NOR2_X1 U2504 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2470)
         );
  INV_X1 U2505 ( .A(IR_REG_3__SCAN_IN), .ZN(n2536) );
  NOR2_X1 U2506 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2468)
         );
  NOR2_X1 U2507 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2467)
         );
  NOR2_X1 U2508 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2466)
         );
  NOR2_X2 U2509 ( .A1(n3437), .A2(n3438), .ZN(n3473) );
  NOR2_X2 U2510 ( .A1(n4096), .A2(n4305), .ZN(n4072) );
  OR2_X2 U2511 ( .A1(n4112), .A2(n3774), .ZN(n4096) );
  BUF_X4 U2512 ( .A(n2551), .Z(n2228) );
  NOR2_X1 U2513 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2464)
         );
  NOR2_X1 U2514 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2408)
         );
  NOR2_X1 U2515 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2407)
         );
  NAND2_X1 U2516 ( .A1(n2434), .A2(n2433), .ZN(n2432) );
  INV_X1 U2517 ( .A(n3020), .ZN(n2434) );
  NAND2_X1 U2518 ( .A1(n2312), .A2(n2311), .ZN(n4070) );
  AOI21_X1 U2519 ( .B1(n2314), .B2(n2316), .A(n2260), .ZN(n2311) );
  AND2_X1 U2520 ( .A1(n2337), .A2(n2687), .ZN(n2336) );
  INV_X1 U2521 ( .A(n4199), .ZN(n2337) );
  NAND2_X1 U2522 ( .A1(n2392), .A2(n2400), .ZN(n2398) );
  INV_X1 U2523 ( .A(n2401), .ZN(n2392) );
  NAND2_X1 U2524 ( .A1(n3334), .A2(n3890), .ZN(n2829) );
  NAND2_X1 U2525 ( .A1(n2540), .A2(n3628), .ZN(n3891) );
  AND2_X1 U2526 ( .A1(n3378), .A2(n3375), .ZN(n3300) );
  OR2_X1 U2527 ( .A1(n3978), .A2(n3351), .ZN(n3882) );
  NAND2_X1 U2528 ( .A1(n2470), .A2(n2301), .ZN(n2300) );
  INV_X1 U2529 ( .A(IR_REG_25__SCAN_IN), .ZN(n2301) );
  NAND2_X1 U2530 ( .A1(n3291), .A2(n3290), .ZN(n2400) );
  NAND2_X1 U2531 ( .A1(n2932), .A2(n2233), .ZN(n2404) );
  NAND2_X1 U2532 ( .A1(n3729), .A2(n2433), .ZN(n2431) );
  NAND2_X1 U2533 ( .A1(n2257), .A2(n2418), .ZN(n2417) );
  INV_X1 U2534 ( .A(n3682), .ZN(n2418) );
  NAND2_X1 U2535 ( .A1(n2381), .A2(n2383), .ZN(n3758) );
  AOI21_X1 U2536 ( .B1(n2386), .B2(n2385), .A(n2384), .ZN(n2383) );
  INV_X1 U2537 ( .A(n3720), .ZN(n2384) );
  NAND2_X1 U2538 ( .A1(n2906), .A2(n2907), .ZN(n2912) );
  INV_X1 U2539 ( .A(n3729), .ZN(n2430) );
  NOR2_X1 U2540 ( .A1(n2499), .A2(n4484), .ZN(n2513) );
  NAND2_X1 U2541 ( .A1(n4534), .A2(n4535), .ZN(n4533) );
  NOR2_X1 U2542 ( .A1(n2600), .A2(n2599), .ZN(n2601) );
  NAND2_X1 U2543 ( .A1(n2832), .A2(n3899), .ZN(n3422) );
  INV_X1 U2544 ( .A(n3975), .ZN(n3478) );
  AND2_X1 U2545 ( .A1(n2808), .A2(n3204), .ZN(n4710) );
  OR2_X1 U2546 ( .A1(n3209), .A2(n4487), .ZN(n4705) );
  INV_X1 U2547 ( .A(IR_REG_28__SCAN_IN), .ZN(n2816) );
  AND2_X1 U2548 ( .A1(n2454), .A2(n2465), .ZN(n2405) );
  INV_X1 U2549 ( .A(IR_REG_13__SCAN_IN), .ZN(n2465) );
  INV_X1 U2550 ( .A(n4108), .ZN(n4157) );
  AOI21_X1 U2551 ( .B1(n3078), .B2(n3832), .A(n2771), .ZN(n2778) );
  AND2_X1 U2552 ( .A1(n3966), .A2(n3653), .ZN(n2771) );
  NOR2_X1 U2553 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2406)
         );
  INV_X1 U2554 ( .A(n3504), .ZN(n2442) );
  INV_X1 U2555 ( .A(n4505), .ZN(n2389) );
  OR2_X1 U2556 ( .A1(n3464), .A2(n3463), .ZN(n2447) );
  AND2_X1 U2557 ( .A1(n2387), .A2(n2268), .ZN(n2385) );
  INV_X1 U2558 ( .A(n3040), .ZN(n2878) );
  INV_X1 U2559 ( .A(n2882), .ZN(n3033) );
  AND2_X1 U2560 ( .A1(n4309), .A2(n3653), .ZN(n3819) );
  NAND2_X1 U2561 ( .A1(n3236), .A2(n3155), .ZN(n3156) );
  NAND2_X1 U2562 ( .A1(n3233), .A2(n2341), .ZN(n2340) );
  NAND2_X1 U2563 ( .A1(n4494), .A2(REG2_REG_2__SCAN_IN), .ZN(n2341) );
  NAND2_X1 U2564 ( .A1(n4491), .A2(REG1_REG_5__SCAN_IN), .ZN(n2361) );
  AND2_X1 U2565 ( .A1(n4092), .A2(n4305), .ZN(n3818) );
  NAND2_X1 U2566 ( .A1(n4104), .A2(n3858), .ZN(n4088) );
  INV_X1 U2567 ( .A(n3807), .ZN(n2287) );
  AND2_X1 U2568 ( .A1(n2707), .A2(n2333), .ZN(n2332) );
  NOR2_X1 U2569 ( .A1(n2706), .A2(n2705), .ZN(n2707) );
  NAND2_X1 U2570 ( .A1(n2334), .A2(n2336), .ZN(n2333) );
  INV_X1 U2571 ( .A(n2336), .ZN(n2335) );
  OAI21_X1 U2572 ( .B1(n2623), .B2(n2305), .A(n2460), .ZN(n2304) );
  AND2_X1 U2573 ( .A1(n3515), .A2(n3918), .ZN(n3591) );
  INV_X1 U2574 ( .A(n3847), .ZN(n2623) );
  INV_X1 U2575 ( .A(n2521), .ZN(n2308) );
  NAND2_X1 U2576 ( .A1(n3891), .A2(n3888), .ZN(n3375) );
  NAND2_X1 U2577 ( .A1(n3882), .A2(n3885), .ZN(n2825) );
  INV_X1 U2578 ( .A(n3254), .ZN(n3206) );
  NAND2_X1 U2579 ( .A1(n2673), .A2(n2672), .ZN(n2683) );
  NOR2_X1 U2580 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2672)
         );
  INV_X1 U2581 ( .A(n2671), .ZN(n2673) );
  INV_X1 U2582 ( .A(IR_REG_4__SCAN_IN), .ZN(n2463) );
  OR3_X1 U2583 ( .A1(n2593), .A2(IR_REG_8__SCAN_IN), .A3(IR_REG_7__SCAN_IN), 
        .ZN(n2610) );
  NOR2_X2 U2584 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2516)
         );
  OAI21_X1 U2585 ( .B1(n3769), .B2(n3772), .A(n3770), .ZN(n3635) );
  NAND2_X1 U2586 ( .A1(n3257), .A2(n2242), .ZN(n2380) );
  AND2_X1 U2587 ( .A1(n2866), .A2(n2870), .ZN(n3030) );
  AND2_X1 U2588 ( .A1(n3464), .A2(n3463), .ZN(n2445) );
  AND2_X1 U2589 ( .A1(n2257), .A2(n3761), .ZN(n2419) );
  NOR2_X1 U2590 ( .A1(n3503), .A2(n2445), .ZN(n2444) );
  OAI22_X1 U2591 ( .A1(n4403), .A2(n2882), .B1(n2955), .B2(n3599), .ZN(n3550)
         );
  INV_X1 U2592 ( .A(n2912), .ZN(n2909) );
  OAI21_X1 U2593 ( .B1(n2428), .B2(n2423), .A(n2425), .ZN(n2422) );
  INV_X1 U2594 ( .A(n2435), .ZN(n2423) );
  AOI21_X1 U2595 ( .B1(n2429), .B2(n2427), .A(n2426), .ZN(n2425) );
  OR3_X1 U2596 ( .A1(n2745), .A2(n3703), .A3(n2744), .ZN(n2753) );
  OR2_X1 U2597 ( .A1(n2641), .A2(n4847), .ZN(n2652) );
  AND2_X1 U2598 ( .A1(n4057), .A2(n4487), .ZN(n3061) );
  NAND3_X1 U2599 ( .A1(n4485), .A2(n3121), .A3(n4486), .ZN(n3119) );
  XNOR2_X1 U2600 ( .A(n2340), .B(n3143), .ZN(n3994) );
  NAND2_X1 U2601 ( .A1(n3271), .A2(REG1_REG_4__SCAN_IN), .ZN(n3270) );
  NAND2_X1 U2602 ( .A1(n2364), .A2(n2363), .ZN(n2362) );
  INV_X1 U2603 ( .A(n3168), .ZN(n2363) );
  XNOR2_X1 U2604 ( .A(n2360), .B(n4490), .ZN(n3183) );
  NAND2_X1 U2605 ( .A1(n2366), .A2(n2365), .ZN(n4030) );
  NAND2_X1 U2606 ( .A1(n2367), .A2(REG1_REG_7__SCAN_IN), .ZN(n2365) );
  OAI21_X1 U2607 ( .B1(n2367), .B2(REG1_REG_7__SCAN_IN), .A(n4489), .ZN(n2366)
         );
  XNOR2_X1 U2608 ( .A(n4004), .B(n4685), .ZN(n4525) );
  NAND2_X1 U2609 ( .A1(n4533), .A2(n4033), .ZN(n4034) );
  NAND2_X1 U2610 ( .A1(n4558), .A2(n4559), .ZN(n4557) );
  XNOR2_X1 U2611 ( .A(n4010), .B(n4037), .ZN(n4568) );
  NAND2_X1 U2612 ( .A1(n4554), .A2(n2259), .ZN(n4038) );
  XNOR2_X1 U2613 ( .A(n4012), .B(n2368), .ZN(n4588) );
  NAND2_X1 U2614 ( .A1(n4581), .A2(n4040), .ZN(n4042) );
  OR2_X1 U2615 ( .A1(n4588), .A2(n3563), .ZN(n2354) );
  INV_X1 U2616 ( .A(n2377), .ZN(n2376) );
  OAI22_X1 U2617 ( .A1(n4070), .A2(n2761), .B1(n4092), .B2(n4075), .ZN(n3078)
         );
  NOR2_X1 U2618 ( .A1(n2742), .A2(n2319), .ZN(n2318) );
  INV_X1 U2619 ( .A(n2734), .ZN(n2319) );
  NAND2_X1 U2620 ( .A1(n2266), .A2(n2321), .ZN(n2317) );
  AOI21_X1 U2621 ( .B1(n4141), .B2(n2726), .A(n2725), .ZN(n4120) );
  AOI21_X1 U2622 ( .B1(n2324), .B2(n2649), .A(n2263), .ZN(n2323) );
  NAND2_X1 U2623 ( .A1(n2327), .A2(n2650), .ZN(n2326) );
  INV_X1 U2624 ( .A(n3588), .ZN(n2327) );
  OR2_X1 U2625 ( .A1(n2639), .A2(n2638), .ZN(n2641) );
  OR2_X1 U2626 ( .A1(n3441), .A2(n3896), .ZN(n2831) );
  NOR2_X1 U2627 ( .A1(n2555), .A2(n3179), .ZN(n2566) );
  NAND2_X1 U2628 ( .A1(n2566), .A2(REG3_REG_7__SCAN_IN), .ZN(n2586) );
  AND2_X1 U2629 ( .A1(n3332), .A2(n2248), .ZN(n2562) );
  NAND2_X1 U2630 ( .A1(n2828), .A2(n3891), .ZN(n3303) );
  NOR2_X1 U2631 ( .A1(n2856), .A2(n2816), .ZN(n2487) );
  AND2_X1 U2632 ( .A1(n3257), .A2(n3206), .ZN(n3250) );
  OR2_X1 U2633 ( .A1(n4705), .A2(n3880), .ZN(n3085) );
  AND2_X1 U2634 ( .A1(n2818), .A2(n3873), .ZN(n3204) );
  INV_X1 U2635 ( .A(n4350), .ZN(n4205) );
  AND2_X1 U2636 ( .A1(n4229), .A2(n4205), .ZN(n4203) );
  OR2_X1 U2637 ( .A1(n4265), .A2(n4248), .ZN(n4244) );
  NOR2_X2 U2638 ( .A1(n4244), .A2(n4224), .ZN(n4229) );
  NAND2_X1 U2639 ( .A1(n4495), .A2(n3134), .ZN(n4402) );
  AND2_X1 U2640 ( .A1(n2803), .A2(n4485), .ZN(n3125) );
  AND2_X1 U2641 ( .A1(n2339), .A2(n2296), .ZN(n2295) );
  AND2_X1 U2642 ( .A1(n2338), .A2(n2816), .ZN(n2296) );
  INV_X1 U2643 ( .A(IR_REG_27__SCAN_IN), .ZN(n2338) );
  NOR2_X1 U2644 ( .A1(n2784), .A2(n2449), .ZN(n2798) );
  INV_X1 U2645 ( .A(IR_REG_23__SCAN_IN), .ZN(n2806) );
  INV_X1 U2646 ( .A(IR_REG_19__SCAN_IN), .ZN(n2779) );
  INV_X1 U2647 ( .A(n2516), .ZN(n2371) );
  NAND2_X1 U2648 ( .A1(n3289), .A2(n2401), .ZN(n2397) );
  AND2_X1 U2649 ( .A1(n2395), .A2(n2926), .ZN(n2394) );
  INV_X1 U2650 ( .A(n4497), .ZN(n3786) );
  NAND2_X1 U2651 ( .A1(n2410), .A2(n2409), .ZN(n3747) );
  AOI21_X1 U2652 ( .B1(n2412), .B2(n2415), .A(n2264), .ZN(n2409) );
  NAND2_X1 U2653 ( .A1(n2417), .A2(n2416), .ZN(n2415) );
  OR2_X1 U2654 ( .A1(n3068), .A2(n3066), .ZN(n3777) );
  NAND2_X1 U2655 ( .A1(n2733), .A2(n2732), .ZN(n4108) );
  INV_X1 U2656 ( .A(n4403), .ZN(n3969) );
  NAND2_X1 U2657 ( .A1(n2234), .A2(n2515), .ZN(n3978) );
  NAND2_X1 U2658 ( .A1(n2499), .A2(n2232), .ZN(n2297) );
  XNOR2_X1 U2659 ( .A(n4034), .B(n2359), .ZN(n4551) );
  NAND2_X1 U2660 ( .A1(n4555), .A2(n4556), .ZN(n4554) );
  XNOR2_X1 U2661 ( .A(n4038), .B(n4037), .ZN(n4566) );
  NAND2_X1 U2662 ( .A1(n4566), .A2(REG1_REG_12__SCAN_IN), .ZN(n4565) );
  NAND2_X1 U2663 ( .A1(n4626), .A2(n4627), .ZN(n2358) );
  OR2_X1 U2664 ( .A1(n4620), .A2(n2377), .ZN(n4630) );
  NOR2_X1 U2665 ( .A1(n4620), .A2(n4050), .ZN(n4632) );
  AOI21_X1 U2666 ( .B1(n4629), .B2(ADDR_REG_18__SCAN_IN), .A(n4628), .ZN(n2355) );
  NOR2_X1 U2667 ( .A1(n4626), .A2(n4627), .ZN(n4625) );
  NAND2_X1 U2668 ( .A1(n3107), .A2(n2289), .ZN(n3108) );
  INV_X1 U2669 ( .A(n2290), .ZN(n2289) );
  OAI21_X1 U2670 ( .B1(n4309), .B2(n4407), .A(n3106), .ZN(n2290) );
  INV_X2 U2671 ( .A(n4711), .ZN(n4713) );
  INV_X1 U2672 ( .A(n3839), .ZN(n2706) );
  INV_X1 U2673 ( .A(n2431), .ZN(n2427) );
  INV_X1 U2674 ( .A(n3699), .ZN(n2426) );
  NAND2_X1 U2675 ( .A1(n4536), .A2(n4006), .ZN(n4007) );
  NOR2_X1 U2676 ( .A1(n2753), .A2(n4981), .ZN(n2762) );
  AOI21_X1 U2677 ( .B1(n2315), .B2(n2317), .A(n2262), .ZN(n2314) );
  INV_X1 U2678 ( .A(n2318), .ZN(n2315) );
  INV_X1 U2679 ( .A(n2317), .ZN(n2316) );
  OR2_X1 U2680 ( .A1(n4366), .A2(n4248), .ZN(n2687) );
  AND2_X1 U2681 ( .A1(n3608), .A2(n3585), .ZN(n3919) );
  OR2_X1 U2682 ( .A1(n3425), .A2(n2600), .ZN(n2595) );
  NAND2_X1 U2683 ( .A1(n2830), .A2(n3900), .ZN(n3440) );
  NAND2_X1 U2684 ( .A1(n2520), .A2(n2825), .ZN(n3347) );
  INV_X1 U2685 ( .A(n3819), .ZN(n2854) );
  NAND2_X1 U2686 ( .A1(n4886), .A2(n2450), .ZN(n2449) );
  INV_X1 U2687 ( .A(IR_REG_21__SCAN_IN), .ZN(n2450) );
  INV_X1 U2688 ( .A(IR_REG_20__SCAN_IN), .ZN(n2782) );
  INV_X1 U2689 ( .A(IR_REG_18__SCAN_IN), .ZN(n5006) );
  INV_X1 U2690 ( .A(IR_REG_17__SCAN_IN), .ZN(n2684) );
  INV_X1 U2691 ( .A(n2683), .ZN(n2685) );
  INV_X1 U2692 ( .A(IR_REG_15__SCAN_IN), .ZN(n2484) );
  INV_X1 U2693 ( .A(IR_REG_14__SCAN_IN), .ZN(n2483) );
  INV_X1 U2694 ( .A(IR_REG_7__SCAN_IN), .ZN(n2579) );
  INV_X1 U2695 ( .A(IR_REG_6__SCAN_IN), .ZN(n2573) );
  OR2_X1 U2696 ( .A1(n3291), .A2(n3290), .ZN(n2401) );
  NOR2_X1 U2697 ( .A1(n2442), .A2(n2438), .ZN(n2437) );
  INV_X1 U2698 ( .A(n2447), .ZN(n2438) );
  INV_X1 U2699 ( .A(n2441), .ZN(n2440) );
  OAI21_X1 U2700 ( .B1(n2444), .B2(n2442), .A(n3551), .ZN(n2441) );
  INV_X1 U2701 ( .A(n4342), .ZN(n3677) );
  XNOR2_X1 U2702 ( .A(n2887), .B(n3038), .ZN(n2898) );
  AND2_X1 U2703 ( .A1(n2398), .A2(n3365), .ZN(n2393) );
  INV_X1 U2704 ( .A(n2400), .ZN(n2399) );
  OR2_X1 U2705 ( .A1(n2708), .A2(n3692), .ZN(n2716) );
  NAND2_X1 U2706 ( .A1(n2265), .A2(n2979), .ZN(n2387) );
  NAND2_X1 U2707 ( .A1(n2267), .A2(n2979), .ZN(n2386) );
  OR2_X1 U2708 ( .A1(n2977), .A2(n2389), .ZN(n2388) );
  INV_X1 U2709 ( .A(n4507), .ZN(n2390) );
  AND2_X1 U2710 ( .A1(n2413), .A2(n2457), .ZN(n2412) );
  INV_X1 U2711 ( .A(n2419), .ZN(n2414) );
  INV_X1 U2712 ( .A(n3689), .ZN(n3005) );
  INV_X1 U2713 ( .A(n3688), .ZN(n3006) );
  NAND2_X1 U2714 ( .A1(n2777), .A2(DATAI_22_), .ZN(n3752) );
  NOR2_X1 U2715 ( .A1(n2403), .A2(n3454), .ZN(n2402) );
  INV_X1 U2716 ( .A(n2943), .ZN(n2403) );
  NAND2_X1 U2717 ( .A1(n2880), .A2(n2879), .ZN(n2881) );
  NAND2_X1 U2718 ( .A1(n3978), .A2(n2877), .ZN(n2880) );
  NAND2_X1 U2719 ( .A1(n2541), .A2(REG3_REG_5__SCAN_IN), .ZN(n2555) );
  INV_X1 U2720 ( .A(n4097), .ZN(n3774) );
  NAND2_X1 U2721 ( .A1(n2978), .A2(n2977), .ZN(n4504) );
  INV_X1 U2722 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2651) );
  INV_X1 U2723 ( .A(n2544), .ZN(n2512) );
  NAND2_X1 U2724 ( .A1(n2502), .A2(n2522), .ZN(n2524) );
  INV_X1 U2725 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2298) );
  NAND2_X1 U2726 ( .A1(n3270), .A2(n3159), .ZN(n2364) );
  AOI21_X1 U2727 ( .B1(n3994), .B2(REG2_REG_3__SCAN_IN), .A(n2246), .ZN(n3144)
         );
  OR2_X1 U2728 ( .A1(n3181), .A2(n2249), .ZN(n2367) );
  AOI21_X1 U2729 ( .B1(REG2_REG_5__SCAN_IN), .B2(n4491), .A(n3170), .ZN(n3146)
         );
  OR2_X1 U2730 ( .A1(n4003), .A2(n4002), .ZN(n4004) );
  NAND2_X1 U2731 ( .A1(n4525), .A2(REG2_REG_8__SCAN_IN), .ZN(n4524) );
  NAND2_X1 U2732 ( .A1(n4529), .A2(n4032), .ZN(n4534) );
  XNOR2_X1 U2733 ( .A(n4007), .B(n2359), .ZN(n4546) );
  NAND2_X1 U2734 ( .A1(n4546), .A2(REG2_REG_10__SCAN_IN), .ZN(n4545) );
  NAND2_X1 U2735 ( .A1(n4557), .A2(n4009), .ZN(n4010) );
  NAND2_X1 U2736 ( .A1(n4568), .A2(REG2_REG_12__SCAN_IN), .ZN(n4567) );
  INV_X1 U2737 ( .A(n4596), .ZN(n2350) );
  OR2_X1 U2738 ( .A1(n4588), .A2(n2352), .ZN(n2351) );
  OR2_X1 U2739 ( .A1(n4596), .A2(n3563), .ZN(n2352) );
  AND2_X1 U2740 ( .A1(n2348), .A2(n2351), .ZN(n4015) );
  AND2_X1 U2741 ( .A1(n2349), .A2(n4014), .ZN(n2348) );
  NAND2_X1 U2742 ( .A1(n4633), .A2(n2378), .ZN(n2377) );
  INV_X1 U2743 ( .A(n4050), .ZN(n2378) );
  NOR2_X1 U2744 ( .A1(n2377), .A2(n2375), .ZN(n2374) );
  INV_X1 U2745 ( .A(n4618), .ZN(n2375) );
  AOI21_X1 U2746 ( .B1(n4088), .B2(n3945), .A(n3834), .ZN(n4068) );
  NOR2_X1 U2747 ( .A1(n3943), .A2(n3818), .ZN(n4071) );
  OR2_X1 U2748 ( .A1(n2287), .A2(n3837), .ZN(n2283) );
  INV_X1 U2749 ( .A(n2286), .ZN(n2285) );
  OAI21_X1 U2750 ( .B1(n2287), .B2(n2848), .A(n3937), .ZN(n2286) );
  NAND2_X1 U2751 ( .A1(n2284), .A2(n3807), .ZN(n4123) );
  NAND2_X1 U2752 ( .A1(n2849), .A2(n2848), .ZN(n2284) );
  NOR2_X1 U2753 ( .A1(n2716), .A2(n3750), .ZN(n2721) );
  NAND2_X1 U2754 ( .A1(n2331), .A2(n2329), .ZN(n4183) );
  AOI21_X1 U2755 ( .B1(n2332), .B2(n2335), .A(n2330), .ZN(n2329) );
  INV_X1 U2756 ( .A(n3840), .ZN(n2330) );
  AND2_X1 U2757 ( .A1(n2688), .A2(REG3_REG_19__SCAN_IN), .ZN(n2697) );
  NAND2_X1 U2758 ( .A1(n4240), .A2(n2687), .ZN(n4215) );
  AND4_X1 U2759 ( .A1(n2682), .A2(n2681), .A3(n2680), .A4(n2679), .ZN(n4228)
         );
  AND4_X1 U2760 ( .A1(n2670), .A2(n2669), .A3(n2668), .A4(n2667), .ZN(n4286)
         );
  NOR2_X1 U2761 ( .A1(n2677), .A2(n4623), .ZN(n2688) );
  INV_X1 U2762 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4623) );
  NAND2_X1 U2763 ( .A1(n4242), .A2(n4241), .ZN(n4240) );
  NAND2_X1 U2764 ( .A1(n2626), .A2(REG3_REG_12__SCAN_IN), .ZN(n2639) );
  NAND2_X1 U2765 ( .A1(n3598), .A2(n4400), .ZN(n2636) );
  INV_X1 U2766 ( .A(n2304), .ZN(n2303) );
  NAND2_X1 U2767 ( .A1(n3535), .A2(n3917), .ZN(n2835) );
  AND2_X1 U2768 ( .A1(n3589), .A2(n3918), .ZN(n3847) );
  OR2_X1 U2769 ( .A1(n2586), .A2(n2475), .ZN(n2603) );
  NOR2_X1 U2770 ( .A1(n2603), .A2(n4848), .ZN(n2613) );
  NAND2_X1 U2771 ( .A1(n3440), .A2(n2583), .ZN(n3425) );
  INV_X1 U2772 ( .A(n2596), .ZN(n2583) );
  AND2_X1 U2773 ( .A1(n2598), .A2(n2597), .ZN(n3426) );
  OR2_X1 U2774 ( .A1(n2596), .A2(n3474), .ZN(n2598) );
  INV_X1 U2775 ( .A(n3440), .ZN(n3846) );
  NAND2_X1 U2776 ( .A1(n2461), .A2(n2554), .ZN(n3332) );
  AND2_X1 U2777 ( .A1(n2307), .A2(n2554), .ZN(n2309) );
  NAND2_X1 U2778 ( .A1(n2308), .A2(n2527), .ZN(n2307) );
  AOI21_X1 U2779 ( .B1(n3280), .B2(n3849), .A(n2827), .ZN(n3376) );
  AND2_X1 U2780 ( .A1(n3887), .A2(n3884), .ZN(n3849) );
  NAND2_X1 U2781 ( .A1(n3347), .A2(n2521), .ZN(n3279) );
  INV_X1 U2782 ( .A(n2825), .ZN(n3851) );
  INV_X1 U2783 ( .A(n4289), .ZN(n3522) );
  INV_X1 U2784 ( .A(n3811), .ZN(n4302) );
  AOI21_X1 U2785 ( .B1(n2292), .B2(n4289), .A(n2291), .ZN(n3107) );
  AND2_X1 U2786 ( .A1(n3964), .A2(n4062), .ZN(n2291) );
  XNOR2_X1 U2787 ( .A(n2294), .B(n2293), .ZN(n2292) );
  OAI21_X1 U2788 ( .B1(n3080), .B2(n3815), .A(n2854), .ZN(n2294) );
  NOR2_X1 U2789 ( .A1(n2228), .A2(n2760), .ZN(n4305) );
  NAND2_X1 U2790 ( .A1(n4127), .A2(n4113), .ZN(n4112) );
  NOR2_X1 U2791 ( .A1(n4158), .A2(n4322), .ZN(n4127) );
  INV_X1 U2792 ( .A(n4134), .ZN(n4322) );
  NAND2_X1 U2793 ( .A1(n2280), .A2(n4159), .ZN(n4158) );
  NAND2_X1 U2794 ( .A1(n4203), .A2(n4190), .ZN(n4185) );
  NOR2_X1 U2795 ( .A1(n2228), .A2(n2704), .ZN(n4350) );
  NAND2_X1 U2796 ( .A1(n4282), .A2(n2258), .ZN(n4265) );
  AND2_X1 U2797 ( .A1(n4282), .A2(n4499), .ZN(n4280) );
  AND4_X1 U2798 ( .A1(n2497), .A2(n2496), .A3(n2495), .A4(n2494), .ZN(n4382)
         );
  AND4_X1 U2799 ( .A1(n2645), .A2(n2644), .A3(n2643), .A4(n2642), .ZN(n4403)
         );
  OR2_X1 U2800 ( .A1(n3530), .A2(n3456), .ZN(n3531) );
  NAND2_X1 U2801 ( .A1(n3471), .A2(n3489), .ZN(n3530) );
  INV_X1 U2802 ( .A(n3429), .ZN(n3489) );
  AND4_X1 U2803 ( .A1(n2578), .A2(n2577), .A3(n2576), .A4(n2575), .ZN(n3493)
         );
  NAND2_X1 U2804 ( .A1(n2279), .A2(n2278), .ZN(n3437) );
  INV_X1 U2805 ( .A(n3978), .ZN(n3312) );
  NAND2_X1 U2806 ( .A1(n3517), .A2(n4705), .ZN(n4411) );
  AND2_X1 U2807 ( .A1(n4488), .A2(n3204), .ZN(n4386) );
  NAND2_X1 U2808 ( .A1(n3226), .A2(n3134), .ZN(n4407) );
  INV_X1 U2809 ( .A(n3089), .ZN(n3098) );
  NAND2_X1 U2810 ( .A1(n2299), .A2(n2470), .ZN(n2448) );
  INV_X1 U2811 ( .A(n2449), .ZN(n2299) );
  AND3_X1 U2812 ( .A1(n2231), .A2(n2518), .A3(n2454), .ZN(n2646) );
  XNOR2_X1 U2813 ( .A(n2923), .B(n2924), .ZN(n3365) );
  NAND2_X1 U2814 ( .A1(n2404), .A2(n2943), .ZN(n3453) );
  NAND2_X1 U2815 ( .A1(n3757), .A2(n3761), .ZN(n3683) );
  NAND2_X1 U2816 ( .A1(n2380), .A2(n2379), .ZN(n2871) );
  AND2_X1 U2817 ( .A1(n3030), .A2(n2230), .ZN(n2379) );
  INV_X1 U2818 ( .A(n2445), .ZN(n2443) );
  NAND2_X1 U2819 ( .A1(n3672), .A2(n2431), .ZN(n2424) );
  AND4_X1 U2820 ( .A1(n2659), .A2(n2658), .A3(n2657), .A4(n2656), .ZN(n4498)
         );
  INV_X1 U2821 ( .A(n2662), .ZN(n4499) );
  NAND2_X1 U2822 ( .A1(n2382), .A2(n2386), .ZN(n3722) );
  OR2_X1 U2823 ( .A1(n2978), .A2(n2387), .ZN(n2382) );
  OAI21_X1 U2824 ( .B1(n3672), .B2(n3020), .A(n3019), .ZN(n3728) );
  NAND2_X1 U2825 ( .A1(n2228), .A2(IR_REG_0__SCAN_IN), .ZN(n2273) );
  NAND2_X1 U2826 ( .A1(n2275), .A2(DATAI_0_), .ZN(n2274) );
  INV_X1 U2827 ( .A(n2227), .ZN(n2275) );
  INV_X1 U2828 ( .A(n3785), .ZN(n4500) );
  NAND2_X1 U2829 ( .A1(n2411), .A2(n2417), .ZN(n3739) );
  NAND2_X1 U2830 ( .A1(n3757), .A2(n2419), .ZN(n2411) );
  NAND2_X1 U2831 ( .A1(n2446), .A2(n2444), .ZN(n2439) );
  OR2_X1 U2832 ( .A1(n3068), .A2(n3065), .ZN(n4497) );
  OR2_X1 U2833 ( .A1(n3625), .A2(n2914), .ZN(n2916) );
  AND2_X1 U2834 ( .A1(n2759), .A2(n2758), .ZN(n4092) );
  INV_X1 U2835 ( .A(n2422), .ZN(n2421) );
  AND2_X1 U2836 ( .A1(n3051), .A2(n3050), .ZN(n4508) );
  INV_X1 U2837 ( .A(n4092), .ZN(n3967) );
  NAND2_X1 U2838 ( .A1(n2752), .A2(n2751), .ZN(n4306) );
  NAND2_X1 U2839 ( .A1(n2741), .A2(n2740), .ZN(n4136) );
  OR2_X1 U2840 ( .A1(n2544), .A2(n4160), .ZN(n2723) );
  NAND4_X1 U2841 ( .A1(n2693), .A2(n2692), .A3(n2691), .A4(n2690), .ZN(n4249)
         );
  INV_X1 U2842 ( .A(n4228), .ZN(n4366) );
  INV_X1 U2843 ( .A(n4286), .ZN(n4502) );
  INV_X1 U2844 ( .A(n4369), .ZN(n4379) );
  INV_X1 U2845 ( .A(n4382), .ZN(n3968) );
  INV_X1 U2846 ( .A(n3493), .ZN(n3974) );
  NAND3_X1 U2847 ( .A1(n2572), .A2(n2571), .A3(n2570), .ZN(n3975) );
  OR2_X1 U2848 ( .A1(n2542), .A2(n3446), .ZN(n2572) );
  NAND4_X1 U2849 ( .A1(n2560), .A2(n2559), .A3(n2558), .A4(n2557), .ZN(n3976)
         );
  OR2_X1 U2850 ( .A1(n2542), .A2(n3211), .ZN(n2509) );
  OR2_X1 U2851 ( .A1(n3119), .A2(n3118), .ZN(n3979) );
  OAI21_X1 U2852 ( .B1(n2347), .B2(n3139), .A(n2342), .ZN(n3985) );
  NAND2_X1 U2853 ( .A1(n3234), .A2(n3235), .ZN(n3233) );
  INV_X1 U2854 ( .A(n2362), .ZN(n3167) );
  INV_X1 U2855 ( .A(n2364), .ZN(n3169) );
  INV_X1 U2856 ( .A(n2367), .ZN(n4029) );
  NOR2_X1 U2857 ( .A1(n3151), .A2(n3150), .ZN(n4003) );
  XOR2_X1 U2858 ( .A(n4031), .B(n4030), .Z(n4530) );
  NAND2_X1 U2859 ( .A1(n4537), .A2(n4538), .ZN(n4536) );
  NAND2_X1 U2860 ( .A1(n4550), .A2(n4035), .ZN(n4555) );
  NAND2_X1 U2861 ( .A1(n4565), .A2(n4039), .ZN(n4582) );
  NAND2_X1 U2862 ( .A1(n4582), .A2(n4583), .ZN(n4581) );
  XNOR2_X1 U2863 ( .A(n4042), .B(n2368), .ZN(n4592) );
  AND2_X1 U2864 ( .A1(n2354), .A2(n2353), .ZN(n4597) );
  XNOR2_X1 U2865 ( .A(n4015), .B(n4045), .ZN(n4606) );
  NAND2_X1 U2866 ( .A1(n4613), .A2(n4615), .ZN(n4614) );
  NOR2_X1 U2867 ( .A1(n2374), .A2(n2271), .ZN(n2373) );
  AND2_X1 U2868 ( .A1(n2770), .A2(n2769), .ZN(n4309) );
  NAND2_X1 U2869 ( .A1(n2313), .A2(n2317), .ZN(n4086) );
  NAND2_X1 U2870 ( .A1(n4120), .A2(n2318), .ZN(n2313) );
  NAND2_X1 U2871 ( .A1(n4120), .A2(n2734), .ZN(n2320) );
  NAND2_X1 U2872 ( .A1(n2777), .A2(DATAI_21_), .ZN(n4190) );
  INV_X1 U2873 ( .A(n4057), .ZN(n4253) );
  INV_X1 U2874 ( .A(n4378), .ZN(n3580) );
  AND2_X1 U2875 ( .A1(n2326), .A2(n2328), .ZN(n3559) );
  NAND2_X1 U2876 ( .A1(n2326), .A2(n2324), .ZN(n3558) );
  AND2_X1 U2877 ( .A1(n3542), .A2(n3541), .ZN(n4642) );
  NAND2_X1 U2878 ( .A1(n4646), .A2(n2821), .ZN(n4233) );
  INV_X1 U2879 ( .A(n2905), .ZN(n3977) );
  AND2_X1 U2880 ( .A1(n4646), .A2(n4323), .ZN(n4267) );
  OR2_X1 U2881 ( .A1(n2544), .A2(n2531), .ZN(n2533) );
  INV_X1 U2882 ( .A(n4295), .ZN(n4264) );
  INV_X1 U2883 ( .A(n4233), .ZN(n4657) );
  NAND2_X1 U2884 ( .A1(n2813), .A2(n3193), .ZN(n4643) );
  INV_X1 U2885 ( .A(n3085), .ZN(n2813) );
  OR2_X1 U2886 ( .A1(n3099), .A2(n3089), .ZN(n4719) );
  INV_X2 U2887 ( .A(n4719), .ZN(n4722) );
  OR2_X1 U2888 ( .A1(n3642), .A2(n2815), .ZN(n2472) );
  XNOR2_X1 U2889 ( .A(n2817), .B(n2816), .ZN(n4495) );
  XNOR2_X1 U2890 ( .A(n2802), .B(IR_REG_26__SCAN_IN), .ZN(n4485) );
  XNOR2_X1 U2891 ( .A(n2800), .B(IR_REG_24__SCAN_IN), .ZN(n4486) );
  AND2_X1 U2892 ( .A1(n3135), .A2(STATE_REG_SCAN_IN), .ZN(n4675) );
  XNOR2_X1 U2893 ( .A(n2786), .B(IR_REG_22__SCAN_IN), .ZN(n4487) );
  XNOR2_X1 U2894 ( .A(n2785), .B(IR_REG_21__SCAN_IN), .ZN(n3880) );
  NAND2_X1 U2895 ( .A1(n2370), .A2(n2369), .ZN(n2519) );
  NAND2_X1 U2896 ( .A1(n2815), .A2(n2462), .ZN(n2369) );
  NAND2_X1 U2897 ( .A1(n2356), .A2(n2238), .ZN(U3258) );
  OR2_X1 U2898 ( .A1(n2357), .A2(n4625), .ZN(n2356) );
  NAND2_X1 U2899 ( .A1(n2358), .A2(n4575), .ZN(n2357) );
  OR2_X1 U2900 ( .A1(n3115), .A2(n4414), .ZN(n3111) );
  NAND2_X1 U2901 ( .A1(n3095), .A2(n3094), .ZN(n3096) );
  NAND2_X1 U2902 ( .A1(n3095), .A2(n3102), .ZN(n3103) );
  NAND2_X1 U2903 ( .A1(n2344), .A2(n2343), .ZN(U3351) );
  NAND2_X1 U2904 ( .A1(U3149), .A2(DATAI_1_), .ZN(n2343) );
  NAND2_X1 U2905 ( .A1(n2502), .A2(REG3_REG_1__SCAN_IN), .ZN(n2229) );
  NAND2_X2 U2906 ( .A1(n2499), .A2(n4484), .ZN(n2542) );
  OR2_X1 U2907 ( .A1(n2526), .A2(n2451), .ZN(n2890) );
  OR2_X1 U2908 ( .A1(n3254), .A2(n3040), .ZN(n2230) );
  AND4_X1 U2909 ( .A1(n2464), .A2(n2408), .A3(n2407), .A4(n2406), .ZN(n2231)
         );
  AND4_X1 U2910 ( .A1(n2547), .A2(n2546), .A3(n2545), .A4(n2247), .ZN(n2905)
         );
  AND2_X1 U2911 ( .A1(n2477), .A2(REG2_REG_2__SCAN_IN), .ZN(n2232) );
  NOR2_X1 U2912 ( .A1(n3412), .A2(n2937), .ZN(n2233) );
  INV_X1 U2913 ( .A(n3336), .ZN(n2278) );
  AND3_X1 U2914 ( .A1(n2514), .A2(n2254), .A3(n2297), .ZN(n2234) );
  AND2_X1 U2915 ( .A1(n2320), .A2(n2256), .ZN(n2235) );
  AND2_X1 U2916 ( .A1(n2251), .A2(n2503), .ZN(n2236) );
  OR2_X1 U2917 ( .A1(n3672), .A2(n2432), .ZN(n2237) );
  AND3_X1 U2918 ( .A1(n4634), .A2(n2355), .A3(n2270), .ZN(n2238) );
  NOR2_X1 U2919 ( .A1(n2456), .A2(n2325), .ZN(n2324) );
  AND2_X1 U2920 ( .A1(n2230), .A2(n2261), .ZN(n2239) );
  INV_X1 U2921 ( .A(n2649), .ZN(n2650) );
  AND2_X1 U2922 ( .A1(n4403), .A2(n3599), .ZN(n2649) );
  NAND2_X1 U2923 ( .A1(n2306), .A2(n2623), .ZN(n3512) );
  AND2_X1 U2924 ( .A1(n2386), .A2(n2268), .ZN(n2240) );
  AND3_X1 U2925 ( .A1(n2282), .A2(n2482), .A3(n2272), .ZN(n2241) );
  OR2_X1 U2926 ( .A1(n2300), .A2(n2449), .ZN(n2243) );
  OR2_X1 U2927 ( .A1(n2499), .A2(n2477), .ZN(n2498) );
  NAND2_X1 U2928 ( .A1(n2362), .A2(n2361), .ZN(n2360) );
  NAND2_X1 U2929 ( .A1(n2424), .A2(n2429), .ZN(n3701) );
  NAND2_X1 U2930 ( .A1(n2516), .A2(n2462), .ZN(n2517) );
  AND2_X1 U2931 ( .A1(n3020), .A2(n3019), .ZN(n2244) );
  OR2_X1 U2932 ( .A1(n2784), .A2(IR_REG_21__SCAN_IN), .ZN(n2245) );
  AND2_X1 U2933 ( .A1(n2340), .A2(n4493), .ZN(n2246) );
  OR2_X1 U2934 ( .A1(n2544), .A2(n2543), .ZN(n2247) );
  NAND2_X1 U2935 ( .A1(n3976), .A2(n3336), .ZN(n2248) );
  AND2_X1 U2936 ( .A1(n2360), .A2(n4490), .ZN(n2249) );
  OR2_X1 U2937 ( .A1(n2784), .A2(n2243), .ZN(n2250) );
  NAND2_X1 U2938 ( .A1(n2696), .A2(IR_REG_31__SCAN_IN), .ZN(n2780) );
  INV_X1 U2939 ( .A(IR_REG_2__SCAN_IN), .ZN(n2462) );
  OR2_X1 U2940 ( .A1(n2501), .A2(n2500), .ZN(n2251) );
  AND2_X1 U2941 ( .A1(n2504), .A2(n3256), .ZN(n2252) );
  INV_X1 U2942 ( .A(n2429), .ZN(n2428) );
  AOI21_X1 U2943 ( .B1(n2432), .B2(n2430), .A(n2244), .ZN(n2429) );
  NAND2_X1 U2944 ( .A1(n3973), .A2(n3429), .ZN(n2253) );
  OR2_X1 U2945 ( .A1(n2542), .A2(n2298), .ZN(n2254) );
  INV_X1 U2946 ( .A(IR_REG_31__SCAN_IN), .ZN(n2815) );
  OR2_X1 U2947 ( .A1(n2784), .A2(n2448), .ZN(n2255) );
  INV_X1 U2948 ( .A(n3868), .ZN(n2325) );
  INV_X1 U2949 ( .A(n3856), .ZN(n2293) );
  NAND2_X1 U2950 ( .A1(n4157), .A2(n4134), .ZN(n2256) );
  NAND2_X1 U2951 ( .A1(n2439), .A2(n3504), .ZN(n3549) );
  NAND2_X1 U2952 ( .A1(n2446), .A2(n2443), .ZN(n3502) );
  NAND2_X1 U2953 ( .A1(n2993), .A2(n2992), .ZN(n2257) );
  INV_X1 U2954 ( .A(n4241), .ZN(n2334) );
  NAND2_X1 U2955 ( .A1(n2482), .A2(n2469), .ZN(n2784) );
  AND2_X1 U2956 ( .A1(n4499), .A2(n4273), .ZN(n2258) );
  INV_X1 U2957 ( .A(n2280), .ZN(n4176) );
  NOR2_X1 U2958 ( .A1(n4185), .A2(n4174), .ZN(n2280) );
  INV_X1 U2959 ( .A(n2624), .ZN(n2305) );
  OR2_X1 U2960 ( .A1(n4682), .A2(n4720), .ZN(n2259) );
  INV_X1 U2961 ( .A(n2742), .ZN(n2321) );
  OR2_X1 U2962 ( .A1(n2978), .A2(n2977), .ZN(n2391) );
  INV_X1 U2963 ( .A(n4408), .ZN(n3971) );
  AND4_X1 U2964 ( .A1(n2619), .A2(n2618), .A3(n2617), .A4(n2616), .ZN(n4408)
         );
  NOR2_X1 U2965 ( .A1(n4306), .A2(n3774), .ZN(n2260) );
  OR2_X1 U2966 ( .A1(n3119), .A2(n2867), .ZN(n2261) );
  NOR2_X1 U2967 ( .A1(n4111), .A2(n4097), .ZN(n2262) );
  NOR2_X1 U2968 ( .A1(n3968), .A2(n4387), .ZN(n2263) );
  AND2_X1 U2969 ( .A1(n3006), .A2(n3005), .ZN(n2264) );
  NAND2_X1 U2970 ( .A1(n2977), .A2(n2389), .ZN(n2265) );
  NAND2_X1 U2971 ( .A1(n2256), .A2(n2743), .ZN(n2266) );
  NAND2_X1 U2972 ( .A1(n2390), .A2(n2388), .ZN(n2267) );
  INV_X1 U2973 ( .A(n3837), .ZN(n2288) );
  NAND2_X1 U2974 ( .A1(n3279), .A2(n2527), .ZN(n3299) );
  INV_X1 U2975 ( .A(n2277), .ZN(n3523) );
  NOR2_X1 U2976 ( .A1(n3531), .A2(n3524), .ZN(n2277) );
  INV_X1 U2977 ( .A(n3736), .ZN(n2416) );
  NAND2_X1 U2978 ( .A1(n3512), .A2(n2624), .ZN(n3610) );
  OAI21_X1 U2979 ( .B1(n3624), .B2(n2916), .A(n2915), .ZN(n3289) );
  NAND2_X1 U2980 ( .A1(n2397), .A2(n2400), .ZN(n3364) );
  NAND2_X1 U2981 ( .A1(n3611), .A2(n3599), .ZN(n3601) );
  INV_X1 U2982 ( .A(n3601), .ZN(n2276) );
  INV_X1 U2983 ( .A(n4159), .ZN(n4154) );
  AOI21_X1 U2984 ( .B1(n3217), .B2(n2901), .A(n2900), .ZN(n3624) );
  NAND2_X1 U2985 ( .A1(n2982), .A2(n2981), .ZN(n2268) );
  INV_X1 U2986 ( .A(n2456), .ZN(n2328) );
  INV_X1 U2987 ( .A(n4041), .ZN(n2368) );
  NAND4_X1 U2988 ( .A1(n2509), .A2(n2508), .A3(n2507), .A4(n2506), .ZN(n3257)
         );
  NAND2_X1 U2989 ( .A1(n3333), .A2(n3332), .ZN(n2269) );
  INV_X1 U2990 ( .A(n3337), .ZN(n2279) );
  OR2_X1 U2991 ( .A1(n4635), .A2(n4676), .ZN(n2270) );
  INV_X1 U2992 ( .A(n4575), .ZN(n4624) );
  AND2_X1 U2993 ( .A1(n4520), .A2(n3959), .ZN(n4575) );
  NOR2_X1 U2994 ( .A1(n4676), .A2(n4051), .ZN(n2271) );
  AND2_X1 U2995 ( .A1(n2339), .A2(n2338), .ZN(n2272) );
  INV_X1 U2996 ( .A(n4544), .ZN(n2359) );
  INV_X1 U2997 ( .A(DATAI_1_), .ZN(n2346) );
  NOR2_X1 U2998 ( .A1(n2473), .A2(IR_REG_29__SCAN_IN), .ZN(n3642) );
  NOR2_X2 U2999 ( .A1(n3359), .A2(n3360), .ZN(n3358) );
  NAND2_X2 U3000 ( .A1(n3253), .A2(n3254), .ZN(n3359) );
  AND2_X2 U3001 ( .A1(n2274), .A2(n2273), .ZN(n3254) );
  NOR2_X2 U3002 ( .A1(n3523), .A2(n3617), .ZN(n3611) );
  NAND3_X1 U3004 ( .A1(n2482), .A2(n2339), .A3(n2282), .ZN(n2281) );
  AND3_X2 U3005 ( .A1(n2405), .A2(n2518), .A3(n2231), .ZN(n2482) );
  NAND3_X1 U3006 ( .A1(n2282), .A2(n2482), .A3(n2295), .ZN(n2473) );
  INV_X1 U3007 ( .A(n3513), .ZN(n2306) );
  NAND2_X1 U3008 ( .A1(n2302), .A2(n2303), .ZN(n2637) );
  NAND2_X1 U3009 ( .A1(n3513), .A2(n2624), .ZN(n2302) );
  NAND3_X1 U3010 ( .A1(n2236), .A2(n2229), .A3(n2504), .ZN(n2510) );
  INV_X1 U3011 ( .A(n2510), .ZN(n3352) );
  OAI22_X1 U3012 ( .A1(n3352), .A2(n2955), .B1(n3040), .B2(n3253), .ZN(n2872)
         );
  NAND3_X1 U3013 ( .A1(n2310), .A2(n2309), .A3(n3300), .ZN(n3333) );
  NAND3_X1 U3014 ( .A1(n2520), .A2(n2527), .A3(n2825), .ZN(n2310) );
  NAND2_X1 U3015 ( .A1(n4120), .A2(n2314), .ZN(n2312) );
  NAND2_X1 U3016 ( .A1(n3588), .A2(n2324), .ZN(n2322) );
  NAND2_X1 U3017 ( .A1(n2322), .A2(n2323), .ZN(n3573) );
  NAND2_X1 U3018 ( .A1(n4242), .A2(n2332), .ZN(n2331) );
  NAND2_X1 U3019 ( .A1(n2347), .A2(n3139), .ZN(n2342) );
  NAND2_X1 U3020 ( .A1(n2347), .A2(REG2_REG_1__SCAN_IN), .ZN(n3141) );
  NAND2_X1 U3021 ( .A1(n2347), .A2(REG1_REG_1__SCAN_IN), .ZN(n3154) );
  NAND2_X1 U3022 ( .A1(n2347), .A2(STATE_REG_SCAN_IN), .ZN(n2344) );
  XNOR2_X1 U3023 ( .A(n2347), .B(n3153), .ZN(n3982) );
  NAND2_X1 U3024 ( .A1(n2228), .A2(n2347), .ZN(n2345) );
  NAND2_X1 U3025 ( .A1(n3992), .A2(n2347), .ZN(n3987) );
  INV_X1 U3026 ( .A(n4013), .ZN(n2353) );
  NAND2_X1 U3027 ( .A1(n2351), .A2(n2349), .ZN(n4595) );
  NAND2_X1 U3028 ( .A1(n4013), .A2(n2350), .ZN(n2349) );
  INV_X1 U3029 ( .A(n2354), .ZN(n4587) );
  NAND3_X1 U3030 ( .A1(n2371), .A2(IR_REG_2__SCAN_IN), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n2370) );
  NAND2_X1 U3031 ( .A1(n2372), .A2(n2373), .ZN(n4054) );
  NAND2_X1 U3032 ( .A1(n4619), .A2(n2376), .ZN(n2372) );
  NOR2_X1 U3033 ( .A1(n4619), .A2(n4618), .ZN(n4620) );
  NAND2_X1 U3034 ( .A1(n2380), .A2(n2239), .ZN(n3190) );
  NAND2_X1 U3035 ( .A1(n2978), .A2(n2240), .ZN(n2381) );
  INV_X1 U3036 ( .A(n2391), .ZN(n3783) );
  NAND3_X1 U3037 ( .A1(n3365), .A2(n2399), .A3(n2398), .ZN(n2395) );
  NAND2_X1 U3038 ( .A1(n3289), .A2(n2393), .ZN(n2396) );
  NAND2_X1 U3039 ( .A1(n2396), .A2(n2394), .ZN(n3390) );
  NAND2_X1 U3040 ( .A1(n2404), .A2(n2402), .ZN(n3451) );
  NAND2_X1 U3041 ( .A1(n2518), .A2(n2454), .ZN(n2548) );
  NAND2_X1 U3042 ( .A1(n3757), .A2(n2412), .ZN(n2410) );
  NAND3_X1 U3043 ( .A1(n2414), .A2(n2417), .A3(n2416), .ZN(n2413) );
  NOR2_X1 U3044 ( .A1(n3746), .A2(n2435), .ZN(n3672) );
  NAND2_X1 U3045 ( .A1(n2420), .A2(n2421), .ZN(n3027) );
  NAND2_X1 U3046 ( .A1(n3746), .A2(n2429), .ZN(n2420) );
  INV_X1 U3047 ( .A(n3019), .ZN(n2433) );
  OR2_X1 U3048 ( .A1(n3673), .A2(n3674), .ZN(n2435) );
  NAND2_X1 U3049 ( .A1(n3462), .A2(n2447), .ZN(n2446) );
  NAND2_X1 U3050 ( .A1(n2436), .A2(n2440), .ZN(n2961) );
  NAND2_X1 U3051 ( .A1(n3462), .A2(n2437), .ZN(n2436) );
  XNOR2_X1 U3052 ( .A(n3078), .B(n3832), .ZN(n3659) );
  OR2_X1 U3053 ( .A1(n2823), .A2(n3261), .ZN(n2824) );
  NAND2_X1 U3054 ( .A1(n2473), .A2(IR_REG_31__SCAN_IN), .ZN(n2474) );
  AOI22_X1 U3055 ( .A1(n3573), .A2(n2661), .B1(n4498), .B2(n3580), .ZN(n4279)
         );
  OR2_X1 U3056 ( .A1(n3075), .A2(n3052), .ZN(n3077) );
  INV_X1 U3057 ( .A(n2540), .ZN(n3322) );
  NOR2_X2 U3058 ( .A1(n3747), .A2(n3748), .ZN(n3746) );
  NOR2_X1 U3059 ( .A1(n2544), .A2(n3993), .ZN(n2451) );
  AND2_X1 U3060 ( .A1(n3054), .A2(n4508), .ZN(n2452) );
  OR2_X1 U3061 ( .A1(n3073), .A2(n3072), .ZN(n2453) );
  AND2_X1 U3062 ( .A1(n2463), .A2(n2536), .ZN(n2454) );
  AND2_X1 U3063 ( .A1(n4502), .A2(n4365), .ZN(n2455) );
  AND2_X1 U3064 ( .A1(n3969), .A2(n3595), .ZN(n2456) );
  INV_X1 U3065 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2638) );
  INV_X1 U3066 ( .A(n4478), .ZN(n3102) );
  INV_X1 U3067 ( .A(n4493), .ZN(n3143) );
  INV_X1 U3068 ( .A(n4414), .ZN(n3094) );
  AND2_X1 U3069 ( .A1(n3004), .A2(n3737), .ZN(n2457) );
  AND2_X1 U3070 ( .A1(n3751), .A2(n4190), .ZN(n2458) );
  OR2_X1 U3071 ( .A1(n3677), .A2(n3752), .ZN(n2459) );
  INV_X1 U3072 ( .A(n2228), .ZN(n2777) );
  OR2_X1 U3073 ( .A1(n3598), .A2(n4400), .ZN(n2460) );
  INV_X1 U3074 ( .A(n3598), .ZN(n3970) );
  AND4_X1 U3075 ( .A1(n2631), .A2(n2630), .A3(n2629), .A4(n2628), .ZN(n3598)
         );
  NAND2_X1 U3076 ( .A1(n3301), .A2(n2553), .ZN(n2461) );
  INV_X1 U3077 ( .A(n3976), .ZN(n2563) );
  NAND2_X1 U3078 ( .A1(n3360), .A2(n2878), .ZN(n2879) );
  NOR2_X1 U3079 ( .A1(n4001), .A2(n4000), .ZN(n4002) );
  INV_X1 U3080 ( .A(n4200), .ZN(n2705) );
  INV_X1 U3081 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4847) );
  INV_X1 U3082 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3179) );
  INV_X1 U3083 ( .A(n4036), .ZN(n4037) );
  NAND2_X1 U3084 ( .A1(n4408), .A2(n3516), .ZN(n2624) );
  NAND2_X1 U3085 ( .A1(n2563), .A2(n2278), .ZN(n2564) );
  INV_X1 U3086 ( .A(IR_REG_26__SCAN_IN), .ZN(n2471) );
  OR2_X1 U3087 ( .A1(n2664), .A2(n2663), .ZN(n2677) );
  INV_X1 U3088 ( .A(n4484), .ZN(n2477) );
  NAND2_X1 U3089 ( .A1(n2697), .A2(REG3_REG_20__SCAN_IN), .ZN(n2708) );
  NAND2_X1 U3090 ( .A1(n2625), .A2(REG1_REG_1__SCAN_IN), .ZN(n2504) );
  NOR2_X1 U3091 ( .A1(n2227), .A2(n4805), .ZN(n3653) );
  AND2_X1 U3092 ( .A1(n4324), .A2(n4154), .ZN(n2725) );
  AND2_X1 U3093 ( .A1(n4195), .A2(n2846), .ZN(n4147) );
  AND2_X1 U3094 ( .A1(n2613), .A2(REG3_REG_11__SCAN_IN), .ZN(n2626) );
  INV_X1 U3095 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4848) );
  NAND2_X1 U3096 ( .A1(n3975), .A2(n3438), .ZN(n3474) );
  INV_X1 U3097 ( .A(n3653), .ZN(n3091) );
  INV_X1 U3098 ( .A(n4400), .ZN(n3617) );
  INV_X1 U3099 ( .A(n3375), .ZN(n3845) );
  INV_X1 U3100 ( .A(n4402), .ZN(n4388) );
  AND2_X1 U3101 ( .A1(n4487), .A2(n3880), .ZN(n3134) );
  NOR2_X1 U3102 ( .A1(n2610), .A2(IR_REG_9__SCAN_IN), .ZN(n2621) );
  NOR2_X1 U3103 ( .A1(n2652), .A2(n2651), .ZN(n2653) );
  NAND2_X1 U3104 ( .A1(n2727), .A2(REG3_REG_24__SCAN_IN), .ZN(n2745) );
  AND2_X1 U3105 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2541) );
  INV_X1 U3106 ( .A(n4495), .ZN(n3226) );
  NAND2_X1 U3107 ( .A1(n3158), .A2(n4492), .ZN(n3159) );
  NAND2_X1 U3108 ( .A1(n4614), .A2(n4018), .ZN(n4626) );
  INV_X1 U3109 ( .A(n4407), .ZN(n4323) );
  INV_X1 U3110 ( .A(n4136), .ZN(n4327) );
  AND2_X1 U3111 ( .A1(n3848), .A2(n4148), .ZN(n4184) );
  AND2_X1 U3112 ( .A1(n3901), .A2(n3899), .ZN(n3842) );
  INV_X1 U3113 ( .A(n4386), .ZN(n4401) );
  INV_X1 U3114 ( .A(n3752), .ZN(n4174) );
  AND2_X1 U3115 ( .A1(n3193), .A2(n3058), .ZN(n3087) );
  OR2_X1 U3116 ( .A1(n3193), .A2(n3137), .ZN(n3148) );
  AND2_X1 U3117 ( .A1(n2721), .A2(REG3_REG_23__SCAN_IN), .ZN(n2727) );
  NOR2_X1 U3118 ( .A1(n3635), .A2(n3037), .ZN(n3075) );
  INV_X1 U3119 ( .A(n3777), .ZN(n4503) );
  AND2_X1 U3120 ( .A1(n2746), .A2(n2753), .ZN(n4099) );
  AND4_X1 U3121 ( .A1(n2481), .A2(n2480), .A3(n2479), .A4(n2478), .ZN(n4369)
         );
  AND2_X1 U3122 ( .A1(n2569), .A2(n2568), .ZN(n2570) );
  AOI22_X1 U3123 ( .A1(n3269), .A2(REG2_REG_4__SCAN_IN), .B1(n4492), .B2(n3145), .ZN(n3172) );
  AND2_X1 U3124 ( .A1(n3149), .A2(n3148), .ZN(n4520) );
  AND2_X1 U3125 ( .A1(n4520), .A2(n3160), .ZN(n4631) );
  INV_X1 U3126 ( .A(n3529), .ZN(n4658) );
  NAND2_X1 U3127 ( .A1(n2811), .A2(n2810), .ZN(n3089) );
  NAND2_X1 U3128 ( .A1(n2777), .A2(DATAI_23_), .ZN(n4159) );
  AND2_X1 U3129 ( .A1(n4642), .A2(n3543), .ZN(n3546) );
  AND2_X1 U3130 ( .A1(n3119), .A2(n4675), .ZN(n3193) );
  AND2_X1 U3131 ( .A1(n3138), .A2(n3148), .ZN(n4629) );
  AND2_X1 U3132 ( .A1(n3064), .A2(n3063), .ZN(n4513) );
  INV_X1 U3133 ( .A(n4508), .ZN(n3781) );
  INV_X1 U3134 ( .A(n4309), .ZN(n3966) );
  OAI211_X1 U3135 ( .C1(n4161), .C2(n2542), .A(n2724), .B(n2723), .ZN(n4324)
         );
  INV_X1 U3136 ( .A(n4498), .ZN(n4389) );
  NAND2_X1 U3137 ( .A1(n4520), .A2(n4495), .ZN(n4635) );
  AND2_X1 U3138 ( .A1(n3512), .A2(n3514), .ZN(n4706) );
  AND2_X2 U3139 ( .A1(n2814), .A2(n4643), .ZN(n4663) );
  NAND2_X1 U3140 ( .A1(n4722), .A2(n4710), .ZN(n4414) );
  OR2_X1 U3141 ( .A1(n3115), .A2(n4478), .ZN(n3116) );
  NAND2_X1 U3142 ( .A1(n4713), .A2(n4710), .ZN(n4478) );
  OR2_X1 U3143 ( .A1(n3099), .A2(n3098), .ZN(n4711) );
  INV_X1 U3144 ( .A(n4049), .ZN(n4677) );
  INV_X1 U3145 ( .A(n4025), .ZN(n4681) );
  INV_X1 U3146 ( .A(n3979), .ZN(U4043) );
  XNOR2_X2 U3147 ( .A(n2472), .B(IR_REG_30__SCAN_IN), .ZN(n2499) );
  NAND2_X1 U31480 ( .A1(n2625), .A2(REG1_REG_16__SCAN_IN), .ZN(n2481) );
  NAND2_X1 U31490 ( .A1(n2735), .A2(REG0_REG_16__SCAN_IN), .ZN(n2480) );
  NAND2_X1 U3150 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2475) );
  NAND2_X1 U3151 ( .A1(n2653), .A2(REG3_REG_16__SCAN_IN), .ZN(n2664) );
  OR2_X1 U3152 ( .A1(n2653), .A2(REG3_REG_16__SCAN_IN), .ZN(n2476) );
  NAND2_X1 U3153 ( .A1(n2664), .A2(n2476), .ZN(n4512) );
  OR2_X1 U3154 ( .A1(n2542), .A2(n4512), .ZN(n2479) );
  INV_X1 U3155 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4283) );
  OR2_X1 U3156 ( .A1(n2544), .A2(n4283), .ZN(n2478) );
  NAND2_X1 U3158 ( .A1(n2489), .A2(n2483), .ZN(n2671) );
  NAND2_X1 U3159 ( .A1(n2671), .A2(IR_REG_31__SCAN_IN), .ZN(n2660) );
  NAND2_X1 U3160 ( .A1(n2660), .A2(n2484), .ZN(n2485) );
  NAND2_X1 U3161 ( .A1(n2485), .A2(IR_REG_31__SCAN_IN), .ZN(n2486) );
  XNOR2_X1 U3162 ( .A(n2486), .B(IR_REG_16__SCAN_IN), .ZN(n4045) );
  MUX2_X2 U3163 ( .A(n2488), .B(n2487), .S(IR_REG_27__SCAN_IN), .Z(n2551) );
  MUX2_X1 U3164 ( .A(DATAI_16_), .B(n4045), .S(n2227), .Z(n2662) );
  NOR2_X1 U3165 ( .A1(n2489), .A2(n2815), .ZN(n2490) );
  MUX2_X1 U3166 ( .A(n2815), .B(n2490), .S(IR_REG_14__SCAN_IN), .Z(n2491) );
  INV_X1 U3167 ( .A(n2491), .ZN(n2492) );
  AND2_X1 U3168 ( .A1(n2492), .A2(n2671), .ZN(n4041) );
  MUX2_X1 U3169 ( .A(DATAI_14_), .B(n4041), .S(n2227), .Z(n4387) );
  NAND2_X1 U3170 ( .A1(n2735), .A2(REG0_REG_14__SCAN_IN), .ZN(n2497) );
  NAND2_X1 U3171 ( .A1(n2625), .A2(REG1_REG_14__SCAN_IN), .ZN(n2496) );
  NAND2_X1 U3172 ( .A1(n2641), .A2(n4847), .ZN(n2493) );
  NAND2_X1 U3173 ( .A1(n2652), .A2(n2493), .ZN(n3668) );
  OR2_X1 U3174 ( .A1(n2542), .A2(n3668), .ZN(n2495) );
  INV_X1 U3175 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3563) );
  OR2_X1 U3176 ( .A1(n2544), .A2(n3563), .ZN(n2494) );
  NAND2_X1 U3177 ( .A1(n2513), .A2(REG0_REG_1__SCAN_IN), .ZN(n2503) );
  INV_X1 U3178 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3139) );
  OR2_X1 U3179 ( .A1(n3139), .A2(n4484), .ZN(n2501) );
  INV_X1 U3180 ( .A(n2499), .ZN(n2500) );
  NAND2_X1 U3181 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2505)
         );
  INV_X2 U3182 ( .A(n3256), .ZN(n3253) );
  NAND2_X1 U3183 ( .A1(n2510), .A2(n3253), .ZN(n3877) );
  NAND2_X1 U3184 ( .A1(n3877), .A2(n3881), .ZN(n2823) );
  INV_X1 U3185 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3211) );
  INV_X1 U3186 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3224) );
  OR2_X1 U3187 ( .A1(n2544), .A2(n3224), .ZN(n2508) );
  NAND2_X1 U3188 ( .A1(n2513), .A2(REG0_REG_0__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U3189 ( .A1(n2625), .A2(REG1_REG_0__SCAN_IN), .ZN(n2506) );
  NAND2_X1 U3190 ( .A1(n2823), .A2(n3250), .ZN(n3252) );
  NAND2_X1 U3191 ( .A1(n2510), .A2(n3256), .ZN(n2511) );
  NAND2_X1 U3192 ( .A1(n3252), .A2(n2511), .ZN(n3349) );
  INV_X1 U3193 ( .A(n3349), .ZN(n2520) );
  NAND2_X1 U3194 ( .A1(n2513), .A2(REG0_REG_2__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U3195 ( .A1(n2625), .A2(REG1_REG_2__SCAN_IN), .ZN(n2515) );
  INV_X1 U3196 ( .A(n2517), .ZN(n2518) );
  MUX2_X1 U3197 ( .A(DATAI_2_), .B(n4494), .S(n2228), .Z(n3360) );
  INV_X1 U3198 ( .A(n3360), .ZN(n3351) );
  NAND2_X1 U3199 ( .A1(n3978), .A2(n3351), .ZN(n3885) );
  NAND2_X1 U3200 ( .A1(n3312), .A2(n3351), .ZN(n2521) );
  NAND2_X1 U3201 ( .A1(n2625), .A2(REG1_REG_3__SCAN_IN), .ZN(n2525) );
  INV_X1 U3202 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2522) );
  NAND2_X1 U3203 ( .A1(n2513), .A2(REG0_REG_3__SCAN_IN), .ZN(n2523) );
  NAND3_X1 U3204 ( .A1(n2525), .A2(n2524), .A3(n2523), .ZN(n2526) );
  INV_X1 U3205 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3993) );
  NAND2_X1 U3206 ( .A1(n2517), .A2(IR_REG_31__SCAN_IN), .ZN(n2537) );
  XNOR2_X1 U3207 ( .A(n2537), .B(IR_REG_3__SCAN_IN), .ZN(n4493) );
  MUX2_X1 U3208 ( .A(DATAI_3_), .B(n4493), .S(n2227), .Z(n3311) );
  NAND2_X1 U3209 ( .A1(n2890), .A2(n3311), .ZN(n2527) );
  INV_X1 U32100 ( .A(n2890), .ZN(n3627) );
  NAND2_X1 U32110 ( .A1(n3627), .A2(n2888), .ZN(n3378) );
  INV_X1 U32120 ( .A(n2541), .ZN(n2530) );
  INV_X1 U32130 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2528) );
  NAND2_X1 U32140 ( .A1(n2522), .A2(n2528), .ZN(n2529) );
  NAND2_X1 U32150 ( .A1(n2530), .A2(n2529), .ZN(n3633) );
  OR2_X1 U32160 ( .A1(n2542), .A2(n3633), .ZN(n2535) );
  NAND2_X1 U32170 ( .A1(n2735), .A2(REG0_REG_4__SCAN_IN), .ZN(n2534) );
  INV_X1 U32180 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U32190 ( .A1(n2625), .A2(REG1_REG_4__SCAN_IN), .ZN(n2532) );
  NAND4_X1 U32200 ( .A1(n2535), .A2(n2534), .A3(n2533), .A4(n2532), .ZN(n2540)
         );
  NAND2_X1 U32210 ( .A1(n2537), .A2(n2536), .ZN(n2538) );
  NAND2_X1 U32220 ( .A1(n2538), .A2(IR_REG_31__SCAN_IN), .ZN(n2539) );
  XNOR2_X1 U32230 ( .A(n2539), .B(IR_REG_4__SCAN_IN), .ZN(n4492) );
  MUX2_X1 U32240 ( .A(DATAI_4_), .B(n4492), .S(n2227), .Z(n3374) );
  INV_X1 U32250 ( .A(n3374), .ZN(n3628) );
  NAND2_X1 U32260 ( .A1(n3322), .A2(n3374), .ZN(n3888) );
  NAND2_X1 U32270 ( .A1(n2735), .A2(REG0_REG_5__SCAN_IN), .ZN(n2547) );
  NAND2_X1 U32280 ( .A1(n2625), .A2(REG1_REG_5__SCAN_IN), .ZN(n2546) );
  OAI21_X1 U32290 ( .B1(n2541), .B2(REG3_REG_5__SCAN_IN), .A(n2555), .ZN(n3715) );
  OR2_X1 U32300 ( .A1(n2542), .A2(n3715), .ZN(n2545) );
  INV_X1 U32310 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2543) );
  INV_X1 U32320 ( .A(DATAI_5_), .ZN(n2552) );
  NAND2_X1 U32330 ( .A1(n2548), .A2(IR_REG_31__SCAN_IN), .ZN(n2550) );
  INV_X1 U32340 ( .A(IR_REG_5__SCAN_IN), .ZN(n2549) );
  XNOR2_X1 U32350 ( .A(n2550), .B(n2549), .ZN(n3174) );
  MUX2_X1 U32360 ( .A(n2552), .B(n3174), .S(n2228), .Z(n2904) );
  NAND2_X1 U32370 ( .A1(n2905), .A2(n2904), .ZN(n2554) );
  NAND2_X1 U32380 ( .A1(n2540), .A2(n3374), .ZN(n3301) );
  INV_X1 U32390 ( .A(n2904), .ZN(n3714) );
  NAND2_X1 U32400 ( .A1(n3977), .A2(n3714), .ZN(n2553) );
  AND2_X1 U32410 ( .A1(n2555), .A2(n3179), .ZN(n2556) );
  OR2_X1 U32420 ( .A1(n2556), .A2(n2566), .ZN(n3339) );
  OR2_X1 U32430 ( .A1(n2542), .A2(n3339), .ZN(n2560) );
  INV_X1 U32440 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3340) );
  OR2_X1 U32450 ( .A1(n2544), .A2(n3340), .ZN(n2559) );
  NAND2_X1 U32460 ( .A1(n2735), .A2(REG0_REG_6__SCAN_IN), .ZN(n2558) );
  NAND2_X1 U32470 ( .A1(n2625), .A2(REG1_REG_6__SCAN_IN), .ZN(n2557) );
  NOR2_X1 U32480 ( .A1(n2548), .A2(IR_REG_5__SCAN_IN), .ZN(n2574) );
  OR2_X1 U32490 ( .A1(n2574), .A2(n2815), .ZN(n2561) );
  XNOR2_X1 U32500 ( .A(n2561), .B(IR_REG_6__SCAN_IN), .ZN(n4490) );
  MUX2_X1 U32510 ( .A(DATAI_6_), .B(n4490), .S(n2227), .Z(n3336) );
  NAND2_X1 U32520 ( .A1(n3333), .A2(n2562), .ZN(n2565) );
  NAND2_X1 U32530 ( .A1(n2565), .A2(n2564), .ZN(n3424) );
  OR2_X1 U32540 ( .A1(n2566), .A2(REG3_REG_7__SCAN_IN), .ZN(n2567) );
  NAND2_X1 U32550 ( .A1(n2586), .A2(n2567), .ZN(n3446) );
  INV_X1 U32560 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4000) );
  OR2_X1 U32570 ( .A1(n2544), .A2(n4000), .ZN(n2571) );
  NAND2_X1 U32580 ( .A1(n2735), .A2(REG0_REG_7__SCAN_IN), .ZN(n2569) );
  NAND2_X1 U32590 ( .A1(n2625), .A2(REG1_REG_7__SCAN_IN), .ZN(n2568) );
  NAND2_X1 U32600 ( .A1(n2574), .A2(n2573), .ZN(n2593) );
  NAND2_X1 U32610 ( .A1(n2593), .A2(IR_REG_31__SCAN_IN), .ZN(n2580) );
  XNOR2_X1 U32620 ( .A(n2580), .B(IR_REG_7__SCAN_IN), .ZN(n4489) );
  MUX2_X1 U32630 ( .A(DATAI_7_), .B(n4489), .S(n2228), .Z(n3438) );
  NAND2_X1 U32640 ( .A1(n3478), .A2(n3438), .ZN(n2830) );
  INV_X1 U32650 ( .A(n3438), .ZN(n3439) );
  NAND2_X1 U32660 ( .A1(n3975), .A2(n3439), .ZN(n3900) );
  NAND2_X1 U32670 ( .A1(n2735), .A2(REG0_REG_8__SCAN_IN), .ZN(n2578) );
  NAND2_X1 U32680 ( .A1(n2625), .A2(REG1_REG_8__SCAN_IN), .ZN(n2577) );
  INV_X1 U32690 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2585) );
  XNOR2_X1 U32700 ( .A(n2586), .B(n2585), .ZN(n4644) );
  OR2_X1 U32710 ( .A1(n2542), .A2(n4644), .ZN(n2576) );
  INV_X1 U32720 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4645) );
  OR2_X1 U32730 ( .A1(n2544), .A2(n4645), .ZN(n2575) );
  INV_X1 U32740 ( .A(DATAI_8_), .ZN(n5055) );
  NAND2_X1 U32750 ( .A1(n2580), .A2(n2579), .ZN(n2581) );
  NAND2_X1 U32760 ( .A1(n2581), .A2(IR_REG_31__SCAN_IN), .ZN(n2582) );
  XNOR2_X1 U32770 ( .A(n2582), .B(IR_REG_8__SCAN_IN), .ZN(n4031) );
  INV_X1 U32780 ( .A(n4031), .ZN(n4685) );
  MUX2_X1 U32790 ( .A(n5055), .B(n4685), .S(n2227), .Z(n3477) );
  AND2_X1 U32800 ( .A1(n3493), .A2(n3477), .ZN(n2596) );
  INV_X1 U32810 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2584) );
  OAI21_X1 U32820 ( .B1(n2586), .B2(n2585), .A(n2584), .ZN(n2587) );
  NAND2_X1 U32830 ( .A1(n2587), .A2(n2603), .ZN(n3431) );
  OR2_X1 U32840 ( .A1(n2542), .A2(n3431), .ZN(n2592) );
  INV_X1 U32850 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2588) );
  OR2_X1 U32860 ( .A1(n2544), .A2(n2588), .ZN(n2591) );
  NAND2_X1 U32870 ( .A1(n2625), .A2(REG1_REG_9__SCAN_IN), .ZN(n2590) );
  NAND2_X1 U32880 ( .A1(n2735), .A2(REG0_REG_9__SCAN_IN), .ZN(n2589) );
  NAND4_X1 U32890 ( .A1(n2592), .A2(n2591), .A3(n2590), .A4(n2589), .ZN(n3973)
         );
  INV_X1 U32900 ( .A(n3973), .ZN(n2833) );
  NAND2_X1 U32910 ( .A1(n2610), .A2(IR_REG_31__SCAN_IN), .ZN(n2594) );
  XNOR2_X1 U32920 ( .A(n2594), .B(IR_REG_9__SCAN_IN), .ZN(n4027) );
  MUX2_X1 U32930 ( .A(DATAI_9_), .B(n4027), .S(n2228), .Z(n3429) );
  AND2_X1 U32940 ( .A1(n2833), .A2(n3489), .ZN(n2600) );
  NOR2_X1 U32950 ( .A1(n3424), .A2(n2595), .ZN(n2602) );
  INV_X1 U32960 ( .A(n3477), .ZN(n3394) );
  NAND2_X1 U32970 ( .A1(n3974), .A2(n3394), .ZN(n2597) );
  AND2_X1 U32980 ( .A1(n2253), .A2(n3426), .ZN(n2599) );
  NOR2_X1 U32990 ( .A1(n2602), .A2(n2601), .ZN(n3534) );
  AND2_X1 U33000 ( .A1(n2603), .A2(n4848), .ZN(n2604) );
  NOR2_X1 U33010 ( .A1(n2613), .A2(n2604), .ZN(n4636) );
  INV_X1 U33020 ( .A(n4636), .ZN(n3459) );
  OR2_X1 U33030 ( .A1(n2542), .A2(n3459), .ZN(n2609) );
  INV_X1 U33040 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2605) );
  OR2_X1 U33050 ( .A1(n2544), .A2(n2605), .ZN(n2608) );
  NAND2_X1 U33060 ( .A1(n2625), .A2(REG1_REG_10__SCAN_IN), .ZN(n2607) );
  NAND2_X1 U33070 ( .A1(n2735), .A2(REG0_REG_10__SCAN_IN), .ZN(n2606) );
  NAND4_X1 U33080 ( .A1(n2609), .A2(n2608), .A3(n2607), .A4(n2606), .ZN(n3972)
         );
  OR2_X1 U33090 ( .A1(n2621), .A2(n2815), .ZN(n2611) );
  XNOR2_X1 U33100 ( .A(n2611), .B(IR_REG_10__SCAN_IN), .ZN(n4544) );
  MUX2_X1 U33110 ( .A(DATAI_10_), .B(n4544), .S(n2228), .Z(n3456) );
  NOR2_X1 U33120 ( .A1(n3972), .A2(n3456), .ZN(n2612) );
  INV_X1 U33130 ( .A(n3972), .ZN(n2834) );
  INV_X1 U33140 ( .A(n3456), .ZN(n3536) );
  OAI22_X1 U33150 ( .A1(n3534), .A2(n2612), .B1(n2834), .B2(n3536), .ZN(n3513)
         );
  NAND2_X1 U33160 ( .A1(n2735), .A2(REG0_REG_11__SCAN_IN), .ZN(n2619) );
  NAND2_X1 U33170 ( .A1(n2625), .A2(REG1_REG_11__SCAN_IN), .ZN(n2618) );
  NOR2_X1 U33180 ( .A1(n2613), .A2(REG3_REG_11__SCAN_IN), .ZN(n2614) );
  OR2_X1 U33190 ( .A1(n2626), .A2(n2614), .ZN(n3525) );
  OR2_X1 U33200 ( .A1(n2542), .A2(n3525), .ZN(n2617) );
  INV_X1 U33210 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2615) );
  OR2_X1 U33220 ( .A1(n2544), .A2(n2615), .ZN(n2616) );
  INV_X1 U33230 ( .A(IR_REG_10__SCAN_IN), .ZN(n2620) );
  NAND2_X1 U33240 ( .A1(n2621), .A2(n2620), .ZN(n2622) );
  NAND2_X1 U33250 ( .A1(n2622), .A2(IR_REG_31__SCAN_IN), .ZN(n2633) );
  XNOR2_X1 U33260 ( .A(n2633), .B(IR_REG_11__SCAN_IN), .ZN(n4026) );
  MUX2_X1 U33270 ( .A(DATAI_11_), .B(n4026), .S(n2227), .Z(n3524) );
  NAND2_X1 U33280 ( .A1(n4408), .A2(n3524), .ZN(n3589) );
  INV_X1 U33290 ( .A(n3524), .ZN(n3516) );
  NAND2_X1 U33300 ( .A1(n3971), .A2(n3516), .ZN(n3918) );
  NAND2_X1 U33310 ( .A1(n2735), .A2(REG0_REG_12__SCAN_IN), .ZN(n2631) );
  NAND2_X1 U33320 ( .A1(n2625), .A2(REG1_REG_12__SCAN_IN), .ZN(n2630) );
  OR2_X1 U33330 ( .A1(n2626), .A2(REG3_REG_12__SCAN_IN), .ZN(n2627) );
  NAND2_X1 U33340 ( .A1(n2639), .A2(n2627), .ZN(n3613) );
  OR2_X1 U33350 ( .A1(n2542), .A2(n3613), .ZN(n2629) );
  INV_X1 U33360 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3614) );
  OR2_X1 U33370 ( .A1(n2544), .A2(n3614), .ZN(n2628) );
  INV_X1 U33380 ( .A(DATAI_12_), .ZN(n4861) );
  INV_X1 U33390 ( .A(IR_REG_11__SCAN_IN), .ZN(n2632) );
  NAND2_X1 U33400 ( .A1(n2633), .A2(n2632), .ZN(n2634) );
  NAND2_X1 U33410 ( .A1(n2634), .A2(IR_REG_31__SCAN_IN), .ZN(n2635) );
  XNOR2_X1 U33420 ( .A(n2635), .B(IR_REG_12__SCAN_IN), .ZN(n4036) );
  MUX2_X1 U33430 ( .A(n4861), .B(n4037), .S(n2228), .Z(n4400) );
  NAND2_X1 U33440 ( .A1(n2637), .A2(n2636), .ZN(n3588) );
  NAND2_X1 U33450 ( .A1(n2625), .A2(REG1_REG_13__SCAN_IN), .ZN(n2645) );
  NAND2_X1 U33460 ( .A1(n2735), .A2(REG0_REG_13__SCAN_IN), .ZN(n2644) );
  NAND2_X1 U33470 ( .A1(n2639), .A2(n2638), .ZN(n2640) );
  NAND2_X1 U33480 ( .A1(n2641), .A2(n2640), .ZN(n3602) );
  OR2_X1 U33490 ( .A1(n2542), .A2(n3602), .ZN(n2643) );
  INV_X1 U33500 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3603) );
  OR2_X1 U33510 ( .A1(n2544), .A2(n3603), .ZN(n2642) );
  INV_X1 U33520 ( .A(DATAI_13_), .ZN(n2648) );
  OR2_X1 U3353 ( .A1(n2646), .A2(n2815), .ZN(n2647) );
  XNOR2_X1 U33540 ( .A(n2647), .B(IR_REG_13__SCAN_IN), .ZN(n4025) );
  MUX2_X1 U3355 ( .A(n2648), .B(n4681), .S(n2228), .Z(n3599) );
  INV_X1 U3356 ( .A(n3599), .ZN(n3595) );
  NAND2_X1 U3357 ( .A1(n4382), .A2(n4387), .ZN(n3796) );
  INV_X1 U3358 ( .A(n4387), .ZN(n3562) );
  NAND2_X1 U3359 ( .A1(n3968), .A2(n3562), .ZN(n3797) );
  NAND2_X1 U3360 ( .A1(n3796), .A2(n3797), .ZN(n3868) );
  NAND2_X1 U3361 ( .A1(n2735), .A2(REG0_REG_15__SCAN_IN), .ZN(n2659) );
  NAND2_X1 U3362 ( .A1(n2625), .A2(REG1_REG_15__SCAN_IN), .ZN(n2658) );
  AND2_X1 U3363 ( .A1(n2652), .A2(n2651), .ZN(n2654) );
  OR2_X1 U3364 ( .A1(n2654), .A2(n2653), .ZN(n3789) );
  OR2_X1 U3365 ( .A1(n2542), .A2(n3789), .ZN(n2657) );
  INV_X1 U3366 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2655) );
  OR2_X1 U3367 ( .A1(n2544), .A2(n2655), .ZN(n2656) );
  XNOR2_X1 U3368 ( .A(n2660), .B(IR_REG_15__SCAN_IN), .ZN(n4023) );
  MUX2_X1 U3369 ( .A(DATAI_15_), .B(n4023), .S(n2228), .Z(n4378) );
  NAND2_X1 U3370 ( .A1(n4389), .A2(n4378), .ZN(n2661) );
  NAND2_X1 U3371 ( .A1(n4369), .A2(n2662), .ZN(n3928) );
  NAND2_X1 U3372 ( .A1(n4379), .A2(n4499), .ZN(n3801) );
  NAND2_X1 U3373 ( .A1(n3928), .A2(n3801), .ZN(n4284) );
  NAND2_X1 U3374 ( .A1(n4279), .A2(n4284), .ZN(n4278) );
  OAI21_X1 U3375 ( .B1(n4369), .B2(n4499), .A(n4278), .ZN(n4263) );
  NAND2_X1 U3376 ( .A1(n2625), .A2(REG1_REG_17__SCAN_IN), .ZN(n2670) );
  NAND2_X1 U3377 ( .A1(n2735), .A2(REG0_REG_17__SCAN_IN), .ZN(n2669) );
  INV_X1 U3378 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2663) );
  NAND2_X1 U3379 ( .A1(n2664), .A2(n2663), .ZN(n2665) );
  NAND2_X1 U3380 ( .A1(n2677), .A2(n2665), .ZN(n4268) );
  OR2_X1 U3381 ( .A1(n2542), .A2(n4268), .ZN(n2668) );
  INV_X1 U3382 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2666) );
  OR2_X1 U3383 ( .A1(n2544), .A2(n2666), .ZN(n2667) );
  INV_X1 U3384 ( .A(DATAI_17_), .ZN(n2675) );
  NAND2_X1 U3385 ( .A1(n2683), .A2(IR_REG_31__SCAN_IN), .ZN(n2674) );
  XNOR2_X1 U3386 ( .A(n2674), .B(IR_REG_17__SCAN_IN), .ZN(n4049) );
  MUX2_X1 U3387 ( .A(n2675), .B(n4677), .S(n2227), .Z(n4273) );
  NAND2_X1 U3388 ( .A1(n4286), .A2(n4273), .ZN(n2676) );
  INV_X1 U3389 ( .A(n4273), .ZN(n4365) );
  AOI21_X1 U3390 ( .B1(n4263), .B2(n2676), .A(n2455), .ZN(n4242) );
  NAND2_X1 U3391 ( .A1(n2735), .A2(REG0_REG_18__SCAN_IN), .ZN(n2682) );
  NAND2_X1 U3392 ( .A1(n2625), .A2(REG1_REG_18__SCAN_IN), .ZN(n2681) );
  AND2_X1 U3393 ( .A1(n2677), .A2(n4623), .ZN(n2678) );
  OR2_X1 U3394 ( .A1(n2678), .A2(n2688), .ZN(n4254) );
  OR2_X1 U3395 ( .A1(n2542), .A2(n4254), .ZN(n2680) );
  INV_X1 U3396 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4255) );
  OR2_X1 U3397 ( .A1(n2544), .A2(n4255), .ZN(n2679) );
  NAND2_X1 U3398 ( .A1(n2685), .A2(n2684), .ZN(n2694) );
  NAND2_X1 U3399 ( .A1(n2694), .A2(IR_REG_31__SCAN_IN), .ZN(n2686) );
  XNOR2_X1 U3400 ( .A(n2686), .B(IR_REG_18__SCAN_IN), .ZN(n4021) );
  MUX2_X1 U3401 ( .A(DATAI_18_), .B(n4021), .S(n2228), .Z(n4248) );
  NAND2_X1 U3402 ( .A1(n4228), .A2(n4248), .ZN(n4218) );
  INV_X1 U3403 ( .A(n4248), .ZN(n4245) );
  NAND2_X1 U3404 ( .A1(n4366), .A2(n4245), .ZN(n4219) );
  NAND2_X1 U3405 ( .A1(n4218), .A2(n4219), .ZN(n4241) );
  NOR2_X1 U3406 ( .A1(n2688), .A2(REG3_REG_19__SCAN_IN), .ZN(n2689) );
  OR2_X1 U3407 ( .A1(n2697), .A2(n2689), .ZN(n4234) );
  OR2_X1 U3408 ( .A1(n4234), .A2(n2542), .ZN(n2693) );
  INV_X1 U3409 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4235) );
  OR2_X1 U3410 ( .A1(n2544), .A2(n4235), .ZN(n2692) );
  NAND2_X1 U3411 ( .A1(n2625), .A2(REG1_REG_19__SCAN_IN), .ZN(n2691) );
  NAND2_X1 U3412 ( .A1(n2735), .A2(REG0_REG_19__SCAN_IN), .ZN(n2690) );
  INV_X1 U3413 ( .A(n2694), .ZN(n2695) );
  NAND2_X1 U3414 ( .A1(n2695), .A2(n5006), .ZN(n2696) );
  XNOR2_X2 U3415 ( .A(n2780), .B(n2779), .ZN(n4057) );
  MUX2_X1 U3416 ( .A(DATAI_19_), .B(n4253), .S(n2227), .Z(n4224) );
  NOR2_X1 U3417 ( .A1(n4249), .A2(n4224), .ZN(n4199) );
  OR2_X1 U3418 ( .A1(n2697), .A2(REG3_REG_20__SCAN_IN), .ZN(n2698) );
  AND2_X1 U3419 ( .A1(n2708), .A2(n2698), .ZN(n4207) );
  NAND2_X1 U3420 ( .A1(n2502), .A2(n4207), .ZN(n2703) );
  INV_X1 U3421 ( .A(REG2_REG_20__SCAN_IN), .ZN(n2699) );
  OR2_X1 U3422 ( .A1(n2544), .A2(n2699), .ZN(n2702) );
  NAND2_X1 U3423 ( .A1(n2735), .A2(REG0_REG_20__SCAN_IN), .ZN(n2701) );
  NAND2_X1 U3424 ( .A1(n2625), .A2(REG1_REG_20__SCAN_IN), .ZN(n2700) );
  NAND4_X1 U3425 ( .A1(n2703), .A2(n2702), .A3(n2701), .A4(n2700), .ZN(n4225)
         );
  INV_X1 U3426 ( .A(DATAI_20_), .ZN(n2704) );
  NAND2_X1 U3427 ( .A1(n4225), .A2(n4350), .ZN(n3839) );
  NAND2_X1 U3428 ( .A1(n4249), .A2(n4224), .ZN(n4200) );
  INV_X1 U3429 ( .A(n4225), .ZN(n4345) );
  NAND2_X1 U3430 ( .A1(n4345), .A2(n4205), .ZN(n3840) );
  INV_X1 U3431 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3692) );
  NAND2_X1 U3432 ( .A1(n2708), .A2(n3692), .ZN(n2709) );
  NAND2_X1 U3433 ( .A1(n2716), .A2(n2709), .ZN(n4186) );
  NAND2_X1 U3434 ( .A1(n2735), .A2(REG0_REG_21__SCAN_IN), .ZN(n2711) );
  NAND2_X1 U3435 ( .A1(n2625), .A2(REG1_REG_21__SCAN_IN), .ZN(n2710) );
  AND2_X1 U3436 ( .A1(n2711), .A2(n2710), .ZN(n2714) );
  INV_X1 U3437 ( .A(REG2_REG_21__SCAN_IN), .ZN(n2712) );
  OR2_X1 U3438 ( .A1(n2544), .A2(n2712), .ZN(n2713) );
  OAI211_X1 U3439 ( .C1(n4186), .C2(n2542), .A(n2714), .B(n2713), .ZN(n4351)
         );
  INV_X1 U3440 ( .A(n4190), .ZN(n4341) );
  NAND2_X1 U3441 ( .A1(n4351), .A2(n4341), .ZN(n2715) );
  INV_X1 U3442 ( .A(n4351), .ZN(n3751) );
  AOI21_X1 U3443 ( .B1(n4183), .B2(n2715), .A(n2458), .ZN(n4167) );
  INV_X1 U3444 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3750) );
  AND2_X1 U3445 ( .A1(n2716), .A2(n3750), .ZN(n2717) );
  OR2_X1 U3446 ( .A1(n2717), .A2(n2721), .ZN(n3749) );
  AOI22_X1 U3447 ( .A1(n2735), .A2(REG0_REG_22__SCAN_IN), .B1(n2625), .B2(
        REG1_REG_22__SCAN_IN), .ZN(n2720) );
  INV_X1 U3448 ( .A(REG2_REG_22__SCAN_IN), .ZN(n2718) );
  OR2_X1 U3449 ( .A1(n2544), .A2(n2718), .ZN(n2719) );
  OAI211_X1 U3450 ( .C1(n3749), .C2(n2542), .A(n2720), .B(n2719), .ZN(n4342)
         );
  OR2_X1 U3451 ( .A1(n4342), .A2(n3752), .ZN(n4150) );
  NAND2_X1 U3452 ( .A1(n4342), .A2(n3752), .ZN(n2850) );
  NAND2_X1 U3453 ( .A1(n4150), .A2(n2850), .ZN(n4168) );
  NAND2_X1 U3454 ( .A1(n4167), .A2(n4168), .ZN(n4166) );
  NAND2_X1 U3455 ( .A1(n4166), .A2(n2459), .ZN(n4141) );
  NOR2_X1 U3456 ( .A1(n2721), .A2(REG3_REG_23__SCAN_IN), .ZN(n2722) );
  OR2_X1 U3457 ( .A1(n2727), .A2(n2722), .ZN(n4161) );
  AOI22_X1 U34580 ( .A1(n2735), .A2(REG0_REG_23__SCAN_IN), .B1(n2625), .B2(
        REG1_REG_23__SCAN_IN), .ZN(n2724) );
  INV_X1 U34590 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4160) );
  INV_X1 U3460 ( .A(n4324), .ZN(n4173) );
  NAND2_X1 U3461 ( .A1(n4173), .A2(n4159), .ZN(n2726) );
  OR2_X1 U3462 ( .A1(n2727), .A2(REG3_REG_24__SCAN_IN), .ZN(n2728) );
  AND2_X1 U3463 ( .A1(n2745), .A2(n2728), .ZN(n4131) );
  NAND2_X1 U3464 ( .A1(n4131), .A2(n2502), .ZN(n2733) );
  INV_X1 U3465 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4129) );
  NAND2_X1 U3466 ( .A1(n2735), .A2(REG0_REG_24__SCAN_IN), .ZN(n2730) );
  NAND2_X1 U34670 ( .A1(n2625), .A2(REG1_REG_24__SCAN_IN), .ZN(n2729) );
  OAI211_X1 U3468 ( .C1(n4129), .C2(n2544), .A(n2730), .B(n2729), .ZN(n2731)
         );
  INV_X1 U34690 ( .A(n2731), .ZN(n2732) );
  NAND2_X1 U3470 ( .A1(n2777), .A2(DATAI_24_), .ZN(n4134) );
  NAND2_X1 U34710 ( .A1(n4108), .A2(n4322), .ZN(n2734) );
  XNOR2_X1 U3472 ( .A(n2745), .B(REG3_REG_25__SCAN_IN), .ZN(n4114) );
  NAND2_X1 U34730 ( .A1(n4114), .A2(n2502), .ZN(n2741) );
  INV_X1 U3474 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2738) );
  NAND2_X1 U34750 ( .A1(n2625), .A2(REG1_REG_25__SCAN_IN), .ZN(n2737) );
  NAND2_X1 U3476 ( .A1(n2735), .A2(REG0_REG_25__SCAN_IN), .ZN(n2736) );
  OAI211_X1 U34770 ( .C1(n2738), .C2(n2544), .A(n2737), .B(n2736), .ZN(n2739)
         );
  INV_X1 U3478 ( .A(n2739), .ZN(n2740) );
  NAND2_X1 U34790 ( .A1(n2777), .A2(DATAI_25_), .ZN(n4113) );
  NAND2_X1 U3480 ( .A1(n4327), .A2(n4113), .ZN(n2743) );
  NOR2_X1 U34810 ( .A1(n4327), .A2(n4113), .ZN(n2742) );
  INV_X1 U3482 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3703) );
  INV_X1 U34830 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2744) );
  OAI21_X1 U3484 ( .B1(n2745), .B2(n3703), .A(n2744), .ZN(n2746) );
  NAND2_X1 U34850 ( .A1(n4099), .A2(n2502), .ZN(n2752) );
  INV_X1 U3486 ( .A(REG2_REG_26__SCAN_IN), .ZN(n2749) );
  NAND2_X1 U34870 ( .A1(n2735), .A2(REG0_REG_26__SCAN_IN), .ZN(n2748) );
  NAND2_X1 U3488 ( .A1(n2625), .A2(REG1_REG_26__SCAN_IN), .ZN(n2747) );
  OAI211_X1 U34890 ( .C1(n2749), .C2(n2544), .A(n2748), .B(n2747), .ZN(n2750)
         );
  INV_X1 U3490 ( .A(n2750), .ZN(n2751) );
  INV_X1 U34910 ( .A(n4306), .ZN(n4111) );
  NAND2_X1 U3492 ( .A1(n2777), .A2(DATAI_26_), .ZN(n4097) );
  INV_X1 U34930 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4981) );
  INV_X1 U3494 ( .A(n2762), .ZN(n2764) );
  NAND2_X1 U34950 ( .A1(n2753), .A2(n4981), .ZN(n2754) );
  NAND2_X1 U3496 ( .A1(n2764), .A2(n2754), .ZN(n4077) );
  OR2_X1 U34970 ( .A1(n4077), .A2(n2542), .ZN(n2759) );
  INV_X1 U3498 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4076) );
  NAND2_X1 U34990 ( .A1(n2625), .A2(REG1_REG_27__SCAN_IN), .ZN(n2756) );
  NAND2_X1 U3500 ( .A1(n2735), .A2(REG0_REG_27__SCAN_IN), .ZN(n2755) );
  OAI211_X1 U35010 ( .C1(n4076), .C2(n2544), .A(n2756), .B(n2755), .ZN(n2757)
         );
  INV_X1 U3502 ( .A(n2757), .ZN(n2758) );
  INV_X1 U35030 ( .A(DATAI_27_), .ZN(n2760) );
  NOR2_X1 U3504 ( .A1(n3967), .A2(n4305), .ZN(n2761) );
  INV_X1 U35050 ( .A(n4305), .ZN(n4075) );
  NAND2_X1 U35060 ( .A1(n2762), .A2(REG3_REG_28__SCAN_IN), .ZN(n2822) );
  INV_X1 U35070 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2763) );
  NAND2_X1 U35080 ( .A1(n2764), .A2(n2763), .ZN(n2765) );
  NAND2_X1 U35090 ( .A1(n2822), .A2(n2765), .ZN(n3649) );
  OR2_X1 U35100 ( .A1(n3649), .A2(n2542), .ZN(n2770) );
  INV_X1 U35110 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3648) );
  NAND2_X1 U35120 ( .A1(n2735), .A2(REG0_REG_28__SCAN_IN), .ZN(n2767) );
  NAND2_X1 U35130 ( .A1(n2625), .A2(REG1_REG_28__SCAN_IN), .ZN(n2766) );
  OAI211_X1 U35140 ( .C1(n3648), .C2(n2544), .A(n2767), .B(n2766), .ZN(n2768)
         );
  INV_X1 U35150 ( .A(n2768), .ZN(n2769) );
  INV_X1 U35160 ( .A(DATAI_28_), .ZN(n4805) );
  NAND2_X1 U35170 ( .A1(n3966), .A2(n3091), .ZN(n2853) );
  NAND2_X1 U35180 ( .A1(n2854), .A2(n2853), .ZN(n3832) );
  OR2_X1 U35190 ( .A1(n2822), .A2(n2542), .ZN(n2776) );
  INV_X1 U35200 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3110) );
  NAND2_X1 U35210 ( .A1(n2735), .A2(REG0_REG_29__SCAN_IN), .ZN(n2773) );
  NAND2_X1 U35220 ( .A1(n2512), .A2(REG2_REG_29__SCAN_IN), .ZN(n2772) );
  OAI211_X1 U35230 ( .C1(n3110), .C2(n2498), .A(n2773), .B(n2772), .ZN(n2774)
         );
  INV_X1 U35240 ( .A(n2774), .ZN(n2775) );
  NAND2_X1 U35250 ( .A1(n2776), .A2(n2775), .ZN(n3965) );
  NAND2_X1 U35260 ( .A1(n2777), .A2(DATAI_29_), .ZN(n3816) );
  XNOR2_X1 U35270 ( .A(n3965), .B(n3816), .ZN(n3856) );
  XNOR2_X1 U35280 ( .A(n2778), .B(n3856), .ZN(n3109) );
  INV_X1 U35290 ( .A(n3109), .ZN(n2864) );
  NAND2_X1 U35300 ( .A1(n2780), .A2(n2779), .ZN(n2781) );
  NAND2_X1 U35310 ( .A1(n2781), .A2(IR_REG_31__SCAN_IN), .ZN(n2783) );
  NAND2_X1 U35320 ( .A1(n2784), .A2(IR_REG_31__SCAN_IN), .ZN(n2785) );
  NAND2_X1 U35330 ( .A1(n2245), .A2(IR_REG_31__SCAN_IN), .ZN(n2786) );
  XNOR2_X1 U35340 ( .A(n2866), .B(n4487), .ZN(n2787) );
  NAND2_X1 U35350 ( .A1(n2787), .A2(n4057), .ZN(n3517) );
  INV_X1 U35360 ( .A(n3517), .ZN(n3561) );
  NOR2_X1 U35370 ( .A1(n2866), .A2(n4057), .ZN(n3210) );
  NOR4_X1 U35380 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n2791) );
  NOR4_X1 U35390 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2790) );
  NOR4_X1 U35400 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2789) );
  NOR4_X1 U35410 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n2788) );
  NAND4_X1 U35420 ( .A1(n2791), .A2(n2790), .A3(n2789), .A4(n2788), .ZN(n2805)
         );
  NOR2_X1 U35430 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_28__SCAN_IN), .ZN(n2795)
         );
  NOR4_X1 U35440 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_23__SCAN_IN), .ZN(n2794) );
  NOR4_X1 U35450 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2793) );
  NOR4_X1 U35460 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2792) );
  NAND4_X1 U35470 ( .A1(n2795), .A2(n2794), .A3(n2793), .A4(n2792), .ZN(n2804)
         );
  NAND2_X1 U35480 ( .A1(n2255), .A2(IR_REG_31__SCAN_IN), .ZN(n2796) );
  MUX2_X1 U35490 ( .A(IR_REG_31__SCAN_IN), .B(n2796), .S(IR_REG_25__SCAN_IN), 
        .Z(n2797) );
  NAND2_X1 U35500 ( .A1(n2797), .A2(n2250), .ZN(n3131) );
  NAND2_X1 U35510 ( .A1(n3131), .A2(B_REG_SCAN_IN), .ZN(n2801) );
  OR2_X1 U35520 ( .A1(n2798), .A2(n2815), .ZN(n2807) );
  NAND2_X1 U35530 ( .A1(n2807), .A2(n2806), .ZN(n2799) );
  NAND2_X1 U35540 ( .A1(n2799), .A2(IR_REG_31__SCAN_IN), .ZN(n2800) );
  MUX2_X1 U35550 ( .A(n2801), .B(B_REG_SCAN_IN), .S(n4486), .Z(n2803) );
  NAND2_X1 U35560 ( .A1(n2250), .A2(IR_REG_31__SCAN_IN), .ZN(n2802) );
  OAI21_X1 U35570 ( .B1(n2805), .B2(n2804), .A(n3125), .ZN(n3086) );
  INV_X1 U35580 ( .A(n4485), .ZN(n3128) );
  NAND2_X1 U35590 ( .A1(n3128), .A2(n3131), .ZN(n3083) );
  AND2_X1 U35600 ( .A1(n3086), .A2(n3083), .ZN(n3045) );
  INV_X1 U35610 ( .A(n3131), .ZN(n3121) );
  XNOR2_X1 U35620 ( .A(n2807), .B(n2806), .ZN(n3135) );
  NAND2_X1 U35630 ( .A1(n2808), .A2(n4057), .ZN(n3046) );
  NAND2_X1 U35640 ( .A1(n3046), .A2(n3134), .ZN(n3058) );
  INV_X1 U35650 ( .A(D_REG_0__SCAN_IN), .ZN(n2809) );
  NAND2_X1 U35660 ( .A1(n3125), .A2(n2809), .ZN(n2811) );
  INV_X1 U35670 ( .A(n4486), .ZN(n3127) );
  NAND2_X1 U35680 ( .A1(n3128), .A2(n3127), .ZN(n2810) );
  INV_X1 U35690 ( .A(D_REG_1__SCAN_IN), .ZN(n2812) );
  NAND2_X1 U35700 ( .A1(n3125), .A2(n2812), .ZN(n3084) );
  NAND4_X1 U35710 ( .A1(n3045), .A2(n3087), .A3(n3089), .A4(n3084), .ZN(n2814)
         );
  NAND2_X1 U35720 ( .A1(n2808), .A2(n4253), .ZN(n3209) );
  OAI21_X2 U35730 ( .B1(n3561), .B2(n3210), .A(n4646), .ZN(n4295) );
  OR2_X1 U35740 ( .A1(n2241), .A2(n2815), .ZN(n2817) );
  INV_X2 U35750 ( .A(n4663), .ZN(n4646) );
  INV_X1 U35760 ( .A(n2808), .ZN(n4488) );
  INV_X1 U35770 ( .A(n4487), .ZN(n2818) );
  INV_X1 U35780 ( .A(n3880), .ZN(n3873) );
  NAND2_X1 U35790 ( .A1(n4646), .A2(n4386), .ZN(n4272) );
  INV_X1 U35800 ( .A(REG2_REG_29__SCAN_IN), .ZN(n2819) );
  OAI22_X1 U35810 ( .A1(n4272), .A2(n3816), .B1(n2819), .B2(n4646), .ZN(n2820)
         );
  AOI21_X1 U3582 ( .B1(n3966), .B2(n4267), .A(n2820), .ZN(n2863) );
  NAND2_X1 U3583 ( .A1(n3358), .A2(n2888), .ZN(n3373) );
  NOR2_X2 U3584 ( .A1(n3373), .A2(n3374), .ZN(n3372) );
  NAND2_X1 U3585 ( .A1(n3372), .A2(n2904), .ZN(n3337) );
  NOR2_X4 U3586 ( .A1(n3574), .A2(n4378), .ZN(n4282) );
  AND2_X2 U3587 ( .A1(n4072), .A2(n3091), .ZN(n3093) );
  OAI21_X1 U3588 ( .B1(n3093), .B2(n3816), .A(n4299), .ZN(n3115) );
  AND2_X1 U3589 ( .A1(n4710), .A2(n4057), .ZN(n2821) );
  OAI22_X1 U3590 ( .A1(n3115), .A2(n4233), .B1(n2822), .B2(n4643), .ZN(n2861)
         );
  INV_X1 U3591 ( .A(n3257), .ZN(n3207) );
  NAND2_X1 U3592 ( .A1(n3207), .A2(n3206), .ZN(n3261) );
  NAND2_X1 U3593 ( .A1(n3350), .A2(n3851), .ZN(n2826) );
  NAND2_X1 U3594 ( .A1(n2826), .A2(n3882), .ZN(n3280) );
  NAND2_X1 U3595 ( .A1(n3627), .A2(n3311), .ZN(n3887) );
  NAND2_X1 U3596 ( .A1(n2890), .A2(n2888), .ZN(n3884) );
  INV_X1 U3597 ( .A(n3887), .ZN(n2827) );
  NAND2_X1 U3598 ( .A1(n3376), .A2(n3888), .ZN(n2828) );
  AND2_X1 U3599 ( .A1(n3977), .A2(n2904), .ZN(n3892) );
  NAND2_X1 U3600 ( .A1(n2905), .A2(n3714), .ZN(n3909) );
  NAND2_X1 U3601 ( .A1(n3976), .A2(n2278), .ZN(n3890) );
  NAND2_X1 U3602 ( .A1(n2563), .A2(n3336), .ZN(n3894) );
  NAND2_X1 U3603 ( .A1(n2829), .A2(n3894), .ZN(n3441) );
  INV_X1 U3604 ( .A(n2830), .ZN(n3896) );
  NAND2_X1 U3605 ( .A1(n2831), .A2(n3900), .ZN(n3476) );
  NAND2_X1 U3606 ( .A1(n3493), .A2(n3394), .ZN(n3901) );
  NAND2_X1 U3607 ( .A1(n3476), .A2(n3901), .ZN(n2832) );
  NAND2_X1 U3608 ( .A1(n3974), .A2(n3477), .ZN(n3899) );
  AND2_X1 U3609 ( .A1(n3973), .A2(n3489), .ZN(n3908) );
  NAND2_X1 U3610 ( .A1(n2833), .A2(n3429), .ZN(n3902) );
  NAND2_X1 U3611 ( .A1(n3972), .A2(n3536), .ZN(n3917) );
  NAND2_X1 U3612 ( .A1(n2834), .A2(n3456), .ZN(n3912) );
  NAND2_X1 U3613 ( .A1(n2835), .A2(n3912), .ZN(n3515) );
  NAND2_X1 U3614 ( .A1(n3970), .A2(n4400), .ZN(n3608) );
  NAND2_X1 U3615 ( .A1(n3969), .A2(n3599), .ZN(n3585) );
  NAND2_X1 U3616 ( .A1(n3591), .A2(n3919), .ZN(n2837) );
  NAND2_X1 U3617 ( .A1(n3598), .A2(n3617), .ZN(n3609) );
  NAND2_X1 U3618 ( .A1(n3589), .A2(n3609), .ZN(n2836) );
  NOR2_X1 U3619 ( .A1(n3969), .A2(n3599), .ZN(n3587) );
  AOI21_X1 U3620 ( .B1(n2836), .B2(n3919), .A(n3587), .ZN(n3921) );
  NAND2_X1 U3621 ( .A1(n2837), .A2(n3921), .ZN(n3800) );
  NAND2_X1 U3622 ( .A1(n3800), .A2(n2325), .ZN(n3569) );
  NAND2_X1 U3623 ( .A1(n4498), .A2(n4378), .ZN(n3799) );
  NAND2_X1 U3624 ( .A1(n4389), .A2(n3580), .ZN(n3798) );
  NAND2_X1 U3625 ( .A1(n3799), .A2(n3798), .ZN(n3867) );
  INV_X1 U3626 ( .A(n3796), .ZN(n2838) );
  NOR2_X1 U3627 ( .A1(n3867), .A2(n2838), .ZN(n2839) );
  NAND2_X1 U3628 ( .A1(n3569), .A2(n2839), .ZN(n2840) );
  NAND2_X1 U3629 ( .A1(n2840), .A2(n3798), .ZN(n4285) );
  INV_X1 U3630 ( .A(n4284), .ZN(n2841) );
  NAND2_X1 U3631 ( .A1(n4285), .A2(n2841), .ZN(n2842) );
  NAND2_X1 U3632 ( .A1(n2842), .A2(n3801), .ZN(n4260) );
  NAND2_X1 U3633 ( .A1(n4286), .A2(n4365), .ZN(n4216) );
  NAND2_X1 U3634 ( .A1(n4218), .A2(n4216), .ZN(n2845) );
  INV_X1 U3635 ( .A(n4224), .ZN(n4231) );
  NAND2_X1 U3636 ( .A1(n4249), .A2(n4231), .ZN(n2843) );
  AND2_X1 U3637 ( .A1(n4219), .A2(n2843), .ZN(n4144) );
  NOR2_X1 U3638 ( .A1(n4249), .A2(n4231), .ZN(n2844) );
  AOI21_X1 U3639 ( .B1(n2845), .B2(n4144), .A(n2844), .ZN(n4195) );
  NAND2_X1 U3640 ( .A1(n4345), .A2(n4350), .ZN(n2846) );
  NAND2_X1 U3641 ( .A1(n4260), .A2(n4147), .ZN(n2847) );
  NAND2_X1 U3642 ( .A1(n4502), .A2(n4273), .ZN(n4142) );
  NAND2_X1 U3643 ( .A1(n4144), .A2(n4142), .ZN(n3929) );
  AND2_X1 U3644 ( .A1(n4225), .A2(n4205), .ZN(n4146) );
  AOI21_X1 U3645 ( .B1(n4147), .B2(n3929), .A(n4146), .ZN(n3803) );
  NAND2_X1 U3646 ( .A1(n2847), .A2(n3803), .ZN(n2849) );
  OR2_X1 U3647 ( .A1(n4351), .A2(n4190), .ZN(n4148) );
  NAND2_X1 U3648 ( .A1(n4150), .A2(n4148), .ZN(n3935) );
  INV_X1 U3649 ( .A(n3935), .ZN(n2848) );
  NAND2_X1 U3650 ( .A1(n4324), .A2(n4159), .ZN(n2851) );
  NAND2_X1 U3651 ( .A1(n2851), .A2(n2850), .ZN(n3938) );
  AND2_X1 U3652 ( .A1(n4351), .A2(n4190), .ZN(n3933) );
  AND2_X1 U3653 ( .A1(n4150), .A2(n3933), .ZN(n2852) );
  NOR2_X1 U3654 ( .A1(n3938), .A2(n2852), .ZN(n3807) );
  NOR2_X1 U3655 ( .A1(n4108), .A2(n4134), .ZN(n3838) );
  NOR2_X1 U3656 ( .A1(n4324), .A2(n4159), .ZN(n4121) );
  NOR2_X1 U3657 ( .A1(n3838), .A2(n4121), .ZN(n3937) );
  AND2_X1 U3658 ( .A1(n4108), .A2(n4134), .ZN(n3837) );
  NAND2_X1 U3659 ( .A1(n4136), .A2(n4113), .ZN(n3858) );
  NOR2_X1 U3660 ( .A1(n4306), .A2(n4097), .ZN(n3833) );
  NOR2_X1 U3661 ( .A1(n4136), .A2(n4113), .ZN(n3857) );
  NOR2_X1 U3662 ( .A1(n3833), .A2(n3857), .ZN(n3945) );
  NAND2_X1 U3663 ( .A1(n4306), .A2(n4097), .ZN(n3817) );
  INV_X1 U3664 ( .A(n3817), .ZN(n3834) );
  NOR2_X1 U3665 ( .A1(n4092), .A2(n4305), .ZN(n3943) );
  AOI21_X1 U3666 ( .B1(n4068), .B2(n4071), .A(n3818), .ZN(n3080) );
  INV_X1 U3667 ( .A(n2853), .ZN(n3815) );
  NAND2_X1 U3668 ( .A1(n4488), .A2(n3880), .ZN(n3955) );
  NAND2_X1 U3669 ( .A1(n4253), .A2(n4487), .ZN(n2855) );
  NAND2_X2 U3670 ( .A1(n3955), .A2(n2855), .ZN(n4289) );
  XNOR2_X1 U3671 ( .A(n2856), .B(IR_REG_27__SCAN_IN), .ZN(n4518) );
  AOI21_X1 U3672 ( .B1(B_REG_SCAN_IN), .B2(n4518), .A(n4402), .ZN(n4062) );
  INV_X1 U3673 ( .A(REG2_REG_30__SCAN_IN), .ZN(n2859) );
  NAND2_X1 U3674 ( .A1(n2625), .A2(REG1_REG_30__SCAN_IN), .ZN(n2858) );
  NAND2_X1 U3675 ( .A1(n2735), .A2(REG0_REG_30__SCAN_IN), .ZN(n2857) );
  OAI211_X1 U3676 ( .C1(n2544), .C2(n2859), .A(n2858), .B(n2857), .ZN(n3964)
         );
  INV_X1 U3677 ( .A(n3107), .ZN(n2860) );
  OAI211_X1 U3678 ( .C1(n2864), .C2(n4295), .A(n2863), .B(n2862), .ZN(U3354)
         );
  INV_X2 U3679 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3680 ( .A(n2866), .ZN(n2865) );
  INV_X1 U3681 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2867) );
  OR2_X2 U3682 ( .A1(n3040), .A2(n4710), .ZN(n2882) );
  NAND2_X1 U3683 ( .A1(n3257), .A2(n3033), .ZN(n2869) );
  INV_X1 U3684 ( .A(n3119), .ZN(n3060) );
  AOI22_X1 U3685 ( .A1(n3206), .A2(n2242), .B1(IR_REG_0__SCAN_IN), .B2(n3060), 
        .ZN(n2868) );
  NAND2_X1 U3686 ( .A1(n2869), .A2(n2868), .ZN(n3189) );
  NAND2_X1 U3687 ( .A1(n3190), .A2(n3189), .ZN(n3188) );
  INV_X1 U3688 ( .A(n3061), .ZN(n2870) );
  NAND2_X1 U3689 ( .A1(n3188), .A2(n2871), .ZN(n3198) );
  XNOR2_X1 U3690 ( .A(n2872), .B(n3030), .ZN(n2873) );
  OAI22_X1 U3691 ( .A1(n3352), .A2(n2882), .B1(n2955), .B2(n3253), .ZN(n2874)
         );
  XNOR2_X1 U3692 ( .A(n2873), .B(n2874), .ZN(n3197) );
  NAND2_X1 U3693 ( .A1(n3198), .A2(n3197), .ZN(n3199) );
  INV_X1 U3694 ( .A(n2873), .ZN(n2875) );
  NAND2_X1 U3695 ( .A1(n2875), .A2(n2874), .ZN(n2876) );
  NAND2_X1 U3696 ( .A1(n3199), .A2(n2876), .ZN(n3216) );
  INV_X1 U3697 ( .A(n3216), .ZN(n2884) );
  XNOR2_X1 U3698 ( .A(n2881), .B(n3038), .ZN(n2892) );
  OAI22_X1 U3699 ( .A1(n3312), .A2(n2882), .B1(n3351), .B2(n2955), .ZN(n2893)
         );
  XNOR2_X1 U3700 ( .A(n2892), .B(n2893), .ZN(n3215) );
  INV_X1 U3701 ( .A(n3215), .ZN(n2883) );
  NAND2_X1 U3702 ( .A1(n2884), .A2(n2883), .ZN(n3217) );
  NAND2_X1 U3703 ( .A1(n2890), .A2(n2242), .ZN(n2886) );
  NAND2_X1 U3704 ( .A1(n3311), .A2(n2878), .ZN(n2885) );
  NAND2_X1 U3705 ( .A1(n2886), .A2(n2885), .ZN(n2887) );
  INV_X1 U3706 ( .A(n2898), .ZN(n2891) );
  NOR2_X1 U3707 ( .A1(n2888), .A2(n2955), .ZN(n2889) );
  AOI21_X1 U3708 ( .B1(n2890), .B2(n3033), .A(n2889), .ZN(n2897) );
  NAND2_X1 U3709 ( .A1(n2891), .A2(n2897), .ZN(n2896) );
  INV_X1 U3710 ( .A(n2892), .ZN(n2895) );
  INV_X1 U3711 ( .A(n2893), .ZN(n2894) );
  NAND2_X1 U3712 ( .A1(n2895), .A2(n2894), .ZN(n3244) );
  AND2_X1 U3713 ( .A1(n2896), .A2(n3244), .ZN(n2901) );
  INV_X1 U3714 ( .A(n2896), .ZN(n2899) );
  XNOR2_X1 U3715 ( .A(n2898), .B(n2897), .ZN(n3243) );
  NOR2_X1 U3716 ( .A1(n2899), .A2(n3243), .ZN(n2900) );
  OAI22_X1 U3717 ( .A1(n3322), .A2(n2955), .B1(n3040), .B2(n3628), .ZN(n2902)
         );
  XNOR2_X1 U3718 ( .A(n2902), .B(n3038), .ZN(n2911) );
  OAI22_X1 U3719 ( .A1(n3322), .A2(n2882), .B1(n2955), .B2(n3628), .ZN(n2910)
         );
  XNOR2_X1 U3720 ( .A(n2911), .B(n2910), .ZN(n3625) );
  OAI22_X1 U3721 ( .A1(n2905), .A2(n2955), .B1(n2904), .B2(n3040), .ZN(n2903)
         );
  XNOR2_X1 U3722 ( .A(n2903), .B(n3030), .ZN(n2908) );
  INV_X1 U3723 ( .A(n2908), .ZN(n2906) );
  OAI22_X1 U3724 ( .A1(n2905), .A2(n2882), .B1(n2904), .B2(n2955), .ZN(n2907)
         );
  XNOR2_X1 U3725 ( .A(n2908), .B(n2907), .ZN(n3710) );
  NOR2_X1 U3726 ( .A1(n2909), .A2(n3710), .ZN(n2914) );
  NAND2_X1 U3727 ( .A1(n2911), .A2(n2910), .ZN(n3708) );
  AND2_X1 U3728 ( .A1(n3708), .A2(n2912), .ZN(n2913) );
  OR2_X1 U3729 ( .A1(n2914), .A2(n2913), .ZN(n2915) );
  NAND2_X1 U3730 ( .A1(n3976), .A2(n3033), .ZN(n2918) );
  NAND2_X1 U3731 ( .A1(n3336), .A2(n2242), .ZN(n2917) );
  NAND2_X1 U3732 ( .A1(n2918), .A2(n2917), .ZN(n3290) );
  NAND2_X1 U3733 ( .A1(n3976), .A2(n2877), .ZN(n2920) );
  NAND2_X1 U3734 ( .A1(n3336), .A2(n2878), .ZN(n2919) );
  NAND2_X1 U3735 ( .A1(n2920), .A2(n2919), .ZN(n2921) );
  XNOR2_X1 U3736 ( .A(n2921), .B(n3038), .ZN(n3291) );
  OAI22_X1 U3737 ( .A1(n3478), .A2(n2955), .B1(n3040), .B2(n3439), .ZN(n2922)
         );
  XNOR2_X1 U3738 ( .A(n2922), .B(n3030), .ZN(n2923) );
  OAI22_X1 U3739 ( .A1(n3478), .A2(n2882), .B1(n2955), .B2(n3439), .ZN(n2924)
         );
  INV_X1 U3740 ( .A(n2923), .ZN(n2925) );
  NAND2_X1 U3741 ( .A1(n2925), .A2(n2924), .ZN(n2926) );
  INV_X1 U3742 ( .A(n3390), .ZN(n2932) );
  OAI22_X1 U3743 ( .A1(n3493), .A2(n2955), .B1(n3040), .B2(n3477), .ZN(n2927)
         );
  XNOR2_X1 U3744 ( .A(n2927), .B(n3038), .ZN(n2933) );
  OAI22_X1 U3745 ( .A1(n3493), .A2(n2882), .B1(n2955), .B2(n3477), .ZN(n2934)
         );
  AND2_X1 U3746 ( .A1(n2933), .A2(n2934), .ZN(n3412) );
  NAND2_X1 U3747 ( .A1(n3973), .A2(n2242), .ZN(n2929) );
  NAND2_X1 U3748 ( .A1(n3429), .A2(n2878), .ZN(n2928) );
  NAND2_X1 U3749 ( .A1(n2929), .A2(n2928), .ZN(n2930) );
  XNOR2_X1 U3750 ( .A(n2930), .B(n3038), .ZN(n2938) );
  NOR2_X1 U3751 ( .A1(n3489), .A2(n2955), .ZN(n2931) );
  AOI21_X1 U3752 ( .B1(n3973), .B2(n3033), .A(n2931), .ZN(n2939) );
  XNOR2_X1 U3753 ( .A(n2938), .B(n2939), .ZN(n3415) );
  INV_X1 U3754 ( .A(n3415), .ZN(n2937) );
  INV_X1 U3755 ( .A(n2933), .ZN(n2936) );
  INV_X1 U3756 ( .A(n2934), .ZN(n2935) );
  NAND2_X1 U3757 ( .A1(n2936), .A2(n2935), .ZN(n3413) );
  OR2_X1 U3758 ( .A1(n2937), .A2(n3413), .ZN(n2942) );
  INV_X1 U3759 ( .A(n2938), .ZN(n2940) );
  NAND2_X1 U3760 ( .A1(n2940), .A2(n2939), .ZN(n2941) );
  AND2_X1 U3761 ( .A1(n2942), .A2(n2941), .ZN(n2943) );
  NAND2_X1 U3762 ( .A1(n3972), .A2(n2877), .ZN(n2945) );
  NAND2_X1 U3763 ( .A1(n3456), .A2(n2878), .ZN(n2944) );
  NAND2_X1 U3764 ( .A1(n2945), .A2(n2944), .ZN(n2946) );
  XNOR2_X1 U3765 ( .A(n2946), .B(n3030), .ZN(n2948) );
  NOR2_X1 U3766 ( .A1(n3536), .A2(n2955), .ZN(n2947) );
  AOI21_X1 U3767 ( .B1(n3972), .B2(n3033), .A(n2947), .ZN(n2949) );
  XNOR2_X1 U3768 ( .A(n2948), .B(n2949), .ZN(n3454) );
  INV_X1 U3769 ( .A(n2948), .ZN(n2951) );
  INV_X1 U3770 ( .A(n2949), .ZN(n2950) );
  NAND2_X1 U3771 ( .A1(n2951), .A2(n2950), .ZN(n2952) );
  NAND2_X1 U3772 ( .A1(n3451), .A2(n2952), .ZN(n3462) );
  OAI22_X1 U3773 ( .A1(n4408), .A2(n2882), .B1(n2955), .B2(n3516), .ZN(n3463)
         );
  OAI22_X1 U3774 ( .A1(n4408), .A2(n2955), .B1(n3040), .B2(n3516), .ZN(n2953)
         );
  XNOR2_X1 U3775 ( .A(n2953), .B(n3038), .ZN(n3464) );
  OAI22_X1 U3776 ( .A1(n3598), .A2(n2955), .B1(n3040), .B2(n4400), .ZN(n2954)
         );
  XNOR2_X1 U3777 ( .A(n2954), .B(n3038), .ZN(n2956) );
  OAI22_X1 U3778 ( .A1(n3598), .A2(n2882), .B1(n2955), .B2(n4400), .ZN(n2957)
         );
  AND2_X1 U3779 ( .A1(n2956), .A2(n2957), .ZN(n3503) );
  INV_X1 U3780 ( .A(n2956), .ZN(n2959) );
  INV_X1 U3781 ( .A(n2957), .ZN(n2958) );
  NAND2_X1 U3782 ( .A1(n2959), .A2(n2958), .ZN(n3504) );
  OAI22_X1 U3783 ( .A1(n4403), .A2(n2955), .B1(n3040), .B2(n3599), .ZN(n2960)
         );
  XNOR2_X1 U3784 ( .A(n2960), .B(n3030), .ZN(n3551) );
  NAND2_X1 U3785 ( .A1(n2961), .A2(n3550), .ZN(n2965) );
  INV_X1 U3786 ( .A(n3549), .ZN(n2963) );
  INV_X1 U3787 ( .A(n3551), .ZN(n2962) );
  NAND2_X1 U3788 ( .A1(n2963), .A2(n2962), .ZN(n2964) );
  NAND2_X1 U3789 ( .A1(n2965), .A2(n2964), .ZN(n3660) );
  OAI22_X1 U3790 ( .A1(n4382), .A2(n2955), .B1(n3040), .B2(n3562), .ZN(n2966)
         );
  XNOR2_X1 U3791 ( .A(n2966), .B(n3038), .ZN(n2967) );
  OAI22_X1 U3792 ( .A1(n4382), .A2(n2882), .B1(n2955), .B2(n3562), .ZN(n2968)
         );
  AND2_X1 U3793 ( .A1(n2967), .A2(n2968), .ZN(n3661) );
  INV_X1 U3794 ( .A(n2967), .ZN(n2970) );
  INV_X1 U3795 ( .A(n2968), .ZN(n2969) );
  NAND2_X1 U3796 ( .A1(n2970), .A2(n2969), .ZN(n3662) );
  OAI22_X1 U3797 ( .A1(n4498), .A2(n2955), .B1(n3580), .B2(n3040), .ZN(n2971)
         );
  XNOR2_X1 U3798 ( .A(n2971), .B(n3030), .ZN(n2977) );
  OAI22_X1 U3799 ( .A1(n4369), .A2(n2955), .B1(n4499), .B2(n3040), .ZN(n2972)
         );
  XNOR2_X1 U3800 ( .A(n2972), .B(n3038), .ZN(n2974) );
  INV_X1 U3801 ( .A(n2974), .ZN(n2976) );
  OAI22_X1 U3802 ( .A1(n4369), .A2(n2882), .B1(n4499), .B2(n2955), .ZN(n2973)
         );
  INV_X1 U3803 ( .A(n2973), .ZN(n2975) );
  OR2_X1 U3804 ( .A1(n2974), .A2(n2973), .ZN(n2979) );
  OAI21_X1 U3805 ( .B1(n2976), .B2(n2975), .A(n2979), .ZN(n4507) );
  OAI22_X1 U3806 ( .A1(n4498), .A2(n2882), .B1(n3580), .B2(n2955), .ZN(n4505)
         );
  OAI22_X1 U3807 ( .A1(n4286), .A2(n2955), .B1(n4273), .B2(n3040), .ZN(n2980)
         );
  XNOR2_X1 U3808 ( .A(n2980), .B(n3038), .ZN(n2982) );
  OAI22_X1 U3809 ( .A1(n4286), .A2(n2882), .B1(n4273), .B2(n2955), .ZN(n2981)
         );
  OR2_X1 U3810 ( .A1(n2982), .A2(n2981), .ZN(n3720) );
  OAI22_X1 U3811 ( .A1(n4228), .A2(n2955), .B1(n4245), .B2(n3040), .ZN(n2983)
         );
  XNOR2_X1 U3812 ( .A(n2983), .B(n3038), .ZN(n2984) );
  OAI22_X1 U3813 ( .A1(n4228), .A2(n2882), .B1(n4245), .B2(n2955), .ZN(n2985)
         );
  NAND2_X1 U3814 ( .A1(n2984), .A2(n2985), .ZN(n3759) );
  NAND2_X1 U3815 ( .A1(n3758), .A2(n3759), .ZN(n3757) );
  INV_X1 U3816 ( .A(n2984), .ZN(n2987) );
  INV_X1 U3817 ( .A(n2985), .ZN(n2986) );
  NAND2_X1 U3818 ( .A1(n2987), .A2(n2986), .ZN(n3761) );
  NAND2_X1 U3819 ( .A1(n4249), .A2(n2877), .ZN(n2989) );
  NAND2_X1 U3820 ( .A1(n4224), .A2(n2878), .ZN(n2988) );
  NAND2_X1 U3821 ( .A1(n2989), .A2(n2988), .ZN(n2990) );
  XNOR2_X1 U3822 ( .A(n2990), .B(n3038), .ZN(n2991) );
  AOI22_X1 U3823 ( .A1(n4249), .A2(n3033), .B1(n2877), .B2(n4224), .ZN(n2992)
         );
  XNOR2_X1 U3824 ( .A(n2991), .B(n2992), .ZN(n3682) );
  INV_X1 U3825 ( .A(n2991), .ZN(n2993) );
  NAND2_X1 U3826 ( .A1(n4225), .A2(n2877), .ZN(n2995) );
  NAND2_X1 U3827 ( .A1(n4350), .A2(n2878), .ZN(n2994) );
  NAND2_X1 U3828 ( .A1(n2995), .A2(n2994), .ZN(n2996) );
  XNOR2_X1 U3829 ( .A(n2996), .B(n3030), .ZN(n3003) );
  AND2_X1 U3830 ( .A1(n4350), .A2(n2242), .ZN(n2997) );
  AOI21_X1 U3831 ( .B1(n4225), .B2(n3033), .A(n2997), .ZN(n3002) );
  NOR2_X1 U3832 ( .A1(n3003), .A2(n3002), .ZN(n3736) );
  NAND2_X1 U3833 ( .A1(n4351), .A2(n2877), .ZN(n2999) );
  NAND2_X1 U3834 ( .A1(n4341), .A2(n2878), .ZN(n2998) );
  NAND2_X1 U3835 ( .A1(n2999), .A2(n2998), .ZN(n3000) );
  XNOR2_X1 U3836 ( .A(n3000), .B(n3030), .ZN(n3688) );
  NOR2_X1 U3837 ( .A1(n4190), .A2(n2955), .ZN(n3001) );
  AOI21_X1 U3838 ( .B1(n4351), .B2(n3033), .A(n3001), .ZN(n3689) );
  NAND2_X1 U3839 ( .A1(n3688), .A2(n3689), .ZN(n3004) );
  NAND2_X1 U3840 ( .A1(n3003), .A2(n3002), .ZN(n3737) );
  OAI22_X1 U3841 ( .A1(n3677), .A2(n2955), .B1(n3752), .B2(n3040), .ZN(n3007)
         );
  XNOR2_X1 U3842 ( .A(n3007), .B(n3038), .ZN(n3009) );
  OAI22_X1 U3843 ( .A1(n3677), .A2(n2882), .B1(n3752), .B2(n2955), .ZN(n3008)
         );
  XNOR2_X1 U3844 ( .A(n3009), .B(n3008), .ZN(n3748) );
  NOR2_X1 U3845 ( .A1(n3009), .A2(n3008), .ZN(n3674) );
  NAND2_X1 U3846 ( .A1(n4324), .A2(n2242), .ZN(n3011) );
  NAND2_X1 U3847 ( .A1(n4154), .A2(n2878), .ZN(n3010) );
  NAND2_X1 U3848 ( .A1(n3011), .A2(n3010), .ZN(n3012) );
  XNOR2_X1 U3849 ( .A(n3012), .B(n3030), .ZN(n3015) );
  NOR2_X1 U3850 ( .A1(n4159), .A2(n2955), .ZN(n3013) );
  AOI21_X1 U3851 ( .B1(n4324), .B2(n3033), .A(n3013), .ZN(n3014) );
  XNOR2_X1 U3852 ( .A(n3015), .B(n3014), .ZN(n3673) );
  NOR2_X1 U3853 ( .A1(n3015), .A2(n3014), .ZN(n3020) );
  NAND2_X1 U3854 ( .A1(n4108), .A2(n3033), .ZN(n3017) );
  NAND2_X1 U3855 ( .A1(n4322), .A2(n2877), .ZN(n3016) );
  NAND2_X1 U3856 ( .A1(n3017), .A2(n3016), .ZN(n3019) );
  OAI22_X1 U3857 ( .A1(n4157), .A2(n2955), .B1(n4134), .B2(n3040), .ZN(n3018)
         );
  XOR2_X1 U3858 ( .A(n3038), .B(n3018), .Z(n3729) );
  NAND2_X1 U3859 ( .A1(n4136), .A2(n2877), .ZN(n3022) );
  INV_X1 U3860 ( .A(n4113), .ZN(n4107) );
  NAND2_X1 U3861 ( .A1(n4107), .A2(n2878), .ZN(n3021) );
  NAND2_X1 U3862 ( .A1(n3022), .A2(n3021), .ZN(n3023) );
  XNOR2_X1 U3863 ( .A(n3023), .B(n3030), .ZN(n3026) );
  NOR2_X1 U3864 ( .A1(n4113), .A2(n2955), .ZN(n3024) );
  AOI21_X1 U3865 ( .B1(n4136), .B2(n3033), .A(n3024), .ZN(n3025) );
  NAND2_X1 U3866 ( .A1(n3026), .A2(n3025), .ZN(n3699) );
  OR2_X1 U3867 ( .A1(n3026), .A2(n3025), .ZN(n3700) );
  NAND2_X1 U3868 ( .A1(n3027), .A2(n3700), .ZN(n3769) );
  NAND2_X1 U3869 ( .A1(n4306), .A2(n2877), .ZN(n3029) );
  NAND2_X1 U3870 ( .A1(n3774), .A2(n2878), .ZN(n3028) );
  NAND2_X1 U3871 ( .A1(n3029), .A2(n3028), .ZN(n3031) );
  XNOR2_X1 U3872 ( .A(n3031), .B(n3030), .ZN(n3035) );
  NOR2_X1 U3873 ( .A1(n4097), .A2(n2955), .ZN(n3032) );
  AOI21_X1 U3874 ( .B1(n4306), .B2(n3033), .A(n3032), .ZN(n3034) );
  NOR2_X1 U3875 ( .A1(n3035), .A2(n3034), .ZN(n3772) );
  NAND2_X1 U3876 ( .A1(n3035), .A2(n3034), .ZN(n3770) );
  OAI22_X1 U3877 ( .A1(n4092), .A2(n2882), .B1(n2955), .B2(n4075), .ZN(n3043)
         );
  OAI22_X1 U3878 ( .A1(n4092), .A2(n2955), .B1(n3040), .B2(n4075), .ZN(n3036)
         );
  XNOR2_X1 U3879 ( .A(n3036), .B(n3038), .ZN(n3044) );
  XOR2_X1 U3880 ( .A(n3043), .B(n3044), .Z(n3634) );
  INV_X1 U3881 ( .A(n3634), .ZN(n3037) );
  OAI22_X1 U3882 ( .A1(n4309), .A2(n2882), .B1(n3091), .B2(n2955), .ZN(n3039)
         );
  XNOR2_X1 U3883 ( .A(n3039), .B(n3038), .ZN(n3042) );
  OAI22_X1 U3884 ( .A1(n4309), .A2(n2955), .B1(n3091), .B2(n3040), .ZN(n3041)
         );
  XNOR2_X1 U3885 ( .A(n3042), .B(n3041), .ZN(n3053) );
  INV_X1 U3886 ( .A(n3053), .ZN(n3055) );
  NAND2_X1 U3887 ( .A1(n3044), .A2(n3043), .ZN(n3054) );
  NAND3_X1 U3888 ( .A1(n3098), .A2(n3045), .A3(n3084), .ZN(n3068) );
  INV_X1 U3889 ( .A(n3068), .ZN(n3051) );
  NAND2_X1 U3890 ( .A1(n3046), .A2(n3204), .ZN(n3048) );
  INV_X1 U3891 ( .A(n3134), .ZN(n3047) );
  NAND2_X1 U3892 ( .A1(n3048), .A2(n3047), .ZN(n3056) );
  INV_X1 U3893 ( .A(n3056), .ZN(n3049) );
  AND2_X1 U3894 ( .A1(n3049), .A2(n3193), .ZN(n3050) );
  NAND2_X1 U3895 ( .A1(n3055), .A2(n2452), .ZN(n3052) );
  AND2_X1 U3896 ( .A1(n3053), .A2(n4508), .ZN(n3074) );
  NOR3_X1 U3897 ( .A1(n3055), .A2(n3781), .A3(n3054), .ZN(n3073) );
  NAND2_X1 U3898 ( .A1(n3056), .A2(n4401), .ZN(n3057) );
  NAND2_X1 U3899 ( .A1(n3068), .A2(n3057), .ZN(n3059) );
  NAND2_X1 U3900 ( .A1(n3059), .A2(n3058), .ZN(n3191) );
  OAI21_X1 U3901 ( .B1(n3191), .B2(n3060), .A(STATE_REG_SCAN_IN), .ZN(n3064)
         );
  NAND2_X1 U3902 ( .A1(n3061), .A2(n4675), .ZN(n3062) );
  NOR2_X1 U3903 ( .A1(n2955), .A2(n3062), .ZN(n3958) );
  NAND2_X1 U3904 ( .A1(n3068), .A2(n3958), .ZN(n3192) );
  OR2_X1 U3905 ( .A1(n3135), .A2(U3149), .ZN(n3962) );
  AND2_X1 U3906 ( .A1(n3192), .A2(n3962), .ZN(n3063) );
  NAND2_X1 U3907 ( .A1(n3958), .A2(n3226), .ZN(n3065) );
  NAND2_X1 U3908 ( .A1(n3958), .A2(n4495), .ZN(n3066) );
  AOI22_X1 U3909 ( .A1(n3967), .A2(n3786), .B1(n4503), .B2(n3965), .ZN(n3071)
         );
  NAND2_X1 U3910 ( .A1(n3193), .A2(n4386), .ZN(n3067) );
  OR2_X1 U3911 ( .A1(n3068), .A2(n3067), .ZN(n3069) );
  NAND2_X1 U3912 ( .A1(n3069), .A2(n4643), .ZN(n3785) );
  AOI22_X1 U3913 ( .A1(n3785), .A2(n3653), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3070) );
  OAI211_X1 U3914 ( .C1(n4513), .C2(n3649), .A(n3071), .B(n3070), .ZN(n3072)
         );
  AOI21_X1 U3915 ( .B1(n3075), .B2(n3074), .A(n2453), .ZN(n3076) );
  NAND2_X1 U3916 ( .A1(n3077), .A2(n3076), .ZN(U3217) );
  INV_X1 U3917 ( .A(n4411), .ZN(n4699) );
  INV_X1 U3918 ( .A(n3965), .ZN(n3650) );
  OAI22_X1 U3919 ( .A1(n3650), .A2(n4402), .B1(n4401), .B2(n3091), .ZN(n3079)
         );
  AOI21_X1 U3920 ( .B1(n4323), .B2(n3967), .A(n3079), .ZN(n3082) );
  XNOR2_X1 U3921 ( .A(n3080), .B(n3832), .ZN(n3081) );
  NAND2_X1 U3922 ( .A1(n3081), .A2(n4289), .ZN(n3647) );
  OAI211_X1 U3923 ( .C1(n3659), .C2(n4699), .A(n3082), .B(n3647), .ZN(n3100)
         );
  NAND2_X1 U3924 ( .A1(n3084), .A2(n3083), .ZN(n3088) );
  NAND4_X1 U3925 ( .A1(n3088), .A2(n3087), .A3(n3086), .A4(n3085), .ZN(n3099)
         );
  MUX2_X1 U3926 ( .A(REG1_REG_28__SCAN_IN), .B(n3100), .S(n4722), .Z(n3090) );
  INV_X1 U3927 ( .A(n3090), .ZN(n3097) );
  NOR2_X1 U3928 ( .A1(n4072), .A2(n3091), .ZN(n3092) );
  NAND2_X1 U3929 ( .A1(n3097), .A2(n3096), .ZN(U3546) );
  MUX2_X1 U3930 ( .A(REG0_REG_28__SCAN_IN), .B(n3100), .S(n4713), .Z(n3101) );
  INV_X1 U3931 ( .A(n3101), .ZN(n3104) );
  NAND2_X1 U3932 ( .A1(n3104), .A2(n3103), .ZN(U3514) );
  INV_X1 U3933 ( .A(n3816), .ZN(n3105) );
  NAND2_X1 U3934 ( .A1(n3105), .A2(n4386), .ZN(n3106) );
  AOI21_X1 U3935 ( .B1(n3109), .B2(n4411), .A(n3108), .ZN(n3113) );
  MUX2_X1 U3936 ( .A(n3110), .B(n3113), .S(n4722), .Z(n3112) );
  NAND2_X1 U3937 ( .A1(n3112), .A2(n3111), .ZN(U3547) );
  INV_X1 U3938 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3114) );
  MUX2_X1 U3939 ( .A(n3114), .B(n3113), .S(n4713), .Z(n3117) );
  NAND2_X1 U3940 ( .A1(n3117), .A2(n3116), .ZN(U3515) );
  INV_X1 U3941 ( .A(n4675), .ZN(n3118) );
  INV_X1 U3942 ( .A(DATAI_21_), .ZN(n4835) );
  NAND2_X1 U3943 ( .A1(n3880), .A2(STATE_REG_SCAN_IN), .ZN(n3120) );
  OAI21_X1 U3944 ( .B1(STATE_REG_SCAN_IN), .B2(n4835), .A(n3120), .ZN(U3331)
         );
  INV_X1 U3945 ( .A(DATAI_25_), .ZN(n4974) );
  NAND2_X1 U3946 ( .A1(n3121), .A2(STATE_REG_SCAN_IN), .ZN(n3122) );
  OAI21_X1 U3947 ( .B1(STATE_REG_SCAN_IN), .B2(n4974), .A(n3122), .ZN(U3327)
         );
  INV_X1 U3948 ( .A(DATAI_19_), .ZN(n5057) );
  MUX2_X1 U3949 ( .A(n5057), .B(n4057), .S(STATE_REG_SCAN_IN), .Z(n3123) );
  INV_X1 U3950 ( .A(n3123), .ZN(U3333) );
  NAND2_X1 U3951 ( .A1(n4518), .A2(STATE_REG_SCAN_IN), .ZN(n3124) );
  OAI21_X1 U3952 ( .B1(STATE_REG_SCAN_IN), .B2(n2760), .A(n3124), .ZN(U3325)
         );
  INV_X1 U3953 ( .A(n3125), .ZN(n3126) );
  AND2_X2 U3954 ( .A1(n3126), .A2(n3193), .ZN(n4674) );
  NAND3_X1 U3955 ( .A1(n3128), .A2(n4675), .A3(n3127), .ZN(n3129) );
  OAI21_X1 U3956 ( .B1(n4674), .B2(D_REG_0__SCAN_IN), .A(n3129), .ZN(n3130) );
  INV_X1 U3957 ( .A(n3130), .ZN(U3458) );
  NAND2_X1 U3958 ( .A1(n4675), .A2(n3131), .ZN(n3132) );
  OAI22_X1 U3959 ( .A1(n4674), .A2(D_REG_1__SCAN_IN), .B1(n4485), .B2(n3132), 
        .ZN(n3133) );
  INV_X1 U3960 ( .A(n3133), .ZN(U3459) );
  AND2_X1 U3961 ( .A1(n3135), .A2(n3134), .ZN(n3136) );
  NOR2_X1 U3962 ( .A1(n2227), .A2(n3136), .ZN(n3149) );
  INV_X1 U3963 ( .A(n3149), .ZN(n3138) );
  INV_X1 U3964 ( .A(n3962), .ZN(n3137) );
  NOR2_X1 U3965 ( .A1(n4629), .A2(U4043), .ZN(U3148) );
  INV_X1 U3966 ( .A(n3174), .ZN(n4491) );
  INV_X1 U3967 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3142) );
  INV_X1 U3968 ( .A(n4494), .ZN(n3232) );
  MUX2_X1 U3969 ( .A(REG2_REG_2__SCAN_IN), .B(n3142), .S(n4494), .Z(n3235) );
  AND2_X1 U3970 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3140)
         );
  NAND2_X1 U3971 ( .A1(n3985), .A2(n3140), .ZN(n3984) );
  NAND2_X1 U3972 ( .A1(n3984), .A2(n3141), .ZN(n3234) );
  XNOR2_X1 U3973 ( .A(n3144), .B(n4492), .ZN(n3269) );
  INV_X1 U3974 ( .A(n3144), .ZN(n3145) );
  MUX2_X1 U3975 ( .A(REG2_REG_5__SCAN_IN), .B(n2543), .S(n3174), .Z(n3171) );
  NOR2_X1 U3976 ( .A1(n3172), .A2(n3171), .ZN(n3170) );
  XNOR2_X1 U3977 ( .A(n3146), .B(n4490), .ZN(n3178) );
  INV_X1 U3978 ( .A(n3146), .ZN(n3147) );
  AOI22_X1 U3979 ( .A1(n3178), .A2(REG2_REG_6__SCAN_IN), .B1(n4490), .B2(n3147), .ZN(n3151) );
  MUX2_X1 U3980 ( .A(n4000), .B(REG2_REG_7__SCAN_IN), .S(n4489), .Z(n3150) );
  INV_X1 U3981 ( .A(n4518), .ZN(n3160) );
  NOR2_X1 U3982 ( .A1(n4495), .A2(n3160), .ZN(n3959) );
  AOI211_X1 U3983 ( .C1(n3151), .C2(n3150), .A(n4624), .B(n4003), .ZN(n3166)
         );
  INV_X1 U3984 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3152) );
  XNOR2_X1 U3985 ( .A(n4494), .B(n3152), .ZN(n3238) );
  INV_X1 U3986 ( .A(REG1_REG_1__SCAN_IN), .ZN(n3153) );
  AND2_X1 U3987 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3981)
         );
  NAND2_X1 U3988 ( .A1(n3982), .A2(n3981), .ZN(n3980) );
  NAND2_X1 U3989 ( .A1(n3980), .A2(n3154), .ZN(n3237) );
  NAND2_X1 U3990 ( .A1(n3238), .A2(n3237), .ZN(n3236) );
  NAND2_X1 U3991 ( .A1(n4494), .A2(REG1_REG_2__SCAN_IN), .ZN(n3155) );
  XNOR2_X1 U3992 ( .A(n3156), .B(n3143), .ZN(n3991) );
  NAND2_X1 U3993 ( .A1(n3991), .A2(REG1_REG_3__SCAN_IN), .ZN(n3990) );
  NAND2_X1 U3994 ( .A1(n3156), .A2(n4493), .ZN(n3157) );
  NAND2_X1 U3995 ( .A1(n3990), .A2(n3157), .ZN(n3158) );
  INV_X1 U3996 ( .A(n4492), .ZN(n3274) );
  XNOR2_X1 U3997 ( .A(n3158), .B(n3274), .ZN(n3271) );
  XNOR2_X1 U3998 ( .A(n4491), .B(REG1_REG_5__SCAN_IN), .ZN(n3168) );
  INV_X1 U3999 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3407) );
  NOR2_X1 U4000 ( .A1(n3183), .A2(n3407), .ZN(n3181) );
  XNOR2_X1 U4001 ( .A(n4489), .B(REG1_REG_7__SCAN_IN), .ZN(n3162) );
  OAI21_X1 U4002 ( .B1(n4029), .B2(n3162), .A(n4631), .ZN(n3161) );
  AOI21_X1 U4003 ( .B1(n4029), .B2(n3162), .A(n3161), .ZN(n3165) );
  INV_X1 U4004 ( .A(n4489), .ZN(n4001) );
  INV_X1 U4005 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4994) );
  NOR2_X1 U4006 ( .A1(STATE_REG_SCAN_IN), .A2(n4994), .ZN(n3366) );
  AOI21_X1 U4007 ( .B1(n4629), .B2(ADDR_REG_7__SCAN_IN), .A(n3366), .ZN(n3163)
         );
  OAI21_X1 U4008 ( .B1(n4001), .B2(n4635), .A(n3163), .ZN(n3164) );
  OR3_X1 U4009 ( .A1(n3166), .A2(n3165), .A3(n3164), .ZN(U3247) );
  INV_X1 U4010 ( .A(n4631), .ZN(n3182) );
  AOI211_X1 U4011 ( .C1(n3169), .C2(n3168), .A(n3167), .B(n3182), .ZN(n3177)
         );
  AOI211_X1 U4012 ( .C1(n3172), .C2(n3171), .A(n3170), .B(n4624), .ZN(n3176)
         );
  INV_X1 U4013 ( .A(REG3_REG_5__SCAN_IN), .ZN(n4995) );
  NOR2_X1 U4014 ( .A1(STATE_REG_SCAN_IN), .A2(n4995), .ZN(n3713) );
  AOI21_X1 U4015 ( .B1(n4629), .B2(ADDR_REG_5__SCAN_IN), .A(n3713), .ZN(n3173)
         );
  OAI21_X1 U4016 ( .B1(n3174), .B2(n4635), .A(n3173), .ZN(n3175) );
  OR3_X1 U4017 ( .A1(n3177), .A2(n3176), .A3(n3175), .ZN(U3245) );
  XNOR2_X1 U4018 ( .A(n3178), .B(REG2_REG_6__SCAN_IN), .ZN(n3187) );
  INV_X1 U4019 ( .A(n4635), .ZN(n3992) );
  NOR2_X1 U4020 ( .A1(STATE_REG_SCAN_IN), .A2(n3179), .ZN(n3293) );
  AOI21_X1 U4021 ( .B1(n4629), .B2(ADDR_REG_6__SCAN_IN), .A(n3293), .ZN(n3180)
         );
  INV_X1 U4022 ( .A(n3180), .ZN(n3185) );
  AOI211_X1 U4023 ( .C1(n3407), .C2(n3183), .A(n3182), .B(n3181), .ZN(n3184)
         );
  AOI211_X1 U4024 ( .C1(n3992), .C2(n4490), .A(n3185), .B(n3184), .ZN(n3186)
         );
  OAI21_X1 U4025 ( .B1(n3187), .B2(n4624), .A(n3186), .ZN(U3246) );
  OAI21_X1 U4026 ( .B1(n3190), .B2(n3189), .A(n3188), .ZN(n3227) );
  INV_X1 U4027 ( .A(n3191), .ZN(n3194) );
  NAND3_X1 U4028 ( .A1(n3194), .A2(n3193), .A3(n3192), .ZN(n3221) );
  OAI22_X1 U4029 ( .A1(n4500), .A2(n3254), .B1(n3352), .B2(n3777), .ZN(n3195)
         );
  AOI21_X1 U4030 ( .B1(REG3_REG_0__SCAN_IN), .B2(n3221), .A(n3195), .ZN(n3196)
         );
  OAI21_X1 U4031 ( .B1(n3227), .B2(n3781), .A(n3196), .ZN(U3229) );
  INV_X1 U4032 ( .A(n3221), .ZN(n3203) );
  INV_X1 U4033 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3255) );
  OAI211_X1 U4034 ( .C1(n3197), .C2(n3198), .A(n3199), .B(n4508), .ZN(n3202)
         );
  OAI22_X1 U4035 ( .A1(n3207), .A2(n4497), .B1(n3312), .B2(n3777), .ZN(n3200)
         );
  AOI21_X1 U4036 ( .B1(n3256), .B2(n3785), .A(n3200), .ZN(n3201) );
  OAI211_X1 U4037 ( .C1(n3203), .C2(n3255), .A(n3202), .B(n3201), .ZN(U3219)
         );
  INV_X1 U4038 ( .A(n3204), .ZN(n3205) );
  NOR2_X1 U4039 ( .A1(n3254), .A2(n3205), .ZN(n4687) );
  NOR2_X1 U4040 ( .A1(n3207), .A2(n3206), .ZN(n3876) );
  INV_X1 U4041 ( .A(n3261), .ZN(n3879) );
  NOR2_X1 U4042 ( .A1(n3876), .A2(n3879), .ZN(n3865) );
  NOR2_X1 U40430 ( .A1(n3561), .A2(n4289), .ZN(n3208) );
  OAI22_X1 U4044 ( .A1(n3865), .A2(n3208), .B1(n3352), .B2(n4402), .ZN(n4686)
         );
  AOI21_X1 U4045 ( .B1(n4687), .B2(n3209), .A(n4686), .ZN(n3214) );
  INV_X1 U4046 ( .A(n3865), .ZN(n4688) );
  NAND2_X1 U4047 ( .A1(n4646), .A2(n3210), .ZN(n3529) );
  OAI22_X1 U4048 ( .A1(n4646), .A2(n3224), .B1(n3211), .B2(n4643), .ZN(n3212)
         );
  AOI21_X1 U4049 ( .B1(n4688), .B2(n4658), .A(n3212), .ZN(n3213) );
  OAI21_X1 U4050 ( .B1(n3214), .B2(n4663), .A(n3213), .ZN(U3290) );
  INV_X1 U4051 ( .A(n3217), .ZN(n3218) );
  AOI21_X1 U4052 ( .B1(n3215), .B2(n3216), .A(n3218), .ZN(n3223) );
  AOI22_X1 U4053 ( .A1(n2510), .A2(n3786), .B1(n4503), .B2(n2890), .ZN(n3219)
         );
  OAI21_X1 U4054 ( .B1(n4500), .B2(n3351), .A(n3219), .ZN(n3220) );
  AOI21_X1 U4055 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3221), .A(n3220), .ZN(n3222)
         );
  OAI21_X1 U4056 ( .B1(n3223), .B2(n3781), .A(n3222), .ZN(U3234) );
  INV_X1 U4057 ( .A(IR_REG_0__SCAN_IN), .ZN(n4986) );
  NAND2_X1 U4058 ( .A1(n4518), .A2(n3224), .ZN(n3225) );
  NAND2_X1 U4059 ( .A1(n3226), .A2(n3225), .ZN(n4519) );
  NAND2_X1 U4060 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3983) );
  NOR2_X1 U4061 ( .A1(n3227), .A2(n4518), .ZN(n3228) );
  AOI211_X1 U4062 ( .C1(n4518), .C2(n3983), .A(n4495), .B(n3228), .ZN(n3229)
         );
  AOI211_X1 U4063 ( .C1(n4986), .C2(n4519), .A(n3979), .B(n3229), .ZN(n3275)
         );
  NAND2_X1 U4064 ( .A1(U3149), .A2(REG3_REG_2__SCAN_IN), .ZN(n3231) );
  NAND2_X1 U4065 ( .A1(n4629), .A2(ADDR_REG_2__SCAN_IN), .ZN(n3230) );
  OAI211_X1 U4066 ( .C1(n4635), .C2(n3232), .A(n3231), .B(n3230), .ZN(n3242)
         );
  OAI211_X1 U4067 ( .C1(n3235), .C2(n3234), .A(n4575), .B(n3233), .ZN(n3240)
         );
  OAI211_X1 U4068 ( .C1(n3238), .C2(n3237), .A(n4631), .B(n3236), .ZN(n3239)
         );
  NAND2_X1 U4069 ( .A1(n3240), .A2(n3239), .ZN(n3241) );
  OR3_X1 U4070 ( .A1(n3275), .A2(n3242), .A3(n3241), .ZN(U3242) );
  NAND2_X1 U4071 ( .A1(n3217), .A2(n3244), .ZN(n3245) );
  XOR2_X1 U4072 ( .A(n3243), .B(n3245), .Z(n3249) );
  OAI22_X1 U4073 ( .A1(n3312), .A2(n4497), .B1(n3322), .B2(n3777), .ZN(n3247)
         );
  INV_X1 U4074 ( .A(n4513), .ZN(n3779) );
  MUX2_X1 U4075 ( .A(n3779), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n3246) );
  AOI211_X1 U4076 ( .C1(n3311), .C2(n3785), .A(n3247), .B(n3246), .ZN(n3248)
         );
  OAI21_X1 U4077 ( .B1(n3249), .B2(n3781), .A(n3248), .ZN(U3215) );
  OR2_X1 U4078 ( .A1(n3250), .A2(n2823), .ZN(n3251) );
  NAND2_X1 U4079 ( .A1(n3252), .A2(n3251), .ZN(n4691) );
  INV_X1 U4080 ( .A(n4691), .ZN(n3267) );
  OAI21_X1 U4081 ( .B1(n3254), .B2(n3253), .A(n3359), .ZN(n4689) );
  OAI22_X1 U4082 ( .A1(n4233), .A2(n4689), .B1(n3255), .B2(n4643), .ZN(n3266)
         );
  NAND2_X1 U4083 ( .A1(n3256), .A2(n4386), .ZN(n3259) );
  NAND2_X1 U4084 ( .A1(n3257), .A2(n4323), .ZN(n3258) );
  OAI211_X1 U4085 ( .C1(n3312), .C2(n4402), .A(n3259), .B(n3258), .ZN(n3260)
         );
  INV_X1 U4086 ( .A(n3260), .ZN(n3264) );
  XNOR2_X1 U4087 ( .A(n2823), .B(n3261), .ZN(n3262) );
  NAND2_X1 U4088 ( .A1(n3262), .A2(n4289), .ZN(n3263) );
  OAI211_X1 U4089 ( .C1(n4691), .C2(n3517), .A(n3264), .B(n3263), .ZN(n4693)
         );
  MUX2_X1 U4090 ( .A(n4693), .B(REG2_REG_1__SCAN_IN), .S(n4663), .Z(n3265) );
  AOI211_X1 U4091 ( .C1(n3267), .C2(n4658), .A(n3266), .B(n3265), .ZN(n3268)
         );
  INV_X1 U4092 ( .A(n3268), .ZN(U3289) );
  XOR2_X1 U4093 ( .A(REG2_REG_4__SCAN_IN), .B(n3269), .Z(n3277) );
  OAI211_X1 U4094 ( .C1(n3271), .C2(REG1_REG_4__SCAN_IN), .A(n4631), .B(n3270), 
        .ZN(n3273) );
  AND2_X1 U4095 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3630) );
  AOI21_X1 U4096 ( .B1(n4629), .B2(ADDR_REG_4__SCAN_IN), .A(n3630), .ZN(n3272)
         );
  OAI211_X1 U4097 ( .C1(n4635), .C2(n3274), .A(n3273), .B(n3272), .ZN(n3276)
         );
  AOI211_X1 U4098 ( .C1(n4575), .C2(n3277), .A(n3276), .B(n3275), .ZN(n3278)
         );
  INV_X1 U4099 ( .A(n3278), .ZN(U3244) );
  XOR2_X1 U4100 ( .A(n3279), .B(n3849), .Z(n3320) );
  XNOR2_X1 U4101 ( .A(n3280), .B(n3849), .ZN(n3281) );
  NAND2_X1 U4102 ( .A1(n3281), .A2(n4289), .ZN(n3318) );
  AOI22_X1 U4103 ( .A1(n2540), .A2(n4388), .B1(n4386), .B2(n3311), .ZN(n3282)
         );
  OAI211_X1 U4104 ( .C1(n3312), .C2(n4407), .A(n3318), .B(n3282), .ZN(n3283)
         );
  AOI21_X1 U4105 ( .B1(n3320), .B2(n4411), .A(n3283), .ZN(n3288) );
  INV_X1 U4106 ( .A(n3358), .ZN(n3285) );
  INV_X1 U4107 ( .A(n3373), .ZN(n3284) );
  AOI21_X1 U4108 ( .B1(n3311), .B2(n3285), .A(n3284), .ZN(n3315) );
  AOI22_X1 U4109 ( .A1(n3315), .A2(n3094), .B1(REG1_REG_3__SCAN_IN), .B2(n4719), .ZN(n3286) );
  OAI21_X1 U4110 ( .B1(n3288), .B2(n4719), .A(n3286), .ZN(U3521) );
  AOI22_X1 U4111 ( .A1(n3315), .A2(n3102), .B1(REG0_REG_3__SCAN_IN), .B2(n4711), .ZN(n3287) );
  OAI21_X1 U4112 ( .B1(n3288), .B2(n4711), .A(n3287), .ZN(U3473) );
  XNOR2_X1 U4113 ( .A(n3291), .B(n3290), .ZN(n3292) );
  XNOR2_X1 U4114 ( .A(n3289), .B(n3292), .ZN(n3297) );
  AOI21_X1 U4115 ( .B1(n3975), .B2(n4503), .A(n3293), .ZN(n3295) );
  AOI22_X1 U4116 ( .A1(n3977), .A2(n3786), .B1(n3336), .B2(n3785), .ZN(n3294)
         );
  OAI211_X1 U4117 ( .C1(n4513), .C2(n3339), .A(n3295), .B(n3294), .ZN(n3296)
         );
  AOI21_X1 U4118 ( .B1(n3297), .B2(n4508), .A(n3296), .ZN(n3298) );
  INV_X1 U4119 ( .A(n3298), .ZN(U3236) );
  XNOR2_X1 U4120 ( .A(n2905), .B(n3714), .ZN(n3866) );
  NAND2_X1 U4121 ( .A1(n3299), .A2(n3300), .ZN(n3381) );
  NAND2_X1 U4122 ( .A1(n3381), .A2(n3301), .ZN(n3302) );
  XOR2_X1 U4123 ( .A(n3866), .B(n3302), .Z(n3330) );
  XNOR2_X1 U4124 ( .A(n3303), .B(n3866), .ZN(n3304) );
  NAND2_X1 U4125 ( .A1(n3304), .A2(n4289), .ZN(n3328) );
  AOI22_X1 U4126 ( .A1(n3976), .A2(n4388), .B1(n4386), .B2(n3714), .ZN(n3305)
         );
  OAI211_X1 U4127 ( .C1(n3322), .C2(n4407), .A(n3328), .B(n3305), .ZN(n3306)
         );
  AOI21_X1 U4128 ( .B1(n3330), .B2(n4411), .A(n3306), .ZN(n3310) );
  INV_X1 U4129 ( .A(n3372), .ZN(n3307) );
  AOI21_X1 U4130 ( .B1(n3714), .B2(n3307), .A(n2279), .ZN(n3325) );
  AOI22_X1 U4131 ( .A1(n3325), .A2(n3102), .B1(REG0_REG_5__SCAN_IN), .B2(n4711), .ZN(n3308) );
  OAI21_X1 U4132 ( .B1(n3310), .B2(n4711), .A(n3308), .ZN(U3477) );
  AOI22_X1 U4133 ( .A1(n3325), .A2(n3094), .B1(REG1_REG_5__SCAN_IN), .B2(n4719), .ZN(n3309) );
  OAI21_X1 U4134 ( .B1(n3310), .B2(n4719), .A(n3309), .ZN(U3523) );
  NAND2_X1 U4135 ( .A1(n4646), .A2(n4388), .ZN(n4081) );
  INV_X1 U4136 ( .A(n4081), .ZN(n4266) );
  INV_X1 U4137 ( .A(n4272), .ZN(n4206) );
  AOI22_X1 U4138 ( .A1(n2540), .A2(n4266), .B1(n4206), .B2(n3311), .ZN(n3317)
         );
  OAI22_X1 U4139 ( .A1(n4646), .A2(n3993), .B1(REG3_REG_3__SCAN_IN), .B2(n4643), .ZN(n3314) );
  INV_X1 U4140 ( .A(n4267), .ZN(n4210) );
  NOR2_X1 U4141 ( .A1(n4210), .A2(n3312), .ZN(n3313) );
  AOI211_X1 U4142 ( .C1(n3315), .C2(n4657), .A(n3314), .B(n3313), .ZN(n3316)
         );
  OAI211_X1 U4143 ( .C1(n3318), .C2(n4663), .A(n3317), .B(n3316), .ZN(n3319)
         );
  AOI21_X1 U4144 ( .B1(n4264), .B2(n3320), .A(n3319), .ZN(n3321) );
  INV_X1 U4145 ( .A(n3321), .ZN(U3287) );
  OAI22_X1 U4146 ( .A1(n4646), .A2(n2543), .B1(n3715), .B2(n4643), .ZN(n3324)
         );
  OAI22_X1 U4147 ( .A1(n4210), .A2(n3322), .B1(n2563), .B2(n4081), .ZN(n3323)
         );
  AOI211_X1 U4148 ( .C1(n3714), .C2(n4206), .A(n3324), .B(n3323), .ZN(n3327)
         );
  NAND2_X1 U4149 ( .A1(n3325), .A2(n4657), .ZN(n3326) );
  OAI211_X1 U4150 ( .C1(n3328), .C2(n4663), .A(n3327), .B(n3326), .ZN(n3329)
         );
  AOI21_X1 U4151 ( .B1(n4264), .B2(n3330), .A(n3329), .ZN(n3331) );
  INV_X1 U4152 ( .A(n3331), .ZN(U3285) );
  NAND2_X1 U4153 ( .A1(n3894), .A2(n3890), .ZN(n3829) );
  XNOR2_X1 U4154 ( .A(n2269), .B(n3829), .ZN(n3403) );
  XNOR2_X1 U4155 ( .A(n3334), .B(n3829), .ZN(n3335) );
  NOR2_X1 U4156 ( .A1(n3335), .A2(n3522), .ZN(n3400) );
  NAND2_X1 U4157 ( .A1(n3337), .A2(n3336), .ZN(n3338) );
  NAND2_X1 U4158 ( .A1(n3437), .A2(n3338), .ZN(n3408) );
  OAI22_X1 U4159 ( .A1(n4646), .A2(n3340), .B1(n3339), .B2(n4643), .ZN(n3341)
         );
  AOI21_X1 U4160 ( .B1(n3977), .B2(n4267), .A(n3341), .ZN(n3344) );
  OAI22_X1 U4161 ( .A1(n3478), .A2(n4081), .B1(n4272), .B2(n2278), .ZN(n3342)
         );
  INV_X1 U4162 ( .A(n3342), .ZN(n3343) );
  OAI211_X1 U4163 ( .C1(n3408), .C2(n4233), .A(n3344), .B(n3343), .ZN(n3345)
         );
  AOI21_X1 U4164 ( .B1(n3400), .B2(n4646), .A(n3345), .ZN(n3346) );
  OAI21_X1 U4165 ( .B1(n4295), .B2(n3403), .A(n3346), .ZN(U3284) );
  INV_X1 U4166 ( .A(n4705), .ZN(n4697) );
  INV_X1 U4167 ( .A(n3347), .ZN(n3348) );
  AOI21_X1 U4168 ( .B1(n3851), .B2(n3349), .A(n3348), .ZN(n3353) );
  INV_X1 U4169 ( .A(n3353), .ZN(n4659) );
  XOR2_X1 U4170 ( .A(n3851), .B(n3350), .Z(n3357) );
  OAI22_X1 U4171 ( .A1(n3352), .A2(n4407), .B1(n3351), .B2(n4401), .ZN(n3355)
         );
  NOR2_X1 U4172 ( .A1(n3353), .A2(n3517), .ZN(n3354) );
  AOI211_X1 U4173 ( .C1(n4388), .C2(n2890), .A(n3355), .B(n3354), .ZN(n3356)
         );
  OAI21_X1 U4174 ( .B1(n3522), .B2(n3357), .A(n3356), .ZN(n4654) );
  AOI21_X1 U4175 ( .B1(n4697), .B2(n4659), .A(n4654), .ZN(n3363) );
  AOI21_X1 U4176 ( .B1(n3360), .B2(n3359), .A(n3358), .ZN(n4656) );
  AOI22_X1 U4177 ( .A1(n4656), .A2(n3094), .B1(REG1_REG_2__SCAN_IN), .B2(n4719), .ZN(n3361) );
  OAI21_X1 U4178 ( .B1(n3363), .B2(n4719), .A(n3361), .ZN(U3520) );
  AOI22_X1 U4179 ( .A1(n4656), .A2(n3102), .B1(n4711), .B2(REG0_REG_2__SCAN_IN), .ZN(n3362) );
  OAI21_X1 U4180 ( .B1(n3363), .B2(n4711), .A(n3362), .ZN(U3471) );
  XOR2_X1 U4181 ( .A(n3364), .B(n3365), .Z(n3370) );
  AOI21_X1 U4182 ( .B1(n3974), .B2(n4503), .A(n3366), .ZN(n3368) );
  AOI22_X1 U4183 ( .A1(n3786), .A2(n3976), .B1(n3785), .B2(n3438), .ZN(n3367)
         );
  OAI211_X1 U4184 ( .C1(n4513), .C2(n3446), .A(n3368), .B(n3367), .ZN(n3369)
         );
  AOI21_X1 U4185 ( .B1(n3370), .B2(n4508), .A(n3369), .ZN(n3371) );
  INV_X1 U4186 ( .A(n3371), .ZN(U3210) );
  INV_X1 U4187 ( .A(n4710), .ZN(n4690) );
  AOI211_X1 U4188 ( .C1(n3374), .C2(n3373), .A(n4690), .B(n3372), .ZN(n4696)
         );
  NOR2_X1 U4189 ( .A1(n4643), .A2(n3633), .ZN(n3386) );
  XNOR2_X1 U4190 ( .A(n3376), .B(n3845), .ZN(n3385) );
  NAND2_X1 U4191 ( .A1(n2890), .A2(n4323), .ZN(n3377) );
  OAI21_X1 U4192 ( .B1(n4401), .B2(n3628), .A(n3377), .ZN(n3383) );
  NAND2_X1 U4193 ( .A1(n3299), .A2(n3378), .ZN(n3379) );
  NAND2_X1 U4194 ( .A1(n3379), .A2(n3845), .ZN(n3380) );
  NAND2_X1 U4195 ( .A1(n3381), .A2(n3380), .ZN(n3387) );
  NOR2_X1 U4196 ( .A1(n3387), .A2(n3517), .ZN(n3382) );
  AOI211_X1 U4197 ( .C1(n4388), .C2(n3977), .A(n3383), .B(n3382), .ZN(n3384)
         );
  OAI21_X1 U4198 ( .B1(n3522), .B2(n3385), .A(n3384), .ZN(n4695) );
  AOI211_X1 U4199 ( .C1(n4696), .C2(n4057), .A(n3386), .B(n4695), .ZN(n3389)
         );
  INV_X1 U4200 ( .A(n3387), .ZN(n4698) );
  AOI22_X1 U4201 ( .A1(n4698), .A2(n4658), .B1(REG2_REG_4__SCAN_IN), .B2(n4663), .ZN(n3388) );
  OAI21_X1 U4202 ( .B1(n3389), .B2(n4663), .A(n3388), .ZN(U3286) );
  INV_X1 U4203 ( .A(n3412), .ZN(n3391) );
  NAND2_X1 U4204 ( .A1(n3391), .A2(n3413), .ZN(n3392) );
  XNOR2_X1 U4205 ( .A(n3390), .B(n3392), .ZN(n3398) );
  NAND2_X1 U4206 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n4526) );
  INV_X1 U4207 ( .A(n4526), .ZN(n3393) );
  AOI21_X1 U4208 ( .B1(n4503), .B2(n3973), .A(n3393), .ZN(n3396) );
  AOI22_X1 U4209 ( .A1(n3975), .A2(n3786), .B1(n3394), .B2(n3785), .ZN(n3395)
         );
  OAI211_X1 U4210 ( .C1(n4513), .C2(n4644), .A(n3396), .B(n3395), .ZN(n3397)
         );
  AOI21_X1 U4211 ( .B1(n3398), .B2(n4508), .A(n3397), .ZN(n3399) );
  INV_X1 U4212 ( .A(n3399), .ZN(U3218) );
  OAI22_X1 U4213 ( .A1(n3478), .A2(n4402), .B1(n4401), .B2(n2278), .ZN(n3401)
         );
  AOI211_X1 U4214 ( .C1(n4323), .C2(n3977), .A(n3401), .B(n3400), .ZN(n3402)
         );
  OAI21_X1 U4215 ( .B1(n4699), .B2(n3403), .A(n3402), .ZN(n3410) );
  INV_X1 U4216 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3404) );
  OAI22_X1 U4217 ( .A1(n3408), .A2(n4478), .B1(n4713), .B2(n3404), .ZN(n3405)
         );
  AOI21_X1 U4218 ( .B1(n3410), .B2(n4713), .A(n3405), .ZN(n3406) );
  INV_X1 U4219 ( .A(n3406), .ZN(U3479) );
  OAI22_X1 U4220 ( .A1(n3408), .A2(n4414), .B1(n4722), .B2(n3407), .ZN(n3409)
         );
  AOI21_X1 U4221 ( .B1(n3410), .B2(n4722), .A(n3409), .ZN(n3411) );
  INV_X1 U4222 ( .A(n3411), .ZN(U3524) );
  OR2_X1 U4223 ( .A1(n3390), .A2(n3412), .ZN(n3414) );
  NAND2_X1 U4224 ( .A1(n3414), .A2(n3413), .ZN(n3416) );
  XNOR2_X1 U4225 ( .A(n3416), .B(n3415), .ZN(n3420) );
  NOR2_X1 U4226 ( .A1(STATE_REG_SCAN_IN), .A2(n2584), .ZN(n4542) );
  AOI21_X1 U4227 ( .B1(n4503), .B2(n3972), .A(n4542), .ZN(n3418) );
  AOI22_X1 U4228 ( .A1(n3974), .A2(n3786), .B1(n3429), .B2(n3785), .ZN(n3417)
         );
  OAI211_X1 U4229 ( .C1(n4513), .C2(n3431), .A(n3418), .B(n3417), .ZN(n3419)
         );
  AOI21_X1 U4230 ( .B1(n3420), .B2(n4508), .A(n3419), .ZN(n3421) );
  INV_X1 U4231 ( .A(n3421), .ZN(U3228) );
  INV_X1 U4232 ( .A(n3908), .ZN(n3905) );
  NAND2_X1 U4233 ( .A1(n3905), .A2(n3902), .ZN(n3830) );
  XNOR2_X1 U4234 ( .A(n3422), .B(n3830), .ZN(n3423) );
  NAND2_X1 U4235 ( .A1(n3423), .A2(n4289), .ZN(n3492) );
  OR2_X1 U4236 ( .A1(n3424), .A2(n3425), .ZN(n3427) );
  NAND2_X1 U4237 ( .A1(n3427), .A2(n3426), .ZN(n3428) );
  XOR2_X1 U4238 ( .A(n3830), .B(n3428), .Z(n3495) );
  NAND2_X1 U4239 ( .A1(n3495), .A2(n4264), .ZN(n3436) );
  OAI21_X1 U4240 ( .B1(n3471), .B2(n3489), .A(n3530), .ZN(n3501) );
  INV_X1 U4241 ( .A(n3501), .ZN(n3434) );
  AOI22_X1 U4242 ( .A1(n4206), .A2(n3429), .B1(n4266), .B2(n3972), .ZN(n3430)
         );
  OAI21_X1 U4243 ( .B1(n3493), .B2(n4210), .A(n3430), .ZN(n3433) );
  OAI22_X1 U4244 ( .A1(n3431), .A2(n4643), .B1(n2588), .B2(n4646), .ZN(n3432)
         );
  AOI211_X1 U4245 ( .C1(n3434), .C2(n4657), .A(n3433), .B(n3432), .ZN(n3435)
         );
  OAI211_X1 U4246 ( .C1(n4663), .C2(n3492), .A(n3436), .B(n3435), .ZN(U3281)
         );
  AOI211_X1 U4247 ( .C1(n3438), .C2(n3437), .A(n4690), .B(n3473), .ZN(n4702)
         );
  OAI22_X1 U4248 ( .A1(n3493), .A2(n4402), .B1(n3439), .B2(n4401), .ZN(n3444)
         );
  XOR2_X1 U4249 ( .A(n3846), .B(n3441), .Z(n3442) );
  NOR2_X1 U4250 ( .A1(n3442), .A2(n3522), .ZN(n3443) );
  AOI211_X1 U4251 ( .C1(n4323), .C2(n3976), .A(n3444), .B(n3443), .ZN(n3445)
         );
  INV_X1 U4252 ( .A(n3445), .ZN(n4701) );
  AOI21_X1 U4253 ( .B1(n4702), .B2(n4057), .A(n4701), .ZN(n3450) );
  AND2_X1 U4254 ( .A1(n3424), .A2(n3846), .ZN(n4700) );
  NOR2_X1 U4255 ( .A1(n4700), .A2(n4295), .ZN(n3448) );
  OR2_X1 U4256 ( .A1(n3424), .A2(n3846), .ZN(n4703) );
  OAI22_X1 U4257 ( .A1(n4646), .A2(n4000), .B1(n3446), .B2(n4643), .ZN(n3447)
         );
  AOI21_X1 U4258 ( .B1(n3448), .B2(n4703), .A(n3447), .ZN(n3449) );
  OAI21_X1 U4259 ( .B1(n3450), .B2(n4663), .A(n3449), .ZN(U3283) );
  INV_X1 U4260 ( .A(n3451), .ZN(n3452) );
  AOI211_X1 U4261 ( .C1(n3454), .C2(n3453), .A(n3781), .B(n3452), .ZN(n3461)
         );
  NAND2_X1 U4262 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4547) );
  INV_X1 U4263 ( .A(n4547), .ZN(n3455) );
  AOI21_X1 U4264 ( .B1(n3786), .B2(n3973), .A(n3455), .ZN(n3458) );
  AOI22_X1 U4265 ( .A1(n3971), .A2(n4503), .B1(n3456), .B2(n3785), .ZN(n3457)
         );
  OAI211_X1 U4266 ( .C1(n4513), .C2(n3459), .A(n3458), .B(n3457), .ZN(n3460)
         );
  OR2_X1 U4267 ( .A1(n3461), .A2(n3460), .ZN(U3214) );
  XNOR2_X1 U4268 ( .A(n3464), .B(n3463), .ZN(n3465) );
  XNOR2_X1 U4269 ( .A(n3462), .B(n3465), .ZN(n3469) );
  AND2_X1 U4270 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4563) );
  AOI21_X1 U4271 ( .B1(n3786), .B2(n3972), .A(n4563), .ZN(n3467) );
  AOI22_X1 U4272 ( .A1(n3970), .A2(n4503), .B1(n3524), .B2(n3785), .ZN(n3466)
         );
  OAI211_X1 U4273 ( .C1(n4513), .C2(n3525), .A(n3467), .B(n3466), .ZN(n3468)
         );
  AOI21_X1 U4274 ( .B1(n3469), .B2(n4508), .A(n3468), .ZN(n3470) );
  INV_X1 U4275 ( .A(n3470), .ZN(U3233) );
  INV_X1 U4276 ( .A(n3471), .ZN(n3472) );
  OAI21_X1 U4277 ( .B1(n3473), .B2(n3477), .A(n3472), .ZN(n4648) );
  INV_X1 U4278 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3484) );
  NAND2_X1 U4279 ( .A1(n4703), .A2(n3474), .ZN(n3475) );
  XNOR2_X1 U4280 ( .A(n3475), .B(n3842), .ZN(n4650) );
  XNOR2_X1 U4281 ( .A(n3476), .B(n3842), .ZN(n3481) );
  OAI22_X1 U4282 ( .A1(n3478), .A2(n4407), .B1(n4401), .B2(n3477), .ZN(n3479)
         );
  AOI21_X1 U4283 ( .B1(n4388), .B2(n3973), .A(n3479), .ZN(n3480) );
  OAI21_X1 U4284 ( .B1(n3481), .B2(n3522), .A(n3480), .ZN(n3482) );
  AOI21_X1 U4285 ( .B1(n3561), .B2(n4650), .A(n3482), .ZN(n4653) );
  INV_X1 U4286 ( .A(n4653), .ZN(n3483) );
  AOI21_X1 U4287 ( .B1(n4697), .B2(n4650), .A(n3483), .ZN(n3486) );
  MUX2_X1 U4288 ( .A(n3484), .B(n3486), .S(n4713), .Z(n3485) );
  OAI21_X1 U4289 ( .B1(n4648), .B2(n4478), .A(n3485), .ZN(U3483) );
  INV_X1 U4290 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3487) );
  MUX2_X1 U4291 ( .A(n3487), .B(n3486), .S(n4722), .Z(n3488) );
  OAI21_X1 U4292 ( .B1(n4648), .B2(n4414), .A(n3488), .ZN(U3526) );
  INV_X1 U4293 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3496) );
  NOR2_X1 U4294 ( .A1(n3489), .A2(n4401), .ZN(n3490) );
  AOI21_X1 U4295 ( .B1(n3972), .B2(n4388), .A(n3490), .ZN(n3491) );
  OAI211_X1 U4296 ( .C1(n3493), .C2(n4407), .A(n3492), .B(n3491), .ZN(n3494)
         );
  AOI21_X1 U4297 ( .B1(n3495), .B2(n4411), .A(n3494), .ZN(n3498) );
  MUX2_X1 U4298 ( .A(n3496), .B(n3498), .S(n4722), .Z(n3497) );
  OAI21_X1 U4299 ( .B1(n4414), .B2(n3501), .A(n3497), .ZN(U3527) );
  INV_X1 U4300 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3499) );
  MUX2_X1 U4301 ( .A(n3499), .B(n3498), .S(n4713), .Z(n3500) );
  OAI21_X1 U4302 ( .B1(n3501), .B2(n4478), .A(n3500), .ZN(U3485) );
  INV_X1 U4303 ( .A(n3503), .ZN(n3505) );
  NAND2_X1 U4304 ( .A1(n3505), .A2(n3504), .ZN(n3506) );
  XNOR2_X1 U4305 ( .A(n3502), .B(n3506), .ZN(n3510) );
  INV_X1 U4306 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4807) );
  NOR2_X1 U4307 ( .A1(STATE_REG_SCAN_IN), .A2(n4807), .ZN(n4572) );
  AOI21_X1 U4308 ( .B1(n3971), .B2(n3786), .A(n4572), .ZN(n3508) );
  AOI22_X1 U4309 ( .A1(n3969), .A2(n4503), .B1(n3617), .B2(n3785), .ZN(n3507)
         );
  OAI211_X1 U4310 ( .C1(n4513), .C2(n3613), .A(n3508), .B(n3507), .ZN(n3509)
         );
  AOI21_X1 U4311 ( .B1(n3510), .B2(n4508), .A(n3509), .ZN(n3511) );
  INV_X1 U4312 ( .A(n3511), .ZN(U3221) );
  NAND2_X1 U4313 ( .A1(n3513), .A2(n3847), .ZN(n3514) );
  XOR2_X1 U4314 ( .A(n3847), .B(n3515), .Z(n3521) );
  OAI22_X1 U4315 ( .A1(n3598), .A2(n4402), .B1(n3516), .B2(n4401), .ZN(n3519)
         );
  NOR2_X1 U4316 ( .A1(n4706), .A2(n3517), .ZN(n3518) );
  AOI211_X1 U4317 ( .C1(n4323), .C2(n3972), .A(n3519), .B(n3518), .ZN(n3520)
         );
  OAI21_X1 U4318 ( .B1(n3522), .B2(n3521), .A(n3520), .ZN(n4707) );
  NAND2_X1 U4319 ( .A1(n4707), .A2(n4646), .ZN(n3528) );
  AOI21_X1 U4320 ( .B1(n3524), .B2(n3531), .A(n2277), .ZN(n4709) );
  OAI22_X1 U4321 ( .A1(n4646), .A2(n2615), .B1(n3525), .B2(n4643), .ZN(n3526)
         );
  AOI21_X1 U4322 ( .B1(n4709), .B2(n4657), .A(n3526), .ZN(n3527) );
  OAI211_X1 U4323 ( .C1(n4706), .C2(n3529), .A(n3528), .B(n3527), .ZN(U3279)
         );
  INV_X1 U4324 ( .A(n3530), .ZN(n3532) );
  OAI21_X1 U4325 ( .B1(n3532), .B2(n3536), .A(n3531), .ZN(n4637) );
  AND2_X1 U4326 ( .A1(n3912), .A2(n3917), .ZN(n3843) );
  INV_X1 U4327 ( .A(n3843), .ZN(n3533) );
  XNOR2_X1 U4328 ( .A(n3534), .B(n3533), .ZN(n4639) );
  NAND2_X1 U4329 ( .A1(n4639), .A2(n3561), .ZN(n3542) );
  XNOR2_X1 U4330 ( .A(n3535), .B(n3843), .ZN(n3540) );
  NOR2_X1 U4331 ( .A1(n3536), .A2(n4401), .ZN(n3537) );
  AOI21_X1 U4332 ( .B1(n3973), .B2(n4323), .A(n3537), .ZN(n3538) );
  OAI21_X1 U4333 ( .B1(n4408), .B2(n4402), .A(n3538), .ZN(n3539) );
  AOI21_X1 U4334 ( .B1(n3540), .B2(n4289), .A(n3539), .ZN(n3541) );
  NAND2_X1 U4335 ( .A1(n4639), .A2(n4697), .ZN(n3543) );
  INV_X1 U4336 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3544) );
  MUX2_X1 U4337 ( .A(n3546), .B(n3544), .S(n4711), .Z(n3545) );
  OAI21_X1 U4338 ( .B1(n4637), .B2(n4478), .A(n3545), .ZN(U3487) );
  INV_X1 U4339 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3547) );
  MUX2_X1 U4340 ( .A(n3547), .B(n3546), .S(n4722), .Z(n3548) );
  OAI21_X1 U4341 ( .B1(n4637), .B2(n4414), .A(n3548), .ZN(U3528) );
  XNOR2_X1 U4342 ( .A(n3551), .B(n3550), .ZN(n3552) );
  XNOR2_X1 U4343 ( .A(n3549), .B(n3552), .ZN(n3556) );
  NOR2_X1 U4344 ( .A1(STATE_REG_SCAN_IN), .A2(n2638), .ZN(n4580) );
  AOI21_X1 U4345 ( .B1(n3970), .B2(n3786), .A(n4580), .ZN(n3554) );
  AOI22_X1 U4346 ( .A1(n3968), .A2(n4503), .B1(n3595), .B2(n3785), .ZN(n3553)
         );
  OAI211_X1 U4347 ( .C1(n4513), .C2(n3602), .A(n3554), .B(n3553), .ZN(n3555)
         );
  AOI21_X1 U4348 ( .B1(n3556), .B2(n4508), .A(n3555), .ZN(n3557) );
  INV_X1 U4349 ( .A(n3557), .ZN(U3231) );
  OAI21_X1 U4350 ( .B1(n3559), .B2(n3868), .A(n3558), .ZN(n4394) );
  OAI21_X1 U4351 ( .B1(n2325), .B2(n3800), .A(n3569), .ZN(n3560) );
  AOI22_X1 U4352 ( .A1(n4394), .A2(n3561), .B1(n4289), .B2(n3560), .ZN(n4391)
         );
  OAI21_X1 U4353 ( .B1(n2276), .B2(n3562), .A(n3574), .ZN(n4474) );
  OAI22_X1 U4354 ( .A1(n4646), .A2(n3563), .B1(n3668), .B2(n4643), .ZN(n3565)
         );
  OAI22_X1 U4355 ( .A1(n4210), .A2(n4403), .B1(n4498), .B2(n4081), .ZN(n3564)
         );
  AOI211_X1 U4356 ( .C1(n4387), .C2(n4206), .A(n3565), .B(n3564), .ZN(n3566)
         );
  OAI21_X1 U4357 ( .B1(n4474), .B2(n4233), .A(n3566), .ZN(n3567) );
  AOI21_X1 U4358 ( .B1(n4394), .B2(n4658), .A(n3567), .ZN(n3568) );
  OAI21_X1 U4359 ( .B1(n4391), .B2(n4663), .A(n3568), .ZN(U3276) );
  NAND2_X1 U4360 ( .A1(n3569), .A2(n3796), .ZN(n3571) );
  INV_X1 U4361 ( .A(n3867), .ZN(n3570) );
  XNOR2_X1 U4362 ( .A(n3571), .B(n3570), .ZN(n3572) );
  NAND2_X1 U4363 ( .A1(n3572), .A2(n4289), .ZN(n4381) );
  XNOR2_X1 U4364 ( .A(n3573), .B(n3867), .ZN(n4384) );
  NAND2_X1 U4365 ( .A1(n4384), .A2(n4264), .ZN(n3584) );
  INV_X1 U4366 ( .A(n3574), .ZN(n3576) );
  INV_X1 U4367 ( .A(n4282), .ZN(n3575) );
  OAI21_X1 U4368 ( .B1(n3576), .B2(n3580), .A(n3575), .ZN(n4470) );
  INV_X1 U4369 ( .A(n4470), .ZN(n3582) );
  AOI22_X1 U4370 ( .A1(n4267), .A2(n3968), .B1(n4379), .B2(n4266), .ZN(n3579)
         );
  INV_X1 U4371 ( .A(n3789), .ZN(n3577) );
  INV_X1 U4372 ( .A(n4643), .ZN(n4655) );
  AOI22_X1 U4373 ( .A1(n4663), .A2(REG2_REG_15__SCAN_IN), .B1(n3577), .B2(
        n4655), .ZN(n3578) );
  OAI211_X1 U4374 ( .C1(n3580), .C2(n4272), .A(n3579), .B(n3578), .ZN(n3581)
         );
  AOI21_X1 U4375 ( .B1(n3582), .B2(n4657), .A(n3581), .ZN(n3583) );
  OAI211_X1 U4376 ( .C1(n4663), .C2(n4381), .A(n3584), .B(n3583), .ZN(U3275)
         );
  INV_X1 U4377 ( .A(n3585), .ZN(n3586) );
  NOR2_X1 U4378 ( .A1(n3587), .A2(n3586), .ZN(n3841) );
  XOR2_X1 U4379 ( .A(n3841), .B(n3588), .Z(n4398) );
  INV_X1 U4380 ( .A(n4398), .ZN(n3607) );
  INV_X1 U4381 ( .A(n3589), .ZN(n3590) );
  NOR2_X1 U4382 ( .A1(n3591), .A2(n3590), .ZN(n3619) );
  INV_X1 U4383 ( .A(n3608), .ZN(n3592) );
  AOI21_X1 U4384 ( .B1(n3619), .B2(n3609), .A(n3592), .ZN(n3593) );
  XNOR2_X1 U4385 ( .A(n3593), .B(n3841), .ZN(n3594) );
  NAND2_X1 U4386 ( .A1(n3594), .A2(n4289), .ZN(n3597) );
  AOI22_X1 U4387 ( .A1(n3968), .A2(n4388), .B1(n4386), .B2(n3595), .ZN(n3596)
         );
  OAI211_X1 U4388 ( .C1(n3598), .C2(n4407), .A(n3597), .B(n3596), .ZN(n4397)
         );
  OR2_X1 U4389 ( .A1(n3611), .A2(n3599), .ZN(n3600) );
  NAND2_X1 U4390 ( .A1(n3601), .A2(n3600), .ZN(n4479) );
  NOR2_X1 U4391 ( .A1(n4479), .A2(n4233), .ZN(n3605) );
  OAI22_X1 U4392 ( .A1(n4646), .A2(n3603), .B1(n3602), .B2(n4643), .ZN(n3604)
         );
  AOI211_X1 U4393 ( .C1(n4397), .C2(n4646), .A(n3605), .B(n3604), .ZN(n3606)
         );
  OAI21_X1 U4394 ( .B1(n3607), .B2(n4295), .A(n3606), .ZN(U3277) );
  AND2_X1 U4395 ( .A1(n3609), .A2(n3608), .ZN(n3844) );
  XOR2_X1 U4396 ( .A(n3844), .B(n3610), .Z(n4410) );
  INV_X1 U4397 ( .A(n3611), .ZN(n3612) );
  OAI21_X1 U4398 ( .B1(n2277), .B2(n4400), .A(n3612), .ZN(n4483) );
  OAI22_X1 U4399 ( .A1(n4646), .A2(n3614), .B1(n3613), .B2(n4643), .ZN(n3616)
         );
  OAI22_X1 U4400 ( .A1(n4210), .A2(n4408), .B1(n4403), .B2(n4081), .ZN(n3615)
         );
  AOI211_X1 U4401 ( .C1(n3617), .C2(n4206), .A(n3616), .B(n3615), .ZN(n3618)
         );
  OAI21_X1 U4402 ( .B1(n4483), .B2(n4233), .A(n3618), .ZN(n3622) );
  XOR2_X1 U4403 ( .A(n3844), .B(n3619), .Z(n3620) );
  NAND2_X1 U4404 ( .A1(n3620), .A2(n4289), .ZN(n4406) );
  NOR2_X1 U4405 ( .A1(n4406), .A2(n4663), .ZN(n3621) );
  AOI211_X1 U4406 ( .C1(n4264), .C2(n4410), .A(n3622), .B(n3621), .ZN(n3623)
         );
  INV_X1 U4407 ( .A(n3623), .ZN(U3278) );
  AOI21_X1 U4408 ( .B1(n3624), .B2(n3625), .A(n3781), .ZN(n3626) );
  OR2_X1 U4409 ( .A1(n3624), .A2(n3625), .ZN(n3709) );
  NAND2_X1 U4410 ( .A1(n3626), .A2(n3709), .ZN(n3632) );
  OAI22_X1 U4411 ( .A1(n4500), .A2(n3628), .B1(n3627), .B2(n4497), .ZN(n3629)
         );
  AOI211_X1 U4412 ( .C1(n4503), .C2(n3977), .A(n3630), .B(n3629), .ZN(n3631)
         );
  OAI211_X1 U4413 ( .C1(n4513), .C2(n3633), .A(n3632), .B(n3631), .ZN(U3227)
         );
  XNOR2_X1 U4414 ( .A(n3635), .B(n3634), .ZN(n3636) );
  NAND2_X1 U4415 ( .A1(n3636), .A2(n4508), .ZN(n3641) );
  NOR2_X1 U4416 ( .A1(n4077), .A2(n4513), .ZN(n3639) );
  AOI22_X1 U4417 ( .A1(n4306), .A2(n3786), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3637) );
  OAI21_X1 U4418 ( .B1(n4500), .B2(n4075), .A(n3637), .ZN(n3638) );
  AOI211_X1 U4419 ( .C1(n4503), .C2(n3966), .A(n3639), .B(n3638), .ZN(n3640)
         );
  NAND2_X1 U4420 ( .A1(n3641), .A2(n3640), .ZN(U3211) );
  INV_X1 U4421 ( .A(n3642), .ZN(n3646) );
  INV_X1 U4422 ( .A(IR_REG_30__SCAN_IN), .ZN(n3643) );
  NAND3_X1 U4423 ( .A1(n3643), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3645) );
  INV_X1 U4424 ( .A(DATAI_31_), .ZN(n3644) );
  OAI22_X1 U4425 ( .A1(n3646), .A2(n3645), .B1(STATE_REG_SCAN_IN), .B2(n3644), 
        .ZN(U3321) );
  INV_X1 U4426 ( .A(n3647), .ZN(n3657) );
  OAI22_X1 U4427 ( .A1(n3649), .A2(n4643), .B1(n3648), .B2(n4646), .ZN(n3652)
         );
  OAI22_X1 U4428 ( .A1(n4092), .A2(n4210), .B1(n3650), .B2(n4081), .ZN(n3651)
         );
  AOI211_X1 U4429 ( .C1(n3653), .C2(n4206), .A(n3652), .B(n3651), .ZN(n3654)
         );
  OAI21_X1 U4430 ( .B1(n3655), .B2(n4233), .A(n3654), .ZN(n3656) );
  AOI21_X1 U4431 ( .B1(n3657), .B2(n4646), .A(n3656), .ZN(n3658) );
  OAI21_X1 U4432 ( .B1(n3659), .B2(n4295), .A(n3658), .ZN(U3262) );
  INV_X1 U4433 ( .A(n3661), .ZN(n3663) );
  NAND2_X1 U4434 ( .A1(n3663), .A2(n3662), .ZN(n3664) );
  XNOR2_X1 U4435 ( .A(n3660), .B(n3664), .ZN(n3670) );
  NAND2_X1 U4436 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4586) );
  OAI21_X1 U4437 ( .B1(n4498), .B2(n3777), .A(n4586), .ZN(n3665) );
  INV_X1 U4438 ( .A(n3665), .ZN(n3667) );
  AOI22_X1 U4439 ( .A1(n3969), .A2(n3786), .B1(n4387), .B2(n3785), .ZN(n3666)
         );
  OAI211_X1 U4440 ( .C1(n4513), .C2(n3668), .A(n3667), .B(n3666), .ZN(n3669)
         );
  AOI21_X1 U4441 ( .B1(n3670), .B2(n4508), .A(n3669), .ZN(n3671) );
  INV_X1 U4442 ( .A(n3671), .ZN(U3212) );
  INV_X1 U4443 ( .A(n3672), .ZN(n3676) );
  OAI21_X1 U4444 ( .B1(n3746), .B2(n3674), .A(n3673), .ZN(n3675) );
  NAND3_X1 U4445 ( .A1(n3676), .A2(n4508), .A3(n3675), .ZN(n3681) );
  OAI22_X1 U4446 ( .A1(n4157), .A2(n3777), .B1(n4500), .B2(n4159), .ZN(n3679)
         );
  INV_X1 U4447 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4864) );
  OAI22_X1 U4448 ( .A1(n3677), .A2(n4497), .B1(STATE_REG_SCAN_IN), .B2(n4864), 
        .ZN(n3678) );
  NOR2_X1 U4449 ( .A1(n3679), .A2(n3678), .ZN(n3680) );
  OAI211_X1 U4450 ( .C1(n4513), .C2(n4161), .A(n3681), .B(n3680), .ZN(U3213)
         );
  XNOR2_X1 U4451 ( .A(n3683), .B(n3682), .ZN(n3684) );
  NAND2_X1 U4452 ( .A1(n3684), .A2(n4508), .ZN(n3687) );
  INV_X1 U4453 ( .A(REG3_REG_19__SCAN_IN), .ZN(n5043) );
  NOR2_X1 U4454 ( .A1(n5043), .A2(STATE_REG_SCAN_IN), .ZN(n4055) );
  OAI22_X1 U4455 ( .A1(n4500), .A2(n4231), .B1(n4345), .B2(n3777), .ZN(n3685)
         );
  AOI211_X1 U4456 ( .C1(n3786), .C2(n4366), .A(n4055), .B(n3685), .ZN(n3686)
         );
  OAI211_X1 U4457 ( .C1(n4513), .C2(n4234), .A(n3687), .B(n3686), .ZN(U3216)
         );
  AOI21_X1 U4458 ( .B1(n3739), .B2(n3737), .A(n3736), .ZN(n3691) );
  XOR2_X1 U4459 ( .A(n3689), .B(n3688), .Z(n3690) );
  XNOR2_X1 U4460 ( .A(n3691), .B(n3690), .ZN(n3697) );
  AOI22_X1 U4461 ( .A1(n4342), .A2(n4503), .B1(n4341), .B2(n3785), .ZN(n3695)
         );
  NOR2_X1 U4462 ( .A1(n3692), .A2(STATE_REG_SCAN_IN), .ZN(n3693) );
  AOI21_X1 U4463 ( .B1(n3786), .B2(n4225), .A(n3693), .ZN(n3694) );
  OAI211_X1 U4464 ( .C1(n4513), .C2(n4186), .A(n3695), .B(n3694), .ZN(n3696)
         );
  AOI21_X1 U4465 ( .B1(n3697), .B2(n4508), .A(n3696), .ZN(n3698) );
  INV_X1 U4466 ( .A(n3698), .ZN(U3220) );
  NAND2_X1 U4467 ( .A1(n3700), .A2(n3699), .ZN(n3702) );
  XOR2_X1 U4468 ( .A(n3702), .B(n3701), .Z(n3707) );
  OAI22_X1 U4469 ( .A1(n4157), .A2(n4497), .B1(STATE_REG_SCAN_IN), .B2(n3703), 
        .ZN(n3705) );
  OAI22_X1 U4470 ( .A1(n4111), .A2(n3777), .B1(n4500), .B2(n4113), .ZN(n3704)
         );
  AOI211_X1 U4471 ( .C1(n4114), .C2(n3779), .A(n3705), .B(n3704), .ZN(n3706)
         );
  OAI21_X1 U4472 ( .B1(n3707), .B2(n3781), .A(n3706), .ZN(U3222) );
  NAND2_X1 U4473 ( .A1(n3709), .A2(n3708), .ZN(n3712) );
  NAND2_X1 U4474 ( .A1(n3712), .A2(n3710), .ZN(n3711) );
  OAI211_X1 U4475 ( .C1(n3712), .C2(n3710), .A(n3711), .B(n4508), .ZN(n3719)
         );
  AOI21_X1 U4476 ( .B1(n2540), .B2(n3786), .A(n3713), .ZN(n3718) );
  AOI22_X1 U4477 ( .A1(n4503), .A2(n3976), .B1(n3785), .B2(n3714), .ZN(n3717)
         );
  OR2_X1 U4478 ( .A1(n4513), .A2(n3715), .ZN(n3716) );
  NAND4_X1 U4479 ( .A1(n3719), .A2(n3718), .A3(n3717), .A4(n3716), .ZN(U3224)
         );
  NAND2_X1 U4480 ( .A1(n2268), .A2(n3720), .ZN(n3721) );
  XNOR2_X1 U4481 ( .A(n3722), .B(n3721), .ZN(n3726) );
  AND2_X1 U4482 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4617) );
  AOI21_X1 U4483 ( .B1(n4379), .B2(n3786), .A(n4617), .ZN(n3724) );
  AOI22_X1 U4484 ( .A1(n4366), .A2(n4503), .B1(n4365), .B2(n3785), .ZN(n3723)
         );
  OAI211_X1 U4485 ( .C1(n4513), .C2(n4268), .A(n3724), .B(n3723), .ZN(n3725)
         );
  AOI21_X1 U4486 ( .B1(n3726), .B2(n4508), .A(n3725), .ZN(n3727) );
  INV_X1 U4487 ( .A(n3727), .ZN(U3225) );
  NAND2_X1 U4488 ( .A1(n2237), .A2(n3728), .ZN(n3730) );
  XNOR2_X1 U4489 ( .A(n3730), .B(n3729), .ZN(n3735) );
  NAND2_X1 U4490 ( .A1(n4136), .A2(n4503), .ZN(n3732) );
  AOI22_X1 U4491 ( .A1(n4324), .A2(n3786), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3731) );
  OAI211_X1 U4492 ( .C1(n4500), .C2(n4134), .A(n3732), .B(n3731), .ZN(n3733)
         );
  AOI21_X1 U4493 ( .B1(n4131), .B2(n3779), .A(n3733), .ZN(n3734) );
  OAI21_X1 U4494 ( .B1(n3735), .B2(n3781), .A(n3734), .ZN(U3226) );
  NAND2_X1 U4495 ( .A1(n2416), .A2(n3737), .ZN(n3738) );
  XNOR2_X1 U4496 ( .A(n3739), .B(n3738), .ZN(n3744) );
  INV_X1 U4497 ( .A(n4207), .ZN(n3742) );
  AOI22_X1 U4498 ( .A1(n3786), .A2(n4249), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n3741) );
  AOI22_X1 U4499 ( .A1(n4351), .A2(n4503), .B1(n3785), .B2(n4350), .ZN(n3740)
         );
  OAI211_X1 U4500 ( .C1(n4513), .C2(n3742), .A(n3741), .B(n3740), .ZN(n3743)
         );
  AOI21_X1 U4501 ( .B1(n3744), .B2(n4508), .A(n3743), .ZN(n3745) );
  INV_X1 U4502 ( .A(n3745), .ZN(U3230) );
  AOI21_X1 U4503 ( .B1(n3748), .B2(n3747), .A(n3746), .ZN(n3756) );
  INV_X1 U4504 ( .A(n3749), .ZN(n4177) );
  OAI22_X1 U4505 ( .A1(n4497), .A2(n3751), .B1(STATE_REG_SCAN_IN), .B2(n3750), 
        .ZN(n3754) );
  OAI22_X1 U4506 ( .A1(n4173), .A2(n3777), .B1(n4500), .B2(n3752), .ZN(n3753)
         );
  AOI211_X1 U4507 ( .C1(n4177), .C2(n3779), .A(n3754), .B(n3753), .ZN(n3755)
         );
  OAI21_X1 U4508 ( .B1(n3756), .B2(n3781), .A(n3755), .ZN(U3232) );
  INV_X1 U4509 ( .A(n3757), .ZN(n3762) );
  AOI21_X1 U4510 ( .B1(n3759), .B2(n3761), .A(n3758), .ZN(n3760) );
  AOI21_X1 U4511 ( .B1(n3762), .B2(n3761), .A(n3760), .ZN(n3768) );
  OAI22_X1 U4512 ( .A1(n4286), .A2(n4497), .B1(STATE_REG_SCAN_IN), .B2(n4623), 
        .ZN(n3763) );
  INV_X1 U4513 ( .A(n3763), .ZN(n3765) );
  AOI22_X1 U4514 ( .A1(n4503), .A2(n4249), .B1(n3785), .B2(n4248), .ZN(n3764)
         );
  OAI211_X1 U4515 ( .C1(n4513), .C2(n4254), .A(n3765), .B(n3764), .ZN(n3766)
         );
  INV_X1 U4516 ( .A(n3766), .ZN(n3767) );
  OAI21_X1 U4517 ( .B1(n3768), .B2(n3781), .A(n3767), .ZN(U3235) );
  INV_X1 U4518 ( .A(n3770), .ZN(n3771) );
  NOR2_X1 U4519 ( .A1(n3772), .A2(n3771), .ZN(n3773) );
  XNOR2_X1 U4520 ( .A(n3769), .B(n3773), .ZN(n3782) );
  AOI22_X1 U4521 ( .A1(n3785), .A2(n3774), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3776) );
  NAND2_X1 U4522 ( .A1(n4136), .A2(n3786), .ZN(n3775) );
  OAI211_X1 U4523 ( .C1(n4092), .C2(n3777), .A(n3776), .B(n3775), .ZN(n3778)
         );
  AOI21_X1 U4524 ( .B1(n4099), .B2(n3779), .A(n3778), .ZN(n3780) );
  OAI21_X1 U4525 ( .B1(n3782), .B2(n3781), .A(n3780), .ZN(U3237) );
  NAND2_X1 U4526 ( .A1(n2391), .A2(n4504), .ZN(n3784) );
  XNOR2_X1 U4527 ( .A(n3784), .B(n4505), .ZN(n3791) );
  AND2_X1 U4528 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4599) );
  AOI21_X1 U4529 ( .B1(n4379), .B2(n4503), .A(n4599), .ZN(n3788) );
  AOI22_X1 U4530 ( .A1(n3968), .A2(n3786), .B1(n4378), .B2(n3785), .ZN(n3787)
         );
  OAI211_X1 U4531 ( .C1(n4513), .C2(n3789), .A(n3788), .B(n3787), .ZN(n3790)
         );
  AOI21_X1 U4532 ( .B1(n3791), .B2(n4508), .A(n3790), .ZN(n3792) );
  INV_X1 U4533 ( .A(n3792), .ZN(U3238) );
  NAND2_X1 U4534 ( .A1(n2777), .A2(DATAI_31_), .ZN(n4064) );
  INV_X1 U4535 ( .A(n4064), .ZN(n3828) );
  INV_X1 U4536 ( .A(n3964), .ZN(n3793) );
  NAND2_X1 U4537 ( .A1(n2777), .A2(DATAI_30_), .ZN(n3811) );
  NOR2_X1 U4538 ( .A1(n3793), .A2(n4302), .ZN(n3860) );
  INV_X1 U4539 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4065) );
  NAND2_X1 U4540 ( .A1(n2625), .A2(REG1_REG_31__SCAN_IN), .ZN(n3795) );
  NAND2_X1 U4541 ( .A1(n2735), .A2(REG0_REG_31__SCAN_IN), .ZN(n3794) );
  OAI211_X1 U4542 ( .C1(n2544), .C2(n4065), .A(n3795), .B(n3794), .ZN(n4063)
         );
  NOR2_X1 U4543 ( .A1(n4063), .A2(n4064), .ZN(n3859) );
  AND2_X1 U4544 ( .A1(n2288), .A2(n3858), .ZN(n3941) );
  INV_X1 U4545 ( .A(n3941), .ZN(n3810) );
  NAND2_X1 U4546 ( .A1(n3796), .A2(n3799), .ZN(n3923) );
  NAND2_X1 U4547 ( .A1(n3798), .A2(n3797), .ZN(n3904) );
  NAND2_X1 U4548 ( .A1(n3904), .A2(n3799), .ZN(n3922) );
  OAI21_X1 U4549 ( .B1(n3800), .B2(n3923), .A(n3922), .ZN(n3802) );
  INV_X1 U4550 ( .A(n3801), .ZN(n3925) );
  AOI21_X1 U4551 ( .B1(n3802), .B2(n3928), .A(n3925), .ZN(n3805) );
  INV_X1 U4552 ( .A(n4147), .ZN(n3804) );
  OAI21_X1 U4553 ( .B1(n3805), .B2(n3804), .A(n3803), .ZN(n3806) );
  INV_X1 U4554 ( .A(n3806), .ZN(n3808) );
  OAI21_X1 U4555 ( .B1(n3808), .B2(n3935), .A(n3807), .ZN(n3809) );
  OAI221_X1 U4556 ( .B1(n3810), .B2(n3937), .C1(n3810), .C2(n3809), .A(n3945), 
        .ZN(n3814) );
  OR2_X1 U4557 ( .A1(n3965), .A2(n3816), .ZN(n3813) );
  OR2_X1 U4558 ( .A1(n3964), .A2(n3811), .ZN(n3812) );
  NAND2_X1 U4559 ( .A1(n4063), .A2(n4064), .ZN(n3949) );
  AND2_X1 U4560 ( .A1(n3812), .A2(n3949), .ZN(n3864) );
  NAND2_X1 U4561 ( .A1(n3813), .A2(n3864), .ZN(n3820) );
  OR4_X1 U4562 ( .A1(n3814), .A2(n3819), .A3(n3818), .A4(n3820), .ZN(n3826) );
  INV_X1 U4563 ( .A(n4071), .ZN(n3823) );
  AOI21_X1 U4564 ( .B1(n3965), .B2(n3816), .A(n3815), .ZN(n3821) );
  NAND2_X1 U4565 ( .A1(n3821), .A2(n3817), .ZN(n3942) );
  OR2_X1 U4566 ( .A1(n3819), .A2(n3818), .ZN(n3822) );
  AOI21_X1 U4567 ( .B1(n3822), .B2(n3821), .A(n3820), .ZN(n3946) );
  OAI21_X1 U4568 ( .B1(n3823), .B2(n3942), .A(n3946), .ZN(n3825) );
  INV_X1 U4569 ( .A(n4063), .ZN(n3824) );
  AOI22_X1 U4570 ( .A1(n3826), .A2(n3825), .B1(n3824), .B2(n4302), .ZN(n3827)
         );
  AOI211_X1 U4571 ( .C1(n3828), .C2(n3860), .A(n3859), .B(n3827), .ZN(n3956)
         );
  XNOR2_X1 U4572 ( .A(n4249), .B(n4224), .ZN(n4222) );
  NOR4_X1 U4573 ( .A1(n4168), .A2(n3830), .A3(n4284), .A4(n3829), .ZN(n3831)
         );
  AND3_X1 U4574 ( .A1(n4071), .A2(n4222), .A3(n3831), .ZN(n3836) );
  INV_X1 U4575 ( .A(n3832), .ZN(n3835) );
  NOR2_X1 U4576 ( .A1(n3834), .A2(n3833), .ZN(n4089) );
  XNOR2_X1 U4577 ( .A(n4324), .B(n4154), .ZN(n4151) );
  NAND4_X1 U4578 ( .A1(n3836), .A2(n3835), .A3(n4089), .A4(n4151), .ZN(n3875)
         );
  OR2_X1 U4579 ( .A1(n3838), .A2(n3837), .ZN(n4119) );
  INV_X1 U4580 ( .A(n4119), .ZN(n4124) );
  NAND2_X1 U4581 ( .A1(n3840), .A2(n3839), .ZN(n4201) );
  NAND3_X1 U4582 ( .A1(n4124), .A2(n3841), .A3(n4201), .ZN(n3855) );
  AND2_X1 U4583 ( .A1(n4216), .A2(n4142), .ZN(n4262) );
  NAND4_X1 U4584 ( .A1(n4262), .A2(n3844), .A3(n3843), .A4(n3842), .ZN(n3854)
         );
  NAND4_X1 U4585 ( .A1(n2334), .A2(n3847), .A3(n3846), .A4(n3845), .ZN(n3853)
         );
  INV_X1 U4586 ( .A(n3933), .ZN(n3848) );
  INV_X1 U4587 ( .A(n2823), .ZN(n3850) );
  NAND4_X1 U4588 ( .A1(n4184), .A2(n3851), .A3(n3850), .A4(n3849), .ZN(n3852)
         );
  NOR4_X1 U4589 ( .A1(n3855), .A2(n3854), .A3(n3853), .A4(n3852), .ZN(n3872)
         );
  INV_X1 U4590 ( .A(n3857), .ZN(n4087) );
  NAND2_X1 U4591 ( .A1(n4087), .A2(n3858), .ZN(n4105) );
  INV_X1 U4592 ( .A(n4105), .ZN(n3871) );
  INV_X1 U4593 ( .A(n3859), .ZN(n3862) );
  INV_X1 U4594 ( .A(n3860), .ZN(n3861) );
  NAND2_X1 U4595 ( .A1(n3862), .A2(n3861), .ZN(n3950) );
  INV_X1 U4596 ( .A(n3950), .ZN(n3863) );
  NAND3_X1 U4597 ( .A1(n3865), .A2(n3864), .A3(n3863), .ZN(n3869) );
  NOR4_X1 U4598 ( .A1(n3869), .A2(n3868), .A3(n3867), .A4(n3866), .ZN(n3870)
         );
  NAND4_X1 U4599 ( .A1(n3872), .A2(n2293), .A3(n3871), .A4(n3870), .ZN(n3874)
         );
  OAI21_X1 U4600 ( .B1(n3875), .B2(n3874), .A(n3873), .ZN(n3953) );
  INV_X1 U4601 ( .A(n3876), .ZN(n3878) );
  OAI211_X1 U4602 ( .C1(n3880), .C2(n3879), .A(n3878), .B(n3877), .ZN(n3883)
         );
  NAND3_X1 U4603 ( .A1(n3883), .A2(n3882), .A3(n3881), .ZN(n3886) );
  NAND3_X1 U4604 ( .A1(n3886), .A2(n3885), .A3(n3884), .ZN(n3889) );
  NAND3_X1 U4605 ( .A1(n3889), .A2(n3888), .A3(n3887), .ZN(n3898) );
  INV_X1 U4606 ( .A(n3890), .ZN(n3911) );
  INV_X1 U4607 ( .A(n3891), .ZN(n3893) );
  NOR3_X1 U4608 ( .A1(n3911), .A2(n3893), .A3(n3892), .ZN(n3897) );
  INV_X1 U4609 ( .A(n3894), .ZN(n3895) );
  AOI211_X1 U4610 ( .C1(n3898), .C2(n3897), .A(n3896), .B(n3895), .ZN(n3903)
         );
  NAND2_X1 U4611 ( .A1(n3900), .A2(n3899), .ZN(n3910) );
  OAI211_X1 U4612 ( .C1(n3903), .C2(n3910), .A(n3902), .B(n3901), .ZN(n3907)
         );
  INV_X1 U4613 ( .A(n3904), .ZN(n3906) );
  NAND3_X1 U4614 ( .A1(n3907), .A2(n3906), .A3(n3905), .ZN(n3916) );
  NOR4_X1 U4615 ( .A1(n3911), .A2(n3910), .A3(n3909), .A4(n3908), .ZN(n3914)
         );
  INV_X1 U4616 ( .A(n3912), .ZN(n3913) );
  OAI21_X1 U4617 ( .B1(n3914), .B2(n3913), .A(n3922), .ZN(n3915) );
  NAND2_X1 U4618 ( .A1(n3916), .A2(n3915), .ZN(n3920) );
  NAND4_X1 U4619 ( .A1(n3920), .A2(n3919), .A3(n3918), .A4(n3917), .ZN(n3927)
         );
  INV_X1 U4620 ( .A(n3921), .ZN(n3924) );
  OAI21_X1 U4621 ( .B1(n3924), .B2(n3923), .A(n3922), .ZN(n3926) );
  AOI21_X1 U4622 ( .B1(n3927), .B2(n3926), .A(n3925), .ZN(n3932) );
  INV_X1 U4623 ( .A(n3928), .ZN(n3931) );
  INV_X1 U4624 ( .A(n3929), .ZN(n3930) );
  OAI21_X1 U4625 ( .B1(n3932), .B2(n3931), .A(n3930), .ZN(n3934) );
  AOI211_X1 U4626 ( .C1(n3934), .C2(n4147), .A(n3933), .B(n4146), .ZN(n3936)
         );
  NOR2_X1 U4627 ( .A1(n3936), .A2(n3935), .ZN(n3939) );
  OAI21_X1 U4628 ( .B1(n3939), .B2(n3938), .A(n3937), .ZN(n3940) );
  NAND2_X1 U4629 ( .A1(n3941), .A2(n3940), .ZN(n3944) );
  AOI211_X1 U4630 ( .C1(n3945), .C2(n3944), .A(n3943), .B(n3942), .ZN(n3948)
         );
  INV_X1 U4631 ( .A(n3946), .ZN(n3947) );
  NOR2_X1 U4632 ( .A1(n3948), .A2(n3947), .ZN(n3951) );
  OAI21_X1 U4633 ( .B1(n3951), .B2(n3950), .A(n3949), .ZN(n3952) );
  MUX2_X1 U4634 ( .A(n3953), .B(n3952), .S(n2808), .Z(n3954) );
  OAI21_X1 U4635 ( .B1(n3956), .B2(n3955), .A(n3954), .ZN(n3957) );
  XNOR2_X1 U4636 ( .A(n3957), .B(n4057), .ZN(n3963) );
  NAND2_X1 U4637 ( .A1(n3959), .A2(n3958), .ZN(n3960) );
  OAI211_X1 U4638 ( .C1(n4487), .C2(n3962), .A(n3960), .B(B_REG_SCAN_IN), .ZN(
        n3961) );
  OAI21_X1 U4639 ( .B1(n3963), .B2(n3962), .A(n3961), .ZN(U3239) );
  MUX2_X1 U4640 ( .A(n4063), .B(DATAO_REG_31__SCAN_IN), .S(n3979), .Z(U3581)
         );
  MUX2_X1 U4641 ( .A(n3964), .B(DATAO_REG_30__SCAN_IN), .S(n3979), .Z(U3580)
         );
  MUX2_X1 U4642 ( .A(n3965), .B(DATAO_REG_29__SCAN_IN), .S(n3979), .Z(U3579)
         );
  MUX2_X1 U4643 ( .A(n3966), .B(DATAO_REG_28__SCAN_IN), .S(n3979), .Z(U3578)
         );
  MUX2_X1 U4644 ( .A(DATAO_REG_27__SCAN_IN), .B(n3967), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4645 ( .A(n4306), .B(DATAO_REG_26__SCAN_IN), .S(n3979), .Z(U3576)
         );
  MUX2_X1 U4646 ( .A(DATAO_REG_25__SCAN_IN), .B(n4136), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4647 ( .A(n4108), .B(DATAO_REG_24__SCAN_IN), .S(n3979), .Z(U3574)
         );
  MUX2_X1 U4648 ( .A(n4324), .B(DATAO_REG_23__SCAN_IN), .S(n3979), .Z(U3573)
         );
  MUX2_X1 U4649 ( .A(n4342), .B(DATAO_REG_22__SCAN_IN), .S(n3979), .Z(U3572)
         );
  MUX2_X1 U4650 ( .A(n4351), .B(DATAO_REG_21__SCAN_IN), .S(n3979), .Z(U3571)
         );
  MUX2_X1 U4651 ( .A(n4225), .B(DATAO_REG_20__SCAN_IN), .S(n3979), .Z(U3570)
         );
  MUX2_X1 U4652 ( .A(n4249), .B(DATAO_REG_19__SCAN_IN), .S(n3979), .Z(U3569)
         );
  MUX2_X1 U4653 ( .A(DATAO_REG_18__SCAN_IN), .B(n4366), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4654 ( .A(DATAO_REG_17__SCAN_IN), .B(n4502), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4655 ( .A(DATAO_REG_16__SCAN_IN), .B(n4379), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4656 ( .A(n4389), .B(DATAO_REG_15__SCAN_IN), .S(n3979), .Z(U3565)
         );
  MUX2_X1 U4657 ( .A(DATAO_REG_14__SCAN_IN), .B(n3968), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4658 ( .A(n3969), .B(DATAO_REG_13__SCAN_IN), .S(n3979), .Z(U3563)
         );
  MUX2_X1 U4659 ( .A(n3970), .B(DATAO_REG_12__SCAN_IN), .S(n3979), .Z(U3562)
         );
  MUX2_X1 U4660 ( .A(DATAO_REG_11__SCAN_IN), .B(n3971), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4661 ( .A(n3972), .B(DATAO_REG_10__SCAN_IN), .S(n3979), .Z(U3560)
         );
  MUX2_X1 U4662 ( .A(n3973), .B(DATAO_REG_9__SCAN_IN), .S(n3979), .Z(U3559) );
  MUX2_X1 U4663 ( .A(DATAO_REG_8__SCAN_IN), .B(n3974), .S(U4043), .Z(U3558) );
  MUX2_X1 U4664 ( .A(DATAO_REG_7__SCAN_IN), .B(n3975), .S(U4043), .Z(U3557) );
  MUX2_X1 U4665 ( .A(n3976), .B(DATAO_REG_6__SCAN_IN), .S(n3979), .Z(U3556) );
  MUX2_X1 U4666 ( .A(DATAO_REG_5__SCAN_IN), .B(n3977), .S(U4043), .Z(U3555) );
  MUX2_X1 U4667 ( .A(DATAO_REG_4__SCAN_IN), .B(n2540), .S(U4043), .Z(U3554) );
  MUX2_X1 U4668 ( .A(n2890), .B(DATAO_REG_3__SCAN_IN), .S(n3979), .Z(U3553) );
  MUX2_X1 U4669 ( .A(DATAO_REG_2__SCAN_IN), .B(n3978), .S(U4043), .Z(U3552) );
  MUX2_X1 U4670 ( .A(DATAO_REG_1__SCAN_IN), .B(n2510), .S(U4043), .Z(U3551) );
  MUX2_X1 U4671 ( .A(n3257), .B(DATAO_REG_0__SCAN_IN), .S(n3979), .Z(U3550) );
  OAI211_X1 U4672 ( .C1(n3982), .C2(n3981), .A(n4631), .B(n3980), .ZN(n3989)
         );
  OAI211_X1 U4673 ( .C1(n3140), .C2(n3985), .A(n4575), .B(n3984), .ZN(n3988)
         );
  AOI22_X1 U4674 ( .A1(n4629), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3986) );
  NAND4_X1 U4675 ( .A1(n3989), .A2(n3988), .A3(n3987), .A4(n3986), .ZN(U3241)
         );
  OAI211_X1 U4676 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3991), .A(n4631), .B(n3990), 
        .ZN(n3999) );
  NAND2_X1 U4677 ( .A1(n3992), .A2(n4493), .ZN(n3998) );
  AOI22_X1 U4678 ( .A1(n4629), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3997) );
  XNOR2_X1 U4679 ( .A(n3994), .B(n3993), .ZN(n3995) );
  NAND2_X1 U4680 ( .A1(n4575), .A2(n3995), .ZN(n3996) );
  NAND4_X1 U4681 ( .A1(n3999), .A2(n3998), .A3(n3997), .A4(n3996), .ZN(U3243)
         );
  MUX2_X1 U4682 ( .A(n4235), .B(REG2_REG_19__SCAN_IN), .S(n4057), .Z(n4020) );
  INV_X1 U4683 ( .A(n4021), .ZN(n4676) );
  AOI22_X1 U4684 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4676), .B1(n4021), .B2(
        n4255), .ZN(n4627) );
  NOR2_X1 U4685 ( .A1(n3603), .A2(n4681), .ZN(n4574) );
  NAND2_X1 U4686 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4026), .ZN(n4009) );
  INV_X1 U4687 ( .A(n4026), .ZN(n4682) );
  AOI22_X1 U4688 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4026), .B1(n4682), .B2(
        n2615), .ZN(n4559) );
  NAND2_X1 U4689 ( .A1(n4027), .A2(REG2_REG_9__SCAN_IN), .ZN(n4006) );
  INV_X1 U4690 ( .A(n4027), .ZN(n4684) );
  AOI22_X1 U4691 ( .A1(n4027), .A2(REG2_REG_9__SCAN_IN), .B1(n2588), .B2(n4684), .ZN(n4538) );
  NAND2_X1 U4692 ( .A1(n4031), .A2(n4004), .ZN(n4005) );
  NAND2_X1 U4693 ( .A1(n4005), .A2(n4524), .ZN(n4537) );
  NAND2_X1 U4694 ( .A1(n4544), .A2(n4007), .ZN(n4008) );
  NAND2_X1 U4695 ( .A1(n4008), .A2(n4545), .ZN(n4558) );
  NAND2_X1 U4696 ( .A1(n4036), .A2(n4010), .ZN(n4011) );
  NAND2_X1 U4697 ( .A1(n4011), .A2(n4567), .ZN(n4577) );
  OAI22_X1 U4698 ( .A1(n4574), .A2(n4577), .B1(REG2_REG_13__SCAN_IN), .B2(
        n4025), .ZN(n4012) );
  NOR2_X1 U4699 ( .A1(n2368), .A2(n4012), .ZN(n4013) );
  NAND2_X1 U4700 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4023), .ZN(n4014) );
  OAI21_X1 U4701 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4023), .A(n4014), .ZN(n4596) );
  INV_X1 U4702 ( .A(n4045), .ZN(n4678) );
  NAND2_X1 U4703 ( .A1(n4015), .A2(n4678), .ZN(n4016) );
  NAND2_X1 U4704 ( .A1(n4606), .A2(n4283), .ZN(n4605) );
  NAND2_X1 U4705 ( .A1(n4016), .A2(n4605), .ZN(n4613) );
  NOR2_X1 U4706 ( .A1(n4049), .A2(REG2_REG_17__SCAN_IN), .ZN(n4017) );
  AOI21_X1 U4707 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4049), .A(n4017), .ZN(n4615) );
  INV_X1 U4708 ( .A(n4017), .ZN(n4018) );
  AOI21_X1 U4709 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4021), .A(n4625), .ZN(n4019) );
  XOR2_X1 U4710 ( .A(n4020), .B(n4019), .Z(n4061) );
  INV_X1 U4711 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U4712 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4021), .B1(n4676), .B2(
        n4051), .ZN(n4633) );
  NOR2_X1 U4713 ( .A1(n4049), .A2(REG1_REG_17__SCAN_IN), .ZN(n4050) );
  NAND2_X1 U4714 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4023), .ZN(n4044) );
  INV_X1 U4715 ( .A(n4023), .ZN(n4679) );
  INV_X1 U4716 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U4717 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4023), .B1(n4679), .B2(
        n4022), .ZN(n4602) );
  NAND2_X1 U4718 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4025), .ZN(n4040) );
  INV_X1 U4719 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U4720 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4025), .B1(n4681), .B2(
        n4024), .ZN(n4583) );
  INV_X1 U4721 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4720) );
  AOI22_X1 U4722 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4026), .B1(n4682), .B2(
        n4720), .ZN(n4556) );
  NAND2_X1 U4723 ( .A1(n4027), .A2(REG1_REG_9__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U4724 ( .A1(n4027), .A2(REG1_REG_9__SCAN_IN), .B1(n3496), .B2(n4684), .ZN(n4535) );
  INV_X1 U4725 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4028) );
  NAND2_X1 U4726 ( .A1(n4031), .A2(n4030), .ZN(n4032) );
  NAND2_X1 U4727 ( .A1(REG1_REG_8__SCAN_IN), .A2(n4530), .ZN(n4529) );
  NAND2_X1 U4728 ( .A1(n4544), .A2(n4034), .ZN(n4035) );
  NAND2_X1 U4729 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4551), .ZN(n4550) );
  NAND2_X1 U4730 ( .A1(n4036), .A2(n4038), .ZN(n4039) );
  NAND2_X1 U4731 ( .A1(n4041), .A2(n4042), .ZN(n4043) );
  NAND2_X1 U4732 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4592), .ZN(n4591) );
  NAND2_X1 U4733 ( .A1(n4043), .A2(n4591), .ZN(n4601) );
  NAND2_X1 U4734 ( .A1(n4602), .A2(n4601), .ZN(n4600) );
  NAND2_X1 U4735 ( .A1(n4044), .A2(n4600), .ZN(n4046) );
  NOR2_X1 U4736 ( .A1(n4045), .A2(n4046), .ZN(n4047) );
  XNOR2_X1 U4737 ( .A(n4046), .B(n4045), .ZN(n4609) );
  NOR2_X1 U4738 ( .A1(REG1_REG_16__SCAN_IN), .A2(n4609), .ZN(n4610) );
  NOR2_X1 U4739 ( .A1(n4047), .A2(n4610), .ZN(n4619) );
  INV_X1 U4740 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U4741 ( .A1(n4049), .A2(n4048), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4677), .ZN(n4618) );
  INV_X1 U4742 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4052) );
  MUX2_X1 U4743 ( .A(REG1_REG_19__SCAN_IN), .B(n4052), .S(n4057), .Z(n4053) );
  XNOR2_X1 U4744 ( .A(n4054), .B(n4053), .ZN(n4059) );
  AOI21_X1 U4745 ( .B1(n4629), .B2(ADDR_REG_19__SCAN_IN), .A(n4055), .ZN(n4056) );
  OAI21_X1 U4746 ( .B1(n4057), .B2(n4635), .A(n4056), .ZN(n4058) );
  AOI21_X1 U4747 ( .B1(n4059), .B2(n4631), .A(n4058), .ZN(n4060) );
  OAI21_X1 U4748 ( .B1(n4061), .B2(n4624), .A(n4060), .ZN(U3259) );
  NOR2_X2 U4749 ( .A1(n4299), .A2(n4302), .ZN(n4298) );
  XNOR2_X1 U4750 ( .A(n4298), .B(n4064), .ZN(n4418) );
  NAND2_X1 U4751 ( .A1(n4063), .A2(n4062), .ZN(n4300) );
  OAI21_X1 U4752 ( .B1(n4064), .B2(n4401), .A(n4300), .ZN(n4415) );
  NOR2_X1 U4753 ( .A1(n4646), .A2(n4065), .ZN(n4066) );
  AOI21_X1 U4754 ( .B1(n4415), .B2(n4646), .A(n4066), .ZN(n4067) );
  OAI21_X1 U4755 ( .B1(n4418), .B2(n4233), .A(n4067), .ZN(U3260) );
  XNOR2_X1 U4756 ( .A(n4068), .B(n4071), .ZN(n4069) );
  NAND2_X1 U4757 ( .A1(n4069), .A2(n4289), .ZN(n4308) );
  XOR2_X1 U4758 ( .A(n4071), .B(n4070), .Z(n4311) );
  NAND2_X1 U4759 ( .A1(n4311), .A2(n4264), .ZN(n4085) );
  INV_X1 U4760 ( .A(n4072), .ZN(n4074) );
  NAND2_X1 U4761 ( .A1(n4096), .A2(n4305), .ZN(n4073) );
  NAND2_X1 U4762 ( .A1(n4074), .A2(n4073), .ZN(n4425) );
  INV_X1 U4763 ( .A(n4425), .ZN(n4083) );
  NOR2_X1 U4764 ( .A1(n4272), .A2(n4075), .ZN(n4079) );
  OAI22_X1 U4765 ( .A1(n4077), .A2(n4643), .B1(n4076), .B2(n4646), .ZN(n4078)
         );
  AOI211_X1 U4766 ( .C1(n4267), .C2(n4306), .A(n4079), .B(n4078), .ZN(n4080)
         );
  OAI21_X1 U4767 ( .B1(n4309), .B2(n4081), .A(n4080), .ZN(n4082) );
  AOI21_X1 U4768 ( .B1(n4083), .B2(n4657), .A(n4082), .ZN(n4084) );
  OAI211_X1 U4769 ( .C1(n4663), .C2(n4308), .A(n4085), .B(n4084), .ZN(U3263)
         );
  XOR2_X1 U4770 ( .A(n4089), .B(n4086), .Z(n4315) );
  INV_X1 U4771 ( .A(n4315), .ZN(n4103) );
  NAND2_X1 U4772 ( .A1(n4088), .A2(n4087), .ZN(n4090) );
  XNOR2_X1 U4773 ( .A(n4090), .B(n4089), .ZN(n4091) );
  NAND2_X1 U4774 ( .A1(n4091), .A2(n4289), .ZN(n4095) );
  OAI22_X1 U4775 ( .A1(n4092), .A2(n4402), .B1(n4401), .B2(n4097), .ZN(n4093)
         );
  INV_X1 U4776 ( .A(n4093), .ZN(n4094) );
  OAI211_X1 U4777 ( .C1(n4327), .C2(n4407), .A(n4095), .B(n4094), .ZN(n4314)
         );
  INV_X1 U4778 ( .A(n4112), .ZN(n4098) );
  OAI21_X1 U4779 ( .B1(n4098), .B2(n4097), .A(n4096), .ZN(n4429) );
  AOI22_X1 U4780 ( .A1(n4099), .A2(n4655), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4663), .ZN(n4100) );
  OAI21_X1 U4781 ( .B1(n4429), .B2(n4233), .A(n4100), .ZN(n4101) );
  AOI21_X1 U4782 ( .B1(n4314), .B2(n4646), .A(n4101), .ZN(n4102) );
  OAI21_X1 U4783 ( .B1(n4103), .B2(n4295), .A(n4102), .ZN(U3264) );
  XOR2_X1 U4784 ( .A(n4105), .B(n2235), .Z(n4319) );
  INV_X1 U4785 ( .A(n4319), .ZN(n4118) );
  XOR2_X1 U4786 ( .A(n4105), .B(n4104), .Z(n4106) );
  NAND2_X1 U4787 ( .A1(n4106), .A2(n4289), .ZN(n4110) );
  AOI22_X1 U4788 ( .A1(n4108), .A2(n4323), .B1(n4107), .B2(n4386), .ZN(n4109)
         );
  OAI211_X1 U4789 ( .C1(n4111), .C2(n4402), .A(n4110), .B(n4109), .ZN(n4318)
         );
  OAI21_X1 U4790 ( .B1(n4127), .B2(n4113), .A(n4112), .ZN(n4433) );
  AOI22_X1 U4791 ( .A1(n4114), .A2(n4655), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4663), .ZN(n4115) );
  OAI21_X1 U4792 ( .B1(n4433), .B2(n4233), .A(n4115), .ZN(n4116) );
  AOI21_X1 U4793 ( .B1(n4318), .B2(n4646), .A(n4116), .ZN(n4117) );
  OAI21_X1 U4794 ( .B1(n4118), .B2(n4295), .A(n4117), .ZN(U3265) );
  XNOR2_X1 U4795 ( .A(n4120), .B(n4119), .ZN(n4329) );
  INV_X1 U4796 ( .A(n4121), .ZN(n4122) );
  NAND2_X1 U4797 ( .A1(n4123), .A2(n4122), .ZN(n4125) );
  XNOR2_X1 U4798 ( .A(n4125), .B(n4124), .ZN(n4126) );
  NAND2_X1 U4799 ( .A1(n4126), .A2(n4289), .ZN(n4326) );
  NOR2_X1 U4800 ( .A1(n4326), .A2(n4663), .ZN(n4139) );
  AND2_X1 U4801 ( .A1(n4158), .A2(n4322), .ZN(n4128) );
  OR2_X1 U4802 ( .A1(n4128), .A2(n4127), .ZN(n4437) );
  NAND2_X1 U4803 ( .A1(n4324), .A2(n4267), .ZN(n4133) );
  NOR2_X1 U4804 ( .A1(n4646), .A2(n4129), .ZN(n4130) );
  AOI21_X1 U4805 ( .B1(n4131), .B2(n4655), .A(n4130), .ZN(n4132) );
  OAI211_X1 U4806 ( .C1(n4272), .C2(n4134), .A(n4133), .B(n4132), .ZN(n4135)
         );
  AOI21_X1 U4807 ( .B1(n4266), .B2(n4136), .A(n4135), .ZN(n4137) );
  OAI21_X1 U4808 ( .B1(n4437), .B2(n4233), .A(n4137), .ZN(n4138) );
  AOI211_X1 U4809 ( .C1(n4329), .C2(n4264), .A(n4139), .B(n4138), .ZN(n4140)
         );
  INV_X1 U4810 ( .A(n4140), .ZN(U3266) );
  XNOR2_X1 U4811 ( .A(n4141), .B(n4151), .ZN(n4333) );
  INV_X1 U4812 ( .A(n4333), .ZN(n4165) );
  INV_X1 U4813 ( .A(n4142), .ZN(n4143) );
  INV_X1 U4814 ( .A(n4144), .ZN(n4145) );
  AOI21_X1 U4815 ( .B1(n4196), .B2(n4147), .A(n4146), .ZN(n4181) );
  INV_X1 U4816 ( .A(n4148), .ZN(n4149) );
  AOI21_X1 U4817 ( .B1(n4181), .B2(n4184), .A(n4149), .ZN(n4169) );
  OAI21_X1 U4818 ( .B1(n4169), .B2(n4168), .A(n4150), .ZN(n4152) );
  XNOR2_X1 U4819 ( .A(n4152), .B(n4151), .ZN(n4153) );
  NAND2_X1 U4820 ( .A1(n4153), .A2(n4289), .ZN(n4156) );
  AOI22_X1 U4821 ( .A1(n4342), .A2(n4323), .B1(n4386), .B2(n4154), .ZN(n4155)
         );
  OAI211_X1 U4822 ( .C1(n4157), .C2(n4402), .A(n4156), .B(n4155), .ZN(n4332)
         );
  OAI21_X1 U4823 ( .B1(n2280), .B2(n4159), .A(n4158), .ZN(n4441) );
  NOR2_X1 U4824 ( .A1(n4441), .A2(n4233), .ZN(n4163) );
  OAI22_X1 U4825 ( .A1(n4161), .A2(n4643), .B1(n4160), .B2(n4646), .ZN(n4162)
         );
  AOI211_X1 U4826 ( .C1(n4332), .C2(n4646), .A(n4163), .B(n4162), .ZN(n4164)
         );
  OAI21_X1 U4827 ( .B1(n4165), .B2(n4295), .A(n4164), .ZN(U3267) );
  OAI21_X1 U4828 ( .B1(n4167), .B2(n4168), .A(n4166), .ZN(n4336) );
  XNOR2_X1 U4829 ( .A(n4169), .B(n4168), .ZN(n4170) );
  NAND2_X1 U4830 ( .A1(n4170), .A2(n4289), .ZN(n4172) );
  AOI22_X1 U4831 ( .A1(n4351), .A2(n4323), .B1(n4174), .B2(n4386), .ZN(n4171)
         );
  OAI211_X1 U4832 ( .C1(n4173), .C2(n4402), .A(n4172), .B(n4171), .ZN(n4337)
         );
  NAND2_X1 U4833 ( .A1(n4185), .A2(n4174), .ZN(n4175) );
  NAND2_X1 U4834 ( .A1(n4176), .A2(n4175), .ZN(n4445) );
  AOI22_X1 U4835 ( .A1(n4177), .A2(n4655), .B1(REG2_REG_22__SCAN_IN), .B2(
        n4663), .ZN(n4178) );
  OAI21_X1 U4836 ( .B1(n4445), .B2(n4233), .A(n4178), .ZN(n4179) );
  AOI21_X1 U4837 ( .B1(n4337), .B2(n4646), .A(n4179), .ZN(n4180) );
  OAI21_X1 U4838 ( .B1(n4336), .B2(n4295), .A(n4180), .ZN(U3268) );
  XNOR2_X1 U4839 ( .A(n4181), .B(n4184), .ZN(n4182) );
  NAND2_X1 U4840 ( .A1(n4182), .A2(n4289), .ZN(n4344) );
  XOR2_X1 U4841 ( .A(n4184), .B(n4183), .Z(n4347) );
  NAND2_X1 U4842 ( .A1(n4347), .A2(n4264), .ZN(n4194) );
  OAI21_X1 U4843 ( .B1(n4203), .B2(n4190), .A(n4185), .ZN(n4449) );
  INV_X1 U4844 ( .A(n4449), .ZN(n4192) );
  AOI22_X1 U4845 ( .A1(n4342), .A2(n4266), .B1(n4267), .B2(n4225), .ZN(n4189)
         );
  INV_X1 U4846 ( .A(n4186), .ZN(n4187) );
  AOI22_X1 U4847 ( .A1(n4663), .A2(REG2_REG_21__SCAN_IN), .B1(n4187), .B2(
        n4655), .ZN(n4188) );
  OAI211_X1 U4848 ( .C1(n4190), .C2(n4272), .A(n4189), .B(n4188), .ZN(n4191)
         );
  AOI21_X1 U4849 ( .B1(n4192), .B2(n4657), .A(n4191), .ZN(n4193) );
  OAI211_X1 U4850 ( .C1(n4663), .C2(n4344), .A(n4194), .B(n4193), .ZN(U3269)
         );
  NAND2_X1 U4851 ( .A1(n4196), .A2(n4195), .ZN(n4197) );
  XNOR2_X1 U4852 ( .A(n4197), .B(n4201), .ZN(n4198) );
  NAND2_X1 U4853 ( .A1(n4198), .A2(n4289), .ZN(n4353) );
  AOI21_X1 U4854 ( .B1(n4215), .B2(n4200), .A(n4199), .ZN(n4202) );
  XNOR2_X1 U4855 ( .A(n4202), .B(n4201), .ZN(n4356) );
  NAND2_X1 U4856 ( .A1(n4356), .A2(n4264), .ZN(n4214) );
  INV_X1 U4857 ( .A(n4203), .ZN(n4204) );
  OAI21_X1 U4858 ( .B1(n4229), .B2(n4205), .A(n4204), .ZN(n4453) );
  INV_X1 U4859 ( .A(n4453), .ZN(n4212) );
  INV_X1 U4860 ( .A(n4249), .ZN(n4354) );
  AOI22_X1 U4861 ( .A1(n4266), .A2(n4351), .B1(n4206), .B2(n4350), .ZN(n4209)
         );
  AOI22_X1 U4862 ( .A1(n4663), .A2(REG2_REG_20__SCAN_IN), .B1(n4207), .B2(
        n4655), .ZN(n4208) );
  OAI211_X1 U4863 ( .C1(n4354), .C2(n4210), .A(n4209), .B(n4208), .ZN(n4211)
         );
  AOI21_X1 U4864 ( .B1(n4212), .B2(n4657), .A(n4211), .ZN(n4213) );
  OAI211_X1 U4865 ( .C1(n4663), .C2(n4353), .A(n4214), .B(n4213), .ZN(U3270)
         );
  XOR2_X1 U4866 ( .A(n4222), .B(n4215), .Z(n4360) );
  INV_X1 U4867 ( .A(n4360), .ZN(n4239) );
  NAND2_X1 U4868 ( .A1(n4217), .A2(n4216), .ZN(n4247) );
  INV_X1 U4869 ( .A(n4218), .ZN(n4220) );
  OAI21_X1 U4870 ( .B1(n4247), .B2(n4220), .A(n4219), .ZN(n4221) );
  XOR2_X1 U4871 ( .A(n4222), .B(n4221), .Z(n4223) );
  NAND2_X1 U4872 ( .A1(n4223), .A2(n4289), .ZN(n4227) );
  AOI22_X1 U4873 ( .A1(n4225), .A2(n4388), .B1(n4386), .B2(n4224), .ZN(n4226)
         );
  OAI211_X1 U4874 ( .C1(n4228), .C2(n4407), .A(n4227), .B(n4226), .ZN(n4359)
         );
  INV_X1 U4875 ( .A(n4244), .ZN(n4232) );
  INV_X1 U4876 ( .A(n4229), .ZN(n4230) );
  OAI21_X1 U4877 ( .B1(n4232), .B2(n4231), .A(n4230), .ZN(n4457) );
  NOR2_X1 U4878 ( .A1(n4457), .A2(n4233), .ZN(n4237) );
  OAI22_X1 U4879 ( .A1(n4646), .A2(n4235), .B1(n4234), .B2(n4643), .ZN(n4236)
         );
  AOI211_X1 U4880 ( .C1(n4359), .C2(n4646), .A(n4237), .B(n4236), .ZN(n4238)
         );
  OAI21_X1 U4881 ( .B1(n4239), .B2(n4295), .A(n4238), .ZN(U3271) );
  OAI21_X1 U4882 ( .B1(n4242), .B2(n4241), .A(n4240), .ZN(n4243) );
  INV_X1 U4883 ( .A(n4243), .ZN(n4364) );
  INV_X1 U4884 ( .A(n4265), .ZN(n4246) );
  OAI211_X1 U4885 ( .C1(n4246), .C2(n4245), .A(n4710), .B(n4244), .ZN(n4362)
         );
  XNOR2_X1 U4886 ( .A(n4247), .B(n2334), .ZN(n4252) );
  AOI22_X1 U4887 ( .A1(n4249), .A2(n4388), .B1(n4386), .B2(n4248), .ZN(n4250)
         );
  OAI21_X1 U4888 ( .B1(n4286), .B2(n4407), .A(n4250), .ZN(n4251) );
  AOI21_X1 U4889 ( .B1(n4252), .B2(n4289), .A(n4251), .ZN(n4363) );
  OAI21_X1 U4890 ( .B1(n4253), .B2(n4362), .A(n4363), .ZN(n4257) );
  OAI22_X1 U4891 ( .A1(n4646), .A2(n4255), .B1(n4254), .B2(n4643), .ZN(n4256)
         );
  AOI21_X1 U4892 ( .B1(n4257), .B2(n4646), .A(n4256), .ZN(n4258) );
  OAI21_X1 U4893 ( .B1(n4364), .B2(n4295), .A(n4258), .ZN(U3272) );
  INV_X1 U4894 ( .A(n4262), .ZN(n4259) );
  XNOR2_X1 U4895 ( .A(n4260), .B(n4259), .ZN(n4261) );
  NAND2_X1 U4896 ( .A1(n4261), .A2(n4289), .ZN(n4368) );
  XNOR2_X1 U4897 ( .A(n4263), .B(n4262), .ZN(n4371) );
  NAND2_X1 U4898 ( .A1(n4371), .A2(n4264), .ZN(n4277) );
  OAI21_X1 U4899 ( .B1(n4280), .B2(n4273), .A(n4265), .ZN(n4462) );
  INV_X1 U4900 ( .A(n4462), .ZN(n4275) );
  AOI22_X1 U4901 ( .A1(n4267), .A2(n4379), .B1(n4366), .B2(n4266), .ZN(n4271)
         );
  INV_X1 U4902 ( .A(n4268), .ZN(n4269) );
  AOI22_X1 U4903 ( .A1(n4663), .A2(REG2_REG_17__SCAN_IN), .B1(n4269), .B2(
        n4655), .ZN(n4270) );
  OAI211_X1 U4904 ( .C1(n4273), .C2(n4272), .A(n4271), .B(n4270), .ZN(n4274)
         );
  AOI21_X1 U4905 ( .B1(n4275), .B2(n4657), .A(n4274), .ZN(n4276) );
  OAI211_X1 U4906 ( .C1(n4663), .C2(n4368), .A(n4277), .B(n4276), .ZN(U3273)
         );
  OAI21_X1 U4907 ( .B1(n4279), .B2(n4284), .A(n4278), .ZN(n4374) );
  INV_X1 U4908 ( .A(n4280), .ZN(n4281) );
  OAI21_X1 U4909 ( .B1(n4282), .B2(n4499), .A(n4281), .ZN(n4466) );
  INV_X1 U4910 ( .A(n4466), .ZN(n4293) );
  OAI22_X1 U4911 ( .A1(n4646), .A2(n4283), .B1(n4512), .B2(n4643), .ZN(n4292)
         );
  XNOR2_X1 U4912 ( .A(n4285), .B(n4284), .ZN(n4290) );
  NOR2_X1 U4913 ( .A1(n4498), .A2(n4407), .ZN(n4288) );
  OAI22_X1 U4914 ( .A1(n4286), .A2(n4402), .B1(n4499), .B2(n4401), .ZN(n4287)
         );
  AOI211_X1 U4915 ( .C1(n4290), .C2(n4289), .A(n4288), .B(n4287), .ZN(n4373)
         );
  NOR2_X1 U4916 ( .A1(n4373), .A2(n4663), .ZN(n4291) );
  AOI211_X1 U4917 ( .C1(n4293), .C2(n4657), .A(n4292), .B(n4291), .ZN(n4294)
         );
  OAI21_X1 U4918 ( .B1(n4374), .B2(n4295), .A(n4294), .ZN(U3274) );
  NAND2_X1 U4919 ( .A1(n4415), .A2(n4722), .ZN(n4297) );
  NAND2_X1 U4920 ( .A1(n4719), .A2(REG1_REG_31__SCAN_IN), .ZN(n4296) );
  OAI211_X1 U4921 ( .C1(n4418), .C2(n4414), .A(n4297), .B(n4296), .ZN(U3549)
         );
  AOI21_X1 U4922 ( .B1(n4302), .B2(n4299), .A(n4298), .ZN(n4514) );
  INV_X1 U4923 ( .A(n4514), .ZN(n4421) );
  INV_X1 U4924 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4303) );
  INV_X1 U4925 ( .A(n4300), .ZN(n4301) );
  AOI21_X1 U4926 ( .B1(n4302), .B2(n4386), .A(n4301), .ZN(n4516) );
  MUX2_X1 U4927 ( .A(n4303), .B(n4516), .S(n4722), .Z(n4304) );
  OAI21_X1 U4928 ( .B1(n4421), .B2(n4414), .A(n4304), .ZN(U3548) );
  INV_X1 U4929 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4312) );
  AOI22_X1 U4930 ( .A1(n4306), .A2(n4323), .B1(n4305), .B2(n4386), .ZN(n4307)
         );
  OAI211_X1 U4931 ( .C1(n4309), .C2(n4402), .A(n4308), .B(n4307), .ZN(n4310)
         );
  AOI21_X1 U4932 ( .B1(n4311), .B2(n4411), .A(n4310), .ZN(n4422) );
  MUX2_X1 U4933 ( .A(n4312), .B(n4422), .S(n4722), .Z(n4313) );
  OAI21_X1 U4934 ( .B1(n4414), .B2(n4425), .A(n4313), .ZN(U3545) );
  INV_X1 U4935 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4316) );
  AOI21_X1 U4936 ( .B1(n4315), .B2(n4411), .A(n4314), .ZN(n4426) );
  MUX2_X1 U4937 ( .A(n4316), .B(n4426), .S(n4722), .Z(n4317) );
  OAI21_X1 U4938 ( .B1(n4414), .B2(n4429), .A(n4317), .ZN(U3544) );
  INV_X1 U4939 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4320) );
  AOI21_X1 U4940 ( .B1(n4319), .B2(n4411), .A(n4318), .ZN(n4430) );
  MUX2_X1 U4941 ( .A(n4320), .B(n4430), .S(n4722), .Z(n4321) );
  OAI21_X1 U4942 ( .B1(n4414), .B2(n4433), .A(n4321), .ZN(U3543) );
  INV_X1 U4943 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4330) );
  AOI22_X1 U4944 ( .A1(n4324), .A2(n4323), .B1(n4322), .B2(n4386), .ZN(n4325)
         );
  OAI211_X1 U4945 ( .C1(n4327), .C2(n4402), .A(n4326), .B(n4325), .ZN(n4328)
         );
  AOI21_X1 U4946 ( .B1(n4329), .B2(n4411), .A(n4328), .ZN(n4434) );
  MUX2_X1 U4947 ( .A(n4330), .B(n4434), .S(n4722), .Z(n4331) );
  OAI21_X1 U4948 ( .B1(n4414), .B2(n4437), .A(n4331), .ZN(U3542) );
  INV_X1 U4949 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4334) );
  AOI21_X1 U4950 ( .B1(n4333), .B2(n4411), .A(n4332), .ZN(n4438) );
  MUX2_X1 U4951 ( .A(n4334), .B(n4438), .S(n4722), .Z(n4335) );
  OAI21_X1 U4952 ( .B1(n4414), .B2(n4441), .A(n4335), .ZN(U3541) );
  INV_X1 U4953 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4339) );
  INV_X1 U4954 ( .A(n4336), .ZN(n4338) );
  AOI21_X1 U4955 ( .B1(n4338), .B2(n4411), .A(n4337), .ZN(n4442) );
  MUX2_X1 U4956 ( .A(n4339), .B(n4442), .S(n4722), .Z(n4340) );
  OAI21_X1 U4957 ( .B1(n4414), .B2(n4445), .A(n4340), .ZN(U3540) );
  INV_X1 U4958 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4348) );
  AOI22_X1 U4959 ( .A1(n4342), .A2(n4388), .B1(n4386), .B2(n4341), .ZN(n4343)
         );
  OAI211_X1 U4960 ( .C1(n4345), .C2(n4407), .A(n4344), .B(n4343), .ZN(n4346)
         );
  AOI21_X1 U4961 ( .B1(n4347), .B2(n4411), .A(n4346), .ZN(n4446) );
  MUX2_X1 U4962 ( .A(n4348), .B(n4446), .S(n4722), .Z(n4349) );
  OAI21_X1 U4963 ( .B1(n4414), .B2(n4449), .A(n4349), .ZN(U3539) );
  INV_X1 U4964 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4357) );
  AOI22_X1 U4965 ( .A1(n4351), .A2(n4388), .B1(n4350), .B2(n4386), .ZN(n4352)
         );
  OAI211_X1 U4966 ( .C1(n4354), .C2(n4407), .A(n4353), .B(n4352), .ZN(n4355)
         );
  AOI21_X1 U4967 ( .B1(n4356), .B2(n4411), .A(n4355), .ZN(n4450) );
  MUX2_X1 U4968 ( .A(n4357), .B(n4450), .S(n4722), .Z(n4358) );
  OAI21_X1 U4969 ( .B1(n4414), .B2(n4453), .A(n4358), .ZN(U3538) );
  AOI21_X1 U4970 ( .B1(n4360), .B2(n4411), .A(n4359), .ZN(n4454) );
  MUX2_X1 U4971 ( .A(n4052), .B(n4454), .S(n4722), .Z(n4361) );
  OAI21_X1 U4972 ( .B1(n4414), .B2(n4457), .A(n4361), .ZN(U3537) );
  OAI211_X1 U4973 ( .C1(n4364), .C2(n4699), .A(n4363), .B(n4362), .ZN(n4458)
         );
  MUX2_X1 U4974 ( .A(REG1_REG_18__SCAN_IN), .B(n4458), .S(n4722), .Z(U3536) );
  AOI22_X1 U4975 ( .A1(n4366), .A2(n4388), .B1(n4386), .B2(n4365), .ZN(n4367)
         );
  OAI211_X1 U4976 ( .C1(n4369), .C2(n4407), .A(n4368), .B(n4367), .ZN(n4370)
         );
  AOI21_X1 U4977 ( .B1(n4371), .B2(n4411), .A(n4370), .ZN(n4459) );
  MUX2_X1 U4978 ( .A(n4048), .B(n4459), .S(n4722), .Z(n4372) );
  OAI21_X1 U4979 ( .B1(n4414), .B2(n4462), .A(n4372), .ZN(U3535) );
  INV_X1 U4980 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4376) );
  OAI21_X1 U4981 ( .B1(n4374), .B2(n4699), .A(n4373), .ZN(n4375) );
  INV_X1 U4982 ( .A(n4375), .ZN(n4463) );
  MUX2_X1 U4983 ( .A(n4376), .B(n4463), .S(n4722), .Z(n4377) );
  OAI21_X1 U4984 ( .B1(n4414), .B2(n4466), .A(n4377), .ZN(U3534) );
  AOI22_X1 U4985 ( .A1(n4379), .A2(n4388), .B1(n4386), .B2(n4378), .ZN(n4380)
         );
  OAI211_X1 U4986 ( .C1(n4382), .C2(n4407), .A(n4381), .B(n4380), .ZN(n4383)
         );
  AOI21_X1 U4987 ( .B1(n4384), .B2(n4411), .A(n4383), .ZN(n4467) );
  MUX2_X1 U4988 ( .A(n4022), .B(n4467), .S(n4722), .Z(n4385) );
  OAI21_X1 U4989 ( .B1(n4414), .B2(n4470), .A(n4385), .ZN(U3533) );
  INV_X1 U4990 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4395) );
  AOI22_X1 U4991 ( .A1(n4389), .A2(n4388), .B1(n4387), .B2(n4386), .ZN(n4390)
         );
  OAI21_X1 U4992 ( .B1(n4403), .B2(n4407), .A(n4390), .ZN(n4393) );
  INV_X1 U4993 ( .A(n4391), .ZN(n4392) );
  AOI211_X1 U4994 ( .C1(n4697), .C2(n4394), .A(n4393), .B(n4392), .ZN(n4471)
         );
  MUX2_X1 U4995 ( .A(n4395), .B(n4471), .S(n4722), .Z(n4396) );
  OAI21_X1 U4996 ( .B1(n4414), .B2(n4474), .A(n4396), .ZN(U3532) );
  AOI21_X1 U4997 ( .B1(n4398), .B2(n4411), .A(n4397), .ZN(n4475) );
  MUX2_X1 U4998 ( .A(n4024), .B(n4475), .S(n4722), .Z(n4399) );
  OAI21_X1 U4999 ( .B1(n4414), .B2(n4479), .A(n4399), .ZN(U3531) );
  INV_X1 U5000 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4412) );
  OAI22_X1 U5001 ( .A1(n4403), .A2(n4402), .B1(n4401), .B2(n4400), .ZN(n4404)
         );
  INV_X1 U5002 ( .A(n4404), .ZN(n4405) );
  OAI211_X1 U5003 ( .C1(n4408), .C2(n4407), .A(n4406), .B(n4405), .ZN(n4409)
         );
  AOI21_X1 U5004 ( .B1(n4411), .B2(n4410), .A(n4409), .ZN(n4480) );
  MUX2_X1 U5005 ( .A(n4412), .B(n4480), .S(n4722), .Z(n4413) );
  OAI21_X1 U5006 ( .B1(n4483), .B2(n4414), .A(n4413), .ZN(U3530) );
  NAND2_X1 U5007 ( .A1(n4415), .A2(n4713), .ZN(n4417) );
  NAND2_X1 U5008 ( .A1(n4711), .A2(REG0_REG_31__SCAN_IN), .ZN(n4416) );
  OAI211_X1 U5009 ( .C1(n4418), .C2(n4478), .A(n4417), .B(n4416), .ZN(U3517)
         );
  INV_X1 U5010 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4419) );
  MUX2_X1 U5011 ( .A(n4419), .B(n4516), .S(n4713), .Z(n4420) );
  OAI21_X1 U5012 ( .B1(n4421), .B2(n4478), .A(n4420), .ZN(U3516) );
  INV_X1 U5013 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4423) );
  MUX2_X1 U5014 ( .A(n4423), .B(n4422), .S(n4713), .Z(n4424) );
  OAI21_X1 U5015 ( .B1(n4425), .B2(n4478), .A(n4424), .ZN(U3513) );
  INV_X1 U5016 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4427) );
  MUX2_X1 U5017 ( .A(n4427), .B(n4426), .S(n4713), .Z(n4428) );
  OAI21_X1 U5018 ( .B1(n4429), .B2(n4478), .A(n4428), .ZN(U3512) );
  INV_X1 U5019 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4431) );
  MUX2_X1 U5020 ( .A(n4431), .B(n4430), .S(n4713), .Z(n4432) );
  OAI21_X1 U5021 ( .B1(n4433), .B2(n4478), .A(n4432), .ZN(U3511) );
  INV_X1 U5022 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4435) );
  MUX2_X1 U5023 ( .A(n4435), .B(n4434), .S(n4713), .Z(n4436) );
  OAI21_X1 U5024 ( .B1(n4437), .B2(n4478), .A(n4436), .ZN(U3510) );
  INV_X1 U5025 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4439) );
  MUX2_X1 U5026 ( .A(n4439), .B(n4438), .S(n4713), .Z(n4440) );
  OAI21_X1 U5027 ( .B1(n4441), .B2(n4478), .A(n4440), .ZN(U3509) );
  INV_X1 U5028 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4443) );
  MUX2_X1 U5029 ( .A(n4443), .B(n4442), .S(n4713), .Z(n4444) );
  OAI21_X1 U5030 ( .B1(n4445), .B2(n4478), .A(n4444), .ZN(U3508) );
  INV_X1 U5031 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4447) );
  MUX2_X1 U5032 ( .A(n4447), .B(n4446), .S(n4713), .Z(n4448) );
  OAI21_X1 U5033 ( .B1(n4449), .B2(n4478), .A(n4448), .ZN(U3507) );
  INV_X1 U5034 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4451) );
  MUX2_X1 U5035 ( .A(n4451), .B(n4450), .S(n4713), .Z(n4452) );
  OAI21_X1 U5036 ( .B1(n4453), .B2(n4478), .A(n4452), .ZN(U3506) );
  INV_X1 U5037 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4455) );
  MUX2_X1 U5038 ( .A(n4455), .B(n4454), .S(n4713), .Z(n4456) );
  OAI21_X1 U5039 ( .B1(n4457), .B2(n4478), .A(n4456), .ZN(U3505) );
  MUX2_X1 U5040 ( .A(REG0_REG_18__SCAN_IN), .B(n4458), .S(n4713), .Z(U3503) );
  INV_X1 U5041 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4460) );
  MUX2_X1 U5042 ( .A(n4460), .B(n4459), .S(n4713), .Z(n4461) );
  OAI21_X1 U5043 ( .B1(n4462), .B2(n4478), .A(n4461), .ZN(U3501) );
  INV_X1 U5044 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4464) );
  MUX2_X1 U5045 ( .A(n4464), .B(n4463), .S(n4713), .Z(n4465) );
  OAI21_X1 U5046 ( .B1(n4466), .B2(n4478), .A(n4465), .ZN(U3499) );
  INV_X1 U5047 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4468) );
  MUX2_X1 U5048 ( .A(n4468), .B(n4467), .S(n4713), .Z(n4469) );
  OAI21_X1 U5049 ( .B1(n4470), .B2(n4478), .A(n4469), .ZN(U3497) );
  INV_X1 U5050 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4472) );
  MUX2_X1 U5051 ( .A(n4472), .B(n4471), .S(n4713), .Z(n4473) );
  OAI21_X1 U5052 ( .B1(n4474), .B2(n4478), .A(n4473), .ZN(U3495) );
  INV_X1 U5053 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4476) );
  MUX2_X1 U5054 ( .A(n4476), .B(n4475), .S(n4713), .Z(n4477) );
  OAI21_X1 U5055 ( .B1(n4479), .B2(n4478), .A(n4477), .ZN(U3493) );
  INV_X1 U5056 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4481) );
  MUX2_X1 U5057 ( .A(n4481), .B(n4480), .S(n4713), .Z(n4482) );
  OAI21_X1 U5058 ( .B1(n4483), .B2(n4478), .A(n4482), .ZN(U3491) );
  MUX2_X1 U5059 ( .A(n2499), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U5060 ( .A(n4484), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5061 ( .A(n4485), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5062 ( .A(n4486), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5063 ( .A(n4487), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5064 ( .A(DATAI_20_), .B(n4488), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5065 ( .A(DATAI_7_), .B(n4489), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U5066 ( .A(n4490), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5067 ( .A(n4491), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5068 ( .A(DATAI_4_), .B(n4492), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5069 ( .A(DATAI_3_), .B(n4493), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5070 ( .A(DATAI_2_), .B(n4494), .S(STATE_REG_SCAN_IN), .Z(U3350) );
  AOI22_X1 U5071 ( .A1(STATE_REG_SCAN_IN), .A2(n4495), .B1(n4805), .B2(U3149), 
        .ZN(U3324) );
  INV_X1 U5072 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4496) );
  NOR2_X1 U5073 ( .A1(STATE_REG_SCAN_IN), .A2(n4496), .ZN(n4608) );
  OAI22_X1 U5074 ( .A1(n4500), .A2(n4499), .B1(n4498), .B2(n4497), .ZN(n4501)
         );
  AOI211_X1 U5075 ( .C1(n4503), .C2(n4502), .A(n4608), .B(n4501), .ZN(n4511)
         );
  OAI21_X1 U5076 ( .B1(n3783), .B2(n4505), .A(n4504), .ZN(n4506) );
  XOR2_X1 U5077 ( .A(n4507), .B(n4506), .Z(n4509) );
  NAND2_X1 U5078 ( .A1(n4509), .A2(n4508), .ZN(n4510) );
  OAI211_X1 U5079 ( .C1(n4513), .C2(n4512), .A(n4511), .B(n4510), .ZN(U3223)
         );
  AOI22_X1 U5080 ( .A1(n4514), .A2(n4657), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4663), .ZN(n4515) );
  OAI21_X1 U5081 ( .B1(n4663), .B2(n4516), .A(n4515), .ZN(U3261) );
  INV_X1 U5082 ( .A(n4519), .ZN(n4517) );
  OAI211_X1 U5083 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4518), .A(n4517), .B(n4520), 
        .ZN(n4523) );
  AOI22_X1 U5084 ( .A1(n4520), .A2(n4519), .B1(n4631), .B2(n2867), .ZN(n4522)
         );
  AOI22_X1 U5085 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4629), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4521) );
  OAI221_X1 U5086 ( .B1(IR_REG_0__SCAN_IN), .B2(n4523), .C1(n4986), .C2(n4522), 
        .A(n4521), .ZN(U3240) );
  OAI211_X1 U5087 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4525), .A(n4575), .B(n4524), 
        .ZN(n4527) );
  NAND2_X1 U5088 ( .A1(n4527), .A2(n4526), .ZN(n4528) );
  AOI21_X1 U5089 ( .B1(n4629), .B2(ADDR_REG_8__SCAN_IN), .A(n4528), .ZN(n4532)
         );
  OAI211_X1 U5090 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4530), .A(n4631), .B(n4529), 
        .ZN(n4531) );
  OAI211_X1 U5091 ( .C1(n4635), .C2(n4685), .A(n4532), .B(n4531), .ZN(U3248)
         );
  OAI211_X1 U5092 ( .C1(n4535), .C2(n4534), .A(n4631), .B(n4533), .ZN(n4540)
         );
  OAI211_X1 U5093 ( .C1(n4538), .C2(n4537), .A(n4575), .B(n4536), .ZN(n4539)
         );
  OAI211_X1 U5094 ( .C1(n4635), .C2(n4684), .A(n4540), .B(n4539), .ZN(n4541)
         );
  AOI211_X1 U5095 ( .C1(n4629), .C2(ADDR_REG_9__SCAN_IN), .A(n4542), .B(n4541), 
        .ZN(n4543) );
  INV_X1 U5096 ( .A(n4543), .ZN(U3249) );
  OAI211_X1 U5097 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4546), .A(n4575), .B(n4545), .ZN(n4548) );
  NAND2_X1 U5098 ( .A1(n4548), .A2(n4547), .ZN(n4549) );
  AOI21_X1 U5099 ( .B1(n4629), .B2(ADDR_REG_10__SCAN_IN), .A(n4549), .ZN(n4553) );
  OAI211_X1 U5100 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4551), .A(n4631), .B(n4550), .ZN(n4552) );
  OAI211_X1 U5101 ( .C1(n4635), .C2(n2359), .A(n4553), .B(n4552), .ZN(U3250)
         );
  OAI211_X1 U5102 ( .C1(n4556), .C2(n4555), .A(n4631), .B(n4554), .ZN(n4561)
         );
  OAI211_X1 U5103 ( .C1(n4559), .C2(n4558), .A(n4575), .B(n4557), .ZN(n4560)
         );
  OAI211_X1 U5104 ( .C1(n4635), .C2(n4682), .A(n4561), .B(n4560), .ZN(n4562)
         );
  AOI211_X1 U5105 ( .C1(n4629), .C2(ADDR_REG_11__SCAN_IN), .A(n4563), .B(n4562), .ZN(n4564) );
  INV_X1 U5106 ( .A(n4564), .ZN(U3251) );
  OAI211_X1 U5107 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4566), .A(n4631), .B(n4565), .ZN(n4570) );
  OAI211_X1 U5108 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4568), .A(n4575), .B(n4567), .ZN(n4569) );
  OAI211_X1 U5109 ( .C1(n4635), .C2(n4037), .A(n4570), .B(n4569), .ZN(n4571)
         );
  AOI211_X1 U5110 ( .C1(n4629), .C2(ADDR_REG_12__SCAN_IN), .A(n4572), .B(n4571), .ZN(n4573) );
  INV_X1 U5111 ( .A(n4573), .ZN(U3252) );
  AOI21_X1 U5112 ( .B1(n3603), .B2(n4681), .A(n4574), .ZN(n4578) );
  OAI21_X1 U5113 ( .B1(n4578), .B2(n4577), .A(n4575), .ZN(n4576) );
  AOI21_X1 U5114 ( .B1(n4578), .B2(n4577), .A(n4576), .ZN(n4579) );
  AOI211_X1 U5115 ( .C1(n4629), .C2(ADDR_REG_13__SCAN_IN), .A(n4580), .B(n4579), .ZN(n4585) );
  OAI211_X1 U5116 ( .C1(n4583), .C2(n4582), .A(n4631), .B(n4581), .ZN(n4584)
         );
  OAI211_X1 U5117 ( .C1(n4635), .C2(n4681), .A(n4585), .B(n4584), .ZN(U3253)
         );
  INV_X1 U5118 ( .A(n4586), .ZN(n4590) );
  AOI211_X1 U5119 ( .C1(n3563), .C2(n4588), .A(n4587), .B(n4624), .ZN(n4589)
         );
  AOI211_X1 U5120 ( .C1(n4629), .C2(ADDR_REG_14__SCAN_IN), .A(n4590), .B(n4589), .ZN(n4594) );
  OAI211_X1 U5121 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4592), .A(n4631), .B(n4591), .ZN(n4593) );
  OAI211_X1 U5122 ( .C1(n4635), .C2(n2368), .A(n4594), .B(n4593), .ZN(U3254)
         );
  AOI211_X1 U5123 ( .C1(n4597), .C2(n4596), .A(n4595), .B(n4624), .ZN(n4598)
         );
  AOI211_X1 U5124 ( .C1(n4629), .C2(ADDR_REG_15__SCAN_IN), .A(n4599), .B(n4598), .ZN(n4604) );
  OAI211_X1 U5125 ( .C1(n4602), .C2(n4601), .A(n4631), .B(n4600), .ZN(n4603)
         );
  OAI211_X1 U5126 ( .C1(n4635), .C2(n4679), .A(n4604), .B(n4603), .ZN(U3255)
         );
  AOI221_X1 U5127 ( .B1(n4606), .B2(n4605), .C1(n4283), .C2(n4605), .A(n4624), 
        .ZN(n4607) );
  AOI211_X1 U5128 ( .C1(n4629), .C2(ADDR_REG_16__SCAN_IN), .A(n4608), .B(n4607), .ZN(n4612) );
  OAI221_X1 U5129 ( .B1(n4610), .B2(REG1_REG_16__SCAN_IN), .C1(n4610), .C2(
        n4609), .A(n4631), .ZN(n4611) );
  OAI211_X1 U5130 ( .C1(n4635), .C2(n4678), .A(n4612), .B(n4611), .ZN(U3256)
         );
  AOI221_X1 U5131 ( .B1(n4615), .B2(n4614), .C1(n4613), .C2(n4614), .A(n4624), 
        .ZN(n4616) );
  AOI211_X1 U5132 ( .C1(n4629), .C2(ADDR_REG_17__SCAN_IN), .A(n4617), .B(n4616), .ZN(n4622) );
  OAI221_X1 U5133 ( .B1(n4620), .B2(n4619), .C1(n4620), .C2(n4618), .A(n4631), 
        .ZN(n4621) );
  OAI211_X1 U5134 ( .C1(n4635), .C2(n4677), .A(n4622), .B(n4621), .ZN(U3257)
         );
  NOR2_X1 U5135 ( .A1(STATE_REG_SCAN_IN), .A2(n4623), .ZN(n4628) );
  OAI211_X1 U5136 ( .C1(n4633), .C2(n4632), .A(n4631), .B(n4630), .ZN(n4634)
         );
  AOI22_X1 U5137 ( .A1(n4636), .A2(n4655), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4663), .ZN(n4641) );
  INV_X1 U5138 ( .A(n4637), .ZN(n4638) );
  AOI22_X1 U5139 ( .A1(n4639), .A2(n4658), .B1(n4657), .B2(n4638), .ZN(n4640)
         );
  OAI211_X1 U5140 ( .C1(n4663), .C2(n4642), .A(n4641), .B(n4640), .ZN(U3280)
         );
  OAI22_X1 U5141 ( .A1(n4646), .A2(n4645), .B1(n4644), .B2(n4643), .ZN(n4647)
         );
  INV_X1 U5142 ( .A(n4647), .ZN(n4652) );
  INV_X1 U5143 ( .A(n4648), .ZN(n4649) );
  AOI22_X1 U5144 ( .A1(n4650), .A2(n4658), .B1(n4657), .B2(n4649), .ZN(n4651)
         );
  OAI211_X1 U5145 ( .C1(n4663), .C2(n4653), .A(n4652), .B(n4651), .ZN(U3282)
         );
  INV_X1 U5146 ( .A(n4654), .ZN(n4662) );
  AOI22_X1 U5147 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4663), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4655), .ZN(n4661) );
  AOI22_X1 U5148 ( .A1(n4659), .A2(n4658), .B1(n4657), .B2(n4656), .ZN(n4660)
         );
  OAI211_X1 U5149 ( .C1(n4663), .C2(n4662), .A(n4661), .B(n4660), .ZN(U3288)
         );
  INV_X1 U5150 ( .A(D_REG_31__SCAN_IN), .ZN(n4859) );
  NOR2_X1 U5151 ( .A1(n4674), .A2(n4859), .ZN(U3291) );
  INV_X1 U5152 ( .A(D_REG_30__SCAN_IN), .ZN(n4664) );
  NOR2_X1 U5153 ( .A1(n4674), .A2(n4664), .ZN(U3292) );
  INV_X1 U5154 ( .A(D_REG_29__SCAN_IN), .ZN(n4819) );
  NOR2_X1 U5155 ( .A1(n4674), .A2(n4819), .ZN(U3293) );
  INV_X1 U5156 ( .A(D_REG_28__SCAN_IN), .ZN(n4665) );
  NOR2_X1 U5157 ( .A1(n4674), .A2(n4665), .ZN(U3294) );
  INV_X1 U5158 ( .A(D_REG_27__SCAN_IN), .ZN(n4882) );
  NOR2_X1 U5159 ( .A1(n4674), .A2(n4882), .ZN(U3295) );
  INV_X1 U5160 ( .A(D_REG_26__SCAN_IN), .ZN(n4808) );
  NOR2_X1 U5161 ( .A1(n4674), .A2(n4808), .ZN(U3296) );
  INV_X1 U5162 ( .A(D_REG_25__SCAN_IN), .ZN(n4666) );
  NOR2_X1 U5163 ( .A1(n4674), .A2(n4666), .ZN(U3297) );
  INV_X1 U5164 ( .A(D_REG_24__SCAN_IN), .ZN(n5034) );
  NOR2_X1 U5165 ( .A1(n4674), .A2(n5034), .ZN(U3298) );
  INV_X1 U5166 ( .A(D_REG_23__SCAN_IN), .ZN(n4667) );
  NOR2_X1 U5167 ( .A1(n4674), .A2(n4667), .ZN(U3299) );
  INV_X1 U5168 ( .A(D_REG_22__SCAN_IN), .ZN(n5013) );
  NOR2_X1 U5169 ( .A1(n4674), .A2(n5013), .ZN(U3300) );
  INV_X1 U5170 ( .A(D_REG_21__SCAN_IN), .ZN(n4668) );
  NOR2_X1 U5171 ( .A1(n4674), .A2(n4668), .ZN(U3301) );
  INV_X1 U5172 ( .A(D_REG_20__SCAN_IN), .ZN(n4800) );
  NOR2_X1 U5173 ( .A1(n4674), .A2(n4800), .ZN(U3302) );
  INV_X1 U5174 ( .A(D_REG_19__SCAN_IN), .ZN(n5026) );
  NOR2_X1 U5175 ( .A1(n4674), .A2(n5026), .ZN(U3303) );
  INV_X1 U5176 ( .A(D_REG_18__SCAN_IN), .ZN(n5025) );
  NOR2_X1 U5177 ( .A1(n4674), .A2(n5025), .ZN(U3304) );
  INV_X1 U5178 ( .A(D_REG_17__SCAN_IN), .ZN(n5031) );
  NOR2_X1 U5179 ( .A1(n4674), .A2(n5031), .ZN(U3305) );
  INV_X1 U5180 ( .A(D_REG_16__SCAN_IN), .ZN(n4669) );
  NOR2_X1 U5181 ( .A1(n4674), .A2(n4669), .ZN(U3306) );
  INV_X1 U5182 ( .A(D_REG_15__SCAN_IN), .ZN(n4670) );
  NOR2_X1 U5183 ( .A1(n4674), .A2(n4670), .ZN(U3307) );
  INV_X1 U5184 ( .A(D_REG_14__SCAN_IN), .ZN(n5032) );
  NOR2_X1 U5185 ( .A1(n4674), .A2(n5032), .ZN(U3308) );
  INV_X1 U5186 ( .A(D_REG_13__SCAN_IN), .ZN(n4671) );
  NOR2_X1 U5187 ( .A1(n4674), .A2(n4671), .ZN(U3309) );
  INV_X1 U5188 ( .A(D_REG_12__SCAN_IN), .ZN(n5028) );
  NOR2_X1 U5189 ( .A1(n4674), .A2(n5028), .ZN(U3310) );
  INV_X1 U5190 ( .A(D_REG_11__SCAN_IN), .ZN(n5012) );
  NOR2_X1 U5191 ( .A1(n4674), .A2(n5012), .ZN(U3311) );
  INV_X1 U5192 ( .A(D_REG_10__SCAN_IN), .ZN(n5035) );
  NOR2_X1 U5193 ( .A1(n4674), .A2(n5035), .ZN(U3312) );
  INV_X1 U5194 ( .A(D_REG_9__SCAN_IN), .ZN(n5029) );
  NOR2_X1 U5195 ( .A1(n4674), .A2(n5029), .ZN(U3313) );
  INV_X1 U5196 ( .A(D_REG_8__SCAN_IN), .ZN(n5015) );
  NOR2_X1 U5197 ( .A1(n4674), .A2(n5015), .ZN(U3314) );
  INV_X1 U5198 ( .A(D_REG_7__SCAN_IN), .ZN(n4672) );
  NOR2_X1 U5199 ( .A1(n4674), .A2(n4672), .ZN(U3315) );
  INV_X1 U5200 ( .A(D_REG_6__SCAN_IN), .ZN(n5007) );
  NOR2_X1 U5201 ( .A1(n4674), .A2(n5007), .ZN(U3316) );
  INV_X1 U5202 ( .A(D_REG_5__SCAN_IN), .ZN(n5016) );
  NOR2_X1 U5203 ( .A1(n4674), .A2(n5016), .ZN(U3317) );
  INV_X1 U5204 ( .A(D_REG_4__SCAN_IN), .ZN(n4673) );
  NOR2_X1 U5205 ( .A1(n4674), .A2(n4673), .ZN(U3318) );
  INV_X1 U5206 ( .A(D_REG_3__SCAN_IN), .ZN(n4857) );
  NOR2_X1 U5207 ( .A1(n4674), .A2(n4857), .ZN(U3319) );
  INV_X1 U5208 ( .A(D_REG_2__SCAN_IN), .ZN(n4817) );
  NOR2_X1 U5209 ( .A1(n4674), .A2(n4817), .ZN(U3320) );
  INV_X1 U5210 ( .A(DATAI_23_), .ZN(n4881) );
  AOI21_X1 U5211 ( .B1(U3149), .B2(n4881), .A(n4675), .ZN(U3329) );
  INV_X1 U5212 ( .A(DATAI_18_), .ZN(n5058) );
  AOI22_X1 U5213 ( .A1(STATE_REG_SCAN_IN), .A2(n4676), .B1(n5058), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5214 ( .A1(STATE_REG_SCAN_IN), .A2(n4677), .B1(n2675), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5215 ( .A(DATAI_16_), .ZN(n4862) );
  AOI22_X1 U5216 ( .A1(STATE_REG_SCAN_IN), .A2(n4678), .B1(n4862), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5217 ( .A(DATAI_15_), .ZN(n5066) );
  AOI22_X1 U5218 ( .A1(STATE_REG_SCAN_IN), .A2(n4679), .B1(n5066), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5219 ( .A(DATAI_14_), .ZN(n4680) );
  AOI22_X1 U5220 ( .A1(STATE_REG_SCAN_IN), .A2(n2368), .B1(n4680), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5221 ( .A1(STATE_REG_SCAN_IN), .A2(n4681), .B1(n2648), .B2(U3149), 
        .ZN(U3339) );
  AOI22_X1 U5222 ( .A1(STATE_REG_SCAN_IN), .A2(n4037), .B1(n4861), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5223 ( .A(DATAI_11_), .ZN(n5044) );
  AOI22_X1 U5224 ( .A1(STATE_REG_SCAN_IN), .A2(n4682), .B1(n5044), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5225 ( .A(DATAI_10_), .ZN(n4683) );
  AOI22_X1 U5226 ( .A1(STATE_REG_SCAN_IN), .A2(n2359), .B1(n4683), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5227 ( .A(DATAI_9_), .ZN(n5005) );
  AOI22_X1 U5228 ( .A1(STATE_REG_SCAN_IN), .A2(n4684), .B1(n5005), .B2(U3149), 
        .ZN(U3343) );
  AOI22_X1 U5229 ( .A1(STATE_REG_SCAN_IN), .A2(n4685), .B1(n5055), .B2(U3149), 
        .ZN(U3344) );
  AOI211_X1 U5230 ( .C1(n4697), .C2(n4688), .A(n4687), .B(n4686), .ZN(n4714)
         );
  INV_X1 U5231 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4773) );
  AOI22_X1 U5232 ( .A1(n4713), .A2(n4714), .B1(n4773), .B2(n4711), .ZN(U3467)
         );
  OAI22_X1 U5233 ( .A1(n4691), .A2(n4705), .B1(n4690), .B2(n4689), .ZN(n4692)
         );
  NOR2_X1 U5234 ( .A1(n4693), .A2(n4692), .ZN(n4715) );
  INV_X1 U5235 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4694) );
  AOI22_X1 U5236 ( .A1(n4713), .A2(n4715), .B1(n4694), .B2(n4711), .ZN(U3469)
         );
  AOI211_X1 U5237 ( .C1(n4698), .C2(n4697), .A(n4696), .B(n4695), .ZN(n4717)
         );
  INV_X1 U5238 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4996) );
  AOI22_X1 U5239 ( .A1(n4713), .A2(n4717), .B1(n4996), .B2(n4711), .ZN(U3475)
         );
  NOR2_X1 U5240 ( .A1(n4700), .A2(n4699), .ZN(n4704) );
  AOI211_X1 U5241 ( .C1(n4704), .C2(n4703), .A(n4702), .B(n4701), .ZN(n4718)
         );
  INV_X1 U5242 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4871) );
  AOI22_X1 U5243 ( .A1(n4713), .A2(n4718), .B1(n4871), .B2(n4711), .ZN(U3481)
         );
  NOR2_X1 U5244 ( .A1(n4706), .A2(n4705), .ZN(n4708) );
  AOI211_X1 U5245 ( .C1(n4710), .C2(n4709), .A(n4708), .B(n4707), .ZN(n4721)
         );
  INV_X1 U5246 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4712) );
  AOI22_X1 U5247 ( .A1(n4713), .A2(n4721), .B1(n4712), .B2(n4711), .ZN(U3489)
         );
  AOI22_X1 U5248 ( .A1(n4722), .A2(n4714), .B1(n2867), .B2(n4719), .ZN(U3518)
         );
  AOI22_X1 U5249 ( .A1(n4722), .A2(n4715), .B1(n3153), .B2(n4719), .ZN(U3519)
         );
  INV_X1 U5250 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4716) );
  AOI22_X1 U5251 ( .A1(n4722), .A2(n4717), .B1(n4716), .B2(n4719), .ZN(U3522)
         );
  AOI22_X1 U5252 ( .A1(n4722), .A2(n4718), .B1(n4028), .B2(n4719), .ZN(U3525)
         );
  AOI22_X1 U5253 ( .A1(n4722), .A2(n4721), .B1(n4720), .B2(n4719), .ZN(U3529)
         );
  OAI22_X1 U5254 ( .A1(IR_REG_19__SCAN_IN), .A2(keyinput_g74), .B1(DATAI_24_), 
        .B2(keyinput_g7), .ZN(n4723) );
  AOI221_X1 U5255 ( .B1(IR_REG_19__SCAN_IN), .B2(keyinput_g74), .C1(
        keyinput_g7), .C2(DATAI_24_), .A(n4723), .ZN(n4730) );
  OAI22_X1 U5256 ( .A1(D_REG_13__SCAN_IN), .A2(keyinput_g100), .B1(keyinput_g5), .B2(DATAI_26_), .ZN(n4724) );
  AOI221_X1 U5257 ( .B1(D_REG_13__SCAN_IN), .B2(keyinput_g100), .C1(DATAI_26_), 
        .C2(keyinput_g5), .A(n4724), .ZN(n4729) );
  OAI22_X1 U5258 ( .A1(D_REG_4__SCAN_IN), .A2(keyinput_g91), .B1(
        REG0_REG_6__SCAN_IN), .B2(keyinput_g125), .ZN(n4725) );
  AOI221_X1 U5259 ( .B1(D_REG_4__SCAN_IN), .B2(keyinput_g91), .C1(
        keyinput_g125), .C2(REG0_REG_6__SCAN_IN), .A(n4725), .ZN(n4728) );
  OAI22_X1 U5260 ( .A1(IR_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(
        REG0_REG_4__SCAN_IN), .B2(keyinput_g123), .ZN(n4726) );
  AOI221_X1 U5261 ( .B1(IR_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(
        keyinput_g123), .C2(REG0_REG_4__SCAN_IN), .A(n4726), .ZN(n4727) );
  NAND4_X1 U5262 ( .A1(n4730), .A2(n4729), .A3(n4728), .A4(n4727), .ZN(n4758)
         );
  OAI22_X1 U5263 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput_g51), .B1(DATAI_27_), 
        .B2(keyinput_g4), .ZN(n4731) );
  AOI221_X1 U5264 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput_g51), .C1(
        keyinput_g4), .C2(DATAI_27_), .A(n4731), .ZN(n4738) );
  OAI22_X1 U5265 ( .A1(REG3_REG_21__SCAN_IN), .A2(keyinput_g43), .B1(
        keyinput_g11), .B2(DATAI_20_), .ZN(n4732) );
  AOI221_X1 U5266 ( .B1(REG3_REG_21__SCAN_IN), .B2(keyinput_g43), .C1(
        DATAI_20_), .C2(keyinput_g11), .A(n4732), .ZN(n4737) );
  OAI22_X1 U5267 ( .A1(D_REG_28__SCAN_IN), .A2(keyinput_g115), .B1(
        keyinput_g38), .B2(REG3_REG_3__SCAN_IN), .ZN(n4733) );
  AOI221_X1 U5268 ( .B1(D_REG_28__SCAN_IN), .B2(keyinput_g115), .C1(
        REG3_REG_3__SCAN_IN), .C2(keyinput_g38), .A(n4733), .ZN(n4736) );
  OAI22_X1 U5269 ( .A1(IR_REG_15__SCAN_IN), .A2(keyinput_g70), .B1(
        keyinput_g110), .B2(D_REG_23__SCAN_IN), .ZN(n4734) );
  AOI221_X1 U5270 ( .B1(IR_REG_15__SCAN_IN), .B2(keyinput_g70), .C1(
        D_REG_23__SCAN_IN), .C2(keyinput_g110), .A(n4734), .ZN(n4735) );
  NAND4_X1 U5271 ( .A1(n4738), .A2(n4737), .A3(n4736), .A4(n4735), .ZN(n4757)
         );
  OAI22_X1 U5272 ( .A1(DATAI_6_), .A2(keyinput_g25), .B1(REG0_REG_1__SCAN_IN), 
        .B2(keyinput_g120), .ZN(n4739) );
  AOI221_X1 U5273 ( .B1(DATAI_6_), .B2(keyinput_g25), .C1(keyinput_g120), .C2(
        REG0_REG_1__SCAN_IN), .A(n4739), .ZN(n4746) );
  OAI22_X1 U5274 ( .A1(REG3_REG_13__SCAN_IN), .A2(keyinput_g54), .B1(
        keyinput_g127), .B2(REG0_REG_8__SCAN_IN), .ZN(n4740) );
  AOI221_X1 U5275 ( .B1(REG3_REG_13__SCAN_IN), .B2(keyinput_g54), .C1(
        REG0_REG_8__SCAN_IN), .C2(keyinput_g127), .A(n4740), .ZN(n4745) );
  OAI22_X1 U5276 ( .A1(REG3_REG_7__SCAN_IN), .A2(keyinput_g33), .B1(
        keyinput_g18), .B2(DATAI_13_), .ZN(n4741) );
  AOI221_X1 U5277 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput_g33), .C1(DATAI_13_), .C2(keyinput_g18), .A(n4741), .ZN(n4744) );
  OAI22_X1 U5278 ( .A1(IR_REG_8__SCAN_IN), .A2(keyinput_g63), .B1(keyinput_g56), .B2(IR_REG_1__SCAN_IN), .ZN(n4742) );
  AOI221_X1 U5279 ( .B1(IR_REG_8__SCAN_IN), .B2(keyinput_g63), .C1(
        IR_REG_1__SCAN_IN), .C2(keyinput_g56), .A(n4742), .ZN(n4743) );
  NAND4_X1 U5280 ( .A1(n4746), .A2(n4745), .A3(n4744), .A4(n4743), .ZN(n4756)
         );
  OAI22_X1 U5281 ( .A1(D_REG_22__SCAN_IN), .A2(keyinput_g109), .B1(
        D_REG_12__SCAN_IN), .B2(keyinput_g99), .ZN(n4747) );
  AOI221_X1 U5282 ( .B1(D_REG_22__SCAN_IN), .B2(keyinput_g109), .C1(
        keyinput_g99), .C2(D_REG_12__SCAN_IN), .A(n4747), .ZN(n4754) );
  OAI22_X1 U5283 ( .A1(D_REG_17__SCAN_IN), .A2(keyinput_g104), .B1(
        REG3_REG_25__SCAN_IN), .B2(keyinput_g45), .ZN(n4748) );
  AOI221_X1 U5284 ( .B1(D_REG_17__SCAN_IN), .B2(keyinput_g104), .C1(
        keyinput_g45), .C2(REG3_REG_25__SCAN_IN), .A(n4748), .ZN(n4753) );
  OAI22_X1 U5285 ( .A1(IR_REG_25__SCAN_IN), .A2(keyinput_g80), .B1(
        keyinput_g75), .B2(IR_REG_20__SCAN_IN), .ZN(n4749) );
  AOI221_X1 U5286 ( .B1(IR_REG_25__SCAN_IN), .B2(keyinput_g80), .C1(
        IR_REG_20__SCAN_IN), .C2(keyinput_g75), .A(n4749), .ZN(n4752) );
  OAI22_X1 U5287 ( .A1(IR_REG_23__SCAN_IN), .A2(keyinput_g78), .B1(
        IR_REG_9__SCAN_IN), .B2(keyinput_g64), .ZN(n4750) );
  AOI221_X1 U5288 ( .B1(IR_REG_23__SCAN_IN), .B2(keyinput_g78), .C1(
        keyinput_g64), .C2(IR_REG_9__SCAN_IN), .A(n4750), .ZN(n4751) );
  NAND4_X1 U5289 ( .A1(n4754), .A2(n4753), .A3(n4752), .A4(n4751), .ZN(n4755)
         );
  NOR4_X1 U5290 ( .A1(n4758), .A2(n4757), .A3(n4756), .A4(n4755), .ZN(n5089)
         );
  OAI22_X1 U5291 ( .A1(IR_REG_24__SCAN_IN), .A2(keyinput_g79), .B1(
        keyinput_g17), .B2(DATAI_14_), .ZN(n4759) );
  AOI221_X1 U5292 ( .B1(IR_REG_24__SCAN_IN), .B2(keyinput_g79), .C1(DATAI_14_), 
        .C2(keyinput_g17), .A(n4759), .ZN(n4766) );
  OAI22_X1 U5293 ( .A1(IR_REG_27__SCAN_IN), .A2(keyinput_g82), .B1(keyinput_g2), .B2(DATAI_29_), .ZN(n4760) );
  AOI221_X1 U5294 ( .B1(IR_REG_27__SCAN_IN), .B2(keyinput_g82), .C1(DATAI_29_), 
        .C2(keyinput_g2), .A(n4760), .ZN(n4765) );
  OAI22_X1 U5295 ( .A1(D_REG_15__SCAN_IN), .A2(keyinput_g102), .B1(
        IR_REG_30__SCAN_IN), .B2(keyinput_g85), .ZN(n4761) );
  AOI221_X1 U5296 ( .B1(D_REG_15__SCAN_IN), .B2(keyinput_g102), .C1(
        keyinput_g85), .C2(IR_REG_30__SCAN_IN), .A(n4761), .ZN(n4764) );
  OAI22_X1 U5297 ( .A1(IR_REG_31__SCAN_IN), .A2(keyinput_g86), .B1(
        REG0_REG_5__SCAN_IN), .B2(keyinput_g124), .ZN(n4762) );
  AOI221_X1 U5298 ( .B1(IR_REG_31__SCAN_IN), .B2(keyinput_g86), .C1(
        keyinput_g124), .C2(REG0_REG_5__SCAN_IN), .A(n4762), .ZN(n4763) );
  NAND4_X1 U5299 ( .A1(n4766), .A2(n4765), .A3(n4764), .A4(n4763), .ZN(n4898)
         );
  OAI22_X1 U5300 ( .A1(IR_REG_17__SCAN_IN), .A2(keyinput_g72), .B1(keyinput_g0), .B2(DATAI_31_), .ZN(n4767) );
  AOI221_X1 U5301 ( .B1(IR_REG_17__SCAN_IN), .B2(keyinput_g72), .C1(DATAI_31_), 
        .C2(keyinput_g0), .A(n4767), .ZN(n4793) );
  OAI22_X1 U5302 ( .A1(DATAI_7_), .A2(keyinput_g24), .B1(keyinput_g26), .B2(
        DATAI_5_), .ZN(n4768) );
  AOI221_X1 U5303 ( .B1(DATAI_7_), .B2(keyinput_g24), .C1(DATAI_5_), .C2(
        keyinput_g26), .A(n4768), .ZN(n4771) );
  OAI22_X1 U5304 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput_g46), .B1(
        keyinput_g21), .B2(DATAI_10_), .ZN(n4769) );
  AOI221_X1 U5305 ( .B1(REG3_REG_16__SCAN_IN), .B2(keyinput_g46), .C1(
        DATAI_10_), .C2(keyinput_g21), .A(n4769), .ZN(n4770) );
  OAI211_X1 U5306 ( .C1(n4773), .C2(keyinput_g119), .A(n4771), .B(n4770), .ZN(
        n4772) );
  AOI21_X1 U5307 ( .B1(n4773), .B2(keyinput_g119), .A(n4772), .ZN(n4792) );
  AOI22_X1 U5308 ( .A1(DATAI_19_), .A2(keyinput_g12), .B1(IR_REG_4__SCAN_IN), 
        .B2(keyinput_g59), .ZN(n4774) );
  OAI221_X1 U5309 ( .B1(DATAI_19_), .B2(keyinput_g12), .C1(IR_REG_4__SCAN_IN), 
        .C2(keyinput_g59), .A(n4774), .ZN(n4781) );
  AOI22_X1 U5310 ( .A1(REG3_REG_24__SCAN_IN), .A2(keyinput_g49), .B1(
        REG3_REG_27__SCAN_IN), .B2(keyinput_g34), .ZN(n4775) );
  OAI221_X1 U5311 ( .B1(REG3_REG_24__SCAN_IN), .B2(keyinput_g49), .C1(
        REG3_REG_27__SCAN_IN), .C2(keyinput_g34), .A(n4775), .ZN(n4780) );
  AOI22_X1 U5312 ( .A1(D_REG_25__SCAN_IN), .A2(keyinput_g112), .B1(
        D_REG_30__SCAN_IN), .B2(keyinput_g117), .ZN(n4776) );
  OAI221_X1 U5313 ( .B1(D_REG_25__SCAN_IN), .B2(keyinput_g112), .C1(
        D_REG_30__SCAN_IN), .C2(keyinput_g117), .A(n4776), .ZN(n4779) );
  AOI22_X1 U5314 ( .A1(D_REG_7__SCAN_IN), .A2(keyinput_g94), .B1(
        D_REG_16__SCAN_IN), .B2(keyinput_g103), .ZN(n4777) );
  OAI221_X1 U5315 ( .B1(D_REG_7__SCAN_IN), .B2(keyinput_g94), .C1(
        D_REG_16__SCAN_IN), .C2(keyinput_g103), .A(n4777), .ZN(n4778) );
  NOR4_X1 U5316 ( .A1(n4781), .A2(n4780), .A3(n4779), .A4(n4778), .ZN(n4791)
         );
  AOI22_X1 U5317 ( .A1(IR_REG_10__SCAN_IN), .A2(keyinput_g65), .B1(
        IR_REG_14__SCAN_IN), .B2(keyinput_g69), .ZN(n4782) );
  OAI221_X1 U5318 ( .B1(IR_REG_10__SCAN_IN), .B2(keyinput_g65), .C1(
        IR_REG_14__SCAN_IN), .C2(keyinput_g69), .A(n4782), .ZN(n4789) );
  AOI22_X1 U5319 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_g42), .B1(
        REG3_REG_17__SCAN_IN), .B2(keyinput_g48), .ZN(n4783) );
  OAI221_X1 U5320 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_g42), .C1(
        REG3_REG_17__SCAN_IN), .C2(keyinput_g48), .A(n4783), .ZN(n4788) );
  AOI22_X1 U5321 ( .A1(IR_REG_3__SCAN_IN), .A2(keyinput_g58), .B1(
        IR_REG_5__SCAN_IN), .B2(keyinput_g60), .ZN(n4784) );
  OAI221_X1 U5322 ( .B1(IR_REG_3__SCAN_IN), .B2(keyinput_g58), .C1(
        IR_REG_5__SCAN_IN), .C2(keyinput_g60), .A(n4784), .ZN(n4787) );
  AOI22_X1 U5323 ( .A1(DATAI_1_), .A2(keyinput_g30), .B1(REG3_REG_8__SCAN_IN), 
        .B2(keyinput_g41), .ZN(n4785) );
  OAI221_X1 U5324 ( .B1(DATAI_1_), .B2(keyinput_g30), .C1(REG3_REG_8__SCAN_IN), 
        .C2(keyinput_g41), .A(n4785), .ZN(n4786) );
  NOR4_X1 U5325 ( .A1(n4789), .A2(n4788), .A3(n4787), .A4(n4786), .ZN(n4790)
         );
  NAND4_X1 U5326 ( .A1(n4793), .A2(n4792), .A3(n4791), .A4(n4790), .ZN(n4897)
         );
  AOI22_X1 U5327 ( .A1(DATAI_4_), .A2(keyinput_g27), .B1(IR_REG_13__SCAN_IN), 
        .B2(keyinput_g68), .ZN(n4794) );
  OAI221_X1 U5328 ( .B1(DATAI_4_), .B2(keyinput_g27), .C1(IR_REG_13__SCAN_IN), 
        .C2(keyinput_g68), .A(n4794), .ZN(n4798) );
  AOI22_X1 U5329 ( .A1(D_REG_21__SCAN_IN), .A2(keyinput_g108), .B1(
        D_REG_1__SCAN_IN), .B2(keyinput_g88), .ZN(n4795) );
  OAI221_X1 U5330 ( .B1(D_REG_21__SCAN_IN), .B2(keyinput_g108), .C1(
        D_REG_1__SCAN_IN), .C2(keyinput_g88), .A(n4795), .ZN(n4797) );
  XOR2_X1 U5331 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_g52), .Z(n4796) );
  OR3_X1 U5332 ( .A1(n4798), .A2(n4797), .A3(n4796), .ZN(n4803) );
  AOI22_X1 U5333 ( .A1(n5066), .A2(keyinput_g16), .B1(n5032), .B2(
        keyinput_g101), .ZN(n4799) );
  OAI221_X1 U5334 ( .B1(n5066), .B2(keyinput_g16), .C1(n5032), .C2(
        keyinput_g101), .A(n4799), .ZN(n4802) );
  XNOR2_X1 U5335 ( .A(n4800), .B(keyinput_g107), .ZN(n4801) );
  NOR3_X1 U5336 ( .A1(n4803), .A2(n4802), .A3(n4801), .ZN(n4843) );
  AOI22_X1 U5337 ( .A1(n4805), .A2(keyinput_g3), .B1(n5034), .B2(keyinput_g111), .ZN(n4804) );
  OAI221_X1 U5338 ( .B1(n4805), .B2(keyinput_g3), .C1(n5034), .C2(
        keyinput_g111), .A(n4804), .ZN(n4815) );
  AOI22_X1 U5339 ( .A1(n4807), .A2(keyinput_g44), .B1(n5043), .B2(keyinput_g39), .ZN(n4806) );
  OAI221_X1 U5340 ( .B1(n4807), .B2(keyinput_g44), .C1(n5043), .C2(
        keyinput_g39), .A(n4806), .ZN(n4814) );
  XNOR2_X1 U5341 ( .A(n4808), .B(keyinput_g113), .ZN(n4813) );
  XNOR2_X1 U5342 ( .A(IR_REG_16__SCAN_IN), .B(keyinput_g71), .ZN(n4811) );
  XNOR2_X1 U5343 ( .A(IR_REG_11__SCAN_IN), .B(keyinput_g66), .ZN(n4810) );
  XNOR2_X1 U5344 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_g67), .ZN(n4809) );
  NAND3_X1 U5345 ( .A1(n4811), .A2(n4810), .A3(n4809), .ZN(n4812) );
  NOR4_X1 U5346 ( .A1(n4815), .A2(n4814), .A3(n4813), .A4(n4812), .ZN(n4842)
         );
  INV_X1 U5347 ( .A(DATAI_0_), .ZN(n4818) );
  AOI22_X1 U5348 ( .A1(n4818), .A2(keyinput_g31), .B1(n4817), .B2(keyinput_g89), .ZN(n4816) );
  OAI221_X1 U5349 ( .B1(n4818), .B2(keyinput_g31), .C1(n4817), .C2(
        keyinput_g89), .A(n4816), .ZN(n4827) );
  XNOR2_X1 U5350 ( .A(n4819), .B(keyinput_g116), .ZN(n4826) );
  XNOR2_X1 U5351 ( .A(n5035), .B(keyinput_g97), .ZN(n4825) );
  XOR2_X1 U5352 ( .A(n2763), .B(keyinput_g40), .Z(n4823) );
  XNOR2_X1 U5353 ( .A(IR_REG_28__SCAN_IN), .B(keyinput_g83), .ZN(n4822) );
  XNOR2_X1 U5354 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_g73), .ZN(n4821) );
  XNOR2_X1 U5355 ( .A(DATAI_2_), .B(keyinput_g29), .ZN(n4820) );
  NAND4_X1 U5356 ( .A1(n4823), .A2(n4822), .A3(n4821), .A4(n4820), .ZN(n4824)
         );
  NOR4_X1 U5357 ( .A1(n4827), .A2(n4826), .A3(n4825), .A4(n4824), .ZN(n4841)
         );
  INV_X1 U5358 ( .A(IR_REG_29__SCAN_IN), .ZN(n4829) );
  AOI22_X1 U5359 ( .A1(n4829), .A2(keyinput_g84), .B1(n5016), .B2(keyinput_g92), .ZN(n4828) );
  OAI221_X1 U5360 ( .B1(n4829), .B2(keyinput_g84), .C1(n5016), .C2(
        keyinput_g92), .A(n4828), .ZN(n4839) );
  INV_X1 U5361 ( .A(DATAI_22_), .ZN(n4831) );
  INV_X1 U5362 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4992) );
  AOI22_X1 U5363 ( .A1(n4831), .A2(keyinput_g9), .B1(keyinput_g122), .B2(n4992), .ZN(n4830) );
  OAI221_X1 U5364 ( .B1(n4831), .B2(keyinput_g9), .C1(n4992), .C2(
        keyinput_g122), .A(n4830), .ZN(n4838) );
  INV_X1 U5365 ( .A(DATAI_30_), .ZN(n4833) );
  AOI22_X1 U5366 ( .A1(n5012), .A2(keyinput_g98), .B1(keyinput_g1), .B2(n4833), 
        .ZN(n4832) );
  OAI221_X1 U5367 ( .B1(n5012), .B2(keyinput_g98), .C1(n4833), .C2(keyinput_g1), .A(n4832), .ZN(n4837) );
  AOI22_X1 U5368 ( .A1(n4835), .A2(keyinput_g10), .B1(keyinput_g22), .B2(n5005), .ZN(n4834) );
  OAI221_X1 U5369 ( .B1(n4835), .B2(keyinput_g10), .C1(n5005), .C2(
        keyinput_g22), .A(n4834), .ZN(n4836) );
  NOR4_X1 U5370 ( .A1(n4839), .A2(n4838), .A3(n4837), .A4(n4836), .ZN(n4840)
         );
  NAND4_X1 U5371 ( .A1(n4843), .A2(n4842), .A3(n4841), .A4(n4840), .ZN(n4896)
         );
  AOI22_X1 U5372 ( .A1(n2809), .A2(keyinput_g87), .B1(keyinput_g6), .B2(n4974), 
        .ZN(n4844) );
  OAI221_X1 U5373 ( .B1(n2809), .B2(keyinput_g87), .C1(n4974), .C2(keyinput_g6), .A(n4844), .ZN(n4854) );
  AOI22_X1 U5374 ( .A1(n5007), .A2(keyinput_g93), .B1(keyinput_g14), .B2(n2675), .ZN(n4845) );
  OAI221_X1 U5375 ( .B1(n5007), .B2(keyinput_g93), .C1(n2675), .C2(
        keyinput_g14), .A(n4845), .ZN(n4853) );
  AOI22_X1 U5376 ( .A1(n4848), .A2(keyinput_g37), .B1(n4847), .B2(keyinput_g35), .ZN(n4846) );
  OAI221_X1 U5377 ( .B1(n4848), .B2(keyinput_g37), .C1(n4847), .C2(
        keyinput_g35), .A(n4846), .ZN(n4852) );
  XOR2_X1 U5378 ( .A(n4986), .B(keyinput_g55), .Z(n4850) );
  XNOR2_X1 U5379 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_g76), .ZN(n4849) );
  NAND2_X1 U5380 ( .A1(n4850), .A2(n4849), .ZN(n4851) );
  NOR4_X1 U5381 ( .A1(n4854), .A2(n4853), .A3(n4852), .A4(n4851), .ZN(n4894)
         );
  INV_X1 U5382 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4856) );
  AOI22_X1 U5383 ( .A1(n4857), .A2(keyinput_g90), .B1(keyinput_g53), .B2(n4856), .ZN(n4855) );
  OAI221_X1 U5384 ( .B1(n4857), .B2(keyinput_g90), .C1(n4856), .C2(
        keyinput_g53), .A(n4855), .ZN(n4868) );
  AOI22_X1 U5385 ( .A1(n5026), .A2(keyinput_g106), .B1(n4859), .B2(
        keyinput_g118), .ZN(n4858) );
  OAI221_X1 U5386 ( .B1(n5026), .B2(keyinput_g106), .C1(n4859), .C2(
        keyinput_g118), .A(n4858), .ZN(n4867) );
  AOI22_X1 U5387 ( .A1(n4862), .A2(keyinput_g15), .B1(keyinput_g19), .B2(n4861), .ZN(n4860) );
  OAI221_X1 U5388 ( .B1(n4862), .B2(keyinput_g15), .C1(n4861), .C2(
        keyinput_g19), .A(n4860), .ZN(n4866) );
  AOI22_X1 U5389 ( .A1(n4864), .A2(keyinput_g36), .B1(keyinput_g47), .B2(n4995), .ZN(n4863) );
  OAI221_X1 U5390 ( .B1(n4864), .B2(keyinput_g36), .C1(n4995), .C2(
        keyinput_g47), .A(n4863), .ZN(n4865) );
  NOR4_X1 U5391 ( .A1(n4868), .A2(n4867), .A3(n4866), .A4(n4865), .ZN(n4893)
         );
  AOI22_X1 U5392 ( .A1(n2462), .A2(keyinput_g57), .B1(n2579), .B2(keyinput_g62), .ZN(n4869) );
  OAI221_X1 U5393 ( .B1(n2462), .B2(keyinput_g57), .C1(n2579), .C2(
        keyinput_g62), .A(n4869), .ZN(n4878) );
  AOI22_X1 U5394 ( .A1(n5058), .A2(keyinput_g13), .B1(n4871), .B2(
        keyinput_g126), .ZN(n4870) );
  OAI221_X1 U5395 ( .B1(n5058), .B2(keyinput_g13), .C1(n4871), .C2(
        keyinput_g126), .A(n4870), .ZN(n4877) );
  INV_X1 U5396 ( .A(REG0_REG_2__SCAN_IN), .ZN(n5054) );
  AOI22_X1 U5397 ( .A1(n5054), .A2(keyinput_g121), .B1(n5055), .B2(
        keyinput_g23), .ZN(n4872) );
  OAI221_X1 U5398 ( .B1(n5054), .B2(keyinput_g121), .C1(n5055), .C2(
        keyinput_g23), .A(n4872), .ZN(n4876) );
  XNOR2_X1 U5399 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_g50), .ZN(n4874) );
  XNOR2_X1 U5400 ( .A(STATE_REG_SCAN_IN), .B(keyinput_g32), .ZN(n4873) );
  NAND2_X1 U5401 ( .A1(n4874), .A2(n4873), .ZN(n4875) );
  NOR4_X1 U5402 ( .A1(n4878), .A2(n4877), .A3(n4876), .A4(n4875), .ZN(n4892)
         );
  AOI22_X1 U5403 ( .A1(n5044), .A2(keyinput_g20), .B1(n5015), .B2(keyinput_g95), .ZN(n4879) );
  OAI221_X1 U5404 ( .B1(n5044), .B2(keyinput_g20), .C1(n5015), .C2(
        keyinput_g95), .A(n4879), .ZN(n4890) );
  AOI22_X1 U5405 ( .A1(n4882), .A2(keyinput_g114), .B1(keyinput_g8), .B2(n4881), .ZN(n4880) );
  OAI221_X1 U5406 ( .B1(n4882), .B2(keyinput_g114), .C1(n4881), .C2(
        keyinput_g8), .A(n4880), .ZN(n4889) );
  INV_X1 U5407 ( .A(DATAI_3_), .ZN(n4884) );
  AOI22_X1 U5408 ( .A1(n4884), .A2(keyinput_g28), .B1(n5029), .B2(keyinput_g96), .ZN(n4883) );
  OAI221_X1 U5409 ( .B1(n4884), .B2(keyinput_g28), .C1(n5029), .C2(
        keyinput_g96), .A(n4883), .ZN(n4888) );
  INV_X1 U5410 ( .A(IR_REG_22__SCAN_IN), .ZN(n4886) );
  AOI22_X1 U5411 ( .A1(n5025), .A2(keyinput_g105), .B1(n4886), .B2(
        keyinput_g77), .ZN(n4885) );
  OAI221_X1 U5412 ( .B1(n5025), .B2(keyinput_g105), .C1(n4886), .C2(
        keyinput_g77), .A(n4885), .ZN(n4887) );
  NOR4_X1 U5413 ( .A1(n4890), .A2(n4889), .A3(n4888), .A4(n4887), .ZN(n4891)
         );
  NAND4_X1 U5414 ( .A1(n4894), .A2(n4893), .A3(n4892), .A4(n4891), .ZN(n4895)
         );
  NOR4_X1 U5415 ( .A1(n4898), .A2(n4897), .A3(n4896), .A4(n4895), .ZN(n5088)
         );
  XOR2_X1 U5416 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_f67), .Z(n4905) );
  AOI22_X1 U5417 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput_f52), .B1(DATAI_29_), 
        .B2(keyinput_f2), .ZN(n4899) );
  OAI221_X1 U5418 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput_f52), .C1(DATAI_29_), .C2(keyinput_f2), .A(n4899), .ZN(n4904) );
  AOI22_X1 U5419 ( .A1(DATAI_20_), .A2(keyinput_f11), .B1(REG3_REG_28__SCAN_IN), .B2(keyinput_f40), .ZN(n4900) );
  OAI221_X1 U5420 ( .B1(DATAI_20_), .B2(keyinput_f11), .C1(
        REG3_REG_28__SCAN_IN), .C2(keyinput_f40), .A(n4900), .ZN(n4903) );
  AOI22_X1 U5421 ( .A1(DATAI_31_), .A2(keyinput_f0), .B1(REG3_REG_21__SCAN_IN), 
        .B2(keyinput_f43), .ZN(n4901) );
  OAI221_X1 U5422 ( .B1(DATAI_31_), .B2(keyinput_f0), .C1(REG3_REG_21__SCAN_IN), .C2(keyinput_f43), .A(n4901), .ZN(n4902) );
  NOR4_X1 U5423 ( .A1(n4905), .A2(n4904), .A3(n4903), .A4(n4902), .ZN(n4933)
         );
  AOI22_X1 U5424 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(DATAI_26_), .B2(
        keyinput_f5), .ZN(n4906) );
  OAI221_X1 U5425 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(DATAI_26_), .C2(
        keyinput_f5), .A(n4906), .ZN(n4913) );
  AOI22_X1 U5426 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_f42), .B1(DATAI_21_), 
        .B2(keyinput_f10), .ZN(n4907) );
  OAI221_X1 U5427 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_f42), .C1(DATAI_21_), .C2(keyinput_f10), .A(n4907), .ZN(n4912) );
  AOI22_X1 U5428 ( .A1(REG3_REG_14__SCAN_IN), .A2(keyinput_f35), .B1(
        REG3_REG_17__SCAN_IN), .B2(keyinput_f48), .ZN(n4908) );
  OAI221_X1 U5429 ( .B1(REG3_REG_14__SCAN_IN), .B2(keyinput_f35), .C1(
        REG3_REG_17__SCAN_IN), .C2(keyinput_f48), .A(n4908), .ZN(n4911) );
  AOI22_X1 U5430 ( .A1(D_REG_28__SCAN_IN), .A2(keyinput_f115), .B1(
        D_REG_30__SCAN_IN), .B2(keyinput_f117), .ZN(n4909) );
  OAI221_X1 U5431 ( .B1(D_REG_28__SCAN_IN), .B2(keyinput_f115), .C1(
        D_REG_30__SCAN_IN), .C2(keyinput_f117), .A(n4909), .ZN(n4910) );
  NOR4_X1 U5432 ( .A1(n4913), .A2(n4912), .A3(n4911), .A4(n4910), .ZN(n4932)
         );
  AOI22_X1 U5433 ( .A1(D_REG_23__SCAN_IN), .A2(keyinput_f110), .B1(
        D_REG_25__SCAN_IN), .B2(keyinput_f112), .ZN(n4914) );
  OAI221_X1 U5434 ( .B1(D_REG_23__SCAN_IN), .B2(keyinput_f110), .C1(
        D_REG_25__SCAN_IN), .C2(keyinput_f112), .A(n4914), .ZN(n4921) );
  AOI22_X1 U5435 ( .A1(D_REG_16__SCAN_IN), .A2(keyinput_f103), .B1(
        D_REG_21__SCAN_IN), .B2(keyinput_f108), .ZN(n4915) );
  OAI221_X1 U5436 ( .B1(D_REG_16__SCAN_IN), .B2(keyinput_f103), .C1(
        D_REG_21__SCAN_IN), .C2(keyinput_f108), .A(n4915), .ZN(n4920) );
  AOI22_X1 U5437 ( .A1(D_REG_13__SCAN_IN), .A2(keyinput_f100), .B1(
        D_REG_15__SCAN_IN), .B2(keyinput_f102), .ZN(n4916) );
  OAI221_X1 U5438 ( .B1(D_REG_13__SCAN_IN), .B2(keyinput_f100), .C1(
        D_REG_15__SCAN_IN), .C2(keyinput_f102), .A(n4916), .ZN(n4919) );
  AOI22_X1 U5439 ( .A1(D_REG_4__SCAN_IN), .A2(keyinput_f91), .B1(
        D_REG_7__SCAN_IN), .B2(keyinput_f94), .ZN(n4917) );
  OAI221_X1 U5440 ( .B1(D_REG_4__SCAN_IN), .B2(keyinput_f91), .C1(
        D_REG_7__SCAN_IN), .C2(keyinput_f94), .A(n4917), .ZN(n4918) );
  NOR4_X1 U5441 ( .A1(n4921), .A2(n4920), .A3(n4919), .A4(n4918), .ZN(n4931)
         );
  AOI22_X1 U5442 ( .A1(IR_REG_30__SCAN_IN), .A2(keyinput_f85), .B1(
        IR_REG_17__SCAN_IN), .B2(keyinput_f72), .ZN(n4922) );
  OAI221_X1 U5443 ( .B1(IR_REG_30__SCAN_IN), .B2(keyinput_f85), .C1(
        IR_REG_17__SCAN_IN), .C2(keyinput_f72), .A(n4922), .ZN(n4929) );
  AOI22_X1 U5444 ( .A1(IR_REG_14__SCAN_IN), .A2(keyinput_f69), .B1(
        IR_REG_16__SCAN_IN), .B2(keyinput_f71), .ZN(n4923) );
  OAI221_X1 U5445 ( .B1(IR_REG_14__SCAN_IN), .B2(keyinput_f69), .C1(
        IR_REG_16__SCAN_IN), .C2(keyinput_f71), .A(n4923), .ZN(n4928) );
  AOI22_X1 U5446 ( .A1(DATAI_10_), .A2(keyinput_f21), .B1(IR_REG_15__SCAN_IN), 
        .B2(keyinput_f70), .ZN(n4924) );
  OAI221_X1 U5447 ( .B1(DATAI_10_), .B2(keyinput_f21), .C1(IR_REG_15__SCAN_IN), 
        .C2(keyinput_f70), .A(n4924), .ZN(n4927) );
  AOI22_X1 U5448 ( .A1(REG0_REG_1__SCAN_IN), .A2(keyinput_f120), .B1(DATAI_6_), 
        .B2(keyinput_f25), .ZN(n4925) );
  OAI221_X1 U5449 ( .B1(REG0_REG_1__SCAN_IN), .B2(keyinput_f120), .C1(DATAI_6_), .C2(keyinput_f25), .A(n4925), .ZN(n4926) );
  NOR4_X1 U5450 ( .A1(n4929), .A2(n4928), .A3(n4927), .A4(n4926), .ZN(n4930)
         );
  NAND4_X1 U5451 ( .A1(n4933), .A2(n4932), .A3(n4931), .A4(n4930), .ZN(n5082)
         );
  AOI22_X1 U5452 ( .A1(REG0_REG_5__SCAN_IN), .A2(keyinput_f124), .B1(
        REG0_REG_6__SCAN_IN), .B2(keyinput_f125), .ZN(n4934) );
  OAI221_X1 U5453 ( .B1(REG0_REG_5__SCAN_IN), .B2(keyinput_f124), .C1(
        REG0_REG_6__SCAN_IN), .C2(keyinput_f125), .A(n4934), .ZN(n4941) );
  AOI22_X1 U5454 ( .A1(REG0_REG_8__SCAN_IN), .A2(keyinput_f127), .B1(
        IR_REG_11__SCAN_IN), .B2(keyinput_f66), .ZN(n4935) );
  OAI221_X1 U5455 ( .B1(REG0_REG_8__SCAN_IN), .B2(keyinput_f127), .C1(
        IR_REG_11__SCAN_IN), .C2(keyinput_f66), .A(n4935), .ZN(n4940) );
  AOI22_X1 U5456 ( .A1(REG0_REG_7__SCAN_IN), .A2(keyinput_f126), .B1(
        IR_REG_10__SCAN_IN), .B2(keyinput_f65), .ZN(n4936) );
  OAI221_X1 U5457 ( .B1(REG0_REG_7__SCAN_IN), .B2(keyinput_f126), .C1(
        IR_REG_10__SCAN_IN), .C2(keyinput_f65), .A(n4936), .ZN(n4939) );
  AOI22_X1 U5458 ( .A1(IR_REG_5__SCAN_IN), .A2(keyinput_f60), .B1(
        IR_REG_6__SCAN_IN), .B2(keyinput_f61), .ZN(n4937) );
  OAI221_X1 U5459 ( .B1(IR_REG_5__SCAN_IN), .B2(keyinput_f60), .C1(
        IR_REG_6__SCAN_IN), .C2(keyinput_f61), .A(n4937), .ZN(n4938) );
  NOR4_X1 U5460 ( .A1(n4941), .A2(n4940), .A3(n4939), .A4(n4938), .ZN(n4969)
         );
  AOI22_X1 U5461 ( .A1(REG0_REG_0__SCAN_IN), .A2(keyinput_f119), .B1(
        REG3_REG_4__SCAN_IN), .B2(keyinput_f50), .ZN(n4942) );
  OAI221_X1 U5462 ( .B1(REG0_REG_0__SCAN_IN), .B2(keyinput_f119), .C1(
        REG3_REG_4__SCAN_IN), .C2(keyinput_f50), .A(n4942), .ZN(n4949) );
  AOI22_X1 U5463 ( .A1(IR_REG_1__SCAN_IN), .A2(keyinput_f56), .B1(
        IR_REG_8__SCAN_IN), .B2(keyinput_f63), .ZN(n4943) );
  OAI221_X1 U5464 ( .B1(IR_REG_1__SCAN_IN), .B2(keyinput_f56), .C1(
        IR_REG_8__SCAN_IN), .C2(keyinput_f63), .A(n4943), .ZN(n4948) );
  AOI22_X1 U5465 ( .A1(D_REG_3__SCAN_IN), .A2(keyinput_f90), .B1(
        D_REG_1__SCAN_IN), .B2(keyinput_f88), .ZN(n4944) );
  OAI221_X1 U5466 ( .B1(D_REG_3__SCAN_IN), .B2(keyinput_f90), .C1(
        D_REG_1__SCAN_IN), .C2(keyinput_f88), .A(n4944), .ZN(n4947) );
  AOI22_X1 U5467 ( .A1(D_REG_29__SCAN_IN), .A2(keyinput_f116), .B1(
        D_REG_31__SCAN_IN), .B2(keyinput_f118), .ZN(n4945) );
  OAI221_X1 U5468 ( .B1(D_REG_29__SCAN_IN), .B2(keyinput_f116), .C1(
        D_REG_31__SCAN_IN), .C2(keyinput_f118), .A(n4945), .ZN(n4946) );
  NOR4_X1 U5469 ( .A1(n4949), .A2(n4948), .A3(n4947), .A4(n4946), .ZN(n4968)
         );
  AOI22_X1 U5470 ( .A1(D_REG_2__SCAN_IN), .A2(keyinput_f89), .B1(
        D_REG_26__SCAN_IN), .B2(keyinput_f113), .ZN(n4950) );
  OAI221_X1 U5471 ( .B1(D_REG_2__SCAN_IN), .B2(keyinput_f89), .C1(
        D_REG_26__SCAN_IN), .C2(keyinput_f113), .A(n4950), .ZN(n4957) );
  AOI22_X1 U5472 ( .A1(D_REG_27__SCAN_IN), .A2(keyinput_f114), .B1(
        D_REG_20__SCAN_IN), .B2(keyinput_f107), .ZN(n4951) );
  OAI221_X1 U5473 ( .B1(D_REG_27__SCAN_IN), .B2(keyinput_f114), .C1(
        D_REG_20__SCAN_IN), .C2(keyinput_f107), .A(n4951), .ZN(n4956) );
  AOI22_X1 U5474 ( .A1(REG3_REG_8__SCAN_IN), .A2(keyinput_f41), .B1(
        REG3_REG_16__SCAN_IN), .B2(keyinput_f46), .ZN(n4952) );
  OAI221_X1 U5475 ( .B1(REG3_REG_8__SCAN_IN), .B2(keyinput_f41), .C1(
        REG3_REG_16__SCAN_IN), .C2(keyinput_f46), .A(n4952), .ZN(n4955) );
  AOI22_X1 U5476 ( .A1(DATAI_16_), .A2(keyinput_f15), .B1(IR_REG_29__SCAN_IN), 
        .B2(keyinput_f84), .ZN(n4953) );
  OAI221_X1 U5477 ( .B1(DATAI_16_), .B2(keyinput_f15), .C1(IR_REG_29__SCAN_IN), 
        .C2(keyinput_f84), .A(n4953), .ZN(n4954) );
  NOR4_X1 U5478 ( .A1(n4957), .A2(n4956), .A3(n4955), .A4(n4954), .ZN(n4967)
         );
  AOI22_X1 U5479 ( .A1(DATAI_12_), .A2(keyinput_f19), .B1(REG3_REG_23__SCAN_IN), .B2(keyinput_f36), .ZN(n4958) );
  OAI221_X1 U5480 ( .B1(DATAI_12_), .B2(keyinput_f19), .C1(
        REG3_REG_23__SCAN_IN), .C2(keyinput_f36), .A(n4958), .ZN(n4965) );
  AOI22_X1 U5481 ( .A1(DATAI_23_), .A2(keyinput_f8), .B1(IR_REG_2__SCAN_IN), 
        .B2(keyinput_f57), .ZN(n4959) );
  OAI221_X1 U5482 ( .B1(DATAI_23_), .B2(keyinput_f8), .C1(IR_REG_2__SCAN_IN), 
        .C2(keyinput_f57), .A(n4959), .ZN(n4964) );
  AOI22_X1 U5483 ( .A1(DATAI_3_), .A2(keyinput_f28), .B1(IR_REG_22__SCAN_IN), 
        .B2(keyinput_f77), .ZN(n4960) );
  OAI221_X1 U5484 ( .B1(DATAI_3_), .B2(keyinput_f28), .C1(IR_REG_22__SCAN_IN), 
        .C2(keyinput_f77), .A(n4960), .ZN(n4963) );
  AOI22_X1 U5485 ( .A1(DATAI_17_), .A2(keyinput_f14), .B1(REG3_REG_10__SCAN_IN), .B2(keyinput_f37), .ZN(n4961) );
  OAI221_X1 U5486 ( .B1(DATAI_17_), .B2(keyinput_f14), .C1(
        REG3_REG_10__SCAN_IN), .C2(keyinput_f37), .A(n4961), .ZN(n4962) );
  NOR4_X1 U5487 ( .A1(n4965), .A2(n4964), .A3(n4963), .A4(n4962), .ZN(n4966)
         );
  NAND4_X1 U5488 ( .A1(n4969), .A2(n4968), .A3(n4967), .A4(n4966), .ZN(n5081)
         );
  AOI22_X1 U5489 ( .A1(DATAI_22_), .A2(keyinput_f9), .B1(IR_REG_25__SCAN_IN), 
        .B2(keyinput_f80), .ZN(n4970) );
  OAI221_X1 U5490 ( .B1(DATAI_22_), .B2(keyinput_f9), .C1(IR_REG_25__SCAN_IN), 
        .C2(keyinput_f80), .A(n4970), .ZN(n4978) );
  AOI22_X1 U5491 ( .A1(DATAI_0_), .A2(keyinput_f31), .B1(IR_REG_28__SCAN_IN), 
        .B2(keyinput_f83), .ZN(n4971) );
  OAI221_X1 U5492 ( .B1(DATAI_0_), .B2(keyinput_f31), .C1(IR_REG_28__SCAN_IN), 
        .C2(keyinput_f83), .A(n4971), .ZN(n4977) );
  AOI22_X1 U5493 ( .A1(DATAI_28_), .A2(keyinput_f3), .B1(REG3_REG_12__SCAN_IN), 
        .B2(keyinput_f44), .ZN(n4972) );
  OAI221_X1 U5494 ( .B1(DATAI_28_), .B2(keyinput_f3), .C1(REG3_REG_12__SCAN_IN), .C2(keyinput_f44), .A(n4972), .ZN(n4976) );
  AOI22_X1 U5495 ( .A1(U3149), .A2(keyinput_f32), .B1(keyinput_f6), .B2(n4974), 
        .ZN(n4973) );
  OAI221_X1 U5496 ( .B1(U3149), .B2(keyinput_f32), .C1(n4974), .C2(keyinput_f6), .A(n4973), .ZN(n4975) );
  NOR4_X1 U5497 ( .A1(n4978), .A2(n4977), .A3(n4976), .A4(n4975), .ZN(n5023)
         );
  INV_X1 U5498 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4980) );
  AOI22_X1 U5499 ( .A1(n4981), .A2(keyinput_f34), .B1(keyinput_f49), .B2(n4980), .ZN(n4979) );
  OAI221_X1 U5500 ( .B1(n4981), .B2(keyinput_f34), .C1(n4980), .C2(
        keyinput_f49), .A(n4979), .ZN(n4990) );
  XNOR2_X1 U5501 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_f53), .ZN(n4985) );
  XNOR2_X1 U5502 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_f38), .ZN(n4984) );
  XNOR2_X1 U5503 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_f86), .ZN(n4983) );
  XNOR2_X1 U5504 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_f82), .ZN(n4982) );
  NAND4_X1 U5505 ( .A1(n4985), .A2(n4984), .A3(n4983), .A4(n4982), .ZN(n4989)
         );
  XNOR2_X1 U5506 ( .A(keyinput_f55), .B(n4986), .ZN(n4988) );
  XNOR2_X1 U5507 ( .A(keyinput_f54), .B(n2638), .ZN(n4987) );
  NOR4_X1 U5508 ( .A1(n4990), .A2(n4989), .A3(n4988), .A4(n4987), .ZN(n5022)
         );
  AOI22_X1 U5509 ( .A1(n4992), .A2(keyinput_f122), .B1(n2579), .B2(
        keyinput_f62), .ZN(n4991) );
  OAI221_X1 U5510 ( .B1(n4992), .B2(keyinput_f122), .C1(n2579), .C2(
        keyinput_f62), .A(n4991), .ZN(n5003) );
  AOI22_X1 U5511 ( .A1(n2648), .A2(keyinput_f18), .B1(n4994), .B2(keyinput_f33), .ZN(n4993) );
  OAI221_X1 U5512 ( .B1(n2648), .B2(keyinput_f18), .C1(n4994), .C2(
        keyinput_f33), .A(n4993), .ZN(n5002) );
  XOR2_X1 U5513 ( .A(n4995), .B(keyinput_f47), .Z(n5000) );
  XOR2_X1 U5514 ( .A(n4996), .B(keyinput_f123), .Z(n4999) );
  XNOR2_X1 U5515 ( .A(DATAI_4_), .B(keyinput_f27), .ZN(n4998) );
  XNOR2_X1 U5516 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_f58), .ZN(n4997) );
  NAND4_X1 U5517 ( .A1(n5000), .A2(n4999), .A3(n4998), .A4(n4997), .ZN(n5001)
         );
  NOR3_X1 U5518 ( .A1(n5003), .A2(n5002), .A3(n5001), .ZN(n5021) );
  AOI22_X1 U5519 ( .A1(n5005), .A2(keyinput_f22), .B1(n2584), .B2(keyinput_f51), .ZN(n5004) );
  OAI221_X1 U5520 ( .B1(n5005), .B2(keyinput_f22), .C1(n2584), .C2(
        keyinput_f51), .A(n5004), .ZN(n5010) );
  XNOR2_X1 U5521 ( .A(n5006), .B(keyinput_f73), .ZN(n5009) );
  XNOR2_X1 U5522 ( .A(n5007), .B(keyinput_f93), .ZN(n5008) );
  OR3_X1 U5523 ( .A1(n5010), .A2(n5009), .A3(n5008), .ZN(n5019) );
  AOI22_X1 U5524 ( .A1(n5013), .A2(keyinput_f109), .B1(keyinput_f98), .B2(
        n5012), .ZN(n5011) );
  OAI221_X1 U5525 ( .B1(n5013), .B2(keyinput_f109), .C1(n5012), .C2(
        keyinput_f98), .A(n5011), .ZN(n5018) );
  AOI22_X1 U5526 ( .A1(n5016), .A2(keyinput_f92), .B1(keyinput_f95), .B2(n5015), .ZN(n5014) );
  OAI221_X1 U5527 ( .B1(n5016), .B2(keyinput_f92), .C1(n5015), .C2(
        keyinput_f95), .A(n5014), .ZN(n5017) );
  NOR3_X1 U5528 ( .A1(n5019), .A2(n5018), .A3(n5017), .ZN(n5020) );
  NAND4_X1 U5529 ( .A1(n5023), .A2(n5022), .A3(n5021), .A4(n5020), .ZN(n5080)
         );
  AOI22_X1 U5530 ( .A1(n5026), .A2(keyinput_f106), .B1(keyinput_f105), .B2(
        n5025), .ZN(n5024) );
  OAI221_X1 U5531 ( .B1(n5026), .B2(keyinput_f106), .C1(n5025), .C2(
        keyinput_f105), .A(n5024), .ZN(n5039) );
  AOI22_X1 U5532 ( .A1(n5029), .A2(keyinput_f96), .B1(keyinput_f99), .B2(n5028), .ZN(n5027) );
  OAI221_X1 U5533 ( .B1(n5029), .B2(keyinput_f96), .C1(n5028), .C2(
        keyinput_f99), .A(n5027), .ZN(n5038) );
  AOI22_X1 U5534 ( .A1(n5032), .A2(keyinput_f101), .B1(keyinput_f104), .B2(
        n5031), .ZN(n5030) );
  OAI221_X1 U5535 ( .B1(n5032), .B2(keyinput_f101), .C1(n5031), .C2(
        keyinput_f104), .A(n5030), .ZN(n5037) );
  AOI22_X1 U5536 ( .A1(n5035), .A2(keyinput_f97), .B1(keyinput_f111), .B2(
        n5034), .ZN(n5033) );
  OAI221_X1 U5537 ( .B1(n5035), .B2(keyinput_f97), .C1(n5034), .C2(
        keyinput_f111), .A(n5033), .ZN(n5036) );
  NOR4_X1 U5538 ( .A1(n5039), .A2(n5038), .A3(n5037), .A4(n5036), .ZN(n5078)
         );
  INV_X1 U5539 ( .A(DATAI_7_), .ZN(n5041) );
  AOI22_X1 U5540 ( .A1(n5041), .A2(keyinput_f24), .B1(keyinput_f26), .B2(n2552), .ZN(n5040) );
  OAI221_X1 U5541 ( .B1(n5041), .B2(keyinput_f24), .C1(n2552), .C2(
        keyinput_f26), .A(n5040), .ZN(n5051) );
  AOI22_X1 U5542 ( .A1(n5043), .A2(keyinput_f39), .B1(n3703), .B2(keyinput_f45), .ZN(n5042) );
  OAI221_X1 U5543 ( .B1(n5043), .B2(keyinput_f39), .C1(n3703), .C2(
        keyinput_f45), .A(n5042), .ZN(n5050) );
  XOR2_X1 U5544 ( .A(n5044), .B(keyinput_f20), .Z(n5048) );
  XNOR2_X1 U5545 ( .A(DATAI_14_), .B(keyinput_f17), .ZN(n5047) );
  XNOR2_X1 U5546 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_f79), .ZN(n5046) );
  XNOR2_X1 U5547 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_f59), .ZN(n5045) );
  NAND4_X1 U5548 ( .A1(n5048), .A2(n5047), .A3(n5046), .A4(n5045), .ZN(n5049)
         );
  NOR3_X1 U5549 ( .A1(n5051), .A2(n5050), .A3(n5049), .ZN(n5077) );
  AOI22_X1 U5550 ( .A1(n2779), .A2(keyinput_f74), .B1(keyinput_f30), .B2(n2346), .ZN(n5052) );
  OAI221_X1 U5551 ( .B1(n2779), .B2(keyinput_f74), .C1(n2346), .C2(
        keyinput_f30), .A(n5052), .ZN(n5064) );
  AOI22_X1 U5552 ( .A1(n5055), .A2(keyinput_f23), .B1(keyinput_f121), .B2(
        n5054), .ZN(n5053) );
  OAI221_X1 U5553 ( .B1(n5055), .B2(keyinput_f23), .C1(n5054), .C2(
        keyinput_f121), .A(n5053), .ZN(n5063) );
  AOI22_X1 U5554 ( .A1(n5058), .A2(keyinput_f13), .B1(n5057), .B2(keyinput_f12), .ZN(n5056) );
  OAI221_X1 U5555 ( .B1(n5058), .B2(keyinput_f13), .C1(n5057), .C2(
        keyinput_f12), .A(n5056), .ZN(n5062) );
  XNOR2_X1 U5556 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_f68), .ZN(n5060) );
  XNOR2_X1 U5557 ( .A(DATAI_24_), .B(keyinput_f7), .ZN(n5059) );
  NAND2_X1 U5558 ( .A1(n5060), .A2(n5059), .ZN(n5061) );
  NOR4_X1 U5559 ( .A1(n5064), .A2(n5063), .A3(n5062), .A4(n5061), .ZN(n5076)
         );
  AOI22_X1 U5560 ( .A1(n5066), .A2(keyinput_f16), .B1(n2760), .B2(keyinput_f4), 
        .ZN(n5065) );
  OAI221_X1 U5561 ( .B1(n5066), .B2(keyinput_f16), .C1(n2760), .C2(keyinput_f4), .A(n5065), .ZN(n5074) );
  AOI22_X1 U5562 ( .A1(n2809), .A2(keyinput_f87), .B1(n2782), .B2(keyinput_f75), .ZN(n5067) );
  OAI221_X1 U5563 ( .B1(n2809), .B2(keyinput_f87), .C1(n2782), .C2(
        keyinput_f75), .A(n5067), .ZN(n5073) );
  XNOR2_X1 U5564 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_f76), .ZN(n5071) );
  XNOR2_X1 U5565 ( .A(IR_REG_23__SCAN_IN), .B(keyinput_f78), .ZN(n5070) );
  XNOR2_X1 U5566 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_f64), .ZN(n5069) );
  XNOR2_X1 U5567 ( .A(DATAI_2_), .B(keyinput_f29), .ZN(n5068) );
  NAND4_X1 U5568 ( .A1(n5071), .A2(n5070), .A3(n5069), .A4(n5068), .ZN(n5072)
         );
  NOR3_X1 U5569 ( .A1(n5074), .A2(n5073), .A3(n5072), .ZN(n5075) );
  NAND4_X1 U5570 ( .A1(n5078), .A2(n5077), .A3(n5076), .A4(n5075), .ZN(n5079)
         );
  OR4_X1 U5571 ( .A1(n5082), .A2(n5081), .A3(n5080), .A4(n5079), .ZN(n5084) );
  AOI21_X1 U5572 ( .B1(keyinput_f81), .B2(n5084), .A(keyinput_g81), .ZN(n5086)
         );
  INV_X1 U5573 ( .A(keyinput_f81), .ZN(n5083) );
  AOI21_X1 U5574 ( .B1(n5084), .B2(n5083), .A(IR_REG_26__SCAN_IN), .ZN(n5085)
         );
  AOI22_X1 U5575 ( .A1(IR_REG_26__SCAN_IN), .A2(n5086), .B1(keyinput_g81), 
        .B2(n5085), .ZN(n5087) );
  AOI21_X1 U5576 ( .B1(n5089), .B2(n5088), .A(n5087), .ZN(n5091) );
  AOI22_X1 U5577 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n5090) );
  XNOR2_X1 U5578 ( .A(n5091), .B(n5090), .ZN(U3352) );
  CLKBUF_X1 U3003 ( .A(n2482), .Z(n2489) );
  NAND2_X1 U3157 ( .A1(n2281), .A2(IR_REG_31__SCAN_IN), .ZN(n2856) );
endmodule

