

module b20_C_AntiSAT_k_256_4 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, ADD_1068_U4, ADD_1068_U55, 
        ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, 
        ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, 
        ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, 
        ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, 
        P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, 
        P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, 
        P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, 
        P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, 
        P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, 
        P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, 
        P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, 
        P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, 
        P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, 
        P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, 
        P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, 
        P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, 
        P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, 
        P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, 
        P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, 
        P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, 
        P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, 
        P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, 
        P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, 
        P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, 
        P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, 
        P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559;

  INV_X1 U5011 ( .A(n8415), .ZN(n8395) );
  CLKBUF_X2 U5012 ( .A(n5634), .Z(n4507) );
  BUF_X1 U5013 ( .A(n6319), .Z(n4505) );
  AOI21_X1 U5014 ( .B1(n4806), .B2(n4805), .A(n4802), .ZN(n8382) );
  NOR2_X1 U5016 ( .A1(n7825), .A2(n7948), .ZN(n7982) );
  AND2_X1 U5017 ( .A1(n6612), .A2(n4610), .ZN(n5220) );
  BUF_X1 U5018 ( .A(n6298), .Z(n6482) );
  OR2_X1 U5019 ( .A1(n9415), .A2(n9414), .ZN(n9416) );
  INV_X1 U5020 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5905) );
  AND2_X1 U5021 ( .A1(n7587), .A2(n7591), .ZN(n7657) );
  NAND2_X1 U5022 ( .A1(n5145), .A2(n5144), .ZN(n7722) );
  XNOR2_X1 U5023 ( .A(n5304), .B(n5303), .ZN(n6640) );
  INV_X2 U5024 ( .A(n4610), .ZN(n6584) );
  AOI21_X1 U5025 ( .B1(n7051), .B2(n8366), .A(n8367), .ZN(n6250) );
  INV_X1 U5026 ( .A(n6804), .ZN(n4768) );
  INV_X1 U5027 ( .A(n9409), .ZN(n9721) );
  BUF_X1 U5028 ( .A(n6294), .Z(n6319) );
  NAND2_X2 U5029 ( .A1(n5751), .A2(n4608), .ZN(n5748) );
  OAI21_X1 U5030 ( .B1(n7627), .B2(n7898), .A(n7900), .ZN(n8530) );
  AOI21_X2 U5031 ( .B1(n8398), .B2(n7809), .A(n7812), .ZN(n8384) );
  NAND2_X2 U5032 ( .A1(n5768), .A2(n5767), .ZN(n6854) );
  NOR2_X2 U5033 ( .A1(n9269), .A2(n6500), .ZN(n8984) );
  OAI22_X2 U5034 ( .A1(n7552), .A2(n6152), .B1(n8232), .B2(n8086), .ZN(n7625)
         );
  OAI21_X2 U5035 ( .B1(n9596), .B2(n7887), .A(n7885), .ZN(n7552) );
  NOR2_X4 U5036 ( .A1(n5788), .A2(n5787), .ZN(n7008) );
  AOI21_X2 U5037 ( .B1(n9388), .B2(n5660), .A(n5659), .ZN(n9376) );
  NAND2_X2 U5038 ( .A1(n8665), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5737) );
  NAND2_X2 U5039 ( .A1(n5308), .A2(n5307), .ZN(n7524) );
  AOI21_X1 U5040 ( .B1(n8530), .B2(n7815), .A(n5973), .ZN(n8522) );
  INV_X2 U5041 ( .A(n9074), .ZN(n6500) );
  NAND2_X1 U5042 ( .A1(n6885), .A2(n10022), .ZN(n8192) );
  INV_X2 U5043 ( .A(n6895), .ZN(n8056) );
  NAND2_X1 U5044 ( .A1(n7070), .A2(n7982), .ZN(n6893) );
  NAND4_X2 U5045 ( .A1(n5785), .A2(n5784), .A3(n5783), .A4(n5782), .ZN(n8244)
         );
  INV_X1 U5046 ( .A(n8243), .ZN(n4735) );
  INV_X2 U5047 ( .A(n7220), .ZN(n5794) );
  NAND2_X2 U5048 ( .A1(n7989), .A2(n8291), .ZN(n5780) );
  XNOR2_X1 U5049 ( .A(n5740), .B(n5739), .ZN(n8670) );
  NAND2_X2 U5050 ( .A1(n6584), .A2(P1_U3086), .ZN(n9572) );
  NAND2_X1 U5051 ( .A1(n4926), .A2(n4925), .ZN(n4927) );
  NAND2_X1 U5052 ( .A1(n4598), .A2(n4595), .ZN(n8547) );
  AND2_X1 U5053 ( .A1(n4917), .A2(n4916), .ZN(n8748) );
  OAI21_X1 U5054 ( .B1(n8004), .B2(n10041), .A(n8003), .ZN(n8375) );
  XNOR2_X1 U5055 ( .A(n6549), .B(n8957), .ZN(n7760) );
  NOR2_X1 U5056 ( .A1(n9241), .A2(n9422), .ZN(n9431) );
  OAI21_X1 U5057 ( .B1(n4870), .B2(n8957), .A(n4869), .ZN(n4868) );
  AND2_X1 U5058 ( .A1(n6550), .A2(n5637), .ZN(n9263) );
  OAI21_X1 U5059 ( .B1(n5011), .B2(n5010), .A(n4580), .ZN(n5009) );
  NOR2_X1 U5060 ( .A1(n8095), .A2(n4556), .ZN(n5007) );
  AND2_X1 U5061 ( .A1(n9267), .A2(n4880), .ZN(n4879) );
  NAND3_X1 U5062 ( .A1(n6409), .A2(n6411), .A3(n7669), .ZN(n7697) );
  NAND2_X1 U5063 ( .A1(n9416), .A2(n8867), .ZN(n4866) );
  INV_X1 U5064 ( .A(n7512), .ZN(n7513) );
  NAND2_X1 U5065 ( .A1(n7599), .A2(n7598), .ZN(n7638) );
  OR2_X1 U5066 ( .A1(n9963), .A2(n9962), .ZN(n4935) );
  OR2_X1 U5067 ( .A1(n7568), .A2(n7569), .ZN(n7597) );
  NOR2_X1 U5068 ( .A1(n7346), .A2(n5302), .ZN(n7418) );
  NAND2_X1 U5069 ( .A1(n5377), .A2(n5376), .ZN(n8860) );
  NAND2_X1 U5070 ( .A1(n5152), .A2(n5151), .ZN(n7620) );
  NAND2_X1 U5071 ( .A1(n5342), .A2(n5341), .ZN(n8845) );
  NAND2_X1 U5072 ( .A1(n5360), .A2(n5359), .ZN(n8824) );
  NAND2_X1 U5073 ( .A1(n7298), .A2(n7961), .ZN(n7297) );
  AND2_X1 U5074 ( .A1(n6134), .A2(n6133), .ZN(n7298) );
  NOR2_X1 U5075 ( .A1(n6977), .A2(n6978), .ZN(n7086) );
  NAND2_X1 U5076 ( .A1(n5882), .A2(n5881), .ZN(n7608) );
  NAND2_X1 U5077 ( .A1(n5279), .A2(n5278), .ZN(n7199) );
  AND2_X1 U5078 ( .A1(n5857), .A2(n5856), .ZN(n10066) );
  NAND2_X1 U5079 ( .A1(n4641), .A2(n5096), .ZN(n5276) );
  INV_X1 U5080 ( .A(n6925), .ZN(n7264) );
  OR2_X1 U5081 ( .A1(n6269), .A2(n6274), .ZN(n6270) );
  AOI21_X1 U5082 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n8277), .A(n8247), .ZN(
        n8248) );
  INV_X1 U5083 ( .A(n10055), .ZN(n7122) );
  INV_X2 U5084 ( .A(n6274), .ZN(n6509) );
  NAND2_X1 U5085 ( .A1(n4769), .A2(n4768), .ZN(n6942) );
  INV_X2 U5086 ( .A(n6621), .ZN(n6731) );
  AND2_X1 U5087 ( .A1(n5759), .A2(n4736), .ZN(n10055) );
  OR2_X1 U5088 ( .A1(n8246), .A2(n6888), .ZN(n7824) );
  NAND4_X2 U5089 ( .A1(n5801), .A2(n5800), .A3(n5799), .A4(n5798), .ZN(n8242)
         );
  AND3_X1 U5090 ( .A1(n5791), .A2(n5790), .A3(n5789), .ZN(n10050) );
  NOR2_X1 U5091 ( .A1(n6791), .A2(n6790), .ZN(n6853) );
  NAND4_X2 U5092 ( .A1(n5764), .A2(n5763), .A3(n5762), .A4(n5761), .ZN(n8245)
         );
  NAND4_X1 U5093 ( .A1(n5206), .A2(n5205), .A3(n5204), .A4(n5203), .ZN(n6285)
         );
  NAND4_X1 U5094 ( .A1(n5775), .A2(n5774), .A3(n5773), .A4(n5772), .ZN(n8246)
         );
  NAND2_X1 U5095 ( .A1(n4684), .A2(n5086), .ZN(n5241) );
  AND2_X4 U5096 ( .A1(n5164), .A2(n5161), .ZN(n5202) );
  NAND2_X2 U5097 ( .A1(n5743), .A2(n8670), .ZN(n7220) );
  NAND2_X2 U5098 ( .A1(n5743), .A2(n5742), .ZN(n5992) );
  INV_X2 U5099 ( .A(n5780), .ZN(n6002) );
  XNOR2_X1 U5100 ( .A(n5442), .B(n5624), .ZN(n5634) );
  NAND2_X1 U5101 ( .A1(n4606), .A2(n4605), .ZN(n5752) );
  NAND2_X1 U5102 ( .A1(n5441), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5442) );
  XNOR2_X1 U5103 ( .A(n5750), .B(n5749), .ZN(n7989) );
  OR2_X1 U5104 ( .A1(n5738), .A2(n5905), .ZN(n5740) );
  AOI21_X1 U5105 ( .B1(n6202), .B2(P2_IR_REG_31__SCAN_IN), .A(n4608), .ZN(
        n4607) );
  OAI21_X1 U5106 ( .B1(n5685), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U5107 ( .A1(n5630), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5632) );
  NAND2_X2 U5108 ( .A1(n4610), .A2(P2_U3151), .ZN(n6582) );
  INV_X1 U5109 ( .A(n5890), .ZN(n5056) );
  INV_X1 U5110 ( .A(n5060), .ZN(n4809) );
  NOR2_X1 U5111 ( .A1(n5623), .A2(n4533), .ZN(n5629) );
  NAND2_X1 U5112 ( .A1(n4645), .A2(n4644), .ZN(n7798) );
  AND2_X1 U5113 ( .A1(n5057), .A2(n5735), .ZN(n4516) );
  CLKBUF_X1 U5114 ( .A(n5755), .Z(n5815) );
  AND4_X1 U5115 ( .A1(n5127), .A2(n5126), .A3(n5125), .A4(n5124), .ZN(n5128)
         );
  NAND2_X1 U5116 ( .A1(n4608), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4605) );
  AND2_X1 U5117 ( .A1(n5906), .A2(n5058), .ZN(n5057) );
  INV_X2 U5118 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X4 U5119 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5120 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n10354) );
  INV_X1 U5121 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5947) );
  INV_X1 U5122 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5726) );
  INV_X1 U5123 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5935) );
  INV_X1 U5124 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5731) );
  OAI22_X2 U5125 ( .A1(n6171), .A2(n6170), .B1(n8395), .B2(n8624), .ZN(n8393)
         );
  NAND2_X4 U5126 ( .A1(n6893), .A2(n6892), .ZN(n6895) );
  NOR2_X2 U5127 ( .A1(n9423), .A2(n9494), .ZN(n9421) );
  XNOR2_X2 U5128 ( .A(n5737), .B(n5736), .ZN(n5741) );
  AOI21_X1 U5129 ( .B1(n8750), .B2(n8677), .A(n8676), .ZN(n8730) );
  NOR2_X2 U5130 ( .A1(n8748), .A2(n8745), .ZN(n8750) );
  NOR2_X2 U5131 ( .A1(n9399), .A2(n9481), .ZN(n4774) );
  INV_X2 U5132 ( .A(n6772), .ZN(n9766) );
  NAND2_X1 U5133 ( .A1(n6612), .A2(n6584), .ZN(n4508) );
  INV_X2 U5134 ( .A(n6545), .ZN(n8910) );
  AOI211_X2 U5135 ( .C1(n6551), .C2(n6550), .A(n9422), .B(n9247), .ZN(n7768)
         );
  NAND2_X1 U5136 ( .A1(n4879), .A2(n8993), .ZN(n4877) );
  INV_X1 U5137 ( .A(n4804), .ZN(n4803) );
  OAI22_X1 U5138 ( .A1(n8385), .A2(n6173), .B1(n8386), .B2(n8223), .ZN(n4804)
         );
  NAND2_X1 U5139 ( .A1(n4738), .A2(n4517), .ZN(n7293) );
  NOR2_X1 U5140 ( .A1(n5116), .A2(n4900), .ZN(n4899) );
  INV_X1 U5141 ( .A(n5111), .ZN(n4900) );
  INV_X1 U5142 ( .A(n5303), .ZN(n5116) );
  NOR2_X1 U5143 ( .A1(n5318), .A2(n4897), .ZN(n4896) );
  NAND2_X1 U5144 ( .A1(n5475), .A2(n4642), .ZN(n5492) );
  NAND2_X1 U5145 ( .A1(n4643), .A2(n5472), .ZN(n4642) );
  NAND2_X1 U5146 ( .A1(n4664), .A2(n4663), .ZN(n5456) );
  AOI21_X1 U5147 ( .B1(n4665), .B2(n4514), .A(n4584), .ZN(n4663) );
  NAND2_X1 U5148 ( .A1(n7174), .A2(n4621), .ZN(n4620) );
  NOR2_X1 U5149 ( .A1(n4622), .A2(n6353), .ZN(n4621) );
  INV_X1 U5150 ( .A(n7175), .ZN(n4622) );
  NOR2_X1 U5151 ( .A1(n7976), .A2(n4733), .ZN(n4732) );
  INV_X1 U5152 ( .A(n5383), .ZN(n5385) );
  NAND2_X1 U5153 ( .A1(n7597), .A2(n7596), .ZN(n7636) );
  INV_X1 U5154 ( .A(n8670), .ZN(n5742) );
  INV_X1 U5155 ( .A(n5741), .ZN(n5743) );
  OR2_X1 U5156 ( .A1(n8386), .A2(n8396), .ZN(n6174) );
  INV_X1 U5157 ( .A(n4798), .ZN(n4797) );
  OAI21_X1 U5158 ( .B1(n4515), .B2(n6169), .A(n4559), .ZN(n4798) );
  OR2_X1 U5159 ( .A1(n8464), .A2(n8478), .ZN(n7917) );
  OR2_X1 U5160 ( .A1(n8470), .A2(n8456), .ZN(n7916) );
  NAND2_X1 U5161 ( .A1(n6008), .A2(n6007), .ZN(n6016) );
  INV_X1 U5162 ( .A(n6009), .ZN(n6008) );
  AND2_X1 U5163 ( .A1(n7909), .A2(n7915), .ZN(n7953) );
  OR2_X1 U5164 ( .A1(n10089), .A2(n9599), .ZN(n7880) );
  AOI21_X1 U5165 ( .B1(n9060), .B2(n9059), .A(n9058), .ZN(n9061) );
  NOR2_X1 U5166 ( .A1(n9057), .A2(n9056), .ZN(n9059) );
  INV_X1 U5167 ( .A(n4879), .ZN(n4878) );
  OR2_X1 U5168 ( .A1(n9500), .A2(n7698), .ZN(n9018) );
  OR2_X1 U5169 ( .A1(n9723), .A2(n6368), .ZN(n8836) );
  NOR2_X1 U5170 ( .A1(n4959), .A2(n5563), .ZN(n4955) );
  NOR2_X1 U5171 ( .A1(n6483), .A2(n9076), .ZN(n5563) );
  INV_X1 U5172 ( .A(n4966), .ZN(n4963) );
  NAND2_X1 U5173 ( .A1(n6251), .A2(n9064), .ZN(n9008) );
  AND2_X1 U5174 ( .A1(n5691), .A2(n5712), .ZN(n6515) );
  AND2_X1 U5175 ( .A1(n5137), .A2(n5129), .ZN(n4990) );
  NAND2_X1 U5176 ( .A1(n5595), .A2(n5594), .ZN(n5606) );
  INV_X1 U5177 ( .A(n4839), .ZN(n4838) );
  OAI21_X1 U5178 ( .B1(n4842), .B2(n4530), .A(n5402), .ZN(n4839) );
  NAND3_X1 U5179 ( .A1(n4928), .A2(n4628), .A3(n5128), .ZN(n5623) );
  AND2_X1 U5180 ( .A1(n5392), .A2(n5129), .ZN(n4628) );
  INV_X1 U5181 ( .A(n4847), .ZN(n4846) );
  OAI21_X1 U5182 ( .B1(n4849), .B2(n5351), .A(n5355), .ZN(n4847) );
  NOR2_X1 U5183 ( .A1(n5337), .A2(n4852), .ZN(n4851) );
  INV_X1 U5184 ( .A(n5121), .ZN(n4852) );
  XNOR2_X1 U5185 ( .A(n5336), .B(n10325), .ZN(n5335) );
  AND2_X1 U5186 ( .A1(n4899), .A2(n5318), .ZN(n4892) );
  NAND2_X1 U5187 ( .A1(n8117), .A2(n5044), .ZN(n5043) );
  INV_X1 U5188 ( .A(n5992), .ZN(n6111) );
  XNOR2_X1 U5189 ( .A(n8066), .B(n8383), .ZN(n8060) );
  NOR2_X1 U5190 ( .A1(n8407), .A2(n8415), .ZN(n6170) );
  INV_X1 U5191 ( .A(n4761), .ZN(n4760) );
  OAI21_X1 U5192 ( .B1(n7928), .B2(n4762), .A(n7951), .ZN(n4761) );
  OR2_X1 U5193 ( .A1(n8489), .A2(n8497), .ZN(n7909) );
  OR2_X1 U5194 ( .A1(n5864), .A2(n4745), .ZN(n4743) );
  NAND2_X1 U5195 ( .A1(n7846), .A2(n7870), .ZN(n4745) );
  INV_X1 U5196 ( .A(n8235), .ZN(n8118) );
  OR2_X1 U5197 ( .A1(n7572), .A2(n7606), .ZN(n7846) );
  INV_X1 U5198 ( .A(n8513), .ZN(n10031) );
  NAND2_X1 U5199 ( .A1(n5780), .A2(n6584), .ZN(n7790) );
  AND2_X1 U5200 ( .A1(n8736), .A2(n6448), .ZN(n4616) );
  INV_X1 U5201 ( .A(n8746), .ZN(n4916) );
  NAND2_X1 U5202 ( .A1(n4618), .A2(n4546), .ZN(n7512) );
  INV_X1 U5203 ( .A(n7514), .ZN(n4617) );
  NOR2_X1 U5204 ( .A1(n4771), .A2(n9251), .ZN(n4770) );
  INV_X1 U5205 ( .A(n4772), .ZN(n4771) );
  NAND2_X1 U5206 ( .A1(n6612), .A2(n6584), .ZN(n6545) );
  AOI21_X1 U5207 ( .B1(n4512), .B2(n5382), .A(n4551), .ZN(n4970) );
  OR2_X1 U5208 ( .A1(n8860), .A2(n9086), .ZN(n4972) );
  AOI21_X1 U5209 ( .B1(n4894), .B2(n4896), .A(n4553), .ZN(n4893) );
  INV_X1 U5210 ( .A(n4899), .ZN(n4894) );
  INV_X1 U5211 ( .A(n4821), .ZN(n4820) );
  NAND2_X1 U5212 ( .A1(n5276), .A2(n4518), .ZN(n4817) );
  OAI21_X1 U5213 ( .B1(n4823), .B2(n4822), .A(n5065), .ZN(n4821) );
  INV_X1 U5214 ( .A(n9752), .ZN(n9710) );
  NAND2_X2 U5215 ( .A1(n5675), .A2(n7722), .ZN(n6612) );
  NAND2_X1 U5216 ( .A1(n4987), .A2(n4986), .ZN(n9341) );
  AOI21_X1 U5217 ( .B1(n4988), .B2(n5469), .A(n4579), .ZN(n4986) );
  XNOR2_X1 U5218 ( .A(n5154), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5164) );
  NAND2_X1 U5219 ( .A1(n5155), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5154) );
  NAND2_X1 U5220 ( .A1(n5606), .A2(n5596), .ZN(n7721) );
  OR2_X1 U5221 ( .A1(n5595), .A2(n5594), .ZN(n5596) );
  OAI21_X1 U5222 ( .B1(n5492), .B2(n5491), .A(n5490), .ZN(n5509) );
  NAND2_X1 U5223 ( .A1(n5004), .A2(n8152), .ZN(n5003) );
  OAI21_X1 U5224 ( .B1(n8805), .B2(n8919), .A(n8806), .ZN(n4785) );
  NOR2_X1 U5225 ( .A1(n8804), .A2(n4789), .ZN(n4784) );
  NAND2_X1 U5226 ( .A1(n7970), .A2(n7897), .ZN(n4700) );
  AND2_X1 U5227 ( .A1(n7893), .A2(n7894), .ZN(n4698) );
  NAND2_X1 U5228 ( .A1(n7912), .A2(n7946), .ZN(n4706) );
  AND2_X1 U5229 ( .A1(n4711), .A2(n4708), .ZN(n4707) );
  NAND2_X1 U5230 ( .A1(n7911), .A2(n4712), .ZN(n4709) );
  NAND2_X1 U5231 ( .A1(n4712), .A2(n7908), .ZN(n4708) );
  AOI21_X1 U5232 ( .B1(n4679), .B2(n4676), .A(n8919), .ZN(n4675) );
  INV_X1 U5233 ( .A(n4681), .ZN(n4676) );
  AOI21_X1 U5234 ( .B1(n4680), .B2(n4520), .A(n4789), .ZN(n4677) );
  INV_X1 U5235 ( .A(n4675), .ZN(n4674) );
  AOI21_X1 U5236 ( .B1(n4677), .B2(n4678), .A(n8984), .ZN(n4673) );
  INV_X1 U5237 ( .A(n4680), .ZN(n4678) );
  AOI21_X1 U5238 ( .B1(n7923), .B2(n8444), .A(n4720), .ZN(n4719) );
  INV_X1 U5239 ( .A(n7926), .ZN(n4720) );
  NOR2_X1 U5240 ( .A1(n7931), .A2(n4718), .ZN(n4717) );
  AND2_X1 U5241 ( .A1(n7928), .A2(n7946), .ZN(n4718) );
  OR2_X1 U5242 ( .A1(n6144), .A2(n6143), .ZN(n6146) );
  AND2_X1 U5243 ( .A1(n7948), .A2(n8353), .ZN(n6891) );
  NAND2_X1 U5244 ( .A1(n4561), .A2(n4781), .ZN(n8902) );
  NAND2_X1 U5245 ( .A1(n9055), .A2(n9054), .ZN(n9060) );
  AND2_X1 U5246 ( .A1(n7762), .A2(n9072), .ZN(n8990) );
  AND2_X1 U5247 ( .A1(n4530), .A2(n4837), .ZN(n4836) );
  NAND2_X1 U5248 ( .A1(n4732), .A2(n4509), .ZN(n4730) );
  OR2_X1 U5249 ( .A1(n8610), .A2(n7805), .ZN(n7978) );
  AOI211_X1 U5250 ( .C1(n7941), .C2(n7940), .A(n7939), .B(n7976), .ZN(n7945)
         );
  NAND2_X1 U5251 ( .A1(n4942), .A2(n7001), .ZN(n4943) );
  AND2_X1 U5252 ( .A1(n9818), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4942) );
  AOI22_X1 U5253 ( .A1(n9825), .A2(n9823), .B1(n6992), .B2(n9827), .ZN(n10141)
         );
  NAND2_X1 U5254 ( .A1(n9828), .A2(n7016), .ZN(n7018) );
  NAND2_X1 U5255 ( .A1(n9864), .A2(n8313), .ZN(n8315) );
  NAND2_X1 U5256 ( .A1(n9889), .A2(n8317), .ZN(n8319) );
  AND3_X1 U5257 ( .A1(n4937), .A2(n4587), .A3(n4936), .ZN(n8254) );
  NAND2_X1 U5258 ( .A1(n9920), .A2(n4639), .ZN(n8322) );
  OR2_X1 U5259 ( .A1(n9919), .A2(n5916), .ZN(n4639) );
  NAND2_X1 U5260 ( .A1(n4935), .A2(n8259), .ZN(n8260) );
  OR2_X1 U5261 ( .A1(n8406), .A2(n8203), .ZN(n7809) );
  AND2_X1 U5262 ( .A1(n8203), .A2(n8406), .ZN(n7812) );
  OR2_X1 U5263 ( .A1(n8421), .A2(n8436), .ZN(n7951) );
  OR2_X1 U5264 ( .A1(n5993), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6009) );
  OR2_X1 U5265 ( .A1(n8503), .A2(n8103), .ZN(n7910) );
  OR2_X1 U5266 ( .A1(n8531), .A2(n8211), .ZN(n7816) );
  NAND2_X1 U5267 ( .A1(n10055), .A2(n8243), .ZN(n7835) );
  AND2_X1 U5268 ( .A1(n6220), .A2(n6604), .ZN(n7070) );
  INV_X1 U5269 ( .A(n6591), .ZN(n4737) );
  INV_X1 U5270 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5058) );
  OR2_X1 U5271 ( .A1(n8701), .A2(n8729), .ZN(n4924) );
  XNOR2_X1 U5272 ( .A(n6305), .B(n6509), .ZN(n6309) );
  NAND2_X1 U5273 ( .A1(n6304), .A2(n6303), .ZN(n6305) );
  XNOR2_X1 U5274 ( .A(n6275), .B(n6509), .ZN(n6277) );
  NAND2_X1 U5275 ( .A1(n6261), .A2(n6262), .ZN(n6266) );
  OAI21_X1 U5276 ( .B1(n7530), .B2(n4908), .A(n4905), .ZN(n6400) );
  INV_X1 U5277 ( .A(n7576), .ZN(n4908) );
  AND2_X1 U5278 ( .A1(n4906), .A2(n6394), .ZN(n4905) );
  INV_X1 U5279 ( .A(n8957), .ZN(n4873) );
  NAND2_X1 U5280 ( .A1(n8957), .A2(n4874), .ZN(n4869) );
  AND2_X1 U5281 ( .A1(n4874), .A2(n4871), .ZN(n4870) );
  INV_X1 U5282 ( .A(n4876), .ZN(n4871) );
  NAND2_X1 U5283 ( .A1(n9284), .A2(n9274), .ZN(n4880) );
  AND2_X1 U5284 ( .A1(n6483), .A2(n5638), .ZN(n8980) );
  NAND2_X1 U5285 ( .A1(n9357), .A2(n8976), .ZN(n4886) );
  INV_X1 U5286 ( .A(n8976), .ZN(n4883) );
  INV_X1 U5287 ( .A(n8889), .ZN(n4882) );
  INV_X1 U5288 ( .A(n5417), .ZN(n4969) );
  OR2_X1 U5289 ( .A1(n7524), .A2(n5316), .ZN(n9033) );
  INV_X1 U5290 ( .A(n4996), .ZN(n4993) );
  NAND2_X1 U5291 ( .A1(n7372), .A2(n5288), .ZN(n4998) );
  OR2_X1 U5292 ( .A1(n6612), .A2(n5187), .ZN(n5188) );
  AND2_X1 U5293 ( .A1(n6251), .A2(n7416), .ZN(n6262) );
  NAND2_X1 U5294 ( .A1(n6551), .A2(n6548), .ZN(n8988) );
  INV_X1 U5295 ( .A(n8980), .ZN(n8893) );
  OR2_X1 U5296 ( .A1(n6483), .A2(n5638), .ZN(n8968) );
  OR2_X1 U5297 ( .A1(n9323), .A2(n5640), .ZN(n9300) );
  NAND2_X1 U5298 ( .A1(n7755), .A2(n8715), .ZN(n9423) );
  AND2_X1 U5299 ( .A1(n5334), .A2(n4978), .ZN(n4977) );
  NAND2_X1 U5300 ( .A1(n4979), .A2(n4981), .ZN(n4978) );
  INV_X1 U5301 ( .A(n4982), .ZN(n4979) );
  NAND2_X1 U5302 ( .A1(n6945), .A2(n9028), .ZN(n8793) );
  NAND2_X1 U5303 ( .A1(n7789), .A2(n7788), .ZN(n7797) );
  INV_X1 U5304 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5124) );
  NOR2_X1 U5305 ( .A1(n5169), .A2(n4824), .ZN(n4823) );
  INV_X1 U5306 ( .A(n5099), .ZN(n4824) );
  NAND2_X1 U5307 ( .A1(n5276), .A2(n5097), .ZN(n4818) );
  XNOR2_X1 U5308 ( .A(n5095), .B(SI_6_), .ZN(n5260) );
  XNOR2_X1 U5309 ( .A(n5088), .B(SI_4_), .ZN(n5240) );
  NAND2_X1 U5310 ( .A1(n5070), .A2(n5069), .ZN(n4645) );
  NAND2_X1 U5311 ( .A1(n5072), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4644) );
  NAND2_X1 U5312 ( .A1(n4813), .A2(n4812), .ZN(n5070) );
  NOR2_X1 U5313 ( .A1(n4577), .A2(n5059), .ZN(n5047) );
  XNOR2_X1 U5314 ( .A(n7636), .B(n7646), .ZN(n7599) );
  INV_X1 U5315 ( .A(n5024), .ZN(n5023) );
  OAI22_X1 U5316 ( .A1(n8071), .A2(n5025), .B1(n8059), .B2(n8396), .ZN(n5024)
         );
  NAND2_X1 U5317 ( .A1(n8196), .A2(n5026), .ZN(n5025) );
  INV_X1 U5318 ( .A(n8195), .ZN(n5026) );
  NAND2_X1 U5319 ( .A1(n5034), .A2(n7161), .ZN(n5033) );
  AOI21_X1 U5320 ( .B1(n7087), .B2(n8243), .A(n7086), .ZN(n7090) );
  AND2_X1 U5321 ( .A1(n4510), .A2(n4535), .ZN(n5013) );
  NAND2_X1 U5322 ( .A1(n5012), .A2(n4535), .ZN(n5011) );
  OR2_X1 U5323 ( .A1(n4513), .A2(n4571), .ZN(n5012) );
  INV_X1 U5324 ( .A(n8095), .ZN(n5014) );
  OR2_X1 U5325 ( .A1(n5883), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U5326 ( .A1(n5040), .A2(n5045), .ZN(n5035) );
  NOR2_X1 U5327 ( .A1(n5042), .A2(n8079), .ZN(n5040) );
  NOR2_X1 U5328 ( .A1(n8015), .A2(n8232), .ZN(n5038) );
  NAND2_X1 U5329 ( .A1(n5794), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U5330 ( .A1(n4638), .A2(n6780), .ZN(n6844) );
  NAND2_X1 U5331 ( .A1(n6854), .A2(n6845), .ZN(n4638) );
  AND2_X1 U5332 ( .A1(n4951), .A2(n5765), .ZN(n5028) );
  NAND2_X1 U5333 ( .A1(n5905), .A2(n4951), .ZN(n4950) );
  OR2_X1 U5334 ( .A1(n7000), .A2(n9798), .ZN(n7001) );
  XNOR2_X1 U5335 ( .A(n7018), .B(n7017), .ZN(n10145) );
  NAND2_X1 U5336 ( .A1(n10145), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10144) );
  OAI21_X1 U5337 ( .B1(n7004), .B2(n4931), .A(n4549), .ZN(n4929) );
  NOR2_X1 U5338 ( .A1(n7017), .A2(n6985), .ZN(n4931) );
  NAND2_X1 U5339 ( .A1(n8307), .A2(n4640), .ZN(n8311) );
  OR2_X1 U5340 ( .A1(n8309), .A2(n8308), .ZN(n4640) );
  XNOR2_X1 U5341 ( .A(n8315), .B(n9872), .ZN(n9874) );
  NAND2_X1 U5342 ( .A1(n9874), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n9873) );
  OR2_X1 U5343 ( .A1(n9882), .A2(n4938), .ZN(n4937) );
  NAND2_X1 U5344 ( .A1(n4939), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4938) );
  NAND2_X1 U5345 ( .A1(n8252), .A2(n4939), .ZN(n4936) );
  OR2_X1 U5346 ( .A1(n9882), .A2(n9881), .ZN(n4941) );
  XNOR2_X1 U5347 ( .A(n8319), .B(n9904), .ZN(n9906) );
  NAND2_X1 U5348 ( .A1(n9906), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9905) );
  XNOR2_X1 U5349 ( .A(n8254), .B(n9904), .ZN(n9913) );
  NOR2_X1 U5350 ( .A1(n5897), .A2(n9913), .ZN(n9912) );
  NAND2_X1 U5351 ( .A1(n5056), .A2(n5057), .ZN(n5922) );
  XNOR2_X1 U5352 ( .A(n8322), .B(n9936), .ZN(n9938) );
  NAND2_X1 U5353 ( .A1(n9938), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n9937) );
  NAND2_X1 U5354 ( .A1(n9990), .A2(n9991), .ZN(n9989) );
  NAND2_X1 U5355 ( .A1(n5974), .A2(n5731), .ZN(n5988) );
  OR2_X1 U5356 ( .A1(n10014), .A2(n10013), .ZN(n4949) );
  XNOR2_X1 U5357 ( .A(n8382), .B(n8385), .ZN(n4599) );
  INV_X1 U5358 ( .A(n6173), .ZN(n4802) );
  NOR2_X1 U5359 ( .A1(n8383), .A2(n10032), .ZN(n4597) );
  AND2_X1 U5360 ( .A1(n6174), .A2(n7936), .ZN(n8385) );
  OAI21_X1 U5361 ( .B1(n4760), .B2(n4758), .A(n7932), .ZN(n4757) );
  INV_X1 U5362 ( .A(n8410), .ZN(n4758) );
  AOI21_X1 U5363 ( .B1(n4797), .B2(n4515), .A(n4558), .ZN(n4795) );
  NOR2_X1 U5364 ( .A1(n8449), .A2(n7928), .ZN(n4759) );
  AND2_X1 U5365 ( .A1(n7932), .A2(n7933), .ZN(n8410) );
  NAND2_X1 U5366 ( .A1(n6065), .A2(n6064), .ZN(n6075) );
  INV_X1 U5367 ( .A(n6066), .ZN(n6065) );
  OR2_X1 U5368 ( .A1(n6043), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6054) );
  NOR2_X1 U5369 ( .A1(n6040), .A2(n4763), .ZN(n4762) );
  AND2_X1 U5370 ( .A1(n7951), .A2(n7950), .ZN(n8426) );
  NAND2_X1 U5371 ( .A1(n8450), .A2(n8444), .ZN(n4764) );
  OR2_X1 U5372 ( .A1(n6033), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6043) );
  AND2_X1 U5373 ( .A1(n7916), .A2(n7909), .ZN(n4748) );
  NAND2_X1 U5374 ( .A1(n8488), .A2(n7953), .ZN(n4749) );
  NOR2_X1 U5375 ( .A1(n6158), .A2(n4808), .ZN(n4807) );
  OR2_X1 U5376 ( .A1(n5967), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5982) );
  AOI21_X1 U5377 ( .B1(n4752), .B2(n7891), .A(n4751), .ZN(n4750) );
  INV_X1 U5378 ( .A(n7896), .ZN(n4751) );
  NAND2_X1 U5379 ( .A1(n5927), .A2(n5926), .ZN(n5940) );
  INV_X1 U5380 ( .A(n5928), .ZN(n5927) );
  NAND2_X1 U5381 ( .A1(n4800), .A2(n4799), .ZN(n9596) );
  OR2_X1 U5382 ( .A1(n10089), .A2(n8234), .ZN(n4799) );
  NAND2_X1 U5383 ( .A1(n4801), .A2(n4544), .ZN(n4800) );
  INV_X1 U5384 ( .A(n5863), .ZN(n4747) );
  OR2_X1 U5385 ( .A1(n5847), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5870) );
  NAND2_X1 U5386 ( .A1(n6138), .A2(n6137), .ZN(n7447) );
  AOI21_X1 U5387 ( .B1(n4528), .B2(n4742), .A(n4741), .ZN(n4740) );
  INV_X1 U5388 ( .A(n7836), .ZN(n4742) );
  INV_X1 U5389 ( .A(n7855), .ZN(n4741) );
  NAND2_X1 U5390 ( .A1(n4739), .A2(n4528), .ZN(n4738) );
  INV_X1 U5391 ( .A(n7053), .ZN(n7957) );
  NAND2_X1 U5392 ( .A1(n7122), .A2(n4735), .ZN(n7849) );
  AND2_X1 U5393 ( .A1(n7946), .A2(n6886), .ZN(n8513) );
  INV_X1 U5394 ( .A(n10032), .ZN(n8511) );
  NAND2_X1 U5395 ( .A1(n5952), .A2(n5951), .ZN(n8016) );
  OR2_X1 U5396 ( .A1(n7296), .A2(n7051), .ZN(n10082) );
  NAND2_X1 U5397 ( .A1(n5051), .A2(n5050), .ZN(n5722) );
  AOI21_X1 U5398 ( .B1(n5053), .B2(n5905), .A(n5905), .ZN(n5050) );
  INV_X1 U5399 ( .A(n5054), .ZN(n5053) );
  NAND2_X1 U5400 ( .A1(n5722), .A2(n10436), .ZN(n6117) );
  AND2_X1 U5401 ( .A1(n5029), .A2(n5765), .ZN(n6784) );
  AND2_X1 U5402 ( .A1(n6363), .A2(n6357), .ZN(n4915) );
  NOR2_X1 U5403 ( .A1(n4924), .A2(n4922), .ZN(n4921) );
  INV_X1 U5404 ( .A(n8677), .ZN(n4922) );
  OR2_X1 U5405 ( .A1(n4924), .A2(n8678), .ZN(n4920) );
  INV_X1 U5406 ( .A(n4626), .ZN(n4625) );
  NAND2_X1 U5407 ( .A1(n7697), .A2(n8717), .ZN(n4623) );
  OAI21_X1 U5408 ( .B1(n8708), .B2(n4627), .A(n8718), .ZN(n4626) );
  AND2_X1 U5409 ( .A1(n6469), .A2(n6468), .ZN(n8745) );
  NAND2_X1 U5410 ( .A1(n4619), .A2(n4620), .ZN(n4618) );
  AND2_X1 U5411 ( .A1(n4569), .A2(n6352), .ZN(n4619) );
  NAND2_X1 U5412 ( .A1(n5631), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U5413 ( .A1(n5201), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5181) );
  OR2_X1 U5414 ( .A1(n9575), .A2(n9574), .ZN(n9577) );
  XNOR2_X1 U5415 ( .A(n9446), .B(n9075), .ZN(n9286) );
  OR2_X1 U5416 ( .A1(n9358), .A2(n9357), .ZN(n9360) );
  AND2_X1 U5417 ( .A1(n8874), .A2(n8877), .ZN(n9400) );
  INV_X1 U5418 ( .A(n8947), .ZN(n4971) );
  OR2_X1 U5419 ( .A1(n7703), .A2(n5382), .ZN(n4973) );
  AOI21_X1 U5420 ( .B1(n4860), .B2(n5656), .A(n4862), .ZN(n4859) );
  AND2_X1 U5421 ( .A1(n9018), .A2(n9015), .ZN(n8947) );
  NOR2_X2 U5422 ( .A1(n7739), .A2(n8860), .ZN(n7755) );
  OR2_X1 U5423 ( .A1(n9723), .A2(n9090), .ZN(n4982) );
  NAND2_X1 U5424 ( .A1(n9723), .A2(n9090), .ZN(n4981) );
  NOR2_X1 U5425 ( .A1(n5652), .A2(n4864), .ZN(n5653) );
  INV_X1 U5426 ( .A(n4896), .ZN(n4895) );
  AND2_X1 U5427 ( .A1(n4890), .A2(n4893), .ZN(n4889) );
  INV_X1 U5428 ( .A(n4892), .ZN(n4890) );
  NOR2_X1 U5429 ( .A1(n7524), .A2(n9091), .ZN(n5317) );
  AND2_X1 U5430 ( .A1(n8811), .A2(n8812), .ZN(n7280) );
  NOR2_X1 U5431 ( .A1(n4997), .A2(n7280), .ZN(n4996) );
  NOR2_X1 U5432 ( .A1(n5287), .A2(n7182), .ZN(n4997) );
  NOR2_X1 U5433 ( .A1(n7199), .A2(n9094), .ZN(n5287) );
  AND2_X1 U5434 ( .A1(n7183), .A2(n7182), .ZN(n7185) );
  OR2_X1 U5435 ( .A1(n6524), .A2(n9064), .ZN(n9422) );
  XNOR2_X1 U5436 ( .A(n6276), .B(n7153), .ZN(n8928) );
  NAND2_X1 U5437 ( .A1(n6252), .A2(n6262), .ZN(n7194) );
  NAND2_X1 U5438 ( .A1(n8913), .A2(n8912), .ZN(n9240) );
  AND2_X1 U5439 ( .A1(n8904), .A2(n8988), .ZN(n8957) );
  NAND2_X1 U5440 ( .A1(n4954), .A2(n4953), .ZN(n9285) );
  AOI21_X1 U5441 ( .B1(n4955), .B2(n4962), .A(n4585), .ZN(n4953) );
  NAND2_X1 U5442 ( .A1(n8968), .A2(n8893), .ZN(n9301) );
  OR2_X1 U5443 ( .A1(n5545), .A2(n4963), .ZN(n4962) );
  OR2_X1 U5444 ( .A1(n5545), .A2(n4961), .ZN(n4960) );
  OR2_X1 U5445 ( .A1(n4964), .A2(n4963), .ZN(n4961) );
  INV_X1 U5446 ( .A(n9323), .ZN(n9454) );
  NAND2_X1 U5447 ( .A1(n9459), .A2(n9078), .ZN(n4966) );
  NOR2_X1 U5448 ( .A1(n4965), .A2(n5528), .ZN(n4964) );
  NOR2_X1 U5449 ( .A1(n9459), .A2(n9078), .ZN(n5528) );
  INV_X1 U5450 ( .A(n5506), .ZN(n4965) );
  AND2_X1 U5451 ( .A1(n9300), .A2(n8974), .ZN(n9311) );
  NAND2_X1 U5452 ( .A1(n5478), .A2(n5477), .ZN(n9367) );
  INV_X2 U5453 ( .A(n6612), .ZN(n5443) );
  AND2_X1 U5454 ( .A1(n5669), .A2(n9008), .ZN(n9752) );
  XNOR2_X1 U5455 ( .A(n7797), .B(n7796), .ZN(n8905) );
  NAND2_X1 U5456 ( .A1(n6107), .A2(SI_29_), .ZN(n7789) );
  INV_X1 U5457 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4765) );
  NAND2_X1 U5458 ( .A1(n5689), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5690) );
  XNOR2_X1 U5459 ( .A(n5586), .B(n5585), .ZN(n7677) );
  XNOR2_X1 U5460 ( .A(n5553), .B(n5567), .ZN(n7666) );
  AND2_X1 U5461 ( .A1(n5548), .A2(n5566), .ZN(n5553) );
  NAND2_X1 U5462 ( .A1(n5629), .A2(n5063), .ZN(n5685) );
  XNOR2_X1 U5463 ( .A(n5534), .B(n5533), .ZN(n7633) );
  NAND2_X1 U5464 ( .A1(n4666), .A2(n4667), .ZN(n5436) );
  OR2_X1 U5465 ( .A1(n5370), .A2(n4514), .ZN(n4666) );
  OAI21_X1 U5466 ( .B1(n5373), .B2(n4530), .A(n4838), .ZN(n5420) );
  NAND2_X1 U5467 ( .A1(n4841), .A2(n5386), .ZN(n5404) );
  NAND2_X1 U5468 ( .A1(n5373), .A2(n4842), .ZN(n4841) );
  NAND2_X1 U5469 ( .A1(n4850), .A2(n4849), .ZN(n5353) );
  NAND2_X1 U5470 ( .A1(n5319), .A2(n4851), .ZN(n4850) );
  NAND2_X1 U5471 ( .A1(n4848), .A2(n5121), .ZN(n5338) );
  OR2_X1 U5472 ( .A1(n5319), .A2(n5318), .ZN(n4848) );
  XNOR2_X1 U5473 ( .A(n4819), .B(n4702), .ZN(n6636) );
  INV_X1 U5474 ( .A(n5065), .ZN(n4702) );
  AOI21_X1 U5475 ( .B1(n4818), .B2(n4823), .A(n4822), .ZN(n4819) );
  NAND2_X1 U5476 ( .A1(n6042), .A2(n6041), .ZN(n8438) );
  AND4_X1 U5477 ( .A1(n5876), .A2(n5875), .A3(n5874), .A4(n5873), .ZN(n7606)
         );
  NAND2_X1 U5478 ( .A1(n6004), .A2(n6003), .ZN(n8489) );
  NAND2_X1 U5479 ( .A1(n8010), .A2(n8009), .ZN(n8117) );
  INV_X1 U5480 ( .A(n8224), .ZN(n8406) );
  AND3_X1 U5481 ( .A1(n6013), .A2(n6012), .A3(n6011), .ZN(n8497) );
  NAND2_X1 U5482 ( .A1(n7638), .A2(n5000), .ZN(n8010) );
  AND2_X1 U5483 ( .A1(n7637), .A2(n5001), .ZN(n5000) );
  INV_X1 U5484 ( .A(n7641), .ZN(n5001) );
  AND4_X1 U5485 ( .A1(n5987), .A2(n5986), .A3(n5985), .A4(n5984), .ZN(n8528)
         );
  NAND2_X1 U5486 ( .A1(n8055), .A2(n8054), .ZN(n8198) );
  NOR2_X1 U5487 ( .A1(n6853), .A2(n4548), .ZN(n6856) );
  NAND2_X1 U5488 ( .A1(n8263), .A2(n4946), .ZN(n4945) );
  INV_X1 U5489 ( .A(n8264), .ZN(n4946) );
  OR2_X1 U5490 ( .A1(n10014), .A2(n4947), .ZN(n4944) );
  OR2_X1 U5491 ( .A1(n8264), .A2(n10013), .ZN(n4947) );
  AND2_X1 U5492 ( .A1(n4593), .A2(n10010), .ZN(n8355) );
  INV_X1 U5493 ( .A(n8349), .ZN(n4594) );
  XNOR2_X1 U5494 ( .A(n7784), .B(n7976), .ZN(n8366) );
  NOR2_X1 U5495 ( .A1(n8002), .A2(n8001), .ZN(n8003) );
  NOR2_X1 U5496 ( .A1(n10031), .A2(n8396), .ZN(n8001) );
  XNOR2_X1 U5497 ( .A(n5725), .B(n5724), .ZN(n8353) );
  NAND2_X1 U5498 ( .A1(n5052), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U5499 ( .A1(n5974), .A2(n5055), .ZN(n5052) );
  NAND2_X1 U5500 ( .A1(n5598), .A2(n5597), .ZN(n9269) );
  NAND2_X1 U5501 ( .A1(n7721), .A2(n8910), .ZN(n5598) );
  INV_X1 U5502 ( .A(n8824), .ZN(n9506) );
  NOR2_X1 U5503 ( .A1(n7771), .A2(n6508), .ZN(n7774) );
  OR2_X1 U5504 ( .A1(n7775), .A2(n7772), .ZN(n6508) );
  NAND2_X1 U5505 ( .A1(n4614), .A2(n4613), .ZN(n8692) );
  AND2_X1 U5506 ( .A1(n4615), .A2(n8693), .ZN(n4613) );
  INV_X1 U5507 ( .A(n9500), .ZN(n8715) );
  NAND2_X1 U5508 ( .A1(n5498), .A2(n5497), .ZN(n9467) );
  XNOR2_X1 U5509 ( .A(n5708), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6254) );
  NAND2_X1 U5510 ( .A1(n4656), .A2(n4662), .ZN(n4655) );
  AND2_X1 U5511 ( .A1(n4661), .A2(n4659), .ZN(n4656) );
  NAND2_X1 U5512 ( .A1(n4660), .A2(n9011), .ZN(n4659) );
  OR2_X1 U5513 ( .A1(n5381), .A2(n5380), .ZN(n9086) );
  NAND2_X1 U5514 ( .A1(n4984), .A2(n4983), .ZN(n9257) );
  AND2_X1 U5515 ( .A1(n8955), .A2(n5604), .ZN(n4983) );
  INV_X1 U5516 ( .A(n9741), .ZN(n9430) );
  INV_X1 U5517 ( .A(n6251), .ZN(n9023) );
  OAI21_X1 U5518 ( .B1(n8793), .B2(n4789), .A(n4788), .ZN(n8801) );
  NAND2_X1 U5519 ( .A1(n8794), .A2(n4789), .ZN(n4788) );
  NAND2_X1 U5520 ( .A1(n4783), .A2(n8813), .ZN(n8834) );
  OAI21_X1 U5521 ( .B1(n4785), .B2(n4784), .A(n8810), .ZN(n4783) );
  NOR2_X1 U5522 ( .A1(n4698), .A2(n4696), .ZN(n4695) );
  NAND2_X1 U5523 ( .A1(n4697), .A2(n7888), .ZN(n4696) );
  INV_X1 U5524 ( .A(n4700), .ZN(n4697) );
  NAND2_X1 U5525 ( .A1(n4692), .A2(n4691), .ZN(n4690) );
  INV_X1 U5526 ( .A(n4698), .ZN(n4692) );
  NOR2_X1 U5527 ( .A1(n4699), .A2(n4700), .ZN(n4691) );
  AND2_X1 U5528 ( .A1(n9595), .A2(n7893), .ZN(n4699) );
  NAND2_X1 U5529 ( .A1(n4694), .A2(n4689), .ZN(n7902) );
  AND2_X1 U5530 ( .A1(n4693), .A2(n4690), .ZN(n4689) );
  NAND2_X1 U5531 ( .A1(n7889), .A2(n4695), .ZN(n4694) );
  AND2_X1 U5532 ( .A1(n7901), .A2(n8529), .ZN(n4693) );
  INV_X1 U5533 ( .A(n8888), .ZN(n4776) );
  NOR2_X1 U5534 ( .A1(n4714), .A2(n4713), .ZN(n4712) );
  INV_X1 U5535 ( .A(n7915), .ZN(n4713) );
  INV_X1 U5536 ( .A(n7907), .ZN(n4714) );
  AND2_X1 U5537 ( .A1(n7916), .A2(n7909), .ZN(n4711) );
  NAND2_X1 U5538 ( .A1(n8882), .A2(n4651), .ZN(n4650) );
  NOR2_X1 U5539 ( .A1(n4519), .A2(n8971), .ZN(n4651) );
  AOI21_X1 U5540 ( .B1(n4775), .B2(n4777), .A(n4778), .ZN(n4653) );
  INV_X1 U5541 ( .A(n9312), .ZN(n4778) );
  NOR2_X1 U5542 ( .A1(n4780), .A2(n4776), .ZN(n4775) );
  NOR2_X1 U5543 ( .A1(n4534), .A2(n9342), .ZN(n4780) );
  NAND2_X1 U5544 ( .A1(n4777), .A2(n8888), .ZN(n4779) );
  AND2_X1 U5545 ( .A1(n4669), .A2(n9274), .ZN(n4680) );
  NAND2_X1 U5546 ( .A1(n4560), .A2(n8896), .ZN(n4669) );
  NAND2_X1 U5547 ( .A1(n4647), .A2(n8919), .ZN(n4646) );
  NAND2_X1 U5548 ( .A1(n4704), .A2(n4706), .ZN(n7918) );
  OAI21_X1 U5549 ( .B1(n4705), .B2(n4703), .A(n4710), .ZN(n7920) );
  AND2_X1 U5550 ( .A1(n7917), .A2(n7916), .ZN(n4710) );
  NAND2_X1 U5551 ( .A1(n4672), .A2(n8898), .ZN(n4670) );
  OAI21_X1 U5552 ( .B1(n4674), .B2(n4679), .A(n4673), .ZN(n4672) );
  INV_X1 U5553 ( .A(n4782), .ZN(n4781) );
  OAI21_X1 U5554 ( .B1(n8898), .B2(n4789), .A(n8985), .ZN(n4782) );
  NAND2_X1 U5555 ( .A1(n4716), .A2(n4715), .ZN(n7935) );
  AND2_X1 U5556 ( .A1(n7930), .A2(n8410), .ZN(n4715) );
  OAI21_X1 U5557 ( .B1(n4719), .B2(n7928), .A(n4717), .ZN(n4716) );
  AND2_X1 U5558 ( .A1(n6166), .A2(n6165), .ZN(n6168) );
  NAND2_X1 U5559 ( .A1(n7576), .A2(n4907), .ZN(n4906) );
  INV_X1 U5560 ( .A(n6386), .ZN(n4907) );
  AND2_X1 U5561 ( .A1(n9514), .A2(n9243), .ZN(n9058) );
  INV_X1 U5562 ( .A(n5456), .ZN(n4811) );
  AND2_X1 U5563 ( .A1(n4667), .A2(n5433), .ZN(n4665) );
  INV_X1 U5564 ( .A(n5419), .ZN(n4837) );
  AND2_X1 U5565 ( .A1(n5352), .A2(n4851), .ZN(n4845) );
  NAND2_X1 U5566 ( .A1(n5114), .A2(SI_10_), .ZN(n5115) );
  INV_X1 U5567 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10271) );
  INV_X1 U5568 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4812) );
  INV_X1 U5569 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4813) );
  NAND2_X1 U5570 ( .A1(n5071), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5072) );
  INV_X1 U5571 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5071) );
  INV_X1 U5572 ( .A(n8177), .ZN(n5010) );
  NAND2_X1 U5573 ( .A1(n4733), .A2(n4727), .ZN(n4726) );
  NOR2_X1 U5574 ( .A1(n4509), .A2(n8383), .ZN(n4727) );
  AOI21_X1 U5575 ( .B1(n4732), .B2(n8383), .A(n4557), .ZN(n4725) );
  INV_X1 U5576 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4755) );
  OAI21_X1 U5577 ( .B1(P2_IR_REG_1__SCAN_IN), .B2(keyinput51), .A(n4636), .ZN(
        n4635) );
  NAND2_X1 U5578 ( .A1(keyinput51), .A2(P2_IR_REG_1__SCAN_IN), .ZN(n4636) );
  XNOR2_X1 U5579 ( .A(keyinput20), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n4637) );
  XNOR2_X1 U5580 ( .A(n4634), .B(P1_REG3_REG_20__SCAN_IN), .ZN(n4633) );
  INV_X1 U5581 ( .A(keyinput209), .ZN(n4634) );
  NAND2_X1 U5582 ( .A1(n5765), .A2(n4631), .ZN(n4630) );
  INV_X1 U5583 ( .A(keyinput179), .ZN(n4631) );
  NAND2_X1 U5584 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(keyinput179), .ZN(n4632) );
  NOR2_X1 U5585 ( .A1(n10156), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4930) );
  INV_X1 U5586 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4734) );
  NOR2_X1 U5587 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5717) );
  NOR2_X1 U5588 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5718) );
  OR2_X1 U5589 ( .A1(n9928), .A2(n4600), .ZN(n8258) );
  NOR2_X1 U5590 ( .A1(n9919), .A2(n8257), .ZN(n4600) );
  NAND2_X1 U5591 ( .A1(n9986), .A2(n4591), .ZN(n8327) );
  OR2_X1 U5592 ( .A1(n6232), .A2(n8062), .ZN(n7943) );
  INV_X1 U5593 ( .A(n6174), .ZN(n7937) );
  OR2_X1 U5594 ( .A1(n6075), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6088) );
  OR2_X1 U5595 ( .A1(n8438), .A2(n8447), .ZN(n7952) );
  INV_X1 U5596 ( .A(n6156), .ZN(n4808) );
  INV_X1 U5597 ( .A(n7892), .ZN(n4754) );
  OR2_X1 U5598 ( .A1(n6141), .A2(n6140), .ZN(n6147) );
  AND2_X1 U5599 ( .A1(n7960), .A2(n6146), .ZN(n6145) );
  OR2_X1 U5600 ( .A1(n5858), .A2(n7843), .ZN(n5860) );
  OAI21_X1 U5601 ( .B1(n5055), .B2(n5905), .A(n5724), .ZN(n5054) );
  OR2_X1 U5602 ( .A1(n5815), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U5603 ( .A1(n6294), .A2(n9755), .ZN(n4612) );
  INV_X1 U5604 ( .A(n6357), .ZN(n4913) );
  INV_X1 U5605 ( .A(n4629), .ZN(n6314) );
  AOI211_X1 U5606 ( .C1(n8994), .C2(n8993), .A(n8992), .B(n8991), .ZN(n9054)
         );
  AND2_X1 U5607 ( .A1(n8915), .A2(n8909), .ZN(n8922) );
  NOR2_X1 U5608 ( .A1(n6551), .A2(n6539), .ZN(n4772) );
  AND2_X1 U5609 ( .A1(n4863), .A2(n8817), .ZN(n4860) );
  INV_X1 U5610 ( .A(n8855), .ZN(n4862) );
  INV_X1 U5611 ( .A(n5115), .ZN(n4897) );
  NAND2_X1 U5612 ( .A1(n8835), .A2(n8836), .ZN(n4864) );
  NAND2_X1 U5613 ( .A1(n7349), .A2(n4766), .ZN(n7419) );
  NOR2_X1 U5614 ( .A1(n7359), .A2(n7524), .ZN(n4766) );
  OR2_X1 U5615 ( .A1(n7359), .A2(n6342), .ZN(n8831) );
  AND2_X1 U5616 ( .A1(n5487), .A2(n5470), .ZN(n4988) );
  NAND2_X1 U5617 ( .A1(n5244), .A2(n6943), .ZN(n8790) );
  INV_X1 U5618 ( .A(n6803), .ZN(n4769) );
  OAI21_X1 U5619 ( .B1(n5606), .B2(n4816), .A(n4814), .ZN(n7787) );
  INV_X1 U5620 ( .A(n4815), .ZN(n4814) );
  OAI21_X1 U5621 ( .B1(n4816), .B2(n5605), .A(n6106), .ZN(n4815) );
  INV_X1 U5622 ( .A(n4829), .ZN(n4828) );
  AOI21_X1 U5623 ( .B1(n4829), .B2(n4831), .A(n4827), .ZN(n4826) );
  INV_X1 U5624 ( .A(n5529), .ZN(n4827) );
  INV_X1 U5625 ( .A(n5490), .ZN(n4833) );
  AOI21_X1 U5626 ( .B1(n5491), .B2(n4832), .A(n4830), .ZN(n4829) );
  INV_X1 U5627 ( .A(n5510), .ZN(n4830) );
  NAND2_X1 U5628 ( .A1(n5422), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5423) );
  INV_X1 U5629 ( .A(n4668), .ZN(n4667) );
  OAI21_X1 U5630 ( .B1(n4514), .B2(n5369), .A(n4834), .ZN(n4668) );
  AOI21_X1 U5631 ( .B1(n4838), .B2(n4836), .A(n4835), .ZN(n4834) );
  INV_X1 U5632 ( .A(n5418), .ZN(n4835) );
  INV_X1 U5633 ( .A(n5386), .ZN(n4840) );
  NOR2_X1 U5634 ( .A1(n5387), .A2(n4843), .ZN(n4842) );
  INV_X1 U5635 ( .A(n5372), .ZN(n4843) );
  AOI21_X1 U5636 ( .B1(n4851), .B2(n5318), .A(n4552), .ZN(n4849) );
  NAND2_X1 U5637 ( .A1(n5118), .A2(n10451), .ZN(n5121) );
  XNOR2_X1 U5638 ( .A(n5113), .B(SI_10_), .ZN(n5303) );
  NAND2_X1 U5639 ( .A1(n5108), .A2(n5107), .ZN(n5111) );
  NAND2_X1 U5640 ( .A1(n5105), .A2(n5104), .ZN(n5169) );
  XNOR2_X1 U5641 ( .A(n5098), .B(SI_7_), .ZN(n5275) );
  INV_X1 U5642 ( .A(n5260), .ZN(n5094) );
  XNOR2_X1 U5643 ( .A(n5079), .B(SI_2_), .ZN(n5207) );
  OAI21_X1 U5644 ( .B1(n7798), .B2(n4686), .A(n4685), .ZN(n5075) );
  INV_X1 U5645 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4686) );
  INV_X1 U5646 ( .A(n8196), .ZN(n5027) );
  AND2_X1 U5647 ( .A1(n8152), .A2(n8447), .ZN(n5002) );
  INV_X1 U5648 ( .A(n8049), .ZN(n5004) );
  NAND2_X1 U5649 ( .A1(n5808), .A2(n5807), .ZN(n5819) );
  INV_X1 U5650 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5807) );
  INV_X1 U5651 ( .A(n5809), .ZN(n5808) );
  OR2_X1 U5652 ( .A1(n8095), .A2(n8134), .ZN(n8146) );
  NAND2_X1 U5653 ( .A1(n7090), .A2(n7089), .ZN(n7164) );
  AND2_X1 U5654 ( .A1(n5033), .A2(n4574), .ZN(n5031) );
  NAND2_X1 U5655 ( .A1(n4728), .A2(n4723), .ZN(n4722) );
  NOR2_X1 U5656 ( .A1(n7944), .A2(n4509), .ZN(n4723) );
  NAND2_X1 U5657 ( .A1(n7218), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5764) );
  NAND2_X1 U5658 ( .A1(n6839), .A2(n6838), .ZN(n6840) );
  NAND2_X1 U5659 ( .A1(n6844), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6846) );
  INV_X1 U5660 ( .A(n4943), .ZN(n9815) );
  NAND2_X1 U5661 ( .A1(n4934), .A2(n7005), .ZN(n10146) );
  NOR2_X1 U5662 ( .A1(n4637), .A2(n4635), .ZN(n10498) );
  NAND2_X1 U5663 ( .A1(n10144), .A2(n7019), .ZN(n7020) );
  NAND2_X1 U5664 ( .A1(n4932), .A2(n4934), .ZN(n10149) );
  NOR2_X1 U5665 ( .A1(n4933), .A2(n6985), .ZN(n4932) );
  INV_X1 U5666 ( .A(n7005), .ZN(n4933) );
  AOI21_X1 U5667 ( .B1(n6994), .B2(n10156), .A(n10139), .ZN(n6996) );
  AOI21_X1 U5668 ( .B1(n8249), .B2(n8310), .A(n9840), .ZN(n9862) );
  NAND2_X1 U5669 ( .A1(n9838), .A2(n8312), .ZN(n9866) );
  OR2_X1 U5670 ( .A1(n5853), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5865) );
  NAND2_X1 U5671 ( .A1(n9873), .A2(n8316), .ZN(n9890) );
  INV_X1 U5672 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U5673 ( .A1(n9905), .A2(n8320), .ZN(n9921) );
  NOR2_X1 U5674 ( .A1(n9912), .A2(n8255), .ZN(n9930) );
  NOR2_X1 U5675 ( .A1(n9930), .A2(n9929), .ZN(n9928) );
  NAND2_X1 U5676 ( .A1(n9937), .A2(n8323), .ZN(n9954) );
  NAND2_X1 U5677 ( .A1(n9987), .A2(n9988), .ZN(n9986) );
  AND2_X1 U5678 ( .A1(n9977), .A2(n8261), .ZN(n9996) );
  XNOR2_X1 U5679 ( .A(n8327), .B(n10003), .ZN(n10005) );
  NAND2_X1 U5680 ( .A1(n10005), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n10004) );
  NAND2_X1 U5681 ( .A1(n9989), .A2(n8288), .ZN(n10007) );
  OR2_X1 U5682 ( .A1(n6097), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8361) );
  INV_X1 U5683 ( .A(n7999), .ZN(n8000) );
  NOR2_X1 U5684 ( .A1(n8062), .A2(n10032), .ZN(n8002) );
  OR2_X1 U5685 ( .A1(n7813), .A2(n7812), .ZN(n8392) );
  NAND2_X1 U5686 ( .A1(n6053), .A2(n6052), .ZN(n6066) );
  INV_X1 U5687 ( .A(n6054), .ZN(n6053) );
  AND3_X1 U5688 ( .A1(n6029), .A2(n6028), .A3(n6027), .ZN(n8478) );
  NAND2_X1 U5689 ( .A1(n6024), .A2(n6023), .ZN(n6033) );
  INV_X1 U5690 ( .A(n6025), .ZN(n6024) );
  OR2_X1 U5691 ( .A1(n6016), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6025) );
  AND2_X1 U5692 ( .A1(n6039), .A2(n6038), .ZN(n8457) );
  INV_X1 U5693 ( .A(n7953), .ZN(n6159) );
  NAND2_X1 U5694 ( .A1(n5981), .A2(n5980), .ZN(n5993) );
  INV_X1 U5695 ( .A(n5982), .ZN(n5981) );
  NAND2_X1 U5696 ( .A1(n8522), .A2(n8521), .ZN(n8520) );
  INV_X1 U5697 ( .A(n6155), .ZN(n8521) );
  AND2_X1 U5698 ( .A1(n7816), .A2(n7815), .ZN(n8529) );
  NAND2_X1 U5699 ( .A1(n5954), .A2(n5953), .ZN(n5967) );
  INV_X1 U5700 ( .A(n5955), .ZN(n5954) );
  OR2_X1 U5701 ( .A1(n5940), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U5702 ( .A1(n5913), .A2(n5912), .ZN(n5928) );
  INV_X1 U5703 ( .A(n5914), .ZN(n5913) );
  OR2_X1 U5704 ( .A1(n5898), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5914) );
  AND4_X1 U5705 ( .A1(n5889), .A2(n5888), .A3(n5887), .A4(n5886), .ZN(n7646)
         );
  AND2_X1 U5706 ( .A1(n7879), .A2(n7877), .ZN(n7964) );
  NAND2_X1 U5707 ( .A1(n5869), .A2(n5868), .ZN(n5883) );
  INV_X1 U5708 ( .A(n5870), .ZN(n5869) );
  NAND2_X1 U5709 ( .A1(n7297), .A2(n6135), .ZN(n7335) );
  OR2_X1 U5710 ( .A1(n5819), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U5711 ( .A1(n5832), .A2(n5831), .ZN(n5847) );
  INV_X1 U5712 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5831) );
  INV_X1 U5713 ( .A(n5845), .ZN(n5832) );
  NAND2_X1 U5714 ( .A1(n5796), .A2(n7121), .ZN(n5809) );
  NAND2_X1 U5715 ( .A1(n10028), .A2(n6123), .ZN(n4790) );
  AND2_X1 U5716 ( .A1(n7135), .A2(n6120), .ZN(n7296) );
  NAND2_X1 U5717 ( .A1(n10020), .A2(n10025), .ZN(n10019) );
  AND2_X1 U5718 ( .A1(n6223), .A2(n6862), .ZN(n7071) );
  AND3_X1 U5719 ( .A1(n5830), .A2(n5829), .A3(n5828), .ZN(n10062) );
  AND2_X1 U5720 ( .A1(n5758), .A2(n5757), .ZN(n5759) );
  NAND2_X1 U5721 ( .A1(n5825), .A2(n4737), .ZN(n4736) );
  NAND2_X1 U5722 ( .A1(n5780), .A2(n4578), .ZN(n5758) );
  NAND2_X1 U5723 ( .A1(n7498), .A2(n7551), .ZN(n10077) );
  AND2_X1 U5724 ( .A1(n6872), .A2(n6883), .ZN(n6906) );
  INV_X1 U5725 ( .A(n10077), .ZN(n10090) );
  XNOR2_X1 U5726 ( .A(n6118), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7825) );
  NAND2_X1 U5727 ( .A1(n6117), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6118) );
  AND2_X1 U5728 ( .A1(n5731), .A2(n5727), .ZN(n5055) );
  NAND2_X1 U5729 ( .A1(n5056), .A2(n4545), .ZN(n5961) );
  NOR2_X2 U5730 ( .A1(n5961), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U5731 ( .A1(n4612), .A2(n6263), .ZN(n6269) );
  NAND2_X1 U5732 ( .A1(n4563), .A2(n8736), .ZN(n4615) );
  OR2_X1 U5733 ( .A1(n8687), .A2(n4904), .ZN(n4903) );
  NAND2_X1 U5734 ( .A1(n7693), .A2(n7697), .ZN(n8707) );
  NAND2_X1 U5735 ( .A1(n4629), .A2(n6318), .ZN(n7041) );
  NAND2_X1 U5736 ( .A1(n8707), .A2(n8708), .ZN(n8716) );
  INV_X1 U5737 ( .A(n8729), .ZN(n4925) );
  INV_X1 U5738 ( .A(n8730), .ZN(n4926) );
  OR2_X1 U5739 ( .A1(n5282), .A2(n5174), .ZN(n5296) );
  INV_X1 U5740 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6684) );
  OR2_X1 U5741 ( .A1(n5344), .A2(n5343), .ZN(n5361) );
  OR2_X1 U5742 ( .A1(n5329), .A2(n5162), .ZN(n5344) );
  NOR2_X1 U5743 ( .A1(n5499), .A2(n8752), .ZN(n5519) );
  INV_X1 U5744 ( .A(n4911), .ZN(n4910) );
  OAI21_X1 U5745 ( .B1(n4915), .B2(n4914), .A(n4912), .ZN(n4911) );
  INV_X1 U5746 ( .A(n7464), .ZN(n4914) );
  NAND2_X1 U5747 ( .A1(n6364), .A2(n4913), .ZN(n4912) );
  AND2_X1 U5748 ( .A1(n6516), .A2(n6633), .ZN(n7028) );
  NAND2_X1 U5749 ( .A1(n6314), .A2(n6317), .ZN(n7096) );
  NAND2_X1 U5750 ( .A1(n5252), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5267) );
  INV_X1 U5751 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5266) );
  NAND2_X1 U5752 ( .A1(n5556), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5578) );
  NOR2_X1 U5753 ( .A1(n10439), .A2(n5578), .ZN(n5614) );
  NAND2_X1 U5754 ( .A1(n6403), .A2(n6402), .ZN(n7669) );
  AND2_X1 U5755 ( .A1(n6254), .A2(n6251), .ZN(n9001) );
  NOR2_X1 U5756 ( .A1(n9063), .A2(n4537), .ZN(n4654) );
  INV_X1 U5757 ( .A(n9063), .ZN(n4660) );
  AND2_X1 U5758 ( .A1(n9577), .A2(n6711), .ZN(n9609) );
  AND2_X1 U5759 ( .A1(n9270), .A2(n4772), .ZN(n9247) );
  NAND2_X1 U5760 ( .A1(n4873), .A2(n4874), .ZN(n4872) );
  INV_X1 U5761 ( .A(n5558), .ZN(n5556) );
  INV_X1 U5762 ( .A(n4885), .ZN(n4884) );
  AOI21_X1 U5763 ( .B1(n4885), .B2(n4883), .A(n4882), .ZN(n4881) );
  AND2_X1 U5764 ( .A1(n5664), .A2(n4886), .ZN(n4885) );
  OAI21_X1 U5765 ( .B1(n4866), .B2(n4865), .A(n8877), .ZN(n9388) );
  INV_X1 U5766 ( .A(n9400), .ZN(n4865) );
  NOR2_X1 U5767 ( .A1(n5413), .A2(n5412), .ZN(n5427) );
  OAI21_X1 U5768 ( .B1(n4970), .B2(n4969), .A(n4581), .ZN(n4968) );
  NAND2_X1 U5769 ( .A1(n7747), .A2(n8947), .ZN(n5657) );
  OR2_X1 U5770 ( .A1(n5396), .A2(n5395), .ZN(n5413) );
  NOR2_X1 U5771 ( .A1(n5361), .A2(n7672), .ZN(n5378) );
  AND2_X1 U5772 ( .A1(n8817), .A2(n8843), .ZN(n8943) );
  AND2_X1 U5773 ( .A1(n5655), .A2(n8841), .ZN(n7734) );
  NOR2_X1 U5774 ( .A1(n5654), .A2(n4857), .ZN(n4856) );
  INV_X1 U5775 ( .A(n8837), .ZN(n4857) );
  NAND2_X1 U5776 ( .A1(n7734), .A2(n8943), .ZN(n7733) );
  NAND2_X1 U5777 ( .A1(n9035), .A2(n5651), .ZN(n9714) );
  INV_X1 U5778 ( .A(n4864), .ZN(n9712) );
  NOR2_X1 U5779 ( .A1(n5296), .A2(n6684), .ZN(n5309) );
  AND2_X1 U5780 ( .A1(n5309), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5327) );
  NOR2_X1 U5781 ( .A1(n9422), .A2(n4507), .ZN(n6525) );
  NOR2_X1 U5782 ( .A1(n7359), .A2(n9092), .ZN(n5302) );
  AND2_X1 U5783 ( .A1(n9033), .A2(n9713), .ZN(n8937) );
  OR2_X1 U5784 ( .A1(n5650), .A2(n8926), .ZN(n9032) );
  NAND2_X1 U5785 ( .A1(n4995), .A2(n4998), .ZN(n4994) );
  NAND2_X1 U5786 ( .A1(n4993), .A2(n4998), .ZN(n4992) );
  INV_X1 U5787 ( .A(n5287), .ZN(n4995) );
  AND2_X1 U5788 ( .A1(n8831), .A2(n8833), .ZN(n7347) );
  NAND2_X1 U5789 ( .A1(n7349), .A2(n7444), .ZN(n7420) );
  AND2_X1 U5790 ( .A1(n7286), .A2(n7372), .ZN(n7349) );
  NOR2_X1 U5791 ( .A1(n7195), .A2(n7199), .ZN(n7286) );
  NOR2_X1 U5792 ( .A1(n5267), .A2(n5266), .ZN(n5280) );
  OR2_X2 U5793 ( .A1(n6961), .A2(n6965), .ZN(n7195) );
  AND2_X1 U5794 ( .A1(n5648), .A2(n9026), .ZN(n6945) );
  NAND2_X1 U5795 ( .A1(n8790), .A2(n9028), .ZN(n6944) );
  NAND2_X1 U5796 ( .A1(n5220), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5189) );
  OAI21_X1 U5797 ( .B1(n4508), .B2(n6586), .A(n5188), .ZN(n4787) );
  NAND2_X1 U5798 ( .A1(n8928), .A2(n7148), .ZN(n7147) );
  INV_X1 U5799 ( .A(n8928), .ZN(n5642) );
  AOI21_X1 U5800 ( .B1(n9279), .B2(n9710), .A(n9278), .ZN(n9440) );
  AND2_X1 U5801 ( .A1(n8899), .A2(n6552), .ZN(n9267) );
  INV_X1 U5802 ( .A(n9286), .ZN(n9284) );
  NAND2_X1 U5803 ( .A1(n7666), .A2(n8910), .ZN(n5555) );
  INV_X1 U5804 ( .A(n4866), .ZN(n9401) );
  NAND2_X1 U5805 ( .A1(n5411), .A2(n5410), .ZN(n9494) );
  AOI21_X1 U5806 ( .B1(n4977), .B2(n4980), .A(n4550), .ZN(n4975) );
  INV_X1 U5807 ( .A(n4981), .ZN(n4980) );
  INV_X1 U5808 ( .A(n8931), .ZN(n6926) );
  AND2_X1 U5809 ( .A1(n6253), .A2(n9756), .ZN(n9499) );
  AND2_X1 U5810 ( .A1(n6255), .A2(n9023), .ZN(n9756) );
  XNOR2_X1 U5811 ( .A(n7802), .B(n7801), .ZN(n8911) );
  XNOR2_X1 U5812 ( .A(n7787), .B(n7785), .ZN(n6107) );
  XNOR2_X1 U5813 ( .A(n6105), .B(n6104), .ZN(n8671) );
  NAND2_X1 U5814 ( .A1(n5606), .A2(n5605), .ZN(n6105) );
  MUX2_X1 U5815 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5143), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5145) );
  XNOR2_X1 U5816 ( .A(n5530), .B(n5529), .ZN(n7611) );
  NAND2_X1 U5817 ( .A1(n4825), .A2(n4829), .ZN(n5530) );
  NAND2_X1 U5818 ( .A1(n5492), .A2(n4832), .ZN(n4825) );
  XNOR2_X1 U5819 ( .A(n5632), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6251) );
  NAND2_X1 U5820 ( .A1(n5373), .A2(n5372), .ZN(n5388) );
  OAI211_X1 U5821 ( .C1(n5112), .C2(n4895), .A(n4893), .B(n4888), .ZN(n6660)
         );
  INV_X1 U5822 ( .A(n5240), .ZN(n5087) );
  XNOR2_X1 U5823 ( .A(n5084), .B(SI_3_), .ZN(n5218) );
  XNOR2_X1 U5824 ( .A(n4687), .B(n4688), .ZN(n5185) );
  INV_X1 U5825 ( .A(n5075), .ZN(n4688) );
  NOR2_X1 U5826 ( .A1(n7313), .A2(n7312), .ZN(n7491) );
  NAND2_X1 U5827 ( .A1(n5022), .A2(n8196), .ZN(n8072) );
  NAND2_X1 U5828 ( .A1(n6085), .A2(n6084), .ZN(n8386) );
  NAND2_X1 U5829 ( .A1(n5939), .A2(n5938), .ZN(n8086) );
  INV_X1 U5830 ( .A(n8225), .ZN(n8436) );
  AND2_X1 U5831 ( .A1(n5017), .A2(n5023), .ZN(n5016) );
  INV_X1 U5832 ( .A(n8061), .ZN(n5017) );
  NAND2_X1 U5833 ( .A1(n5020), .A2(n5019), .ZN(n5018) );
  OR2_X1 U5834 ( .A1(n8061), .A2(n5023), .ZN(n5019) );
  OAI21_X1 U5835 ( .B1(n8061), .B2(n4531), .A(n5023), .ZN(n5020) );
  NAND2_X1 U5836 ( .A1(n8061), .A2(n4531), .ZN(n5021) );
  AOI21_X1 U5837 ( .B1(n5014), .B2(n4510), .A(n4513), .ZN(n8108) );
  NAND2_X1 U5838 ( .A1(n6022), .A2(n6021), .ZN(n8464) );
  NAND2_X1 U5839 ( .A1(n5966), .A2(n5965), .ZN(n8531) );
  NAND2_X1 U5840 ( .A1(n5032), .A2(n5033), .ZN(n7236) );
  NAND2_X1 U5841 ( .A1(n6015), .A2(n6014), .ZN(n8470) );
  INV_X1 U5842 ( .A(n5059), .ZN(n5046) );
  NAND2_X1 U5843 ( .A1(n8117), .A2(n8116), .ZN(n5048) );
  NAND2_X1 U5844 ( .A1(n5924), .A2(n5923), .ZN(n9591) );
  NAND2_X1 U5845 ( .A1(n5014), .A2(n5013), .ZN(n5008) );
  NAND2_X1 U5846 ( .A1(n7638), .A2(n7637), .ZN(n7640) );
  NAND2_X1 U5847 ( .A1(n5991), .A2(n5990), .ZN(n8503) );
  NAND2_X1 U5848 ( .A1(n5032), .A2(n5030), .ZN(n7309) );
  AND2_X1 U5849 ( .A1(n5031), .A2(n7239), .ZN(n5030) );
  NAND2_X1 U5850 ( .A1(n6083), .A2(n6082), .ZN(n8203) );
  AND4_X1 U5851 ( .A1(n5972), .A2(n5971), .A3(n5970), .A4(n5969), .ZN(n8211)
         );
  OAI21_X1 U5852 ( .B1(n8117), .B2(n5036), .A(n4521), .ZN(n8209) );
  INV_X1 U5853 ( .A(n5040), .ZN(n5036) );
  NAND2_X1 U5854 ( .A1(n5039), .A2(n5037), .ZN(n8208) );
  INV_X1 U5855 ( .A(n5038), .ZN(n5037) );
  NAND2_X1 U5856 ( .A1(n5043), .A2(n5040), .ZN(n5039) );
  OAI21_X1 U5857 ( .B1(n8291), .B2(n6783), .A(n4609), .ZN(n6760) );
  NAND2_X1 U5858 ( .A1(n8291), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4609) );
  OR2_X1 U5859 ( .A1(n6786), .A2(n5760), .ZN(n6839) );
  OAI21_X1 U5860 ( .B1(n6784), .B2(n4952), .A(n4950), .ZN(n5788) );
  NAND2_X1 U5861 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4952) );
  AOI21_X1 U5862 ( .B1(n6989), .B2(n6988), .A(n6987), .ZN(n9811) );
  NAND2_X1 U5863 ( .A1(n7001), .A2(n9818), .ZN(n9803) );
  XNOR2_X1 U5864 ( .A(n8311), .B(n9843), .ZN(n9839) );
  NAND2_X1 U5865 ( .A1(n9839), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9838) );
  NAND2_X1 U5866 ( .A1(n4936), .A2(n4937), .ZN(n9897) );
  OAI21_X1 U5867 ( .B1(n10012), .B2(n4601), .A(n9980), .ZN(n10015) );
  NAND2_X1 U5868 ( .A1(n4604), .A2(n4602), .ZN(n8300) );
  NAND2_X1 U5869 ( .A1(n4603), .A2(n8340), .ZN(n4602) );
  NAND2_X1 U5870 ( .A1(n8299), .A2(n8344), .ZN(n4604) );
  OAI21_X1 U5871 ( .B1(n8298), .B2(n8297), .A(n10157), .ZN(n4603) );
  INV_X1 U5872 ( .A(n9837), .ZN(n10159) );
  NAND2_X1 U5873 ( .A1(n4945), .A2(n4944), .ZN(n8336) );
  AOI22_X1 U5874 ( .A1(n8911), .A2(n7804), .B1(n7803), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n8363) );
  NOR2_X1 U5875 ( .A1(n4597), .A2(n4596), .ZN(n4595) );
  NAND2_X1 U5876 ( .A1(n4599), .A2(n8516), .ZN(n4598) );
  NOR2_X1 U5877 ( .A1(n8406), .A2(n10031), .ZN(n4596) );
  NAND2_X1 U5878 ( .A1(n6063), .A2(n6062), .ZN(n8407) );
  NAND2_X1 U5879 ( .A1(n4756), .A2(n4760), .ZN(n8409) );
  NAND2_X1 U5880 ( .A1(n8450), .A2(n4759), .ZN(n4756) );
  NAND2_X1 U5881 ( .A1(n6051), .A2(n6050), .ZN(n8421) );
  AND2_X1 U5882 ( .A1(n4764), .A2(n4762), .ZN(n8425) );
  NAND2_X1 U5883 ( .A1(n6032), .A2(n6031), .ZN(n8568) );
  NAND2_X1 U5884 ( .A1(n4749), .A2(n7909), .ZN(n8469) );
  NAND2_X1 U5885 ( .A1(n6157), .A2(n6156), .ZN(n8495) );
  NAND2_X1 U5886 ( .A1(n5979), .A2(n5978), .ZN(n8590) );
  INV_X1 U5887 ( .A(n4801), .ZN(n7541) );
  NAND2_X1 U5888 ( .A1(n5911), .A2(n5910), .ZN(n10089) );
  NAND2_X1 U5889 ( .A1(n4744), .A2(n7846), .ZN(n7453) );
  NAND2_X1 U5890 ( .A1(n5864), .A2(n5863), .ZN(n7379) );
  NAND2_X1 U5891 ( .A1(n4738), .A2(n4740), .ZN(n7270) );
  NAND2_X1 U5892 ( .A1(n7073), .A2(n4528), .ZN(n7075) );
  NAND2_X1 U5893 ( .A1(n7052), .A2(n7836), .ZN(n7073) );
  INV_X1 U5894 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7121) );
  OR2_X1 U5895 ( .A1(n10077), .A2(n7076), .ZN(n10023) );
  OR2_X1 U5896 ( .A1(n7077), .A2(n10023), .ZN(n8532) );
  INV_X1 U5897 ( .A(n8363), .ZN(n8605) );
  NAND2_X1 U5898 ( .A1(n7792), .A2(n7791), .ZN(n8610) );
  AND2_X1 U5899 ( .A1(n8379), .A2(n10082), .ZN(n4794) );
  INV_X1 U5900 ( .A(n8203), .ZN(n8621) );
  NAND2_X1 U5901 ( .A1(n4701), .A2(n5866), .ZN(n7572) );
  NAND2_X1 U5902 ( .A1(n6636), .A2(n7804), .ZN(n4701) );
  AND2_X1 U5903 ( .A1(n6864), .A2(n6606), .ZN(n6883) );
  AND2_X1 U5904 ( .A1(n6871), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6606) );
  INV_X1 U5905 ( .A(n6215), .ZN(n7692) );
  NAND2_X1 U5906 ( .A1(n5723), .A2(n6117), .ZN(n7948) );
  INV_X1 U5907 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6642) );
  INV_X1 U5908 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6639) );
  INV_X1 U5909 ( .A(n9855), .ZN(n8306) );
  INV_X1 U5910 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10288) );
  INV_X1 U5911 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6587) );
  INV_X1 U5912 ( .A(n7011), .ZN(n9798) );
  NOR2_X1 U5913 ( .A1(n5711), .A2(n7635), .ZN(n4901) );
  NAND2_X1 U5914 ( .A1(n4909), .A2(n6364), .ZN(n7462) );
  NAND2_X1 U5915 ( .A1(n7434), .A2(n6357), .ZN(n4909) );
  NAND2_X1 U5916 ( .A1(n5445), .A2(n5444), .ZN(n9481) );
  INV_X1 U5917 ( .A(n7153), .ZN(n5190) );
  AND2_X1 U5918 ( .A1(n4614), .A2(n4615), .ZN(n8694) );
  NAND2_X1 U5919 ( .A1(n4611), .A2(n4547), .ZN(n8773) );
  NAND2_X1 U5920 ( .A1(n8750), .A2(n4921), .ZN(n4611) );
  OR2_X1 U5921 ( .A1(n8701), .A2(n6481), .ZN(n4923) );
  INV_X1 U5922 ( .A(n4927), .ZN(n8728) );
  NAND2_X1 U5923 ( .A1(n5536), .A2(n5535), .ZN(n9323) );
  NAND2_X1 U5924 ( .A1(n4620), .A2(n6352), .ZN(n7434) );
  INV_X1 U5925 ( .A(n4902), .ZN(n8738) );
  AOI21_X1 U5926 ( .B1(n8686), .B2(n8687), .A(n4904), .ZN(n4902) );
  NAND2_X1 U5927 ( .A1(n7575), .A2(n7576), .ZN(n7574) );
  NAND2_X1 U5928 ( .A1(n7530), .A2(n6386), .ZN(n7575) );
  NOR2_X1 U5929 ( .A1(n6468), .A2(n4919), .ZN(n4918) );
  INV_X1 U5930 ( .A(n6464), .ZN(n4919) );
  NAND2_X1 U5931 ( .A1(n5426), .A2(n5425), .ZN(n9487) );
  INV_X1 U5932 ( .A(n8769), .ZN(n8775) );
  INV_X1 U5933 ( .A(n8765), .ZN(n8782) );
  NAND4_X1 U5934 ( .A1(n5257), .A2(n5256), .A3(n5255), .A4(n5254), .ZN(n9096)
         );
  NAND4_X1 U5935 ( .A1(n5232), .A2(n5231), .A3(n5230), .A4(n5229), .ZN(n9097)
         );
  NAND4_X1 U5936 ( .A1(n5217), .A2(n5216), .A3(n5215), .A4(n5214), .ZN(n9098)
         );
  NAND2_X1 U5937 ( .A1(n5201), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5205) );
  OR2_X1 U5938 ( .A1(n5180), .A2(n6663), .ZN(n5184) );
  NAND2_X1 U5939 ( .A1(n5200), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5183) );
  OR2_X1 U5940 ( .A1(n6679), .A2(n6680), .ZN(n6709) );
  XNOR2_X1 U5941 ( .A(n9248), .B(n9240), .ZN(n9241) );
  AND2_X1 U5942 ( .A1(n6547), .A2(n6546), .ZN(n7762) );
  AOI21_X1 U5943 ( .B1(n5676), .B2(n9710), .A(n6532), .ZN(n9266) );
  OR3_X1 U5944 ( .A1(n9271), .A2(n9270), .A3(n9422), .ZN(n9439) );
  NAND2_X1 U5945 ( .A1(n5577), .A2(n5576), .ZN(n9446) );
  NAND2_X1 U5946 ( .A1(n7677), .A2(n8910), .ZN(n5577) );
  NAND2_X1 U5947 ( .A1(n9360), .A2(n8976), .ZN(n9343) );
  NAND2_X1 U5948 ( .A1(n7703), .A2(n4512), .ZN(n4967) );
  NAND2_X1 U5949 ( .A1(n4973), .A2(n4512), .ZN(n9498) );
  NAND2_X1 U5950 ( .A1(n4973), .A2(n4972), .ZN(n7753) );
  NAND2_X1 U5951 ( .A1(n5394), .A2(n5393), .ZN(n9500) );
  INV_X1 U5952 ( .A(n7755), .ZN(n7708) );
  NAND2_X1 U5953 ( .A1(n7582), .A2(n8837), .ZN(n4858) );
  INV_X1 U5954 ( .A(n7620), .ZN(n7591) );
  NAND2_X1 U5955 ( .A1(n4976), .A2(n4981), .ZN(n7581) );
  NAND2_X1 U5956 ( .A1(n9709), .A2(n4982), .ZN(n4976) );
  NAND2_X1 U5957 ( .A1(n5326), .A2(n5325), .ZN(n9723) );
  NAND2_X1 U5958 ( .A1(n4893), .A2(n4895), .ZN(n4891) );
  NAND2_X1 U5959 ( .A1(n9749), .A2(n6525), .ZN(n9405) );
  NOR2_X1 U5960 ( .A1(n7185), .A2(n5287), .ZN(n7279) );
  OAI21_X1 U5961 ( .B1(n7183), .B2(n5287), .A(n4996), .ZN(n4999) );
  NOR2_X1 U5962 ( .A1(n9721), .A2(n7126), .ZN(n9741) );
  INV_X1 U5963 ( .A(n9737), .ZN(n9722) );
  AND2_X1 U5964 ( .A1(n9797), .A2(n9768), .ZN(n7727) );
  INV_X1 U5965 ( .A(n9240), .ZN(n9514) );
  INV_X1 U5966 ( .A(n7762), .ZN(n6551) );
  NAND2_X1 U5967 ( .A1(n9257), .A2(n6544), .ZN(n6549) );
  INV_X1 U5968 ( .A(n9269), .ZN(n9519) );
  XOR2_X1 U5969 ( .A(n9301), .B(n9296), .Z(n9528) );
  OR2_X1 U5970 ( .A1(n5507), .A2(n4962), .ZN(n4956) );
  NAND2_X1 U5971 ( .A1(n4957), .A2(n4966), .ZN(n9310) );
  NAND2_X1 U5972 ( .A1(n5507), .A2(n4964), .ZN(n4957) );
  NAND2_X1 U5973 ( .A1(n5507), .A2(n5506), .ZN(n9328) );
  INV_X1 U5974 ( .A(n9367), .ZN(n9544) );
  AND2_X1 U5975 ( .A1(n4989), .A2(n5470), .ZN(n9356) );
  OR2_X1 U5976 ( .A1(n9374), .A2(n5469), .ZN(n4989) );
  NOR2_X1 U5977 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n4985) );
  NAND2_X1 U5978 ( .A1(n7789), .A2(n6108), .ZN(n9568) );
  OR2_X1 U5979 ( .A1(n6107), .A2(SI_29_), .ZN(n6108) );
  INV_X1 U5980 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5069) );
  AND3_X1 U5981 ( .A1(n4944), .A2(n4592), .A3(n4945), .ZN(n8338) );
  NOR2_X1 U5982 ( .A1(n5062), .A2(n6248), .ZN(n6249) );
  NAND2_X1 U5983 ( .A1(n4793), .A2(n4791), .ZN(P2_U3455) );
  INV_X1 U5984 ( .A(n4792), .ZN(n4791) );
  OR2_X1 U5985 ( .A1(n8544), .A2(n10093), .ZN(n4793) );
  OAI22_X1 U5986 ( .A1(n4731), .A2(n8662), .B1(n10091), .B2(n8005), .ZN(n4792)
         );
  OR2_X1 U5987 ( .A1(n8960), .A2(n4658), .ZN(n4657) );
  INV_X1 U5988 ( .A(n5200), .ZN(n5253) );
  AND2_X4 U5989 ( .A1(n7996), .A2(n9567), .ZN(n5200) );
  AND2_X1 U5990 ( .A1(n4731), .A2(n7946), .ZN(n4509) );
  NOR2_X1 U5991 ( .A1(n8158), .A2(n8039), .ZN(n4510) );
  OR3_X1 U5992 ( .A1(n9007), .A2(n7416), .A3(n9070), .ZN(n4511) );
  INV_X2 U5993 ( .A(n5289), .ZN(n8906) );
  AND2_X4 U5994 ( .A1(n7996), .A2(n5161), .ZN(n5201) );
  AND2_X1 U5995 ( .A1(n4971), .A2(n4972), .ZN(n4512) );
  NOR2_X1 U5996 ( .A1(n8039), .A2(n8159), .ZN(n4513) );
  NAND2_X1 U5997 ( .A1(n4838), .A2(n4837), .ZN(n4514) );
  NOR2_X1 U5998 ( .A1(n6168), .A2(n6167), .ZN(n4515) );
  INV_X1 U5999 ( .A(n9898), .ZN(n4939) );
  NAND2_X1 U6000 ( .A1(n6103), .A2(n6102), .ZN(n8222) );
  INV_X1 U6001 ( .A(n7944), .ZN(n4733) );
  AND2_X1 U6002 ( .A1(n4740), .A2(n7854), .ZN(n4517) );
  INV_X1 U6003 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5129) );
  INV_X1 U6004 ( .A(n7359), .ZN(n7444) );
  NAND2_X1 U6005 ( .A1(n4991), .A2(n4990), .ZN(n5142) );
  AND2_X1 U6006 ( .A1(n5105), .A2(n5097), .ZN(n4518) );
  AND2_X1 U6007 ( .A1(n8881), .A2(n8880), .ZN(n4519) );
  NAND2_X1 U6008 ( .A1(n8896), .A2(n8968), .ZN(n4520) );
  AND2_X1 U6009 ( .A1(n4583), .A2(n5035), .ZN(n4521) );
  NOR2_X1 U6010 ( .A1(n9003), .A2(n4507), .ZN(n4522) );
  NAND2_X1 U6011 ( .A1(n5518), .A2(n5517), .ZN(n9459) );
  AND2_X1 U6012 ( .A1(n4764), .A2(n7925), .ZN(n4523) );
  AND2_X1 U6013 ( .A1(n7097), .A2(n6317), .ZN(n4524) );
  AND2_X1 U6014 ( .A1(n4522), .A2(n9064), .ZN(n4525) );
  AND2_X1 U6015 ( .A1(n4927), .A2(n6481), .ZN(n4526) );
  INV_X1 U6016 ( .A(n6232), .ZN(n8368) );
  OAI21_X1 U6017 ( .B1(n9568), .B2(n6110), .A(n6109), .ZN(n6232) );
  AND2_X1 U6018 ( .A1(n5459), .A2(SI_20_), .ZN(n4527) );
  NAND2_X1 U6019 ( .A1(n4589), .A2(n7096), .ZN(n7042) );
  INV_X1 U6020 ( .A(n9070), .ZN(n4662) );
  AND2_X1 U6021 ( .A1(n7855), .A2(n7851), .ZN(n4528) );
  INV_X1 U6022 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U6023 ( .A1(n5712), .A2(n4901), .ZN(n6261) );
  OR2_X1 U6024 ( .A1(n9297), .A2(n9446), .ZN(n4529) );
  INV_X1 U6025 ( .A(n5180), .ZN(n5213) );
  NAND2_X1 U6026 ( .A1(n4956), .A2(n4958), .ZN(n9296) );
  OR2_X1 U6027 ( .A1(n4840), .A2(n5403), .ZN(n4530) );
  INV_X1 U6028 ( .A(n4928), .ZN(n5146) );
  INV_X1 U6029 ( .A(n7961), .ZN(n7859) );
  NOR2_X1 U6030 ( .A1(n8071), .A2(n5027), .ZN(n4531) );
  AND2_X1 U6031 ( .A1(n7978), .A2(n7943), .ZN(n4532) );
  NAND4_X1 U6032 ( .A1(n5627), .A2(n5626), .A3(n5625), .A4(n5624), .ZN(n4533)
         );
  INV_X1 U6033 ( .A(n7017), .ZN(n10156) );
  NAND2_X1 U6034 ( .A1(n5008), .A2(n5011), .ZN(n8176) );
  AND2_X1 U6035 ( .A1(n8962), .A2(n8919), .ZN(n4534) );
  OR2_X1 U6036 ( .A1(n8043), .A2(n8110), .ZN(n4535) );
  AOI21_X1 U6037 ( .B1(n8455), .B2(n6169), .A(n4515), .ZN(n8414) );
  NAND2_X1 U6038 ( .A1(n6440), .A2(n8758), .ZN(n8686) );
  AND2_X1 U6039 ( .A1(n7089), .A2(n5034), .ZN(n4536) );
  AND2_X1 U6040 ( .A1(n9057), .A2(n4789), .ZN(n4537) );
  INV_X1 U6041 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5765) );
  AND4_X1 U6042 ( .A1(n5719), .A2(n5718), .A3(n5717), .A4(n5877), .ZN(n4538)
         );
  NOR3_X1 U6043 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n4539) );
  AND2_X1 U6044 ( .A1(n4759), .A2(n8410), .ZN(n4540) );
  NOR2_X1 U6045 ( .A1(n9287), .A2(n9284), .ZN(n4541) );
  AND3_X1 U6046 ( .A1(n5935), .A2(n5726), .A3(n5947), .ZN(n4542) );
  AND2_X1 U6047 ( .A1(n7097), .A2(n7044), .ZN(n4543) );
  NAND2_X1 U6048 ( .A1(n7943), .A2(n7793), .ZN(n7976) );
  INV_X1 U6049 ( .A(n8449), .ZN(n8444) );
  NAND2_X1 U6050 ( .A1(n7925), .A2(n7924), .ZN(n8449) );
  INV_X1 U6051 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4608) );
  NAND2_X1 U6052 ( .A1(n10089), .A2(n8234), .ZN(n4544) );
  AND2_X1 U6053 ( .A1(n5057), .A2(n4542), .ZN(n4545) );
  NAND2_X1 U6054 ( .A1(n8692), .A2(n4918), .ZN(n4917) );
  AND2_X1 U6055 ( .A1(n4910), .A2(n4617), .ZN(n4546) );
  INV_X1 U6056 ( .A(n5042), .ZN(n5041) );
  NOR2_X1 U6057 ( .A1(n5047), .A2(n8013), .ZN(n5042) );
  INV_X1 U6058 ( .A(n7524), .ZN(n4767) );
  NAND2_X1 U6059 ( .A1(n5197), .A2(n5778), .ZN(n4687) );
  AND2_X1 U6060 ( .A1(n4920), .A2(n4923), .ZN(n4547) );
  OR2_X1 U6061 ( .A1(n8240), .A2(n10062), .ZN(n7854) );
  OR2_X1 U6062 ( .A1(n7608), .A2(n7646), .ZN(n7870) );
  AND2_X1 U6063 ( .A1(n6855), .A2(n6854), .ZN(n4548) );
  INV_X1 U6064 ( .A(n5045), .ZN(n5044) );
  NAND2_X1 U6065 ( .A1(n5049), .A2(n8116), .ZN(n5045) );
  NOR2_X1 U6066 ( .A1(n7006), .A2(n4930), .ZN(n4549) );
  NOR2_X1 U6067 ( .A1(n7591), .A2(n6378), .ZN(n4550) );
  NOR2_X1 U6068 ( .A1(n8715), .A2(n7698), .ZN(n4551) );
  AND2_X1 U6069 ( .A1(n5613), .A2(n5612), .ZN(n9260) );
  AOI21_X1 U6070 ( .B1(n4681), .B2(n8894), .A(n8981), .ZN(n4679) );
  INV_X1 U6071 ( .A(n4959), .ZN(n4958) );
  NAND2_X1 U6072 ( .A1(n4960), .A2(n5544), .ZN(n4959) );
  AND2_X1 U6073 ( .A1(n5336), .A2(SI_12_), .ZN(n4552) );
  AND2_X1 U6074 ( .A1(n5318), .A2(n4897), .ZN(n4553) );
  OR2_X1 U6075 ( .A1(n5922), .A2(n5060), .ZN(n4554) );
  AND2_X1 U6076 ( .A1(n4724), .A2(n4722), .ZN(n4555) );
  NAND2_X1 U6077 ( .A1(n5013), .A2(n8177), .ZN(n4556) );
  INV_X1 U6078 ( .A(n6172), .ZN(n4805) );
  INV_X1 U6079 ( .A(n4705), .ZN(n4704) );
  AOI21_X1 U6080 ( .B1(n4709), .B2(n4707), .A(n7946), .ZN(n4705) );
  NAND2_X1 U6081 ( .A1(n7793), .A2(n7977), .ZN(n4557) );
  AND2_X1 U6082 ( .A1(n8628), .A2(n8436), .ZN(n4558) );
  NAND2_X1 U6083 ( .A1(n8421), .A2(n8225), .ZN(n4559) );
  AND2_X1 U6084 ( .A1(n8980), .A2(n8968), .ZN(n4560) );
  OR2_X1 U6085 ( .A1(n8407), .A2(n8395), .ZN(n7932) );
  AND2_X1 U6086 ( .A1(n4671), .A2(n4670), .ZN(n4561) );
  AND2_X1 U6087 ( .A1(n9260), .A2(n9073), .ZN(n8961) );
  INV_X1 U6088 ( .A(n8961), .ZN(n8985) );
  NAND2_X1 U6089 ( .A1(n5028), .A2(n5029), .ZN(n5753) );
  INV_X1 U6090 ( .A(n5105), .ZN(n4822) );
  NAND2_X1 U6091 ( .A1(n5102), .A2(n5101), .ZN(n5105) );
  INV_X1 U6092 ( .A(n5825), .ZN(n6110) );
  OR2_X1 U6093 ( .A1(n4532), .A2(n7947), .ZN(n4562) );
  NAND2_X1 U6094 ( .A1(n4903), .A2(n8737), .ZN(n4563) );
  INV_X1 U6095 ( .A(n9251), .ZN(n9518) );
  NAND2_X1 U6096 ( .A1(n8908), .A2(n8907), .ZN(n9251) );
  AND3_X1 U6097 ( .A1(n4516), .A2(n4539), .A3(n4755), .ZN(n4564) );
  AND2_X1 U6098 ( .A1(n8460), .A2(n7915), .ZN(n4565) );
  OR2_X1 U6099 ( .A1(n4675), .A2(n4677), .ZN(n4566) );
  AND2_X1 U6100 ( .A1(n8258), .A2(n8321), .ZN(n4567) );
  AND2_X1 U6101 ( .A1(n9311), .A2(n4646), .ZN(n4568) );
  OR2_X1 U6102 ( .A1(n6364), .A2(n7464), .ZN(n4569) );
  AND2_X1 U6103 ( .A1(n4512), .A2(n5417), .ZN(n4570) );
  NAND2_X1 U6104 ( .A1(n5121), .A2(n5120), .ZN(n5318) );
  NAND2_X1 U6105 ( .A1(n8107), .A2(n8041), .ZN(n4571) );
  AND2_X1 U6106 ( .A1(n4728), .A2(n4725), .ZN(n4572) );
  OR2_X1 U6107 ( .A1(n8385), .A2(n6172), .ZN(n4573) );
  NAND2_X1 U6108 ( .A1(n7237), .A2(n7245), .ZN(n4574) );
  AND2_X1 U6109 ( .A1(n4949), .A2(n4948), .ZN(n4575) );
  NAND2_X1 U6110 ( .A1(n8978), .A2(n8919), .ZN(n4576) );
  INV_X1 U6111 ( .A(n4753), .ZN(n4752) );
  OAI21_X1 U6112 ( .B1(n4754), .B2(n7891), .A(n7895), .ZN(n4753) );
  INV_X1 U6113 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4951) );
  INV_X1 U6114 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5153) );
  INV_X1 U6115 ( .A(n4729), .ZN(n4728) );
  NAND2_X1 U6116 ( .A1(n4562), .A2(n4730), .ZN(n4729) );
  XNOR2_X1 U6117 ( .A(n5690), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U6118 ( .A1(n6096), .A2(n6095), .ZN(n8066) );
  INV_X1 U6119 ( .A(n8066), .ZN(n4731) );
  INV_X1 U6120 ( .A(n9888), .ZN(n8305) );
  NOR2_X1 U6121 ( .A1(n5890), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U6122 ( .A1(n5462), .A2(n5461), .ZN(n9476) );
  INV_X1 U6123 ( .A(n9476), .ZN(n4773) );
  NAND2_X1 U6124 ( .A1(n7174), .A2(n7175), .ZN(n7173) );
  INV_X1 U6125 ( .A(n9092), .ZN(n6342) );
  INV_X1 U6126 ( .A(n9091), .ZN(n5316) );
  NAND2_X1 U6127 ( .A1(n5043), .A2(n5041), .ZN(n8078) );
  OAI21_X1 U6128 ( .B1(n8525), .B2(n8529), .A(n6154), .ZN(n8510) );
  NAND2_X1 U6129 ( .A1(n5623), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5408) );
  NAND2_X1 U6130 ( .A1(n5409), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U6131 ( .A1(n4967), .A2(n4970), .ZN(n9413) );
  AND2_X1 U6132 ( .A1(n8168), .A2(n8233), .ZN(n4577) );
  NAND2_X1 U6133 ( .A1(n4928), .A2(n5128), .ZN(n5356) );
  INV_X1 U6134 ( .A(n4832), .ZN(n4831) );
  NOR2_X1 U6135 ( .A1(n5508), .A2(n4833), .ZN(n4832) );
  INV_X1 U6136 ( .A(n4774), .ZN(n9391) );
  AND2_X1 U6137 ( .A1(n6584), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4578) );
  AND2_X1 U6138 ( .A1(n9367), .A2(n9080), .ZN(n4579) );
  OR2_X1 U6139 ( .A1(n8568), .A2(n8457), .ZN(n7925) );
  OR2_X1 U6140 ( .A1(n8045), .A2(n8227), .ZN(n4580) );
  OR2_X1 U6141 ( .A1(n9427), .A2(n7751), .ZN(n4581) );
  NOR2_X1 U6142 ( .A1(n8503), .A2(n8512), .ZN(n4582) );
  NOR2_X1 U6143 ( .A1(n8207), .A2(n5038), .ZN(n4583) );
  AND2_X1 U6144 ( .A1(n5435), .A2(SI_18_), .ZN(n4584) );
  INV_X1 U6145 ( .A(n6483), .ZN(n9527) );
  NAND2_X1 U6146 ( .A1(n5555), .A2(n5554), .ZN(n6483) );
  AND2_X1 U6147 ( .A1(n6483), .A2(n9076), .ZN(n4585) );
  AND2_X1 U6148 ( .A1(n5048), .A2(n5046), .ZN(n4586) );
  INV_X1 U6149 ( .A(n8226), .ZN(n8447) );
  INV_X1 U6150 ( .A(n6448), .ZN(n4904) );
  OR2_X1 U6151 ( .A1(n9888), .A2(n7451), .ZN(n4587) );
  NAND2_X1 U6152 ( .A1(n7946), .A2(n6903), .ZN(n10032) );
  NAND2_X1 U6153 ( .A1(n7090), .A2(n4536), .ZN(n5032) );
  INV_X1 U6154 ( .A(n8919), .ZN(n4789) );
  INV_X1 U6155 ( .A(n8717), .ZN(n4627) );
  NAND2_X1 U6156 ( .A1(n4618), .A2(n4910), .ZN(n7511) );
  NAND2_X1 U6157 ( .A1(n7434), .A2(n4915), .ZN(n7461) );
  INV_X1 U6158 ( .A(n7947), .ZN(n7946) );
  NAND2_X1 U6159 ( .A1(n7825), .A2(n7991), .ZN(n7947) );
  AND2_X1 U6160 ( .A1(n5032), .A2(n5031), .ZN(n4588) );
  AOI22_X1 U6161 ( .A1(n7041), .A2(n4543), .B1(n6314), .B2(n4524), .ZN(n7100)
         );
  AND2_X1 U6162 ( .A1(n7041), .A2(n7044), .ZN(n4589) );
  AND2_X1 U6163 ( .A1(n4941), .A2(n4940), .ZN(n4590) );
  NAND2_X1 U6164 ( .A1(n5141), .A2(n5156), .ZN(n5675) );
  OR2_X1 U6165 ( .A1(n7004), .A2(n10156), .ZN(n4934) );
  NAND2_X1 U6166 ( .A1(n7004), .A2(n10156), .ZN(n7005) );
  OR2_X1 U6167 ( .A1(n9985), .A2(n10323), .ZN(n4591) );
  INV_X1 U6168 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5796) );
  OR2_X1 U6169 ( .A1(n8340), .A2(n5995), .ZN(n4592) );
  INV_X1 U6170 ( .A(n8763), .ZN(n8780) );
  XNOR2_X1 U6171 ( .A(n8350), .B(n4594), .ZN(n4593) );
  NAND2_X1 U6172 ( .A1(n5720), .A2(n4538), .ZN(n5890) );
  INV_X1 U6173 ( .A(n8296), .ZN(n8342) );
  NAND2_X1 U6174 ( .A1(n9346), .A2(n9353), .ZN(n9347) );
  NAND2_X1 U6175 ( .A1(n4774), .A2(n4773), .ZN(n9363) );
  NAND2_X1 U6176 ( .A1(n9766), .A2(n7208), .ZN(n6803) );
  NOR2_X2 U6177 ( .A1(n7419), .A2(n9723), .ZN(n7587) );
  AOI211_X2 U6178 ( .C1(n9251), .C2(n9250), .A(n9422), .B(n9249), .ZN(n9435)
         );
  NAND2_X1 U6179 ( .A1(n6151), .A2(n6150), .ZN(n4801) );
  MUX2_X1 U6180 ( .A(n8549), .B(n8614), .S(n10105), .Z(n8550) );
  MUX2_X1 U6181 ( .A(n8615), .B(n8614), .S(n10091), .Z(n8616) );
  NAND2_X1 U6182 ( .A1(n8484), .A2(n6159), .ZN(n8483) );
  NAND2_X1 U6183 ( .A1(n5261), .A2(n5094), .ZN(n4641) );
  NAND2_X1 U6184 ( .A1(n4796), .A2(n4795), .ZN(n6171) );
  NAND2_X1 U6185 ( .A1(n4943), .A2(n9818), .ZN(n7002) );
  AND2_X1 U6186 ( .A1(n10014), .A2(n10013), .ZN(n4601) );
  INV_X1 U6187 ( .A(n4607), .ZN(n4606) );
  NAND2_X1 U6188 ( .A1(n8292), .A2(n8293), .ZN(n8296) );
  NAND2_X1 U6189 ( .A1(n5077), .A2(n5076), .ZN(n4682) );
  BUF_X2 U6190 ( .A(n7798), .Z(n4610) );
  NAND2_X1 U6191 ( .A1(n4875), .A2(n4879), .ZN(n9276) );
  NAND2_X1 U6192 ( .A1(n5093), .A2(n5092), .ZN(n5261) );
  NAND2_X1 U6193 ( .A1(n4818), .A2(n5099), .ZN(n5170) );
  NAND2_X1 U6194 ( .A1(n4683), .A2(n5089), .ZN(n5247) );
  OAI21_X1 U6195 ( .B1(n9358), .B2(n4884), .A(n4881), .ZN(n9330) );
  AOI21_X2 U6196 ( .B1(n5666), .B2(n9315), .A(n8980), .ZN(n9287) );
  NOR2_X1 U6197 ( .A1(n8773), .A2(n6495), .ZN(n7771) );
  NAND3_X1 U6198 ( .A1(n5064), .A2(n4612), .A3(n6263), .ZN(n6644) );
  NAND3_X1 U6199 ( .A1(n6440), .A2(n4616), .A3(n8758), .ZN(n4614) );
  INV_X1 U6200 ( .A(n7693), .ZN(n4624) );
  OAI21_X1 U6201 ( .B1(n4624), .B2(n4623), .A(n4625), .ZN(n8720) );
  NAND3_X1 U6202 ( .A1(n4928), .A2(n5128), .A3(n5129), .ZN(n5391) );
  NAND2_X1 U6203 ( .A1(n6826), .A2(n6310), .ZN(n4629) );
  NAND3_X1 U6204 ( .A1(n4633), .A2(n4632), .A3(n4630), .ZN(n10226) );
  NAND2_X1 U6205 ( .A1(n4810), .A2(n5459), .ZN(n5474) );
  NAND2_X1 U6206 ( .A1(n4810), .A2(n4527), .ZN(n4643) );
  INV_X2 U6207 ( .A(n7798), .ZN(n5082) );
  NAND2_X1 U6208 ( .A1(n4648), .A2(n4568), .ZN(n8892) );
  INV_X1 U6209 ( .A(n8890), .ZN(n4647) );
  NAND3_X1 U6210 ( .A1(n4652), .A2(n4649), .A3(n4576), .ZN(n4648) );
  NAND2_X1 U6211 ( .A1(n4653), .A2(n4650), .ZN(n4649) );
  NAND2_X1 U6212 ( .A1(n4653), .A2(n4779), .ZN(n4652) );
  NAND2_X1 U6213 ( .A1(n9012), .A2(n4654), .ZN(n4661) );
  NAND4_X1 U6214 ( .A1(n4657), .A2(n9069), .A3(n4655), .A4(n4511), .ZN(
        P1_U3242) );
  NAND2_X1 U6215 ( .A1(n4525), .A2(n4662), .ZN(n4658) );
  NAND2_X1 U6216 ( .A1(n5370), .A2(n4665), .ZN(n4664) );
  NAND2_X1 U6217 ( .A1(n5370), .A2(n5369), .ZN(n5373) );
  NAND3_X1 U6218 ( .A1(n8897), .A2(n8898), .A3(n4566), .ZN(n4671) );
  AND2_X1 U6219 ( .A1(n8893), .A2(n9274), .ZN(n4681) );
  NAND2_X1 U6220 ( .A1(n4682), .A2(n5078), .ZN(n5081) );
  XNOR2_X1 U6221 ( .A(n4682), .B(n5207), .ZN(n5786) );
  NAND2_X1 U6222 ( .A1(n5241), .A2(n5087), .ZN(n4683) );
  NAND2_X1 U6223 ( .A1(n5219), .A2(n5218), .ZN(n4684) );
  NAND2_X1 U6224 ( .A1(n7798), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4685) );
  NAND2_X1 U6225 ( .A1(n7798), .A2(n5073), .ZN(n5778) );
  NAND2_X1 U6226 ( .A1(n4706), .A2(n4565), .ZN(n4703) );
  OR2_X1 U6227 ( .A1(n7945), .A2(n4729), .ZN(n4724) );
  NAND2_X1 U6228 ( .A1(n4721), .A2(n4572), .ZN(n4855) );
  NAND2_X1 U6229 ( .A1(n7945), .A2(n4726), .ZN(n4721) );
  NAND4_X1 U6230 ( .A1(n5765), .A2(n5029), .A3(n4951), .A4(n4734), .ZN(n5755)
         );
  INV_X2 U6231 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5029) );
  NAND2_X1 U6232 ( .A1(n7849), .A2(n7835), .ZN(n7955) );
  INV_X1 U6233 ( .A(n7052), .ZN(n4739) );
  OAI211_X1 U6234 ( .C1(n4745), .C2(n4746), .A(n4743), .B(n7868), .ZN(n7506)
         );
  NAND2_X1 U6235 ( .A1(n4746), .A2(n5864), .ZN(n4744) );
  NOR2_X1 U6236 ( .A1(n4747), .A2(n7960), .ZN(n4746) );
  NAND2_X1 U6237 ( .A1(n4749), .A2(n4748), .ZN(n8461) );
  OAI21_X1 U6238 ( .B1(n9590), .B2(n4753), .A(n4750), .ZN(n7627) );
  OAI21_X1 U6239 ( .B1(n9590), .B2(n7892), .A(n7890), .ZN(n7555) );
  INV_X4 U6240 ( .A(n7790), .ZN(n7803) );
  AND3_X2 U6241 ( .A1(n4809), .A2(n5056), .A3(n4564), .ZN(n5751) );
  NAND4_X1 U6242 ( .A1(n4809), .A2(n5056), .A3(n4516), .A4(n4539), .ZN(n6199)
         );
  NAND3_X1 U6243 ( .A1(n4809), .A2(n5056), .A3(n4516), .ZN(n6190) );
  AOI21_X2 U6244 ( .B1(n8450), .B2(n4540), .A(n4757), .ZN(n8398) );
  INV_X1 U6245 ( .A(n7952), .ZN(n4763) );
  NAND3_X1 U6246 ( .A1(n4991), .A2(n4990), .A3(n4765), .ZN(n5144) );
  NOR2_X2 U6247 ( .A1(n6942), .A2(n6943), .ZN(n6941) );
  NOR2_X2 U6248 ( .A1(n7153), .A2(n9755), .ZN(n7208) );
  NAND2_X1 U6249 ( .A1(n9270), .A2(n4770), .ZN(n9248) );
  NAND2_X1 U6250 ( .A1(n9270), .A2(n9260), .ZN(n6550) );
  NOR2_X2 U6251 ( .A1(n9363), .A2(n9367), .ZN(n9346) );
  NAND2_X1 U6252 ( .A1(n5664), .A2(n8885), .ZN(n4777) );
  NAND2_X2 U6253 ( .A1(n4786), .A2(n5189), .ZN(n7153) );
  INV_X1 U6254 ( .A(n4787), .ZN(n4786) );
  NAND2_X1 U6255 ( .A1(n4790), .A2(n6124), .ZN(n7055) );
  XNOR2_X1 U6256 ( .A(n4790), .B(n7955), .ZN(n7119) );
  NOR2_X1 U6257 ( .A1(n8375), .A2(n4794), .ZN(n8544) );
  NAND2_X1 U6258 ( .A1(n8455), .A2(n4797), .ZN(n4796) );
  INV_X1 U6259 ( .A(n6171), .ZN(n8404) );
  INV_X1 U6260 ( .A(n8393), .ZN(n4806) );
  OAI21_X1 U6261 ( .B1(n8393), .B2(n4573), .A(n4803), .ZN(n7999) );
  AOI21_X2 U6262 ( .B1(n6157), .B2(n4807), .A(n4582), .ZN(n8484) );
  NAND2_X1 U6263 ( .A1(n5474), .A2(n5473), .ZN(n5475) );
  NAND2_X1 U6264 ( .A1(n4811), .A2(n5458), .ZN(n4810) );
  INV_X1 U6265 ( .A(n6104), .ZN(n4816) );
  NAND2_X2 U6266 ( .A1(n4817), .A2(n4820), .ZN(n5112) );
  OAI21_X1 U6267 ( .B1(n5492), .B2(n4828), .A(n4826), .ZN(n5571) );
  NAND2_X1 U6268 ( .A1(n5319), .A2(n4845), .ZN(n4844) );
  NAND2_X1 U6269 ( .A1(n4844), .A2(n4846), .ZN(n5370) );
  MUX2_X1 U6270 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5082), .Z(n5079) );
  OAI211_X1 U6271 ( .C1(n4555), .C2(n7947), .A(n7949), .B(n4853), .ZN(n7985)
         );
  NAND2_X1 U6272 ( .A1(n4855), .A2(n4854), .ZN(n4853) );
  AND2_X1 U6273 ( .A1(n7978), .A2(n7947), .ZN(n4854) );
  AOI21_X1 U6274 ( .B1(n5571), .B2(n5570), .A(n5068), .ZN(n5586) );
  NAND2_X1 U6275 ( .A1(n5185), .A2(SI_1_), .ZN(n5077) );
  NAND2_X1 U6276 ( .A1(n5588), .A2(n5587), .ZN(n5595) );
  NAND2_X1 U6277 ( .A1(n4898), .A2(n5115), .ZN(n5319) );
  OR2_X2 U6278 ( .A1(n8245), .A2(n10047), .ZN(n7820) );
  NAND2_X2 U6279 ( .A1(n8475), .A2(n8474), .ZN(n8473) );
  NAND2_X1 U6280 ( .A1(n5082), .A2(n5074), .ZN(n5197) );
  NAND2_X1 U6281 ( .A1(n4856), .A2(n7582), .ZN(n5655) );
  XNOR2_X1 U6282 ( .A(n4858), .B(n8941), .ZN(n7656) );
  OAI21_X1 U6283 ( .B1(n7734), .B2(n4861), .A(n4859), .ZN(n7747) );
  NAND2_X1 U6284 ( .A1(n5656), .A2(n8817), .ZN(n4861) );
  INV_X1 U6285 ( .A(n8943), .ZN(n4863) );
  NAND3_X1 U6286 ( .A1(n8957), .A2(n4876), .A3(n9287), .ZN(n4867) );
  OAI211_X1 U6287 ( .C1(n4872), .C2(n9287), .A(n4868), .B(n4867), .ZN(n6560)
         );
  NAND2_X1 U6288 ( .A1(n9287), .A2(n9274), .ZN(n4875) );
  AOI21_X2 U6289 ( .B1(n4876), .B2(n4878), .A(n8961), .ZN(n4874) );
  AND2_X2 U6290 ( .A1(n4877), .A2(n8898), .ZN(n4876) );
  NAND2_X1 U6291 ( .A1(n5112), .A2(n4889), .ZN(n4887) );
  NAND2_X1 U6292 ( .A1(n5112), .A2(n4892), .ZN(n4888) );
  OAI211_X1 U6293 ( .C1(n5112), .C2(n4891), .A(n8910), .B(n4887), .ZN(n5326)
         );
  NAND2_X1 U6294 ( .A1(n5112), .A2(n4899), .ZN(n4898) );
  NAND2_X1 U6295 ( .A1(n5112), .A2(n5111), .ZN(n5304) );
  INV_X1 U6296 ( .A(n5629), .ZN(n5680) );
  INV_X4 U6297 ( .A(n6266), .ZN(n6496) );
  INV_X1 U6298 ( .A(n6400), .ZN(n6403) );
  NAND2_X1 U6299 ( .A1(n8692), .A2(n6464), .ZN(n6469) );
  AND4_X2 U6300 ( .A1(n5122), .A2(n5123), .A3(n5208), .A4(n5233), .ZN(n4928)
         );
  INV_X1 U6301 ( .A(n4929), .ZN(n8247) );
  INV_X1 U6302 ( .A(n4935), .ZN(n9961) );
  NOR2_X1 U6303 ( .A1(n9947), .A2(n4567), .ZN(n9963) );
  INV_X1 U6304 ( .A(n4941), .ZN(n9880) );
  INV_X1 U6305 ( .A(n8252), .ZN(n4940) );
  INV_X1 U6306 ( .A(n4949), .ZN(n10012) );
  INV_X1 U6307 ( .A(n8263), .ZN(n4948) );
  NAND3_X1 U6308 ( .A1(n5122), .A2(n5208), .A3(n5233), .ZN(n5262) );
  NAND2_X1 U6309 ( .A1(n5507), .A2(n4955), .ZN(n4954) );
  AOI21_X1 U6310 ( .B1(n7703), .B2(n4570), .A(n4968), .ZN(n9398) );
  NAND2_X1 U6311 ( .A1(n9709), .A2(n4977), .ZN(n4974) );
  NAND2_X1 U6312 ( .A1(n4974), .A2(n4975), .ZN(n7654) );
  NAND2_X1 U6313 ( .A1(n9268), .A2(n9275), .ZN(n4984) );
  NAND2_X1 U6314 ( .A1(n4984), .A2(n5604), .ZN(n5622) );
  NAND2_X1 U6315 ( .A1(n5140), .A2(n5139), .ZN(n5156) );
  NAND2_X1 U6316 ( .A1(n5140), .A2(n4985), .ZN(n5155) );
  NAND2_X1 U6317 ( .A1(n9374), .A2(n4988), .ZN(n4987) );
  INV_X1 U6318 ( .A(n5356), .ZN(n4991) );
  OAI21_X1 U6319 ( .B1(n7183), .B2(n4994), .A(n4992), .ZN(n7348) );
  INV_X1 U6320 ( .A(n4999), .ZN(n7278) );
  NAND2_X1 U6321 ( .A1(n8089), .A2(n5002), .ZN(n5005) );
  NAND3_X1 U6322 ( .A1(n5005), .A2(n8051), .A3(n5003), .ZN(n8126) );
  NAND2_X1 U6323 ( .A1(n5006), .A2(n8049), .ZN(n8151) );
  NAND2_X1 U6324 ( .A1(n8089), .A2(n8447), .ZN(n5006) );
  NOR2_X1 U6325 ( .A1(n5009), .A2(n5007), .ZN(n8046) );
  NAND2_X1 U6326 ( .A1(n8198), .A2(n5016), .ZN(n5015) );
  OAI211_X1 U6327 ( .C1(n8198), .C2(n5021), .A(n5018), .B(n5015), .ZN(n8068)
         );
  NAND2_X1 U6328 ( .A1(n8198), .A2(n8195), .ZN(n5022) );
  INV_X1 U6329 ( .A(n7163), .ZN(n5034) );
  INV_X1 U6330 ( .A(n8013), .ZN(n5049) );
  NAND2_X1 U6331 ( .A1(n5974), .A2(n5053), .ZN(n5051) );
  INV_X1 U6332 ( .A(n7956), .ZN(n10025) );
  XNOR2_X1 U6333 ( .A(n8000), .B(n8060), .ZN(n8004) );
  NAND2_X1 U6334 ( .A1(n6280), .A2(n6279), .ZN(n6748) );
  OAI21_X1 U6335 ( .B1(n7954), .B2(n7824), .A(n7820), .ZN(n10020) );
  OAI22_X1 U6336 ( .A1(n7998), .A2(n8060), .B1(n8383), .B2(n8066), .ZN(n7784)
         );
  NAND2_X1 U6337 ( .A1(n7954), .A2(n7139), .ZN(n10026) );
  OR2_X1 U6338 ( .A1(n7217), .A2(n10095), .ZN(n5763) );
  NAND2_X1 U6339 ( .A1(n6766), .A2(n6293), .ZN(n6815) );
  NOR2_X1 U6340 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5122) );
  INV_X1 U6341 ( .A(n6436), .ZN(n6439) );
  NAND2_X2 U6342 ( .A1(n8473), .A2(n6161), .ZN(n8455) );
  INV_X1 U6343 ( .A(n7217), .ZN(n6068) );
  NAND2_X1 U6344 ( .A1(n6808), .A2(n6807), .ZN(n6806) );
  AOI21_X1 U6345 ( .B1(n7776), .B2(n7775), .A(n7774), .ZN(n7783) );
  INV_X1 U6346 ( .A(n5755), .ZN(n5720) );
  INV_X1 U6347 ( .A(n6277), .ZN(n6280) );
  INV_X1 U6348 ( .A(n4505), .ZN(n6320) );
  INV_X1 U6349 ( .A(n9543), .ZN(n6562) );
  AND2_X1 U6350 ( .A1(n8012), .A2(n8234), .ZN(n5059) );
  OR2_X1 U6351 ( .A1(n5733), .A2(n5732), .ZN(n5060) );
  AND3_X1 U6352 ( .A1(n6536), .A2(n8775), .A3(n6535), .ZN(n5061) );
  NOR2_X1 U6353 ( .A1(n8368), .A2(n8662), .ZN(n5062) );
  AND4_X1 U6354 ( .A1(n5628), .A2(n5707), .A3(n5681), .A4(n10370), .ZN(n5063)
         );
  OR2_X1 U6355 ( .A1(n6261), .A2(n6264), .ZN(n5064) );
  INV_X1 U6356 ( .A(n8955), .ZN(n5667) );
  NAND2_X1 U6357 ( .A1(n8985), .A2(n6553), .ZN(n8955) );
  AND2_X1 U6358 ( .A1(n5111), .A2(n5110), .ZN(n5065) );
  INV_X1 U6359 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5174) );
  AND2_X1 U6360 ( .A1(n10035), .A2(n10034), .ZN(n8536) );
  AND2_X1 U6361 ( .A1(n6574), .A2(n6573), .ZN(n5066) );
  AND2_X1 U6362 ( .A1(n6564), .A2(n6563), .ZN(n5067) );
  INV_X1 U6363 ( .A(n9260), .ZN(n6539) );
  NOR2_X1 U6364 ( .A1(n7417), .A2(n5317), .ZN(n9709) );
  INV_X1 U6365 ( .A(n5220), .ZN(n5289) );
  NOR2_X1 U6366 ( .A1(n5569), .A2(n5568), .ZN(n5068) );
  NOR2_X1 U6367 ( .A1(n5136), .A2(n5135), .ZN(n5137) );
  INV_X1 U6368 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5123) );
  AND2_X1 U6369 ( .A1(n8203), .A2(n8224), .ZN(n6172) );
  OR2_X1 U6370 ( .A1(n6149), .A2(n6148), .ZN(n6150) );
  AND2_X1 U6371 ( .A1(n8994), .A2(n8963), .ZN(n9053) );
  INV_X1 U6372 ( .A(n9088), .ZN(n8846) );
  OR2_X1 U6373 ( .A1(n7595), .A2(n7606), .ZN(n7596) );
  NAND2_X1 U6374 ( .A1(n8621), .A2(n8406), .ZN(n6173) );
  OR2_X1 U6375 ( .A1(n5862), .A2(n5861), .ZN(n5863) );
  INV_X1 U6376 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5906) );
  INV_X1 U6377 ( .A(n6278), .ZN(n6279) );
  AND2_X1 U6378 ( .A1(n9581), .A2(n6724), .ZN(n9614) );
  INV_X1 U6379 ( .A(n9267), .ZN(n9275) );
  NAND2_X1 U6380 ( .A1(n7591), .A2(n6378), .ZN(n5334) );
  NOR2_X1 U6381 ( .A1(n9098), .A2(n4768), .ZN(n5647) );
  INV_X1 U6382 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5682) );
  INV_X1 U6383 ( .A(n5400), .ZN(n5401) );
  INV_X1 U6384 ( .A(n5275), .ZN(n5097) );
  AND2_X1 U6385 ( .A1(n6896), .A2(n8245), .ZN(n6897) );
  NAND2_X1 U6386 ( .A1(n7002), .A2(n9816), .ZN(n9820) );
  NAND2_X1 U6387 ( .A1(n8260), .A2(n8324), .ZN(n8261) );
  AOI21_X1 U6388 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8302), .A(n9994), .ZN(
        n8262) );
  AND2_X1 U6389 ( .A1(n6507), .A2(n6506), .ZN(n7772) );
  INV_X1 U6390 ( .A(n6437), .ZN(n6438) );
  OR2_X1 U6391 ( .A1(n8771), .A2(n8772), .ZN(n6495) );
  OR2_X1 U6392 ( .A1(n5480), .A2(n5479), .ZN(n5499) );
  OR2_X1 U6393 ( .A1(n9579), .A2(n9578), .ZN(n9581) );
  OR2_X1 U6394 ( .A1(n9697), .A2(n9696), .ZN(n9700) );
  OR2_X1 U6395 ( .A1(n9568), .A2(n6545), .ZN(n6547) );
  INV_X1 U6396 ( .A(n9093), .ZN(n5288) );
  INV_X1 U6397 ( .A(n9469), .ZN(n6572) );
  INV_X1 U6398 ( .A(n8990), .ZN(n8904) );
  NAND2_X1 U6399 ( .A1(n5455), .A2(n5454), .ZN(n9374) );
  INV_X1 U6400 ( .A(n9756), .ZN(n6524) );
  OR2_X1 U6401 ( .A1(n7787), .A2(n7786), .ZN(n7788) );
  INV_X1 U6402 ( .A(n5335), .ZN(n5337) );
  OR2_X1 U6403 ( .A1(n8008), .A2(n8118), .ZN(n8009) );
  NAND2_X1 U6404 ( .A1(n5748), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U6405 ( .A1(n9978), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n9977) );
  INV_X1 U6406 ( .A(n8222), .ZN(n8383) );
  NAND2_X1 U6407 ( .A1(n7506), .A2(n7964), .ZN(n7505) );
  OR2_X1 U6408 ( .A1(n7947), .A2(n6119), .ZN(n6904) );
  INV_X1 U6409 ( .A(n8232), .ZN(n9598) );
  AND2_X1 U6410 ( .A1(n7986), .A2(n6239), .ZN(n10041) );
  AND2_X1 U6411 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5252) );
  NAND2_X1 U6412 ( .A1(n5446), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5480) );
  NAND2_X1 U6413 ( .A1(n6439), .A2(n6438), .ZN(n8758) );
  NOR2_X1 U6414 ( .A1(n6494), .A2(n6493), .ZN(n8772) );
  AND2_X1 U6415 ( .A1(n5670), .A2(n5617), .ZN(n9258) );
  AND2_X1 U6416 ( .A1(n5427), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5446) );
  OR2_X1 U6417 ( .A1(n6700), .A2(n6699), .ZN(n6721) );
  NAND2_X1 U6418 ( .A1(n8786), .A2(n8895), .ZN(n5583) );
  INV_X1 U6419 ( .A(n9467), .ZN(n9353) );
  AND2_X1 U6420 ( .A1(n8867), .A2(n8876), .ZN(n9417) );
  NAND2_X1 U6421 ( .A1(n5327), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5329) );
  AOI21_X1 U6422 ( .B1(n9398), .B2(n5432), .A(n5431), .ZN(n9386) );
  OAI22_X1 U6423 ( .A1(n7732), .A2(n5367), .B1(n8821), .B2(n9506), .ZN(n7703)
         );
  INV_X1 U6424 ( .A(n7375), .ZN(n7372) );
  NAND2_X1 U6425 ( .A1(n6927), .A2(n6926), .ZN(n6929) );
  NAND2_X1 U6426 ( .A1(n5153), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5158) );
  INV_X1 U6427 ( .A(n8212), .ZN(n8187) );
  AND2_X1 U6428 ( .A1(n6094), .A2(n6093), .ZN(n8396) );
  AND3_X1 U6429 ( .A1(n6020), .A2(n6019), .A3(n6018), .ZN(n8456) );
  INV_X1 U6430 ( .A(n10140), .ZN(n10010) );
  AND2_X1 U6431 ( .A1(n6787), .A2(n8291), .ZN(n10153) );
  NAND2_X1 U6432 ( .A1(n6884), .A2(n6883), .ZN(n10022) );
  INV_X1 U6433 ( .A(n10041), .ZN(n8516) );
  AND2_X1 U6434 ( .A1(n6230), .A2(n6229), .ZN(n6231) );
  AND2_X1 U6435 ( .A1(n8360), .A2(n8359), .ZN(n8606) );
  AND2_X1 U6436 ( .A1(n6222), .A2(n6221), .ZN(n7069) );
  INV_X1 U6437 ( .A(n5202), .ZN(n5521) );
  INV_X1 U6438 ( .A(n9649), .ZN(n9699) );
  AND2_X1 U6439 ( .A1(n5677), .A2(n9266), .ZN(n5678) );
  INV_X1 U6440 ( .A(n8950), .ZN(n9331) );
  AND2_X1 U6441 ( .A1(n9788), .A2(n9768), .ZN(n7714) );
  MUX2_X1 U6442 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9573), .S(n6612), .Z(n9755) );
  AND2_X1 U6443 ( .A1(n5324), .A2(n5339), .ZN(n9607) );
  XNOR2_X1 U6444 ( .A(n5090), .B(SI_5_), .ZN(n5246) );
  INV_X1 U6445 ( .A(n8199), .ZN(n8214) );
  AND2_X1 U6446 ( .A1(n6880), .A2(n6879), .ZN(n8206) );
  AND2_X1 U6447 ( .A1(n7226), .A2(n6116), .ZN(n8062) );
  INV_X1 U6448 ( .A(n8457), .ZN(n8227) );
  NAND2_X1 U6449 ( .A1(n7077), .A2(n10022), .ZN(n10035) );
  AOI21_X1 U6450 ( .B1(n6232), .B2(n8539), .A(n6234), .ZN(n6235) );
  NAND2_X1 U6451 ( .A1(n10105), .A2(n10090), .ZN(n8604) );
  INV_X1 U6452 ( .A(n10105), .ZN(n10103) );
  OR2_X1 U6453 ( .A1(n10093), .A2(n10077), .ZN(n8662) );
  AND2_X1 U6454 ( .A1(n6246), .A2(n6245), .ZN(n10093) );
  INV_X1 U6455 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10453) );
  INV_X1 U6456 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6597) );
  AND2_X1 U6457 ( .A1(n7612), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6579) );
  INV_X1 U6458 ( .A(n9494), .ZN(n9427) );
  INV_X1 U6459 ( .A(n8845), .ZN(n8849) );
  INV_X1 U6460 ( .A(n8767), .ZN(n8785) );
  INV_X1 U6461 ( .A(n9670), .ZN(n9708) );
  NAND2_X1 U6462 ( .A1(n9409), .A2(n7031), .ZN(n9737) );
  AND2_X1 U6463 ( .A1(n7032), .A2(n9405), .ZN(n9744) );
  INV_X1 U6464 ( .A(n7727), .ZN(n9484) );
  INV_X1 U6465 ( .A(n9797), .ZN(n9795) );
  NAND2_X1 U6466 ( .A1(n9786), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5715) );
  INV_X1 U6467 ( .A(n7714), .ZN(n9555) );
  INV_X1 U6468 ( .A(n9788), .ZN(n9786) );
  AND2_X1 U6469 ( .A1(n6579), .A2(n6261), .ZN(n9749) );
  INV_X1 U6470 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6641) );
  INV_X1 U6471 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10284) );
  INV_X1 U6472 ( .A(n8297), .ZN(P2_U3893) );
  NAND2_X1 U6473 ( .A1(n5716), .A2(n5715), .ZN(P1_U3518) );
  AND2_X1 U6474 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5073) );
  AND2_X1 U6475 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5074) );
  NAND2_X1 U6476 ( .A1(n5075), .A2(n4687), .ZN(n5076) );
  INV_X1 U6477 ( .A(n5207), .ZN(n5078) );
  NAND2_X1 U6478 ( .A1(n5079), .A2(SI_2_), .ZN(n5080) );
  NAND2_X1 U6479 ( .A1(n5081), .A2(n5080), .ZN(n5219) );
  INV_X1 U6480 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n5083) );
  MUX2_X1 U6481 ( .A(n6587), .B(n5083), .S(n5082), .Z(n5084) );
  INV_X1 U6482 ( .A(n5084), .ZN(n5085) );
  NAND2_X1 U6483 ( .A1(n5085), .A2(SI_3_), .ZN(n5086) );
  MUX2_X1 U6484 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5082), .Z(n5088) );
  NAND2_X1 U6485 ( .A1(n5088), .A2(SI_4_), .ZN(n5089) );
  MUX2_X1 U6486 ( .A(n6597), .B(n10271), .S(n6584), .Z(n5090) );
  NAND2_X1 U6487 ( .A1(n5247), .A2(n5246), .ZN(n5093) );
  INV_X1 U6488 ( .A(n5090), .ZN(n5091) );
  NAND2_X1 U6489 ( .A1(n5091), .A2(SI_5_), .ZN(n5092) );
  MUX2_X1 U6490 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6584), .Z(n5095) );
  NAND2_X1 U6491 ( .A1(n5095), .A2(SI_6_), .ZN(n5096) );
  MUX2_X1 U6492 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6584), .Z(n5098) );
  NAND2_X1 U6493 ( .A1(n5098), .A2(SI_7_), .ZN(n5099) );
  INV_X1 U6494 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5100) );
  MUX2_X1 U6495 ( .A(n10288), .B(n5100), .S(n6584), .Z(n5102) );
  INV_X1 U6496 ( .A(SI_8_), .ZN(n5101) );
  INV_X1 U6497 ( .A(n5102), .ZN(n5103) );
  NAND2_X1 U6498 ( .A1(n5103), .A2(SI_8_), .ZN(n5104) );
  INV_X1 U6499 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5106) );
  MUX2_X1 U6500 ( .A(n6639), .B(n5106), .S(n6584), .Z(n5108) );
  INV_X1 U6501 ( .A(SI_9_), .ZN(n5107) );
  INV_X1 U6502 ( .A(n5108), .ZN(n5109) );
  NAND2_X1 U6503 ( .A1(n5109), .A2(SI_9_), .ZN(n5110) );
  MUX2_X1 U6504 ( .A(n6642), .B(n6641), .S(n6584), .Z(n5113) );
  INV_X1 U6505 ( .A(n5113), .ZN(n5114) );
  INV_X1 U6506 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5117) );
  MUX2_X1 U6507 ( .A(n10453), .B(n5117), .S(n6584), .Z(n5118) );
  INV_X1 U6508 ( .A(SI_11_), .ZN(n10451) );
  INV_X1 U6509 ( .A(n5118), .ZN(n5119) );
  NAND2_X1 U6510 ( .A1(n5119), .A2(SI_11_), .ZN(n5120) );
  MUX2_X1 U6511 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6584), .Z(n5336) );
  INV_X1 U6512 ( .A(SI_12_), .ZN(n10325) );
  XNOR2_X1 U6513 ( .A(n5338), .B(n5335), .ZN(n6776) );
  NOR2_X2 U6514 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5208) );
  NOR2_X2 U6515 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5233) );
  NOR2_X1 U6516 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5127) );
  NOR2_X1 U6517 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5126) );
  NOR2_X1 U6518 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5125) );
  NOR2_X1 U6519 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5133) );
  NOR2_X1 U6520 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5132) );
  NOR2_X1 U6521 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5131) );
  NOR2_X1 U6522 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5130) );
  NAND4_X1 U6523 ( .A1(n5133), .A2(n5132), .A3(n5131), .A4(n5130), .ZN(n5136)
         );
  INV_X2 U6524 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10370) );
  INV_X1 U6525 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5134) );
  NAND4_X1 U6526 ( .A1(n10370), .A2(n5682), .A3(n10354), .A4(n5134), .ZN(n5135) );
  NAND2_X1 U6527 ( .A1(n5144), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5138) );
  MUX2_X1 U6528 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5138), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5141) );
  INV_X1 U6529 ( .A(n5144), .ZN(n5140) );
  INV_X1 U6530 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5139) );
  NAND2_X1 U6531 ( .A1(n5142), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U6532 ( .A1(n6776), .A2(n8910), .ZN(n5152) );
  NOR2_X1 U6533 ( .A1(n5146), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5171) );
  NOR2_X1 U6534 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5147) );
  AND2_X1 U6535 ( .A1(n5171), .A2(n5147), .ZN(n5305) );
  INV_X1 U6536 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5148) );
  AND2_X1 U6537 ( .A1(n5305), .A2(n5148), .ZN(n5320) );
  INV_X1 U6538 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5149) );
  NAND2_X1 U6539 ( .A1(n5320), .A2(n5149), .ZN(n5339) );
  NAND2_X1 U6540 ( .A1(n5339), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5150) );
  XNOR2_X1 U6541 ( .A(n5150), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9216) );
  AOI22_X1 U6542 ( .A1(n8906), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5443), .B2(
        n9216), .ZN(n5151) );
  INV_X1 U6543 ( .A(n5164), .ZN(n7996) );
  NAND2_X1 U6544 ( .A1(n5156), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5157) );
  NAND2_X1 U6545 ( .A1(n5157), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n5159) );
  NAND2_X1 U6546 ( .A1(n5159), .A2(n5158), .ZN(n5160) );
  NAND2_X1 U6547 ( .A1(n5155), .A2(n5160), .ZN(n9567) );
  INV_X1 U6548 ( .A(n9567), .ZN(n5161) );
  NAND2_X1 U6549 ( .A1(n5201), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U6550 ( .A1(n5200), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6551 ( .A1(n5280), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5282) );
  INV_X1 U6552 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5162) );
  NAND2_X1 U6553 ( .A1(n5329), .A2(n5162), .ZN(n5163) );
  AND2_X1 U6554 ( .A1(n5344), .A2(n5163), .ZN(n7588) );
  NAND2_X1 U6555 ( .A1(n5202), .A2(n7588), .ZN(n5166) );
  NAND2_X1 U6556 ( .A1(n5164), .A2(n9567), .ZN(n5180) );
  INV_X2 U6557 ( .A(n5180), .ZN(n6554) );
  NAND2_X1 U6558 ( .A1(n6554), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5165) );
  NAND4_X1 U6559 ( .A1(n5168), .A2(n5167), .A3(n5166), .A4(n5165), .ZN(n9089)
         );
  INV_X1 U6560 ( .A(n9089), .ZN(n6378) );
  XNOR2_X1 U6561 ( .A(n5170), .B(n5169), .ZN(n6618) );
  NAND2_X1 U6562 ( .A1(n6618), .A2(n8910), .ZN(n5173) );
  OR2_X1 U6563 ( .A1(n5171), .A2(n5322), .ZN(n5291) );
  XNOR2_X1 U6564 ( .A(n5291), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9199) );
  AOI22_X1 U6565 ( .A1(n8906), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5443), .B2(
        n9199), .ZN(n5172) );
  NAND2_X2 U6566 ( .A1(n5173), .A2(n5172), .ZN(n7375) );
  NAND2_X1 U6567 ( .A1(n6554), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5179) );
  NAND2_X1 U6568 ( .A1(n5201), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5178) );
  NAND2_X1 U6569 ( .A1(n5282), .A2(n5174), .ZN(n5175) );
  AND2_X1 U6570 ( .A1(n5296), .A2(n5175), .ZN(n7328) );
  NAND2_X1 U6571 ( .A1(n5202), .A2(n7328), .ZN(n5177) );
  NAND2_X1 U6572 ( .A1(n5200), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5176) );
  NAND4_X1 U6573 ( .A1(n5179), .A2(n5178), .A3(n5177), .A4(n5176), .ZN(n9093)
         );
  INV_X1 U6574 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6663) );
  NAND2_X1 U6575 ( .A1(n5202), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5182) );
  NAND4_X2 U6576 ( .A1(n5184), .A2(n5183), .A3(n5182), .A4(n5181), .ZN(n6276)
         );
  XNOR2_X1 U6577 ( .A(n5185), .B(SI_1_), .ZN(n6586) );
  NAND2_X1 U6578 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5186) );
  XNOR2_X1 U6579 ( .A(n5186), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9105) );
  INV_X1 U6580 ( .A(n9105), .ZN(n5187) );
  NAND2_X1 U6581 ( .A1(n5213), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U6582 ( .A1(n5200), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5193) );
  NAND2_X1 U6583 ( .A1(n5202), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6584 ( .A1(n5201), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5191) );
  NAND4_X1 U6585 ( .A1(n5194), .A2(n5193), .A3(n5192), .A4(n5191), .ZN(n6265)
         );
  INV_X1 U6586 ( .A(SI_0_), .ZN(n5196) );
  INV_X1 U6587 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5195) );
  OAI21_X1 U6588 ( .B1(n4610), .B2(n5196), .A(n5195), .ZN(n5198) );
  AND2_X1 U6589 ( .A1(n5198), .A2(n5197), .ZN(n9573) );
  NAND2_X1 U6590 ( .A1(n6265), .A2(n9755), .ZN(n7152) );
  NAND2_X1 U6591 ( .A1(n5642), .A2(n7152), .ZN(n7151) );
  INV_X1 U6592 ( .A(n6276), .ZN(n5643) );
  NAND2_X1 U6593 ( .A1(n5643), .A2(n5190), .ZN(n5199) );
  NAND2_X1 U6594 ( .A1(n7151), .A2(n5199), .ZN(n7206) );
  NAND2_X1 U6595 ( .A1(n5200), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5206) );
  NAND2_X1 U6596 ( .A1(n5202), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5204) );
  NAND2_X1 U6597 ( .A1(n5213), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5203) );
  INV_X1 U6598 ( .A(n5786), .ZN(n6589) );
  NAND2_X1 U6599 ( .A1(n5220), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5210) );
  OR2_X1 U6600 ( .A1(n5208), .A2(n5322), .ZN(n5235) );
  XNOR2_X1 U6601 ( .A(n5235), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9118) );
  NAND2_X1 U6602 ( .A1(n5443), .A2(n9118), .ZN(n5209) );
  OAI211_X2 U6603 ( .C1(n6545), .C2(n6589), .A(n5210), .B(n5209), .ZN(n6772)
         );
  XNOR2_X1 U6604 ( .A(n6285), .B(n6772), .ZN(n8930) );
  INV_X1 U6605 ( .A(n8930), .ZN(n7207) );
  NAND2_X1 U6606 ( .A1(n7206), .A2(n7207), .ZN(n5212) );
  INV_X1 U6607 ( .A(n6285), .ZN(n6752) );
  NAND2_X1 U6608 ( .A1(n6752), .A2(n9766), .ZN(n5211) );
  NAND2_X1 U6609 ( .A1(n5212), .A2(n5211), .ZN(n6808) );
  INV_X1 U6610 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7127) );
  NAND2_X1 U6611 ( .A1(n5202), .A2(n7127), .ZN(n5217) );
  NAND2_X1 U6612 ( .A1(n5201), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U6613 ( .A1(n5200), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5215) );
  NAND2_X1 U6614 ( .A1(n5213), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5214) );
  XNOR2_X1 U6615 ( .A(n5219), .B(n5218), .ZN(n6591) );
  NAND2_X1 U6616 ( .A1(n5220), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5225) );
  INV_X1 U6617 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5221) );
  NAND2_X1 U6618 ( .A1(n5235), .A2(n5221), .ZN(n5222) );
  NAND2_X1 U6619 ( .A1(n5222), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5223) );
  XNOR2_X1 U6620 ( .A(n5223), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9131) );
  NAND2_X1 U6621 ( .A1(n5443), .A2(n9131), .ZN(n5224) );
  OAI211_X1 U6622 ( .C1(n6545), .C2(n6591), .A(n5225), .B(n5224), .ZN(n6804)
         );
  INV_X1 U6623 ( .A(n5647), .ZN(n8927) );
  NAND2_X1 U6624 ( .A1(n9098), .A2(n4768), .ZN(n9026) );
  NAND2_X1 U6625 ( .A1(n8927), .A2(n9026), .ZN(n6807) );
  INV_X1 U6626 ( .A(n9098), .ZN(n5226) );
  NAND2_X1 U6627 ( .A1(n5226), .A2(n4768), .ZN(n5227) );
  NAND2_X1 U6628 ( .A1(n6806), .A2(n5227), .ZN(n6939) );
  NAND2_X1 U6629 ( .A1(n6554), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5232) );
  NAND2_X1 U6630 ( .A1(n5201), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5231) );
  NOR2_X1 U6631 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5228) );
  NOR2_X1 U6632 ( .A1(n5252), .A2(n5228), .ZN(n9734) );
  NAND2_X1 U6633 ( .A1(n5202), .A2(n9734), .ZN(n5230) );
  NAND2_X1 U6634 ( .A1(n5200), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5229) );
  INV_X1 U6635 ( .A(n9097), .ZN(n5244) );
  OR2_X1 U6636 ( .A1(n5233), .A2(n5322), .ZN(n5234) );
  AND2_X1 U6637 ( .A1(n5235), .A2(n5234), .ZN(n5237) );
  INV_X1 U6638 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5236) );
  NAND2_X1 U6639 ( .A1(n5237), .A2(n5236), .ZN(n5248) );
  INV_X1 U6640 ( .A(n5237), .ZN(n5238) );
  NAND2_X1 U6641 ( .A1(n5238), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5239) );
  AND2_X1 U6642 ( .A1(n5248), .A2(n5239), .ZN(n9143) );
  AOI22_X1 U6643 ( .A1(n8906), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n5443), .B2(
        n9143), .ZN(n5243) );
  XNOR2_X1 U6644 ( .A(n5241), .B(n5240), .ZN(n6592) );
  NAND2_X1 U6645 ( .A1(n6592), .A2(n8910), .ZN(n5242) );
  NAND2_X1 U6646 ( .A1(n5243), .A2(n5242), .ZN(n6943) );
  INV_X1 U6647 ( .A(n6943), .ZN(n9738) );
  NAND2_X1 U6648 ( .A1(n9738), .A2(n9097), .ZN(n9028) );
  NAND2_X1 U6649 ( .A1(n6939), .A2(n6944), .ZN(n6940) );
  NAND2_X1 U6650 ( .A1(n5244), .A2(n9738), .ZN(n5245) );
  NAND2_X1 U6651 ( .A1(n6940), .A2(n5245), .ZN(n6927) );
  XNOR2_X1 U6652 ( .A(n5247), .B(n5246), .ZN(n6598) );
  OR2_X1 U6653 ( .A1(n6598), .A2(n4508), .ZN(n5251) );
  NAND2_X1 U6654 ( .A1(n5248), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5249) );
  XNOR2_X1 U6655 ( .A(n5249), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9156) );
  AOI22_X1 U6656 ( .A1(n8906), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5443), .B2(
        n9156), .ZN(n5250) );
  NAND2_X1 U6657 ( .A1(n5251), .A2(n5250), .ZN(n6925) );
  NAND2_X1 U6658 ( .A1(n6554), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5257) );
  NAND2_X1 U6659 ( .A1(n5201), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5256) );
  OAI21_X1 U6660 ( .B1(n5252), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5267), .ZN(
        n7263) );
  INV_X1 U6661 ( .A(n7263), .ZN(n7048) );
  NAND2_X1 U6662 ( .A1(n5202), .A2(n7048), .ZN(n5255) );
  NAND2_X1 U6663 ( .A1(n5200), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6664 ( .A1(n7264), .A2(n9096), .ZN(n9022) );
  INV_X1 U6665 ( .A(n9096), .ZN(n5258) );
  NAND2_X1 U6666 ( .A1(n5258), .A2(n6925), .ZN(n8795) );
  AND2_X1 U6667 ( .A1(n9022), .A2(n8795), .ZN(n8931) );
  NAND2_X1 U6668 ( .A1(n7264), .A2(n5258), .ZN(n5259) );
  NAND2_X1 U6669 ( .A1(n6929), .A2(n5259), .ZN(n6964) );
  XNOR2_X1 U6670 ( .A(n5261), .B(n5260), .ZN(n6599) );
  NAND2_X1 U6671 ( .A1(n6599), .A2(n8910), .ZN(n5265) );
  NAND2_X1 U6672 ( .A1(n5262), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5263) );
  XNOR2_X1 U6673 ( .A(n5263), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9169) );
  AOI22_X1 U6674 ( .A1(n8906), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5443), .B2(
        n9169), .ZN(n5264) );
  NAND2_X1 U6675 ( .A1(n5265), .A2(n5264), .ZN(n6965) );
  NAND2_X1 U6676 ( .A1(n6554), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U6677 ( .A1(n5201), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5271) );
  AND2_X1 U6678 ( .A1(n5267), .A2(n5266), .ZN(n5268) );
  NOR2_X1 U6679 ( .A1(n5280), .A2(n5268), .ZN(n7252) );
  NAND2_X1 U6680 ( .A1(n5202), .A2(n7252), .ZN(n5270) );
  NAND2_X1 U6681 ( .A1(n5200), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5269) );
  NAND4_X1 U6682 ( .A1(n5272), .A2(n5271), .A3(n5270), .A4(n5269), .ZN(n9095)
         );
  INV_X1 U6683 ( .A(n9095), .ZN(n5273) );
  AND2_X1 U6684 ( .A1(n6965), .A2(n5273), .ZN(n8796) );
  INV_X1 U6685 ( .A(n8796), .ZN(n8802) );
  OR2_X1 U6686 ( .A1(n6965), .A2(n5273), .ZN(n7186) );
  NAND2_X1 U6687 ( .A1(n8802), .A2(n7186), .ZN(n6963) );
  NAND2_X1 U6688 ( .A1(n6964), .A2(n6963), .ZN(n6962) );
  OR2_X1 U6689 ( .A1(n6965), .A2(n9095), .ZN(n5274) );
  NAND2_X1 U6690 ( .A1(n6962), .A2(n5274), .ZN(n7183) );
  XNOR2_X1 U6691 ( .A(n5276), .B(n5275), .ZN(n6614) );
  NAND2_X1 U6692 ( .A1(n6614), .A2(n8910), .ZN(n5279) );
  NAND2_X1 U6693 ( .A1(n5146), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5277) );
  XNOR2_X1 U6694 ( .A(n5277), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6696) );
  AOI22_X1 U6695 ( .A1(n8906), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5443), .B2(
        n6696), .ZN(n5278) );
  NAND2_X1 U6696 ( .A1(n6554), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6697 ( .A1(n5201), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5285) );
  OR2_X1 U6698 ( .A1(n5280), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5281) );
  AND2_X1 U6699 ( .A1(n5282), .A2(n5281), .ZN(n7198) );
  NAND2_X1 U6700 ( .A1(n5202), .A2(n7198), .ZN(n5284) );
  NAND2_X1 U6701 ( .A1(n5200), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5283) );
  NAND4_X1 U6702 ( .A1(n5286), .A2(n5285), .A3(n5284), .A4(n5283), .ZN(n9094)
         );
  XNOR2_X1 U6703 ( .A(n7199), .B(n9094), .ZN(n8806) );
  INV_X1 U6704 ( .A(n8806), .ZN(n7182) );
  INV_X1 U6705 ( .A(n7199), .ZN(n9772) );
  INV_X1 U6706 ( .A(n9094), .ZN(n6332) );
  OR2_X1 U6707 ( .A1(n7375), .A2(n5288), .ZN(n8811) );
  NAND2_X1 U6708 ( .A1(n7375), .A2(n5288), .ZN(n8812) );
  NAND2_X1 U6709 ( .A1(n6636), .A2(n8910), .ZN(n5295) );
  INV_X1 U6710 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U6711 ( .A1(n5291), .A2(n5290), .ZN(n5292) );
  NAND2_X1 U6712 ( .A1(n5292), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5293) );
  XNOR2_X1 U6713 ( .A(n5293), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6719) );
  AOI22_X1 U6714 ( .A1(n8906), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5443), .B2(
        n6719), .ZN(n5294) );
  NAND2_X2 U6715 ( .A1(n5295), .A2(n5294), .ZN(n7359) );
  NAND2_X1 U6716 ( .A1(n5201), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5301) );
  NAND2_X1 U6717 ( .A1(n6554), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5300) );
  AND2_X1 U6718 ( .A1(n5296), .A2(n6684), .ZN(n5297) );
  NOR2_X1 U6719 ( .A1(n5309), .A2(n5297), .ZN(n7441) );
  NAND2_X1 U6720 ( .A1(n5202), .A2(n7441), .ZN(n5299) );
  NAND2_X1 U6721 ( .A1(n5200), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5298) );
  NAND4_X1 U6722 ( .A1(n5301), .A2(n5300), .A3(n5299), .A4(n5298), .ZN(n9092)
         );
  NAND2_X1 U6723 ( .A1(n7359), .A2(n6342), .ZN(n8833) );
  NOR2_X1 U6724 ( .A1(n7348), .A2(n7347), .ZN(n7346) );
  NAND2_X1 U6725 ( .A1(n6640), .A2(n8910), .ZN(n5308) );
  OR2_X1 U6726 ( .A1(n5305), .A2(n5322), .ZN(n5306) );
  XNOR2_X1 U6727 ( .A(n5306), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6723) );
  AOI22_X1 U6728 ( .A1(n8906), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5443), .B2(
        n6723), .ZN(n5307) );
  NAND2_X1 U6729 ( .A1(n5201), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5315) );
  NOR2_X1 U6730 ( .A1(n5309), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5310) );
  OR2_X1 U6731 ( .A1(n5327), .A2(n5310), .ZN(n7467) );
  INV_X1 U6732 ( .A(n7467), .ZN(n5311) );
  NAND2_X1 U6733 ( .A1(n5202), .A2(n5311), .ZN(n5314) );
  NAND2_X1 U6734 ( .A1(n5200), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U6735 ( .A1(n6554), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5312) );
  NAND4_X1 U6736 ( .A1(n5315), .A2(n5314), .A3(n5313), .A4(n5312), .ZN(n9091)
         );
  NAND2_X1 U6737 ( .A1(n7524), .A2(n5316), .ZN(n9713) );
  NOR2_X1 U6738 ( .A1(n7418), .A2(n8937), .ZN(n7417) );
  NOR2_X1 U6739 ( .A1(n5320), .A2(n5322), .ZN(n5321) );
  MUX2_X1 U6740 ( .A(n5322), .B(n5321), .S(P1_IR_REG_11__SCAN_IN), .Z(n5323)
         );
  INV_X1 U6741 ( .A(n5323), .ZN(n5324) );
  AOI22_X1 U6742 ( .A1(n8906), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5443), .B2(
        n9607), .ZN(n5325) );
  NAND2_X1 U6743 ( .A1(n5201), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U6744 ( .A1(n6554), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5332) );
  OR2_X1 U6745 ( .A1(n5327), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5328) );
  AND2_X1 U6746 ( .A1(n5329), .A2(n5328), .ZN(n9720) );
  NAND2_X1 U6747 ( .A1(n5202), .A2(n9720), .ZN(n5331) );
  NAND2_X1 U6748 ( .A1(n5200), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5330) );
  NAND4_X1 U6749 ( .A1(n5333), .A2(n5332), .A3(n5331), .A4(n5330), .ZN(n9090)
         );
  MUX2_X1 U6750 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6584), .Z(n5354) );
  XNOR2_X1 U6751 ( .A(n5354), .B(SI_13_), .ZN(n5351) );
  XNOR2_X1 U6752 ( .A(n5353), .B(n5351), .ZN(n6800) );
  NAND2_X1 U6753 ( .A1(n6800), .A2(n8910), .ZN(n5342) );
  OAI21_X1 U6754 ( .B1(n5339), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5340) );
  XNOR2_X1 U6755 ( .A(n5340), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9633) );
  AOI22_X1 U6756 ( .A1(n8906), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5443), .B2(
        n9633), .ZN(n5341) );
  NAND2_X1 U6757 ( .A1(n6554), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U6758 ( .A1(n5201), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5348) );
  INV_X1 U6759 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U6760 ( .A1(n5344), .A2(n5343), .ZN(n5345) );
  AND2_X1 U6761 ( .A1(n5361), .A2(n5345), .ZN(n7660) );
  NAND2_X1 U6762 ( .A1(n5202), .A2(n7660), .ZN(n5347) );
  NAND2_X1 U6763 ( .A1(n5200), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5346) );
  NAND4_X1 U6764 ( .A1(n5349), .A2(n5348), .A3(n5347), .A4(n5346), .ZN(n9088)
         );
  NOR2_X1 U6765 ( .A1(n8849), .A2(n8846), .ZN(n5350) );
  OAI22_X1 U6766 ( .A1(n7654), .A2(n5350), .B1(n9088), .B2(n8845), .ZN(n7732)
         );
  INV_X1 U6767 ( .A(n5351), .ZN(n5352) );
  NAND2_X1 U6768 ( .A1(n5354), .A2(SI_13_), .ZN(n5355) );
  MUX2_X1 U6769 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6584), .Z(n5371) );
  XNOR2_X1 U6770 ( .A(n5371), .B(SI_14_), .ZN(n5368) );
  XNOR2_X1 U6771 ( .A(n5370), .B(n5368), .ZN(n6822) );
  NAND2_X1 U6772 ( .A1(n6822), .A2(n8910), .ZN(n5360) );
  NAND2_X1 U6773 ( .A1(n5356), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5357) );
  MUX2_X1 U6774 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5357), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n5358) );
  AND2_X1 U6775 ( .A1(n5391), .A2(n5358), .ZN(n9645) );
  AOI22_X1 U6776 ( .A1(n8906), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5443), .B2(
        n9645), .ZN(n5359) );
  INV_X1 U6777 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7672) );
  AND2_X1 U6778 ( .A1(n5361), .A2(n7672), .ZN(n5362) );
  NOR2_X1 U6779 ( .A1(n5378), .A2(n5362), .ZN(n7741) );
  NAND2_X1 U6780 ( .A1(n7741), .A2(n5202), .ZN(n5366) );
  NAND2_X1 U6781 ( .A1(n5201), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5365) );
  NAND2_X1 U6782 ( .A1(n5200), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U6783 ( .A1(n6554), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5363) );
  NAND4_X1 U6784 ( .A1(n5366), .A2(n5365), .A3(n5364), .A4(n5363), .ZN(n9087)
         );
  NOR2_X1 U6785 ( .A1(n8824), .A2(n9087), .ZN(n5367) );
  INV_X1 U6786 ( .A(n9087), .ZN(n8821) );
  INV_X1 U6787 ( .A(n5368), .ZN(n5369) );
  NAND2_X1 U6788 ( .A1(n5371), .A2(SI_14_), .ZN(n5372) );
  MUX2_X1 U6789 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6584), .Z(n5383) );
  XNOR2_X1 U6790 ( .A(n5383), .B(SI_15_), .ZN(n5374) );
  XNOR2_X1 U6791 ( .A(n5388), .B(n5374), .ZN(n6936) );
  NAND2_X1 U6792 ( .A1(n6936), .A2(n8910), .ZN(n5377) );
  NAND2_X1 U6793 ( .A1(n5391), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5375) );
  INV_X1 U6794 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5392) );
  XNOR2_X1 U6795 ( .A(n5375), .B(n5392), .ZN(n9218) );
  INV_X1 U6796 ( .A(n9218), .ZN(n9658) );
  AOI22_X1 U6797 ( .A1(n8906), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5443), .B2(
        n9658), .ZN(n5376) );
  INV_X1 U6798 ( .A(n8860), .ZN(n7718) );
  NAND2_X1 U6799 ( .A1(n5378), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5396) );
  OR2_X1 U6800 ( .A1(n5378), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6801 ( .A1(n5396), .A2(n5379), .ZN(n7707) );
  INV_X1 U6802 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n7717) );
  OAI22_X1 U6803 ( .A1(n7707), .A2(n5521), .B1(n5253), .B2(n7717), .ZN(n5381)
         );
  INV_X1 U6804 ( .A(n5201), .ZN(n5524) );
  INV_X1 U6805 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9651) );
  INV_X1 U6806 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9654) );
  OAI22_X1 U6807 ( .A1(n5524), .A2(n9651), .B1(n5180), .B2(n9654), .ZN(n5380)
         );
  INV_X1 U6808 ( .A(n9086), .ZN(n7749) );
  NOR2_X1 U6809 ( .A1(n7718), .A2(n7749), .ZN(n5382) );
  INV_X1 U6810 ( .A(SI_15_), .ZN(n5384) );
  NOR2_X1 U6811 ( .A1(n5385), .A2(n5384), .ZN(n5387) );
  NAND2_X1 U6812 ( .A1(n5385), .A2(n5384), .ZN(n5386) );
  INV_X1 U6813 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10341) );
  INV_X1 U6814 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5389) );
  MUX2_X1 U6815 ( .A(n10341), .B(n5389), .S(n6584), .Z(n5400) );
  XNOR2_X1 U6816 ( .A(n5400), .B(SI_16_), .ZN(n5390) );
  XNOR2_X1 U6817 ( .A(n5404), .B(n5390), .ZN(n6956) );
  NAND2_X1 U6818 ( .A1(n6956), .A2(n8910), .ZN(n5394) );
  XNOR2_X1 U6819 ( .A(n5408), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9674) );
  AOI22_X1 U6820 ( .A1(n8906), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5443), .B2(
        n9674), .ZN(n5393) );
  INV_X1 U6821 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U6822 ( .A1(n5396), .A2(n5395), .ZN(n5397) );
  NAND2_X1 U6823 ( .A1(n5413), .A2(n5397), .ZN(n8710) );
  AOI22_X1 U6824 ( .A1(n5201), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n6554), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n5399) );
  NAND2_X1 U6825 ( .A1(n5200), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5398) );
  OAI211_X1 U6826 ( .C1(n8710), .C2(n5521), .A(n5399), .B(n5398), .ZN(n9085)
         );
  INV_X1 U6827 ( .A(n9085), .ZN(n7698) );
  NAND2_X1 U6828 ( .A1(n9500), .A2(n7698), .ZN(n9015) );
  NOR2_X1 U6829 ( .A1(n5401), .A2(SI_16_), .ZN(n5403) );
  NAND2_X1 U6830 ( .A1(n5401), .A2(SI_16_), .ZN(n5402) );
  INV_X1 U6831 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7084) );
  INV_X1 U6832 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7083) );
  MUX2_X1 U6833 ( .A(n7084), .B(n7083), .S(n6584), .Z(n5405) );
  INV_X1 U6834 ( .A(SI_17_), .ZN(n10454) );
  NAND2_X1 U6835 ( .A1(n5405), .A2(n10454), .ZN(n5418) );
  INV_X1 U6836 ( .A(n5405), .ZN(n5406) );
  NAND2_X1 U6837 ( .A1(n5406), .A2(SI_17_), .ZN(n5407) );
  NAND2_X1 U6838 ( .A1(n5418), .A2(n5407), .ZN(n5419) );
  XNOR2_X1 U6839 ( .A(n5420), .B(n5419), .ZN(n7082) );
  NAND2_X1 U6840 ( .A1(n7082), .A2(n8910), .ZN(n5411) );
  INV_X1 U6841 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U6842 ( .A1(n5408), .A2(n5625), .ZN(n5409) );
  XNOR2_X1 U6843 ( .A(n5421), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9224) );
  AOI22_X1 U6844 ( .A1(n8906), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5443), .B2(
        n9224), .ZN(n5410) );
  INV_X1 U6845 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5412) );
  AND2_X1 U6846 ( .A1(n5413), .A2(n5412), .ZN(n5414) );
  OR2_X1 U6847 ( .A1(n5414), .A2(n5427), .ZN(n8723) );
  AOI22_X1 U6848 ( .A1(n5201), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n6554), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U6849 ( .A1(n5200), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5415) );
  OAI211_X1 U6850 ( .C1(n8723), .C2(n5521), .A(n5416), .B(n5415), .ZN(n9084)
         );
  INV_X1 U6851 ( .A(n9084), .ZN(n7751) );
  NAND2_X1 U6852 ( .A1(n9427), .A2(n7751), .ZN(n5417) );
  INV_X1 U6853 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7204) );
  INV_X1 U6854 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7146) );
  MUX2_X1 U6855 ( .A(n7204), .B(n7146), .S(n6584), .Z(n5434) );
  XNOR2_X1 U6856 ( .A(n5434), .B(SI_18_), .ZN(n5433) );
  XNOR2_X1 U6857 ( .A(n5436), .B(n5433), .ZN(n7145) );
  NAND2_X1 U6858 ( .A1(n7145), .A2(n8910), .ZN(n5426) );
  INV_X1 U6859 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U6860 ( .A1(n5421), .A2(n5626), .ZN(n5422) );
  INV_X1 U6861 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U6862 ( .A1(n5423), .A2(n5627), .ZN(n5441) );
  OR2_X1 U6863 ( .A1(n5423), .A2(n5627), .ZN(n5424) );
  AND2_X1 U6864 ( .A1(n5441), .A2(n5424), .ZN(n9227) );
  AOI22_X1 U6865 ( .A1(n8906), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5443), .B2(
        n9227), .ZN(n5425) );
  NOR2_X1 U6866 ( .A1(n5427), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5428) );
  OR2_X1 U6867 ( .A1(n5446), .A2(n5428), .ZN(n9406) );
  AOI22_X1 U6868 ( .A1(n5201), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n5200), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U6869 ( .A1(n6554), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5429) );
  OAI211_X1 U6870 ( .C1(n9406), .C2(n5521), .A(n5430), .B(n5429), .ZN(n9083)
         );
  NAND2_X1 U6871 ( .A1(n9487), .A2(n9083), .ZN(n5432) );
  NOR2_X1 U6872 ( .A1(n9487), .A2(n9083), .ZN(n5431) );
  INV_X1 U6873 ( .A(n5434), .ZN(n5435) );
  INV_X1 U6874 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7307) );
  INV_X1 U6875 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8007) );
  MUX2_X1 U6876 ( .A(n7307), .B(n8007), .S(n6584), .Z(n5438) );
  INV_X1 U6877 ( .A(SI_19_), .ZN(n5437) );
  NAND2_X1 U6878 ( .A1(n5438), .A2(n5437), .ZN(n5459) );
  INV_X1 U6879 ( .A(n5438), .ZN(n5439) );
  NAND2_X1 U6880 ( .A1(n5439), .A2(SI_19_), .ZN(n5440) );
  NAND2_X1 U6881 ( .A1(n5459), .A2(n5440), .ZN(n5457) );
  XNOR2_X1 U6882 ( .A(n5456), .B(n5457), .ZN(n7306) );
  NAND2_X1 U6883 ( .A1(n7306), .A2(n8910), .ZN(n5445) );
  INV_X1 U6884 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5624) );
  INV_X1 U6885 ( .A(n4507), .ZN(n6252) );
  AOI22_X1 U6886 ( .A1(n6252), .A2(n5443), .B1(n8906), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n5444) );
  INV_X1 U6887 ( .A(n9481), .ZN(n9395) );
  OR2_X1 U6888 ( .A1(n5446), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5447) );
  AND2_X1 U6889 ( .A1(n5480), .A2(n5447), .ZN(n9392) );
  NAND2_X1 U6890 ( .A1(n9392), .A2(n5202), .ZN(n5452) );
  INV_X1 U6891 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10372) );
  NAND2_X1 U6892 ( .A1(n5201), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U6893 ( .A1(n6554), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5448) );
  OAI211_X1 U6894 ( .C1(n5253), .C2(n10372), .A(n5449), .B(n5448), .ZN(n5450)
         );
  INV_X1 U6895 ( .A(n5450), .ZN(n5451) );
  NAND2_X1 U6896 ( .A1(n5452), .A2(n5451), .ZN(n9082) );
  INV_X1 U6897 ( .A(n9082), .ZN(n8787) );
  NAND2_X1 U6898 ( .A1(n9395), .A2(n8787), .ZN(n5453) );
  NAND2_X1 U6899 ( .A1(n9386), .A2(n5453), .ZN(n5455) );
  NAND2_X1 U6900 ( .A1(n9481), .A2(n9082), .ZN(n5454) );
  INV_X1 U6901 ( .A(n5457), .ZN(n5458) );
  MUX2_X1 U6902 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n5082), .Z(n5471) );
  INV_X1 U6903 ( .A(SI_20_), .ZN(n5473) );
  XNOR2_X1 U6904 ( .A(n5471), .B(n5473), .ZN(n5460) );
  XNOR2_X1 U6905 ( .A(n5474), .B(n5460), .ZN(n7414) );
  NAND2_X1 U6906 ( .A1(n7414), .A2(n8910), .ZN(n5462) );
  NAND2_X1 U6907 ( .A1(n8906), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5461) );
  XNOR2_X1 U6908 ( .A(n5480), .B(P1_REG3_REG_20__SCAN_IN), .ZN(n9381) );
  NAND2_X1 U6909 ( .A1(n9381), .A2(n5202), .ZN(n5468) );
  INV_X1 U6910 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U6911 ( .A1(n5200), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U6912 ( .A1(n5201), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5463) );
  OAI211_X1 U6913 ( .C1(n5180), .C2(n5465), .A(n5464), .B(n5463), .ZN(n5466)
         );
  INV_X1 U6914 ( .A(n5466), .ZN(n5467) );
  NAND2_X1 U6915 ( .A1(n5468), .A2(n5467), .ZN(n9081) );
  INV_X1 U6916 ( .A(n9081), .ZN(n5661) );
  NOR2_X1 U6917 ( .A1(n4773), .A2(n5661), .ZN(n5469) );
  NAND2_X1 U6918 ( .A1(n4773), .A2(n5661), .ZN(n5470) );
  INV_X1 U6919 ( .A(n5471), .ZN(n5472) );
  INV_X1 U6920 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10376) );
  INV_X1 U6921 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7475) );
  MUX2_X1 U6922 ( .A(n10376), .B(n7475), .S(n6584), .Z(n5488) );
  XNOR2_X1 U6923 ( .A(n5488), .B(SI_21_), .ZN(n5476) );
  XNOR2_X1 U6924 ( .A(n5492), .B(n5476), .ZN(n7474) );
  NAND2_X1 U6925 ( .A1(n7474), .A2(n8910), .ZN(n5478) );
  NAND2_X1 U6926 ( .A1(n8906), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5477) );
  INV_X1 U6927 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8740) );
  INV_X1 U6928 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8697) );
  OAI21_X1 U6929 ( .B1(n5480), .B2(n8740), .A(n8697), .ZN(n5481) );
  NAND2_X1 U6930 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .ZN(n5479) );
  NAND2_X1 U6931 ( .A1(n5481), .A2(n5499), .ZN(n9365) );
  OR2_X1 U6932 ( .A1(n9365), .A2(n5521), .ZN(n5486) );
  INV_X1 U6933 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10447) );
  NAND2_X1 U6934 ( .A1(n6554), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U6935 ( .A1(n5200), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5482) );
  OAI211_X1 U6936 ( .C1(n5524), .C2(n10447), .A(n5483), .B(n5482), .ZN(n5484)
         );
  INV_X1 U6937 ( .A(n5484), .ZN(n5485) );
  NAND2_X1 U6938 ( .A1(n5486), .A2(n5485), .ZN(n9080) );
  INV_X1 U6939 ( .A(n9080), .ZN(n8873) );
  NAND2_X1 U6940 ( .A1(n9544), .A2(n8873), .ZN(n5487) );
  INV_X1 U6941 ( .A(n5488), .ZN(n5489) );
  NOR2_X1 U6942 ( .A1(n5489), .A2(SI_21_), .ZN(n5491) );
  NAND2_X1 U6943 ( .A1(n5489), .A2(SI_21_), .ZN(n5490) );
  INV_X1 U6944 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7549) );
  INV_X1 U6945 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7548) );
  MUX2_X1 U6946 ( .A(n7549), .B(n7548), .S(n6584), .Z(n5494) );
  INV_X1 U6947 ( .A(SI_22_), .ZN(n5493) );
  NAND2_X1 U6948 ( .A1(n5494), .A2(n5493), .ZN(n5510) );
  INV_X1 U6949 ( .A(n5494), .ZN(n5495) );
  NAND2_X1 U6950 ( .A1(n5495), .A2(SI_22_), .ZN(n5496) );
  NAND2_X1 U6951 ( .A1(n5510), .A2(n5496), .ZN(n5508) );
  XNOR2_X1 U6952 ( .A(n5509), .B(n5508), .ZN(n7547) );
  NAND2_X1 U6953 ( .A1(n7547), .A2(n8910), .ZN(n5498) );
  NAND2_X1 U6954 ( .A1(n8906), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5497) );
  INV_X1 U6955 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8752) );
  AND2_X1 U6956 ( .A1(n5499), .A2(n8752), .ZN(n5500) );
  OR2_X1 U6957 ( .A1(n5500), .A2(n5519), .ZN(n9349) );
  INV_X1 U6958 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10394) );
  NAND2_X1 U6959 ( .A1(n5200), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5502) );
  NAND2_X1 U6960 ( .A1(n6554), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5501) );
  OAI211_X1 U6961 ( .C1(n5524), .C2(n10394), .A(n5502), .B(n5501), .ZN(n5503)
         );
  INV_X1 U6962 ( .A(n5503), .ZN(n5504) );
  OAI21_X1 U6963 ( .B1(n9349), .B2(n5521), .A(n5504), .ZN(n9079) );
  INV_X1 U6964 ( .A(n9079), .ZN(n8886) );
  NOR2_X1 U6965 ( .A1(n9353), .A2(n8886), .ZN(n5505) );
  OR2_X1 U6966 ( .A1(n9341), .A2(n5505), .ZN(n5507) );
  NAND2_X1 U6967 ( .A1(n9353), .A2(n8886), .ZN(n5506) );
  INV_X1 U6968 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5512) );
  INV_X1 U6969 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5511) );
  MUX2_X1 U6970 ( .A(n5512), .B(n5511), .S(n6584), .Z(n5514) );
  INV_X1 U6971 ( .A(SI_23_), .ZN(n5513) );
  NAND2_X1 U6972 ( .A1(n5514), .A2(n5513), .ZN(n5547) );
  INV_X1 U6973 ( .A(n5514), .ZN(n5515) );
  NAND2_X1 U6974 ( .A1(n5515), .A2(SI_23_), .ZN(n5516) );
  AND2_X1 U6975 ( .A1(n5547), .A2(n5516), .ZN(n5529) );
  NAND2_X1 U6976 ( .A1(n7611), .A2(n8910), .ZN(n5518) );
  NAND2_X1 U6977 ( .A1(n8906), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5517) );
  OR2_X1 U6978 ( .A1(n5519), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U6979 ( .A1(n5519), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U6980 ( .A1(n5520), .A2(n5538), .ZN(n9335) );
  OR2_X1 U6981 ( .A1(n9335), .A2(n5521), .ZN(n5527) );
  INV_X1 U6982 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10409) );
  NAND2_X1 U6983 ( .A1(n6554), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U6984 ( .A1(n5200), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5522) );
  OAI211_X1 U6985 ( .C1(n5524), .C2(n10409), .A(n5523), .B(n5522), .ZN(n5525)
         );
  INV_X1 U6986 ( .A(n5525), .ZN(n5526) );
  NAND2_X1 U6987 ( .A1(n5527), .A2(n5526), .ZN(n9078) );
  INV_X1 U6988 ( .A(n9078), .ZN(n5665) );
  NAND2_X1 U6989 ( .A1(n5571), .A2(n5547), .ZN(n5534) );
  INV_X1 U6990 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7651) );
  INV_X1 U6991 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7634) );
  MUX2_X1 U6992 ( .A(n7651), .B(n7634), .S(n6584), .Z(n5531) );
  NAND2_X1 U6993 ( .A1(n5531), .A2(n10267), .ZN(n5546) );
  INV_X1 U6994 ( .A(n5531), .ZN(n5532) );
  NAND2_X1 U6995 ( .A1(n5532), .A2(SI_24_), .ZN(n5566) );
  AND2_X1 U6996 ( .A1(n5546), .A2(n5566), .ZN(n5533) );
  NAND2_X1 U6997 ( .A1(n7633), .A2(n8910), .ZN(n5536) );
  NAND2_X1 U6998 ( .A1(n8906), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U6999 ( .A1(n6554), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U7000 ( .A1(n5201), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5542) );
  INV_X1 U7001 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5539) );
  INV_X1 U7002 ( .A(n5538), .ZN(n5537) );
  NAND2_X1 U7003 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n5537), .ZN(n5558) );
  AOI21_X1 U7004 ( .B1(n5539), .B2(n5538), .A(n5556), .ZN(n9322) );
  NAND2_X1 U7005 ( .A1(n5202), .A2(n9322), .ZN(n5541) );
  NAND2_X1 U7006 ( .A1(n5200), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5540) );
  NAND4_X1 U7007 ( .A1(n5543), .A2(n5542), .A3(n5541), .A4(n5540), .ZN(n9077)
         );
  INV_X1 U7008 ( .A(n9077), .ZN(n5640) );
  NOR2_X1 U7009 ( .A1(n9454), .A2(n5640), .ZN(n5545) );
  NAND2_X1 U7010 ( .A1(n9454), .A2(n5640), .ZN(n5544) );
  AND2_X1 U7011 ( .A1(n5547), .A2(n5546), .ZN(n5564) );
  NAND2_X1 U7012 ( .A1(n5571), .A2(n5564), .ZN(n5548) );
  INV_X1 U7013 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7688) );
  INV_X1 U7014 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7667) );
  MUX2_X1 U7015 ( .A(n7688), .B(n7667), .S(n6584), .Z(n5550) );
  INV_X1 U7016 ( .A(SI_25_), .ZN(n5549) );
  NAND2_X1 U7017 ( .A1(n5550), .A2(n5549), .ZN(n5565) );
  INV_X1 U7018 ( .A(n5550), .ZN(n5551) );
  NAND2_X1 U7019 ( .A1(n5551), .A2(SI_25_), .ZN(n5552) );
  AND2_X1 U7020 ( .A1(n5565), .A2(n5552), .ZN(n5567) );
  NAND2_X1 U7021 ( .A1(n8906), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U7022 ( .A1(n5201), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U7023 ( .A1(n5200), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5561) );
  INV_X1 U7024 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8702) );
  INV_X1 U7025 ( .A(n5578), .ZN(n5557) );
  AOI21_X1 U7026 ( .B1(n8702), .B2(n5558), .A(n5557), .ZN(n9298) );
  NAND2_X1 U7027 ( .A1(n5202), .A2(n9298), .ZN(n5560) );
  NAND2_X1 U7028 ( .A1(n6554), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5559) );
  NAND4_X1 U7029 ( .A1(n5562), .A2(n5561), .A3(n5560), .A4(n5559), .ZN(n9076)
         );
  INV_X1 U7030 ( .A(n9076), .ZN(n5638) );
  AND2_X1 U7031 ( .A1(n5564), .A2(n5565), .ZN(n5570) );
  INV_X1 U7032 ( .A(n5565), .ZN(n5569) );
  AND2_X1 U7033 ( .A1(n5567), .A2(n5566), .ZN(n5568) );
  INV_X1 U7034 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n10246) );
  INV_X1 U7035 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7678) );
  MUX2_X1 U7036 ( .A(n10246), .B(n7678), .S(n6584), .Z(n5573) );
  INV_X1 U7037 ( .A(SI_26_), .ZN(n5572) );
  NAND2_X1 U7038 ( .A1(n5573), .A2(n5572), .ZN(n5587) );
  INV_X1 U7039 ( .A(n5573), .ZN(n5574) );
  NAND2_X1 U7040 ( .A1(n5574), .A2(SI_26_), .ZN(n5575) );
  AND2_X1 U7041 ( .A1(n5587), .A2(n5575), .ZN(n5585) );
  NAND2_X1 U7042 ( .A1(n8906), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5576) );
  INV_X1 U7043 ( .A(n9446), .ZN(n8786) );
  NAND2_X1 U7044 ( .A1(n6554), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U7045 ( .A1(n5201), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5581) );
  INV_X1 U7046 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n10439) );
  AOI21_X1 U7047 ( .B1(n10439), .B2(n5578), .A(n5614), .ZN(n9291) );
  NAND2_X1 U7048 ( .A1(n5202), .A2(n9291), .ZN(n5580) );
  NAND2_X1 U7049 ( .A1(n5200), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5579) );
  NAND4_X1 U7050 ( .A1(n5582), .A2(n5581), .A3(n5580), .A4(n5579), .ZN(n9075)
         );
  INV_X1 U7051 ( .A(n9075), .ZN(n8895) );
  NOR2_X1 U7052 ( .A1(n8786), .A2(n8895), .ZN(n5584) );
  OAI21_X1 U7053 ( .B1(n9285), .B2(n5584), .A(n5583), .ZN(n9268) );
  NAND2_X1 U7054 ( .A1(n5586), .A2(n5585), .ZN(n5588) );
  INV_X1 U7055 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n10424) );
  INV_X1 U7056 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5589) );
  MUX2_X1 U7057 ( .A(n10424), .B(n5589), .S(n6584), .Z(n5591) );
  INV_X1 U7058 ( .A(SI_27_), .ZN(n5590) );
  NAND2_X1 U7059 ( .A1(n5591), .A2(n5590), .ZN(n5605) );
  INV_X1 U7060 ( .A(n5591), .ZN(n5592) );
  NAND2_X1 U7061 ( .A1(n5592), .A2(SI_27_), .ZN(n5593) );
  AND2_X1 U7062 ( .A1(n5605), .A2(n5593), .ZN(n5594) );
  NAND2_X1 U7063 ( .A1(n8906), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U7064 ( .A1(n5201), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U7065 ( .A1(n5200), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5602) );
  INV_X1 U7066 ( .A(n5614), .ZN(n5599) );
  XNOR2_X1 U7067 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n5599), .ZN(n9272) );
  NAND2_X1 U7068 ( .A1(n5202), .A2(n9272), .ZN(n5601) );
  NAND2_X1 U7069 ( .A1(n6554), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5600) );
  NAND4_X1 U7070 ( .A1(n5603), .A2(n5602), .A3(n5601), .A4(n5600), .ZN(n9074)
         );
  INV_X1 U7071 ( .A(n8984), .ZN(n8899) );
  NAND2_X1 U7072 ( .A1(n9269), .A2(n6500), .ZN(n6552) );
  NAND2_X1 U7073 ( .A1(n9519), .A2(n6500), .ZN(n5604) );
  INV_X1 U7074 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5607) );
  INV_X1 U7075 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9570) );
  MUX2_X1 U7076 ( .A(n5607), .B(n9570), .S(n6584), .Z(n5609) );
  INV_X1 U7077 ( .A(SI_28_), .ZN(n5608) );
  NAND2_X1 U7078 ( .A1(n5609), .A2(n5608), .ZN(n6106) );
  INV_X1 U7079 ( .A(n5609), .ZN(n5610) );
  NAND2_X1 U7080 ( .A1(n5610), .A2(SI_28_), .ZN(n5611) );
  AND2_X1 U7081 ( .A1(n6106), .A2(n5611), .ZN(n6104) );
  NAND2_X1 U7082 ( .A1(n8671), .A2(n8910), .ZN(n5613) );
  NAND2_X1 U7083 ( .A1(n8906), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U7084 ( .A1(n6554), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U7085 ( .A1(n5201), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5620) );
  AND2_X1 U7086 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n5614), .ZN(n5615) );
  NAND2_X1 U7087 ( .A1(n5615), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n5670) );
  INV_X1 U7088 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n10361) );
  INV_X1 U7089 ( .A(n5615), .ZN(n5616) );
  NAND2_X1 U7090 ( .A1(n10361), .A2(n5616), .ZN(n5617) );
  NAND2_X1 U7091 ( .A1(n5202), .A2(n9258), .ZN(n5619) );
  NAND2_X1 U7092 ( .A1(n5200), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5618) );
  NAND4_X1 U7093 ( .A1(n5621), .A2(n5620), .A3(n5619), .A4(n5618), .ZN(n9073)
         );
  INV_X1 U7094 ( .A(n9073), .ZN(n6543) );
  NAND2_X1 U7095 ( .A1(n6539), .A2(n6543), .ZN(n6553) );
  NAND2_X1 U7096 ( .A1(n5622), .A2(n5667), .ZN(n9256) );
  INV_X1 U7097 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5628) );
  NAND2_X1 U7098 ( .A1(n5629), .A2(n5628), .ZN(n5630) );
  INV_X1 U7099 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5681) );
  NAND2_X1 U7100 ( .A1(n5632), .A2(n5681), .ZN(n5631) );
  OR2_X1 U7101 ( .A1(n9001), .A2(n9756), .ZN(n7036) );
  INV_X1 U7102 ( .A(n7036), .ZN(n5636) );
  NAND2_X1 U7103 ( .A1(n5680), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5633) );
  XNOR2_X1 U7104 ( .A(n5633), .B(n5628), .ZN(n7416) );
  NAND2_X1 U7105 ( .A1(n4507), .A2(n7416), .ZN(n6253) );
  NAND2_X1 U7106 ( .A1(n6254), .A2(n5634), .ZN(n6258) );
  NAND2_X1 U7107 ( .A1(n6253), .A2(n6258), .ZN(n5635) );
  NAND2_X1 U7108 ( .A1(n5636), .A2(n5635), .ZN(n7737) );
  OR2_X1 U7109 ( .A1(n4507), .A2(n6254), .ZN(n8919) );
  INV_X1 U7110 ( .A(n7416), .ZN(n9064) );
  OR2_X1 U7111 ( .A1(n8919), .A2(n9064), .ZN(n7366) );
  NAND2_X1 U7112 ( .A1(n7737), .A2(n7366), .ZN(n9768) );
  NAND3_X1 U7113 ( .A1(n9257), .A2(n9256), .A3(n9768), .ZN(n5679) );
  INV_X1 U7114 ( .A(n9487), .ZN(n9404) );
  NAND2_X1 U7115 ( .A1(n6941), .A2(n7264), .ZN(n6961) );
  NAND2_X1 U7116 ( .A1(n7657), .A2(n8849), .ZN(n7658) );
  OR2_X1 U7117 ( .A1(n7658), .A2(n8824), .ZN(n7739) );
  NAND2_X1 U7118 ( .A1(n9404), .A2(n9421), .ZN(n9399) );
  OR2_X2 U7119 ( .A1(n9347), .A2(n9459), .ZN(n9334) );
  NOR2_X2 U7120 ( .A1(n9323), .A2(n9334), .ZN(n9321) );
  NAND2_X1 U7121 ( .A1(n9321), .A2(n9527), .ZN(n9297) );
  NOR2_X2 U7122 ( .A1(n4529), .A2(n9269), .ZN(n9270) );
  OR2_X1 U7123 ( .A1(n9260), .A2(n9270), .ZN(n5637) );
  INV_X1 U7124 ( .A(n9422), .ZN(n9724) );
  AOI22_X1 U7125 ( .A1(n9263), .A2(n9724), .B1(n9499), .B2(n6539), .ZN(n5677)
         );
  INV_X1 U7126 ( .A(n9300), .ZN(n5639) );
  NOR2_X1 U7127 ( .A1(n9301), .A2(n5639), .ZN(n5666) );
  NAND2_X1 U7128 ( .A1(n9323), .A2(n5640), .ZN(n8974) );
  XNOR2_X1 U7129 ( .A(n9467), .B(n8886), .ZN(n9342) );
  INV_X1 U7130 ( .A(n9342), .ZN(n5664) );
  NAND2_X1 U7131 ( .A1(n7199), .A2(n6332), .ZN(n7282) );
  NAND2_X1 U7132 ( .A1(n8812), .A2(n7282), .ZN(n8807) );
  AND2_X1 U7133 ( .A1(n8811), .A2(n8807), .ZN(n7341) );
  NAND2_X1 U7134 ( .A1(n7341), .A2(n8831), .ZN(n5641) );
  NAND2_X1 U7135 ( .A1(n5641), .A2(n8833), .ZN(n5650) );
  NOR2_X1 U7136 ( .A1(n5650), .A2(n8796), .ZN(n8938) );
  INV_X1 U7137 ( .A(n9755), .ZN(n7033) );
  NOR2_X1 U7138 ( .A1(n6265), .A2(n7033), .ZN(n7148) );
  NAND2_X1 U7139 ( .A1(n5643), .A2(n7153), .ZN(n5644) );
  NAND2_X1 U7140 ( .A1(n7147), .A2(n5644), .ZN(n7209) );
  NAND2_X1 U7141 ( .A1(n6285), .A2(n9766), .ZN(n9024) );
  NAND2_X1 U7142 ( .A1(n7209), .A2(n9024), .ZN(n5646) );
  NAND2_X1 U7143 ( .A1(n6752), .A2(n6772), .ZN(n5645) );
  NAND2_X1 U7144 ( .A1(n5646), .A2(n5645), .ZN(n8789) );
  OR2_X1 U7145 ( .A1(n8789), .A2(n5647), .ZN(n5648) );
  AND2_X1 U7146 ( .A1(n8790), .A2(n8795), .ZN(n8798) );
  NAND2_X1 U7147 ( .A1(n8793), .A2(n8798), .ZN(n7187) );
  NAND2_X1 U7148 ( .A1(n7187), .A2(n9022), .ZN(n6958) );
  NAND2_X1 U7149 ( .A1(n8938), .A2(n6958), .ZN(n9035) );
  OR2_X1 U7150 ( .A1(n7199), .A2(n6332), .ZN(n5649) );
  AND2_X1 U7151 ( .A1(n8811), .A2(n5649), .ZN(n8808) );
  AND3_X1 U7152 ( .A1(n8831), .A2(n8808), .A3(n7186), .ZN(n8926) );
  AND2_X1 U7153 ( .A1(n9032), .A2(n8937), .ZN(n5651) );
  INV_X1 U7154 ( .A(n9090), .ZN(n6368) );
  NAND2_X1 U7155 ( .A1(n9723), .A2(n6368), .ZN(n8835) );
  INV_X1 U7156 ( .A(n9713), .ZN(n5652) );
  NAND2_X1 U7157 ( .A1(n9714), .A2(n5653), .ZN(n9711) );
  NAND2_X1 U7158 ( .A1(n9711), .A2(n8836), .ZN(n7584) );
  OR2_X1 U7159 ( .A1(n7620), .A2(n6378), .ZN(n8837) );
  AND2_X1 U7160 ( .A1(n7620), .A2(n6378), .ZN(n9039) );
  INV_X1 U7161 ( .A(n9039), .ZN(n8842) );
  NAND2_X1 U7162 ( .A1(n8837), .A2(n8842), .ZN(n8940) );
  INV_X1 U7163 ( .A(n8940), .ZN(n7583) );
  NAND2_X1 U7164 ( .A1(n7584), .A2(n7583), .ZN(n7582) );
  XNOR2_X1 U7165 ( .A(n8845), .B(n9088), .ZN(n8941) );
  INV_X1 U7166 ( .A(n8941), .ZN(n5654) );
  AND2_X1 U7167 ( .A1(n8845), .A2(n8846), .ZN(n9040) );
  INV_X1 U7168 ( .A(n9040), .ZN(n8841) );
  NOR2_X1 U7169 ( .A1(n8824), .A2(n8821), .ZN(n9021) );
  INV_X1 U7170 ( .A(n9021), .ZN(n8817) );
  AND2_X1 U7171 ( .A1(n8824), .A2(n8821), .ZN(n9013) );
  INV_X1 U7172 ( .A(n9013), .ZN(n8843) );
  OR2_X1 U7173 ( .A1(n8860), .A2(n7749), .ZN(n9017) );
  NAND2_X1 U7174 ( .A1(n8860), .A2(n7749), .ZN(n8855) );
  NAND2_X1 U7175 ( .A1(n9017), .A2(n8855), .ZN(n8945) );
  INV_X1 U7176 ( .A(n8945), .ZN(n5656) );
  NAND2_X1 U7177 ( .A1(n5657), .A2(n9015), .ZN(n9415) );
  NOR2_X1 U7178 ( .A1(n9494), .A2(n7751), .ZN(n9019) );
  INV_X1 U7179 ( .A(n9019), .ZN(n8867) );
  NAND2_X1 U7180 ( .A1(n9494), .A2(n7751), .ZN(n8876) );
  INV_X1 U7181 ( .A(n9417), .ZN(n9414) );
  INV_X1 U7182 ( .A(n9083), .ZN(n5658) );
  OR2_X1 U7183 ( .A1(n9487), .A2(n5658), .ZN(n8874) );
  NAND2_X1 U7184 ( .A1(n9487), .A2(n5658), .ZN(n8877) );
  OR2_X1 U7185 ( .A1(n9481), .A2(n8787), .ZN(n8875) );
  NAND2_X1 U7186 ( .A1(n9481), .A2(n8787), .ZN(n9048) );
  NAND2_X1 U7187 ( .A1(n8875), .A2(n9048), .ZN(n9387) );
  INV_X1 U7188 ( .A(n9387), .ZN(n5660) );
  INV_X1 U7189 ( .A(n9048), .ZN(n5659) );
  OR2_X1 U7190 ( .A1(n9476), .A2(n5661), .ZN(n8883) );
  NAND2_X1 U7191 ( .A1(n9476), .A2(n5661), .ZN(n8975) );
  NAND2_X1 U7192 ( .A1(n8883), .A2(n8975), .ZN(n9375) );
  INV_X1 U7193 ( .A(n9375), .ZN(n5662) );
  NAND2_X1 U7194 ( .A1(n9376), .A2(n5662), .ZN(n5663) );
  NAND2_X1 U7195 ( .A1(n5663), .A2(n8883), .ZN(n9358) );
  XNOR2_X1 U7196 ( .A(n9367), .B(n8873), .ZN(n9357) );
  NAND2_X1 U7197 ( .A1(n9367), .A2(n8873), .ZN(n8976) );
  NAND2_X1 U7198 ( .A1(n9467), .A2(n8886), .ZN(n8889) );
  OR2_X1 U7199 ( .A1(n9459), .A2(n5665), .ZN(n8890) );
  NAND2_X1 U7200 ( .A1(n9459), .A2(n5665), .ZN(n9312) );
  NAND2_X1 U7201 ( .A1(n8890), .A2(n9312), .ZN(n8950) );
  NAND2_X1 U7202 ( .A1(n9330), .A2(n9331), .ZN(n9329) );
  NAND3_X1 U7203 ( .A1(n9311), .A2(n9329), .A3(n9312), .ZN(n9315) );
  AND2_X1 U7204 ( .A1(n9446), .A2(n8895), .ZN(n8993) );
  NAND2_X1 U7205 ( .A1(n9276), .A2(n6552), .ZN(n5668) );
  XNOR2_X1 U7206 ( .A(n5668), .B(n5667), .ZN(n5676) );
  OR2_X1 U7207 ( .A1(n6255), .A2(n4507), .ZN(n5669) );
  NAND2_X1 U7208 ( .A1(n6554), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U7209 ( .A1(n5201), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5673) );
  INV_X1 U7210 ( .A(n5670), .ZN(n7764) );
  NAND2_X1 U7211 ( .A1(n5202), .A2(n7764), .ZN(n5672) );
  NAND2_X1 U7212 ( .A1(n5200), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5671) );
  NAND4_X1 U7213 ( .A1(n5674), .A2(n5673), .A3(n5672), .A4(n5671), .ZN(n9072)
         );
  INV_X1 U7214 ( .A(n9072), .ZN(n6548) );
  AND2_X2 U7215 ( .A1(n9001), .A2(n5675), .ZN(n8777) );
  INV_X1 U7216 ( .A(n8777), .ZN(n7750) );
  INV_X1 U7217 ( .A(n5675), .ZN(n6682) );
  AND2_X2 U7218 ( .A1(n9001), .A2(n6682), .ZN(n9066) );
  INV_X1 U7219 ( .A(n9066), .ZN(n7748) );
  OAI22_X1 U7220 ( .A1(n6548), .A2(n7750), .B1(n6500), .B2(n7748), .ZN(n6532)
         );
  NAND2_X1 U7221 ( .A1(n5679), .A2(n5678), .ZN(n9438) );
  INV_X1 U7222 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U7223 ( .A1(n5683), .A2(n5682), .ZN(n5689) );
  OR2_X1 U7224 ( .A1(n5683), .A2(n5682), .ZN(n5684) );
  NAND2_X1 U7225 ( .A1(n5689), .A2(n5684), .ZN(n5711) );
  NAND2_X1 U7226 ( .A1(n5711), .A2(P1_B_REG_SCAN_IN), .ZN(n5688) );
  NAND2_X1 U7227 ( .A1(n5685), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5686) );
  XNOR2_X1 U7228 ( .A(n5686), .B(n10354), .ZN(n7635) );
  INV_X1 U7229 ( .A(n7635), .ZN(n5687) );
  MUX2_X1 U7230 ( .A(n5688), .B(P1_B_REG_SCAN_IN), .S(n5687), .Z(n5691) );
  INV_X1 U7231 ( .A(n6515), .ZN(n6632) );
  NOR4_X1 U7232 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5695) );
  NOR4_X1 U7233 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n5694) );
  NOR4_X1 U7234 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5693) );
  NOR4_X1 U7235 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5692) );
  NAND4_X1 U7236 ( .A1(n5695), .A2(n5694), .A3(n5693), .A4(n5692), .ZN(n5701)
         );
  NOR2_X1 U7237 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .ZN(
        n5699) );
  NOR4_X1 U7238 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5698) );
  NOR4_X1 U7239 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5697) );
  NOR4_X1 U7240 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5696) );
  NAND4_X1 U7241 ( .A1(n5699), .A2(n5698), .A3(n5697), .A4(n5696), .ZN(n5700)
         );
  NOR2_X1 U7242 ( .A1(n5701), .A2(n5700), .ZN(n6513) );
  INV_X1 U7243 ( .A(n6525), .ZN(n5705) );
  INV_X1 U7244 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6635) );
  NAND2_X1 U7245 ( .A1(n6515), .A2(n6635), .ZN(n5703) );
  INV_X1 U7246 ( .A(n5711), .ZN(n5702) );
  OR2_X1 U7247 ( .A1(n5712), .A2(n5702), .ZN(n6633) );
  NAND2_X1 U7248 ( .A1(n5703), .A2(n6633), .ZN(n5704) );
  OAI211_X1 U7249 ( .C1(n6632), .C2(n6513), .A(n5705), .B(n5704), .ZN(n6568)
         );
  INV_X1 U7250 ( .A(n6568), .ZN(n5714) );
  INV_X1 U7251 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9748) );
  INV_X1 U7252 ( .A(n5712), .ZN(n7679) );
  AND2_X1 U7253 ( .A1(n7679), .A2(n7635), .ZN(n5706) );
  AOI21_X1 U7254 ( .B1(n6515), .B2(n9748), .A(n5706), .ZN(n6527) );
  NAND2_X1 U7255 ( .A1(n5708), .A2(n5707), .ZN(n5709) );
  NAND2_X1 U7256 ( .A1(n5709), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5710) );
  XNOR2_X1 U7257 ( .A(n5710), .B(n10370), .ZN(n7612) );
  NAND2_X1 U7258 ( .A1(n6253), .A2(n9001), .ZN(n6566) );
  NAND2_X1 U7259 ( .A1(n9749), .A2(n6566), .ZN(n5713) );
  NOR2_X1 U7260 ( .A1(n6527), .A2(n5713), .ZN(n7029) );
  AND2_X2 U7261 ( .A1(n5714), .A2(n7029), .ZN(n9788) );
  NAND2_X1 U7262 ( .A1(n9438), .A2(n9788), .ZN(n5716) );
  NOR2_X1 U7263 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5719) );
  INV_X1 U7264 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5724) );
  INV_X1 U7265 ( .A(n5722), .ZN(n5721) );
  NAND2_X1 U7266 ( .A1(n5721), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n5723) );
  INV_X1 U7267 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n10436) );
  INV_X1 U7268 ( .A(n8353), .ZN(n6178) );
  NAND2_X1 U7269 ( .A1(n7948), .A2(n6178), .ZN(n9592) );
  NOR2_X1 U7270 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5728) );
  INV_X1 U7271 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5727) );
  NAND4_X1 U7272 ( .A1(n5728), .A2(n5727), .A3(n5726), .A4(n5935), .ZN(n5733)
         );
  INV_X1 U7273 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5730) );
  INV_X1 U7274 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5729) );
  NAND4_X1 U7275 ( .A1(n5731), .A2(n5730), .A3(n5947), .A4(n5729), .ZN(n5732)
         );
  NAND2_X1 U7276 ( .A1(n4554), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5734) );
  XNOR2_X1 U7277 ( .A(n5734), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7991) );
  OR2_X1 U7278 ( .A1(n9592), .A2(n7991), .ZN(n10067) );
  INV_X1 U7279 ( .A(n10067), .ZN(n7051) );
  INV_X1 U7280 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5735) );
  NOR2_X2 U7281 ( .A1(n5748), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5738) );
  INV_X1 U7282 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5739) );
  NAND2_X1 U7283 ( .A1(n5738), .A2(n5739), .ZN(n8665) );
  INV_X1 U7284 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5736) );
  NAND2_X2 U7285 ( .A1(n5741), .A2(n8670), .ZN(n6071) );
  INV_X4 U7286 ( .A(n6071), .ZN(n7218) );
  NAND2_X1 U7287 ( .A1(n7218), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5747) );
  OR2_X1 U7288 ( .A1(n5992), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5746) );
  NAND2_X4 U7289 ( .A1(n5741), .A2(n5742), .ZN(n7217) );
  INV_X1 U7290 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6986) );
  OR2_X1 U7291 ( .A1(n7217), .A2(n6986), .ZN(n5745) );
  INV_X1 U7292 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7120) );
  OR2_X1 U7293 ( .A1(n7220), .A2(n7120), .ZN(n5744) );
  NAND4_X1 U7294 ( .A1(n5747), .A2(n5746), .A3(n5745), .A4(n5744), .ZN(n8243)
         );
  INV_X1 U7295 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5749) );
  INV_X1 U7296 ( .A(n5751), .ZN(n6202) );
  NAND2_X4 U7297 ( .A1(n5752), .A2(n5748), .ZN(n8291) );
  AND2_X1 U7298 ( .A1(n5780), .A2(n4610), .ZN(n5825) );
  NAND2_X1 U7299 ( .A1(n5753), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5754) );
  MUX2_X1 U7300 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5754), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5756) );
  AND2_X1 U7301 ( .A1(n5756), .A2(n5815), .ZN(n7011) );
  NAND2_X1 U7302 ( .A1(n6002), .A2(n7011), .ZN(n5757) );
  INV_X1 U7303 ( .A(n7955), .ZN(n5793) );
  INV_X1 U7304 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7141) );
  OR2_X1 U7305 ( .A1(n5992), .A2(n7141), .ZN(n5762) );
  INV_X1 U7306 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5760) );
  OR2_X1 U7307 ( .A1(n7220), .A2(n5760), .ZN(n5761) );
  NAND2_X1 U7308 ( .A1(n5825), .A2(n6586), .ZN(n5770) );
  NAND2_X1 U7309 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5766) );
  MUX2_X1 U7310 ( .A(n5766), .B(P2_IR_REG_31__SCAN_IN), .S(n5765), .Z(n5768)
         );
  INV_X1 U7311 ( .A(n6784), .ZN(n5767) );
  NAND2_X1 U7312 ( .A1(n6002), .A2(n6854), .ZN(n5769) );
  OAI211_X2 U7313 ( .C1(n7790), .C2(P1_DATAO_REG_1__SCAN_IN), .A(n5770), .B(
        n5769), .ZN(n10047) );
  NAND2_X1 U7314 ( .A1(n8245), .A2(n10047), .ZN(n7817) );
  NAND2_X2 U7315 ( .A1(n7820), .A2(n7817), .ZN(n7954) );
  NAND2_X1 U7316 ( .A1(n7218), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5775) );
  INV_X1 U7317 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10385) );
  OR2_X1 U7318 ( .A1(n5992), .A2(n10385), .ZN(n5774) );
  INV_X1 U7319 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5771) );
  OR2_X1 U7320 ( .A1(n7217), .A2(n5771), .ZN(n5773) );
  INV_X1 U7321 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6783) );
  OR2_X1 U7322 ( .A1(n7220), .A2(n6783), .ZN(n5772) );
  NAND2_X1 U7323 ( .A1(n4610), .A2(SI_0_), .ZN(n5777) );
  INV_X1 U7324 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5776) );
  NAND2_X1 U7325 ( .A1(n5777), .A2(n5776), .ZN(n5779) );
  AND2_X1 U7326 ( .A1(n5779), .A2(n5778), .ZN(n8675) );
  MUX2_X1 U7327 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8675), .S(n5780), .Z(n10044)
         );
  INV_X1 U7328 ( .A(n10044), .ZN(n6888) );
  INV_X1 U7329 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5781) );
  OR2_X1 U7330 ( .A1(n6071), .A2(n5781), .ZN(n5784) );
  INV_X1 U7331 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10021) );
  OR2_X1 U7332 ( .A1(n5992), .A2(n10021), .ZN(n5783) );
  INV_X1 U7333 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6843) );
  OR2_X1 U7334 ( .A1(n7217), .A2(n6843), .ZN(n5782) );
  NAND2_X1 U7335 ( .A1(n7803), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5791) );
  NAND2_X1 U7336 ( .A1(n5825), .A2(n5786), .ZN(n5790) );
  INV_X1 U7337 ( .A(n5753), .ZN(n5787) );
  NAND2_X1 U7338 ( .A1(n6002), .A2(n7008), .ZN(n5789) );
  OR2_X2 U7339 ( .A1(n8244), .A2(n10050), .ZN(n7828) );
  NAND2_X1 U7340 ( .A1(n8244), .A2(n10050), .ZN(n7829) );
  NAND2_X1 U7341 ( .A1(n7828), .A2(n7829), .ZN(n7956) );
  NAND2_X1 U7342 ( .A1(n10019), .A2(n7828), .ZN(n5792) );
  NAND2_X1 U7343 ( .A1(n5793), .A2(n5792), .ZN(n7118) );
  NAND2_X1 U7344 ( .A1(n7118), .A2(n7849), .ZN(n5806) );
  NAND2_X1 U7345 ( .A1(n5794), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5801) );
  INV_X1 U7346 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5795) );
  OR2_X1 U7347 ( .A1(n6071), .A2(n5795), .ZN(n5800) );
  NAND2_X1 U7348 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5797) );
  AND2_X1 U7349 ( .A1(n5809), .A2(n5797), .ZN(n7229) );
  OR2_X1 U7350 ( .A1(n5992), .A2(n7229), .ZN(n5799) );
  INV_X1 U7351 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7014) );
  OR2_X1 U7352 ( .A1(n7217), .A2(n7014), .ZN(n5798) );
  NAND2_X1 U7353 ( .A1(n5825), .A2(n6592), .ZN(n5805) );
  NAND2_X1 U7354 ( .A1(n7803), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U7355 ( .A1(n5815), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5802) );
  XNOR2_X1 U7356 ( .A(n5802), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7015) );
  NAND2_X1 U7357 ( .A1(n6002), .A2(n7015), .ZN(n5803) );
  AND3_X2 U7358 ( .A1(n5805), .A2(n5804), .A3(n5803), .ZN(n7230) );
  OR2_X1 U7359 ( .A1(n8242), .A2(n7230), .ZN(n7836) );
  NAND2_X1 U7360 ( .A1(n8242), .A2(n7230), .ZN(n7852) );
  NAND2_X1 U7361 ( .A1(n7836), .A2(n7852), .ZN(n7053) );
  NAND2_X1 U7362 ( .A1(n5806), .A2(n7957), .ZN(n7052) );
  NAND2_X1 U7363 ( .A1(n7218), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5814) );
  INV_X1 U7364 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6985) );
  OR2_X1 U7365 ( .A1(n7220), .A2(n6985), .ZN(n5813) );
  NAND2_X1 U7366 ( .A1(n5809), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5810) );
  AND2_X1 U7367 ( .A1(n5819), .A2(n5810), .ZN(n7172) );
  OR2_X1 U7368 ( .A1(n5992), .A2(n7172), .ZN(n5812) );
  INV_X1 U7369 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6984) );
  OR2_X1 U7370 ( .A1(n7217), .A2(n6984), .ZN(n5811) );
  NAND4_X1 U7371 ( .A1(n5814), .A2(n5813), .A3(n5812), .A4(n5811), .ZN(n8241)
         );
  NAND2_X1 U7372 ( .A1(n7803), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U7373 ( .A1(n5826), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5816) );
  XNOR2_X1 U7374 ( .A(n5816), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7017) );
  NAND2_X1 U7375 ( .A1(n6002), .A2(n7017), .ZN(n5817) );
  OAI211_X1 U7376 ( .C1(n6110), .C2(n6598), .A(n5818), .B(n5817), .ZN(n7169)
         );
  INV_X1 U7377 ( .A(n7169), .ZN(n7113) );
  OR2_X1 U7378 ( .A1(n8241), .A2(n7113), .ZN(n7855) );
  NAND2_X1 U7379 ( .A1(n8241), .A2(n7113), .ZN(n7851) );
  NAND2_X1 U7380 ( .A1(n7218), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5824) );
  INV_X1 U7381 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7273) );
  OR2_X1 U7382 ( .A1(n7220), .A2(n7273), .ZN(n5823) );
  NAND2_X1 U7383 ( .A1(n5819), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5820) );
  AND2_X1 U7384 ( .A1(n5845), .A2(n5820), .ZN(n7242) );
  OR2_X1 U7385 ( .A1(n5992), .A2(n7242), .ZN(n5822) );
  INV_X1 U7386 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n8308) );
  OR2_X1 U7387 ( .A1(n7217), .A2(n8308), .ZN(n5821) );
  NAND4_X1 U7388 ( .A1(n5824), .A2(n5823), .A3(n5822), .A4(n5821), .ZN(n8240)
         );
  NAND2_X1 U7389 ( .A1(n5825), .A2(n6599), .ZN(n5830) );
  NAND2_X1 U7390 ( .A1(n7803), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5829) );
  NOR2_X1 U7391 ( .A1(n5826), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5840) );
  OR2_X1 U7392 ( .A1(n5840), .A2(n5905), .ZN(n5827) );
  XNOR2_X1 U7393 ( .A(n5827), .B(P2_IR_REG_6__SCAN_IN), .ZN(n8309) );
  NAND2_X1 U7394 ( .A1(n6002), .A2(n8309), .ZN(n5828) );
  NAND2_X1 U7395 ( .A1(n8240), .A2(n10062), .ZN(n7857) );
  NAND2_X1 U7396 ( .A1(n7218), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5838) );
  INV_X1 U7397 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7337) );
  OR2_X1 U7398 ( .A1(n7220), .A2(n7337), .ZN(n5837) );
  NAND2_X1 U7399 ( .A1(n5847), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5833) );
  AND2_X1 U7400 ( .A1(n5870), .A2(n5833), .ZN(n7338) );
  OR2_X1 U7401 ( .A1(n5992), .A2(n7338), .ZN(n5836) );
  INV_X1 U7402 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5834) );
  OR2_X1 U7403 ( .A1(n7217), .A2(n5834), .ZN(n5835) );
  NAND4_X1 U7404 ( .A1(n5838), .A2(n5837), .A3(n5836), .A4(n5835), .ZN(n8238)
         );
  INV_X1 U7405 ( .A(n8238), .ZN(n7563) );
  INV_X2 U7406 ( .A(n6110), .ZN(n7804) );
  NAND2_X1 U7407 ( .A1(n6618), .A2(n7804), .ZN(n5843) );
  INV_X1 U7408 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U7409 ( .A1(n5840), .A2(n5839), .ZN(n5853) );
  NAND2_X1 U7410 ( .A1(n5865), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5841) );
  XNOR2_X1 U7411 ( .A(n5841), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9855) );
  AOI22_X1 U7412 ( .A1(n7803), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6002), .B2(
        n9855), .ZN(n5842) );
  NAND2_X1 U7413 ( .A1(n5843), .A2(n5842), .ZN(n7495) );
  NAND2_X1 U7414 ( .A1(n7563), .A2(n7495), .ZN(n7863) );
  INV_X1 U7415 ( .A(n7863), .ZN(n5858) );
  INV_X1 U7416 ( .A(n7495), .ZN(n10072) );
  NAND2_X1 U7417 ( .A1(n10072), .A2(n8238), .ZN(n7839) );
  NAND2_X1 U7418 ( .A1(n7218), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5852) );
  INV_X1 U7419 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5844) );
  OR2_X1 U7420 ( .A1(n7217), .A2(n5844), .ZN(n5851) );
  NAND2_X1 U7421 ( .A1(n5845), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5846) );
  AND2_X1 U7422 ( .A1(n5847), .A2(n5846), .ZN(n7314) );
  OR2_X1 U7423 ( .A1(n5992), .A2(n7314), .ZN(n5850) );
  INV_X1 U7424 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5848) );
  OR2_X1 U7425 ( .A1(n7220), .A2(n5848), .ZN(n5849) );
  NAND4_X1 U7426 ( .A1(n5852), .A2(n5851), .A3(n5850), .A4(n5849), .ZN(n8239)
         );
  NAND2_X1 U7427 ( .A1(n5853), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5855) );
  INV_X1 U7428 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5854) );
  XNOR2_X1 U7429 ( .A(n5855), .B(n5854), .ZN(n8310) );
  INV_X1 U7430 ( .A(n8310), .ZN(n9843) );
  AOI22_X1 U7431 ( .A1(n7803), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6002), .B2(
        n9843), .ZN(n5857) );
  NAND2_X1 U7432 ( .A1(n6614), .A2(n7804), .ZN(n5856) );
  NAND2_X1 U7433 ( .A1(n8239), .A2(n10066), .ZN(n7332) );
  AND2_X1 U7434 ( .A1(n7839), .A2(n7332), .ZN(n7843) );
  AND2_X1 U7435 ( .A1(n7857), .A2(n5860), .ZN(n5859) );
  NAND2_X1 U7436 ( .A1(n7293), .A2(n5859), .ZN(n5864) );
  INV_X1 U7437 ( .A(n5860), .ZN(n5862) );
  OR2_X1 U7438 ( .A1(n8239), .A2(n10066), .ZN(n7862) );
  NAND2_X1 U7439 ( .A1(n7862), .A2(n7332), .ZN(n7961) );
  AND2_X1 U7440 ( .A1(n7859), .A2(n7863), .ZN(n5861) );
  OAI21_X1 U7441 ( .B1(n5865), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5878) );
  XNOR2_X1 U7442 ( .A(n5878), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9872) );
  AOI22_X1 U7443 ( .A1(n7803), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6002), .B2(
        n9872), .ZN(n5866) );
  NAND2_X1 U7444 ( .A1(n5794), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5876) );
  INV_X1 U7445 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5867) );
  OR2_X1 U7446 ( .A1(n6071), .A2(n5867), .ZN(n5875) );
  INV_X1 U7447 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7448 ( .A1(n5870), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5871) );
  AND2_X1 U7449 ( .A1(n5883), .A2(n5871), .ZN(n7559) );
  OR2_X1 U7450 ( .A1(n5992), .A2(n7559), .ZN(n5874) );
  INV_X1 U7451 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5872) );
  OR2_X1 U7452 ( .A1(n7217), .A2(n5872), .ZN(n5873) );
  NAND2_X1 U7453 ( .A1(n7572), .A2(n7606), .ZN(n7867) );
  NAND2_X1 U7454 ( .A1(n7846), .A2(n7867), .ZN(n7960) );
  NAND2_X1 U7455 ( .A1(n6640), .A2(n7804), .ZN(n5882) );
  NAND2_X1 U7456 ( .A1(n5878), .A2(n5877), .ZN(n5879) );
  NAND2_X1 U7457 ( .A1(n5879), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5880) );
  XNOR2_X1 U7458 ( .A(n5880), .B(P2_IR_REG_10__SCAN_IN), .ZN(n9888) );
  AOI22_X1 U7459 ( .A1(n7803), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6002), .B2(
        n9888), .ZN(n5881) );
  NAND2_X1 U7460 ( .A1(n7218), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5889) );
  INV_X1 U7461 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7451) );
  OR2_X1 U7462 ( .A1(n7220), .A2(n7451), .ZN(n5888) );
  NAND2_X1 U7463 ( .A1(n5883), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5884) );
  AND2_X1 U7464 ( .A1(n5898), .A2(n5884), .ZN(n7602) );
  OR2_X1 U7465 ( .A1(n5992), .A2(n7602), .ZN(n5887) );
  INV_X1 U7466 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5885) );
  OR2_X1 U7467 ( .A1(n7217), .A2(n5885), .ZN(n5886) );
  NAND2_X1 U7468 ( .A1(n7608), .A2(n7646), .ZN(n7868) );
  NAND2_X1 U7469 ( .A1(n6660), .A2(n7804), .ZN(n5896) );
  NAND2_X1 U7470 ( .A1(n5890), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5891) );
  MUX2_X1 U7471 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5891), .S(
        P2_IR_REG_11__SCAN_IN), .Z(n5892) );
  INV_X1 U7472 ( .A(n5892), .ZN(n5894) );
  NOR2_X1 U7473 ( .A1(n5894), .A2(n5893), .ZN(n9904) );
  AOI22_X1 U7474 ( .A1(n7803), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6002), .B2(
        n9904), .ZN(n5895) );
  NAND2_X1 U7475 ( .A1(n5896), .A2(n5895), .ZN(n7639) );
  NAND2_X1 U7476 ( .A1(n7218), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5904) );
  INV_X1 U7477 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5897) );
  OR2_X1 U7478 ( .A1(n7220), .A2(n5897), .ZN(n5903) );
  NAND2_X1 U7479 ( .A1(n5898), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5899) );
  AND2_X1 U7480 ( .A1(n5914), .A2(n5899), .ZN(n7643) );
  OR2_X1 U7481 ( .A1(n5992), .A2(n7643), .ZN(n5902) );
  INV_X1 U7482 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5900) );
  OR2_X1 U7483 ( .A1(n7217), .A2(n5900), .ZN(n5901) );
  NAND4_X1 U7484 ( .A1(n5904), .A2(n5903), .A3(n5902), .A4(n5901), .ZN(n8235)
         );
  OR2_X1 U7485 ( .A1(n7639), .A2(n8118), .ZN(n7879) );
  NAND2_X1 U7486 ( .A1(n7639), .A2(n8118), .ZN(n7877) );
  NAND2_X1 U7487 ( .A1(n6776), .A2(n7804), .ZN(n5911) );
  NOR2_X1 U7488 ( .A1(n5893), .A2(n5905), .ZN(n5907) );
  MUX2_X1 U7489 ( .A(n5907), .B(n5905), .S(n5906), .Z(n5908) );
  INV_X1 U7490 ( .A(n5908), .ZN(n5909) );
  AND2_X1 U7491 ( .A1(n5909), .A2(n5922), .ZN(n9919) );
  AOI22_X1 U7492 ( .A1(n7803), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6002), .B2(
        n9919), .ZN(n5910) );
  NAND2_X1 U7493 ( .A1(n7218), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5920) );
  INV_X1 U7494 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U7495 ( .A1(n5914), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5915) );
  AND2_X1 U7496 ( .A1(n5928), .A2(n5915), .ZN(n8122) );
  OR2_X1 U7497 ( .A1(n5992), .A2(n8122), .ZN(n5919) );
  INV_X1 U7498 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n5916) );
  OR2_X1 U7499 ( .A1(n7217), .A2(n5916), .ZN(n5918) );
  INV_X1 U7500 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8257) );
  OR2_X1 U7501 ( .A1(n7220), .A2(n8257), .ZN(n5917) );
  NAND4_X1 U7502 ( .A1(n5920), .A2(n5919), .A3(n5918), .A4(n5917), .ZN(n8234)
         );
  INV_X1 U7503 ( .A(n8234), .ZN(n9599) );
  NAND2_X1 U7504 ( .A1(n10089), .A2(n9599), .ZN(n7881) );
  NAND2_X1 U7505 ( .A1(n7880), .A2(n7881), .ZN(n7968) );
  INV_X1 U7506 ( .A(n7877), .ZN(n7537) );
  NOR2_X1 U7507 ( .A1(n7968), .A2(n7537), .ZN(n5921) );
  NAND2_X1 U7508 ( .A1(n7505), .A2(n5921), .ZN(n7539) );
  NAND2_X1 U7509 ( .A1(n7539), .A2(n7880), .ZN(n9590) );
  NAND2_X1 U7510 ( .A1(n6800), .A2(n7804), .ZN(n5924) );
  NAND2_X1 U7511 ( .A1(n5922), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5936) );
  XNOR2_X1 U7512 ( .A(n5936), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9936) );
  AOI22_X1 U7513 ( .A1(n7803), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6002), .B2(
        n9936), .ZN(n5923) );
  NAND2_X1 U7514 ( .A1(n7218), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5934) );
  INV_X1 U7515 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5925) );
  OR2_X1 U7516 ( .A1(n7220), .A2(n5925), .ZN(n5933) );
  INV_X1 U7517 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U7518 ( .A1(n5928), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5929) );
  AND2_X1 U7519 ( .A1(n5940), .A2(n5929), .ZN(n9594) );
  OR2_X1 U7520 ( .A1(n5992), .A2(n9594), .ZN(n5932) );
  INV_X1 U7521 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5930) );
  OR2_X1 U7522 ( .A1(n7217), .A2(n5930), .ZN(n5931) );
  NAND4_X1 U7523 ( .A1(n5934), .A2(n5933), .A3(n5932), .A4(n5931), .ZN(n8233)
         );
  INV_X1 U7524 ( .A(n8233), .ZN(n8081) );
  NOR2_X1 U7525 ( .A1(n9591), .A2(n8081), .ZN(n7892) );
  NAND2_X1 U7526 ( .A1(n9591), .A2(n8081), .ZN(n7890) );
  NAND2_X1 U7527 ( .A1(n6822), .A2(n7804), .ZN(n5939) );
  NAND2_X1 U7528 ( .A1(n5936), .A2(n5935), .ZN(n5937) );
  NAND2_X1 U7529 ( .A1(n5937), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5948) );
  XNOR2_X1 U7530 ( .A(n5948), .B(P2_IR_REG_14__SCAN_IN), .ZN(n9952) );
  AOI22_X1 U7531 ( .A1(n7803), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6002), .B2(
        n9952), .ZN(n5938) );
  NAND2_X1 U7532 ( .A1(n7218), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5946) );
  INV_X1 U7533 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n10418) );
  OR2_X1 U7534 ( .A1(n7220), .A2(n10418), .ZN(n5945) );
  NAND2_X1 U7535 ( .A1(n5940), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5941) );
  AND2_X1 U7536 ( .A1(n5955), .A2(n5941), .ZN(n8084) );
  OR2_X1 U7537 ( .A1(n5992), .A2(n8084), .ZN(n5944) );
  INV_X1 U7538 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5942) );
  OR2_X1 U7539 ( .A1(n7217), .A2(n5942), .ZN(n5943) );
  NAND4_X1 U7540 ( .A1(n5946), .A2(n5945), .A3(n5944), .A4(n5943), .ZN(n8232)
         );
  OR2_X1 U7541 ( .A1(n8086), .A2(n9598), .ZN(n7895) );
  NAND2_X1 U7542 ( .A1(n8086), .A2(n9598), .ZN(n7896) );
  NAND2_X1 U7543 ( .A1(n6936), .A2(n7804), .ZN(n5952) );
  NAND2_X1 U7544 ( .A1(n5948), .A2(n5947), .ZN(n5949) );
  NAND2_X1 U7545 ( .A1(n5949), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5950) );
  XNOR2_X1 U7546 ( .A(n5950), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9969) );
  AOI22_X1 U7547 ( .A1(n7803), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6002), .B2(
        n9969), .ZN(n5951) );
  NAND2_X1 U7548 ( .A1(n7218), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5960) );
  INV_X1 U7549 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8599) );
  OR2_X1 U7550 ( .A1(n7217), .A2(n8599), .ZN(n5959) );
  INV_X1 U7551 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U7552 ( .A1(n5955), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5956) );
  AND2_X1 U7553 ( .A1(n5967), .A2(n5956), .ZN(n8213) );
  OR2_X1 U7554 ( .A1(n5992), .A2(n8213), .ZN(n5958) );
  INV_X1 U7555 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7628) );
  OR2_X1 U7556 ( .A1(n7220), .A2(n7628), .ZN(n5957) );
  NAND4_X1 U7557 ( .A1(n5960), .A2(n5959), .A3(n5958), .A4(n5957), .ZN(n8231)
         );
  INV_X1 U7558 ( .A(n8231), .ZN(n8527) );
  AND2_X1 U7559 ( .A1(n8016), .A2(n8527), .ZN(n7898) );
  OR2_X1 U7560 ( .A1(n8016), .A2(n8527), .ZN(n7900) );
  NAND2_X1 U7561 ( .A1(n6956), .A2(n7804), .ZN(n5966) );
  NAND2_X1 U7562 ( .A1(n5961), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5962) );
  MUX2_X1 U7563 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5962), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5964) );
  INV_X1 U7564 ( .A(n5974), .ZN(n5963) );
  NAND2_X1 U7565 ( .A1(n5964), .A2(n5963), .ZN(n8302) );
  INV_X1 U7566 ( .A(n8302), .ZN(n9985) );
  AOI22_X1 U7567 ( .A1(n7803), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6002), .B2(
        n9985), .ZN(n5965) );
  NAND2_X1 U7568 ( .A1(n7218), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5972) );
  INV_X1 U7569 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n10375) );
  OR2_X1 U7570 ( .A1(n7220), .A2(n10375), .ZN(n5971) );
  NAND2_X1 U7571 ( .A1(n5967), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5968) );
  AND2_X1 U7572 ( .A1(n5982), .A2(n5968), .ZN(n8533) );
  OR2_X1 U7573 ( .A1(n5992), .A2(n8533), .ZN(n5970) );
  INV_X1 U7574 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n10323) );
  OR2_X1 U7575 ( .A1(n7217), .A2(n10323), .ZN(n5969) );
  NAND2_X1 U7576 ( .A1(n8531), .A2(n8211), .ZN(n7815) );
  INV_X1 U7577 ( .A(n7816), .ZN(n5973) );
  NAND2_X1 U7578 ( .A1(n7082), .A2(n7804), .ZN(n5979) );
  NOR2_X1 U7579 ( .A1(n5974), .A2(n5905), .ZN(n5975) );
  MUX2_X1 U7580 ( .A(n5905), .B(n5975), .S(P2_IR_REG_17__SCAN_IN), .Z(n5976)
         );
  INV_X1 U7581 ( .A(n5976), .ZN(n5977) );
  AND2_X1 U7582 ( .A1(n5977), .A2(n5988), .ZN(n10003) );
  AOI22_X1 U7583 ( .A1(n7803), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6002), .B2(
        n10003), .ZN(n5978) );
  NAND2_X1 U7584 ( .A1(n7218), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5987) );
  INV_X1 U7585 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n10013) );
  OR2_X1 U7586 ( .A1(n7220), .A2(n10013), .ZN(n5986) );
  INV_X1 U7587 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U7588 ( .A1(n5982), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5983) );
  AND2_X1 U7589 ( .A1(n5993), .A2(n5983), .ZN(n8517) );
  OR2_X1 U7590 ( .A1(n5992), .A2(n8517), .ZN(n5985) );
  INV_X1 U7591 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8265) );
  OR2_X1 U7592 ( .A1(n7217), .A2(n8265), .ZN(n5984) );
  OR2_X1 U7593 ( .A1(n8590), .A2(n8528), .ZN(n7906) );
  NAND2_X1 U7594 ( .A1(n8590), .A2(n8528), .ZN(n8498) );
  NAND2_X1 U7595 ( .A1(n7906), .A2(n8498), .ZN(n6155) );
  NAND2_X1 U7596 ( .A1(n7145), .A2(n7804), .ZN(n5991) );
  NAND2_X1 U7597 ( .A1(n5988), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5989) );
  XNOR2_X1 U7598 ( .A(n5989), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8340) );
  AOI22_X1 U7599 ( .A1(n7803), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6002), .B2(
        n8340), .ZN(n5990) );
  NAND2_X1 U7600 ( .A1(n5993), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U7601 ( .A1(n6009), .A2(n5994), .ZN(n8504) );
  NAND2_X1 U7602 ( .A1(n6111), .A2(n8504), .ZN(n5999) );
  INV_X1 U7603 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n5995) );
  OR2_X1 U7604 ( .A1(n7220), .A2(n5995), .ZN(n5998) );
  INV_X1 U7605 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n10487) );
  OR2_X1 U7606 ( .A1(n6071), .A2(n10487), .ZN(n5997) );
  INV_X1 U7607 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8588) );
  OR2_X1 U7608 ( .A1(n7217), .A2(n8588), .ZN(n5996) );
  NAND4_X1 U7609 ( .A1(n5999), .A2(n5998), .A3(n5997), .A4(n5996), .ZN(n8512)
         );
  INV_X1 U7610 ( .A(n8512), .ZN(n8103) );
  NAND2_X1 U7611 ( .A1(n8503), .A2(n8103), .ZN(n7907) );
  NAND2_X1 U7612 ( .A1(n7910), .A2(n7907), .ZN(n8502) );
  INV_X1 U7613 ( .A(n8498), .ZN(n6000) );
  NOR2_X1 U7614 ( .A1(n8502), .A2(n6000), .ZN(n6001) );
  NAND2_X1 U7615 ( .A1(n8520), .A2(n6001), .ZN(n8499) );
  NAND2_X1 U7616 ( .A1(n8499), .A2(n7910), .ZN(n8488) );
  NAND2_X1 U7617 ( .A1(n7306), .A2(n7804), .ZN(n6004) );
  AOI22_X1 U7618 ( .A1(n7803), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6178), .B2(
        n6002), .ZN(n6003) );
  INV_X1 U7619 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8337) );
  OR2_X1 U7620 ( .A1(n7220), .A2(n8337), .ZN(n6006) );
  INV_X1 U7621 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n10388) );
  OR2_X1 U7622 ( .A1(n6071), .A2(n10388), .ZN(n6005) );
  AND2_X1 U7623 ( .A1(n6006), .A2(n6005), .ZN(n6013) );
  INV_X1 U7624 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7625 ( .A1(n6009), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7626 ( .A1(n6016), .A2(n6010), .ZN(n8490) );
  NAND2_X1 U7627 ( .A1(n8490), .A2(n6111), .ZN(n6012) );
  NAND2_X1 U7628 ( .A1(n6068), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7629 ( .A1(n8489), .A2(n8497), .ZN(n7915) );
  NAND2_X1 U7630 ( .A1(n7414), .A2(n7804), .ZN(n6015) );
  NAND2_X1 U7631 ( .A1(n7803), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7632 ( .A1(n6016), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7633 ( .A1(n6025), .A2(n6017), .ZN(n8471) );
  NAND2_X1 U7634 ( .A1(n8471), .A2(n6111), .ZN(n6020) );
  AOI22_X1 U7635 ( .A1(n5794), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n7218), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n6019) );
  INV_X1 U7636 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n10234) );
  OR2_X1 U7637 ( .A1(n7217), .A2(n10234), .ZN(n6018) );
  NAND2_X1 U7638 ( .A1(n8470), .A2(n8456), .ZN(n8460) );
  NAND2_X1 U7639 ( .A1(n7474), .A2(n7804), .ZN(n6022) );
  NAND2_X1 U7640 ( .A1(n7803), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6021) );
  INV_X1 U7641 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7642 ( .A1(n6025), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U7643 ( .A1(n6033), .A2(n6026), .ZN(n8465) );
  NAND2_X1 U7644 ( .A1(n8465), .A2(n6111), .ZN(n6029) );
  AOI22_X1 U7645 ( .A1(n6068), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n7218), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U7646 ( .A1(n5794), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6027) );
  NAND2_X1 U7647 ( .A1(n8464), .A2(n8478), .ZN(n7919) );
  AND2_X1 U7648 ( .A1(n8460), .A2(n7919), .ZN(n7913) );
  NAND2_X1 U7649 ( .A1(n8461), .A2(n7913), .ZN(n6030) );
  NAND2_X1 U7650 ( .A1(n6030), .A2(n7917), .ZN(n8450) );
  NAND2_X1 U7651 ( .A1(n7547), .A2(n7804), .ZN(n6032) );
  NAND2_X1 U7652 ( .A1(n7803), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7653 ( .A1(n6033), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7654 ( .A1(n6043), .A2(n6034), .ZN(n8448) );
  NAND2_X1 U7655 ( .A1(n8448), .A2(n6111), .ZN(n6039) );
  INV_X1 U7656 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8634) );
  NAND2_X1 U7657 ( .A1(n5794), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7658 ( .A1(n6068), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6035) );
  OAI211_X1 U7659 ( .C1(n6071), .C2(n8634), .A(n6036), .B(n6035), .ZN(n6037)
         );
  INV_X1 U7660 ( .A(n6037), .ZN(n6038) );
  NAND2_X1 U7661 ( .A1(n8568), .A2(n8457), .ZN(n7924) );
  INV_X1 U7662 ( .A(n7925), .ZN(n6040) );
  NAND2_X1 U7663 ( .A1(n7611), .A2(n7804), .ZN(n6042) );
  NAND2_X1 U7664 ( .A1(n7803), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U7665 ( .A1(n6043), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U7666 ( .A1(n6054), .A2(n6044), .ZN(n8439) );
  NAND2_X1 U7667 ( .A1(n8439), .A2(n6111), .ZN(n6049) );
  INV_X1 U7668 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8566) );
  NAND2_X1 U7669 ( .A1(n7218), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6046) );
  NAND2_X1 U7670 ( .A1(n5794), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6045) );
  OAI211_X1 U7671 ( .C1(n7217), .C2(n8566), .A(n6046), .B(n6045), .ZN(n6047)
         );
  INV_X1 U7672 ( .A(n6047), .ZN(n6048) );
  NAND2_X1 U7673 ( .A1(n6049), .A2(n6048), .ZN(n8226) );
  NAND2_X1 U7674 ( .A1(n7633), .A2(n7804), .ZN(n6051) );
  NAND2_X1 U7675 ( .A1(n7803), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6050) );
  INV_X1 U7676 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7677 ( .A1(n6054), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U7678 ( .A1(n6066), .A2(n6055), .ZN(n8419) );
  NAND2_X1 U7679 ( .A1(n8419), .A2(n6111), .ZN(n6061) );
  INV_X1 U7680 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7681 ( .A1(n7218), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U7682 ( .A1(n6068), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6056) );
  OAI211_X1 U7683 ( .C1(n6058), .C2(n7220), .A(n6057), .B(n6056), .ZN(n6059)
         );
  INV_X1 U7684 ( .A(n6059), .ZN(n6060) );
  NAND2_X1 U7685 ( .A1(n6061), .A2(n6060), .ZN(n8225) );
  NAND2_X1 U7686 ( .A1(n8421), .A2(n8436), .ZN(n7950) );
  NAND2_X1 U7687 ( .A1(n8438), .A2(n8447), .ZN(n8423) );
  NAND2_X1 U7688 ( .A1(n7950), .A2(n8423), .ZN(n7928) );
  NAND2_X1 U7689 ( .A1(n7666), .A2(n7804), .ZN(n6063) );
  NAND2_X1 U7690 ( .A1(n7803), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6062) );
  INV_X1 U7691 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7692 ( .A1(n6066), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7693 ( .A1(n6075), .A2(n6067), .ZN(n8408) );
  NAND2_X1 U7694 ( .A1(n8408), .A2(n6111), .ZN(n6074) );
  INV_X1 U7695 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n10297) );
  NAND2_X1 U7696 ( .A1(n5794), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7697 ( .A1(n6068), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6069) );
  OAI211_X1 U7698 ( .C1(n6071), .C2(n10297), .A(n6070), .B(n6069), .ZN(n6072)
         );
  INV_X1 U7699 ( .A(n6072), .ZN(n6073) );
  NAND2_X1 U7700 ( .A1(n6074), .A2(n6073), .ZN(n8415) );
  NAND2_X1 U7701 ( .A1(n8407), .A2(n8395), .ZN(n7933) );
  NAND2_X1 U7702 ( .A1(n6075), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7703 ( .A1(n6088), .A2(n6076), .ZN(n8399) );
  NAND2_X1 U7704 ( .A1(n8399), .A2(n6111), .ZN(n6081) );
  INV_X1 U7705 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8553) );
  NAND2_X1 U7706 ( .A1(n5794), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7707 ( .A1(n7218), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6077) );
  OAI211_X1 U7708 ( .C1(n8553), .C2(n7217), .A(n6078), .B(n6077), .ZN(n6079)
         );
  INV_X1 U7709 ( .A(n6079), .ZN(n6080) );
  NAND2_X1 U7710 ( .A1(n6081), .A2(n6080), .ZN(n8224) );
  NAND2_X1 U7711 ( .A1(n7677), .A2(n7804), .ZN(n6083) );
  NAND2_X1 U7712 ( .A1(n7803), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6082) );
  NAND2_X1 U7713 ( .A1(n7721), .A2(n7804), .ZN(n6085) );
  NAND2_X1 U7714 ( .A1(n7803), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6084) );
  INV_X1 U7715 ( .A(n6088), .ZN(n6087) );
  INV_X1 U7716 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7717 ( .A1(n6087), .A2(n6086), .ZN(n6097) );
  NAND2_X1 U7718 ( .A1(n6088), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7719 ( .A1(n6097), .A2(n6089), .ZN(n8387) );
  NAND2_X1 U7720 ( .A1(n8387), .A2(n6111), .ZN(n6094) );
  INV_X1 U7721 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U7722 ( .A1(n5794), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7723 ( .A1(n7218), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6090) );
  OAI211_X1 U7724 ( .C1(n8549), .C2(n7217), .A(n6091), .B(n6090), .ZN(n6092)
         );
  INV_X1 U7725 ( .A(n6092), .ZN(n6093) );
  NAND2_X1 U7726 ( .A1(n8386), .A2(n8396), .ZN(n7936) );
  AOI21_X2 U7727 ( .B1(n8384), .B2(n7936), .A(n7937), .ZN(n7998) );
  NAND2_X1 U7728 ( .A1(n8671), .A2(n7804), .ZN(n6096) );
  NAND2_X1 U7729 ( .A1(n7803), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7730 ( .A1(n6097), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7731 ( .A1(n8361), .A2(n6098), .ZN(n8376) );
  NAND2_X1 U7732 ( .A1(n8376), .A2(n6111), .ZN(n6103) );
  INV_X1 U7733 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U7734 ( .A1(n7218), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U7735 ( .A1(n5794), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6099) );
  OAI211_X1 U7736 ( .C1(n7217), .C2(n8545), .A(n6100), .B(n6099), .ZN(n6101)
         );
  INV_X1 U7737 ( .A(n6101), .ZN(n6102) );
  MUX2_X1 U7738 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n5082), .Z(n7785) );
  NAND2_X1 U7739 ( .A1(n7803), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6109) );
  INV_X1 U7740 ( .A(n8361), .ZN(n6112) );
  NAND2_X1 U7741 ( .A1(n6112), .A2(n6111), .ZN(n7226) );
  INV_X1 U7742 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6233) );
  NAND2_X1 U7743 ( .A1(n7218), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7744 ( .A1(n5794), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6113) );
  OAI211_X1 U7745 ( .C1(n7217), .C2(n6233), .A(n6114), .B(n6113), .ZN(n6115)
         );
  INV_X1 U7746 ( .A(n6115), .ZN(n6116) );
  NAND2_X1 U7747 ( .A1(n6232), .A2(n8062), .ZN(n7793) );
  INV_X1 U7748 ( .A(n6891), .ZN(n6119) );
  INV_X1 U7749 ( .A(n7825), .ZN(n7498) );
  INV_X1 U7750 ( .A(n7991), .ZN(n7551) );
  AND2_X1 U7751 ( .A1(n6904), .A2(n10077), .ZN(n7135) );
  NAND2_X1 U7752 ( .A1(n8353), .A2(n7991), .ZN(n6224) );
  NAND2_X1 U7753 ( .A1(n6119), .A2(n6224), .ZN(n6120) );
  NAND2_X1 U7754 ( .A1(n8366), .A2(n7296), .ZN(n6189) );
  INV_X1 U7755 ( .A(n8421), .ZN(n8628) );
  NAND2_X1 U7756 ( .A1(n8246), .A2(n10044), .ZN(n7139) );
  INV_X1 U7757 ( .A(n10047), .ZN(n6121) );
  OR2_X1 U7758 ( .A1(n8245), .A2(n6121), .ZN(n10024) );
  NAND2_X1 U7759 ( .A1(n10026), .A2(n10024), .ZN(n6122) );
  NAND2_X1 U7760 ( .A1(n6122), .A2(n7956), .ZN(n10028) );
  INV_X1 U7761 ( .A(n10050), .ZN(n6894) );
  OR2_X1 U7762 ( .A1(n8244), .A2(n6894), .ZN(n6123) );
  NAND2_X1 U7763 ( .A1(n8243), .A2(n7122), .ZN(n6124) );
  OR2_X1 U7764 ( .A1(n8243), .A2(n7122), .ZN(n7056) );
  INV_X1 U7765 ( .A(n7230), .ZN(n7093) );
  OR2_X1 U7766 ( .A1(n8242), .A2(n7093), .ZN(n6127) );
  AND2_X1 U7767 ( .A1(n7056), .A2(n6127), .ZN(n7063) );
  NOR2_X1 U7768 ( .A1(n8241), .A2(n7169), .ZN(n6129) );
  INV_X1 U7769 ( .A(n6129), .ZN(n6125) );
  AND2_X1 U7770 ( .A1(n7063), .A2(n6125), .ZN(n6126) );
  NAND2_X1 U7771 ( .A1(n7055), .A2(n6126), .ZN(n6132) );
  INV_X1 U7772 ( .A(n6127), .ZN(n6128) );
  OR2_X1 U7773 ( .A1(n6128), .A2(n7053), .ZN(n7064) );
  OR2_X1 U7774 ( .A1(n6129), .A2(n7064), .ZN(n6131) );
  NAND2_X1 U7775 ( .A1(n8241), .A2(n7169), .ZN(n6130) );
  NAND3_X1 U7776 ( .A1(n6132), .A2(n6131), .A3(n6130), .ZN(n7271) );
  NAND2_X1 U7777 ( .A1(n7854), .A2(n7857), .ZN(n7959) );
  NAND2_X1 U7778 ( .A1(n7271), .A2(n7959), .ZN(n6134) );
  INV_X1 U7779 ( .A(n10062), .ZN(n7275) );
  NAND2_X1 U7780 ( .A1(n8240), .A2(n7275), .ZN(n6133) );
  INV_X1 U7781 ( .A(n8239), .ZN(n7487) );
  NAND2_X1 U7782 ( .A1(n7487), .A2(n10066), .ZN(n6135) );
  NAND2_X1 U7783 ( .A1(n7495), .A2(n8238), .ZN(n6136) );
  NAND2_X1 U7784 ( .A1(n7335), .A2(n6136), .ZN(n6138) );
  OR2_X1 U7785 ( .A1(n8238), .A2(n7495), .ZN(n6137) );
  NAND2_X1 U7786 ( .A1(n7639), .A2(n8235), .ZN(n6142) );
  INV_X1 U7787 ( .A(n6142), .ZN(n6141) );
  OR2_X1 U7788 ( .A1(n7639), .A2(n8235), .ZN(n6139) );
  INV_X1 U7789 ( .A(n7646), .ZN(n8236) );
  OR2_X1 U7790 ( .A1(n7608), .A2(n8236), .ZN(n7501) );
  AND2_X1 U7791 ( .A1(n6139), .A2(n7501), .ZN(n6140) );
  INV_X1 U7792 ( .A(n6147), .ZN(n6144) );
  NAND2_X1 U7793 ( .A1(n7870), .A2(n7868), .ZN(n7499) );
  AND2_X1 U7794 ( .A1(n7499), .A2(n6142), .ZN(n6143) );
  NAND2_X1 U7795 ( .A1(n7447), .A2(n6145), .ZN(n6151) );
  INV_X1 U7796 ( .A(n6146), .ZN(n6149) );
  INV_X1 U7797 ( .A(n7606), .ZN(n8237) );
  OR2_X1 U7798 ( .A1(n7572), .A2(n8237), .ZN(n7448) );
  AND2_X1 U7799 ( .A1(n7448), .A2(n6147), .ZN(n6148) );
  NOR2_X1 U7800 ( .A1(n9591), .A2(n8233), .ZN(n7887) );
  NAND2_X1 U7801 ( .A1(n9591), .A2(n8233), .ZN(n7885) );
  AND2_X1 U7802 ( .A1(n8086), .A2(n8232), .ZN(n6152) );
  NAND2_X1 U7803 ( .A1(n8016), .A2(n8231), .ZN(n7623) );
  NAND2_X1 U7804 ( .A1(n7625), .A2(n7623), .ZN(n6153) );
  OR2_X1 U7805 ( .A1(n8016), .A2(n8231), .ZN(n7624) );
  NAND2_X1 U7806 ( .A1(n6153), .A2(n7624), .ZN(n8525) );
  INV_X1 U7807 ( .A(n8211), .ZN(n8514) );
  NAND2_X1 U7808 ( .A1(n8531), .A2(n8514), .ZN(n6154) );
  NAND2_X1 U7809 ( .A1(n8510), .A2(n6155), .ZN(n6157) );
  INV_X1 U7810 ( .A(n8528), .ZN(n8230) );
  NAND2_X1 U7811 ( .A1(n8590), .A2(n8230), .ZN(n6156) );
  AND2_X1 U7812 ( .A1(n8503), .A2(n8512), .ZN(n6158) );
  INV_X1 U7813 ( .A(n8497), .ZN(n8229) );
  NAND2_X1 U7814 ( .A1(n8489), .A2(n8229), .ZN(n6160) );
  AND2_X2 U7815 ( .A1(n8483), .A2(n6160), .ZN(n8475) );
  NAND2_X1 U7816 ( .A1(n7916), .A2(n8460), .ZN(n8474) );
  INV_X1 U7817 ( .A(n8456), .ZN(n8485) );
  OR2_X1 U7818 ( .A1(n8470), .A2(n8485), .ZN(n6161) );
  NAND2_X1 U7819 ( .A1(n7917), .A2(n7919), .ZN(n8454) );
  INV_X1 U7820 ( .A(n8454), .ZN(n8462) );
  OR2_X1 U7821 ( .A1(n8438), .A2(n8226), .ZN(n6162) );
  OR2_X1 U7822 ( .A1(n8568), .A2(n8227), .ZN(n8432) );
  NAND2_X1 U7823 ( .A1(n6162), .A2(n8432), .ZN(n6163) );
  NAND2_X1 U7824 ( .A1(n8438), .A2(n8226), .ZN(n6164) );
  NAND2_X1 U7825 ( .A1(n6163), .A2(n6164), .ZN(n6166) );
  NAND2_X1 U7826 ( .A1(n8449), .A2(n6164), .ZN(n6165) );
  NOR2_X1 U7827 ( .A1(n8462), .A2(n6168), .ZN(n6169) );
  INV_X1 U7828 ( .A(n8478), .ZN(n8228) );
  OR2_X1 U7829 ( .A1(n8464), .A2(n8228), .ZN(n8430) );
  AND2_X1 U7830 ( .A1(n8430), .A2(n6166), .ZN(n6167) );
  INV_X1 U7831 ( .A(n8407), .ZN(n8624) );
  INV_X1 U7832 ( .A(n8396), .ZN(n8223) );
  NOR2_X1 U7833 ( .A1(n8066), .A2(n8222), .ZN(n6175) );
  OAI22_X1 U7834 ( .A1(n7999), .A2(n6175), .B1(n8383), .B2(n4731), .ZN(n6176)
         );
  XNOR2_X1 U7835 ( .A(n6176), .B(n7976), .ZN(n6186) );
  INV_X1 U7836 ( .A(n7948), .ZN(n6177) );
  NAND2_X1 U7837 ( .A1(n7825), .A2(n6177), .ZN(n7986) );
  NAND2_X1 U7838 ( .A1(n6178), .A2(n7991), .ZN(n6239) );
  INV_X1 U7839 ( .A(n7989), .ZN(n6759) );
  INV_X1 U7840 ( .A(n8291), .ZN(n8346) );
  NAND2_X1 U7841 ( .A1(n6759), .A2(n8346), .ZN(n6179) );
  NAND2_X1 U7842 ( .A1(n5780), .A2(n6179), .ZN(n6903) );
  INV_X1 U7843 ( .A(n6903), .ZN(n6886) );
  INV_X1 U7844 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n10269) );
  NAND2_X1 U7845 ( .A1(n5794), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U7846 ( .A1(n7218), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6180) );
  OAI211_X1 U7847 ( .C1(n10269), .C2(n7217), .A(n6181), .B(n6180), .ZN(n6182)
         );
  INV_X1 U7848 ( .A(n6182), .ZN(n6183) );
  NAND2_X1 U7849 ( .A1(n7226), .A2(n6183), .ZN(n8221) );
  AND2_X1 U7850 ( .A1(n5780), .A2(P2_B_REG_SCAN_IN), .ZN(n6184) );
  NOR2_X1 U7851 ( .A1(n10032), .A2(n6184), .ZN(n8359) );
  AOI22_X1 U7852 ( .A1(n8513), .A2(n8222), .B1(n8221), .B2(n8359), .ZN(n6185)
         );
  OAI21_X1 U7853 ( .B1(n6186), .B2(n10041), .A(n6185), .ZN(n6187) );
  INV_X1 U7854 ( .A(n6187), .ZN(n6188) );
  NAND2_X1 U7855 ( .A1(n6189), .A2(n6188), .ZN(n8367) );
  NAND2_X1 U7856 ( .A1(n6190), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6219) );
  INV_X1 U7857 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U7858 ( .A1(n6219), .A2(n6218), .ZN(n6191) );
  NAND2_X1 U7859 ( .A1(n6191), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6195) );
  INV_X1 U7860 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7861 ( .A1(n6195), .A2(n6194), .ZN(n6197) );
  NAND2_X1 U7862 ( .A1(n6197), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6193) );
  INV_X1 U7863 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6192) );
  XNOR2_X1 U7864 ( .A(n6193), .B(n6192), .ZN(n7690) );
  OR2_X1 U7865 ( .A1(n6195), .A2(n6194), .ZN(n6196) );
  NAND2_X1 U7866 ( .A1(n6197), .A2(n6196), .ZN(n7653) );
  XNOR2_X1 U7867 ( .A(n7653), .B(P2_B_REG_SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7868 ( .A1(n7690), .A2(n6198), .ZN(n6203) );
  NAND2_X1 U7869 ( .A1(n6199), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6200) );
  MUX2_X1 U7870 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6200), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6201) );
  AND2_X1 U7871 ( .A1(n6202), .A2(n6201), .ZN(n6215) );
  NAND2_X1 U7872 ( .A1(n6203), .A2(n6215), .ZN(n6603) );
  NOR2_X1 U7873 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6207) );
  NOR4_X1 U7874 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n6206) );
  NOR4_X1 U7875 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6205) );
  NOR4_X1 U7876 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n6204) );
  NAND4_X1 U7877 ( .A1(n6207), .A2(n6206), .A3(n6205), .A4(n6204), .ZN(n6213)
         );
  NOR4_X1 U7878 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6211) );
  NOR4_X1 U7879 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6210) );
  NOR4_X1 U7880 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6209) );
  NOR4_X1 U7881 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6208) );
  NAND4_X1 U7882 ( .A1(n6211), .A2(n6210), .A3(n6209), .A4(n6208), .ZN(n6212)
         );
  NOR2_X1 U7883 ( .A1(n6213), .A2(n6212), .ZN(n6214) );
  OR2_X1 U7884 ( .A1(n6603), .A2(n6214), .ZN(n6236) );
  INV_X1 U7885 ( .A(n7690), .ZN(n6217) );
  NOR2_X1 U7886 ( .A1(n7653), .A2(n7692), .ZN(n6216) );
  NAND2_X1 U7887 ( .A1(n6217), .A2(n6216), .ZN(n6864) );
  XNOR2_X1 U7888 ( .A(n6219), .B(n6218), .ZN(n6871) );
  AND2_X1 U7889 ( .A1(n6236), .A2(n6883), .ZN(n6242) );
  OR2_X1 U7890 ( .A1(n7947), .A2(n6891), .ZN(n6865) );
  AND2_X1 U7891 ( .A1(n6242), .A2(n6865), .ZN(n6223) );
  OR2_X1 U7892 ( .A1(n6603), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7893 ( .A1(n7653), .A2(n7692), .ZN(n6604) );
  OR2_X1 U7894 ( .A1(n6603), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6222) );
  NAND2_X1 U7895 ( .A1(n7690), .A2(n7692), .ZN(n6221) );
  NAND2_X1 U7896 ( .A1(n7070), .A2(n7069), .ZN(n6862) );
  OR2_X1 U7897 ( .A1(n10067), .A2(n7825), .ZN(n6882) );
  NAND2_X1 U7898 ( .A1(n7070), .A2(n6882), .ZN(n6226) );
  OR2_X1 U7899 ( .A1(n7948), .A2(n6224), .ZN(n6225) );
  AND2_X1 U7900 ( .A1(n7947), .A2(n6225), .ZN(n7068) );
  NAND2_X1 U7901 ( .A1(n6226), .A2(n7068), .ZN(n6230) );
  INV_X1 U7902 ( .A(n7068), .ZN(n6228) );
  INV_X1 U7903 ( .A(n7069), .ZN(n6227) );
  NAND2_X1 U7904 ( .A1(n6228), .A2(n6227), .ZN(n6229) );
  AND2_X2 U7905 ( .A1(n7071), .A2(n6231), .ZN(n10105) );
  NOR2_X1 U7906 ( .A1(n10105), .A2(n6233), .ZN(n6234) );
  OAI21_X1 U7907 ( .B1(n6250), .B2(n10103), .A(n6235), .ZN(P2_U3488) );
  INV_X1 U7908 ( .A(n6236), .ZN(n6863) );
  NOR2_X1 U7909 ( .A1(n7069), .A2(n6863), .ZN(n6238) );
  INV_X1 U7910 ( .A(n7070), .ZN(n6237) );
  AND2_X1 U7911 ( .A1(n6238), .A2(n6237), .ZN(n6872) );
  INV_X1 U7912 ( .A(n6239), .ZN(n6240) );
  NAND2_X1 U7913 ( .A1(n7982), .A2(n6240), .ZN(n6868) );
  AND2_X1 U7914 ( .A1(n10077), .A2(n7947), .ZN(n6241) );
  NAND2_X1 U7915 ( .A1(n6868), .A2(n6241), .ZN(n6877) );
  INV_X1 U7916 ( .A(n9592), .ZN(n7076) );
  NAND2_X1 U7917 ( .A1(n6877), .A2(n10023), .ZN(n6861) );
  NAND2_X1 U7918 ( .A1(n6906), .A2(n6861), .ZN(n6246) );
  INV_X1 U7919 ( .A(n6868), .ZN(n6876) );
  INV_X1 U7920 ( .A(n6904), .ZN(n6244) );
  INV_X1 U7921 ( .A(n6242), .ZN(n6243) );
  NOR2_X1 U7922 ( .A1(n6862), .A2(n6243), .ZN(n6881) );
  OAI21_X1 U7923 ( .B1(n6876), .B2(n6244), .A(n6881), .ZN(n6245) );
  INV_X2 U7924 ( .A(n10093), .ZN(n10091) );
  INV_X1 U7925 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6247) );
  NOR2_X1 U7926 ( .A1(n10091), .A2(n6247), .ZN(n6248) );
  OAI21_X1 U7927 ( .B1(n6250), .B2(n10093), .A(n6249), .ZN(P2_U3456) );
  INV_X1 U7928 ( .A(n6253), .ZN(n6256) );
  INV_X1 U7929 ( .A(n6254), .ZN(n6255) );
  NAND2_X1 U7930 ( .A1(n6256), .A2(n6255), .ZN(n6257) );
  NAND3_X2 U7931 ( .A1(n7194), .A2(n6257), .A3(n6261), .ZN(n6331) );
  NAND2_X1 U7932 ( .A1(n6258), .A2(n9023), .ZN(n6259) );
  NAND2_X1 U7933 ( .A1(n6259), .A2(n9008), .ZN(n6260) );
  NAND2_X2 U7934 ( .A1(n6260), .A2(n6261), .ZN(n6274) );
  NAND2_X2 U7935 ( .A1(n6331), .A2(n6274), .ZN(n6294) );
  INV_X2 U7936 ( .A(n6266), .ZN(n6484) );
  NAND2_X1 U7937 ( .A1(n6484), .A2(n6265), .ZN(n6263) );
  INV_X1 U7938 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6264) );
  INV_X1 U7939 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6656) );
  INV_X1 U7940 ( .A(n6331), .ZN(n6298) );
  NAND2_X1 U7941 ( .A1(n6298), .A2(n6265), .ZN(n6268) );
  NAND2_X1 U7942 ( .A1(n6496), .A2(n9755), .ZN(n6267) );
  OAI211_X1 U7943 ( .C1(n6656), .C2(n6261), .A(n6268), .B(n6267), .ZN(n6645)
         );
  NAND2_X1 U7944 ( .A1(n6644), .A2(n6645), .ZN(n6271) );
  NAND2_X1 U7945 ( .A1(n6271), .A2(n6270), .ZN(n6746) );
  NAND2_X1 U7946 ( .A1(n6294), .A2(n7153), .ZN(n6273) );
  NAND2_X1 U7947 ( .A1(n6276), .A2(n6496), .ZN(n6272) );
  NAND2_X1 U7948 ( .A1(n6273), .A2(n6272), .ZN(n6275) );
  AOI22_X1 U7949 ( .A1(n6298), .A2(n6276), .B1(n6484), .B2(n7153), .ZN(n6278)
         );
  NAND2_X1 U7950 ( .A1(n6277), .A2(n6278), .ZN(n6747) );
  NAND2_X1 U7951 ( .A1(n6746), .A2(n6747), .ZN(n6281) );
  NAND2_X1 U7952 ( .A1(n6281), .A2(n6748), .ZN(n6765) );
  INV_X1 U7953 ( .A(n6765), .ZN(n6292) );
  NAND2_X1 U7954 ( .A1(n6294), .A2(n6772), .ZN(n6283) );
  NAND2_X1 U7955 ( .A1(n6484), .A2(n6285), .ZN(n6282) );
  NAND2_X1 U7956 ( .A1(n6283), .A2(n6282), .ZN(n6284) );
  XNOR2_X1 U7957 ( .A(n6284), .B(n6509), .ZN(n6286) );
  AOI22_X1 U7958 ( .A1(n6298), .A2(n6285), .B1(n6484), .B2(n6772), .ZN(n6287)
         );
  NAND2_X1 U7959 ( .A1(n6286), .A2(n6287), .ZN(n6293) );
  INV_X1 U7960 ( .A(n6286), .ZN(n6289) );
  INV_X1 U7961 ( .A(n6287), .ZN(n6288) );
  NAND2_X1 U7962 ( .A1(n6289), .A2(n6288), .ZN(n6290) );
  NAND2_X1 U7963 ( .A1(n6293), .A2(n6290), .ZN(n6768) );
  INV_X1 U7964 ( .A(n6768), .ZN(n6291) );
  NAND2_X1 U7965 ( .A1(n6292), .A2(n6291), .ZN(n6766) );
  NAND2_X1 U7966 ( .A1(n6319), .A2(n6804), .ZN(n6296) );
  NAND2_X1 U7967 ( .A1(n9098), .A2(n6496), .ZN(n6295) );
  NAND2_X1 U7968 ( .A1(n6296), .A2(n6295), .ZN(n6297) );
  XNOR2_X1 U7969 ( .A(n6297), .B(n6274), .ZN(n6299) );
  AOI22_X1 U7970 ( .A1(n6482), .A2(n9098), .B1(n6484), .B2(n6804), .ZN(n6300)
         );
  XNOR2_X1 U7971 ( .A(n6299), .B(n6300), .ZN(n6816) );
  NAND2_X1 U7972 ( .A1(n6815), .A2(n6816), .ZN(n6814) );
  INV_X1 U7973 ( .A(n6299), .ZN(n6301) );
  NAND2_X1 U7974 ( .A1(n6301), .A2(n6300), .ZN(n6302) );
  NAND2_X1 U7975 ( .A1(n6814), .A2(n6302), .ZN(n6824) );
  INV_X1 U7976 ( .A(n6824), .ZN(n6307) );
  NAND2_X1 U7977 ( .A1(n6496), .A2(n9097), .ZN(n6304) );
  NAND2_X1 U7978 ( .A1(n4505), .A2(n6943), .ZN(n6303) );
  AOI22_X1 U7979 ( .A1(n6482), .A2(n9097), .B1(n6484), .B2(n6943), .ZN(n6308)
         );
  XNOR2_X1 U7980 ( .A(n6309), .B(n6308), .ZN(n6825) );
  INV_X1 U7981 ( .A(n6825), .ZN(n6306) );
  NAND2_X1 U7982 ( .A1(n6307), .A2(n6306), .ZN(n6826) );
  OR2_X1 U7983 ( .A1(n6309), .A2(n6308), .ZN(n6310) );
  NAND2_X1 U7984 ( .A1(n4506), .A2(n6925), .ZN(n6312) );
  NAND2_X1 U7985 ( .A1(n6496), .A2(n9096), .ZN(n6311) );
  NAND2_X1 U7986 ( .A1(n6312), .A2(n6311), .ZN(n6313) );
  XNOR2_X1 U7987 ( .A(n6313), .B(n6509), .ZN(n6317) );
  NAND2_X1 U7988 ( .A1(n6482), .A2(n9096), .ZN(n6316) );
  NAND2_X1 U7989 ( .A1(n6925), .A2(n6484), .ZN(n6315) );
  AND2_X1 U7990 ( .A1(n6316), .A2(n6315), .ZN(n7044) );
  INV_X1 U7991 ( .A(n6317), .ZN(n6318) );
  NAND2_X1 U7992 ( .A1(n6965), .A2(n4505), .ZN(n6322) );
  NAND2_X1 U7993 ( .A1(n6496), .A2(n9095), .ZN(n6321) );
  NAND2_X1 U7994 ( .A1(n6322), .A2(n6321), .ZN(n6323) );
  XNOR2_X1 U7995 ( .A(n6323), .B(n6509), .ZN(n6325) );
  AOI22_X1 U7996 ( .A1(n6965), .A2(n6496), .B1(n6482), .B2(n9095), .ZN(n6324)
         );
  NAND2_X1 U7997 ( .A1(n6325), .A2(n6324), .ZN(n6327) );
  OR2_X1 U7998 ( .A1(n6325), .A2(n6324), .ZN(n6326) );
  AND2_X1 U7999 ( .A1(n6327), .A2(n6326), .ZN(n7097) );
  NAND2_X1 U8000 ( .A1(n7100), .A2(n6327), .ZN(n7174) );
  NAND2_X1 U8001 ( .A1(n7199), .A2(n4505), .ZN(n6329) );
  NAND2_X1 U8002 ( .A1(n6496), .A2(n9094), .ZN(n6328) );
  NAND2_X1 U8003 ( .A1(n6329), .A2(n6328), .ZN(n6330) );
  XNOR2_X1 U8004 ( .A(n6330), .B(n6274), .ZN(n6345) );
  NOR2_X1 U8005 ( .A1(n6332), .A2(n6331), .ZN(n6333) );
  AOI21_X1 U8006 ( .B1(n7199), .B2(n6484), .A(n6333), .ZN(n6346) );
  XNOR2_X1 U8007 ( .A(n6345), .B(n6346), .ZN(n7175) );
  NAND2_X1 U8008 ( .A1(n7375), .A2(n4506), .ZN(n6335) );
  NAND2_X1 U8009 ( .A1(n6496), .A2(n9093), .ZN(n6334) );
  NAND2_X1 U8010 ( .A1(n6335), .A2(n6334), .ZN(n6336) );
  XNOR2_X1 U8011 ( .A(n6336), .B(n6274), .ZN(n6344) );
  NAND2_X1 U8012 ( .A1(n7375), .A2(n6496), .ZN(n6338) );
  NAND2_X1 U8013 ( .A1(n6482), .A2(n9093), .ZN(n6337) );
  NAND2_X1 U8014 ( .A1(n6338), .A2(n6337), .ZN(n7324) );
  AND2_X1 U8015 ( .A1(n6344), .A2(n7324), .ZN(n6353) );
  NAND2_X1 U8016 ( .A1(n7359), .A2(n4506), .ZN(n6340) );
  NAND2_X1 U8017 ( .A1(n6496), .A2(n9092), .ZN(n6339) );
  NAND2_X1 U8018 ( .A1(n6340), .A2(n6339), .ZN(n6341) );
  XNOR2_X1 U8019 ( .A(n6341), .B(n6274), .ZN(n6356) );
  NOR2_X1 U8020 ( .A1(n6342), .A2(n6331), .ZN(n6343) );
  AOI21_X1 U8021 ( .B1(n7359), .B2(n6496), .A(n6343), .ZN(n6354) );
  XNOR2_X1 U8022 ( .A(n6356), .B(n6354), .ZN(n7435) );
  INV_X1 U8023 ( .A(n6344), .ZN(n7433) );
  INV_X1 U8024 ( .A(n6345), .ZN(n6347) );
  NAND2_X1 U8025 ( .A1(n6347), .A2(n6346), .ZN(n7323) );
  NAND2_X1 U8026 ( .A1(n7323), .A2(n7324), .ZN(n6350) );
  INV_X1 U8027 ( .A(n7323), .ZN(n6349) );
  INV_X1 U8028 ( .A(n7324), .ZN(n6348) );
  AOI22_X1 U8029 ( .A1(n7433), .A2(n6350), .B1(n6349), .B2(n6348), .ZN(n6351)
         );
  AND2_X1 U8030 ( .A1(n7435), .A2(n6351), .ZN(n6352) );
  INV_X1 U8031 ( .A(n6354), .ZN(n6355) );
  NAND2_X1 U8032 ( .A1(n6356), .A2(n6355), .ZN(n6357) );
  NAND2_X1 U8033 ( .A1(n7524), .A2(n4506), .ZN(n6359) );
  NAND2_X1 U8034 ( .A1(n6484), .A2(n9091), .ZN(n6358) );
  NAND2_X1 U8035 ( .A1(n6359), .A2(n6358), .ZN(n6360) );
  XNOR2_X1 U8036 ( .A(n6360), .B(n6509), .ZN(n6363) );
  NAND2_X1 U8037 ( .A1(n7524), .A2(n6484), .ZN(n6362) );
  NAND2_X1 U8038 ( .A1(n6482), .A2(n9091), .ZN(n6361) );
  NAND2_X1 U8039 ( .A1(n6362), .A2(n6361), .ZN(n7464) );
  INV_X1 U8040 ( .A(n6363), .ZN(n6364) );
  NAND2_X1 U8041 ( .A1(n9723), .A2(n4505), .ZN(n6366) );
  NAND2_X1 U8042 ( .A1(n6496), .A2(n9090), .ZN(n6365) );
  NAND2_X1 U8043 ( .A1(n6366), .A2(n6365), .ZN(n6367) );
  XNOR2_X1 U8044 ( .A(n6367), .B(n6509), .ZN(n6370) );
  NOR2_X1 U8045 ( .A1(n6368), .A2(n6331), .ZN(n6369) );
  AOI21_X1 U8046 ( .B1(n9723), .B2(n6496), .A(n6369), .ZN(n6371) );
  NAND2_X1 U8047 ( .A1(n6370), .A2(n6371), .ZN(n7527) );
  INV_X1 U8048 ( .A(n6370), .ZN(n6373) );
  INV_X1 U8049 ( .A(n6371), .ZN(n6372) );
  NAND2_X1 U8050 ( .A1(n6373), .A2(n6372), .ZN(n6374) );
  NAND2_X1 U8051 ( .A1(n7527), .A2(n6374), .ZN(n7514) );
  NAND2_X1 U8052 ( .A1(n7512), .A2(n7527), .ZN(n6385) );
  NAND2_X1 U8053 ( .A1(n7620), .A2(n4505), .ZN(n6376) );
  NAND2_X1 U8054 ( .A1(n6496), .A2(n9089), .ZN(n6375) );
  NAND2_X1 U8055 ( .A1(n6376), .A2(n6375), .ZN(n6377) );
  XNOR2_X1 U8056 ( .A(n6377), .B(n6509), .ZN(n6380) );
  NOR2_X1 U8057 ( .A1(n6378), .A2(n6331), .ZN(n6379) );
  AOI21_X1 U8058 ( .B1(n7620), .B2(n6496), .A(n6379), .ZN(n6381) );
  NAND2_X1 U8059 ( .A1(n6380), .A2(n6381), .ZN(n6386) );
  INV_X1 U8060 ( .A(n6380), .ZN(n6383) );
  INV_X1 U8061 ( .A(n6381), .ZN(n6382) );
  NAND2_X1 U8062 ( .A1(n6383), .A2(n6382), .ZN(n6384) );
  AND2_X1 U8063 ( .A1(n6386), .A2(n6384), .ZN(n7528) );
  NAND2_X1 U8064 ( .A1(n6385), .A2(n7528), .ZN(n7530) );
  NAND2_X1 U8065 ( .A1(n8845), .A2(n4506), .ZN(n6388) );
  NAND2_X1 U8066 ( .A1(n6484), .A2(n9088), .ZN(n6387) );
  NAND2_X1 U8067 ( .A1(n6388), .A2(n6387), .ZN(n6389) );
  XNOR2_X1 U8068 ( .A(n6389), .B(n6274), .ZN(n6391) );
  NOR2_X1 U8069 ( .A1(n8846), .A2(n6331), .ZN(n6390) );
  AOI21_X1 U8070 ( .B1(n8845), .B2(n6496), .A(n6390), .ZN(n6392) );
  XNOR2_X1 U8071 ( .A(n6391), .B(n6392), .ZN(n7576) );
  INV_X1 U8072 ( .A(n6391), .ZN(n6393) );
  NAND2_X1 U8073 ( .A1(n6393), .A2(n6392), .ZN(n6394) );
  NAND2_X1 U8074 ( .A1(n8824), .A2(n4506), .ZN(n6396) );
  NAND2_X1 U8075 ( .A1(n6496), .A2(n9087), .ZN(n6395) );
  NAND2_X1 U8076 ( .A1(n6396), .A2(n6395), .ZN(n6397) );
  XNOR2_X1 U8077 ( .A(n6397), .B(n6509), .ZN(n6401) );
  NAND2_X1 U8078 ( .A1(n6400), .A2(n6401), .ZN(n7668) );
  NAND2_X1 U8079 ( .A1(n8824), .A2(n6484), .ZN(n6399) );
  NAND2_X1 U8080 ( .A1(n6482), .A2(n9087), .ZN(n6398) );
  NAND2_X1 U8081 ( .A1(n6399), .A2(n6398), .ZN(n7671) );
  NAND2_X1 U8082 ( .A1(n7668), .A2(n7671), .ZN(n6409) );
  INV_X1 U8083 ( .A(n6401), .ZN(n6402) );
  NAND2_X1 U8084 ( .A1(n6409), .A2(n7669), .ZN(n6407) );
  NAND2_X1 U8085 ( .A1(n8860), .A2(n4506), .ZN(n6405) );
  NAND2_X1 U8086 ( .A1(n6496), .A2(n9086), .ZN(n6404) );
  NAND2_X1 U8087 ( .A1(n6405), .A2(n6404), .ZN(n6406) );
  XNOR2_X1 U8088 ( .A(n6406), .B(n6274), .ZN(n6410) );
  NAND2_X1 U8089 ( .A1(n6407), .A2(n6410), .ZN(n7694) );
  AND2_X1 U8090 ( .A1(n6482), .A2(n9086), .ZN(n6408) );
  AOI21_X1 U8091 ( .B1(n8860), .B2(n6484), .A(n6408), .ZN(n7695) );
  NAND2_X1 U8092 ( .A1(n7694), .A2(n7695), .ZN(n7693) );
  INV_X1 U8093 ( .A(n6410), .ZN(n6411) );
  NAND2_X1 U8094 ( .A1(n9500), .A2(n4505), .ZN(n6413) );
  NAND2_X1 U8095 ( .A1(n9085), .A2(n6496), .ZN(n6412) );
  NAND2_X1 U8096 ( .A1(n6413), .A2(n6412), .ZN(n6414) );
  XNOR2_X1 U8097 ( .A(n6414), .B(n6509), .ZN(n6416) );
  AND2_X1 U8098 ( .A1(n9085), .A2(n6482), .ZN(n6415) );
  AOI21_X1 U8099 ( .B1(n9500), .B2(n6496), .A(n6415), .ZN(n6417) );
  NAND2_X1 U8100 ( .A1(n6416), .A2(n6417), .ZN(n8717) );
  INV_X1 U8101 ( .A(n6416), .ZN(n6419) );
  INV_X1 U8102 ( .A(n6417), .ZN(n6418) );
  NAND2_X1 U8103 ( .A1(n6419), .A2(n6418), .ZN(n6420) );
  AND2_X1 U8104 ( .A1(n8717), .A2(n6420), .ZN(n8708) );
  NAND2_X1 U8105 ( .A1(n9494), .A2(n4506), .ZN(n6422) );
  NAND2_X1 U8106 ( .A1(n9084), .A2(n6484), .ZN(n6421) );
  NAND2_X1 U8107 ( .A1(n6422), .A2(n6421), .ZN(n6423) );
  XNOR2_X1 U8108 ( .A(n6423), .B(n6509), .ZN(n6425) );
  AND2_X1 U8109 ( .A1(n9084), .A2(n6482), .ZN(n6424) );
  AOI21_X1 U8110 ( .B1(n9494), .B2(n6484), .A(n6424), .ZN(n6426) );
  NAND2_X1 U8111 ( .A1(n6425), .A2(n6426), .ZN(n6430) );
  INV_X1 U8112 ( .A(n6425), .ZN(n6428) );
  INV_X1 U8113 ( .A(n6426), .ZN(n6427) );
  NAND2_X1 U8114 ( .A1(n6428), .A2(n6427), .ZN(n6429) );
  AND2_X1 U8115 ( .A1(n6430), .A2(n6429), .ZN(n8718) );
  NAND2_X1 U8116 ( .A1(n8720), .A2(n6430), .ZN(n6436) );
  NAND2_X1 U8117 ( .A1(n9487), .A2(n4506), .ZN(n6432) );
  NAND2_X1 U8118 ( .A1(n9083), .A2(n6484), .ZN(n6431) );
  NAND2_X1 U8119 ( .A1(n6432), .A2(n6431), .ZN(n6433) );
  XNOR2_X1 U8120 ( .A(n6433), .B(n6509), .ZN(n6437) );
  NAND2_X1 U8121 ( .A1(n6436), .A2(n6437), .ZN(n8757) );
  NAND2_X1 U8122 ( .A1(n9487), .A2(n6496), .ZN(n6435) );
  NAND2_X1 U8123 ( .A1(n9083), .A2(n6482), .ZN(n6434) );
  NAND2_X1 U8124 ( .A1(n6435), .A2(n6434), .ZN(n8760) );
  NAND2_X1 U8125 ( .A1(n8757), .A2(n8760), .ZN(n6440) );
  NAND2_X1 U8126 ( .A1(n9481), .A2(n4505), .ZN(n6442) );
  NAND2_X1 U8127 ( .A1(n9082), .A2(n6496), .ZN(n6441) );
  NAND2_X1 U8128 ( .A1(n6442), .A2(n6441), .ZN(n6443) );
  XNOR2_X1 U8129 ( .A(n6443), .B(n6274), .ZN(n6447) );
  AND2_X1 U8130 ( .A1(n9082), .A2(n6482), .ZN(n6444) );
  AOI21_X1 U8131 ( .B1(n9481), .B2(n6496), .A(n6444), .ZN(n6445) );
  XNOR2_X1 U8132 ( .A(n6447), .B(n6445), .ZN(n8687) );
  INV_X1 U8133 ( .A(n6445), .ZN(n6446) );
  NAND2_X1 U8134 ( .A1(n6447), .A2(n6446), .ZN(n6448) );
  NAND2_X1 U8135 ( .A1(n9476), .A2(n4506), .ZN(n6450) );
  NAND2_X1 U8136 ( .A1(n9081), .A2(n6496), .ZN(n6449) );
  NAND2_X1 U8137 ( .A1(n6450), .A2(n6449), .ZN(n6451) );
  XNOR2_X1 U8138 ( .A(n6451), .B(n6509), .ZN(n6453) );
  AND2_X1 U8139 ( .A1(n9081), .A2(n6482), .ZN(n6452) );
  AOI21_X1 U8140 ( .B1(n9476), .B2(n6496), .A(n6452), .ZN(n6454) );
  NAND2_X1 U8141 ( .A1(n6453), .A2(n6454), .ZN(n8737) );
  INV_X1 U8142 ( .A(n6453), .ZN(n6456) );
  INV_X1 U8143 ( .A(n6454), .ZN(n6455) );
  NAND2_X1 U8144 ( .A1(n6456), .A2(n6455), .ZN(n8736) );
  NAND2_X1 U8145 ( .A1(n9367), .A2(n4505), .ZN(n6458) );
  NAND2_X1 U8146 ( .A1(n9080), .A2(n6496), .ZN(n6457) );
  NAND2_X1 U8147 ( .A1(n6458), .A2(n6457), .ZN(n6459) );
  XNOR2_X1 U8148 ( .A(n6459), .B(n6274), .ZN(n6463) );
  AND2_X1 U8149 ( .A1(n9080), .A2(n6482), .ZN(n6460) );
  AOI21_X1 U8150 ( .B1(n9367), .B2(n6496), .A(n6460), .ZN(n6461) );
  XNOR2_X1 U8151 ( .A(n6463), .B(n6461), .ZN(n8693) );
  INV_X1 U8152 ( .A(n6461), .ZN(n6462) );
  NAND2_X1 U8153 ( .A1(n6463), .A2(n6462), .ZN(n6464) );
  NAND2_X1 U8154 ( .A1(n9467), .A2(n6294), .ZN(n6466) );
  NAND2_X1 U8155 ( .A1(n9079), .A2(n6496), .ZN(n6465) );
  NAND2_X1 U8156 ( .A1(n6466), .A2(n6465), .ZN(n6467) );
  XNOR2_X1 U8157 ( .A(n6467), .B(n6274), .ZN(n6468) );
  AOI22_X1 U8158 ( .A1(n9467), .A2(n6496), .B1(n6482), .B2(n9079), .ZN(n8746)
         );
  NAND2_X1 U8159 ( .A1(n9459), .A2(n4505), .ZN(n6471) );
  NAND2_X1 U8160 ( .A1(n9078), .A2(n6484), .ZN(n6470) );
  NAND2_X1 U8161 ( .A1(n6471), .A2(n6470), .ZN(n6472) );
  XNOR2_X1 U8162 ( .A(n6472), .B(n6509), .ZN(n6477) );
  INV_X1 U8163 ( .A(n6477), .ZN(n6475) );
  AND2_X1 U8164 ( .A1(n9078), .A2(n6482), .ZN(n6473) );
  AOI21_X1 U8165 ( .B1(n9459), .B2(n6484), .A(n6473), .ZN(n6476) );
  INV_X1 U8166 ( .A(n6476), .ZN(n6474) );
  NAND2_X1 U8167 ( .A1(n6475), .A2(n6474), .ZN(n8677) );
  AND2_X1 U8168 ( .A1(n6477), .A2(n6476), .ZN(n8676) );
  AOI22_X1 U8169 ( .A1(n9323), .A2(n4506), .B1(n6484), .B2(n9077), .ZN(n6478)
         );
  XNOR2_X1 U8170 ( .A(n6478), .B(n6274), .ZN(n6480) );
  AOI22_X1 U8171 ( .A1(n9323), .A2(n6496), .B1(n6482), .B2(n9077), .ZN(n6479)
         );
  NAND2_X1 U8172 ( .A1(n6480), .A2(n6479), .ZN(n6481) );
  OAI21_X1 U8173 ( .B1(n6480), .B2(n6479), .A(n6481), .ZN(n8729) );
  AOI22_X1 U8174 ( .A1(n6483), .A2(n6496), .B1(n6482), .B2(n9076), .ZN(n6492)
         );
  NAND2_X1 U8175 ( .A1(n6483), .A2(n4505), .ZN(n6486) );
  NAND2_X1 U8176 ( .A1(n6484), .A2(n9076), .ZN(n6485) );
  NAND2_X1 U8177 ( .A1(n6486), .A2(n6485), .ZN(n6487) );
  XNOR2_X1 U8178 ( .A(n6487), .B(n6274), .ZN(n6494) );
  XOR2_X1 U8179 ( .A(n6492), .B(n6494), .Z(n8701) );
  NAND2_X1 U8180 ( .A1(n9446), .A2(n4506), .ZN(n6489) );
  NAND2_X1 U8181 ( .A1(n6496), .A2(n9075), .ZN(n6488) );
  NAND2_X1 U8182 ( .A1(n6489), .A2(n6488), .ZN(n6490) );
  XNOR2_X1 U8183 ( .A(n6490), .B(n6509), .ZN(n6504) );
  NOR2_X1 U8184 ( .A1(n8895), .A2(n6331), .ZN(n6491) );
  AOI21_X1 U8185 ( .B1(n9446), .B2(n6496), .A(n6491), .ZN(n6505) );
  XNOR2_X1 U8186 ( .A(n6504), .B(n6505), .ZN(n8771) );
  INV_X1 U8187 ( .A(n6492), .ZN(n6493) );
  NAND2_X1 U8188 ( .A1(n9269), .A2(n6294), .ZN(n6498) );
  NAND2_X1 U8189 ( .A1(n6496), .A2(n9074), .ZN(n6497) );
  NAND2_X1 U8190 ( .A1(n6498), .A2(n6497), .ZN(n6499) );
  XNOR2_X1 U8191 ( .A(n6499), .B(n6509), .ZN(n6503) );
  NOR2_X1 U8192 ( .A1(n6500), .A2(n6331), .ZN(n6501) );
  AOI21_X1 U8193 ( .B1(n9269), .B2(n6496), .A(n6501), .ZN(n6502) );
  NAND2_X1 U8194 ( .A1(n6503), .A2(n6502), .ZN(n6535) );
  OAI21_X1 U8195 ( .B1(n6503), .B2(n6502), .A(n6535), .ZN(n7775) );
  INV_X1 U8196 ( .A(n6504), .ZN(n6507) );
  INV_X1 U8197 ( .A(n6505), .ZN(n6506) );
  INV_X1 U8198 ( .A(n7774), .ZN(n6521) );
  OAI22_X1 U8199 ( .A1(n9260), .A2(n6266), .B1(n6543), .B2(n6331), .ZN(n6510)
         );
  XNOR2_X1 U8200 ( .A(n6510), .B(n6509), .ZN(n6512) );
  OAI22_X1 U8201 ( .A1(n9260), .A2(n6320), .B1(n6543), .B2(n6266), .ZN(n6511)
         );
  XNOR2_X1 U8202 ( .A(n6512), .B(n6511), .ZN(n6522) );
  INV_X1 U8203 ( .A(n6522), .ZN(n6536) );
  NAND2_X1 U8204 ( .A1(n6527), .A2(n9749), .ZN(n9747) );
  NAND2_X1 U8205 ( .A1(n6513), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U8206 ( .A1(n6515), .A2(n6514), .ZN(n6516) );
  INV_X1 U8207 ( .A(n7028), .ZN(n6517) );
  OR2_X1 U8208 ( .A1(n9747), .A2(n6517), .ZN(n6526) );
  INV_X1 U8209 ( .A(n6526), .ZN(n6520) );
  INV_X1 U8210 ( .A(n9499), .ZN(n9779) );
  INV_X1 U8211 ( .A(n9001), .ZN(n6518) );
  AND2_X1 U8212 ( .A1(n9779), .A2(n6518), .ZN(n6519) );
  NAND2_X1 U8213 ( .A1(n6520), .A2(n6519), .ZN(n8769) );
  NAND2_X1 U8214 ( .A1(n6521), .A2(n5061), .ZN(n6542) );
  AND2_X1 U8215 ( .A1(n6522), .A2(n8775), .ZN(n6523) );
  NAND2_X1 U8216 ( .A1(n7774), .A2(n6523), .ZN(n6541) );
  OR2_X1 U8217 ( .A1(n6524), .A2(n7416), .ZN(n7030) );
  OAI21_X2 U8218 ( .B1(n6526), .B2(n7030), .A(n9405), .ZN(n8767) );
  INV_X1 U8219 ( .A(n9258), .ZN(n6534) );
  NAND2_X1 U8220 ( .A1(n6527), .A2(n7028), .ZN(n6529) );
  NAND2_X1 U8221 ( .A1(n9499), .A2(n7030), .ZN(n6528) );
  NAND2_X1 U8222 ( .A1(n6529), .A2(n6528), .ZN(n6530) );
  AND3_X1 U8223 ( .A1(n6261), .A2(n6566), .A3(n7612), .ZN(n9067) );
  NAND2_X1 U8224 ( .A1(n6530), .A2(n9067), .ZN(n6646) );
  NAND2_X1 U8225 ( .A1(n6646), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8765) );
  NAND2_X1 U8226 ( .A1(n7028), .A2(n6256), .ZN(n6531) );
  NOR2_X1 U8227 ( .A1(n9747), .A2(n6531), .ZN(n8763) );
  AOI22_X1 U8228 ( .A1(n8763), .A2(n6532), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6533) );
  OAI21_X1 U8229 ( .B1(n6534), .B2(n8765), .A(n6533), .ZN(n6538) );
  NOR3_X1 U8230 ( .A1(n6536), .A2(n6535), .A3(n8769), .ZN(n6537) );
  AOI211_X1 U8231 ( .C1(n6539), .C2(n8767), .A(n6538), .B(n6537), .ZN(n6540)
         );
  NAND3_X1 U8232 ( .A1(n6542), .A2(n6541), .A3(n6540), .ZN(P1_U3220) );
  NAND2_X1 U8233 ( .A1(n6539), .A2(n9073), .ZN(n6544) );
  NAND2_X1 U8234 ( .A1(n8906), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U8235 ( .A1(n7760), .A2(n7714), .ZN(n6565) );
  INV_X1 U8236 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6561) );
  NAND2_X1 U8237 ( .A1(n6553), .A2(n6552), .ZN(n8986) );
  INV_X1 U8238 ( .A(n8986), .ZN(n8898) );
  NAND2_X1 U8239 ( .A1(n5201), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6557) );
  NAND2_X1 U8240 ( .A1(n6554), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U8241 ( .A1(n5200), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6555) );
  AND3_X1 U8242 ( .A1(n6557), .A2(n6556), .A3(n6555), .ZN(n8925) );
  INV_X1 U8243 ( .A(n8925), .ZN(n9071) );
  INV_X1 U8244 ( .A(n7722), .ZN(n9110) );
  NAND2_X1 U8245 ( .A1(n9110), .A2(P1_B_REG_SCAN_IN), .ZN(n6558) );
  AND2_X1 U8246 ( .A1(n8777), .A2(n6558), .ZN(n9242) );
  AOI22_X1 U8247 ( .A1(n9071), .A2(n9242), .B1(n9066), .B2(n9073), .ZN(n6559)
         );
  OAI21_X1 U8248 ( .B1(n6560), .B2(n9752), .A(n6559), .ZN(n7763) );
  NOR2_X1 U8249 ( .A1(n7768), .A2(n7763), .ZN(n6571) );
  MUX2_X1 U8250 ( .A(n6561), .B(n6571), .S(n9788), .Z(n6564) );
  NAND2_X1 U8251 ( .A1(n9788), .A2(n9499), .ZN(n9543) );
  NAND2_X1 U8252 ( .A1(n6551), .A2(n6562), .ZN(n6563) );
  NAND2_X1 U8253 ( .A1(n6565), .A2(n5067), .ZN(P1_U3519) );
  INV_X1 U8254 ( .A(n6566), .ZN(n6567) );
  NOR2_X1 U8255 ( .A1(n6568), .A2(n6567), .ZN(n6570) );
  INV_X1 U8256 ( .A(n9747), .ZN(n6569) );
  AND2_X2 U8257 ( .A1(n6570), .A2(n6569), .ZN(n9797) );
  NAND2_X1 U8258 ( .A1(n7760), .A2(n7727), .ZN(n6575) );
  INV_X1 U8259 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n10270) );
  MUX2_X1 U8260 ( .A(n10270), .B(n6571), .S(n9797), .Z(n6574) );
  NAND2_X1 U8261 ( .A1(n9797), .A2(n9499), .ZN(n9469) );
  NAND2_X1 U8262 ( .A1(n6551), .A2(n6572), .ZN(n6573) );
  NAND2_X1 U8263 ( .A1(n6575), .A2(n5066), .ZN(P1_U3551) );
  INV_X1 U8264 ( .A(n6606), .ZN(n6576) );
  OR2_X2 U8265 ( .A1(n6864), .A2(n6576), .ZN(n8297) );
  NAND2_X1 U8266 ( .A1(n7947), .A2(n6864), .ZN(n6577) );
  NAND2_X1 U8267 ( .A1(n6577), .A2(n6871), .ZN(n6758) );
  NAND2_X1 U8268 ( .A1(n6758), .A2(n5780), .ZN(n6578) );
  NAND2_X1 U8269 ( .A1(n6578), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8270 ( .A(n6261), .ZN(n6580) );
  AND2_X2 U8271 ( .A1(n6580), .A2(n6579), .ZN(P1_U3973) );
  INV_X1 U8272 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6581) );
  NOR2_X1 U8273 ( .A1(n4610), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8673) );
  INV_X2 U8274 ( .A(n8673), .ZN(n8668) );
  OAI222_X1 U8275 ( .A1(P2_U3151), .A2(n6854), .B1(n6582), .B2(n6586), .C1(
        n6581), .C2(n8668), .ZN(P2_U3294) );
  INV_X1 U8276 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6583) );
  INV_X1 U8277 ( .A(n7008), .ZN(n6988) );
  OAI222_X1 U8278 ( .A1(n8668), .A2(n6583), .B1(n6582), .B2(n6589), .C1(n6988), 
        .C2(P2_U3151), .ZN(P2_U3293) );
  NAND2_X1 U8279 ( .A1(n4610), .A2(P1_U3086), .ZN(n9569) );
  INV_X1 U8280 ( .A(n9569), .ZN(n9563) );
  AOI22_X1 U8281 ( .A1(n9563), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n9105), .ZN(n6585) );
  OAI21_X1 U8282 ( .B1(n6586), .B2(n9572), .A(n6585), .ZN(P1_U3354) );
  OAI222_X1 U8283 ( .A1(n9798), .A2(P2_U3151), .B1(n6582), .B2(n6591), .C1(
        n6587), .C2(n8668), .ZN(P2_U3292) );
  AOI22_X1 U8284 ( .A1(n9563), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n9118), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6588) );
  OAI21_X1 U8285 ( .B1(n6589), .B2(n9572), .A(n6588), .ZN(P1_U3353) );
  AOI22_X1 U8286 ( .A1(n9131), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n9563), .ZN(n6590) );
  OAI21_X1 U8287 ( .B1(n6591), .B2(n9572), .A(n6590), .ZN(P1_U3352) );
  INV_X1 U8288 ( .A(n6592), .ZN(n6596) );
  AOI22_X1 U8289 ( .A1(n9143), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n9563), .ZN(n6593) );
  OAI21_X1 U8290 ( .B1(n6596), .B2(n9572), .A(n6593), .ZN(P1_U3351) );
  AOI22_X1 U8291 ( .A1(n9156), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9563), .ZN(n6594) );
  OAI21_X1 U8292 ( .B1(n6598), .B2(n9572), .A(n6594), .ZN(P1_U3350) );
  INV_X1 U8293 ( .A(n7015), .ZN(n9827) );
  INV_X1 U8294 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6595) );
  OAI222_X1 U8295 ( .A1(n9827), .A2(P2_U3151), .B1(n6582), .B2(n6596), .C1(
        n6595), .C2(n8668), .ZN(P2_U3291) );
  OAI222_X1 U8296 ( .A1(n10156), .A2(P2_U3151), .B1(n6582), .B2(n6598), .C1(
        n6597), .C2(n8668), .ZN(P2_U3290) );
  INV_X1 U8297 ( .A(n6599), .ZN(n6609) );
  AOI22_X1 U8298 ( .A1(n9169), .A2(P1_STATE_REG_SCAN_IN), .B1(n9563), .B2(
        P2_DATAO_REG_6__SCAN_IN), .ZN(n6600) );
  OAI21_X1 U8299 ( .B1(n6609), .B2(n9572), .A(n6600), .ZN(P1_U3349) );
  INV_X1 U8300 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6602) );
  NAND2_X1 U8301 ( .A1(n7069), .A2(n6883), .ZN(n6601) );
  OAI21_X1 U8302 ( .B1(n6883), .B2(n6602), .A(n6601), .ZN(P2_U3377) );
  NAND2_X1 U8303 ( .A1(n6883), .A2(n6603), .ZN(n6621) );
  INV_X1 U8304 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6607) );
  INV_X1 U8305 ( .A(n6604), .ZN(n6605) );
  AOI22_X1 U8306 ( .A1(n6621), .A2(n6607), .B1(n6606), .B2(n6605), .ZN(
        P2_U3376) );
  INV_X1 U8307 ( .A(n8309), .ZN(n8277) );
  INV_X1 U8308 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6608) );
  OAI222_X1 U8309 ( .A1(n8277), .A2(P2_U3151), .B1(n6582), .B2(n6609), .C1(
        n6608), .C2(n8668), .ZN(P2_U3289) );
  INV_X1 U8310 ( .A(n7612), .ZN(n6610) );
  OR2_X1 U8311 ( .A1(n6261), .A2(n6610), .ZN(n6611) );
  AND2_X1 U8312 ( .A1(n6611), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6649) );
  NAND2_X1 U8313 ( .A1(n9001), .A2(n7612), .ZN(n6613) );
  NAND2_X1 U8314 ( .A1(n6613), .A2(n6612), .ZN(n6650) );
  AND2_X1 U8315 ( .A1(n6649), .A2(n6650), .ZN(n9670) );
  NOR2_X1 U8316 ( .A1(n9670), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8317 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6615) );
  INV_X1 U8318 ( .A(n6614), .ZN(n6617) );
  INV_X1 U8319 ( .A(n6696), .ZN(n9187) );
  OAI222_X1 U8320 ( .A1(n9569), .A2(n6615), .B1(n9572), .B2(n6617), .C1(
        P1_U3086), .C2(n9187), .ZN(P1_U3348) );
  INV_X1 U8321 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6616) );
  OAI222_X1 U8322 ( .A1(n8310), .A2(P2_U3151), .B1(n6582), .B2(n6617), .C1(
        n6616), .C2(n8668), .ZN(P2_U3288) );
  INV_X1 U8323 ( .A(n6618), .ZN(n6620) );
  AOI22_X1 U8324 ( .A1(n9199), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9563), .ZN(n6619) );
  OAI21_X1 U8325 ( .B1(n6620), .B2(n9572), .A(n6619), .ZN(P1_U3347) );
  OAI222_X1 U8326 ( .A1(n8306), .A2(P2_U3151), .B1(n6582), .B2(n6620), .C1(
        n10288), .C2(n8668), .ZN(P2_U3287) );
  INV_X1 U8327 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10404) );
  NOR2_X1 U8328 ( .A1(n6731), .A2(n10404), .ZN(P2_U3250) );
  INV_X1 U8329 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n6622) );
  NOR2_X1 U8330 ( .A1(n6731), .A2(n6622), .ZN(P2_U3251) );
  INV_X1 U8331 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n10287) );
  NOR2_X1 U8332 ( .A1(n6731), .A2(n10287), .ZN(P2_U3247) );
  INV_X1 U8333 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n6623) );
  NOR2_X1 U8334 ( .A1(n6731), .A2(n6623), .ZN(P2_U3254) );
  INV_X1 U8335 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n6624) );
  NOR2_X1 U8336 ( .A1(n6731), .A2(n6624), .ZN(P2_U3256) );
  INV_X1 U8337 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n6625) );
  NOR2_X1 U8338 ( .A1(n6731), .A2(n6625), .ZN(P2_U3257) );
  INV_X1 U8339 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n6626) );
  NOR2_X1 U8340 ( .A1(n6731), .A2(n6626), .ZN(P2_U3249) );
  INV_X1 U8341 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n6627) );
  NOR2_X1 U8342 ( .A1(n6731), .A2(n6627), .ZN(P2_U3253) );
  INV_X1 U8343 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n6628) );
  NOR2_X1 U8344 ( .A1(n6731), .A2(n6628), .ZN(P2_U3248) );
  INV_X1 U8345 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n6629) );
  NOR2_X1 U8346 ( .A1(n6731), .A2(n6629), .ZN(P2_U3246) );
  INV_X1 U8347 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n6630) );
  NOR2_X1 U8348 ( .A1(n6731), .A2(n6630), .ZN(P2_U3252) );
  INV_X1 U8349 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n6631) );
  NOR2_X1 U8350 ( .A1(n6731), .A2(n6631), .ZN(P2_U3255) );
  NAND2_X1 U8351 ( .A1(n9749), .A2(n6632), .ZN(n9746) );
  INV_X1 U8352 ( .A(n9746), .ZN(n9745) );
  OAI21_X1 U8353 ( .B1(n9745), .B2(P1_D_REG_1__SCAN_IN), .A(n6633), .ZN(n6634)
         );
  OAI21_X1 U8354 ( .B1(n9749), .B2(n6635), .A(n6634), .ZN(P1_U3440) );
  INV_X1 U8355 ( .A(n6636), .ZN(n6638) );
  AOI22_X1 U8356 ( .A1(n6719), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9563), .ZN(n6637) );
  OAI21_X1 U8357 ( .B1(n6638), .B2(n9572), .A(n6637), .ZN(P1_U3346) );
  INV_X1 U8358 ( .A(n9872), .ZN(n8314) );
  OAI222_X1 U8359 ( .A1(n8668), .A2(n6639), .B1(n6582), .B2(n6638), .C1(
        P2_U3151), .C2(n8314), .ZN(P2_U3286) );
  INV_X1 U8360 ( .A(n6640), .ZN(n6643) );
  INV_X1 U8361 ( .A(n6723), .ZN(n9584) );
  OAI222_X1 U8362 ( .A1(n9572), .A2(n6643), .B1(n9584), .B2(P1_U3086), .C1(
        n6641), .C2(n9569), .ZN(P1_U3345) );
  OAI222_X1 U8363 ( .A1(P2_U3151), .A2(n8305), .B1(n6582), .B2(n6643), .C1(
        n6642), .C2(n8668), .ZN(P2_U3285) );
  XNOR2_X1 U8364 ( .A(n6645), .B(n6644), .ZN(n9111) );
  OR2_X1 U8365 ( .A1(n6646), .A2(P1_U3086), .ZN(n6771) );
  AND2_X1 U8366 ( .A1(n6276), .A2(n8777), .ZN(n9754) );
  AOI22_X1 U8367 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n6771), .B1(n8763), .B2(
        n9754), .ZN(n6648) );
  NAND2_X1 U8368 ( .A1(n8767), .A2(n9755), .ZN(n6647) );
  OAI211_X1 U8369 ( .C1(n9111), .C2(n8769), .A(n6648), .B(n6647), .ZN(P1_U3232) );
  INV_X1 U8370 ( .A(n6649), .ZN(n6651) );
  OR2_X1 U8371 ( .A1(n6651), .A2(n6650), .ZN(n6681) );
  NOR2_X1 U8372 ( .A1(n7722), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6652) );
  NOR2_X1 U8373 ( .A1(n5675), .A2(n6652), .ZN(n9114) );
  OAI21_X1 U8374 ( .B1(n9110), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9114), .ZN(
        n6653) );
  MUX2_X1 U8375 ( .A(n6653), .B(n9114), .S(P1_IR_REG_0__SCAN_IN), .Z(n6655) );
  INV_X1 U8376 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6654) );
  OAI22_X1 U8377 ( .A1(n6681), .A2(n6655), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6654), .ZN(n6658) );
  INV_X1 U8378 ( .A(n6681), .ZN(n6683) );
  NAND2_X1 U8379 ( .A1(n6683), .A2(n7722), .ZN(n9649) );
  NOR3_X1 U8380 ( .A1(n9649), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n6656), .ZN(
        n6657) );
  AOI211_X1 U8381 ( .C1(n9670), .C2(P1_ADDR_REG_0__SCAN_IN), .A(n6658), .B(
        n6657), .ZN(n6659) );
  INV_X1 U8382 ( .A(n6659), .ZN(P1_U3243) );
  INV_X1 U8383 ( .A(n6660), .ZN(n6706) );
  AOI22_X1 U8384 ( .A1(n9607), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9563), .ZN(n6661) );
  OAI21_X1 U8385 ( .B1(n6706), .B2(n9572), .A(n6661), .ZN(P1_U3344) );
  XNOR2_X1 U8386 ( .A(n6719), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n6680) );
  INV_X1 U8387 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6662) );
  MUX2_X1 U8388 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6662), .S(n9118), .Z(n9121)
         );
  XNOR2_X1 U8389 ( .A(n9105), .B(n6663), .ZN(n9101) );
  AND2_X1 U8390 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9100) );
  NAND2_X1 U8391 ( .A1(n9101), .A2(n9100), .ZN(n9099) );
  NAND2_X1 U8392 ( .A1(n9105), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6664) );
  NAND2_X1 U8393 ( .A1(n9099), .A2(n6664), .ZN(n9120) );
  NAND2_X1 U8394 ( .A1(n9121), .A2(n9120), .ZN(n9119) );
  NAND2_X1 U8395 ( .A1(n9118), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6665) );
  NAND2_X1 U8396 ( .A1(n9119), .A2(n6665), .ZN(n9133) );
  INV_X1 U8397 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6666) );
  XNOR2_X1 U8398 ( .A(n9131), .B(n6666), .ZN(n9134) );
  NAND2_X1 U8399 ( .A1(n9133), .A2(n9134), .ZN(n9132) );
  NAND2_X1 U8400 ( .A1(n9131), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6667) );
  NAND2_X1 U8401 ( .A1(n9132), .A2(n6667), .ZN(n9145) );
  INV_X1 U8402 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6668) );
  XNOR2_X1 U8403 ( .A(n9143), .B(n6668), .ZN(n9146) );
  NAND2_X1 U8404 ( .A1(n9145), .A2(n9146), .ZN(n9144) );
  NAND2_X1 U8405 ( .A1(n9143), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U8406 ( .A1(n9144), .A2(n6669), .ZN(n9158) );
  INV_X1 U8407 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6670) );
  MUX2_X1 U8408 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6670), .S(n9156), .Z(n9159)
         );
  NAND2_X1 U8409 ( .A1(n9158), .A2(n9159), .ZN(n9157) );
  NAND2_X1 U8410 ( .A1(n9156), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6671) );
  NAND2_X1 U8411 ( .A1(n9157), .A2(n6671), .ZN(n9171) );
  INV_X1 U8412 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6672) );
  MUX2_X1 U8413 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6672), .S(n9169), .Z(n9172)
         );
  NAND2_X1 U8414 ( .A1(n9171), .A2(n9172), .ZN(n9170) );
  NAND2_X1 U8415 ( .A1(n9169), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U8416 ( .A1(n9170), .A2(n6673), .ZN(n9180) );
  INV_X1 U8417 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6674) );
  MUX2_X1 U8418 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n6674), .S(n6696), .Z(n9181)
         );
  NAND2_X1 U8419 ( .A1(n9180), .A2(n9181), .ZN(n9179) );
  NAND2_X1 U8420 ( .A1(n6696), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6675) );
  NAND2_X1 U8421 ( .A1(n9179), .A2(n6675), .ZN(n9193) );
  INV_X1 U8422 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6676) );
  MUX2_X1 U8423 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n6676), .S(n9199), .Z(n9194)
         );
  NAND2_X1 U8424 ( .A1(n9193), .A2(n9194), .ZN(n9192) );
  NAND2_X1 U8425 ( .A1(n9199), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6677) );
  NAND2_X1 U8426 ( .A1(n9192), .A2(n6677), .ZN(n6679) );
  INV_X1 U8427 ( .A(n6709), .ZN(n6678) );
  AOI21_X1 U8428 ( .B1(n6680), .B2(n6679), .A(n6678), .ZN(n6705) );
  NOR2_X1 U8429 ( .A1(n6681), .A2(n7722), .ZN(n9231) );
  NAND2_X1 U8430 ( .A1(n9231), .A2(n6682), .ZN(n9665) );
  NAND2_X1 U8431 ( .A1(n6683), .A2(n5675), .ZN(n9704) );
  INV_X1 U8432 ( .A(n9704), .ZN(n9673) );
  INV_X1 U8433 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6686) );
  NOR2_X1 U8434 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6684), .ZN(n7440) );
  INV_X1 U8435 ( .A(n7440), .ZN(n6685) );
  OAI21_X1 U8436 ( .B1(n9708), .B2(n6686), .A(n6685), .ZN(n6703) );
  INV_X1 U8437 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9791) );
  MUX2_X1 U8438 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9791), .S(n9118), .Z(n9124)
         );
  INV_X1 U8439 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6687) );
  XNOR2_X1 U8440 ( .A(n9105), .B(n6687), .ZN(n9104) );
  AND2_X1 U8441 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9103) );
  NAND2_X1 U8442 ( .A1(n9104), .A2(n9103), .ZN(n9102) );
  NAND2_X1 U8443 ( .A1(n9105), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6688) );
  NAND2_X1 U8444 ( .A1(n9102), .A2(n6688), .ZN(n9123) );
  NAND2_X1 U8445 ( .A1(n9124), .A2(n9123), .ZN(n9122) );
  NAND2_X1 U8446 ( .A1(n9118), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6689) );
  NAND2_X1 U8447 ( .A1(n9122), .A2(n6689), .ZN(n9136) );
  INV_X1 U8448 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6690) );
  XNOR2_X1 U8449 ( .A(n9131), .B(n6690), .ZN(n9137) );
  NAND2_X1 U8450 ( .A1(n9136), .A2(n9137), .ZN(n9135) );
  NAND2_X1 U8451 ( .A1(n9131), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6691) );
  NAND2_X1 U8452 ( .A1(n9135), .A2(n6691), .ZN(n9148) );
  INV_X1 U8453 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6692) );
  XNOR2_X1 U8454 ( .A(n9143), .B(n6692), .ZN(n9149) );
  NAND2_X1 U8455 ( .A1(n9148), .A2(n9149), .ZN(n9147) );
  NAND2_X1 U8456 ( .A1(n9143), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6693) );
  NAND2_X1 U8457 ( .A1(n9147), .A2(n6693), .ZN(n9161) );
  INV_X1 U8458 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10360) );
  MUX2_X1 U8459 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10360), .S(n9156), .Z(n9162)
         );
  NAND2_X1 U8460 ( .A1(n9161), .A2(n9162), .ZN(n9160) );
  NAND2_X1 U8461 ( .A1(n9156), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6694) );
  NAND2_X1 U8462 ( .A1(n9160), .A2(n6694), .ZN(n9174) );
  INV_X1 U8463 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6966) );
  MUX2_X1 U8464 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6966), .S(n9169), .Z(n9175)
         );
  NAND2_X1 U8465 ( .A1(n9174), .A2(n9175), .ZN(n9173) );
  NAND2_X1 U8466 ( .A1(n9169), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6695) );
  NAND2_X1 U8467 ( .A1(n9173), .A2(n6695), .ZN(n9185) );
  INV_X1 U8468 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9793) );
  MUX2_X1 U8469 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9793), .S(n6696), .Z(n9186)
         );
  NAND2_X1 U8470 ( .A1(n9185), .A2(n9186), .ZN(n9184) );
  NAND2_X1 U8471 ( .A1(n6696), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6697) );
  NAND2_X1 U8472 ( .A1(n9184), .A2(n6697), .ZN(n9197) );
  INV_X1 U8473 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10343) );
  MUX2_X1 U8474 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10343), .S(n9199), .Z(n9198)
         );
  NAND2_X1 U8475 ( .A1(n9197), .A2(n9198), .ZN(n9196) );
  NAND2_X1 U8476 ( .A1(n9199), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6698) );
  NAND2_X1 U8477 ( .A1(n9196), .A2(n6698), .ZN(n6700) );
  XNOR2_X1 U8478 ( .A(n6719), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U8479 ( .A1(n6700), .A2(n6699), .ZN(n6701) );
  AOI21_X1 U8480 ( .B1(n6721), .B2(n6701), .A(n9649), .ZN(n6702) );
  AOI211_X1 U8481 ( .C1(n9673), .C2(n6719), .A(n6703), .B(n6702), .ZN(n6704)
         );
  OAI21_X1 U8482 ( .B1(n6705), .B2(n9665), .A(n6704), .ZN(P1_U3252) );
  INV_X1 U8483 ( .A(n9904), .ZN(n8318) );
  OAI222_X1 U8484 ( .A1(n8318), .A2(P2_U3151), .B1(n6582), .B2(n6706), .C1(
        n10453), .C2(n8668), .ZN(P2_U3284) );
  NOR2_X1 U8485 ( .A1(n9216), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6707) );
  AOI21_X1 U8486 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9216), .A(n6707), .ZN(
        n6715) );
  OR2_X1 U8487 ( .A1(n6719), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U8488 ( .A1(n6709), .A2(n6708), .ZN(n9575) );
  INV_X1 U8489 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6710) );
  MUX2_X1 U8490 ( .A(n6710), .B(P1_REG2_REG_10__SCAN_IN), .S(n6723), .Z(n9574)
         );
  NAND2_X1 U8491 ( .A1(n6723), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6711) );
  OR2_X1 U8492 ( .A1(n9607), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6713) );
  NAND2_X1 U8493 ( .A1(n9607), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6712) );
  NAND2_X1 U8494 ( .A1(n6713), .A2(n6712), .ZN(n9608) );
  NOR2_X1 U8495 ( .A1(n9609), .A2(n9608), .ZN(n9610) );
  AOI21_X1 U8496 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9607), .A(n9610), .ZN(
        n6714) );
  NAND2_X1 U8497 ( .A1(n6715), .A2(n6714), .ZN(n9205) );
  OAI21_X1 U8498 ( .B1(n6715), .B2(n6714), .A(n9205), .ZN(n6718) );
  INV_X1 U8499 ( .A(n9665), .ZN(n9692) );
  INV_X1 U8500 ( .A(n9216), .ZN(n6778) );
  NAND2_X1 U8501 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7533) );
  NAND2_X1 U8502 ( .A1(n9670), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6716) );
  OAI211_X1 U8503 ( .C1(n9704), .C2(n6778), .A(n7533), .B(n6716), .ZN(n6717)
         );
  AOI21_X1 U8504 ( .B1(n6718), .B2(n9692), .A(n6717), .ZN(n6730) );
  OR2_X1 U8505 ( .A1(n6719), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6720) );
  NAND2_X1 U8506 ( .A1(n6721), .A2(n6720), .ZN(n9579) );
  INV_X1 U8507 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6722) );
  MUX2_X1 U8508 ( .A(n6722), .B(P1_REG1_REG_10__SCAN_IN), .S(n6723), .Z(n9578)
         );
  NAND2_X1 U8509 ( .A1(n6723), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6724) );
  INV_X1 U8510 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6725) );
  MUX2_X1 U8511 ( .A(n6725), .B(P1_REG1_REG_11__SCAN_IN), .S(n9607), .Z(n9613)
         );
  NOR2_X1 U8512 ( .A1(n9614), .A2(n9613), .ZN(n9615) );
  AOI21_X1 U8513 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9607), .A(n9615), .ZN(
        n6727) );
  INV_X1 U8514 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U8515 ( .A1(n9216), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n10319), .B2(
        n6778), .ZN(n6726) );
  NAND2_X1 U8516 ( .A1(n6727), .A2(n6726), .ZN(n9215) );
  OAI21_X1 U8517 ( .B1(n6727), .B2(n6726), .A(n9215), .ZN(n6728) );
  NAND2_X1 U8518 ( .A1(n6728), .A2(n9699), .ZN(n6729) );
  NAND2_X1 U8519 ( .A1(n6730), .A2(n6729), .ZN(P1_U3255) );
  INV_X1 U8520 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n6732) );
  NOR2_X1 U8521 ( .A1(n6731), .A2(n6732), .ZN(P2_U3234) );
  INV_X1 U8522 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n6733) );
  NOR2_X1 U8523 ( .A1(n6731), .A2(n6733), .ZN(P2_U3263) );
  INV_X1 U8524 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n6734) );
  NOR2_X1 U8525 ( .A1(n6731), .A2(n6734), .ZN(P2_U3262) );
  INV_X1 U8526 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n6735) );
  NOR2_X1 U8527 ( .A1(n6731), .A2(n6735), .ZN(P2_U3258) );
  INV_X1 U8528 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n6736) );
  NOR2_X1 U8529 ( .A1(n6731), .A2(n6736), .ZN(P2_U3260) );
  INV_X1 U8530 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n6737) );
  NOR2_X1 U8531 ( .A1(n6731), .A2(n6737), .ZN(P2_U3259) );
  INV_X1 U8532 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10435) );
  NOR2_X1 U8533 ( .A1(n6731), .A2(n10435), .ZN(P2_U3245) );
  INV_X1 U8534 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n6738) );
  NOR2_X1 U8535 ( .A1(n6731), .A2(n6738), .ZN(P2_U3243) );
  INV_X1 U8536 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n6739) );
  NOR2_X1 U8537 ( .A1(n6731), .A2(n6739), .ZN(P2_U3242) );
  INV_X1 U8538 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n6740) );
  NOR2_X1 U8539 ( .A1(n6731), .A2(n6740), .ZN(P2_U3241) );
  INV_X1 U8540 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n6741) );
  NOR2_X1 U8541 ( .A1(n6731), .A2(n6741), .ZN(P2_U3240) );
  INV_X1 U8542 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10389) );
  NOR2_X1 U8543 ( .A1(n6731), .A2(n10389), .ZN(P2_U3239) );
  INV_X1 U8544 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n6742) );
  NOR2_X1 U8545 ( .A1(n6731), .A2(n6742), .ZN(P2_U3238) );
  INV_X1 U8546 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n6743) );
  NOR2_X1 U8547 ( .A1(n6731), .A2(n6743), .ZN(P2_U3237) );
  INV_X1 U8548 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n6744) );
  NOR2_X1 U8549 ( .A1(n6731), .A2(n6744), .ZN(P2_U3236) );
  INV_X1 U8550 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n6745) );
  NOR2_X1 U8551 ( .A1(n6731), .A2(n6745), .ZN(P2_U3235) );
  INV_X1 U8552 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n10373) );
  NOR2_X1 U8553 ( .A1(n6731), .A2(n10373), .ZN(P2_U3261) );
  INV_X1 U8554 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10369) );
  NOR2_X1 U8555 ( .A1(n6731), .A2(n10369), .ZN(P2_U3244) );
  NAND2_X1 U8556 ( .A1(n6748), .A2(n6747), .ZN(n6749) );
  XNOR2_X1 U8557 ( .A(n6746), .B(n6749), .ZN(n6750) );
  NAND2_X1 U8558 ( .A1(n6750), .A2(n8775), .ZN(n6754) );
  INV_X1 U8559 ( .A(n6265), .ZN(n6751) );
  OAI22_X1 U8560 ( .A1(n6752), .A2(n7750), .B1(n6751), .B2(n7748), .ZN(n7149)
         );
  AOI22_X1 U8561 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(n6771), .B1(n8763), .B2(
        n7149), .ZN(n6753) );
  OAI211_X1 U8562 ( .C1(n5190), .C2(n8785), .A(n6754), .B(n6753), .ZN(P1_U3222) );
  NOR2_X1 U8563 ( .A1(n8291), .A2(P2_U3151), .ZN(n7724) );
  NAND2_X1 U8564 ( .A1(n6758), .A2(n7724), .ZN(n6755) );
  MUX2_X1 U8565 ( .A(n8297), .B(n6755), .S(n7989), .Z(n10157) );
  INV_X1 U8566 ( .A(n6871), .ZN(n6756) );
  NOR2_X1 U8567 ( .A1(n6864), .A2(n6756), .ZN(n6757) );
  OR2_X1 U8568 ( .A1(P2_U3150), .A2(n6757), .ZN(n9837) );
  NOR2_X1 U8569 ( .A1(n7989), .A2(P2_U3151), .ZN(n8672) );
  AND2_X1 U8570 ( .A1(n6758), .A2(n8672), .ZN(n6787) );
  OR2_X1 U8571 ( .A1(n8297), .A2(n6759), .ZN(n10140) );
  NOR2_X1 U8572 ( .A1(n6787), .A2(n10010), .ZN(n6762) );
  NOR2_X1 U8573 ( .A1(n6760), .A2(n5029), .ZN(n6790) );
  AOI21_X1 U8574 ( .B1(n5029), .B2(n6760), .A(n6790), .ZN(n6761) );
  OAI22_X1 U8575 ( .A1(n6762), .A2(n6761), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10385), .ZN(n6763) );
  AOI21_X1 U8576 ( .B1(n10159), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n6763), .ZN(
        n6764) );
  OAI21_X1 U8577 ( .B1(n5029), .B2(n10157), .A(n6764), .ZN(P2_U3182) );
  INV_X1 U8578 ( .A(n6766), .ZN(n6767) );
  AOI21_X1 U8579 ( .B1(n6765), .B2(n6768), .A(n6767), .ZN(n6775) );
  NAND2_X1 U8580 ( .A1(n6276), .A2(n9066), .ZN(n6770) );
  NAND2_X1 U8581 ( .A1(n9098), .A2(n8777), .ZN(n6769) );
  NAND2_X1 U8582 ( .A1(n6770), .A2(n6769), .ZN(n7210) );
  AOI22_X1 U8583 ( .A1(P1_REG3_REG_2__SCAN_IN), .A2(n6771), .B1(n8763), .B2(
        n7210), .ZN(n6774) );
  NAND2_X1 U8584 ( .A1(n8767), .A2(n6772), .ZN(n6773) );
  OAI211_X1 U8585 ( .C1(n6775), .C2(n8769), .A(n6774), .B(n6773), .ZN(P1_U3237) );
  INV_X1 U8586 ( .A(n6776), .ZN(n6799) );
  INV_X1 U8587 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6777) );
  OAI222_X1 U8588 ( .A1(n9572), .A2(n6799), .B1(n6778), .B2(P1_U3086), .C1(
        n6777), .C2(n9569), .ZN(P1_U3343) );
  INV_X1 U8589 ( .A(n10153), .ZN(n6782) );
  NAND2_X1 U8590 ( .A1(n6784), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6845) );
  NAND2_X1 U8591 ( .A1(n5029), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6779) );
  OR2_X1 U8592 ( .A1(n6779), .A2(n6784), .ZN(n6780) );
  XOR2_X1 U8593 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6844), .Z(n6781) );
  OAI22_X1 U8594 ( .A1(n6782), .A2(n6781), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7141), .ZN(n6796) );
  NOR2_X1 U8595 ( .A1(n6783), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6785) );
  NAND2_X1 U8596 ( .A1(n6784), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6838) );
  OAI21_X1 U8597 ( .B1(n6854), .B2(n6785), .A(n6838), .ZN(n6786) );
  NAND2_X1 U8598 ( .A1(n6786), .A2(n5760), .ZN(n6789) );
  INV_X1 U8599 ( .A(n6787), .ZN(n6788) );
  OR2_X1 U8600 ( .A1(n6788), .A2(n8291), .ZN(n10147) );
  AOI21_X1 U8601 ( .B1(n6839), .B2(n6789), .A(n10147), .ZN(n6795) );
  MUX2_X1 U8602 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8291), .Z(n6855) );
  XNOR2_X1 U8603 ( .A(n6855), .B(n6854), .ZN(n6791) );
  AOI21_X1 U8604 ( .B1(n6791), .B2(n6790), .A(n10140), .ZN(n6792) );
  INV_X1 U8605 ( .A(n6792), .ZN(n6793) );
  OAI22_X1 U8606 ( .A1(n9837), .A2(n10284), .B1(n6853), .B2(n6793), .ZN(n6794)
         );
  NOR3_X1 U8607 ( .A1(n6796), .A2(n6795), .A3(n6794), .ZN(n6797) );
  OAI21_X1 U8608 ( .B1(n6854), .B2(n10157), .A(n6797), .ZN(P2_U3183) );
  INV_X1 U8609 ( .A(n9919), .ZN(n8304) );
  INV_X1 U8610 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6798) );
  OAI222_X1 U8611 ( .A1(P2_U3151), .A2(n8304), .B1(n6582), .B2(n6799), .C1(
        n6798), .C2(n8668), .ZN(P2_U3283) );
  INV_X1 U8612 ( .A(n6800), .ZN(n6813) );
  AOI22_X1 U8613 ( .A1(n9633), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9563), .ZN(n6801) );
  OAI21_X1 U8614 ( .B1(n6813), .B2(n9572), .A(n6801), .ZN(P1_U3342) );
  XNOR2_X1 U8615 ( .A(n8789), .B(n6807), .ZN(n6802) );
  AOI22_X1 U8616 ( .A1(n9066), .A2(n6285), .B1(n9097), .B2(n8777), .ZN(n6818)
         );
  OAI21_X1 U8617 ( .B1(n6802), .B2(n9752), .A(n6818), .ZN(n7125) );
  AOI21_X1 U8618 ( .B1(n6803), .B2(n6804), .A(n9422), .ZN(n6805) );
  AND2_X1 U8619 ( .A1(n6942), .A2(n6805), .ZN(n7128) );
  NOR2_X1 U8620 ( .A1(n7125), .A2(n7128), .ZN(n6835) );
  OAI21_X1 U8621 ( .B1(n6808), .B2(n6807), .A(n6806), .ZN(n7132) );
  INV_X1 U8622 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6809) );
  OAI22_X1 U8623 ( .A1(n9543), .A2(n4768), .B1(n9788), .B2(n6809), .ZN(n6810)
         );
  AOI21_X1 U8624 ( .B1(n7132), .B2(n7714), .A(n6810), .ZN(n6811) );
  OAI21_X1 U8625 ( .B1(n6835), .B2(n9786), .A(n6811), .ZN(P1_U3462) );
  INV_X1 U8626 ( .A(n9936), .ZN(n8321) );
  INV_X1 U8627 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6812) );
  OAI222_X1 U8628 ( .A1(n8321), .A2(P2_U3151), .B1(n6582), .B2(n6813), .C1(
        n6812), .C2(n8668), .ZN(P2_U3282) );
  OAI21_X1 U8629 ( .B1(n6816), .B2(n6815), .A(n6814), .ZN(n6817) );
  NAND2_X1 U8630 ( .A1(n6817), .A2(n8775), .ZN(n6821) );
  OAI22_X1 U8631 ( .A1(n8780), .A2(n6818), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7127), .ZN(n6819) );
  AOI21_X1 U8632 ( .B1(n8782), .B2(n7127), .A(n6819), .ZN(n6820) );
  OAI211_X1 U8633 ( .C1(n4768), .C2(n8785), .A(n6821), .B(n6820), .ZN(P1_U3218) );
  INV_X1 U8634 ( .A(n6822), .ZN(n6837) );
  AOI22_X1 U8635 ( .A1(n9645), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9563), .ZN(n6823) );
  OAI21_X1 U8636 ( .B1(n6837), .B2(n9572), .A(n6823), .ZN(P1_U3341) );
  AOI21_X1 U8637 ( .B1(n6824), .B2(n6825), .A(n8769), .ZN(n6827) );
  NAND2_X1 U8638 ( .A1(n6827), .A2(n6826), .ZN(n6832) );
  NAND2_X1 U8639 ( .A1(n9098), .A2(n9066), .ZN(n6829) );
  NAND2_X1 U8640 ( .A1(n9096), .A2(n8777), .ZN(n6828) );
  AND2_X1 U8641 ( .A1(n6829), .A2(n6828), .ZN(n6946) );
  INV_X1 U8642 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n10296) );
  OAI22_X1 U8643 ( .A1(n8780), .A2(n6946), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10296), .ZN(n6830) );
  AOI21_X1 U8644 ( .B1(n9734), .B2(n8782), .A(n6830), .ZN(n6831) );
  OAI211_X1 U8645 ( .C1(n9738), .C2(n8785), .A(n6832), .B(n6831), .ZN(P1_U3230) );
  OAI22_X1 U8646 ( .A1(n9469), .A2(n4768), .B1(n9797), .B2(n6690), .ZN(n6833)
         );
  AOI21_X1 U8647 ( .B1(n7132), .B2(n7727), .A(n6833), .ZN(n6834) );
  OAI21_X1 U8648 ( .B1(n6835), .B2(n9795), .A(n6834), .ZN(P1_U3525) );
  INV_X1 U8649 ( .A(n9952), .ZN(n8303) );
  INV_X1 U8650 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6836) );
  OAI222_X1 U8651 ( .A1(n8303), .A2(P2_U3151), .B1(n6582), .B2(n6837), .C1(
        n6836), .C2(n8668), .ZN(P2_U3281) );
  INV_X1 U8652 ( .A(n10157), .ZN(n10002) );
  INV_X1 U8653 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6852) );
  INV_X1 U8654 ( .A(n10147), .ZN(n9980) );
  INV_X1 U8655 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10037) );
  MUX2_X1 U8656 ( .A(n10037), .B(P2_REG2_REG_2__SCAN_IN), .S(n7008), .Z(n6841)
         );
  NAND2_X1 U8657 ( .A1(n6841), .A2(n6840), .ZN(n6999) );
  OAI21_X1 U8658 ( .B1(n6841), .B2(n6840), .A(n6999), .ZN(n6842) );
  AOI22_X1 U8659 ( .A1(n9980), .A2(n6842), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n6851) );
  MUX2_X1 U8660 ( .A(n6843), .B(P2_REG1_REG_2__SCAN_IN), .S(n7008), .Z(n6848)
         );
  NAND2_X1 U8661 ( .A1(n6846), .A2(n6845), .ZN(n6847) );
  NAND2_X1 U8662 ( .A1(n6848), .A2(n6847), .ZN(n7010) );
  OAI21_X1 U8663 ( .B1(n6848), .B2(n6847), .A(n7010), .ZN(n6849) );
  NAND2_X1 U8664 ( .A1(n10153), .A2(n6849), .ZN(n6850) );
  OAI211_X1 U8665 ( .C1(n6852), .C2(n9837), .A(n6851), .B(n6850), .ZN(n6859)
         );
  MUX2_X1 U8666 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8291), .Z(n6989) );
  XOR2_X1 U8667 ( .A(n7008), .B(n6989), .Z(n6857) );
  NOR2_X1 U8668 ( .A1(n6856), .A2(n6857), .ZN(n6987) );
  AOI211_X1 U8669 ( .C1(n6857), .C2(n6856), .A(n10140), .B(n6987), .ZN(n6858)
         );
  AOI211_X1 U8670 ( .C1(n10002), .C2(n7008), .A(n6859), .B(n6858), .ZN(n6860)
         );
  INV_X1 U8671 ( .A(n6860), .ZN(P2_U3184) );
  OAI21_X1 U8672 ( .B1(n6863), .B2(n6862), .A(n6861), .ZN(n6867) );
  AND2_X1 U8673 ( .A1(n6865), .A2(n6864), .ZN(n6866) );
  OAI211_X1 U8674 ( .C1(n6872), .C2(n6868), .A(n6867), .B(n6866), .ZN(n6869)
         );
  NAND2_X1 U8675 ( .A1(n6869), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6875) );
  INV_X1 U8676 ( .A(n6883), .ZN(n6870) );
  OR2_X1 U8677 ( .A1(n6904), .A2(n6870), .ZN(n7990) );
  OR2_X1 U8678 ( .A1(n6871), .A2(P2_U3151), .ZN(n7994) );
  OAI21_X1 U8679 ( .B1(n6872), .B2(n7990), .A(n7994), .ZN(n6873) );
  INV_X1 U8680 ( .A(n6873), .ZN(n6874) );
  NAND2_X1 U8681 ( .A1(n6875), .A2(n6874), .ZN(n8199) );
  NOR2_X1 U8682 ( .A1(n8199), .A2(P2_U3151), .ZN(n6918) );
  NAND2_X1 U8683 ( .A1(n6906), .A2(n6876), .ZN(n6880) );
  INV_X1 U8684 ( .A(n6877), .ZN(n6878) );
  NAND2_X1 U8685 ( .A1(n6881), .A2(n6878), .ZN(n6879) );
  INV_X1 U8686 ( .A(n8206), .ZN(n7238) );
  NAND2_X1 U8687 ( .A1(n8246), .A2(n6888), .ZN(n7818) );
  NAND2_X1 U8688 ( .A1(n7824), .A2(n7818), .ZN(n10039) );
  NAND2_X1 U8689 ( .A1(n6881), .A2(n10090), .ZN(n6885) );
  INV_X1 U8690 ( .A(n6882), .ZN(n6884) );
  INV_X1 U8691 ( .A(n8192), .ZN(n8220) );
  NOR2_X1 U8692 ( .A1(n6904), .A2(n6886), .ZN(n6887) );
  NAND2_X1 U8693 ( .A1(n6906), .A2(n6887), .ZN(n8212) );
  INV_X1 U8694 ( .A(n8245), .ZN(n10030) );
  OAI22_X1 U8695 ( .A1(n8220), .A2(n6888), .B1(n8212), .B2(n10030), .ZN(n6889)
         );
  AOI21_X1 U8696 ( .B1(n7238), .B2(n10039), .A(n6889), .ZN(n6890) );
  OAI21_X1 U8697 ( .B1(n6918), .B2(n10385), .A(n6890), .ZN(P2_U3172) );
  AOI21_X1 U8698 ( .B1(n7825), .B2(n7948), .A(n6891), .ZN(n6892) );
  XNOR2_X1 U8699 ( .A(n6894), .B(n6895), .ZN(n6974) );
  XNOR2_X1 U8700 ( .A(n6974), .B(n8244), .ZN(n6901) );
  XNOR2_X1 U8701 ( .A(n6895), .B(n10047), .ZN(n6896) );
  NOR2_X1 U8702 ( .A1(n6896), .A2(n8245), .ZN(n6898) );
  NOR2_X1 U8703 ( .A1(n6898), .A2(n6897), .ZN(n6912) );
  OAI21_X1 U8704 ( .B1(n10044), .B2(n8052), .A(n7824), .ZN(n6911) );
  NAND2_X1 U8705 ( .A1(n6912), .A2(n6911), .ZN(n6910) );
  INV_X1 U8706 ( .A(n6898), .ZN(n6899) );
  NAND2_X1 U8707 ( .A1(n6910), .A2(n6899), .ZN(n6900) );
  NAND2_X1 U8708 ( .A1(n6900), .A2(n6901), .ZN(n6975) );
  OAI21_X1 U8709 ( .B1(n6901), .B2(n6900), .A(n6975), .ZN(n6902) );
  NAND2_X1 U8710 ( .A1(n6902), .A2(n7238), .ZN(n6909) );
  NOR2_X1 U8711 ( .A1(n6904), .A2(n6903), .ZN(n6905) );
  NAND2_X1 U8712 ( .A1(n6906), .A2(n6905), .ZN(n8190) );
  OAI22_X1 U8713 ( .A1(n8220), .A2(n10050), .B1(n8190), .B2(n10030), .ZN(n6907) );
  AOI21_X1 U8714 ( .B1(n8187), .B2(n8243), .A(n6907), .ZN(n6908) );
  OAI211_X1 U8715 ( .C1(n6918), .C2(n10021), .A(n6909), .B(n6908), .ZN(
        P2_U3177) );
  OAI21_X1 U8716 ( .B1(n6912), .B2(n6911), .A(n6910), .ZN(n6913) );
  NAND2_X1 U8717 ( .A1(n6913), .A2(n7238), .ZN(n6917) );
  INV_X1 U8718 ( .A(n8246), .ZN(n6914) );
  OAI22_X1 U8719 ( .A1(n8220), .A2(n10047), .B1(n8190), .B2(n6914), .ZN(n6915)
         );
  AOI21_X1 U8720 ( .B1(n8187), .B2(n8244), .A(n6915), .ZN(n6916) );
  OAI211_X1 U8721 ( .C1(n6918), .C2(n7141), .A(n6917), .B(n6916), .ZN(P2_U3162) );
  NAND2_X1 U8722 ( .A1(n8793), .A2(n8790), .ZN(n6919) );
  XNOR2_X1 U8723 ( .A(n6919), .B(n6926), .ZN(n6922) );
  NAND2_X1 U8724 ( .A1(n9097), .A2(n9066), .ZN(n6921) );
  NAND2_X1 U8725 ( .A1(n9095), .A2(n8777), .ZN(n6920) );
  AND2_X1 U8726 ( .A1(n6921), .A2(n6920), .ZN(n7046) );
  OAI21_X1 U8727 ( .B1(n6922), .B2(n9752), .A(n7046), .ZN(n7261) );
  INV_X1 U8728 ( .A(n6941), .ZN(n6924) );
  INV_X1 U8729 ( .A(n6961), .ZN(n6923) );
  AOI211_X1 U8730 ( .C1(n6925), .C2(n6924), .A(n9422), .B(n6923), .ZN(n7266)
         );
  NOR2_X1 U8731 ( .A1(n7261), .A2(n7266), .ZN(n6935) );
  OR2_X1 U8732 ( .A1(n6927), .A2(n6926), .ZN(n6928) );
  NAND2_X1 U8733 ( .A1(n6929), .A2(n6928), .ZN(n7260) );
  OAI22_X1 U8734 ( .A1(n9469), .A2(n7264), .B1(n9797), .B2(n10360), .ZN(n6930)
         );
  AOI21_X1 U8735 ( .B1(n7260), .B2(n7727), .A(n6930), .ZN(n6931) );
  OAI21_X1 U8736 ( .B1(n6935), .B2(n9795), .A(n6931), .ZN(P1_U3527) );
  INV_X1 U8737 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6932) );
  OAI22_X1 U8738 ( .A1(n9543), .A2(n7264), .B1(n9788), .B2(n6932), .ZN(n6933)
         );
  AOI21_X1 U8739 ( .B1(n7260), .B2(n7714), .A(n6933), .ZN(n6934) );
  OAI21_X1 U8740 ( .B1(n6935), .B2(n9786), .A(n6934), .ZN(P1_U3468) );
  INV_X1 U8741 ( .A(n9969), .ZN(n8324) );
  INV_X1 U8742 ( .A(n6936), .ZN(n6938) );
  INV_X1 U8743 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6937) );
  OAI222_X1 U8744 ( .A1(n8324), .A2(P2_U3151), .B1(n6582), .B2(n6938), .C1(
        n6937), .C2(n8668), .ZN(P2_U3280) );
  INV_X1 U8745 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10484) );
  OAI222_X1 U8746 ( .A1(n9569), .A2(n10484), .B1(n9572), .B2(n6938), .C1(
        P1_U3086), .C2(n9218), .ZN(P1_U3340) );
  OAI21_X1 U8747 ( .B1(n6939), .B2(n6944), .A(n6940), .ZN(n9740) );
  AOI211_X1 U8748 ( .C1(n6943), .C2(n6942), .A(n9422), .B(n6941), .ZN(n9732)
         );
  INV_X1 U8749 ( .A(n6944), .ZN(n8932) );
  XNOR2_X1 U8750 ( .A(n6945), .B(n8932), .ZN(n6948) );
  INV_X1 U8751 ( .A(n6946), .ZN(n6947) );
  AOI21_X1 U8752 ( .B1(n6948), .B2(n9710), .A(n6947), .ZN(n9743) );
  INV_X1 U8753 ( .A(n9743), .ZN(n6949) );
  AOI211_X1 U8754 ( .C1(n9768), .C2(n9740), .A(n9732), .B(n6949), .ZN(n6955)
         );
  INV_X1 U8755 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6950) );
  OAI22_X1 U8756 ( .A1(n9543), .A2(n9738), .B1(n9788), .B2(n6950), .ZN(n6951)
         );
  INV_X1 U8757 ( .A(n6951), .ZN(n6952) );
  OAI21_X1 U8758 ( .B1(n6955), .B2(n9786), .A(n6952), .ZN(P1_U3465) );
  OAI22_X1 U8759 ( .A1(n9469), .A2(n9738), .B1(n9797), .B2(n6692), .ZN(n6953)
         );
  INV_X1 U8760 ( .A(n6953), .ZN(n6954) );
  OAI21_X1 U8761 ( .B1(n6955), .B2(n9795), .A(n6954), .ZN(P1_U3526) );
  INV_X1 U8762 ( .A(n6956), .ZN(n6973) );
  AOI22_X1 U8763 ( .A1(n9674), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9563), .ZN(n6957) );
  OAI21_X1 U8764 ( .B1(n6973), .B2(n9572), .A(n6957), .ZN(P1_U3339) );
  XOR2_X1 U8765 ( .A(n6963), .B(n6958), .Z(n6959) );
  AOI22_X1 U8766 ( .A1(n9066), .A2(n9096), .B1(n9094), .B2(n8777), .ZN(n7103)
         );
  OAI21_X1 U8767 ( .B1(n6959), .B2(n9752), .A(n7103), .ZN(n7250) );
  INV_X1 U8768 ( .A(n7195), .ZN(n6960) );
  AOI211_X1 U8769 ( .C1(n6965), .C2(n6961), .A(n9422), .B(n6960), .ZN(n7256)
         );
  NOR2_X1 U8770 ( .A1(n7250), .A2(n7256), .ZN(n6972) );
  OAI21_X1 U8771 ( .B1(n6964), .B2(n6963), .A(n6962), .ZN(n7249) );
  INV_X1 U8772 ( .A(n6965), .ZN(n7254) );
  OAI22_X1 U8773 ( .A1(n9469), .A2(n7254), .B1(n9797), .B2(n6966), .ZN(n6967)
         );
  AOI21_X1 U8774 ( .B1(n7249), .B2(n7727), .A(n6967), .ZN(n6968) );
  OAI21_X1 U8775 ( .B1(n6972), .B2(n9795), .A(n6968), .ZN(P1_U3528) );
  INV_X1 U8776 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6969) );
  OAI22_X1 U8777 ( .A1(n9543), .A2(n7254), .B1(n9788), .B2(n6969), .ZN(n6970)
         );
  AOI21_X1 U8778 ( .B1(n7249), .B2(n7714), .A(n6970), .ZN(n6971) );
  OAI21_X1 U8779 ( .B1(n6972), .B2(n9786), .A(n6971), .ZN(P1_U3471) );
  OAI222_X1 U8780 ( .A1(P2_U3151), .A2(n8302), .B1(n6582), .B2(n6973), .C1(
        n10341), .C2(n8668), .ZN(P2_U3279) );
  INV_X2 U8781 ( .A(n8056), .ZN(n8052) );
  XNOR2_X1 U8782 ( .A(n10055), .B(n8052), .ZN(n7087) );
  XNOR2_X1 U8783 ( .A(n7087), .B(n8243), .ZN(n6978) );
  INV_X1 U8784 ( .A(n6974), .ZN(n6976) );
  OAI21_X1 U8785 ( .B1(n6976), .B2(n8244), .A(n6975), .ZN(n6977) );
  AOI211_X1 U8786 ( .C1(n6978), .C2(n6977), .A(n8206), .B(n7086), .ZN(n6979)
         );
  INV_X1 U8787 ( .A(n6979), .ZN(n6983) );
  AND2_X1 U8788 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9802) );
  INV_X1 U8789 ( .A(n8244), .ZN(n6980) );
  INV_X1 U8790 ( .A(n8242), .ZN(n7167) );
  OAI22_X1 U8791 ( .A1(n6980), .A2(n8190), .B1(n8212), .B2(n7167), .ZN(n6981)
         );
  AOI211_X1 U8792 ( .C1(n7122), .C2(n8192), .A(n9802), .B(n6981), .ZN(n6982)
         );
  OAI211_X1 U8793 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8214), .A(n6983), .B(
        n6982), .ZN(P2_U3158) );
  MUX2_X1 U8794 ( .A(n6985), .B(n6984), .S(n8291), .Z(n6993) );
  INV_X1 U8795 ( .A(n6993), .ZN(n6994) );
  MUX2_X1 U8796 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8291), .Z(n6992) );
  XNOR2_X1 U8797 ( .A(n6992), .B(n7015), .ZN(n9825) );
  MUX2_X1 U8798 ( .A(n7120), .B(n6986), .S(n8291), .Z(n6991) );
  XNOR2_X1 U8799 ( .A(n6991), .B(n9798), .ZN(n9810) );
  NAND2_X1 U8800 ( .A1(n9810), .A2(n9811), .ZN(n9809) );
  INV_X1 U8801 ( .A(n9809), .ZN(n6990) );
  AOI21_X1 U8802 ( .B1(n6991), .B2(n7011), .A(n6990), .ZN(n9823) );
  XNOR2_X1 U8803 ( .A(n6993), .B(n7017), .ZN(n10142) );
  NOR2_X1 U8804 ( .A1(n10141), .A2(n10142), .ZN(n10139) );
  MUX2_X1 U8805 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8291), .Z(n8278) );
  XNOR2_X1 U8806 ( .A(n8278), .B(n8309), .ZN(n6995) );
  NAND2_X1 U8807 ( .A1(n6996), .A2(n6995), .ZN(n8276) );
  OAI21_X1 U8808 ( .B1(n6996), .B2(n6995), .A(n8276), .ZN(n6997) );
  NAND2_X1 U8809 ( .A1(n6997), .A2(n10010), .ZN(n7027) );
  OR2_X1 U8810 ( .A1(n7008), .A2(n10037), .ZN(n6998) );
  NAND2_X1 U8811 ( .A1(n6999), .A2(n6998), .ZN(n7000) );
  NAND2_X1 U8812 ( .A1(n7000), .A2(n9798), .ZN(n9818) );
  INV_X1 U8813 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10379) );
  MUX2_X1 U8814 ( .A(n10379), .B(P2_REG2_REG_4__SCAN_IN), .S(n7015), .Z(n9816)
         );
  OR2_X1 U8815 ( .A1(n7015), .A2(n10379), .ZN(n7003) );
  NAND2_X1 U8816 ( .A1(n9820), .A2(n7003), .ZN(n7004) );
  XNOR2_X1 U8817 ( .A(n8309), .B(n7273), .ZN(n7006) );
  AND3_X1 U8818 ( .A1(n10149), .A2(n7006), .A3(n7005), .ZN(n7007) );
  NOR2_X1 U8819 ( .A1(n8247), .A2(n7007), .ZN(n7024) );
  MUX2_X1 U8820 ( .A(n8308), .B(P2_REG1_REG_6__SCAN_IN), .S(n8309), .Z(n7021)
         );
  OR2_X1 U8821 ( .A1(n7008), .A2(n6843), .ZN(n7009) );
  NAND2_X1 U8822 ( .A1(n7010), .A2(n7009), .ZN(n7012) );
  NAND2_X1 U8823 ( .A1(n7012), .A2(n9798), .ZN(n7013) );
  XNOR2_X1 U8824 ( .A(n7012), .B(n7011), .ZN(n9800) );
  NAND2_X1 U8825 ( .A1(P2_REG1_REG_3__SCAN_IN), .A2(n9800), .ZN(n9799) );
  NAND2_X1 U8826 ( .A1(n7013), .A2(n9799), .ZN(n9829) );
  MUX2_X1 U8827 ( .A(n7014), .B(P2_REG1_REG_4__SCAN_IN), .S(n7015), .Z(n9830)
         );
  NAND2_X1 U8828 ( .A1(n9829), .A2(n9830), .ZN(n9828) );
  OR2_X1 U8829 ( .A1(n7015), .A2(n7014), .ZN(n7016) );
  NAND2_X1 U8830 ( .A1(n7018), .A2(n10156), .ZN(n7019) );
  NAND2_X1 U8831 ( .A1(n7020), .A2(n7021), .ZN(n8307) );
  OAI21_X1 U8832 ( .B1(n7021), .B2(n7020), .A(n8307), .ZN(n7022) );
  NAND2_X1 U8833 ( .A1(n10153), .A2(n7022), .ZN(n7023) );
  NAND2_X1 U8834 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7240) );
  OAI211_X1 U8835 ( .C1(n7024), .C2(n10147), .A(n7023), .B(n7240), .ZN(n7025)
         );
  AOI21_X1 U8836 ( .B1(n10159), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n7025), .ZN(
        n7026) );
  OAI211_X1 U8837 ( .C1(n10157), .C2(n8277), .A(n7027), .B(n7026), .ZN(
        P2_U3188) );
  INV_X1 U8838 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7040) );
  NAND2_X1 U8839 ( .A1(n7029), .A2(n7028), .ZN(n7032) );
  INV_X2 U8840 ( .A(n9744), .ZN(n9409) );
  INV_X1 U8841 ( .A(n7030), .ZN(n7031) );
  NOR2_X2 U8842 ( .A1(n7032), .A2(n6252), .ZN(n9731) );
  AND2_X1 U8843 ( .A1(n9731), .A2(n9724), .ZN(n9262) );
  OAI21_X1 U8844 ( .B1(n9722), .B2(n9262), .A(n9755), .ZN(n7039) );
  INV_X1 U8845 ( .A(n7148), .ZN(n7034) );
  NAND2_X1 U8846 ( .A1(n6265), .A2(n7033), .ZN(n9025) );
  AND2_X1 U8847 ( .A1(n7034), .A2(n9025), .ZN(n9750) );
  INV_X1 U8848 ( .A(n9405), .ZN(n9733) );
  AOI21_X1 U8849 ( .B1(n9733), .B2(P1_REG3_REG_0__SCAN_IN), .A(n9754), .ZN(
        n7035) );
  OAI21_X1 U8850 ( .B1(n9750), .B2(n7036), .A(n7035), .ZN(n7037) );
  NAND2_X1 U8851 ( .A1(n9409), .A2(n7037), .ZN(n7038) );
  OAI211_X1 U8852 ( .C1(n7040), .C2(n9409), .A(n7039), .B(n7038), .ZN(P1_U3293) );
  AND2_X1 U8853 ( .A1(n7096), .A2(n7041), .ZN(n7043) );
  OAI21_X1 U8854 ( .B1(n7044), .B2(n7043), .A(n7042), .ZN(n7045) );
  NAND2_X1 U8855 ( .A1(n7045), .A2(n8775), .ZN(n7050) );
  NAND2_X1 U8856 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9154) );
  OAI21_X1 U8857 ( .B1(n8780), .B2(n7046), .A(n9154), .ZN(n7047) );
  AOI21_X1 U8858 ( .B1(n7048), .B2(n8782), .A(n7047), .ZN(n7049) );
  OAI211_X1 U8859 ( .C1(n7264), .C2(n8785), .A(n7050), .B(n7049), .ZN(P1_U3227) );
  NAND3_X1 U8860 ( .A1(n7118), .A2(n7849), .A3(n7053), .ZN(n7054) );
  NAND2_X1 U8861 ( .A1(n7052), .A2(n7054), .ZN(n7234) );
  INV_X1 U8862 ( .A(n8241), .ZN(n7245) );
  NAND2_X1 U8863 ( .A1(n7055), .A2(n7056), .ZN(n7057) );
  XNOR2_X1 U8864 ( .A(n7057), .B(n7957), .ZN(n7058) );
  OAI222_X1 U8865 ( .A1(n10032), .A2(n7245), .B1(n10031), .B2(n4735), .C1(
        n10041), .C2(n7058), .ZN(n7231) );
  AOI21_X1 U8866 ( .B1(n10082), .B2(n7234), .A(n7231), .ZN(n7062) );
  INV_X1 U8867 ( .A(n8604), .ZN(n8539) );
  AOI22_X1 U8868 ( .A1(n8539), .A2(n7093), .B1(n10103), .B2(
        P2_REG1_REG_4__SCAN_IN), .ZN(n7059) );
  OAI21_X1 U8869 ( .B1(n7062), .B2(n10103), .A(n7059), .ZN(P2_U3463) );
  OAI22_X1 U8870 ( .A1(n7230), .A2(n8662), .B1(n10091), .B2(n5795), .ZN(n7060)
         );
  INV_X1 U8871 ( .A(n7060), .ZN(n7061) );
  OAI21_X1 U8872 ( .B1(n7062), .B2(n10093), .A(n7061), .ZN(P2_U3402) );
  INV_X1 U8873 ( .A(n8240), .ZN(n7318) );
  NAND2_X1 U8874 ( .A1(n7055), .A2(n7063), .ZN(n7065) );
  AND2_X1 U8875 ( .A1(n7065), .A2(n7064), .ZN(n7066) );
  XNOR2_X1 U8876 ( .A(n7066), .B(n4528), .ZN(n7067) );
  OAI222_X1 U8877 ( .A1(n10032), .A2(n7318), .B1(n10031), .B2(n7167), .C1(
        n10041), .C2(n7067), .ZN(n7108) );
  INV_X1 U8878 ( .A(n7108), .ZN(n7081) );
  MUX2_X1 U8879 ( .A(n7070), .B(n7069), .S(n7068), .Z(n7072) );
  NAND2_X1 U8880 ( .A1(n7072), .A2(n7071), .ZN(n7077) );
  INV_X2 U8881 ( .A(n10035), .ZN(n10038) );
  OR2_X1 U8882 ( .A1(n7073), .A2(n4528), .ZN(n7074) );
  NAND2_X1 U8883 ( .A1(n7075), .A2(n7074), .ZN(n7109) );
  AND2_X1 U8884 ( .A1(n7076), .A2(n7825), .ZN(n7295) );
  OR2_X1 U8885 ( .A1(n7296), .A2(n7295), .ZN(n10034) );
  NOR2_X1 U8886 ( .A1(n8532), .A2(n7113), .ZN(n7079) );
  OAI22_X1 U8887 ( .A1(n10035), .A2(n6985), .B1(n7172), .B2(n10022), .ZN(n7078) );
  AOI211_X1 U8888 ( .C1(n7109), .C2(n8536), .A(n7079), .B(n7078), .ZN(n7080)
         );
  OAI21_X1 U8889 ( .B1(n7081), .B2(n10038), .A(n7080), .ZN(P2_U3228) );
  INV_X1 U8890 ( .A(n7082), .ZN(n7085) );
  INV_X1 U8891 ( .A(n9224), .ZN(n9687) );
  OAI222_X1 U8892 ( .A1(n9569), .A2(n7083), .B1(n9572), .B2(n7085), .C1(
        P1_U3086), .C2(n9687), .ZN(P1_U3338) );
  INV_X1 U8893 ( .A(n10003), .ZN(n8328) );
  OAI222_X1 U8894 ( .A1(n8328), .A2(P2_U3151), .B1(n6582), .B2(n7085), .C1(
        n7084), .C2(n8668), .ZN(P2_U3278) );
  XNOR2_X1 U8895 ( .A(n7230), .B(n8052), .ZN(n7088) );
  NOR2_X1 U8896 ( .A1(n7088), .A2(n8242), .ZN(n7161) );
  AOI21_X1 U8897 ( .B1(n7088), .B2(n8242), .A(n7161), .ZN(n7089) );
  OAI21_X1 U8898 ( .B1(n7090), .B2(n7089), .A(n7164), .ZN(n7091) );
  NAND2_X1 U8899 ( .A1(n7091), .A2(n7238), .ZN(n7095) );
  NOR2_X1 U8900 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5796), .ZN(n9821) );
  OAI22_X1 U8901 ( .A1(n4735), .A2(n8190), .B1(n8212), .B2(n7245), .ZN(n7092)
         );
  AOI211_X1 U8902 ( .C1(n7093), .C2(n8192), .A(n9821), .B(n7092), .ZN(n7094)
         );
  OAI211_X1 U8903 ( .C1(n7229), .C2(n8214), .A(n7095), .B(n7094), .ZN(P2_U3170) );
  INV_X1 U8904 ( .A(n7042), .ZN(n7099) );
  INV_X1 U8905 ( .A(n7096), .ZN(n7098) );
  NOR3_X1 U8906 ( .A1(n7099), .A2(n7098), .A3(n7097), .ZN(n7102) );
  INV_X1 U8907 ( .A(n7100), .ZN(n7101) );
  OAI21_X1 U8908 ( .B1(n7102), .B2(n7101), .A(n8775), .ZN(n7107) );
  NAND2_X1 U8909 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9166) );
  INV_X1 U8910 ( .A(n9166), .ZN(n7105) );
  NOR2_X1 U8911 ( .A1(n8780), .A2(n7103), .ZN(n7104) );
  AOI211_X1 U8912 ( .C1(n8782), .C2(n7252), .A(n7105), .B(n7104), .ZN(n7106)
         );
  OAI211_X1 U8913 ( .C1(n7254), .C2(n8785), .A(n7107), .B(n7106), .ZN(P1_U3239) );
  AOI21_X1 U8914 ( .B1(n10082), .B2(n7109), .A(n7108), .ZN(n7116) );
  INV_X1 U8915 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7110) );
  OAI22_X1 U8916 ( .A1(n7113), .A2(n8662), .B1(n10091), .B2(n7110), .ZN(n7111)
         );
  INV_X1 U8917 ( .A(n7111), .ZN(n7112) );
  OAI21_X1 U8918 ( .B1(n7116), .B2(n10093), .A(n7112), .ZN(P2_U3405) );
  OAI22_X1 U8919 ( .A1(n8604), .A2(n7113), .B1(n10105), .B2(n6984), .ZN(n7114)
         );
  INV_X1 U8920 ( .A(n7114), .ZN(n7115) );
  OAI21_X1 U8921 ( .B1(n7116), .B2(n10103), .A(n7115), .ZN(P2_U3464) );
  NAND3_X1 U8922 ( .A1(n10019), .A2(n7828), .A3(n7955), .ZN(n7117) );
  AND2_X1 U8923 ( .A1(n7118), .A2(n7117), .ZN(n10056) );
  INV_X1 U8924 ( .A(n8536), .ZN(n7546) );
  AOI222_X1 U8925 ( .A1(n8516), .A2(n7119), .B1(n8242), .B2(n8511), .C1(n8244), 
        .C2(n8513), .ZN(n10054) );
  MUX2_X1 U8926 ( .A(n7120), .B(n10054), .S(n10035), .Z(n7124) );
  INV_X1 U8927 ( .A(n8532), .ZN(n8519) );
  INV_X1 U8928 ( .A(n10022), .ZN(n8505) );
  AOI22_X1 U8929 ( .A1(n8519), .A2(n7122), .B1(n8505), .B2(n7121), .ZN(n7123)
         );
  OAI211_X1 U8930 ( .C1(n10056), .C2(n7546), .A(n7124), .B(n7123), .ZN(
        P2_U3230) );
  INV_X1 U8931 ( .A(n7125), .ZN(n7134) );
  AND2_X1 U8932 ( .A1(n7737), .A2(n7194), .ZN(n7126) );
  AOI22_X1 U8933 ( .A1(n9744), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9733), .B2(
        n7127), .ZN(n7130) );
  NAND2_X1 U8934 ( .A1(n9731), .A2(n7128), .ZN(n7129) );
  OAI211_X1 U8935 ( .C1(n9737), .C2(n4768), .A(n7130), .B(n7129), .ZN(n7131)
         );
  AOI21_X1 U8936 ( .B1(n9741), .B2(n7132), .A(n7131), .ZN(n7133) );
  OAI21_X1 U8937 ( .B1(n9744), .B2(n7134), .A(n7133), .ZN(P1_U3290) );
  NOR2_X1 U8938 ( .A1(n10030), .A2(n10032), .ZN(n10043) );
  AOI21_X1 U8939 ( .B1(n7135), .B2(n10039), .A(n10043), .ZN(n7138) );
  AOI22_X1 U8940 ( .A1(n8519), .A2(n10044), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n8505), .ZN(n7137) );
  OR2_X1 U8941 ( .A1(n10035), .A2(n6783), .ZN(n7136) );
  OAI211_X1 U8942 ( .C1(n7138), .C2(n10038), .A(n7137), .B(n7136), .ZN(
        P2_U3233) );
  OAI21_X1 U8943 ( .B1(n7139), .B2(n7954), .A(n10026), .ZN(n7140) );
  AOI222_X1 U8944 ( .A1(n8516), .A2(n7140), .B1(n8244), .B2(n8511), .C1(n8246), 
        .C2(n8513), .ZN(n10046) );
  OAI22_X1 U8945 ( .A1(n8532), .A2(n10047), .B1(n7141), .B2(n10022), .ZN(n7142) );
  AOI21_X1 U8946 ( .B1(n10038), .B2(P2_REG2_REG_1__SCAN_IN), .A(n7142), .ZN(
        n7144) );
  XNOR2_X1 U8947 ( .A(n7954), .B(n7824), .ZN(n10049) );
  NAND2_X1 U8948 ( .A1(n10049), .A2(n8536), .ZN(n7143) );
  OAI211_X1 U8949 ( .C1(n10046), .C2(n10038), .A(n7144), .B(n7143), .ZN(
        P2_U3232) );
  INV_X1 U8950 ( .A(n7145), .ZN(n7205) );
  INV_X1 U8951 ( .A(n9227), .ZN(n9703) );
  OAI222_X1 U8952 ( .A1(n9572), .A2(n7205), .B1(n9703), .B2(P1_U3086), .C1(
        n7146), .C2(n9569), .ZN(P1_U3337) );
  OAI21_X1 U8953 ( .B1(n7148), .B2(n8928), .A(n7147), .ZN(n7150) );
  AOI21_X1 U8954 ( .B1(n7150), .B2(n9710), .A(n7149), .ZN(n9760) );
  OAI21_X1 U8955 ( .B1(n5642), .B2(n7152), .A(n7151), .ZN(n9763) );
  NAND2_X1 U8956 ( .A1(n9722), .A2(n7153), .ZN(n7157) );
  NAND2_X1 U8957 ( .A1(n9755), .A2(n7153), .ZN(n7154) );
  NAND2_X1 U8958 ( .A1(n9724), .A2(n7154), .ZN(n7155) );
  NOR2_X1 U8959 ( .A1(n7208), .A2(n7155), .ZN(n9758) );
  AOI22_X1 U8960 ( .A1(n9731), .A2(n9758), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n9733), .ZN(n7156) );
  OAI211_X1 U8961 ( .C1(n6663), .C2(n9409), .A(n7157), .B(n7156), .ZN(n7158)
         );
  AOI21_X1 U8962 ( .B1(n9741), .B2(n9763), .A(n7158), .ZN(n7159) );
  OAI21_X1 U8963 ( .B1(n9744), .B2(n9760), .A(n7159), .ZN(P1_U3292) );
  NAND2_X1 U8964 ( .A1(n8297), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7160) );
  OAI21_X1 U8965 ( .B1(n8062), .B2(n8297), .A(n7160), .ZN(P2_U3520) );
  INV_X1 U8966 ( .A(n7161), .ZN(n7162) );
  XNOR2_X1 U8967 ( .A(n8052), .B(n7169), .ZN(n7237) );
  XNOR2_X1 U8968 ( .A(n7237), .B(n7245), .ZN(n7163) );
  AND3_X1 U8969 ( .A1(n7164), .A2(n7163), .A3(n7162), .ZN(n7165) );
  OAI21_X1 U8970 ( .B1(n7236), .B2(n7165), .A(n7238), .ZN(n7171) );
  AND2_X1 U8971 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10151) );
  AOI21_X1 U8972 ( .B1(n8187), .B2(n8240), .A(n10151), .ZN(n7166) );
  OAI21_X1 U8973 ( .B1(n7167), .B2(n8190), .A(n7166), .ZN(n7168) );
  AOI21_X1 U8974 ( .B1(n7169), .B2(n8192), .A(n7168), .ZN(n7170) );
  OAI211_X1 U8975 ( .C1(n7172), .C2(n8214), .A(n7171), .B(n7170), .ZN(P2_U3167) );
  OAI21_X1 U8976 ( .B1(n7175), .B2(n7174), .A(n7173), .ZN(n7176) );
  NAND2_X1 U8977 ( .A1(n7176), .A2(n8775), .ZN(n7181) );
  NAND2_X1 U8978 ( .A1(n9095), .A2(n9066), .ZN(n7178) );
  NAND2_X1 U8979 ( .A1(n9093), .A2(n8777), .ZN(n7177) );
  AND2_X1 U8980 ( .A1(n7178), .A2(n7177), .ZN(n7191) );
  NAND2_X1 U8981 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9182) );
  OAI21_X1 U8982 ( .B1(n8780), .B2(n7191), .A(n9182), .ZN(n7179) );
  AOI21_X1 U8983 ( .B1(n7198), .B2(n8782), .A(n7179), .ZN(n7180) );
  OAI211_X1 U8984 ( .C1(n9772), .C2(n8785), .A(n7181), .B(n7180), .ZN(P1_U3213) );
  NOR2_X1 U8985 ( .A1(n7183), .A2(n7182), .ZN(n7184) );
  OR2_X1 U8986 ( .A1(n7185), .A2(n7184), .ZN(n9774) );
  INV_X1 U8987 ( .A(n7737), .ZN(n9719) );
  AND2_X1 U8988 ( .A1(n7186), .A2(n9022), .ZN(n8799) );
  NAND2_X1 U8989 ( .A1(n7187), .A2(n8799), .ZN(n7188) );
  NAND2_X1 U8990 ( .A1(n7188), .A2(n8802), .ZN(n7189) );
  NAND2_X1 U8991 ( .A1(n7189), .A2(n8806), .ZN(n7283) );
  OAI21_X1 U8992 ( .B1(n7189), .B2(n8806), .A(n7283), .ZN(n7190) );
  NAND2_X1 U8993 ( .A1(n7190), .A2(n9710), .ZN(n7192) );
  NAND2_X1 U8994 ( .A1(n7192), .A2(n7191), .ZN(n7193) );
  AOI21_X1 U8995 ( .B1(n9774), .B2(n9719), .A(n7193), .ZN(n9776) );
  NOR2_X1 U8996 ( .A1(n9721), .A2(n7194), .ZN(n9728) );
  NAND2_X1 U8997 ( .A1(n7195), .A2(n7199), .ZN(n7196) );
  NAND2_X1 U8998 ( .A1(n7196), .A2(n9724), .ZN(n7197) );
  OR2_X1 U8999 ( .A1(n7197), .A2(n7286), .ZN(n9771) );
  INV_X1 U9000 ( .A(n9731), .ZN(n9370) );
  AOI22_X1 U9001 ( .A1(n9744), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7198), .B2(
        n9733), .ZN(n7201) );
  NAND2_X1 U9002 ( .A1(n9722), .A2(n7199), .ZN(n7200) );
  OAI211_X1 U9003 ( .C1(n9771), .C2(n9370), .A(n7201), .B(n7200), .ZN(n7202)
         );
  AOI21_X1 U9004 ( .B1(n9774), .B2(n9728), .A(n7202), .ZN(n7203) );
  OAI21_X1 U9005 ( .B1(n9776), .B2(n9721), .A(n7203), .ZN(P1_U3286) );
  INV_X1 U9006 ( .A(n8340), .ZN(n8344) );
  OAI222_X1 U9007 ( .A1(P2_U3151), .A2(n8344), .B1(n6582), .B2(n7205), .C1(
        n7204), .C2(n8668), .ZN(P2_U3277) );
  XNOR2_X1 U9008 ( .A(n7207), .B(n7206), .ZN(n9769) );
  OAI211_X1 U9009 ( .C1(n7208), .C2(n9766), .A(n6803), .B(n9724), .ZN(n9764)
         );
  OAI22_X1 U9010 ( .A1(n9737), .A2(n9766), .B1(n9370), .B2(n9764), .ZN(n7215)
         );
  INV_X1 U9011 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9115) );
  NAND2_X1 U9012 ( .A1(n9769), .A2(n9719), .ZN(n7212) );
  XNOR2_X1 U9013 ( .A(n8930), .B(n7209), .ZN(n7211) );
  AOI21_X1 U9014 ( .B1(n7211), .B2(n9710), .A(n7210), .ZN(n9765) );
  OAI211_X1 U9015 ( .C1(n9405), .C2(n9115), .A(n7212), .B(n9765), .ZN(n7213)
         );
  MUX2_X1 U9016 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n7213), .S(n9409), .Z(n7214)
         );
  AOI211_X1 U9017 ( .C1(n9769), .C2(n9728), .A(n7215), .B(n7214), .ZN(n7216)
         );
  INV_X1 U9018 ( .A(n7216), .ZN(P1_U3291) );
  INV_X1 U9019 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7228) );
  INV_X1 U9020 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7223) );
  NAND2_X1 U9021 ( .A1(n7218), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7222) );
  INV_X1 U9022 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7219) );
  OR2_X1 U9023 ( .A1(n7220), .A2(n7219), .ZN(n7221) );
  OAI211_X1 U9024 ( .C1(n7217), .C2(n7223), .A(n7222), .B(n7221), .ZN(n7224)
         );
  INV_X1 U9025 ( .A(n7224), .ZN(n7225) );
  NAND2_X1 U9026 ( .A1(n7226), .A2(n7225), .ZN(n8360) );
  NAND2_X1 U9027 ( .A1(n8360), .A2(P2_U3893), .ZN(n7227) );
  OAI21_X1 U9028 ( .B1(P2_U3893), .B2(n7228), .A(n7227), .ZN(P2_U3522) );
  OAI22_X1 U9029 ( .A1(n8532), .A2(n7230), .B1(n7229), .B2(n10022), .ZN(n7233)
         );
  MUX2_X1 U9030 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7231), .S(n10035), .Z(n7232)
         );
  AOI211_X1 U9031 ( .C1(n8536), .C2(n7234), .A(n7233), .B(n7232), .ZN(n7235)
         );
  INV_X1 U9032 ( .A(n7235), .ZN(P2_U3229) );
  XNOR2_X1 U9033 ( .A(n10062), .B(n8052), .ZN(n7308) );
  XOR2_X1 U9034 ( .A(n8240), .B(n7308), .Z(n7239) );
  OAI211_X1 U9035 ( .C1(n4588), .C2(n7239), .A(n7309), .B(n7238), .ZN(n7248)
         );
  INV_X1 U9036 ( .A(n7240), .ZN(n7241) );
  AOI21_X1 U9037 ( .B1(n8187), .B2(n8239), .A(n7241), .ZN(n7244) );
  INV_X1 U9038 ( .A(n7242), .ZN(n7274) );
  NAND2_X1 U9039 ( .A1(n8199), .A2(n7274), .ZN(n7243) );
  OAI211_X1 U9040 ( .C1(n7245), .C2(n8190), .A(n7244), .B(n7243), .ZN(n7246)
         );
  AOI21_X1 U9041 ( .B1(n7275), .B2(n8192), .A(n7246), .ZN(n7247) );
  NAND2_X1 U9042 ( .A1(n7248), .A2(n7247), .ZN(P2_U3179) );
  INV_X1 U9043 ( .A(n7249), .ZN(n7259) );
  INV_X1 U9044 ( .A(n7250), .ZN(n7251) );
  MUX2_X1 U9045 ( .A(n6672), .B(n7251), .S(n9409), .Z(n7258) );
  INV_X1 U9046 ( .A(n7252), .ZN(n7253) );
  OAI22_X1 U9047 ( .A1(n9737), .A2(n7254), .B1(n7253), .B2(n9405), .ZN(n7255)
         );
  AOI21_X1 U9048 ( .B1(n7256), .B2(n9731), .A(n7255), .ZN(n7257) );
  OAI211_X1 U9049 ( .C1(n7259), .C2(n9430), .A(n7258), .B(n7257), .ZN(P1_U3287) );
  INV_X1 U9050 ( .A(n7260), .ZN(n7269) );
  INV_X1 U9051 ( .A(n7261), .ZN(n7262) );
  MUX2_X1 U9052 ( .A(n6670), .B(n7262), .S(n9409), .Z(n7268) );
  OAI22_X1 U9053 ( .A1(n9737), .A2(n7264), .B1(n9405), .B2(n7263), .ZN(n7265)
         );
  AOI21_X1 U9054 ( .B1(n7266), .B2(n9731), .A(n7265), .ZN(n7267) );
  OAI211_X1 U9055 ( .C1(n7269), .C2(n9430), .A(n7268), .B(n7267), .ZN(P1_U3288) );
  XNOR2_X1 U9056 ( .A(n7270), .B(n7959), .ZN(n10060) );
  XOR2_X1 U9057 ( .A(n7959), .B(n7271), .Z(n7272) );
  AOI222_X1 U9058 ( .A1(n8516), .A2(n7272), .B1(n8239), .B2(n8511), .C1(n8241), 
        .C2(n8513), .ZN(n10061) );
  MUX2_X1 U9059 ( .A(n7273), .B(n10061), .S(n10035), .Z(n7277) );
  AOI22_X1 U9060 ( .A1(n8519), .A2(n7275), .B1(n8505), .B2(n7274), .ZN(n7276)
         );
  OAI211_X1 U9061 ( .C1(n7546), .C2(n10060), .A(n7277), .B(n7276), .ZN(
        P2_U3227) );
  AOI21_X1 U9062 ( .B1(n7279), .B2(n7280), .A(n7278), .ZN(n7367) );
  INV_X1 U9063 ( .A(n9728), .ZN(n7292) );
  AOI22_X1 U9064 ( .A1(n9066), .A2(n9094), .B1(n9092), .B2(n8777), .ZN(n7326)
         );
  INV_X1 U9065 ( .A(n7280), .ZN(n7281) );
  AOI21_X1 U9066 ( .B1(n7283), .B2(n7282), .A(n7281), .ZN(n7342) );
  AND3_X1 U9067 ( .A1(n7283), .A2(n7282), .A3(n7281), .ZN(n7284) );
  OAI21_X1 U9068 ( .B1(n7342), .B2(n7284), .A(n9710), .ZN(n7285) );
  OAI211_X1 U9069 ( .C1(n7367), .C2(n7737), .A(n7326), .B(n7285), .ZN(n7368)
         );
  NAND2_X1 U9070 ( .A1(n7368), .A2(n9409), .ZN(n7291) );
  INV_X1 U9071 ( .A(n7286), .ZN(n7287) );
  AOI211_X1 U9072 ( .C1(n7375), .C2(n7287), .A(n9422), .B(n7349), .ZN(n7369)
         );
  AOI22_X1 U9073 ( .A1(n9744), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7328), .B2(
        n9733), .ZN(n7288) );
  OAI21_X1 U9074 ( .B1(n9737), .B2(n7372), .A(n7288), .ZN(n7289) );
  AOI21_X1 U9075 ( .B1(n7369), .B2(n9731), .A(n7289), .ZN(n7290) );
  OAI211_X1 U9076 ( .C1(n7367), .C2(n7292), .A(n7291), .B(n7290), .ZN(P1_U3285) );
  NAND2_X1 U9077 ( .A1(n7293), .A2(n7857), .ZN(n7294) );
  NAND2_X1 U9078 ( .A1(n7294), .A2(n7859), .ZN(n7333) );
  OAI21_X1 U9079 ( .B1(n7294), .B2(n7859), .A(n7333), .ZN(n10068) );
  NAND2_X1 U9080 ( .A1(n10035), .A2(n7295), .ZN(n8373) );
  INV_X1 U9081 ( .A(n7296), .ZN(n7302) );
  OAI21_X1 U9082 ( .B1(n7298), .B2(n7961), .A(n7297), .ZN(n7300) );
  OAI22_X1 U9083 ( .A1(n7318), .A2(n10031), .B1(n7563), .B2(n10032), .ZN(n7299) );
  AOI21_X1 U9084 ( .B1(n7300), .B2(n8516), .A(n7299), .ZN(n7301) );
  OAI21_X1 U9085 ( .B1(n10068), .B2(n7302), .A(n7301), .ZN(n10070) );
  NAND2_X1 U9086 ( .A1(n10070), .A2(n10035), .ZN(n7305) );
  INV_X1 U9087 ( .A(n10066), .ZN(n7320) );
  OAI22_X1 U9088 ( .A1(n10035), .A2(n5848), .B1(n7314), .B2(n10022), .ZN(n7303) );
  AOI21_X1 U9089 ( .B1(n8519), .B2(n7320), .A(n7303), .ZN(n7304) );
  OAI211_X1 U9090 ( .C1(n10068), .C2(n8373), .A(n7305), .B(n7304), .ZN(
        P2_U3226) );
  INV_X1 U9091 ( .A(n7306), .ZN(n8006) );
  OAI222_X1 U9092 ( .A1(P2_U3151), .A2(n8353), .B1(n6582), .B2(n8006), .C1(
        n7307), .C2(n8668), .ZN(P2_U3276) );
  INV_X1 U9093 ( .A(n7308), .ZN(n7310) );
  OAI21_X1 U9094 ( .B1(n7318), .B2(n7310), .A(n7309), .ZN(n7313) );
  XNOR2_X1 U9095 ( .A(n8056), .B(n10066), .ZN(n7311) );
  NAND2_X1 U9096 ( .A1(n7311), .A2(n7487), .ZN(n7488) );
  OAI21_X1 U9097 ( .B1(n7311), .B2(n7487), .A(n7488), .ZN(n7312) );
  AOI21_X1 U9098 ( .B1(n7313), .B2(n7312), .A(n7491), .ZN(n7322) );
  AND2_X1 U9099 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9842) );
  AOI21_X1 U9100 ( .B1(n8187), .B2(n8238), .A(n9842), .ZN(n7317) );
  INV_X1 U9101 ( .A(n7314), .ZN(n7315) );
  NAND2_X1 U9102 ( .A1(n8199), .A2(n7315), .ZN(n7316) );
  OAI211_X1 U9103 ( .C1(n7318), .C2(n8190), .A(n7317), .B(n7316), .ZN(n7319)
         );
  AOI21_X1 U9104 ( .B1(n7320), .B2(n8192), .A(n7319), .ZN(n7321) );
  OAI21_X1 U9105 ( .B1(n7322), .B2(n8206), .A(n7321), .ZN(P2_U3153) );
  NAND2_X1 U9106 ( .A1(n7173), .A2(n7323), .ZN(n7432) );
  XNOR2_X1 U9107 ( .A(n7432), .B(n7433), .ZN(n7325) );
  NOR2_X1 U9108 ( .A1(n7325), .A2(n7324), .ZN(n7431) );
  AOI21_X1 U9109 ( .B1(n7325), .B2(n7324), .A(n7431), .ZN(n7331) );
  NOR2_X1 U9110 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5174), .ZN(n9195) );
  NOR2_X1 U9111 ( .A1(n8780), .A2(n7326), .ZN(n7327) );
  AOI211_X1 U9112 ( .C1(n8782), .C2(n7328), .A(n9195), .B(n7327), .ZN(n7330)
         );
  NAND2_X1 U9113 ( .A1(n8767), .A2(n7375), .ZN(n7329) );
  OAI211_X1 U9114 ( .C1(n7331), .C2(n8769), .A(n7330), .B(n7329), .ZN(P1_U3221) );
  NAND2_X1 U9115 ( .A1(n7333), .A2(n7332), .ZN(n7334) );
  XNOR2_X1 U9116 ( .A(n7495), .B(n8238), .ZN(n7963) );
  XNOR2_X1 U9117 ( .A(n7334), .B(n7963), .ZN(n10073) );
  XOR2_X1 U9118 ( .A(n7963), .B(n7335), .Z(n7336) );
  AOI222_X1 U9119 ( .A1(n8516), .A2(n7336), .B1(n8237), .B2(n8511), .C1(n8239), 
        .C2(n8513), .ZN(n10071) );
  MUX2_X1 U9120 ( .A(n7337), .B(n10071), .S(n10035), .Z(n7340) );
  INV_X1 U9121 ( .A(n7338), .ZN(n7484) );
  AOI22_X1 U9122 ( .A1(n8519), .A2(n7495), .B1(n8505), .B2(n7484), .ZN(n7339)
         );
  OAI211_X1 U9123 ( .C1(n7546), .C2(n10073), .A(n7340), .B(n7339), .ZN(
        P2_U3225) );
  NOR2_X1 U9124 ( .A1(n7342), .A2(n7341), .ZN(n7343) );
  XOR2_X1 U9125 ( .A(n7347), .B(n7343), .Z(n7345) );
  NAND2_X1 U9126 ( .A1(n9093), .A2(n9066), .ZN(n7437) );
  INV_X1 U9127 ( .A(n7437), .ZN(n7344) );
  AOI21_X1 U9128 ( .B1(n7345), .B2(n9710), .A(n7344), .ZN(n7357) );
  AOI21_X1 U9129 ( .B1(n7348), .B2(n7347), .A(n7346), .ZN(n7358) );
  INV_X1 U9130 ( .A(n7358), .ZN(n7354) );
  OAI211_X1 U9131 ( .C1(n7444), .C2(n7349), .A(n7420), .B(n9724), .ZN(n7350)
         );
  NAND2_X1 U9132 ( .A1(n9091), .A2(n8777), .ZN(n7438) );
  AND2_X1 U9133 ( .A1(n7350), .A2(n7438), .ZN(n7356) );
  AOI22_X1 U9134 ( .A1(n9744), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7441), .B2(
        n9733), .ZN(n7352) );
  NAND2_X1 U9135 ( .A1(n9722), .A2(n7359), .ZN(n7351) );
  OAI211_X1 U9136 ( .C1(n7356), .C2(n9370), .A(n7352), .B(n7351), .ZN(n7353)
         );
  AOI21_X1 U9137 ( .B1(n7354), .B2(n9741), .A(n7353), .ZN(n7355) );
  OAI21_X1 U9138 ( .B1(n9744), .B2(n7357), .A(n7355), .ZN(P1_U3284) );
  INV_X1 U9139 ( .A(n9768), .ZN(n9751) );
  OAI211_X1 U9140 ( .C1(n7358), .C2(n9751), .A(n7357), .B(n7356), .ZN(n7364)
         );
  INV_X1 U9141 ( .A(n7364), .ZN(n7361) );
  AOI22_X1 U9142 ( .A1(n6562), .A2(n7359), .B1(n9786), .B2(
        P1_REG0_REG_9__SCAN_IN), .ZN(n7360) );
  OAI21_X1 U9143 ( .B1(n7361), .B2(n9786), .A(n7360), .ZN(P1_U3480) );
  INV_X1 U9144 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7362) );
  OAI22_X1 U9145 ( .A1(n7444), .A2(n9469), .B1(n9797), .B2(n7362), .ZN(n7363)
         );
  AOI21_X1 U9146 ( .B1(n7364), .B2(n9797), .A(n7363), .ZN(n7365) );
  INV_X1 U9147 ( .A(n7365), .ZN(P1_U3531) );
  INV_X1 U9148 ( .A(n7366), .ZN(n9785) );
  INV_X1 U9149 ( .A(n7367), .ZN(n7370) );
  AOI211_X1 U9150 ( .C1(n9785), .C2(n7370), .A(n7369), .B(n7368), .ZN(n7377)
         );
  INV_X1 U9151 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7371) );
  OAI22_X1 U9152 ( .A1(n9543), .A2(n7372), .B1(n9788), .B2(n7371), .ZN(n7373)
         );
  INV_X1 U9153 ( .A(n7373), .ZN(n7374) );
  OAI21_X1 U9154 ( .B1(n7377), .B2(n9786), .A(n7374), .ZN(P1_U3477) );
  AOI22_X1 U9155 ( .A1(n6572), .A2(n7375), .B1(n9795), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n7376) );
  OAI21_X1 U9156 ( .B1(n7377), .B2(n9795), .A(n7376), .ZN(P1_U3530) );
  XNOR2_X1 U9157 ( .A(n7447), .B(n7960), .ZN(n7378) );
  AOI222_X1 U9158 ( .A1(n8516), .A2(n7378), .B1(n8236), .B2(n8511), .C1(n8238), 
        .C2(n8513), .ZN(n7457) );
  INV_X1 U9159 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9881) );
  OAI22_X1 U9160 ( .A1(n10035), .A2(n9881), .B1(n7559), .B2(n10022), .ZN(n7381) );
  XNOR2_X1 U9161 ( .A(n7379), .B(n7960), .ZN(n7458) );
  NOR2_X1 U9162 ( .A1(n7458), .A2(n7546), .ZN(n7380) );
  AOI211_X1 U9163 ( .C1(n8519), .C2(n7572), .A(n7381), .B(n7380), .ZN(n7382)
         );
  OAI21_X1 U9164 ( .B1(n10038), .B2(n7457), .A(n7382), .ZN(P2_U3224) );
  INV_X1 U9165 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10419) );
  NOR2_X1 U9166 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7383) );
  AOI21_X1 U9167 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7383), .ZN(n10116) );
  NOR2_X1 U9168 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7384) );
  AOI21_X1 U9169 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7384), .ZN(n10119) );
  NOR2_X1 U9170 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7385) );
  AOI21_X1 U9171 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7385), .ZN(n10122) );
  NOR2_X1 U9172 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7386) );
  AOI21_X1 U9173 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7386), .ZN(n10125) );
  NOR2_X1 U9174 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7387) );
  AOI21_X1 U9175 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7387), .ZN(n10128) );
  NOR2_X1 U9176 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7388) );
  AOI21_X1 U9177 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7388), .ZN(n10131) );
  INV_X1 U9178 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10322) );
  INV_X1 U9179 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9588) );
  NAND2_X1 U9180 ( .A1(n10322), .A2(n9588), .ZN(n10136) );
  NOR2_X1 U9181 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7394) );
  INV_X1 U9182 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10307) );
  XOR2_X1 U9183 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n10307), .Z(n10559) );
  NAND2_X1 U9184 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7392) );
  INV_X1 U9185 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9129) );
  XNOR2_X1 U9186 ( .A(n9129), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(n10557) );
  NAND2_X1 U9187 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7390) );
  XOR2_X1 U9188 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10555) );
  AOI21_X1 U9189 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10106) );
  NAND3_X1 U9190 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10108) );
  OAI21_X1 U9191 ( .B1(n10106), .B2(n10284), .A(n10108), .ZN(n10554) );
  NAND2_X1 U9192 ( .A1(n10555), .A2(n10554), .ZN(n7389) );
  NAND2_X1 U9193 ( .A1(n7390), .A2(n7389), .ZN(n10556) );
  NAND2_X1 U9194 ( .A1(n10557), .A2(n10556), .ZN(n7391) );
  NAND2_X1 U9195 ( .A1(n7392), .A2(n7391), .ZN(n10558) );
  NOR2_X1 U9196 ( .A1(n10559), .A2(n10558), .ZN(n7393) );
  NOR2_X1 U9197 ( .A1(n7394), .A2(n7393), .ZN(n7395) );
  NOR2_X1 U9198 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7395), .ZN(n10549) );
  AND2_X1 U9199 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7395), .ZN(n10548) );
  NOR2_X1 U9200 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10548), .ZN(n7396) );
  NOR2_X1 U9201 ( .A1(n10549), .A2(n7396), .ZN(n7397) );
  NAND2_X1 U9202 ( .A1(n7397), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7399) );
  INV_X1 U9203 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9167) );
  XNOR2_X1 U9204 ( .A(n7397), .B(n9167), .ZN(n10547) );
  NAND2_X1 U9205 ( .A1(n10547), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7398) );
  NAND2_X1 U9206 ( .A1(n7399), .A2(n7398), .ZN(n7400) );
  NAND2_X1 U9207 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7400), .ZN(n7403) );
  INV_X1 U9208 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7401) );
  XNOR2_X1 U9209 ( .A(n7401), .B(n7400), .ZN(n10552) );
  NAND2_X1 U9210 ( .A1(n10552), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7402) );
  NAND2_X1 U9211 ( .A1(n7403), .A2(n7402), .ZN(n7404) );
  NAND2_X1 U9212 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7404), .ZN(n7406) );
  XOR2_X1 U9213 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7404), .Z(n10553) );
  NAND2_X1 U9214 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10553), .ZN(n7405) );
  NAND2_X1 U9215 ( .A1(n7406), .A2(n7405), .ZN(n7407) );
  NAND2_X1 U9216 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n7407), .ZN(n7409) );
  XOR2_X1 U9217 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n7407), .Z(n10551) );
  NAND2_X1 U9218 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10551), .ZN(n7408) );
  NAND2_X1 U9219 ( .A1(n7409), .A2(n7408), .ZN(n10137) );
  AOI22_X1 U9220 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .B1(n10136), .B2(n10137), .ZN(n10134) );
  NAND2_X1 U9221 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7410) );
  OAI21_X1 U9222 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7410), .ZN(n10133) );
  NOR2_X1 U9223 ( .A1(n10134), .A2(n10133), .ZN(n10132) );
  AOI21_X1 U9224 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10132), .ZN(n10130) );
  NAND2_X1 U9225 ( .A1(n10131), .A2(n10130), .ZN(n10129) );
  OAI21_X1 U9226 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10129), .ZN(n10127) );
  NAND2_X1 U9227 ( .A1(n10128), .A2(n10127), .ZN(n10126) );
  OAI21_X1 U9228 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10126), .ZN(n10124) );
  NAND2_X1 U9229 ( .A1(n10125), .A2(n10124), .ZN(n10123) );
  OAI21_X1 U9230 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10123), .ZN(n10121) );
  NAND2_X1 U9231 ( .A1(n10122), .A2(n10121), .ZN(n10120) );
  OAI21_X1 U9232 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10120), .ZN(n10118) );
  NAND2_X1 U9233 ( .A1(n10119), .A2(n10118), .ZN(n10117) );
  OAI21_X1 U9234 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10117), .ZN(n10115) );
  NAND2_X1 U9235 ( .A1(n10116), .A2(n10115), .ZN(n10114) );
  OAI21_X1 U9236 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10114), .ZN(n10112) );
  NAND2_X1 U9237 ( .A1(n10419), .A2(n10112), .ZN(n7411) );
  NOR2_X1 U9238 ( .A1(n10419), .A2(n10112), .ZN(n10111) );
  AOI21_X1 U9239 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7411), .A(n10111), .ZN(
        n7413) );
  XNOR2_X1 U9240 ( .A(n5069), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7412) );
  XNOR2_X1 U9241 ( .A(n7413), .B(n7412), .ZN(ADD_1068_U4) );
  INV_X1 U9242 ( .A(n7414), .ZN(n7446) );
  INV_X1 U9243 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7415) );
  OAI222_X1 U9244 ( .A1(n9572), .A2(n7446), .B1(P1_U3086), .B2(n7416), .C1(
        n7415), .C2(n9569), .ZN(P1_U3335) );
  AOI21_X1 U9245 ( .B1(n7418), .B2(n8937), .A(n7417), .ZN(n7519) );
  INV_X1 U9246 ( .A(n7419), .ZN(n9726) );
  AOI211_X1 U9247 ( .C1(n7524), .C2(n7420), .A(n9422), .B(n9726), .ZN(n7521)
         );
  NOR2_X1 U9248 ( .A1(n4767), .A2(n9737), .ZN(n7422) );
  OAI22_X1 U9249 ( .A1(n9409), .A2(n6710), .B1(n7467), .B2(n9405), .ZN(n7421)
         );
  AOI211_X1 U9250 ( .C1(n7521), .C2(n9731), .A(n7422), .B(n7421), .ZN(n7430)
         );
  INV_X1 U9251 ( .A(n9714), .ZN(n7424) );
  AOI21_X1 U9252 ( .B1(n9035), .B2(n9032), .A(n8937), .ZN(n7423) );
  OAI21_X1 U9253 ( .B1(n7424), .B2(n7423), .A(n9710), .ZN(n7428) );
  NAND2_X1 U9254 ( .A1(n9092), .A2(n9066), .ZN(n7426) );
  NAND2_X1 U9255 ( .A1(n9090), .A2(n8777), .ZN(n7425) );
  NAND2_X1 U9256 ( .A1(n7426), .A2(n7425), .ZN(n7465) );
  INV_X1 U9257 ( .A(n7465), .ZN(n7427) );
  NAND2_X1 U9258 ( .A1(n7428), .A2(n7427), .ZN(n7520) );
  NAND2_X1 U9259 ( .A1(n7520), .A2(n9409), .ZN(n7429) );
  OAI211_X1 U9260 ( .C1(n7519), .C2(n9430), .A(n7430), .B(n7429), .ZN(P1_U3283) );
  AOI21_X1 U9261 ( .B1(n7433), .B2(n7432), .A(n7431), .ZN(n7436) );
  OAI211_X1 U9262 ( .C1(n7436), .C2(n7435), .A(n8775), .B(n7434), .ZN(n7443)
         );
  AOI21_X1 U9263 ( .B1(n7438), .B2(n7437), .A(n8780), .ZN(n7439) );
  AOI211_X1 U9264 ( .C1(n8782), .C2(n7441), .A(n7440), .B(n7439), .ZN(n7442)
         );
  OAI211_X1 U9265 ( .C1(n7444), .C2(n8785), .A(n7443), .B(n7442), .ZN(P1_U3231) );
  INV_X1 U9266 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7445) );
  OAI222_X1 U9267 ( .A1(n7948), .A2(P2_U3151), .B1(n6582), .B2(n7446), .C1(
        n7445), .C2(n8668), .ZN(P2_U3275) );
  NAND2_X1 U9268 ( .A1(n7447), .A2(n7960), .ZN(n7449) );
  NAND2_X1 U9269 ( .A1(n7449), .A2(n7448), .ZN(n7500) );
  INV_X1 U9270 ( .A(n7499), .ZN(n7965) );
  XNOR2_X1 U9271 ( .A(n7500), .B(n7965), .ZN(n7450) );
  OAI222_X1 U9272 ( .A1(n10032), .A2(n8118), .B1(n10031), .B2(n7606), .C1(
        n10041), .C2(n7450), .ZN(n7476) );
  INV_X1 U9273 ( .A(n7476), .ZN(n7456) );
  OAI22_X1 U9274 ( .A1(n10035), .A2(n7451), .B1(n7602), .B2(n10022), .ZN(n7452) );
  AOI21_X1 U9275 ( .B1(n8519), .B2(n7608), .A(n7452), .ZN(n7455) );
  XNOR2_X1 U9276 ( .A(n7499), .B(n7453), .ZN(n7477) );
  NAND2_X1 U9277 ( .A1(n7477), .A2(n8536), .ZN(n7454) );
  OAI211_X1 U9278 ( .C1(n7456), .C2(n10038), .A(n7455), .B(n7454), .ZN(
        P2_U3223) );
  INV_X1 U9279 ( .A(n10082), .ZN(n10084) );
  OAI21_X1 U9280 ( .B1(n10084), .B2(n7458), .A(n7457), .ZN(n7471) );
  INV_X1 U9281 ( .A(n7471), .ZN(n7460) );
  INV_X1 U9282 ( .A(n8662), .ZN(n8609) );
  AOI22_X1 U9283 ( .A1(n8609), .A2(n7572), .B1(n10093), .B2(
        P2_REG0_REG_9__SCAN_IN), .ZN(n7459) );
  OAI21_X1 U9284 ( .B1(n7460), .B2(n10093), .A(n7459), .ZN(P2_U3417) );
  NAND2_X1 U9285 ( .A1(n7461), .A2(n7462), .ZN(n7463) );
  XOR2_X1 U9286 ( .A(n7464), .B(n7463), .Z(n7470) );
  AOI22_X1 U9287 ( .A1(n8763), .A2(n7465), .B1(P1_REG3_REG_10__SCAN_IN), .B2(
        P1_U3086), .ZN(n7466) );
  OAI21_X1 U9288 ( .B1(n7467), .B2(n8765), .A(n7466), .ZN(n7468) );
  AOI21_X1 U9289 ( .B1(n7524), .B2(n8767), .A(n7468), .ZN(n7469) );
  OAI21_X1 U9290 ( .B1(n7470), .B2(n8769), .A(n7469), .ZN(P1_U3217) );
  NAND2_X1 U9291 ( .A1(n7471), .A2(n10105), .ZN(n7473) );
  NAND2_X1 U9292 ( .A1(n8539), .A2(n7572), .ZN(n7472) );
  OAI211_X1 U9293 ( .C1(n10105), .C2(n5872), .A(n7473), .B(n7472), .ZN(
        P2_U3468) );
  INV_X1 U9294 ( .A(n7474), .ZN(n7497) );
  OAI222_X1 U9295 ( .A1(n9572), .A2(n7497), .B1(P1_U3086), .B2(n9023), .C1(
        n7475), .C2(n9569), .ZN(P1_U3334) );
  AOI21_X1 U9296 ( .B1(n10082), .B2(n7477), .A(n7476), .ZN(n7482) );
  INV_X1 U9297 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7478) );
  NOR2_X1 U9298 ( .A1(n10091), .A2(n7478), .ZN(n7479) );
  AOI21_X1 U9299 ( .B1(n8609), .B2(n7608), .A(n7479), .ZN(n7480) );
  OAI21_X1 U9300 ( .B1(n7482), .B2(n10093), .A(n7480), .ZN(P2_U3420) );
  AOI22_X1 U9301 ( .A1(n7608), .A2(n8539), .B1(n10103), .B2(
        P2_REG1_REG_10__SCAN_IN), .ZN(n7481) );
  OAI21_X1 U9302 ( .B1(n7482), .B2(n10103), .A(n7481), .ZN(P2_U3469) );
  INV_X1 U9303 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7483) );
  NOR2_X1 U9304 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7483), .ZN(n9854) );
  AOI21_X1 U9305 ( .B1(n8187), .B2(n8237), .A(n9854), .ZN(n7486) );
  NAND2_X1 U9306 ( .A1(n8199), .A2(n7484), .ZN(n7485) );
  OAI211_X1 U9307 ( .C1(n7487), .C2(n8190), .A(n7486), .B(n7485), .ZN(n7494)
         );
  INV_X1 U9308 ( .A(n7488), .ZN(n7490) );
  XNOR2_X1 U9309 ( .A(n7495), .B(n8052), .ZN(n7564) );
  XNOR2_X1 U9310 ( .A(n7564), .B(n8238), .ZN(n7489) );
  OAI21_X1 U9311 ( .B1(n7491), .B2(n7490), .A(n7489), .ZN(n7565) );
  OR3_X1 U9312 ( .A1(n7491), .A2(n7490), .A3(n7489), .ZN(n7492) );
  AOI21_X1 U9313 ( .B1(n7565), .B2(n7492), .A(n8206), .ZN(n7493) );
  AOI211_X1 U9314 ( .C1(n7495), .C2(n8192), .A(n7494), .B(n7493), .ZN(n7496)
         );
  INV_X1 U9315 ( .A(n7496), .ZN(P2_U3161) );
  OAI222_X1 U9316 ( .A1(n7498), .A2(P2_U3151), .B1(n6582), .B2(n7497), .C1(
        n10376), .C2(n8668), .ZN(P2_U3274) );
  NAND2_X1 U9317 ( .A1(n7500), .A2(n7499), .ZN(n7502) );
  NAND2_X1 U9318 ( .A1(n7502), .A2(n7501), .ZN(n7503) );
  XNOR2_X1 U9319 ( .A(n7503), .B(n7964), .ZN(n7504) );
  OAI222_X1 U9320 ( .A1(n10031), .A2(n7646), .B1(n10032), .B2(n9599), .C1(
        n10041), .C2(n7504), .ZN(n10079) );
  INV_X1 U9321 ( .A(n10079), .ZN(n7510) );
  OAI21_X1 U9322 ( .B1(n7506), .B2(n7964), .A(n7505), .ZN(n10081) );
  INV_X1 U9323 ( .A(n7639), .ZN(n10078) );
  NOR2_X1 U9324 ( .A1(n10078), .A2(n8532), .ZN(n7508) );
  OAI22_X1 U9325 ( .A1(n10035), .A2(n5897), .B1(n7643), .B2(n10022), .ZN(n7507) );
  AOI211_X1 U9326 ( .C1(n10081), .C2(n8536), .A(n7508), .B(n7507), .ZN(n7509)
         );
  OAI21_X1 U9327 ( .B1(n7510), .B2(n10038), .A(n7509), .ZN(P2_U3222) );
  AOI21_X1 U9328 ( .B1(n7511), .B2(n7514), .A(n7513), .ZN(n7518) );
  AOI22_X1 U9329 ( .A1(n9066), .A2(n9091), .B1(n9089), .B2(n8777), .ZN(n9715)
         );
  NAND2_X1 U9330 ( .A1(n8782), .A2(n9720), .ZN(n7515) );
  NAND2_X1 U9331 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9622) );
  OAI211_X1 U9332 ( .C1(n8780), .C2(n9715), .A(n7515), .B(n9622), .ZN(n7516)
         );
  AOI21_X1 U9333 ( .B1(n9723), .B2(n8767), .A(n7516), .ZN(n7517) );
  OAI21_X1 U9334 ( .B1(n7518), .B2(n8769), .A(n7517), .ZN(P1_U3236) );
  INV_X1 U9335 ( .A(n7519), .ZN(n7522) );
  AOI211_X1 U9336 ( .C1(n7522), .C2(n9768), .A(n7521), .B(n7520), .ZN(n7526)
         );
  AOI22_X1 U9337 ( .A1(n7524), .A2(n6572), .B1(n9795), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7523) );
  OAI21_X1 U9338 ( .B1(n7526), .B2(n9795), .A(n7523), .ZN(P1_U3532) );
  AOI22_X1 U9339 ( .A1(n7524), .A2(n6562), .B1(n9786), .B2(
        P1_REG0_REG_10__SCAN_IN), .ZN(n7525) );
  OAI21_X1 U9340 ( .B1(n7526), .B2(n9786), .A(n7525), .ZN(P1_U3483) );
  INV_X1 U9341 ( .A(n7527), .ZN(n7529) );
  NOR3_X1 U9342 ( .A1(n7513), .A2(n7529), .A3(n7528), .ZN(n7532) );
  INV_X1 U9343 ( .A(n7530), .ZN(n7531) );
  OAI21_X1 U9344 ( .B1(n7532), .B2(n7531), .A(n8775), .ZN(n7536) );
  AOI22_X1 U9345 ( .A1(n9066), .A2(n9090), .B1(n9088), .B2(n8777), .ZN(n7585)
         );
  OAI21_X1 U9346 ( .B1(n8780), .B2(n7585), .A(n7533), .ZN(n7534) );
  AOI21_X1 U9347 ( .B1(n7588), .B2(n8782), .A(n7534), .ZN(n7535) );
  OAI211_X1 U9348 ( .C1(n7591), .C2(n8785), .A(n7536), .B(n7535), .ZN(P1_U3224) );
  INV_X1 U9349 ( .A(n7505), .ZN(n7538) );
  OAI21_X1 U9350 ( .B1(n7538), .B2(n7537), .A(n7968), .ZN(n7540) );
  NAND2_X1 U9351 ( .A1(n7540), .A2(n7539), .ZN(n10085) );
  XOR2_X1 U9352 ( .A(n7968), .B(n7541), .Z(n7542) );
  AOI222_X1 U9353 ( .A1(n8516), .A2(n7542), .B1(n8233), .B2(n8511), .C1(n8235), 
        .C2(n8513), .ZN(n10086) );
  OAI21_X1 U9354 ( .B1(n8122), .B2(n10022), .A(n10086), .ZN(n7543) );
  NAND2_X1 U9355 ( .A1(n7543), .A2(n10035), .ZN(n7545) );
  AOI22_X1 U9356 ( .A1(n10089), .A2(n8519), .B1(P2_REG2_REG_12__SCAN_IN), .B2(
        n10038), .ZN(n7544) );
  OAI211_X1 U9357 ( .C1(n7546), .C2(n10085), .A(n7545), .B(n7544), .ZN(
        P2_U3221) );
  INV_X1 U9358 ( .A(n7547), .ZN(n7550) );
  OAI222_X1 U9359 ( .A1(n9569), .A2(n7548), .B1(n9572), .B2(n7550), .C1(n6255), 
        .C2(P1_U3086), .ZN(P1_U3333) );
  OAI222_X1 U9360 ( .A1(P2_U3151), .A2(n7551), .B1(n6582), .B2(n7550), .C1(
        n7549), .C2(n8668), .ZN(P2_U3273) );
  AND2_X1 U9361 ( .A1(n7895), .A2(n7896), .ZN(n7893) );
  INV_X1 U9362 ( .A(n7893), .ZN(n7969) );
  XNOR2_X1 U9363 ( .A(n7552), .B(n7969), .ZN(n7553) );
  OAI222_X1 U9364 ( .A1(n10032), .A2(n8527), .B1(n10031), .B2(n8081), .C1(
        n7553), .C2(n10041), .ZN(n8601) );
  INV_X1 U9365 ( .A(n8086), .ZN(n8663) );
  OAI22_X1 U9366 ( .A1(n8663), .A2(n10023), .B1(n8084), .B2(n10022), .ZN(n7554) );
  OAI21_X1 U9367 ( .B1(n8601), .B2(n7554), .A(n10035), .ZN(n7557) );
  XNOR2_X1 U9368 ( .A(n7555), .B(n7893), .ZN(n8602) );
  AOI22_X1 U9369 ( .A1(n8602), .A2(n8536), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n10038), .ZN(n7556) );
  NAND2_X1 U9370 ( .A1(n7557), .A2(n7556), .ZN(P2_U3219) );
  NAND2_X1 U9371 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n9885) );
  INV_X1 U9372 ( .A(n9885), .ZN(n7558) );
  AOI21_X1 U9373 ( .B1(n8187), .B2(n8236), .A(n7558), .ZN(n7562) );
  INV_X1 U9374 ( .A(n7559), .ZN(n7560) );
  NAND2_X1 U9375 ( .A1(n8199), .A2(n7560), .ZN(n7561) );
  OAI211_X1 U9376 ( .C1(n7563), .C2(n8190), .A(n7562), .B(n7561), .ZN(n7571)
         );
  XNOR2_X1 U9377 ( .A(n7572), .B(n6895), .ZN(n7595) );
  XNOR2_X1 U9378 ( .A(n7595), .B(n7606), .ZN(n7569) );
  INV_X1 U9379 ( .A(n7564), .ZN(n7566) );
  OAI21_X1 U9380 ( .B1(n7566), .B2(n8238), .A(n7565), .ZN(n7568) );
  INV_X1 U9381 ( .A(n7597), .ZN(n7567) );
  AOI211_X1 U9382 ( .C1(n7569), .C2(n7568), .A(n8206), .B(n7567), .ZN(n7570)
         );
  AOI211_X1 U9383 ( .C1(n7572), .C2(n8192), .A(n7571), .B(n7570), .ZN(n7573)
         );
  INV_X1 U9384 ( .A(n7573), .ZN(P2_U3171) );
  OAI21_X1 U9385 ( .B1(n7576), .B2(n7575), .A(n7574), .ZN(n7577) );
  NAND2_X1 U9386 ( .A1(n7577), .A2(n8775), .ZN(n7580) );
  AOI22_X1 U9387 ( .A1(n9066), .A2(n9089), .B1(n9087), .B2(n8777), .ZN(n7655)
         );
  NAND2_X1 U9388 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9634) );
  OAI21_X1 U9389 ( .B1(n8780), .B2(n7655), .A(n9634), .ZN(n7578) );
  AOI21_X1 U9390 ( .B1(n7660), .B2(n8782), .A(n7578), .ZN(n7579) );
  OAI211_X1 U9391 ( .C1(n8849), .C2(n8785), .A(n7580), .B(n7579), .ZN(P1_U3234) );
  XNOR2_X1 U9392 ( .A(n7581), .B(n7583), .ZN(n7618) );
  INV_X1 U9393 ( .A(n7618), .ZN(n7594) );
  OAI211_X1 U9394 ( .C1(n7584), .C2(n7583), .A(n7582), .B(n9710), .ZN(n7586)
         );
  NAND2_X1 U9395 ( .A1(n7586), .A2(n7585), .ZN(n7616) );
  INV_X1 U9396 ( .A(n7587), .ZN(n9725) );
  AOI211_X1 U9397 ( .C1(n7620), .C2(n9725), .A(n9422), .B(n7657), .ZN(n7617)
         );
  NAND2_X1 U9398 ( .A1(n7617), .A2(n9731), .ZN(n7590) );
  AOI22_X1 U9399 ( .A1(n9744), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7588), .B2(
        n9733), .ZN(n7589) );
  OAI211_X1 U9400 ( .C1(n7591), .C2(n9737), .A(n7590), .B(n7589), .ZN(n7592)
         );
  AOI21_X1 U9401 ( .B1(n9409), .B2(n7616), .A(n7592), .ZN(n7593) );
  OAI21_X1 U9402 ( .B1(n7594), .B2(n9430), .A(n7593), .ZN(P1_U3281) );
  XNOR2_X1 U9403 ( .A(n7608), .B(n8052), .ZN(n7598) );
  OAI21_X1 U9404 ( .B1(n7599), .B2(n7598), .A(n7638), .ZN(n7600) );
  INV_X1 U9405 ( .A(n7600), .ZN(n7610) );
  NAND2_X1 U9406 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9901) );
  INV_X1 U9407 ( .A(n9901), .ZN(n7601) );
  AOI21_X1 U9408 ( .B1(n8187), .B2(n8235), .A(n7601), .ZN(n7605) );
  INV_X1 U9409 ( .A(n7602), .ZN(n7603) );
  NAND2_X1 U9410 ( .A1(n8199), .A2(n7603), .ZN(n7604) );
  OAI211_X1 U9411 ( .C1(n7606), .C2(n8190), .A(n7605), .B(n7604), .ZN(n7607)
         );
  AOI21_X1 U9412 ( .B1(n7608), .B2(n8192), .A(n7607), .ZN(n7609) );
  OAI21_X1 U9413 ( .B1(n7610), .B2(n8206), .A(n7609), .ZN(P2_U3157) );
  INV_X1 U9414 ( .A(n7611), .ZN(n7615) );
  OR2_X1 U9415 ( .A1(n7612), .A2(P1_U3086), .ZN(n9070) );
  NAND2_X1 U9416 ( .A1(n9563), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7613) );
  OAI211_X1 U9417 ( .C1(n7615), .C2(n9572), .A(n9070), .B(n7613), .ZN(P1_U3332) );
  NAND2_X1 U9418 ( .A1(n8673), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7614) );
  OAI211_X1 U9419 ( .C1(n7615), .C2(n6582), .A(n7994), .B(n7614), .ZN(P2_U3272) );
  AOI211_X1 U9420 ( .C1(n7618), .C2(n9768), .A(n7617), .B(n7616), .ZN(n7622)
         );
  AOI22_X1 U9421 ( .A1(n7620), .A2(n6562), .B1(n9786), .B2(
        P1_REG0_REG_12__SCAN_IN), .ZN(n7619) );
  OAI21_X1 U9422 ( .B1(n7622), .B2(n9786), .A(n7619), .ZN(P1_U3489) );
  AOI22_X1 U9423 ( .A1(n7620), .A2(n6572), .B1(n9795), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7621) );
  OAI21_X1 U9424 ( .B1(n7622), .B2(n9795), .A(n7621), .ZN(P1_U3534) );
  NAND2_X1 U9425 ( .A1(n7624), .A2(n7623), .ZN(n7970) );
  XNOR2_X1 U9426 ( .A(n7625), .B(n7970), .ZN(n7626) );
  OAI222_X1 U9427 ( .A1(n10032), .A2(n8211), .B1(n10031), .B2(n9598), .C1(
        n7626), .C2(n10041), .ZN(n8597) );
  INV_X1 U9428 ( .A(n8597), .ZN(n7632) );
  XNOR2_X1 U9429 ( .A(n7627), .B(n7970), .ZN(n8598) );
  INV_X1 U9430 ( .A(n8016), .ZN(n8658) );
  NOR2_X1 U9431 ( .A1(n8658), .A2(n8532), .ZN(n7630) );
  OAI22_X1 U9432 ( .A1(n10035), .A2(n7628), .B1(n8213), .B2(n10022), .ZN(n7629) );
  AOI211_X1 U9433 ( .C1(n8598), .C2(n8536), .A(n7630), .B(n7629), .ZN(n7631)
         );
  OAI21_X1 U9434 ( .B1(n7632), .B2(n10038), .A(n7631), .ZN(P2_U3218) );
  INV_X1 U9435 ( .A(n7633), .ZN(n7652) );
  OAI222_X1 U9436 ( .A1(n9572), .A2(n7652), .B1(P1_U3086), .B2(n7635), .C1(
        n7634), .C2(n9569), .ZN(P1_U3331) );
  OR2_X1 U9437 ( .A1(n7636), .A2(n8236), .ZN(n7637) );
  XNOR2_X1 U9438 ( .A(n7639), .B(n8052), .ZN(n8008) );
  XNOR2_X1 U9439 ( .A(n8008), .B(n8118), .ZN(n7641) );
  AOI21_X1 U9440 ( .B1(n7640), .B2(n7641), .A(n8206), .ZN(n7642) );
  NAND2_X1 U9441 ( .A1(n7642), .A2(n8010), .ZN(n7650) );
  INV_X1 U9442 ( .A(n7643), .ZN(n7648) );
  NAND2_X1 U9443 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n9916) );
  INV_X1 U9444 ( .A(n9916), .ZN(n7644) );
  AOI21_X1 U9445 ( .B1(n8187), .B2(n8234), .A(n7644), .ZN(n7645) );
  OAI21_X1 U9446 ( .B1(n7646), .B2(n8190), .A(n7645), .ZN(n7647) );
  AOI21_X1 U9447 ( .B1(n7648), .B2(n8199), .A(n7647), .ZN(n7649) );
  OAI211_X1 U9448 ( .C1(n10078), .C2(n8220), .A(n7650), .B(n7649), .ZN(
        P2_U3176) );
  OAI222_X1 U9449 ( .A1(n7653), .A2(P2_U3151), .B1(n6582), .B2(n7652), .C1(
        n7651), .C2(n8668), .ZN(P2_U3271) );
  XNOR2_X1 U9450 ( .A(n7654), .B(n8941), .ZN(n7684) );
  INV_X1 U9451 ( .A(n7684), .ZN(n7665) );
  OAI21_X1 U9452 ( .B1(n7656), .B2(n9752), .A(n7655), .ZN(n7680) );
  INV_X1 U9453 ( .A(n7657), .ZN(n7659) );
  INV_X1 U9454 ( .A(n7658), .ZN(n7740) );
  AOI211_X1 U9455 ( .C1(n8845), .C2(n7659), .A(n9422), .B(n7740), .ZN(n7681)
         );
  NAND2_X1 U9456 ( .A1(n7681), .A2(n9731), .ZN(n7662) );
  AOI22_X1 U9457 ( .A1(n9744), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7660), .B2(
        n9733), .ZN(n7661) );
  OAI211_X1 U9458 ( .C1(n8849), .C2(n9737), .A(n7662), .B(n7661), .ZN(n7663)
         );
  AOI21_X1 U9459 ( .B1(n9409), .B2(n7680), .A(n7663), .ZN(n7664) );
  OAI21_X1 U9460 ( .B1(n7665), .B2(n9430), .A(n7664), .ZN(P1_U3280) );
  INV_X1 U9461 ( .A(n7666), .ZN(n7689) );
  OAI222_X1 U9462 ( .A1(n9572), .A2(n7689), .B1(P1_U3086), .B2(n5711), .C1(
        n7667), .C2(n9569), .ZN(P1_U3330) );
  NAND2_X1 U9463 ( .A1(n7669), .A2(n7668), .ZN(n7670) );
  XOR2_X1 U9464 ( .A(n7671), .B(n7670), .Z(n7676) );
  AOI22_X1 U9465 ( .A1(n9086), .A2(n8777), .B1(n9088), .B2(n9066), .ZN(n7736)
         );
  OAI22_X1 U9466 ( .A1(n8780), .A2(n7736), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7672), .ZN(n7674) );
  NOR2_X1 U9467 ( .A1(n9506), .A2(n8785), .ZN(n7673) );
  AOI211_X1 U9468 ( .C1(n8782), .C2(n7741), .A(n7674), .B(n7673), .ZN(n7675)
         );
  OAI21_X1 U9469 ( .B1(n7676), .B2(n8769), .A(n7675), .ZN(P1_U3215) );
  INV_X1 U9470 ( .A(n7677), .ZN(n7691) );
  OAI222_X1 U9471 ( .A1(n9572), .A2(n7691), .B1(P1_U3086), .B2(n7679), .C1(
        n7678), .C2(n9569), .ZN(P1_U3329) );
  NOR2_X1 U9472 ( .A1(n7681), .A2(n7680), .ZN(n7687) );
  NAND2_X1 U9473 ( .A1(n7684), .A2(n7714), .ZN(n7683) );
  AOI22_X1 U9474 ( .A1(n8845), .A2(n6562), .B1(P1_REG0_REG_13__SCAN_IN), .B2(
        n9786), .ZN(n7682) );
  OAI211_X1 U9475 ( .C1(n7687), .C2(n9786), .A(n7683), .B(n7682), .ZN(P1_U3492) );
  NAND2_X1 U9476 ( .A1(n7684), .A2(n7727), .ZN(n7686) );
  AOI22_X1 U9477 ( .A1(n8845), .A2(n6572), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n9795), .ZN(n7685) );
  OAI211_X1 U9478 ( .C1(n7687), .C2(n9795), .A(n7686), .B(n7685), .ZN(P1_U3535) );
  OAI222_X1 U9479 ( .A1(n7690), .A2(P2_U3151), .B1(n6582), .B2(n7689), .C1(
        n7688), .C2(n8668), .ZN(P2_U3270) );
  OAI222_X1 U9480 ( .A1(n7692), .A2(P2_U3151), .B1(n6582), .B2(n7691), .C1(
        n10246), .C2(n8668), .ZN(P2_U3269) );
  AOI21_X1 U9481 ( .B1(n7694), .B2(n7697), .A(n7695), .ZN(n7696) );
  AOI21_X1 U9482 ( .B1(n4624), .B2(n7697), .A(n7696), .ZN(n7702) );
  OAI22_X1 U9483 ( .A1(n7698), .A2(n7750), .B1(n8821), .B2(n7748), .ZN(n7705)
         );
  AOI22_X1 U9484 ( .A1(n8763), .A2(n7705), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n7699) );
  OAI21_X1 U9485 ( .B1(n7707), .B2(n8765), .A(n7699), .ZN(n7700) );
  AOI21_X1 U9486 ( .B1(n8860), .B2(n8767), .A(n7700), .ZN(n7701) );
  OAI21_X1 U9487 ( .B1(n7702), .B2(n8769), .A(n7701), .ZN(P1_U3241) );
  XNOR2_X1 U9488 ( .A(n7703), .B(n8945), .ZN(n7731) );
  NAND2_X1 U9489 ( .A1(n7733), .A2(n8817), .ZN(n7704) );
  XNOR2_X1 U9490 ( .A(n7704), .B(n8945), .ZN(n7706) );
  AOI21_X1 U9491 ( .B1(n7706), .B2(n9710), .A(n7705), .ZN(n7716) );
  OAI21_X1 U9492 ( .B1(n7707), .B2(n9405), .A(n7716), .ZN(n7712) );
  INV_X1 U9493 ( .A(n7739), .ZN(n7709) );
  OAI211_X1 U9494 ( .C1(n7718), .C2(n7709), .A(n9724), .B(n7708), .ZN(n7715)
         );
  AOI22_X1 U9495 ( .A1(n8860), .A2(n9722), .B1(n9721), .B2(
        P1_REG2_REG_15__SCAN_IN), .ZN(n7710) );
  OAI21_X1 U9496 ( .B1(n7715), .B2(n9370), .A(n7710), .ZN(n7711) );
  AOI21_X1 U9497 ( .B1(n7712), .B2(n9409), .A(n7711), .ZN(n7713) );
  OAI21_X1 U9498 ( .B1(n7731), .B2(n9430), .A(n7713), .ZN(P1_U3278) );
  NAND2_X1 U9499 ( .A1(n7716), .A2(n7715), .ZN(n7728) );
  OAI22_X1 U9500 ( .A1(n7718), .A2(n9543), .B1(n9788), .B2(n7717), .ZN(n7719)
         );
  AOI21_X1 U9501 ( .B1(n7728), .B2(n9788), .A(n7719), .ZN(n7720) );
  OAI21_X1 U9502 ( .B1(n7731), .B2(n9555), .A(n7720), .ZN(P1_U3498) );
  INV_X1 U9503 ( .A(n7721), .ZN(n7726) );
  NOR2_X1 U9504 ( .A1(n7722), .A2(P1_U3086), .ZN(n9065) );
  AOI21_X1 U9505 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(n9563), .A(n9065), .ZN(
        n7723) );
  OAI21_X1 U9506 ( .B1(n7726), .B2(n9572), .A(n7723), .ZN(P1_U3328) );
  AOI21_X1 U9507 ( .B1(n8673), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7724), .ZN(
        n7725) );
  OAI21_X1 U9508 ( .B1(n7726), .B2(n6582), .A(n7725), .ZN(P2_U3268) );
  AOI22_X1 U9509 ( .A1(n8860), .A2(n6572), .B1(P1_REG1_REG_15__SCAN_IN), .B2(
        n9795), .ZN(n7730) );
  NAND2_X1 U9510 ( .A1(n7728), .A2(n9797), .ZN(n7729) );
  OAI211_X1 U9511 ( .C1(n7731), .C2(n9484), .A(n7730), .B(n7729), .ZN(P1_U3537) );
  XNOR2_X1 U9512 ( .A(n7732), .B(n8943), .ZN(n7738) );
  OAI211_X1 U9513 ( .C1(n8943), .C2(n7734), .A(n7733), .B(n9710), .ZN(n7735)
         );
  OAI211_X1 U9514 ( .C1(n7738), .C2(n7737), .A(n7736), .B(n7735), .ZN(n9507)
         );
  INV_X1 U9515 ( .A(n9507), .ZN(n7746) );
  INV_X1 U9516 ( .A(n7738), .ZN(n9509) );
  OAI211_X1 U9517 ( .C1(n9506), .C2(n7740), .A(n7739), .B(n9724), .ZN(n9505)
         );
  AOI22_X1 U9518 ( .A1(n9744), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7741), .B2(
        n9733), .ZN(n7743) );
  NAND2_X1 U9519 ( .A1(n8824), .A2(n9722), .ZN(n7742) );
  OAI211_X1 U9520 ( .C1(n9505), .C2(n9370), .A(n7743), .B(n7742), .ZN(n7744)
         );
  AOI21_X1 U9521 ( .B1(n9509), .B2(n9728), .A(n7744), .ZN(n7745) );
  OAI21_X1 U9522 ( .B1(n7746), .B2(n9721), .A(n7745), .ZN(P1_U3279) );
  XNOR2_X1 U9523 ( .A(n7747), .B(n8947), .ZN(n7752) );
  OAI22_X1 U9524 ( .A1(n7751), .A2(n7750), .B1(n7749), .B2(n7748), .ZN(n8712)
         );
  AOI21_X1 U9525 ( .B1(n7752), .B2(n9710), .A(n8712), .ZN(n9503) );
  NAND2_X1 U9526 ( .A1(n7753), .A2(n8947), .ZN(n9497) );
  NAND3_X1 U9527 ( .A1(n9498), .A2(n9497), .A3(n9741), .ZN(n7759) );
  INV_X1 U9528 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7754) );
  OAI22_X1 U9529 ( .A1(n9409), .A2(n7754), .B1(n8710), .B2(n9405), .ZN(n7757)
         );
  OAI211_X1 U9530 ( .C1(n8715), .C2(n7755), .A(n9724), .B(n9423), .ZN(n9502)
         );
  NOR2_X1 U9531 ( .A1(n9502), .A2(n9370), .ZN(n7756) );
  AOI211_X1 U9532 ( .C1(n9722), .C2(n9500), .A(n7757), .B(n7756), .ZN(n7758)
         );
  OAI211_X1 U9533 ( .C1(n9744), .C2(n9503), .A(n7759), .B(n7758), .ZN(P1_U3277) );
  NAND2_X1 U9534 ( .A1(n7760), .A2(n9741), .ZN(n7770) );
  INV_X1 U9535 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n7761) );
  OAI22_X1 U9536 ( .A1(n7762), .A2(n9737), .B1(n7761), .B2(n9409), .ZN(n7767)
         );
  AOI21_X1 U9537 ( .B1(n7764), .B2(n9733), .A(n7763), .ZN(n7765) );
  NOR2_X1 U9538 ( .A1(n7765), .A2(n9721), .ZN(n7766) );
  AOI211_X1 U9539 ( .C1(n9731), .C2(n7768), .A(n7767), .B(n7766), .ZN(n7769)
         );
  NAND2_X1 U9540 ( .A1(n7770), .A2(n7769), .ZN(P1_U3356) );
  INV_X1 U9541 ( .A(n7771), .ZN(n8776) );
  INV_X1 U9542 ( .A(n7772), .ZN(n7773) );
  NAND2_X1 U9543 ( .A1(n8776), .A2(n7773), .ZN(n7776) );
  INV_X1 U9544 ( .A(n9272), .ZN(n7780) );
  NAND2_X1 U9545 ( .A1(n9073), .A2(n8777), .ZN(n7778) );
  NAND2_X1 U9546 ( .A1(n9075), .A2(n9066), .ZN(n7777) );
  NAND2_X1 U9547 ( .A1(n7778), .A2(n7777), .ZN(n9278) );
  AOI22_X1 U9548 ( .A1(n8763), .A2(n9278), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n7779) );
  OAI21_X1 U9549 ( .B1(n7780), .B2(n8765), .A(n7779), .ZN(n7781) );
  AOI21_X1 U9550 ( .B1(n9269), .B2(n8767), .A(n7781), .ZN(n7782) );
  OAI21_X1 U9551 ( .B1(n7783), .B2(n8769), .A(n7782), .ZN(P1_U3214) );
  INV_X1 U9552 ( .A(n7784), .ZN(n7794) );
  INV_X1 U9553 ( .A(n7976), .ZN(n7942) );
  INV_X1 U9554 ( .A(n7785), .ZN(n7786) );
  MUX2_X1 U9555 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n4610), .Z(n7795) );
  XNOR2_X1 U9556 ( .A(n7795), .B(SI_30_), .ZN(n7796) );
  NAND2_X1 U9557 ( .A1(n8905), .A2(n7804), .ZN(n7792) );
  INV_X1 U9558 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8069) );
  OR2_X1 U9559 ( .A1(n7790), .A2(n8069), .ZN(n7791) );
  INV_X1 U9560 ( .A(n8221), .ZN(n7805) );
  NAND2_X1 U9561 ( .A1(n8610), .A2(n7805), .ZN(n7977) );
  AOI21_X1 U9562 ( .B1(n7794), .B2(n7942), .A(n4557), .ZN(n7808) );
  OAI22_X1 U9563 ( .A1(n7797), .A2(n7796), .B1(SI_30_), .B2(n7795), .ZN(n7802)
         );
  INV_X1 U9564 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n7799) );
  MUX2_X1 U9565 ( .A(n7228), .B(n7799), .S(n4610), .Z(n7800) );
  XNOR2_X1 U9566 ( .A(n7800), .B(SI_31_), .ZN(n7801) );
  OAI21_X1 U9567 ( .B1(n8610), .B2(n8360), .A(n8363), .ZN(n7807) );
  INV_X1 U9568 ( .A(n7978), .ZN(n7806) );
  AOI22_X1 U9569 ( .A1(n7808), .A2(n7807), .B1(n7806), .B2(n8605), .ZN(n7987)
         );
  MUX2_X1 U9570 ( .A(n8222), .B(n8066), .S(n7947), .Z(n7944) );
  INV_X1 U9571 ( .A(n8385), .ZN(n7811) );
  INV_X1 U9572 ( .A(n7809), .ZN(n7813) );
  MUX2_X1 U9573 ( .A(n7812), .B(n7813), .S(n7946), .Z(n7810) );
  NOR2_X1 U9574 ( .A1(n7811), .A2(n7810), .ZN(n7941) );
  INV_X1 U9575 ( .A(n8392), .ZN(n8397) );
  NAND2_X1 U9576 ( .A1(n7907), .A2(n8498), .ZN(n7814) );
  NAND2_X1 U9577 ( .A1(n7814), .A2(n7946), .ZN(n7905) );
  MUX2_X1 U9578 ( .A(n7816), .B(n7815), .S(n7947), .Z(n7903) );
  MUX2_X1 U9579 ( .A(n7820), .B(n7817), .S(n7947), .Z(n7827) );
  NAND2_X1 U9580 ( .A1(n7818), .A2(n7991), .ZN(n7822) );
  NAND2_X1 U9581 ( .A1(n7818), .A2(n7825), .ZN(n7819) );
  NAND3_X1 U9582 ( .A1(n7820), .A2(n7819), .A3(n7947), .ZN(n7821) );
  OAI21_X1 U9583 ( .B1(n7954), .B2(n7822), .A(n7821), .ZN(n7823) );
  OAI21_X1 U9584 ( .B1(n7825), .B2(n7824), .A(n7823), .ZN(n7826) );
  NAND3_X1 U9585 ( .A1(n7827), .A2(n10025), .A3(n7826), .ZN(n7834) );
  NAND2_X1 U9586 ( .A1(n7849), .A2(n7828), .ZN(n7831) );
  NAND2_X1 U9587 ( .A1(n7835), .A2(n7829), .ZN(n7830) );
  MUX2_X1 U9588 ( .A(n7831), .B(n7830), .S(n7946), .Z(n7832) );
  INV_X1 U9589 ( .A(n7832), .ZN(n7833) );
  NAND2_X1 U9590 ( .A1(n7834), .A2(n7833), .ZN(n7850) );
  NAND3_X1 U9591 ( .A1(n7850), .A2(n7957), .A3(n7835), .ZN(n7837) );
  NAND3_X1 U9592 ( .A1(n7837), .A2(n7836), .A3(n7855), .ZN(n7838) );
  NAND3_X1 U9593 ( .A1(n7838), .A2(n7857), .A3(n7851), .ZN(n7842) );
  AND2_X1 U9594 ( .A1(n7839), .A2(n7946), .ZN(n7840) );
  NAND2_X1 U9595 ( .A1(n7846), .A2(n7840), .ZN(n7861) );
  NAND3_X1 U9596 ( .A1(n7867), .A2(n7947), .A3(n7863), .ZN(n7841) );
  NAND2_X1 U9597 ( .A1(n7861), .A2(n7841), .ZN(n7858) );
  NAND4_X1 U9598 ( .A1(n7842), .A2(n7859), .A3(n7858), .A4(n7854), .ZN(n7847)
         );
  INV_X1 U9599 ( .A(n7843), .ZN(n7844) );
  NAND2_X1 U9600 ( .A1(n7858), .A2(n7844), .ZN(n7845) );
  NAND4_X1 U9601 ( .A1(n7847), .A2(n7846), .A3(n7845), .A4(n7870), .ZN(n7848)
         );
  NAND2_X1 U9602 ( .A1(n7848), .A2(n7868), .ZN(n7873) );
  NAND3_X1 U9603 ( .A1(n7850), .A2(n7957), .A3(n7849), .ZN(n7853) );
  NAND3_X1 U9604 ( .A1(n7853), .A2(n7852), .A3(n7851), .ZN(n7856) );
  NAND3_X1 U9605 ( .A1(n7856), .A2(n7855), .A3(n7854), .ZN(n7860) );
  NAND4_X1 U9606 ( .A1(n7860), .A2(n7859), .A3(n7858), .A4(n7857), .ZN(n7869)
         );
  INV_X1 U9607 ( .A(n7861), .ZN(n7865) );
  NAND2_X1 U9608 ( .A1(n7863), .A2(n7862), .ZN(n7864) );
  NAND2_X1 U9609 ( .A1(n7865), .A2(n7864), .ZN(n7866) );
  NAND4_X1 U9610 ( .A1(n7869), .A2(n7868), .A3(n7867), .A4(n7866), .ZN(n7871)
         );
  NAND2_X1 U9611 ( .A1(n7871), .A2(n7870), .ZN(n7872) );
  MUX2_X1 U9612 ( .A(n7873), .B(n7872), .S(n7946), .Z(n7876) );
  INV_X1 U9613 ( .A(n7964), .ZN(n7874) );
  NOR2_X1 U9614 ( .A1(n7968), .A2(n7874), .ZN(n7875) );
  NAND2_X1 U9615 ( .A1(n7876), .A2(n7875), .ZN(n7889) );
  NAND2_X1 U9616 ( .A1(n7881), .A2(n7877), .ZN(n7878) );
  NAND2_X1 U9617 ( .A1(n7878), .A2(n7880), .ZN(n7884) );
  NAND2_X1 U9618 ( .A1(n7880), .A2(n7879), .ZN(n7882) );
  NAND2_X1 U9619 ( .A1(n7882), .A2(n7881), .ZN(n7883) );
  MUX2_X1 U9620 ( .A(n7884), .B(n7883), .S(n7946), .Z(n7888) );
  INV_X1 U9621 ( .A(n7885), .ZN(n7886) );
  OR2_X1 U9622 ( .A1(n7887), .A2(n7886), .ZN(n9595) );
  INV_X1 U9623 ( .A(n9595), .ZN(n9589) );
  INV_X1 U9624 ( .A(n7890), .ZN(n7891) );
  MUX2_X1 U9625 ( .A(n7892), .B(n7891), .S(n7947), .Z(n7894) );
  MUX2_X1 U9626 ( .A(n7896), .B(n7895), .S(n7946), .Z(n7897) );
  INV_X1 U9627 ( .A(n7898), .ZN(n7899) );
  MUX2_X1 U9628 ( .A(n7900), .B(n7899), .S(n7946), .Z(n7901) );
  NAND3_X1 U9629 ( .A1(n8521), .A2(n7903), .A3(n7902), .ZN(n7904) );
  NAND2_X1 U9630 ( .A1(n7905), .A2(n7904), .ZN(n7911) );
  NAND2_X1 U9631 ( .A1(n7910), .A2(n7906), .ZN(n7908) );
  AND3_X1 U9632 ( .A1(n7953), .A2(n7911), .A3(n7910), .ZN(n7912) );
  NAND2_X1 U9633 ( .A1(n7913), .A2(n7918), .ZN(n7914) );
  NAND2_X1 U9634 ( .A1(n7914), .A2(n7917), .ZN(n7922) );
  NAND2_X1 U9635 ( .A1(n7920), .A2(n7919), .ZN(n7921) );
  MUX2_X1 U9636 ( .A(n7922), .B(n7921), .S(n7946), .Z(n7923) );
  MUX2_X1 U9637 ( .A(n7925), .B(n7924), .S(n7946), .Z(n7926) );
  INV_X1 U9638 ( .A(n7950), .ZN(n7927) );
  AOI21_X1 U9639 ( .B1(n7951), .B2(n7952), .A(n7927), .ZN(n7931) );
  OAI21_X1 U9640 ( .B1(n7928), .B2(n7952), .A(n7951), .ZN(n7929) );
  NAND2_X1 U9641 ( .A1(n7929), .A2(n7946), .ZN(n7930) );
  MUX2_X1 U9642 ( .A(n7933), .B(n7932), .S(n7947), .Z(n7934) );
  NAND3_X1 U9643 ( .A1(n8397), .A2(n7935), .A3(n7934), .ZN(n7940) );
  INV_X1 U9644 ( .A(n7936), .ZN(n7938) );
  MUX2_X1 U9645 ( .A(n7938), .B(n7937), .S(n7947), .Z(n7939) );
  NAND2_X1 U9646 ( .A1(n8363), .A2(n8360), .ZN(n7980) );
  AND3_X1 U9647 ( .A1(n7980), .A2(n7948), .A3(n7977), .ZN(n7949) );
  NAND2_X1 U9648 ( .A1(n7952), .A2(n8423), .ZN(n8437) );
  NOR4_X1 U9649 ( .A1(n7956), .A2(n7955), .A3(n10039), .A4(n7954), .ZN(n7958)
         );
  NAND3_X1 U9650 ( .A1(n7958), .A2(n7957), .A3(n4528), .ZN(n7962) );
  NOR4_X1 U9651 ( .A1(n7962), .A2(n7961), .A3(n7960), .A4(n7959), .ZN(n7966)
         );
  NAND4_X1 U9652 ( .A1(n7966), .A2(n7965), .A3(n7964), .A4(n7963), .ZN(n7967)
         );
  NOR4_X1 U9653 ( .A1(n9589), .A2(n7969), .A3(n7968), .A4(n7967), .ZN(n7971)
         );
  NAND4_X1 U9654 ( .A1(n8521), .A2(n8529), .A3(n7971), .A4(n7970), .ZN(n7972)
         );
  OR4_X1 U9655 ( .A1(n8474), .A2(n6159), .A3(n8502), .A4(n7972), .ZN(n7973) );
  NOR4_X1 U9656 ( .A1(n8437), .A2(n8449), .A3(n8454), .A4(n7973), .ZN(n7974)
         );
  NAND4_X1 U9657 ( .A1(n8385), .A2(n8410), .A3(n8426), .A4(n7974), .ZN(n7975)
         );
  NOR4_X1 U9658 ( .A1(n7976), .A2(n8060), .A3(n8392), .A4(n7975), .ZN(n7979)
         );
  NAND4_X1 U9659 ( .A1(n7980), .A2(n7979), .A3(n7978), .A4(n7977), .ZN(n7983)
         );
  INV_X1 U9660 ( .A(n8360), .ZN(n7981) );
  AOI22_X1 U9661 ( .A1(n7983), .A2(n7982), .B1(n7981), .B2(n8605), .ZN(n7984)
         );
  OAI211_X1 U9662 ( .C1(n7987), .C2(n7986), .A(n7985), .B(n7984), .ZN(n7988)
         );
  XNOR2_X1 U9663 ( .A(n7988), .B(n8353), .ZN(n7995) );
  NOR3_X1 U9664 ( .A1(n7990), .A2(n8346), .A3(n7989), .ZN(n7993) );
  OAI21_X1 U9665 ( .B1(n7994), .B2(n7991), .A(P2_B_REG_SCAN_IN), .ZN(n7992) );
  OAI22_X1 U9666 ( .A1(n7995), .A2(n7994), .B1(n7993), .B2(n7992), .ZN(
        P2_U3296) );
  INV_X1 U9667 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7997) );
  INV_X1 U9668 ( .A(n8905), .ZN(n8070) );
  OAI222_X1 U9669 ( .A1(n9569), .A2(n7997), .B1(n9572), .B2(n8070), .C1(
        P1_U3086), .C2(n7996), .ZN(P1_U3325) );
  INV_X1 U9670 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8005) );
  XOR2_X1 U9671 ( .A(n8060), .B(n7998), .Z(n8379) );
  OAI222_X1 U9672 ( .A1(n9569), .A2(n8007), .B1(n9572), .B2(n8006), .C1(n4507), 
        .C2(P1_U3086), .ZN(P1_U3336) );
  XNOR2_X1 U9673 ( .A(n10089), .B(n8052), .ZN(n8011) );
  XNOR2_X1 U9674 ( .A(n8011), .B(n8234), .ZN(n8116) );
  INV_X1 U9675 ( .A(n8011), .ZN(n8012) );
  XNOR2_X1 U9676 ( .A(n9591), .B(n8056), .ZN(n8168) );
  NOR2_X1 U9677 ( .A1(n8168), .A2(n8233), .ZN(n8013) );
  XNOR2_X1 U9678 ( .A(n8086), .B(n6895), .ZN(n8014) );
  XNOR2_X1 U9679 ( .A(n8014), .B(n9598), .ZN(n8079) );
  INV_X1 U9680 ( .A(n8014), .ZN(n8015) );
  XNOR2_X1 U9681 ( .A(n8016), .B(n6895), .ZN(n8017) );
  XNOR2_X1 U9682 ( .A(n8017), .B(n8527), .ZN(n8207) );
  INV_X1 U9683 ( .A(n8017), .ZN(n8018) );
  NAND2_X1 U9684 ( .A1(n8018), .A2(n8231), .ZN(n8019) );
  NAND2_X1 U9685 ( .A1(n8209), .A2(n8019), .ZN(n8095) );
  XNOR2_X1 U9686 ( .A(n8531), .B(n6895), .ZN(n8033) );
  XNOR2_X1 U9687 ( .A(n8033), .B(n8211), .ZN(n8134) );
  XNOR2_X1 U9688 ( .A(n8489), .B(n6895), .ZN(n8020) );
  NAND2_X1 U9689 ( .A1(n8020), .A2(n8497), .ZN(n8035) );
  INV_X1 U9690 ( .A(n8035), .ZN(n8032) );
  XNOR2_X1 U9691 ( .A(n8020), .B(n8229), .ZN(n8100) );
  INV_X1 U9692 ( .A(n8100), .ZN(n8026) );
  XNOR2_X1 U9693 ( .A(n8503), .B(n8052), .ZN(n8021) );
  NAND2_X1 U9694 ( .A1(n8021), .A2(n8103), .ZN(n8023) );
  INV_X1 U9695 ( .A(n8023), .ZN(n8022) );
  XNOR2_X1 U9696 ( .A(n8021), .B(n8512), .ZN(n8186) );
  OR2_X1 U9697 ( .A1(n8022), .A2(n8186), .ZN(n8028) );
  INV_X1 U9698 ( .A(n8028), .ZN(n8025) );
  XNOR2_X1 U9699 ( .A(n8590), .B(n6895), .ZN(n8027) );
  NAND2_X1 U9700 ( .A1(n8027), .A2(n8528), .ZN(n8183) );
  AND2_X1 U9701 ( .A1(n8183), .A2(n8023), .ZN(n8024) );
  OR2_X1 U9702 ( .A1(n8025), .A2(n8024), .ZN(n8097) );
  OR2_X1 U9703 ( .A1(n8026), .A2(n8097), .ZN(n8034) );
  INV_X1 U9704 ( .A(n8034), .ZN(n8030) );
  XNOR2_X1 U9705 ( .A(n8027), .B(n8230), .ZN(n8143) );
  AND2_X1 U9706 ( .A1(n8143), .A2(n8028), .ZN(n8096) );
  AND2_X1 U9707 ( .A1(n8096), .A2(n8100), .ZN(n8029) );
  OR2_X1 U9708 ( .A1(n8030), .A2(n8029), .ZN(n8031) );
  NOR2_X1 U9709 ( .A1(n8032), .A2(n8031), .ZN(n8038) );
  OR2_X1 U9710 ( .A1(n8134), .A2(n8038), .ZN(n8158) );
  XNOR2_X1 U9711 ( .A(n8470), .B(n6895), .ZN(n8040) );
  XNOR2_X1 U9712 ( .A(n8040), .B(n8485), .ZN(n8162) );
  INV_X1 U9713 ( .A(n8162), .ZN(n8039) );
  NAND2_X1 U9714 ( .A1(n8033), .A2(n8211), .ZN(n8144) );
  AND2_X1 U9715 ( .A1(n8144), .A2(n8034), .ZN(n8036) );
  AND2_X1 U9716 ( .A1(n8036), .A2(n8035), .ZN(n8037) );
  OR2_X1 U9717 ( .A1(n8038), .A2(n8037), .ZN(n8159) );
  NAND2_X1 U9718 ( .A1(n8040), .A2(n8456), .ZN(n8107) );
  XNOR2_X1 U9719 ( .A(n8464), .B(n6895), .ZN(n8042) );
  NAND2_X1 U9720 ( .A1(n8042), .A2(n8478), .ZN(n8041) );
  INV_X1 U9721 ( .A(n8041), .ZN(n8043) );
  XNOR2_X1 U9722 ( .A(n8042), .B(n8228), .ZN(n8110) );
  XOR2_X1 U9723 ( .A(n8052), .B(n8568), .Z(n8045) );
  INV_X1 U9724 ( .A(n8045), .ZN(n8044) );
  XNOR2_X1 U9725 ( .A(n8044), .B(n8227), .ZN(n8177) );
  XNOR2_X1 U9726 ( .A(n8438), .B(n8052), .ZN(n8047) );
  XNOR2_X1 U9727 ( .A(n8046), .B(n8047), .ZN(n8089) );
  INV_X1 U9728 ( .A(n8046), .ZN(n8048) );
  NAND2_X1 U9729 ( .A1(n8048), .A2(n8047), .ZN(n8049) );
  XNOR2_X1 U9730 ( .A(n8421), .B(n6895), .ZN(n8050) );
  XNOR2_X1 U9731 ( .A(n8050), .B(n8225), .ZN(n8152) );
  NAND2_X1 U9732 ( .A1(n8050), .A2(n8436), .ZN(n8051) );
  XNOR2_X1 U9733 ( .A(n8407), .B(n6895), .ZN(n8053) );
  XNOR2_X1 U9734 ( .A(n8053), .B(n8415), .ZN(n8127) );
  NAND2_X1 U9735 ( .A1(n8126), .A2(n8127), .ZN(n8055) );
  NAND2_X1 U9736 ( .A1(n8053), .A2(n8395), .ZN(n8054) );
  XNOR2_X1 U9737 ( .A(n8203), .B(n8056), .ZN(n8057) );
  NAND2_X1 U9738 ( .A1(n8057), .A2(n8224), .ZN(n8195) );
  INV_X1 U9739 ( .A(n8057), .ZN(n8058) );
  NAND2_X1 U9740 ( .A1(n8058), .A2(n8406), .ZN(n8196) );
  XNOR2_X1 U9741 ( .A(n8386), .B(n6895), .ZN(n8059) );
  XNOR2_X1 U9742 ( .A(n8059), .B(n8396), .ZN(n8071) );
  XOR2_X1 U9743 ( .A(n6895), .B(n8060), .Z(n8061) );
  NOR2_X1 U9744 ( .A1(n8062), .A2(n8212), .ZN(n8065) );
  AOI22_X1 U9745 ( .A1(n8376), .A2(n8199), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8063) );
  OAI21_X1 U9746 ( .B1(n8396), .B2(n8190), .A(n8063), .ZN(n8064) );
  AOI211_X1 U9747 ( .C1(n8066), .C2(n8192), .A(n8065), .B(n8064), .ZN(n8067)
         );
  OAI21_X1 U9748 ( .B1(n8068), .B2(n8206), .A(n8067), .ZN(P2_U3160) );
  OAI222_X1 U9749 ( .A1(n5741), .A2(P2_U3151), .B1(n6582), .B2(n8070), .C1(
        n8069), .C2(n8668), .ZN(P2_U3265) );
  XNOR2_X1 U9750 ( .A(n8072), .B(n8071), .ZN(n8077) );
  NOR2_X1 U9751 ( .A1(n8383), .A2(n8212), .ZN(n8075) );
  AOI22_X1 U9752 ( .A1(n8387), .A2(n8199), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8073) );
  OAI21_X1 U9753 ( .B1(n8406), .B2(n8190), .A(n8073), .ZN(n8074) );
  AOI211_X1 U9754 ( .C1(n8386), .C2(n8192), .A(n8075), .B(n8074), .ZN(n8076)
         );
  OAI21_X1 U9755 ( .B1(n8077), .B2(n8206), .A(n8076), .ZN(P2_U3154) );
  XOR2_X1 U9756 ( .A(n8079), .B(n8078), .Z(n8088) );
  INV_X1 U9757 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8080) );
  OAI22_X1 U9758 ( .A1(n8190), .A2(n8081), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8080), .ZN(n8082) );
  AOI21_X1 U9759 ( .B1(n8187), .B2(n8231), .A(n8082), .ZN(n8083) );
  OAI21_X1 U9760 ( .B1(n8084), .B2(n8214), .A(n8083), .ZN(n8085) );
  AOI21_X1 U9761 ( .B1(n8086), .B2(n8192), .A(n8085), .ZN(n8087) );
  OAI21_X1 U9762 ( .B1(n8088), .B2(n8206), .A(n8087), .ZN(P2_U3155) );
  XNOR2_X1 U9763 ( .A(n8089), .B(n8226), .ZN(n8094) );
  INV_X1 U9764 ( .A(n8190), .ZN(n8217) );
  AOI22_X1 U9765 ( .A1(n8227), .A2(n8217), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8091) );
  NAND2_X1 U9766 ( .A1(n8199), .A2(n8439), .ZN(n8090) );
  OAI211_X1 U9767 ( .C1(n8436), .C2(n8212), .A(n8091), .B(n8090), .ZN(n8092)
         );
  AOI21_X1 U9768 ( .B1(n8438), .B2(n8192), .A(n8092), .ZN(n8093) );
  OAI21_X1 U9769 ( .B1(n8094), .B2(n8206), .A(n8093), .ZN(P2_U3156) );
  NAND2_X1 U9770 ( .A1(n8146), .A2(n8144), .ZN(n8142) );
  NAND2_X1 U9771 ( .A1(n8142), .A2(n8096), .ZN(n8098) );
  NAND2_X1 U9772 ( .A1(n8098), .A2(n8097), .ZN(n8099) );
  XOR2_X1 U9773 ( .A(n8100), .B(n8099), .Z(n8106) );
  AOI22_X1 U9774 ( .A1(n8187), .A2(n8485), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3151), .ZN(n8102) );
  NAND2_X1 U9775 ( .A1(n8199), .A2(n8490), .ZN(n8101) );
  OAI211_X1 U9776 ( .C1(n8103), .C2(n8190), .A(n8102), .B(n8101), .ZN(n8104)
         );
  AOI21_X1 U9777 ( .B1(n8489), .B2(n8192), .A(n8104), .ZN(n8105) );
  OAI21_X1 U9778 ( .B1(n8106), .B2(n8206), .A(n8105), .ZN(P2_U3159) );
  NAND2_X1 U9779 ( .A1(n8108), .A2(n8107), .ZN(n8109) );
  XOR2_X1 U9780 ( .A(n8110), .B(n8109), .Z(n8115) );
  AOI22_X1 U9781 ( .A1(n8227), .A2(n8187), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8112) );
  NAND2_X1 U9782 ( .A1(n8199), .A2(n8465), .ZN(n8111) );
  OAI211_X1 U9783 ( .C1(n8456), .C2(n8190), .A(n8112), .B(n8111), .ZN(n8113)
         );
  AOI21_X1 U9784 ( .B1(n8464), .B2(n8192), .A(n8113), .ZN(n8114) );
  OAI21_X1 U9785 ( .B1(n8115), .B2(n8206), .A(n8114), .ZN(P2_U3163) );
  XNOR2_X1 U9786 ( .A(n8117), .B(n8116), .ZN(n8125) );
  NAND2_X1 U9787 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9933) );
  INV_X1 U9788 ( .A(n9933), .ZN(n8120) );
  NOR2_X1 U9789 ( .A1(n8190), .A2(n8118), .ZN(n8119) );
  AOI211_X1 U9790 ( .C1(n8187), .C2(n8233), .A(n8120), .B(n8119), .ZN(n8121)
         );
  OAI21_X1 U9791 ( .B1(n8122), .B2(n8214), .A(n8121), .ZN(n8123) );
  AOI21_X1 U9792 ( .B1(n10089), .B2(n8192), .A(n8123), .ZN(n8124) );
  OAI21_X1 U9793 ( .B1(n8125), .B2(n8206), .A(n8124), .ZN(P2_U3164) );
  XOR2_X1 U9794 ( .A(n8127), .B(n8126), .Z(n8132) );
  AOI22_X1 U9795 ( .A1(n8225), .A2(n8217), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8129) );
  NAND2_X1 U9796 ( .A1(n8408), .A2(n8199), .ZN(n8128) );
  OAI211_X1 U9797 ( .C1(n8406), .C2(n8212), .A(n8129), .B(n8128), .ZN(n8130)
         );
  AOI21_X1 U9798 ( .B1(n8407), .B2(n8192), .A(n8130), .ZN(n8131) );
  OAI21_X1 U9799 ( .B1(n8132), .B2(n8206), .A(n8131), .ZN(P2_U3165) );
  INV_X1 U9800 ( .A(n8146), .ZN(n8133) );
  AOI21_X1 U9801 ( .B1(n8134), .B2(n8095), .A(n8133), .ZN(n8139) );
  AOI22_X1 U9802 ( .A1(n8187), .A2(n8230), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3151), .ZN(n8136) );
  NAND2_X1 U9803 ( .A1(n8217), .A2(n8231), .ZN(n8135) );
  OAI211_X1 U9804 ( .C1(n8214), .C2(n8533), .A(n8136), .B(n8135), .ZN(n8137)
         );
  AOI21_X1 U9805 ( .B1(n8531), .B2(n8192), .A(n8137), .ZN(n8138) );
  OAI21_X1 U9806 ( .B1(n8139), .B2(n8206), .A(n8138), .ZN(P2_U3166) );
  AOI22_X1 U9807 ( .A1(n8187), .A2(n8512), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n8141) );
  NAND2_X1 U9808 ( .A1(n8217), .A2(n8514), .ZN(n8140) );
  OAI211_X1 U9809 ( .C1(n8214), .C2(n8517), .A(n8141), .B(n8140), .ZN(n8149)
         );
  NAND2_X1 U9810 ( .A1(n8142), .A2(n8143), .ZN(n8184) );
  INV_X1 U9811 ( .A(n8143), .ZN(n8145) );
  NAND3_X1 U9812 ( .A1(n8146), .A2(n8145), .A3(n8144), .ZN(n8147) );
  AOI21_X1 U9813 ( .B1(n8184), .B2(n8147), .A(n8206), .ZN(n8148) );
  AOI211_X1 U9814 ( .C1(n8590), .C2(n8192), .A(n8149), .B(n8148), .ZN(n8150)
         );
  INV_X1 U9815 ( .A(n8150), .ZN(P2_U3168) );
  XOR2_X1 U9816 ( .A(n8152), .B(n8151), .Z(n8157) );
  AOI22_X1 U9817 ( .A1(n8226), .A2(n8217), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8154) );
  NAND2_X1 U9818 ( .A1(n8419), .A2(n8199), .ZN(n8153) );
  OAI211_X1 U9819 ( .C1(n8395), .C2(n8212), .A(n8154), .B(n8153), .ZN(n8155)
         );
  AOI21_X1 U9820 ( .B1(n8421), .B2(n8192), .A(n8155), .ZN(n8156) );
  OAI21_X1 U9821 ( .B1(n8157), .B2(n8206), .A(n8156), .ZN(P2_U3169) );
  OR2_X1 U9822 ( .A1(n8095), .A2(n8158), .ZN(n8160) );
  NAND2_X1 U9823 ( .A1(n8160), .A2(n8159), .ZN(n8161) );
  XOR2_X1 U9824 ( .A(n8162), .B(n8161), .Z(n8167) );
  AOI22_X1 U9825 ( .A1(n8228), .A2(n8187), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8164) );
  NAND2_X1 U9826 ( .A1(n8199), .A2(n8471), .ZN(n8163) );
  OAI211_X1 U9827 ( .C1(n8497), .C2(n8190), .A(n8164), .B(n8163), .ZN(n8165)
         );
  AOI21_X1 U9828 ( .B1(n8470), .B2(n8192), .A(n8165), .ZN(n8166) );
  OAI21_X1 U9829 ( .B1(n8167), .B2(n8206), .A(n8166), .ZN(P2_U3173) );
  XNOR2_X1 U9830 ( .A(n8168), .B(n8233), .ZN(n8169) );
  XNOR2_X1 U9831 ( .A(n4586), .B(n8169), .ZN(n8175) );
  NAND2_X1 U9832 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9949) );
  INV_X1 U9833 ( .A(n9949), .ZN(n8171) );
  NOR2_X1 U9834 ( .A1(n8212), .A2(n9598), .ZN(n8170) );
  AOI211_X1 U9835 ( .C1(n8217), .C2(n8234), .A(n8171), .B(n8170), .ZN(n8172)
         );
  OAI21_X1 U9836 ( .B1(n9594), .B2(n8214), .A(n8172), .ZN(n8173) );
  AOI21_X1 U9837 ( .B1(n9591), .B2(n8192), .A(n8173), .ZN(n8174) );
  OAI21_X1 U9838 ( .B1(n8175), .B2(n8206), .A(n8174), .ZN(P2_U3174) );
  XOR2_X1 U9839 ( .A(n8177), .B(n8176), .Z(n8182) );
  AOI22_X1 U9840 ( .A1(n8228), .A2(n8217), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8179) );
  NAND2_X1 U9841 ( .A1(n8199), .A2(n8448), .ZN(n8178) );
  OAI211_X1 U9842 ( .C1(n8447), .C2(n8212), .A(n8179), .B(n8178), .ZN(n8180)
         );
  AOI21_X1 U9843 ( .B1(n8568), .B2(n8192), .A(n8180), .ZN(n8181) );
  OAI21_X1 U9844 ( .B1(n8182), .B2(n8206), .A(n8181), .ZN(P2_U3175) );
  NAND2_X1 U9845 ( .A1(n8184), .A2(n8183), .ZN(n8185) );
  XOR2_X1 U9846 ( .A(n8186), .B(n8185), .Z(n8194) );
  AND2_X1 U9847 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8301) );
  AOI21_X1 U9848 ( .B1(n8187), .B2(n8229), .A(n8301), .ZN(n8189) );
  NAND2_X1 U9849 ( .A1(n8199), .A2(n8504), .ZN(n8188) );
  OAI211_X1 U9850 ( .C1(n8528), .C2(n8190), .A(n8189), .B(n8188), .ZN(n8191)
         );
  AOI21_X1 U9851 ( .B1(n8503), .B2(n8192), .A(n8191), .ZN(n8193) );
  OAI21_X1 U9852 ( .B1(n8194), .B2(n8206), .A(n8193), .ZN(P2_U3178) );
  NAND2_X1 U9853 ( .A1(n8196), .A2(n8195), .ZN(n8197) );
  XNOR2_X1 U9854 ( .A(n8198), .B(n8197), .ZN(n8205) );
  AOI22_X1 U9855 ( .A1(n8415), .A2(n8217), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8201) );
  NAND2_X1 U9856 ( .A1(n8399), .A2(n8199), .ZN(n8200) );
  OAI211_X1 U9857 ( .C1(n8396), .C2(n8212), .A(n8201), .B(n8200), .ZN(n8202)
         );
  AOI21_X1 U9858 ( .B1(n8203), .B2(n8192), .A(n8202), .ZN(n8204) );
  OAI21_X1 U9859 ( .B1(n8205), .B2(n8206), .A(n8204), .ZN(P2_U3180) );
  AOI21_X1 U9860 ( .B1(n8208), .B2(n8207), .A(n8206), .ZN(n8210) );
  NAND2_X1 U9861 ( .A1(n8210), .A2(n8209), .ZN(n8219) );
  NAND2_X1 U9862 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9982) );
  OAI21_X1 U9863 ( .B1(n8212), .B2(n8211), .A(n9982), .ZN(n8216) );
  NOR2_X1 U9864 ( .A1(n8214), .A2(n8213), .ZN(n8215) );
  AOI211_X1 U9865 ( .C1(n8217), .C2(n8232), .A(n8216), .B(n8215), .ZN(n8218)
         );
  OAI211_X1 U9866 ( .C1(n8658), .C2(n8220), .A(n8219), .B(n8218), .ZN(P2_U3181) );
  MUX2_X1 U9867 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8221), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9868 ( .A(n8222), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8297), .Z(
        P2_U3519) );
  MUX2_X1 U9869 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8223), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9870 ( .A(n8224), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8297), .Z(
        P2_U3517) );
  MUX2_X1 U9871 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8415), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9872 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8225), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9873 ( .A(n8226), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8297), .Z(
        P2_U3514) );
  MUX2_X1 U9874 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8227), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9875 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8228), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9876 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8485), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9877 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8229), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9878 ( .A(n8512), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8297), .Z(
        P2_U3509) );
  MUX2_X1 U9879 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8230), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9880 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8514), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9881 ( .A(n8231), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8297), .Z(
        P2_U3506) );
  MUX2_X1 U9882 ( .A(n8232), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8297), .Z(
        P2_U3505) );
  MUX2_X1 U9883 ( .A(n8233), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8297), .Z(
        P2_U3504) );
  MUX2_X1 U9884 ( .A(n8234), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8297), .Z(
        P2_U3503) );
  MUX2_X1 U9885 ( .A(n8235), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8297), .Z(
        P2_U3502) );
  MUX2_X1 U9886 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8236), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U9887 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8237), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U9888 ( .A(n8238), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8297), .Z(
        P2_U3499) );
  MUX2_X1 U9889 ( .A(n8239), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8297), .Z(
        P2_U3498) );
  MUX2_X1 U9890 ( .A(n8240), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8297), .Z(
        P2_U3497) );
  MUX2_X1 U9891 ( .A(n8241), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8297), .Z(
        P2_U3496) );
  MUX2_X1 U9892 ( .A(n8242), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8297), .Z(
        P2_U3495) );
  MUX2_X1 U9893 ( .A(n8243), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8297), .Z(
        P2_U3494) );
  MUX2_X1 U9894 ( .A(n8244), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8297), .Z(
        P2_U3493) );
  MUX2_X1 U9895 ( .A(n8245), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8297), .Z(
        P2_U3492) );
  MUX2_X1 U9896 ( .A(n8246), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8297), .Z(
        P2_U3491) );
  OR2_X1 U9897 ( .A1(n9952), .A2(n10418), .ZN(n8259) );
  INV_X1 U9898 ( .A(n8248), .ZN(n8249) );
  XNOR2_X1 U9899 ( .A(n8248), .B(n9843), .ZN(n9841) );
  NOR2_X1 U9900 ( .A1(n9841), .A2(n5848), .ZN(n9840) );
  NAND2_X1 U9901 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n8306), .ZN(n8250) );
  OAI21_X1 U9902 ( .B1(n8306), .B2(P2_REG2_REG_8__SCAN_IN), .A(n8250), .ZN(
        n9861) );
  NOR2_X1 U9903 ( .A1(n9862), .A2(n9861), .ZN(n9860) );
  AOI21_X2 U9904 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n8306), .A(n9860), .ZN(
        n8251) );
  NOR2_X1 U9905 ( .A1(n9872), .A2(n8251), .ZN(n8252) );
  XNOR2_X1 U9906 ( .A(n9872), .B(n8251), .ZN(n9882) );
  NAND2_X1 U9907 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n8305), .ZN(n8253) );
  OAI21_X1 U9908 ( .B1(n8305), .B2(P2_REG2_REG_10__SCAN_IN), .A(n8253), .ZN(
        n9898) );
  NOR2_X1 U9909 ( .A1(n9904), .A2(n8254), .ZN(n8255) );
  MUX2_X1 U9910 ( .A(n8257), .B(P2_REG2_REG_12__SCAN_IN), .S(n9919), .Z(n8256)
         );
  INV_X1 U9911 ( .A(n8256), .ZN(n9929) );
  XNOR2_X1 U9912 ( .A(n8258), .B(n8321), .ZN(n9944) );
  NOR2_X1 U9913 ( .A1(n9944), .A2(n5925), .ZN(n9947) );
  XNOR2_X1 U9914 ( .A(n8303), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n9962) );
  XNOR2_X1 U9915 ( .A(n8260), .B(n9969), .ZN(n9978) );
  XNOR2_X1 U9916 ( .A(n8302), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n9995) );
  NOR2_X1 U9917 ( .A1(n9996), .A2(n9995), .ZN(n9994) );
  NOR2_X1 U9918 ( .A1(n10003), .A2(n8262), .ZN(n8263) );
  XNOR2_X1 U9919 ( .A(n10003), .B(n8262), .ZN(n10014) );
  AOI22_X1 U9920 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8340), .B1(n8344), .B2(
        n5995), .ZN(n8264) );
  AOI21_X1 U9921 ( .B1(n4575), .B2(n8264), .A(n8336), .ZN(n8335) );
  MUX2_X1 U9922 ( .A(n10013), .B(n8265), .S(n8291), .Z(n8290) );
  XNOR2_X1 U9923 ( .A(n8290), .B(n8328), .ZN(n10008) );
  MUX2_X1 U9924 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8291), .Z(n8266) );
  OR2_X1 U9925 ( .A1(n8266), .A2(n8302), .ZN(n8288) );
  XNOR2_X1 U9926 ( .A(n8266), .B(n9985), .ZN(n9991) );
  MUX2_X1 U9927 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8291), .Z(n8267) );
  OR2_X1 U9928 ( .A1(n8267), .A2(n8324), .ZN(n8287) );
  XNOR2_X1 U9929 ( .A(n8267), .B(n9969), .ZN(n9974) );
  MUX2_X1 U9930 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8291), .Z(n8268) );
  OR2_X1 U9931 ( .A1(n8268), .A2(n8303), .ZN(n8286) );
  XNOR2_X1 U9932 ( .A(n8268), .B(n9952), .ZN(n9958) );
  MUX2_X1 U9933 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8291), .Z(n8269) );
  OR2_X1 U9934 ( .A1(n8269), .A2(n8321), .ZN(n8285) );
  XNOR2_X1 U9935 ( .A(n8269), .B(n9936), .ZN(n9941) );
  MUX2_X1 U9936 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8291), .Z(n8270) );
  OR2_X1 U9937 ( .A1(n8270), .A2(n8304), .ZN(n8284) );
  XNOR2_X1 U9938 ( .A(n8270), .B(n9919), .ZN(n9925) );
  MUX2_X1 U9939 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8291), .Z(n8271) );
  OR2_X1 U9940 ( .A1(n8271), .A2(n8318), .ZN(n8283) );
  XNOR2_X1 U9941 ( .A(n8271), .B(n9904), .ZN(n9909) );
  MUX2_X1 U9942 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8291), .Z(n8272) );
  OR2_X1 U9943 ( .A1(n8272), .A2(n8305), .ZN(n8282) );
  XNOR2_X1 U9944 ( .A(n8272), .B(n9888), .ZN(n9894) );
  MUX2_X1 U9945 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8291), .Z(n8273) );
  OR2_X1 U9946 ( .A1(n8273), .A2(n8314), .ZN(n8281) );
  XNOR2_X1 U9947 ( .A(n8273), .B(n9872), .ZN(n9877) );
  MUX2_X1 U9948 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8291), .Z(n8274) );
  OR2_X1 U9949 ( .A1(n8274), .A2(n8306), .ZN(n8280) );
  XNOR2_X1 U9950 ( .A(n8274), .B(n9855), .ZN(n9858) );
  MUX2_X1 U9951 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8291), .Z(n8275) );
  OR2_X1 U9952 ( .A1(n8275), .A2(n8310), .ZN(n8279) );
  XNOR2_X1 U9953 ( .A(n8275), .B(n9843), .ZN(n9849) );
  OAI21_X1 U9954 ( .B1(n8278), .B2(n8277), .A(n8276), .ZN(n9850) );
  NAND2_X1 U9955 ( .A1(n9849), .A2(n9850), .ZN(n9848) );
  NAND2_X1 U9956 ( .A1(n8279), .A2(n9848), .ZN(n9857) );
  NAND2_X1 U9957 ( .A1(n9858), .A2(n9857), .ZN(n9856) );
  NAND2_X1 U9958 ( .A1(n8280), .A2(n9856), .ZN(n9876) );
  NAND2_X1 U9959 ( .A1(n9877), .A2(n9876), .ZN(n9875) );
  NAND2_X1 U9960 ( .A1(n8281), .A2(n9875), .ZN(n9893) );
  NAND2_X1 U9961 ( .A1(n9894), .A2(n9893), .ZN(n9892) );
  NAND2_X1 U9962 ( .A1(n8282), .A2(n9892), .ZN(n9908) );
  NAND2_X1 U9963 ( .A1(n9909), .A2(n9908), .ZN(n9907) );
  NAND2_X1 U9964 ( .A1(n8283), .A2(n9907), .ZN(n9924) );
  NAND2_X1 U9965 ( .A1(n9925), .A2(n9924), .ZN(n9923) );
  NAND2_X1 U9966 ( .A1(n8284), .A2(n9923), .ZN(n9940) );
  NAND2_X1 U9967 ( .A1(n9941), .A2(n9940), .ZN(n9939) );
  NAND2_X1 U9968 ( .A1(n8285), .A2(n9939), .ZN(n9957) );
  NAND2_X1 U9969 ( .A1(n9958), .A2(n9957), .ZN(n9956) );
  NAND2_X1 U9970 ( .A1(n8286), .A2(n9956), .ZN(n9973) );
  NAND2_X1 U9971 ( .A1(n9974), .A2(n9973), .ZN(n9972) );
  NAND2_X1 U9972 ( .A1(n8287), .A2(n9972), .ZN(n9990) );
  NAND2_X1 U9973 ( .A1(n10008), .A2(n10007), .ZN(n10006) );
  INV_X1 U9974 ( .A(n10006), .ZN(n8289) );
  AOI21_X1 U9975 ( .B1(n8290), .B2(n10003), .A(n8289), .ZN(n8292) );
  MUX2_X1 U9976 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8291), .Z(n8293) );
  INV_X1 U9977 ( .A(n8292), .ZN(n8295) );
  INV_X1 U9978 ( .A(n8293), .ZN(n8294) );
  NAND2_X1 U9979 ( .A1(n8295), .A2(n8294), .ZN(n8343) );
  NAND2_X1 U9980 ( .A1(n8296), .A2(n8343), .ZN(n8298) );
  AND2_X1 U9981 ( .A1(n8298), .A2(n10010), .ZN(n8299) );
  AOI211_X1 U9982 ( .C1(n10159), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8301), .B(
        n8300), .ZN(n8334) );
  AOI22_X1 U9983 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n8344), .B1(n8340), .B2(
        n8588), .ZN(n8331) );
  AOI22_X1 U9984 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8302), .B1(n9985), .B2(
        n10323), .ZN(n9988) );
  AOI22_X1 U9985 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8303), .B1(n9952), .B2(
        n5942), .ZN(n9955) );
  AOI22_X1 U9986 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8304), .B1(n9919), .B2(
        n5916), .ZN(n9922) );
  NAND2_X1 U9987 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n8305), .ZN(n8317) );
  AOI22_X1 U9988 ( .A1(n9888), .A2(n5885), .B1(P2_REG1_REG_10__SCAN_IN), .B2(
        n8305), .ZN(n9891) );
  NAND2_X1 U9989 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n8306), .ZN(n8313) );
  AOI22_X1 U9990 ( .A1(n9855), .A2(n5834), .B1(P2_REG1_REG_8__SCAN_IN), .B2(
        n8306), .ZN(n9865) );
  NAND2_X1 U9991 ( .A1(n8310), .A2(n8311), .ZN(n8312) );
  NAND2_X1 U9992 ( .A1(n9865), .A2(n9866), .ZN(n9864) );
  NAND2_X1 U9993 ( .A1(n8314), .A2(n8315), .ZN(n8316) );
  NAND2_X1 U9994 ( .A1(n9891), .A2(n9890), .ZN(n9889) );
  NAND2_X1 U9995 ( .A1(n8318), .A2(n8319), .ZN(n8320) );
  NAND2_X1 U9996 ( .A1(n9922), .A2(n9921), .ZN(n9920) );
  NAND2_X1 U9997 ( .A1(n8322), .A2(n8321), .ZN(n8323) );
  NAND2_X1 U9998 ( .A1(n9955), .A2(n9954), .ZN(n9953) );
  OAI21_X1 U9999 ( .B1(n9952), .B2(n5942), .A(n9953), .ZN(n8325) );
  NAND2_X1 U10000 ( .A1(n8325), .A2(n8324), .ZN(n8326) );
  XNOR2_X1 U10001 ( .A(n8325), .B(n9969), .ZN(n9971) );
  NAND2_X1 U10002 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n9971), .ZN(n9970) );
  NAND2_X1 U10003 ( .A1(n8326), .A2(n9970), .ZN(n9987) );
  NAND2_X1 U10004 ( .A1(n8328), .A2(n8327), .ZN(n8329) );
  NAND2_X1 U10005 ( .A1(n8329), .A2(n10004), .ZN(n8330) );
  NAND2_X1 U10006 ( .A1(n8331), .A2(n8330), .ZN(n8339) );
  OAI21_X1 U10007 ( .B1(n8331), .B2(n8330), .A(n8339), .ZN(n8332) );
  NAND2_X1 U10008 ( .A1(n8332), .A2(n10153), .ZN(n8333) );
  OAI211_X1 U10009 ( .C1(n8335), .C2(n10147), .A(n8334), .B(n8333), .ZN(
        P2_U3200) );
  XNOR2_X1 U10010 ( .A(n8353), .B(n8337), .ZN(n8345) );
  XNOR2_X1 U10011 ( .A(n8338), .B(n8345), .ZN(n8358) );
  XNOR2_X1 U10012 ( .A(n8353), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8348) );
  OAI21_X1 U10013 ( .B1(n8340), .B2(n8588), .A(n8339), .ZN(n8341) );
  XOR2_X1 U10014 ( .A(n8348), .B(n8341), .Z(n8356) );
  AOI21_X1 U10015 ( .B1(n8344), .B2(n8343), .A(n8342), .ZN(n8350) );
  INV_X1 U10016 ( .A(n8345), .ZN(n8347) );
  MUX2_X1 U10017 ( .A(n8348), .B(n8347), .S(n8346), .Z(n8349) );
  NAND2_X1 U10018 ( .A1(n10159), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8352) );
  NAND2_X1 U10019 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3151), .ZN(n8351) );
  OAI211_X1 U10020 ( .C1(n10157), .C2(n8353), .A(n8352), .B(n8351), .ZN(n8354)
         );
  AOI211_X1 U10021 ( .C1(n8356), .C2(n10153), .A(n8355), .B(n8354), .ZN(n8357)
         );
  OAI21_X1 U10022 ( .B1(n8358), .B2(n10147), .A(n8357), .ZN(P2_U3201) );
  NOR2_X1 U10023 ( .A1(n8361), .A2(n10022), .ZN(n8370) );
  AOI21_X1 U10024 ( .B1(n8606), .B2(n10035), .A(n8370), .ZN(n8365) );
  NAND2_X1 U10025 ( .A1(n10038), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8362) );
  OAI211_X1 U10026 ( .C1(n8363), .C2(n8532), .A(n8365), .B(n8362), .ZN(
        P2_U3202) );
  INV_X1 U10027 ( .A(n8610), .ZN(n8543) );
  NAND2_X1 U10028 ( .A1(n10038), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8364) );
  OAI211_X1 U10029 ( .C1(n8543), .C2(n8532), .A(n8365), .B(n8364), .ZN(
        P2_U3203) );
  INV_X1 U10030 ( .A(n8366), .ZN(n8374) );
  NAND2_X1 U10031 ( .A1(n8367), .A2(n10035), .ZN(n8372) );
  NOR2_X1 U10032 ( .A1(n8368), .A2(n8532), .ZN(n8369) );
  AOI211_X1 U10033 ( .C1(n10038), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8370), .B(
        n8369), .ZN(n8371) );
  OAI211_X1 U10034 ( .C1(n8374), .C2(n8373), .A(n8372), .B(n8371), .ZN(
        P2_U3204) );
  INV_X1 U10035 ( .A(n8375), .ZN(n8381) );
  AOI22_X1 U10036 ( .A1(n8376), .A2(n8505), .B1(n10038), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8377) );
  OAI21_X1 U10037 ( .B1(n4731), .B2(n8532), .A(n8377), .ZN(n8378) );
  AOI21_X1 U10038 ( .B1(n8379), .B2(n8536), .A(n8378), .ZN(n8380) );
  OAI21_X1 U10039 ( .B1(n8381), .B2(n10038), .A(n8380), .ZN(P2_U3205) );
  INV_X1 U10040 ( .A(n8547), .ZN(n8391) );
  XOR2_X1 U10041 ( .A(n8385), .B(n8384), .Z(n8548) );
  INV_X1 U10042 ( .A(n8386), .ZN(n8617) );
  AOI22_X1 U10043 ( .A1(n8387), .A2(n8505), .B1(n10038), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8388) );
  OAI21_X1 U10044 ( .B1(n8617), .B2(n8532), .A(n8388), .ZN(n8389) );
  AOI21_X1 U10045 ( .B1(n8548), .B2(n8536), .A(n8389), .ZN(n8390) );
  OAI21_X1 U10046 ( .B1(n8391), .B2(n10038), .A(n8390), .ZN(P2_U3206) );
  XNOR2_X1 U10047 ( .A(n8393), .B(n8392), .ZN(n8394) );
  OAI222_X1 U10048 ( .A1(n10032), .A2(n8396), .B1(n10031), .B2(n8395), .C1(
        n8394), .C2(n10041), .ZN(n8551) );
  INV_X1 U10049 ( .A(n8551), .ZN(n8403) );
  XNOR2_X1 U10050 ( .A(n8398), .B(n8397), .ZN(n8552) );
  AOI22_X1 U10051 ( .A1(n8399), .A2(n8505), .B1(n10038), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8400) );
  OAI21_X1 U10052 ( .B1(n8621), .B2(n8532), .A(n8400), .ZN(n8401) );
  AOI21_X1 U10053 ( .B1(n8552), .B2(n8536), .A(n8401), .ZN(n8402) );
  OAI21_X1 U10054 ( .B1(n8403), .B2(n10038), .A(n8402), .ZN(P2_U3207) );
  INV_X1 U10055 ( .A(n10023), .ZN(n8420) );
  XOR2_X1 U10056 ( .A(n8404), .B(n8410), .Z(n8405) );
  OAI222_X1 U10057 ( .A1(n10032), .A2(n8406), .B1(n10031), .B2(n8436), .C1(
        n10041), .C2(n8405), .ZN(n8555) );
  AOI21_X1 U10058 ( .B1(n8420), .B2(n8407), .A(n8555), .ZN(n8413) );
  AOI22_X1 U10059 ( .A1(n8408), .A2(n8505), .B1(n10038), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8412) );
  XOR2_X1 U10060 ( .A(n8410), .B(n8409), .Z(n8556) );
  NAND2_X1 U10061 ( .A1(n8556), .A2(n8536), .ZN(n8411) );
  OAI211_X1 U10062 ( .C1(n8413), .C2(n10038), .A(n8412), .B(n8411), .ZN(
        P2_U3208) );
  XNOR2_X1 U10063 ( .A(n8414), .B(n8426), .ZN(n8418) );
  NAND2_X1 U10064 ( .A1(n8415), .A2(n8511), .ZN(n8416) );
  OAI21_X1 U10065 ( .B1(n8447), .B2(n10031), .A(n8416), .ZN(n8417) );
  AOI21_X1 U10066 ( .B1(n8418), .B2(n8516), .A(n8417), .ZN(n8561) );
  AOI22_X1 U10067 ( .A1(n8421), .A2(n8420), .B1(n8505), .B2(n8419), .ZN(n8422)
         );
  AND2_X1 U10068 ( .A1(n8561), .A2(n8422), .ZN(n8429) );
  INV_X1 U10069 ( .A(n8423), .ZN(n8424) );
  OR2_X1 U10070 ( .A1(n8425), .A2(n8424), .ZN(n8427) );
  XNOR2_X1 U10071 ( .A(n8427), .B(n8426), .ZN(n8559) );
  AOI22_X1 U10072 ( .A1(n8559), .A2(n8536), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n10038), .ZN(n8428) );
  OAI21_X1 U10073 ( .B1(n8429), .B2(n10038), .A(n8428), .ZN(P2_U3209) );
  NAND2_X1 U10074 ( .A1(n8455), .A2(n8454), .ZN(n8431) );
  NAND2_X1 U10075 ( .A1(n8431), .A2(n8430), .ZN(n8445) );
  NAND2_X1 U10076 ( .A1(n8445), .A2(n8449), .ZN(n8433) );
  NAND2_X1 U10077 ( .A1(n8433), .A2(n8432), .ZN(n8434) );
  XOR2_X1 U10078 ( .A(n8437), .B(n8434), .Z(n8435) );
  OAI222_X1 U10079 ( .A1(n10031), .A2(n8457), .B1(n10032), .B2(n8436), .C1(
        n10041), .C2(n8435), .ZN(n8564) );
  INV_X1 U10080 ( .A(n8564), .ZN(n8443) );
  XOR2_X1 U10081 ( .A(n8437), .B(n4523), .Z(n8565) );
  INV_X1 U10082 ( .A(n8438), .ZN(n8632) );
  AOI22_X1 U10083 ( .A1(n10038), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8439), 
        .B2(n8505), .ZN(n8440) );
  OAI21_X1 U10084 ( .B1(n8632), .B2(n8532), .A(n8440), .ZN(n8441) );
  AOI21_X1 U10085 ( .B1(n8565), .B2(n8536), .A(n8441), .ZN(n8442) );
  OAI21_X1 U10086 ( .B1(n8443), .B2(n10038), .A(n8442), .ZN(P2_U3210) );
  XNOR2_X1 U10087 ( .A(n8445), .B(n8444), .ZN(n8446) );
  OAI222_X1 U10088 ( .A1(n10032), .A2(n8447), .B1(n10031), .B2(n8478), .C1(
        n10041), .C2(n8446), .ZN(n8569) );
  AOI21_X1 U10089 ( .B1(n8505), .B2(n8448), .A(n8569), .ZN(n8453) );
  AOI22_X1 U10090 ( .A1(n8568), .A2(n8519), .B1(P2_REG2_REG_22__SCAN_IN), .B2(
        n10038), .ZN(n8452) );
  XNOR2_X1 U10091 ( .A(n8450), .B(n8449), .ZN(n8570) );
  NAND2_X1 U10092 ( .A1(n8570), .A2(n8536), .ZN(n8451) );
  OAI211_X1 U10093 ( .C1(n8453), .C2(n10038), .A(n8452), .B(n8451), .ZN(
        P2_U3211) );
  XNOR2_X1 U10094 ( .A(n8455), .B(n8454), .ZN(n8459) );
  OAI22_X1 U10095 ( .A1(n8457), .A2(n10032), .B1(n8456), .B2(n10031), .ZN(
        n8458) );
  AOI21_X1 U10096 ( .B1(n8459), .B2(n8516), .A(n8458), .ZN(n8575) );
  NAND2_X1 U10097 ( .A1(n8461), .A2(n8460), .ZN(n8463) );
  XNOR2_X1 U10098 ( .A(n8463), .B(n8462), .ZN(n8573) );
  INV_X1 U10099 ( .A(n8464), .ZN(n8639) );
  AOI22_X1 U10100 ( .A1(n10038), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8505), 
        .B2(n8465), .ZN(n8466) );
  OAI21_X1 U10101 ( .B1(n8639), .B2(n8532), .A(n8466), .ZN(n8467) );
  AOI21_X1 U10102 ( .B1(n8573), .B2(n8536), .A(n8467), .ZN(n8468) );
  OAI21_X1 U10103 ( .B1(n8575), .B2(n10038), .A(n8468), .ZN(P2_U3212) );
  XNOR2_X1 U10104 ( .A(n8469), .B(n8474), .ZN(n8578) );
  INV_X1 U10105 ( .A(n8470), .ZN(n8643) );
  AOI22_X1 U10106 ( .A1(n10038), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8505), 
        .B2(n8471), .ZN(n8472) );
  OAI21_X1 U10107 ( .B1(n8643), .B2(n8532), .A(n8472), .ZN(n8481) );
  OAI21_X1 U10108 ( .B1(n8475), .B2(n8474), .A(n8473), .ZN(n8477) );
  NOR2_X1 U10109 ( .A1(n8497), .A2(n10031), .ZN(n8476) );
  AOI21_X1 U10110 ( .B1(n8477), .B2(n8516), .A(n8476), .ZN(n8580) );
  NOR2_X1 U10111 ( .A1(n8478), .A2(n10032), .ZN(n8577) );
  INV_X1 U10112 ( .A(n8577), .ZN(n8479) );
  AOI21_X1 U10113 ( .B1(n8580), .B2(n8479), .A(n10038), .ZN(n8480) );
  AOI211_X1 U10114 ( .C1(n8536), .C2(n8578), .A(n8481), .B(n8480), .ZN(n8482)
         );
  INV_X1 U10115 ( .A(n8482), .ZN(P2_U3213) );
  OAI211_X1 U10116 ( .C1(n8484), .C2(n6159), .A(n8483), .B(n8516), .ZN(n8487)
         );
  AOI22_X1 U10117 ( .A1(n8485), .A2(n8511), .B1(n8513), .B2(n8512), .ZN(n8486)
         );
  NAND2_X1 U10118 ( .A1(n8487), .A2(n8486), .ZN(n8582) );
  INV_X1 U10119 ( .A(n8582), .ZN(n8494) );
  XNOR2_X1 U10120 ( .A(n8488), .B(n6159), .ZN(n8583) );
  INV_X1 U10121 ( .A(n8489), .ZN(n8646) );
  AOI22_X1 U10122 ( .A1(n10038), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8505), 
        .B2(n8490), .ZN(n8491) );
  OAI21_X1 U10123 ( .B1(n8646), .B2(n8532), .A(n8491), .ZN(n8492) );
  AOI21_X1 U10124 ( .B1(n8583), .B2(n8536), .A(n8492), .ZN(n8493) );
  OAI21_X1 U10125 ( .B1(n8494), .B2(n10038), .A(n8493), .ZN(P2_U3214) );
  XNOR2_X1 U10126 ( .A(n8495), .B(n8502), .ZN(n8496) );
  OAI222_X1 U10127 ( .A1(n10031), .A2(n8528), .B1(n10032), .B2(n8497), .C1(
        n8496), .C2(n10041), .ZN(n8586) );
  INV_X1 U10128 ( .A(n8586), .ZN(n8509) );
  NAND2_X1 U10129 ( .A1(n8520), .A2(n8498), .ZN(n8501) );
  INV_X1 U10130 ( .A(n8499), .ZN(n8500) );
  AOI21_X1 U10131 ( .B1(n8502), .B2(n8501), .A(n8500), .ZN(n8587) );
  INV_X1 U10132 ( .A(n8503), .ZN(n8649) );
  AOI22_X1 U10133 ( .A1(n10038), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8505), 
        .B2(n8504), .ZN(n8506) );
  OAI21_X1 U10134 ( .B1(n8649), .B2(n8532), .A(n8506), .ZN(n8507) );
  AOI21_X1 U10135 ( .B1(n8587), .B2(n8536), .A(n8507), .ZN(n8508) );
  OAI21_X1 U10136 ( .B1(n8509), .B2(n10038), .A(n8508), .ZN(P2_U3215) );
  XNOR2_X1 U10137 ( .A(n8510), .B(n8521), .ZN(n8515) );
  AOI222_X1 U10138 ( .A1(n8516), .A2(n8515), .B1(n8514), .B2(n8513), .C1(n8512), .C2(n8511), .ZN(n8593) );
  OAI22_X1 U10139 ( .A1(n10035), .A2(n10013), .B1(n8517), .B2(n10022), .ZN(
        n8518) );
  AOI21_X1 U10140 ( .B1(n8590), .B2(n8519), .A(n8518), .ZN(n8524) );
  OAI21_X1 U10141 ( .B1(n8522), .B2(n8521), .A(n8520), .ZN(n8591) );
  NAND2_X1 U10142 ( .A1(n8591), .A2(n8536), .ZN(n8523) );
  OAI211_X1 U10143 ( .C1(n8593), .C2(n10038), .A(n8524), .B(n8523), .ZN(
        P2_U3216) );
  XNOR2_X1 U10144 ( .A(n8525), .B(n8529), .ZN(n8526) );
  OAI222_X1 U10145 ( .A1(n10032), .A2(n8528), .B1(n10031), .B2(n8527), .C1(
        n10041), .C2(n8526), .ZN(n8594) );
  INV_X1 U10146 ( .A(n8594), .ZN(n8538) );
  XOR2_X1 U10147 ( .A(n8530), .B(n8529), .Z(n8595) );
  INV_X1 U10148 ( .A(n8531), .ZN(n8654) );
  NOR2_X1 U10149 ( .A1(n8654), .A2(n8532), .ZN(n8535) );
  OAI22_X1 U10150 ( .A1(n10035), .A2(n10375), .B1(n8533), .B2(n10022), .ZN(
        n8534) );
  AOI211_X1 U10151 ( .C1(n8595), .C2(n8536), .A(n8535), .B(n8534), .ZN(n8537)
         );
  OAI21_X1 U10152 ( .B1(n8538), .B2(n10038), .A(n8537), .ZN(P2_U3217) );
  NAND2_X1 U10153 ( .A1(n8605), .A2(n8539), .ZN(n8540) );
  NAND2_X1 U10154 ( .A1(n8606), .A2(n10105), .ZN(n8541) );
  OAI211_X1 U10155 ( .C1(n10105), .C2(n7223), .A(n8540), .B(n8541), .ZN(
        P2_U3490) );
  NAND2_X1 U10156 ( .A1(n10103), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8542) );
  OAI211_X1 U10157 ( .C1(n8543), .C2(n8604), .A(n8542), .B(n8541), .ZN(
        P2_U3489) );
  MUX2_X1 U10158 ( .A(n8545), .B(n8544), .S(n10105), .Z(n8546) );
  OAI21_X1 U10159 ( .B1(n4731), .B2(n8604), .A(n8546), .ZN(P2_U3487) );
  AOI21_X1 U10160 ( .B1(n8548), .B2(n10082), .A(n8547), .ZN(n8614) );
  OAI21_X1 U10161 ( .B1(n8617), .B2(n8604), .A(n8550), .ZN(P2_U3486) );
  AOI21_X1 U10162 ( .B1(n10082), .B2(n8552), .A(n8551), .ZN(n8618) );
  MUX2_X1 U10163 ( .A(n8553), .B(n8618), .S(n10105), .Z(n8554) );
  OAI21_X1 U10164 ( .B1(n8621), .B2(n8604), .A(n8554), .ZN(P2_U3485) );
  INV_X1 U10165 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8557) );
  AOI21_X1 U10166 ( .B1(n10082), .B2(n8556), .A(n8555), .ZN(n8622) );
  MUX2_X1 U10167 ( .A(n8557), .B(n8622), .S(n10105), .Z(n8558) );
  OAI21_X1 U10168 ( .B1(n8624), .B2(n8604), .A(n8558), .ZN(P2_U3484) );
  INV_X1 U10169 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8562) );
  NAND2_X1 U10170 ( .A1(n8559), .A2(n10082), .ZN(n8560) );
  AND2_X1 U10171 ( .A1(n8561), .A2(n8560), .ZN(n8625) );
  MUX2_X1 U10172 ( .A(n8562), .B(n8625), .S(n10105), .Z(n8563) );
  OAI21_X1 U10173 ( .B1(n8628), .B2(n8604), .A(n8563), .ZN(P2_U3483) );
  AOI21_X1 U10174 ( .B1(n10082), .B2(n8565), .A(n8564), .ZN(n8629) );
  MUX2_X1 U10175 ( .A(n8566), .B(n8629), .S(n10105), .Z(n8567) );
  OAI21_X1 U10176 ( .B1(n8632), .B2(n8604), .A(n8567), .ZN(P2_U3482) );
  INV_X1 U10177 ( .A(n8568), .ZN(n8636) );
  INV_X1 U10178 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8571) );
  AOI21_X1 U10179 ( .B1(n10082), .B2(n8570), .A(n8569), .ZN(n8633) );
  MUX2_X1 U10180 ( .A(n8571), .B(n8633), .S(n10105), .Z(n8572) );
  OAI21_X1 U10181 ( .B1(n8636), .B2(n8604), .A(n8572), .ZN(P2_U3481) );
  INV_X1 U10182 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n10310) );
  NAND2_X1 U10183 ( .A1(n8573), .A2(n10082), .ZN(n8574) );
  AND2_X1 U10184 ( .A1(n8575), .A2(n8574), .ZN(n8637) );
  MUX2_X1 U10185 ( .A(n10310), .B(n8637), .S(n10105), .Z(n8576) );
  OAI21_X1 U10186 ( .B1(n8639), .B2(n8604), .A(n8576), .ZN(P2_U3480) );
  AOI21_X1 U10187 ( .B1(n8578), .B2(n10082), .A(n8577), .ZN(n8579) );
  AND2_X1 U10188 ( .A1(n8580), .A2(n8579), .ZN(n8640) );
  MUX2_X1 U10189 ( .A(n10234), .B(n8640), .S(n10105), .Z(n8581) );
  OAI21_X1 U10190 ( .B1(n8643), .B2(n8604), .A(n8581), .ZN(P2_U3479) );
  INV_X1 U10191 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8584) );
  AOI21_X1 U10192 ( .B1(n10082), .B2(n8583), .A(n8582), .ZN(n8644) );
  MUX2_X1 U10193 ( .A(n8584), .B(n8644), .S(n10105), .Z(n8585) );
  OAI21_X1 U10194 ( .B1(n8646), .B2(n8604), .A(n8585), .ZN(P2_U3478) );
  AOI21_X1 U10195 ( .B1(n8587), .B2(n10082), .A(n8586), .ZN(n8647) );
  MUX2_X1 U10196 ( .A(n8588), .B(n8647), .S(n10105), .Z(n8589) );
  OAI21_X1 U10197 ( .B1(n8649), .B2(n8604), .A(n8589), .ZN(P2_U3477) );
  AOI22_X1 U10198 ( .A1(n8591), .A2(n10082), .B1(n10090), .B2(n8590), .ZN(
        n8592) );
  NAND2_X1 U10199 ( .A1(n8593), .A2(n8592), .ZN(n8650) );
  MUX2_X1 U10200 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8650), .S(n10105), .Z(
        P2_U3476) );
  AOI21_X1 U10201 ( .B1(n10082), .B2(n8595), .A(n8594), .ZN(n8651) );
  MUX2_X1 U10202 ( .A(n10323), .B(n8651), .S(n10105), .Z(n8596) );
  OAI21_X1 U10203 ( .B1(n8654), .B2(n8604), .A(n8596), .ZN(P2_U3475) );
  AOI21_X1 U10204 ( .B1(n10082), .B2(n8598), .A(n8597), .ZN(n8655) );
  MUX2_X1 U10205 ( .A(n8599), .B(n8655), .S(n10105), .Z(n8600) );
  OAI21_X1 U10206 ( .B1(n8658), .B2(n8604), .A(n8600), .ZN(P2_U3474) );
  AOI21_X1 U10207 ( .B1(n8602), .B2(n10082), .A(n8601), .ZN(n8659) );
  MUX2_X1 U10208 ( .A(n5942), .B(n8659), .S(n10105), .Z(n8603) );
  OAI21_X1 U10209 ( .B1(n8663), .B2(n8604), .A(n8603), .ZN(P2_U3473) );
  INV_X1 U10210 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U10211 ( .A1(n8605), .A2(n8609), .ZN(n8607) );
  NAND2_X1 U10212 ( .A1(n8606), .A2(n10091), .ZN(n8611) );
  OAI211_X1 U10213 ( .C1(n8608), .C2(n10091), .A(n8607), .B(n8611), .ZN(
        P2_U3458) );
  INV_X1 U10214 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8613) );
  NAND2_X1 U10215 ( .A1(n8610), .A2(n8609), .ZN(n8612) );
  OAI211_X1 U10216 ( .C1(n8613), .C2(n10091), .A(n8612), .B(n8611), .ZN(
        P2_U3457) );
  INV_X1 U10217 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8615) );
  OAI21_X1 U10218 ( .B1(n8617), .B2(n8662), .A(n8616), .ZN(P2_U3454) );
  INV_X1 U10219 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8619) );
  MUX2_X1 U10220 ( .A(n8619), .B(n8618), .S(n10091), .Z(n8620) );
  OAI21_X1 U10221 ( .B1(n8621), .B2(n8662), .A(n8620), .ZN(P2_U3453) );
  MUX2_X1 U10222 ( .A(n10297), .B(n8622), .S(n10091), .Z(n8623) );
  OAI21_X1 U10223 ( .B1(n8624), .B2(n8662), .A(n8623), .ZN(P2_U3452) );
  INV_X1 U10224 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8626) );
  MUX2_X1 U10225 ( .A(n8626), .B(n8625), .S(n10091), .Z(n8627) );
  OAI21_X1 U10226 ( .B1(n8628), .B2(n8662), .A(n8627), .ZN(P2_U3451) );
  INV_X1 U10227 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8630) );
  MUX2_X1 U10228 ( .A(n8630), .B(n8629), .S(n10091), .Z(n8631) );
  OAI21_X1 U10229 ( .B1(n8632), .B2(n8662), .A(n8631), .ZN(P2_U3450) );
  MUX2_X1 U10230 ( .A(n8634), .B(n8633), .S(n10091), .Z(n8635) );
  OAI21_X1 U10231 ( .B1(n8636), .B2(n8662), .A(n8635), .ZN(P2_U3449) );
  INV_X1 U10232 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n10410) );
  MUX2_X1 U10233 ( .A(n10410), .B(n8637), .S(n10091), .Z(n8638) );
  OAI21_X1 U10234 ( .B1(n8639), .B2(n8662), .A(n8638), .ZN(P2_U3448) );
  INV_X1 U10235 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8641) );
  MUX2_X1 U10236 ( .A(n8641), .B(n8640), .S(n10091), .Z(n8642) );
  OAI21_X1 U10237 ( .B1(n8643), .B2(n8662), .A(n8642), .ZN(P2_U3447) );
  MUX2_X1 U10238 ( .A(n10388), .B(n8644), .S(n10091), .Z(n8645) );
  OAI21_X1 U10239 ( .B1(n8646), .B2(n8662), .A(n8645), .ZN(P2_U3446) );
  MUX2_X1 U10240 ( .A(n10487), .B(n8647), .S(n10091), .Z(n8648) );
  OAI21_X1 U10241 ( .B1(n8649), .B2(n8662), .A(n8648), .ZN(P2_U3444) );
  MUX2_X1 U10242 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8650), .S(n10091), .Z(
        P2_U3441) );
  INV_X1 U10243 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8652) );
  MUX2_X1 U10244 ( .A(n8652), .B(n8651), .S(n10091), .Z(n8653) );
  OAI21_X1 U10245 ( .B1(n8654), .B2(n8662), .A(n8653), .ZN(P2_U3438) );
  INV_X1 U10246 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8656) );
  MUX2_X1 U10247 ( .A(n8656), .B(n8655), .S(n10091), .Z(n8657) );
  OAI21_X1 U10248 ( .B1(n8658), .B2(n8662), .A(n8657), .ZN(P2_U3435) );
  INV_X1 U10249 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8660) );
  MUX2_X1 U10250 ( .A(n8660), .B(n8659), .S(n10091), .Z(n8661) );
  OAI21_X1 U10251 ( .B1(n8663), .B2(n8662), .A(n8661), .ZN(P2_U3432) );
  INV_X1 U10252 ( .A(n8911), .ZN(n9565) );
  NOR4_X1 U10253 ( .A1(n8665), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n5905), .ZN(n8666) );
  AOI21_X1 U10254 ( .B1(n8673), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8666), .ZN(
        n8667) );
  OAI21_X1 U10255 ( .B1(n9565), .B2(n6582), .A(n8667), .ZN(P2_U3264) );
  INV_X1 U10256 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8669) );
  OAI222_X1 U10257 ( .A1(P2_U3151), .A2(n8670), .B1(n6582), .B2(n9568), .C1(
        n8669), .C2(n8668), .ZN(P2_U3266) );
  INV_X1 U10258 ( .A(n8671), .ZN(n9571) );
  AOI21_X1 U10259 ( .B1(n8673), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8672), .ZN(
        n8674) );
  OAI21_X1 U10260 ( .B1(n9571), .B2(n6582), .A(n8674), .ZN(P2_U3267) );
  MUX2_X1 U10261 ( .A(n8675), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10262 ( .A(n8676), .ZN(n8678) );
  NAND2_X1 U10263 ( .A1(n8678), .A2(n8677), .ZN(n8679) );
  XNOR2_X1 U10264 ( .A(n8750), .B(n8679), .ZN(n8685) );
  NAND2_X1 U10265 ( .A1(n9079), .A2(n9066), .ZN(n8681) );
  NAND2_X1 U10266 ( .A1(n9077), .A2(n8777), .ZN(n8680) );
  NAND2_X1 U10267 ( .A1(n8681), .A2(n8680), .ZN(n9458) );
  AOI22_X1 U10268 ( .A1(n9458), .A2(n8763), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n8682) );
  OAI21_X1 U10269 ( .B1(n9335), .B2(n8765), .A(n8682), .ZN(n8683) );
  AOI21_X1 U10270 ( .B1(n9459), .B2(n8767), .A(n8683), .ZN(n8684) );
  OAI21_X1 U10271 ( .B1(n8685), .B2(n8769), .A(n8684), .ZN(P1_U3216) );
  XNOR2_X1 U10272 ( .A(n8686), .B(n8687), .ZN(n8691) );
  AOI22_X1 U10273 ( .A1(n9081), .A2(n8777), .B1(n9066), .B2(n9083), .ZN(n9389)
         );
  NAND2_X1 U10274 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9238) );
  NAND2_X1 U10275 ( .A1(n8782), .A2(n9392), .ZN(n8688) );
  OAI211_X1 U10276 ( .C1(n9389), .C2(n8780), .A(n9238), .B(n8688), .ZN(n8689)
         );
  AOI21_X1 U10277 ( .B1(n9481), .B2(n8767), .A(n8689), .ZN(n8690) );
  OAI21_X1 U10278 ( .B1(n8691), .B2(n8769), .A(n8690), .ZN(P1_U3219) );
  OAI211_X1 U10279 ( .C1(n8694), .C2(n8693), .A(n8692), .B(n8775), .ZN(n8700)
         );
  NAND2_X1 U10280 ( .A1(n9079), .A2(n8777), .ZN(n8696) );
  NAND2_X1 U10281 ( .A1(n9081), .A2(n9066), .ZN(n8695) );
  NAND2_X1 U10282 ( .A1(n8696), .A2(n8695), .ZN(n9361) );
  OAI22_X1 U10283 ( .A1(n8765), .A2(n9365), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8697), .ZN(n8698) );
  AOI21_X1 U10284 ( .B1(n9361), .B2(n8763), .A(n8698), .ZN(n8699) );
  OAI211_X1 U10285 ( .C1(n9544), .C2(n8785), .A(n8700), .B(n8699), .ZN(
        P1_U3223) );
  AOI21_X1 U10286 ( .B1(n4526), .B2(n8701), .A(n8773), .ZN(n8706) );
  AOI22_X1 U10287 ( .A1(n9066), .A2(n9077), .B1(n9075), .B2(n8777), .ZN(n9303)
         );
  OAI22_X1 U10288 ( .A1(n8780), .A2(n9303), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8702), .ZN(n8704) );
  NOR2_X1 U10289 ( .A1(n9527), .A2(n8785), .ZN(n8703) );
  AOI211_X1 U10290 ( .C1(n8782), .C2(n9298), .A(n8704), .B(n8703), .ZN(n8705)
         );
  OAI21_X1 U10291 ( .B1(n8706), .B2(n8769), .A(n8705), .ZN(P1_U3225) );
  OAI21_X1 U10292 ( .B1(n8708), .B2(n8707), .A(n8716), .ZN(n8709) );
  NAND2_X1 U10293 ( .A1(n8709), .A2(n8775), .ZN(n8714) );
  AND2_X1 U10294 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9669) );
  NOR2_X1 U10295 ( .A1(n8765), .A2(n8710), .ZN(n8711) );
  AOI211_X1 U10296 ( .C1(n8763), .C2(n8712), .A(n9669), .B(n8711), .ZN(n8713)
         );
  OAI211_X1 U10297 ( .C1(n8715), .C2(n8785), .A(n8714), .B(n8713), .ZN(
        P1_U3226) );
  INV_X1 U10298 ( .A(n8716), .ZN(n8719) );
  NOR3_X1 U10299 ( .A1(n8719), .A2(n4627), .A3(n8718), .ZN(n8722) );
  INV_X1 U10300 ( .A(n8720), .ZN(n8721) );
  OAI21_X1 U10301 ( .B1(n8722), .B2(n8721), .A(n8775), .ZN(n8727) );
  INV_X1 U10302 ( .A(n8723), .ZN(n9424) );
  AND2_X1 U10303 ( .A1(n9085), .A2(n9066), .ZN(n8724) );
  AOI21_X1 U10304 ( .B1(n9083), .B2(n8777), .A(n8724), .ZN(n9419) );
  NAND2_X1 U10305 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9689) );
  OAI21_X1 U10306 ( .B1(n9419), .B2(n8780), .A(n9689), .ZN(n8725) );
  AOI21_X1 U10307 ( .B1(n9424), .B2(n8782), .A(n8725), .ZN(n8726) );
  OAI211_X1 U10308 ( .C1(n9427), .C2(n8785), .A(n8727), .B(n8726), .ZN(
        P1_U3228) );
  AOI21_X1 U10309 ( .B1(n8730), .B2(n8729), .A(n8728), .ZN(n8735) );
  AND2_X1 U10310 ( .A1(n9076), .A2(n8777), .ZN(n8731) );
  AOI21_X1 U10311 ( .B1(n9078), .B2(n9066), .A(n8731), .ZN(n9317) );
  AOI22_X1 U10312 ( .A1(n8782), .A2(n9322), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8732) );
  OAI21_X1 U10313 ( .B1(n9317), .B2(n8780), .A(n8732), .ZN(n8733) );
  AOI21_X1 U10314 ( .B1(n9323), .B2(n8767), .A(n8733), .ZN(n8734) );
  OAI21_X1 U10315 ( .B1(n8735), .B2(n8769), .A(n8734), .ZN(P1_U3229) );
  NAND2_X1 U10316 ( .A1(n8737), .A2(n8736), .ZN(n8739) );
  XOR2_X1 U10317 ( .A(n8739), .B(n8738), .Z(n8744) );
  AOI22_X1 U10318 ( .A1(n9080), .A2(n8777), .B1(n9066), .B2(n9082), .ZN(n9378)
         );
  OAI22_X1 U10319 ( .A1(n9378), .A2(n8780), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8740), .ZN(n8742) );
  NOR2_X1 U10320 ( .A1(n4773), .A2(n8785), .ZN(n8741) );
  AOI211_X1 U10321 ( .C1(n8782), .C2(n9381), .A(n8742), .B(n8741), .ZN(n8743)
         );
  OAI21_X1 U10322 ( .B1(n8744), .B2(n8769), .A(n8743), .ZN(P1_U3233) );
  INV_X1 U10323 ( .A(n8745), .ZN(n8747) );
  AOI21_X1 U10324 ( .B1(n8748), .B2(n8747), .A(n8746), .ZN(n8749) );
  AOI21_X1 U10325 ( .B1(n8750), .B2(n4917), .A(n8749), .ZN(n8756) );
  AND2_X1 U10326 ( .A1(n9080), .A2(n9066), .ZN(n8751) );
  AOI21_X1 U10327 ( .B1(n9078), .B2(n8777), .A(n8751), .ZN(n9344) );
  NOR2_X1 U10328 ( .A1(n9344), .A2(n8780), .ZN(n8754) );
  OAI22_X1 U10329 ( .A1(n9349), .A2(n8765), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8752), .ZN(n8753) );
  AOI211_X1 U10330 ( .C1(n9467), .C2(n8767), .A(n8754), .B(n8753), .ZN(n8755)
         );
  OAI21_X1 U10331 ( .B1(n8756), .B2(n8769), .A(n8755), .ZN(P1_U3235) );
  NAND2_X1 U10332 ( .A1(n8758), .A2(n8757), .ZN(n8759) );
  XOR2_X1 U10333 ( .A(n8760), .B(n8759), .Z(n8770) );
  NAND2_X1 U10334 ( .A1(n9082), .A2(n8777), .ZN(n8762) );
  NAND2_X1 U10335 ( .A1(n9084), .A2(n9066), .ZN(n8761) );
  NAND2_X1 U10336 ( .A1(n8762), .A2(n8761), .ZN(n9486) );
  AOI22_X1 U10337 ( .A1(n9486), .A2(n8763), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n8764) );
  OAI21_X1 U10338 ( .B1(n9406), .B2(n8765), .A(n8764), .ZN(n8766) );
  AOI21_X1 U10339 ( .B1(n9487), .B2(n8767), .A(n8766), .ZN(n8768) );
  OAI21_X1 U10340 ( .B1(n8770), .B2(n8769), .A(n8768), .ZN(P1_U3238) );
  OAI21_X1 U10341 ( .B1(n8773), .B2(n8772), .A(n8771), .ZN(n8774) );
  NAND3_X1 U10342 ( .A1(n8776), .A2(n8775), .A3(n8774), .ZN(n8784) );
  NAND2_X1 U10343 ( .A1(n9074), .A2(n8777), .ZN(n8779) );
  NAND2_X1 U10344 ( .A1(n9076), .A2(n9066), .ZN(n8778) );
  AND2_X1 U10345 ( .A1(n8779), .A2(n8778), .ZN(n9288) );
  OAI22_X1 U10346 ( .A1(n8780), .A2(n9288), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10439), .ZN(n8781) );
  AOI21_X1 U10347 ( .B1(n9291), .B2(n8782), .A(n8781), .ZN(n8783) );
  OAI211_X1 U10348 ( .C1(n8786), .C2(n8785), .A(n8784), .B(n8783), .ZN(
        P1_U3240) );
  INV_X1 U10349 ( .A(n8975), .ZN(n8788) );
  OAI22_X1 U10350 ( .A1(n9375), .A2(n9481), .B1(n8788), .B2(n8787), .ZN(n8872)
         );
  NAND2_X1 U10351 ( .A1(n8789), .A2(n9026), .ZN(n8791) );
  NAND3_X1 U10352 ( .A1(n8791), .A2(n8790), .A3(n8927), .ZN(n8792) );
  NAND2_X1 U10353 ( .A1(n8792), .A2(n9028), .ZN(n8794) );
  NAND2_X1 U10354 ( .A1(n8801), .A2(n8795), .ZN(n8797) );
  AOI21_X1 U10355 ( .B1(n8797), .B2(n8799), .A(n8796), .ZN(n8805) );
  INV_X1 U10356 ( .A(n8798), .ZN(n8800) );
  OAI21_X1 U10357 ( .B1(n8801), .B2(n8800), .A(n8799), .ZN(n8803) );
  NAND2_X1 U10358 ( .A1(n8803), .A2(n8802), .ZN(n8804) );
  INV_X1 U10359 ( .A(n8807), .ZN(n8809) );
  MUX2_X1 U10360 ( .A(n8809), .B(n8808), .S(n4789), .Z(n8810) );
  MUX2_X1 U10361 ( .A(n8812), .B(n8811), .S(n8919), .Z(n8813) );
  NAND2_X1 U10362 ( .A1(n8834), .A2(n8831), .ZN(n8814) );
  NAND3_X1 U10363 ( .A1(n8814), .A2(n8833), .A3(n9713), .ZN(n8815) );
  NAND3_X1 U10364 ( .A1(n8815), .A2(n8836), .A3(n9033), .ZN(n8820) );
  AND2_X1 U10365 ( .A1(n8842), .A2(n8835), .ZN(n8819) );
  NOR2_X1 U10366 ( .A1(n8845), .A2(n8846), .ZN(n9044) );
  INV_X1 U10367 ( .A(n9044), .ZN(n8816) );
  NAND4_X1 U10368 ( .A1(n8817), .A2(n4789), .A3(n8837), .A4(n8816), .ZN(n8818)
         );
  AOI21_X1 U10369 ( .B1(n8820), .B2(n8819), .A(n8818), .ZN(n8830) );
  NAND3_X1 U10370 ( .A1(n8845), .A2(n8846), .A3(n4789), .ZN(n8822) );
  NAND2_X1 U10371 ( .A1(n8821), .A2(n4789), .ZN(n8825) );
  NAND2_X1 U10372 ( .A1(n8822), .A2(n8825), .ZN(n8823) );
  NAND2_X1 U10373 ( .A1(n8824), .A2(n8823), .ZN(n8828) );
  INV_X1 U10374 ( .A(n8825), .ZN(n8826) );
  NAND3_X1 U10375 ( .A1(n8845), .A2(n8846), .A3(n8826), .ZN(n8827) );
  NAND2_X1 U10376 ( .A1(n8828), .A2(n8827), .ZN(n8829) );
  OAI21_X1 U10377 ( .B1(n8830), .B2(n8829), .A(n9018), .ZN(n8858) );
  NAND2_X1 U10378 ( .A1(n9033), .A2(n8831), .ZN(n8832) );
  AOI21_X1 U10379 ( .B1(n8834), .B2(n8833), .A(n8832), .ZN(n8840) );
  AND2_X1 U10380 ( .A1(n8835), .A2(n9713), .ZN(n9037) );
  INV_X1 U10381 ( .A(n9037), .ZN(n8839) );
  NAND2_X1 U10382 ( .A1(n8837), .A2(n8836), .ZN(n9036) );
  INV_X1 U10383 ( .A(n9036), .ZN(n8838) );
  OAI21_X1 U10384 ( .B1(n8840), .B2(n8839), .A(n8838), .ZN(n8854) );
  AND4_X1 U10385 ( .A1(n8843), .A2(n8842), .A3(n8841), .A4(n8919), .ZN(n8853)
         );
  NAND2_X1 U10386 ( .A1(n9088), .A2(n8919), .ZN(n8844) );
  NAND2_X1 U10387 ( .A1(n9087), .A2(n8919), .ZN(n8847) );
  OAI21_X1 U10388 ( .B1(n8845), .B2(n8844), .A(n8847), .ZN(n8850) );
  NOR2_X1 U10389 ( .A1(n8847), .A2(n8846), .ZN(n8848) );
  AOI22_X1 U10390 ( .A1(n9506), .A2(n8850), .B1(n8849), .B2(n8848), .ZN(n8851)
         );
  NAND2_X1 U10391 ( .A1(n8851), .A2(n9017), .ZN(n8852) );
  AOI21_X1 U10392 ( .B1(n8854), .B2(n8853), .A(n8852), .ZN(n8857) );
  NAND2_X1 U10393 ( .A1(n9015), .A2(n8855), .ZN(n9014) );
  NAND2_X1 U10394 ( .A1(n9014), .A2(n9018), .ZN(n8859) );
  OR2_X1 U10395 ( .A1(n9018), .A2(n4789), .ZN(n8856) );
  NAND4_X1 U10396 ( .A1(n8858), .A2(n8857), .A3(n8859), .A4(n8856), .ZN(n8865)
         );
  OAI21_X1 U10397 ( .B1(n8919), .B2(n8860), .A(n8859), .ZN(n8863) );
  NAND2_X1 U10398 ( .A1(n9015), .A2(n9086), .ZN(n8861) );
  NAND2_X1 U10399 ( .A1(n8861), .A2(n4789), .ZN(n8862) );
  NAND2_X1 U10400 ( .A1(n8863), .A2(n8862), .ZN(n8864) );
  NAND2_X1 U10401 ( .A1(n8865), .A2(n8864), .ZN(n8866) );
  NAND2_X1 U10402 ( .A1(n8866), .A2(n9417), .ZN(n8878) );
  NAND3_X1 U10403 ( .A1(n8878), .A2(n8874), .A3(n8867), .ZN(n8868) );
  NAND3_X1 U10404 ( .A1(n8868), .A2(n9048), .A3(n8877), .ZN(n8869) );
  NAND3_X1 U10405 ( .A1(n8883), .A2(n8875), .A3(n8869), .ZN(n8870) );
  NAND3_X1 U10406 ( .A1(n8976), .A2(n8975), .A3(n8870), .ZN(n8871) );
  MUX2_X1 U10407 ( .A(n8872), .B(n8871), .S(n4789), .Z(n8882) );
  NOR2_X1 U10408 ( .A1(n9367), .A2(n8873), .ZN(n8971) );
  INV_X1 U10409 ( .A(n8971), .ZN(n8884) );
  NAND2_X1 U10410 ( .A1(n8875), .A2(n8874), .ZN(n9049) );
  INV_X1 U10411 ( .A(n9049), .ZN(n8881) );
  NAND2_X1 U10412 ( .A1(n8877), .A2(n8876), .ZN(n9045) );
  INV_X1 U10413 ( .A(n9045), .ZN(n8879) );
  AOI21_X1 U10414 ( .B1(n8879), .B2(n8878), .A(n4789), .ZN(n8880) );
  NAND2_X1 U10415 ( .A1(n8884), .A2(n8883), .ZN(n8962) );
  NOR2_X1 U10416 ( .A1(n8976), .A2(n4789), .ZN(n8885) );
  OR2_X1 U10417 ( .A1(n9467), .A2(n8886), .ZN(n8887) );
  NAND2_X1 U10418 ( .A1(n8890), .A2(n8887), .ZN(n8964) );
  NAND2_X1 U10419 ( .A1(n8964), .A2(n4789), .ZN(n8888) );
  AND2_X1 U10420 ( .A1(n9312), .A2(n8889), .ZN(n8972) );
  INV_X1 U10421 ( .A(n8972), .ZN(n8978) );
  MUX2_X1 U10422 ( .A(n9300), .B(n8974), .S(n8919), .Z(n8891) );
  NAND2_X1 U10423 ( .A1(n8892), .A2(n8891), .ZN(n8897) );
  INV_X1 U10424 ( .A(n8968), .ZN(n8894) );
  INV_X1 U10425 ( .A(n8993), .ZN(n9274) );
  NOR2_X1 U10426 ( .A1(n9446), .A2(n8895), .ZN(n8981) );
  INV_X1 U10427 ( .A(n8981), .ZN(n8896) );
  OAI21_X1 U10428 ( .B1(n8986), .B2(n8899), .A(n8985), .ZN(n8900) );
  NAND2_X1 U10429 ( .A1(n8900), .A2(n8919), .ZN(n8901) );
  NAND2_X1 U10430 ( .A1(n8902), .A2(n8901), .ZN(n8903) );
  NAND2_X1 U10431 ( .A1(n8903), .A2(n8957), .ZN(n8915) );
  MUX2_X1 U10432 ( .A(n8904), .B(n8988), .S(n4789), .Z(n8914) );
  NAND2_X1 U10433 ( .A1(n8905), .A2(n8910), .ZN(n8908) );
  NAND2_X1 U10434 ( .A1(n8906), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8907) );
  AND2_X1 U10435 ( .A1(n8914), .A2(n9251), .ZN(n8909) );
  NAND2_X1 U10436 ( .A1(n8911), .A2(n8910), .ZN(n8913) );
  NAND2_X1 U10437 ( .A1(n8906), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8912) );
  OAI211_X1 U10438 ( .C1(n9251), .C2(n8919), .A(n9240), .B(n9071), .ZN(n8924)
         );
  NAND2_X1 U10439 ( .A1(n8915), .A2(n8914), .ZN(n8921) );
  NAND2_X1 U10440 ( .A1(n5201), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8918) );
  NAND2_X1 U10441 ( .A1(n6554), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8917) );
  NAND2_X1 U10442 ( .A1(n5200), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8916) );
  AND3_X1 U10443 ( .A1(n8918), .A2(n8917), .A3(n8916), .ZN(n8996) );
  INV_X1 U10444 ( .A(n8996), .ZN(n9243) );
  AOI22_X1 U10445 ( .A1(n9251), .A2(n8919), .B1(n9243), .B2(n9071), .ZN(n8920)
         );
  INV_X1 U10446 ( .A(n9058), .ZN(n9010) );
  OAI211_X1 U10447 ( .C1(n8922), .C2(n8921), .A(n8920), .B(n9010), .ZN(n8923)
         );
  AND2_X1 U10448 ( .A1(n9240), .A2(n8996), .ZN(n9057) );
  INV_X1 U10449 ( .A(n9057), .ZN(n9000) );
  OAI211_X1 U10450 ( .C1(n8922), .C2(n8924), .A(n8923), .B(n9000), .ZN(n9012)
         );
  AOI21_X1 U10451 ( .B1(n9012), .B2(n6254), .A(n9023), .ZN(n8960) );
  NOR2_X1 U10452 ( .A1(n9251), .A2(n8925), .ZN(n9056) );
  INV_X1 U10453 ( .A(n9056), .ZN(n8995) );
  AND2_X1 U10454 ( .A1(n9251), .A2(n8925), .ZN(n8992) );
  INV_X1 U10455 ( .A(n8992), .ZN(n8958) );
  INV_X1 U10456 ( .A(n8926), .ZN(n8935) );
  AND2_X1 U10457 ( .A1(n8927), .A2(n9026), .ZN(n8929) );
  AND4_X1 U10458 ( .A1(n8929), .A2(n9750), .A3(n9023), .A4(n8928), .ZN(n8933)
         );
  NAND4_X1 U10459 ( .A1(n8933), .A2(n8932), .A3(n8931), .A4(n8930), .ZN(n8934)
         );
  NOR2_X1 U10460 ( .A1(n8935), .A2(n8934), .ZN(n8936) );
  NAND4_X1 U10461 ( .A1(n9712), .A2(n8938), .A3(n8937), .A4(n8936), .ZN(n8939)
         );
  NOR2_X1 U10462 ( .A1(n8940), .A2(n8939), .ZN(n8942) );
  NAND3_X1 U10463 ( .A1(n8943), .A2(n8942), .A3(n8941), .ZN(n8944) );
  NOR2_X1 U10464 ( .A1(n8945), .A2(n8944), .ZN(n8946) );
  NAND4_X1 U10465 ( .A1(n9400), .A2(n9417), .A3(n8947), .A4(n8946), .ZN(n8948)
         );
  OR4_X1 U10466 ( .A1(n9375), .A2(n9357), .A3(n9387), .A4(n8948), .ZN(n8949)
         );
  NOR3_X1 U10467 ( .A1(n8950), .A2(n9342), .A3(n8949), .ZN(n8951) );
  NAND2_X1 U10468 ( .A1(n8951), .A2(n9311), .ZN(n8952) );
  NOR2_X1 U10469 ( .A1(n9301), .A2(n8952), .ZN(n8953) );
  NAND3_X1 U10470 ( .A1(n9267), .A2(n8953), .A3(n9286), .ZN(n8954) );
  NOR2_X1 U10471 ( .A1(n8955), .A2(n8954), .ZN(n8956) );
  AND4_X1 U10472 ( .A1(n8995), .A2(n8958), .A3(n8957), .A4(n8956), .ZN(n8959)
         );
  AND3_X1 U10473 ( .A1(n9010), .A2(n8959), .A3(n9000), .ZN(n9003) );
  NOR4_X1 U10474 ( .A1(n8990), .A2(n8961), .A3(n8984), .A4(n8981), .ZN(n8994)
         );
  INV_X1 U10475 ( .A(n8962), .ZN(n8963) );
  INV_X1 U10476 ( .A(n9053), .ZN(n8970) );
  NAND2_X1 U10477 ( .A1(n8964), .A2(n9312), .ZN(n8965) );
  NAND2_X1 U10478 ( .A1(n9300), .A2(n8965), .ZN(n8966) );
  NAND2_X1 U10479 ( .A1(n8966), .A2(n8974), .ZN(n8967) );
  AND2_X1 U10480 ( .A1(n8968), .A2(n8967), .ZN(n9052) );
  INV_X1 U10481 ( .A(n9052), .ZN(n8969) );
  NOR3_X1 U10482 ( .A1(n8970), .A2(n9376), .A3(n8969), .ZN(n8998) );
  NAND3_X1 U10483 ( .A1(n8974), .A2(n8972), .A3(n8971), .ZN(n8973) );
  AOI21_X1 U10484 ( .B1(n9052), .B2(n8973), .A(n8980), .ZN(n8983) );
  INV_X1 U10485 ( .A(n8974), .ZN(n8979) );
  NAND2_X1 U10486 ( .A1(n8976), .A2(n8975), .ZN(n8977) );
  NOR4_X1 U10487 ( .A1(n8980), .A2(n8979), .A3(n8978), .A4(n8977), .ZN(n8982)
         );
  NOR4_X1 U10488 ( .A1(n8984), .A2(n8983), .A3(n8982), .A4(n8981), .ZN(n8987)
         );
  OAI21_X1 U10489 ( .B1(n8987), .B2(n8986), .A(n8985), .ZN(n8989) );
  OAI21_X1 U10490 ( .B1(n8990), .B2(n8989), .A(n8988), .ZN(n8991) );
  INV_X1 U10491 ( .A(n9054), .ZN(n8997) );
  OAI22_X1 U10492 ( .A1(n8998), .A2(n8997), .B1(n8996), .B2(n8995), .ZN(n8999)
         );
  OAI211_X1 U10493 ( .C1(n9518), .C2(n9243), .A(n8999), .B(n9010), .ZN(n9002)
         );
  NAND3_X1 U10494 ( .A1(n9002), .A2(n9001), .A3(n9000), .ZN(n9005) );
  INV_X1 U10495 ( .A(n9003), .ZN(n9004) );
  NAND2_X1 U10496 ( .A1(n9005), .A2(n9004), .ZN(n9006) );
  NAND2_X1 U10497 ( .A1(n9006), .A2(n4507), .ZN(n9007) );
  INV_X1 U10498 ( .A(n9008), .ZN(n9009) );
  OAI211_X1 U10499 ( .C1(n9010), .C2(n4507), .A(n9009), .B(n6255), .ZN(n9011)
         );
  NOR2_X1 U10500 ( .A1(n4507), .A2(n9064), .ZN(n9062) );
  NOR2_X1 U10501 ( .A1(n9014), .A2(n9013), .ZN(n9042) );
  INV_X1 U10502 ( .A(n9015), .ZN(n9016) );
  AOI21_X1 U10503 ( .B1(n9018), .B2(n9017), .A(n9016), .ZN(n9020) );
  AOI211_X1 U10504 ( .C1(n9021), .C2(n9042), .A(n9020), .B(n9019), .ZN(n9047)
         );
  INV_X1 U10505 ( .A(n9022), .ZN(n9031) );
  AOI21_X1 U10506 ( .B1(n6276), .B2(n5190), .A(n9023), .ZN(n9027) );
  NAND4_X1 U10507 ( .A1(n9027), .A2(n9026), .A3(n9025), .A4(n9024), .ZN(n9030)
         );
  INV_X1 U10508 ( .A(n9028), .ZN(n9029) );
  NOR3_X1 U10509 ( .A1(n9031), .A2(n9030), .A3(n9029), .ZN(n9034) );
  OAI211_X1 U10510 ( .C1(n9035), .C2(n9034), .A(n9033), .B(n9032), .ZN(n9038)
         );
  AOI21_X1 U10511 ( .B1(n9038), .B2(n9037), .A(n9036), .ZN(n9041) );
  NOR3_X1 U10512 ( .A1(n9041), .A2(n9040), .A3(n9039), .ZN(n9043) );
  OAI21_X1 U10513 ( .B1(n9044), .B2(n9043), .A(n9042), .ZN(n9046) );
  AOI21_X1 U10514 ( .B1(n9047), .B2(n9046), .A(n9045), .ZN(n9050) );
  OAI21_X1 U10515 ( .B1(n9050), .B2(n9049), .A(n9048), .ZN(n9051) );
  NAND3_X1 U10516 ( .A1(n9053), .A2(n9052), .A3(n9051), .ZN(n9055) );
  MUX2_X1 U10517 ( .A(n6256), .B(n9062), .S(n9061), .Z(n9063) );
  NAND3_X1 U10518 ( .A1(n9067), .A2(n9066), .A3(n9065), .ZN(n9068) );
  OAI211_X1 U10519 ( .C1(n6254), .C2(n9070), .A(n9068), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9069) );
  MUX2_X1 U10520 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9243), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10521 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9071), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10522 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9072), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10523 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9073), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10524 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9074), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10525 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9075), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10526 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9076), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10527 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9077), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10528 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9078), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10529 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9079), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10530 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9080), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10531 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9081), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10532 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9082), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10533 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9083), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10534 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9084), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10535 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9085), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10536 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9086), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10537 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9087), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10538 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9088), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10539 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9089), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10540 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9090), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10541 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9091), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10542 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9092), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10543 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9093), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10544 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9094), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10545 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9095), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10546 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9096), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10547 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9097), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10548 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9098), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10549 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n6285), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10550 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6276), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10551 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6265), .S(P1_U3973), .Z(
        P1_U3554) );
  OAI211_X1 U10552 ( .C1(n9101), .C2(n9100), .A(n9692), .B(n9099), .ZN(n9109)
         );
  AOI22_X1 U10553 ( .A1(n9670), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9108) );
  OAI211_X1 U10554 ( .C1(n9104), .C2(n9103), .A(n9699), .B(n9102), .ZN(n9107)
         );
  NAND2_X1 U10555 ( .A1(n9673), .A2(n9105), .ZN(n9106) );
  NAND4_X1 U10556 ( .A1(n9109), .A2(n9108), .A3(n9107), .A4(n9106), .ZN(
        P1_U3244) );
  MUX2_X1 U10557 ( .A(n9111), .B(P1_IR_REG_0__SCAN_IN), .S(n9110), .Z(n9112)
         );
  NAND2_X1 U10558 ( .A1(n9112), .A2(n9114), .ZN(n9113) );
  OAI211_X1 U10559 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9114), .A(n9113), .B(
        P1_U3973), .ZN(n9153) );
  INV_X1 U10560 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9116) );
  OAI22_X1 U10561 ( .A1(n9708), .A2(n9116), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9115), .ZN(n9117) );
  AOI21_X1 U10562 ( .B1(n9118), .B2(n9673), .A(n9117), .ZN(n9127) );
  OAI211_X1 U10563 ( .C1(n9121), .C2(n9120), .A(n9692), .B(n9119), .ZN(n9126)
         );
  OAI211_X1 U10564 ( .C1(n9124), .C2(n9123), .A(n9699), .B(n9122), .ZN(n9125)
         );
  NAND4_X1 U10565 ( .A1(n9153), .A2(n9127), .A3(n9126), .A4(n9125), .ZN(
        P1_U3245) );
  NAND2_X1 U10566 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9128) );
  OAI21_X1 U10567 ( .B1(n9708), .B2(n9129), .A(n9128), .ZN(n9130) );
  AOI21_X1 U10568 ( .B1(n9131), .B2(n9673), .A(n9130), .ZN(n9140) );
  OAI211_X1 U10569 ( .C1(n9134), .C2(n9133), .A(n9692), .B(n9132), .ZN(n9139)
         );
  OAI211_X1 U10570 ( .C1(n9137), .C2(n9136), .A(n9699), .B(n9135), .ZN(n9138)
         );
  NAND3_X1 U10571 ( .A1(n9140), .A2(n9139), .A3(n9138), .ZN(P1_U3246) );
  INV_X1 U10572 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9141) );
  OAI22_X1 U10573 ( .A1(n9708), .A2(n9141), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10296), .ZN(n9142) );
  AOI21_X1 U10574 ( .B1(n9143), .B2(n9673), .A(n9142), .ZN(n9152) );
  OAI211_X1 U10575 ( .C1(n9146), .C2(n9145), .A(n9692), .B(n9144), .ZN(n9151)
         );
  OAI211_X1 U10576 ( .C1(n9149), .C2(n9148), .A(n9699), .B(n9147), .ZN(n9150)
         );
  NAND4_X1 U10577 ( .A1(n9153), .A2(n9152), .A3(n9151), .A4(n9150), .ZN(
        P1_U3247) );
  INV_X1 U10578 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10311) );
  OAI21_X1 U10579 ( .B1(n9708), .B2(n10311), .A(n9154), .ZN(n9155) );
  AOI21_X1 U10580 ( .B1(n9156), .B2(n9673), .A(n9155), .ZN(n9165) );
  OAI211_X1 U10581 ( .C1(n9159), .C2(n9158), .A(n9692), .B(n9157), .ZN(n9164)
         );
  OAI211_X1 U10582 ( .C1(n9162), .C2(n9161), .A(n9699), .B(n9160), .ZN(n9163)
         );
  NAND3_X1 U10583 ( .A1(n9165), .A2(n9164), .A3(n9163), .ZN(P1_U3248) );
  OAI21_X1 U10584 ( .B1(n9708), .B2(n9167), .A(n9166), .ZN(n9168) );
  AOI21_X1 U10585 ( .B1(n9169), .B2(n9673), .A(n9168), .ZN(n9178) );
  OAI211_X1 U10586 ( .C1(n9172), .C2(n9171), .A(n9692), .B(n9170), .ZN(n9177)
         );
  OAI211_X1 U10587 ( .C1(n9175), .C2(n9174), .A(n9699), .B(n9173), .ZN(n9176)
         );
  NAND3_X1 U10588 ( .A1(n9178), .A2(n9177), .A3(n9176), .ZN(P1_U3249) );
  OAI211_X1 U10589 ( .C1(n9181), .C2(n9180), .A(n9692), .B(n9179), .ZN(n9191)
         );
  INV_X1 U10590 ( .A(n9182), .ZN(n9183) );
  AOI21_X1 U10591 ( .B1(n9670), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n9183), .ZN(
        n9190) );
  OAI211_X1 U10592 ( .C1(n9186), .C2(n9185), .A(n9699), .B(n9184), .ZN(n9189)
         );
  OR2_X1 U10593 ( .A1(n9704), .A2(n9187), .ZN(n9188) );
  NAND4_X1 U10594 ( .A1(n9191), .A2(n9190), .A3(n9189), .A4(n9188), .ZN(
        P1_U3250) );
  OAI211_X1 U10595 ( .C1(n9194), .C2(n9193), .A(n9692), .B(n9192), .ZN(n9203)
         );
  AOI21_X1 U10596 ( .B1(n9670), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n9195), .ZN(
        n9202) );
  OAI211_X1 U10597 ( .C1(n9198), .C2(n9197), .A(n9699), .B(n9196), .ZN(n9201)
         );
  NAND2_X1 U10598 ( .A1(n9673), .A2(n9199), .ZN(n9200) );
  NAND4_X1 U10599 ( .A1(n9203), .A2(n9202), .A3(n9201), .A4(n9200), .ZN(
        P1_U3251) );
  NAND2_X1 U10600 ( .A1(n9633), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9204) );
  OAI21_X1 U10601 ( .B1(n9633), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9204), .ZN(
        n9626) );
  OAI21_X1 U10602 ( .B1(n9216), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9205), .ZN(
        n9627) );
  NOR2_X1 U10603 ( .A1(n9626), .A2(n9627), .ZN(n9625) );
  AOI21_X1 U10604 ( .B1(n9633), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9625), .ZN(
        n9642) );
  NAND2_X1 U10605 ( .A1(n9645), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9206) );
  OAI21_X1 U10606 ( .B1(n9645), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9206), .ZN(
        n9641) );
  NOR2_X1 U10607 ( .A1(n9642), .A2(n9641), .ZN(n9640) );
  AOI21_X1 U10608 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9645), .A(n9640), .ZN(
        n9207) );
  NOR2_X1 U10609 ( .A1(n9207), .A2(n9218), .ZN(n9208) );
  XNOR2_X1 U10610 ( .A(n9218), .B(n9207), .ZN(n9655) );
  NOR2_X1 U10611 ( .A1(n9654), .A2(n9655), .ZN(n9653) );
  NOR2_X1 U10612 ( .A1(n9208), .A2(n9653), .ZN(n9667) );
  XNOR2_X1 U10613 ( .A(n9674), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9666) );
  OR2_X1 U10614 ( .A1(n9667), .A2(n9666), .ZN(n9663) );
  NAND2_X1 U10615 ( .A1(n9674), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9209) );
  AND2_X1 U10616 ( .A1(n9663), .A2(n9209), .ZN(n9679) );
  INV_X1 U10617 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9210) );
  XNOR2_X1 U10618 ( .A(n9224), .B(n9210), .ZN(n9680) );
  NAND2_X1 U10619 ( .A1(n9679), .A2(n9680), .ZN(n9678) );
  OR2_X1 U10620 ( .A1(n9224), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9211) );
  AND2_X1 U10621 ( .A1(n9678), .A2(n9211), .ZN(n9695) );
  NAND2_X1 U10622 ( .A1(n9227), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9213) );
  OAI21_X1 U10623 ( .B1(n9227), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9213), .ZN(
        n9212) );
  INV_X1 U10624 ( .A(n9212), .ZN(n9694) );
  NAND2_X1 U10625 ( .A1(n9695), .A2(n9694), .ZN(n9693) );
  NAND2_X1 U10626 ( .A1(n9693), .A2(n9213), .ZN(n9214) );
  XNOR2_X1 U10627 ( .A(n9214), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9232) );
  XNOR2_X1 U10628 ( .A(n9633), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9629) );
  OAI21_X1 U10629 ( .B1(n9216), .B2(P1_REG1_REG_12__SCAN_IN), .A(n9215), .ZN(
        n9630) );
  NOR2_X1 U10630 ( .A1(n9629), .A2(n9630), .ZN(n9628) );
  AOI21_X1 U10631 ( .B1(n9633), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9628), .ZN(
        n9639) );
  XNOR2_X1 U10632 ( .A(n9645), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9638) );
  NOR2_X1 U10633 ( .A1(n9639), .A2(n9638), .ZN(n9637) );
  AOI21_X1 U10634 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9645), .A(n9637), .ZN(
        n9217) );
  NOR2_X1 U10635 ( .A1(n9217), .A2(n9218), .ZN(n9219) );
  XNOR2_X1 U10636 ( .A(n9218), .B(n9217), .ZN(n9652) );
  NOR2_X1 U10637 ( .A1(n9651), .A2(n9652), .ZN(n9650) );
  NOR2_X1 U10638 ( .A1(n9219), .A2(n9650), .ZN(n9672) );
  INV_X1 U10639 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9220) );
  XNOR2_X1 U10640 ( .A(n9674), .B(n9220), .ZN(n9671) );
  NAND2_X1 U10641 ( .A1(n9672), .A2(n9671), .ZN(n9222) );
  OR2_X1 U10642 ( .A1(n9674), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9221) );
  NAND2_X1 U10643 ( .A1(n9222), .A2(n9221), .ZN(n9683) );
  INV_X1 U10644 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9223) );
  XNOR2_X1 U10645 ( .A(n9224), .B(n9223), .ZN(n9682) );
  NAND2_X1 U10646 ( .A1(n9683), .A2(n9682), .ZN(n9226) );
  OR2_X1 U10647 ( .A1(n9224), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9225) );
  NAND2_X1 U10648 ( .A1(n9226), .A2(n9225), .ZN(n9697) );
  NAND2_X1 U10649 ( .A1(n9227), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9228) );
  OAI21_X1 U10650 ( .B1(n9227), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9228), .ZN(
        n9696) );
  NAND2_X1 U10651 ( .A1(n9700), .A2(n9228), .ZN(n9229) );
  INV_X1 U10652 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9482) );
  XNOR2_X1 U10653 ( .A(n9229), .B(n9482), .ZN(n9234) );
  INV_X1 U10654 ( .A(n9234), .ZN(n9230) );
  OAI22_X1 U10655 ( .A1(n9232), .A2(n9665), .B1(n9230), .B2(n9649), .ZN(n9236)
         );
  NAND2_X1 U10656 ( .A1(n9232), .A2(n9231), .ZN(n9233) );
  OAI211_X1 U10657 ( .C1(n9649), .C2(n9234), .A(n9233), .B(n9704), .ZN(n9235)
         );
  MUX2_X1 U10658 ( .A(n9236), .B(n9235), .S(n6252), .Z(n9237) );
  INV_X1 U10659 ( .A(n9237), .ZN(n9239) );
  OAI211_X1 U10660 ( .C1(n5069), .C2(n9708), .A(n9239), .B(n9238), .ZN(
        P1_U3262) );
  NAND2_X1 U10661 ( .A1(n9431), .A2(n9731), .ZN(n9246) );
  AND2_X1 U10662 ( .A1(n9243), .A2(n9242), .ZN(n9434) );
  INV_X1 U10663 ( .A(n9434), .ZN(n9244) );
  NOR2_X1 U10664 ( .A1(n9744), .A2(n9244), .ZN(n9253) );
  AOI21_X1 U10665 ( .B1(n9721), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9253), .ZN(
        n9245) );
  OAI211_X1 U10666 ( .C1(n9514), .C2(n9737), .A(n9246), .B(n9245), .ZN(
        P1_U3263) );
  INV_X1 U10667 ( .A(n9247), .ZN(n9250) );
  INV_X1 U10668 ( .A(n9248), .ZN(n9249) );
  NAND2_X1 U10669 ( .A1(n9435), .A2(n9731), .ZN(n9255) );
  AND2_X1 U10670 ( .A1(n9721), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9252) );
  NOR2_X1 U10671 ( .A1(n9253), .A2(n9252), .ZN(n9254) );
  OAI211_X1 U10672 ( .C1(n9518), .C2(n9737), .A(n9255), .B(n9254), .ZN(
        P1_U3264) );
  NAND3_X1 U10673 ( .A1(n9257), .A2(n9256), .A3(n9741), .ZN(n9265) );
  AOI22_X1 U10674 ( .A1(n9721), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9258), .B2(
        n9733), .ZN(n9259) );
  OAI21_X1 U10675 ( .B1(n9260), .B2(n9737), .A(n9259), .ZN(n9261) );
  AOI21_X1 U10676 ( .B1(n9263), .B2(n9262), .A(n9261), .ZN(n9264) );
  OAI211_X1 U10677 ( .C1(n9744), .C2(n9266), .A(n9265), .B(n9264), .ZN(
        P1_U3265) );
  XNOR2_X1 U10678 ( .A(n9268), .B(n9267), .ZN(n9520) );
  AND2_X1 U10679 ( .A1(n4529), .A2(n9269), .ZN(n9271) );
  INV_X1 U10680 ( .A(n9439), .ZN(n9282) );
  AOI22_X1 U10681 ( .A1(n9721), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9272), .B2(
        n9733), .ZN(n9273) );
  OAI21_X1 U10682 ( .B1(n9519), .B2(n9737), .A(n9273), .ZN(n9281) );
  NAND2_X1 U10683 ( .A1(n9275), .A2(n9274), .ZN(n9277) );
  OAI21_X1 U10684 ( .B1(n4541), .B2(n9277), .A(n9276), .ZN(n9279) );
  NOR2_X1 U10685 ( .A1(n9440), .A2(n9721), .ZN(n9280) );
  AOI211_X1 U10686 ( .C1(n9282), .C2(n9731), .A(n9281), .B(n9280), .ZN(n9283)
         );
  OAI21_X1 U10687 ( .B1(n9520), .B2(n9430), .A(n9283), .ZN(P1_U3266) );
  XNOR2_X1 U10688 ( .A(n9285), .B(n9284), .ZN(n9526) );
  AOI22_X1 U10689 ( .A1(n9446), .A2(n9722), .B1(n9721), .B2(
        P1_REG2_REG_26__SCAN_IN), .ZN(n9295) );
  XNOR2_X1 U10690 ( .A(n9287), .B(n9286), .ZN(n9289) );
  OAI21_X1 U10691 ( .B1(n9289), .B2(n9752), .A(n9288), .ZN(n9444) );
  AOI21_X1 U10692 ( .B1(n9297), .B2(n9446), .A(n9422), .ZN(n9290) );
  NAND2_X1 U10693 ( .A1(n9290), .A2(n4529), .ZN(n9443) );
  INV_X1 U10694 ( .A(n9291), .ZN(n9292) );
  OAI22_X1 U10695 ( .A1(n9443), .A2(n6252), .B1(n9405), .B2(n9292), .ZN(n9293)
         );
  OAI21_X1 U10696 ( .B1(n9444), .B2(n9293), .A(n9409), .ZN(n9294) );
  OAI211_X1 U10697 ( .C1(n9526), .C2(n9430), .A(n9295), .B(n9294), .ZN(
        P1_U3267) );
  OAI211_X1 U10698 ( .C1(n9527), .C2(n9321), .A(n9724), .B(n9297), .ZN(n9449)
         );
  INV_X1 U10699 ( .A(n9449), .ZN(n9308) );
  AOI22_X1 U10700 ( .A1(n9721), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9298), .B2(
        n9733), .ZN(n9299) );
  OAI21_X1 U10701 ( .B1(n9527), .B2(n9737), .A(n9299), .ZN(n9307) );
  NAND2_X1 U10702 ( .A1(n9315), .A2(n9300), .ZN(n9302) );
  XNOR2_X1 U10703 ( .A(n9302), .B(n9301), .ZN(n9305) );
  INV_X1 U10704 ( .A(n9303), .ZN(n9304) );
  AOI21_X1 U10705 ( .B1(n9305), .B2(n9710), .A(n9304), .ZN(n9450) );
  NOR2_X1 U10706 ( .A1(n9450), .A2(n9721), .ZN(n9306) );
  AOI211_X1 U10707 ( .C1(n9308), .C2(n9731), .A(n9307), .B(n9306), .ZN(n9309)
         );
  OAI21_X1 U10708 ( .B1(n9528), .B2(n9430), .A(n9309), .ZN(P1_U3268) );
  XOR2_X1 U10709 ( .A(n9310), .B(n9311), .Z(n9534) );
  INV_X1 U10710 ( .A(n9311), .ZN(n9314) );
  NAND2_X1 U10711 ( .A1(n9329), .A2(n9312), .ZN(n9313) );
  NAND2_X1 U10712 ( .A1(n9314), .A2(n9313), .ZN(n9316) );
  NAND3_X1 U10713 ( .A1(n9316), .A2(n9710), .A3(n9315), .ZN(n9318) );
  NAND2_X1 U10714 ( .A1(n9318), .A2(n9317), .ZN(n9456) );
  NAND2_X1 U10715 ( .A1(n9323), .A2(n9334), .ZN(n9319) );
  NAND2_X1 U10716 ( .A1(n9319), .A2(n9724), .ZN(n9320) );
  OR2_X1 U10717 ( .A1(n9321), .A2(n9320), .ZN(n9453) );
  AOI22_X1 U10718 ( .A1(n9721), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9322), .B2(
        n9733), .ZN(n9325) );
  NAND2_X1 U10719 ( .A1(n9323), .A2(n9722), .ZN(n9324) );
  OAI211_X1 U10720 ( .C1(n9453), .C2(n9370), .A(n9325), .B(n9324), .ZN(n9326)
         );
  AOI21_X1 U10721 ( .B1(n9456), .B2(n9409), .A(n9326), .ZN(n9327) );
  OAI21_X1 U10722 ( .B1(n9534), .B2(n9430), .A(n9327), .ZN(P1_U3269) );
  XNOR2_X1 U10723 ( .A(n9328), .B(n9331), .ZN(n9538) );
  AOI22_X1 U10724 ( .A1(n9459), .A2(n9722), .B1(n9721), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n9340) );
  OAI21_X1 U10725 ( .B1(n9331), .B2(n9330), .A(n9329), .ZN(n9332) );
  AND2_X1 U10726 ( .A1(n9332), .A2(n9710), .ZN(n9463) );
  NAND2_X1 U10727 ( .A1(n9347), .A2(n9459), .ZN(n9333) );
  NAND3_X1 U10728 ( .A1(n9334), .A2(n9724), .A3(n9333), .ZN(n9461) );
  INV_X1 U10729 ( .A(n9335), .ZN(n9336) );
  AOI21_X1 U10730 ( .B1(n9336), .B2(n9733), .A(n9458), .ZN(n9337) );
  OAI21_X1 U10731 ( .B1(n9461), .B2(n6252), .A(n9337), .ZN(n9338) );
  OAI21_X1 U10732 ( .B1(n9463), .B2(n9338), .A(n9409), .ZN(n9339) );
  OAI211_X1 U10733 ( .C1(n9538), .C2(n9430), .A(n9340), .B(n9339), .ZN(
        P1_U3270) );
  XNOR2_X1 U10734 ( .A(n9341), .B(n9342), .ZN(n9542) );
  XNOR2_X1 U10735 ( .A(n9343), .B(n9342), .ZN(n9345) );
  OAI21_X1 U10736 ( .B1(n9345), .B2(n9752), .A(n9344), .ZN(n9466) );
  INV_X1 U10737 ( .A(n9346), .ZN(n9364) );
  INV_X1 U10738 ( .A(n9347), .ZN(n9348) );
  AOI211_X1 U10739 ( .C1(n9467), .C2(n9364), .A(n9422), .B(n9348), .ZN(n9465)
         );
  NAND2_X1 U10740 ( .A1(n9465), .A2(n9731), .ZN(n9352) );
  INV_X1 U10741 ( .A(n9349), .ZN(n9350) );
  AOI22_X1 U10742 ( .A1(n9350), .A2(n9733), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9721), .ZN(n9351) );
  OAI211_X1 U10743 ( .C1(n9353), .C2(n9737), .A(n9352), .B(n9351), .ZN(n9354)
         );
  AOI21_X1 U10744 ( .B1(n9409), .B2(n9466), .A(n9354), .ZN(n9355) );
  OAI21_X1 U10745 ( .B1(n9542), .B2(n9430), .A(n9355), .ZN(P1_U3271) );
  XNOR2_X1 U10746 ( .A(n9356), .B(n9357), .ZN(n9545) );
  NAND2_X1 U10747 ( .A1(n9358), .A2(n9357), .ZN(n9359) );
  NAND2_X1 U10748 ( .A1(n9360), .A2(n9359), .ZN(n9362) );
  AOI21_X1 U10749 ( .B1(n9362), .B2(n9710), .A(n9361), .ZN(n9471) );
  INV_X1 U10750 ( .A(n9471), .ZN(n9372) );
  INV_X1 U10751 ( .A(n9363), .ZN(n9380) );
  OAI211_X1 U10752 ( .C1(n9544), .C2(n9380), .A(n9364), .B(n9724), .ZN(n9470)
         );
  INV_X1 U10753 ( .A(n9365), .ZN(n9366) );
  AOI22_X1 U10754 ( .A1(n9721), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9366), .B2(
        n9733), .ZN(n9369) );
  NAND2_X1 U10755 ( .A1(n9367), .A2(n9722), .ZN(n9368) );
  OAI211_X1 U10756 ( .C1(n9470), .C2(n9370), .A(n9369), .B(n9368), .ZN(n9371)
         );
  AOI21_X1 U10757 ( .B1(n9372), .B2(n9409), .A(n9371), .ZN(n9373) );
  OAI21_X1 U10758 ( .B1(n9545), .B2(n9430), .A(n9373), .ZN(P1_U3272) );
  XNOR2_X1 U10759 ( .A(n9374), .B(n9375), .ZN(n9552) );
  XNOR2_X1 U10760 ( .A(n9376), .B(n9375), .ZN(n9377) );
  NAND2_X1 U10761 ( .A1(n9377), .A2(n9710), .ZN(n9379) );
  NAND2_X1 U10762 ( .A1(n9379), .A2(n9378), .ZN(n9474) );
  AOI211_X1 U10763 ( .C1(n9476), .C2(n9391), .A(n9422), .B(n9380), .ZN(n9475)
         );
  NAND2_X1 U10764 ( .A1(n9475), .A2(n9731), .ZN(n9383) );
  AOI22_X1 U10765 ( .A1(n9721), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9381), .B2(
        n9733), .ZN(n9382) );
  OAI211_X1 U10766 ( .C1(n4773), .C2(n9737), .A(n9383), .B(n9382), .ZN(n9384)
         );
  AOI21_X1 U10767 ( .B1(n9409), .B2(n9474), .A(n9384), .ZN(n9385) );
  OAI21_X1 U10768 ( .B1(n9552), .B2(n9430), .A(n9385), .ZN(P1_U3273) );
  XNOR2_X1 U10769 ( .A(n9386), .B(n9387), .ZN(n9556) );
  XNOR2_X1 U10770 ( .A(n9388), .B(n9387), .ZN(n9390) );
  OAI21_X1 U10771 ( .B1(n9390), .B2(n9752), .A(n9389), .ZN(n9479) );
  AOI211_X1 U10772 ( .C1(n9481), .C2(n9399), .A(n9422), .B(n4774), .ZN(n9480)
         );
  NAND2_X1 U10773 ( .A1(n9480), .A2(n9731), .ZN(n9394) );
  AOI22_X1 U10774 ( .A1(n9721), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9392), .B2(
        n9733), .ZN(n9393) );
  OAI211_X1 U10775 ( .C1(n9395), .C2(n9737), .A(n9394), .B(n9393), .ZN(n9396)
         );
  AOI21_X1 U10776 ( .B1(n9409), .B2(n9479), .A(n9396), .ZN(n9397) );
  OAI21_X1 U10777 ( .B1(n9556), .B2(n9430), .A(n9397), .ZN(P1_U3274) );
  XOR2_X1 U10778 ( .A(n9398), .B(n9400), .Z(n9485) );
  INV_X1 U10779 ( .A(n9485), .ZN(n9412) );
  OAI211_X1 U10780 ( .C1(n9404), .C2(n9421), .A(n9724), .B(n9399), .ZN(n9488)
         );
  XNOR2_X1 U10781 ( .A(n9401), .B(n9400), .ZN(n9402) );
  NAND2_X1 U10782 ( .A1(n9402), .A2(n9710), .ZN(n9489) );
  INV_X1 U10783 ( .A(n9486), .ZN(n9403) );
  OAI211_X1 U10784 ( .C1(n6252), .C2(n9488), .A(n9489), .B(n9403), .ZN(n9410)
         );
  NOR2_X1 U10785 ( .A1(n9404), .A2(n9737), .ZN(n9408) );
  INV_X1 U10786 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10421) );
  OAI22_X1 U10787 ( .A1(n9409), .A2(n10421), .B1(n9406), .B2(n9405), .ZN(n9407) );
  AOI211_X1 U10788 ( .C1(n9410), .C2(n9409), .A(n9408), .B(n9407), .ZN(n9411)
         );
  OAI21_X1 U10789 ( .B1(n9412), .B2(n9430), .A(n9411), .ZN(P1_U3275) );
  XNOR2_X1 U10790 ( .A(n9413), .B(n9414), .ZN(n9496) );
  INV_X1 U10791 ( .A(n9415), .ZN(n9418) );
  OAI211_X1 U10792 ( .C1(n9418), .C2(n9417), .A(n9710), .B(n9416), .ZN(n9420)
         );
  NAND2_X1 U10793 ( .A1(n9420), .A2(n9419), .ZN(n9493) );
  AOI211_X1 U10794 ( .C1(n9494), .C2(n9423), .A(n9422), .B(n9421), .ZN(n9492)
         );
  NAND2_X1 U10795 ( .A1(n9492), .A2(n9731), .ZN(n9426) );
  AOI22_X1 U10796 ( .A1(n9744), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9424), .B2(
        n9733), .ZN(n9425) );
  OAI211_X1 U10797 ( .C1(n9427), .C2(n9737), .A(n9426), .B(n9425), .ZN(n9428)
         );
  AOI21_X1 U10798 ( .B1(n9409), .B2(n9493), .A(n9428), .ZN(n9429) );
  OAI21_X1 U10799 ( .B1(n9496), .B2(n9430), .A(n9429), .ZN(P1_U3276) );
  INV_X1 U10800 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9432) );
  NOR2_X1 U10801 ( .A1(n9431), .A2(n9434), .ZN(n9511) );
  MUX2_X1 U10802 ( .A(n9432), .B(n9511), .S(n9797), .Z(n9433) );
  OAI21_X1 U10803 ( .B1(n9514), .B2(n9469), .A(n9433), .ZN(P1_U3553) );
  INV_X1 U10804 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9436) );
  NOR2_X1 U10805 ( .A1(n9435), .A2(n9434), .ZN(n9515) );
  MUX2_X1 U10806 ( .A(n9436), .B(n9515), .S(n9797), .Z(n9437) );
  OAI21_X1 U10807 ( .B1(n9518), .B2(n9469), .A(n9437), .ZN(P1_U3552) );
  MUX2_X1 U10808 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9438), .S(n9797), .Z(
        P1_U3550) );
  OAI22_X1 U10809 ( .A1(n9520), .A2(n9484), .B1(n9519), .B2(n9469), .ZN(n9442)
         );
  NAND2_X1 U10810 ( .A1(n9440), .A2(n9439), .ZN(n9521) );
  MUX2_X1 U10811 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9521), .S(n9797), .Z(n9441) );
  OR2_X1 U10812 ( .A1(n9442), .A2(n9441), .ZN(P1_U3549) );
  INV_X1 U10813 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9447) );
  INV_X1 U10814 ( .A(n9443), .ZN(n9445) );
  AOI211_X1 U10815 ( .C1(n9499), .C2(n9446), .A(n9445), .B(n9444), .ZN(n9524)
         );
  MUX2_X1 U10816 ( .A(n9447), .B(n9524), .S(n9797), .Z(n9448) );
  OAI21_X1 U10817 ( .B1(n9526), .B2(n9484), .A(n9448), .ZN(P1_U3548) );
  OAI22_X1 U10818 ( .A1(n9528), .A2(n9484), .B1(n9527), .B2(n9469), .ZN(n9452)
         );
  NAND2_X1 U10819 ( .A1(n9450), .A2(n9449), .ZN(n9529) );
  MUX2_X1 U10820 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9529), .S(n9797), .Z(n9451) );
  OR2_X1 U10821 ( .A1(n9452), .A2(n9451), .ZN(P1_U3547) );
  INV_X1 U10822 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10433) );
  OAI21_X1 U10823 ( .B1(n9454), .B2(n9779), .A(n9453), .ZN(n9455) );
  NOR2_X1 U10824 ( .A1(n9456), .A2(n9455), .ZN(n9532) );
  MUX2_X1 U10825 ( .A(n10433), .B(n9532), .S(n9797), .Z(n9457) );
  OAI21_X1 U10826 ( .B1(n9534), .B2(n9484), .A(n9457), .ZN(P1_U3546) );
  AOI21_X1 U10827 ( .B1(n9459), .B2(n9499), .A(n9458), .ZN(n9460) );
  NAND2_X1 U10828 ( .A1(n9461), .A2(n9460), .ZN(n9462) );
  NOR2_X1 U10829 ( .A1(n9463), .A2(n9462), .ZN(n9535) );
  MUX2_X1 U10830 ( .A(n10409), .B(n9535), .S(n9797), .Z(n9464) );
  OAI21_X1 U10831 ( .B1(n9538), .B2(n9484), .A(n9464), .ZN(P1_U3545) );
  AOI211_X1 U10832 ( .C1(n9499), .C2(n9467), .A(n9466), .B(n9465), .ZN(n9539)
         );
  MUX2_X1 U10833 ( .A(n10394), .B(n9539), .S(n9797), .Z(n9468) );
  OAI21_X1 U10834 ( .B1(n9542), .B2(n9484), .A(n9468), .ZN(P1_U3544) );
  OAI22_X1 U10835 ( .A1(n9545), .A2(n9484), .B1(n9544), .B2(n9469), .ZN(n9473)
         );
  NAND2_X1 U10836 ( .A1(n9471), .A2(n9470), .ZN(n9546) );
  MUX2_X1 U10837 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9546), .S(n9797), .Z(n9472) );
  OR2_X1 U10838 ( .A1(n9473), .A2(n9472), .ZN(P1_U3543) );
  INV_X1 U10839 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9477) );
  AOI211_X1 U10840 ( .C1(n9499), .C2(n9476), .A(n9475), .B(n9474), .ZN(n9549)
         );
  MUX2_X1 U10841 ( .A(n9477), .B(n9549), .S(n9797), .Z(n9478) );
  OAI21_X1 U10842 ( .B1(n9552), .B2(n9484), .A(n9478), .ZN(P1_U3542) );
  AOI211_X1 U10843 ( .C1(n9499), .C2(n9481), .A(n9480), .B(n9479), .ZN(n9553)
         );
  MUX2_X1 U10844 ( .A(n9482), .B(n9553), .S(n9797), .Z(n9483) );
  OAI21_X1 U10845 ( .B1(n9556), .B2(n9484), .A(n9483), .ZN(P1_U3541) );
  NAND2_X1 U10846 ( .A1(n9485), .A2(n9768), .ZN(n9491) );
  AOI21_X1 U10847 ( .B1(n9487), .B2(n9499), .A(n9486), .ZN(n9490) );
  NAND4_X1 U10848 ( .A1(n9491), .A2(n9490), .A3(n9489), .A4(n9488), .ZN(n9557)
         );
  MUX2_X1 U10849 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9557), .S(n9797), .Z(
        P1_U3540) );
  AOI211_X1 U10850 ( .C1(n9499), .C2(n9494), .A(n9493), .B(n9492), .ZN(n9495)
         );
  OAI21_X1 U10851 ( .B1(n9496), .B2(n9751), .A(n9495), .ZN(n9558) );
  MUX2_X1 U10852 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9558), .S(n9797), .Z(
        P1_U3539) );
  NAND3_X1 U10853 ( .A1(n9498), .A2(n9497), .A3(n9768), .ZN(n9504) );
  NAND2_X1 U10854 ( .A1(n9500), .A2(n9499), .ZN(n9501) );
  NAND4_X1 U10855 ( .A1(n9504), .A2(n9503), .A3(n9502), .A4(n9501), .ZN(n9559)
         );
  MUX2_X1 U10856 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9559), .S(n9797), .Z(
        P1_U3538) );
  OAI21_X1 U10857 ( .B1(n9506), .B2(n9779), .A(n9505), .ZN(n9508) );
  AOI211_X1 U10858 ( .C1(n9785), .C2(n9509), .A(n9508), .B(n9507), .ZN(n9561)
         );
  NAND2_X1 U10859 ( .A1(n9795), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9510) );
  OAI21_X1 U10860 ( .B1(n9561), .B2(n9795), .A(n9510), .ZN(P1_U3536) );
  INV_X1 U10861 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9512) );
  MUX2_X1 U10862 ( .A(n9512), .B(n9511), .S(n9788), .Z(n9513) );
  OAI21_X1 U10863 ( .B1(n9514), .B2(n9543), .A(n9513), .ZN(P1_U3521) );
  INV_X1 U10864 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9516) );
  MUX2_X1 U10865 ( .A(n9516), .B(n9515), .S(n9788), .Z(n9517) );
  OAI21_X1 U10866 ( .B1(n9518), .B2(n9543), .A(n9517), .ZN(P1_U3520) );
  OAI22_X1 U10867 ( .A1(n9520), .A2(n9555), .B1(n9519), .B2(n9543), .ZN(n9523)
         );
  MUX2_X1 U10868 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9521), .S(n9788), .Z(n9522) );
  OR2_X1 U10869 ( .A1(n9523), .A2(n9522), .ZN(P1_U3517) );
  INV_X1 U10870 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10248) );
  MUX2_X1 U10871 ( .A(n10248), .B(n9524), .S(n9788), .Z(n9525) );
  OAI21_X1 U10872 ( .B1(n9526), .B2(n9555), .A(n9525), .ZN(P1_U3516) );
  OAI22_X1 U10873 ( .A1(n9528), .A2(n9555), .B1(n9527), .B2(n9543), .ZN(n9531)
         );
  MUX2_X1 U10874 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9529), .S(n9788), .Z(n9530) );
  OR2_X1 U10875 ( .A1(n9531), .A2(n9530), .ZN(P1_U3515) );
  INV_X1 U10876 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10391) );
  MUX2_X1 U10877 ( .A(n10391), .B(n9532), .S(n9788), .Z(n9533) );
  OAI21_X1 U10878 ( .B1(n9534), .B2(n9555), .A(n9533), .ZN(P1_U3514) );
  INV_X1 U10879 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9536) );
  MUX2_X1 U10880 ( .A(n9536), .B(n9535), .S(n9788), .Z(n9537) );
  OAI21_X1 U10881 ( .B1(n9538), .B2(n9555), .A(n9537), .ZN(P1_U3513) );
  INV_X1 U10882 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9540) );
  MUX2_X1 U10883 ( .A(n9540), .B(n9539), .S(n9788), .Z(n9541) );
  OAI21_X1 U10884 ( .B1(n9542), .B2(n9555), .A(n9541), .ZN(P1_U3512) );
  OAI22_X1 U10885 ( .A1(n9545), .A2(n9555), .B1(n9544), .B2(n9543), .ZN(n9548)
         );
  MUX2_X1 U10886 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9546), .S(n9788), .Z(n9547) );
  OR2_X1 U10887 ( .A1(n9548), .A2(n9547), .ZN(P1_U3511) );
  INV_X1 U10888 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9550) );
  MUX2_X1 U10889 ( .A(n9550), .B(n9549), .S(n9788), .Z(n9551) );
  OAI21_X1 U10890 ( .B1(n9552), .B2(n9555), .A(n9551), .ZN(P1_U3510) );
  MUX2_X1 U10891 ( .A(n10372), .B(n9553), .S(n9788), .Z(n9554) );
  OAI21_X1 U10892 ( .B1(n9556), .B2(n9555), .A(n9554), .ZN(P1_U3509) );
  MUX2_X1 U10893 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9557), .S(n9788), .Z(
        P1_U3507) );
  MUX2_X1 U10894 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9558), .S(n9788), .Z(
        P1_U3504) );
  MUX2_X1 U10895 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9559), .S(n9788), .Z(
        P1_U3501) );
  NAND2_X1 U10896 ( .A1(n9786), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9560) );
  OAI21_X1 U10897 ( .B1(n9561), .B2(n9786), .A(n9560), .ZN(P1_U3495) );
  NOR4_X1 U10898 ( .A1(n5155), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n5322), .ZN(n9562) );
  AOI21_X1 U10899 ( .B1(n9563), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9562), .ZN(
        n9564) );
  OAI21_X1 U10900 ( .B1(n9565), .B2(n9572), .A(n9564), .ZN(P1_U3324) );
  INV_X1 U10901 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9566) );
  OAI222_X1 U10902 ( .A1(n9572), .A2(n9568), .B1(n9567), .B2(P1_U3086), .C1(
        n9566), .C2(n9569), .ZN(P1_U3326) );
  OAI222_X1 U10903 ( .A1(n9572), .A2(n9571), .B1(P1_U3086), .B2(n5675), .C1(
        n9570), .C2(n9569), .ZN(P1_U3327) );
  MUX2_X1 U10904 ( .A(n9573), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NAND2_X1 U10905 ( .A1(n9575), .A2(n9574), .ZN(n9576) );
  NAND3_X1 U10906 ( .A1(n9692), .A2(n9577), .A3(n9576), .ZN(n9583) );
  NAND2_X1 U10907 ( .A1(n9579), .A2(n9578), .ZN(n9580) );
  NAND3_X1 U10908 ( .A1(n9581), .A2(n9699), .A3(n9580), .ZN(n9582) );
  OAI211_X1 U10909 ( .C1(n9704), .C2(n9584), .A(n9583), .B(n9582), .ZN(n9585)
         );
  INV_X1 U10910 ( .A(n9585), .ZN(n9587) );
  NAND2_X1 U10911 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9586) );
  OAI211_X1 U10912 ( .C1(n9588), .C2(n9708), .A(n9587), .B(n9586), .ZN(
        P1_U3253) );
  XNOR2_X1 U10913 ( .A(n9590), .B(n9589), .ZN(n9604) );
  AND2_X1 U10914 ( .A1(n9591), .A2(n10090), .ZN(n9603) );
  NAND2_X1 U10915 ( .A1(n9603), .A2(n9592), .ZN(n9593) );
  OAI21_X1 U10916 ( .B1(n9594), .B2(n10022), .A(n9593), .ZN(n9600) );
  XNOR2_X1 U10917 ( .A(n9596), .B(n9595), .ZN(n9597) );
  OAI222_X1 U10918 ( .A1(n10031), .A2(n9599), .B1(n10032), .B2(n9598), .C1(
        n9597), .C2(n10041), .ZN(n9602) );
  AOI211_X1 U10919 ( .C1(n9604), .C2(n10034), .A(n9600), .B(n9602), .ZN(n9601)
         );
  AOI22_X1 U10920 ( .A1(n10038), .A2(n5925), .B1(n9601), .B2(n10035), .ZN(
        P2_U3220) );
  AOI211_X1 U10921 ( .C1(n9604), .C2(n10082), .A(n9603), .B(n9602), .ZN(n9605)
         );
  AOI22_X1 U10922 ( .A1(n10105), .A2(n9605), .B1(n5930), .B2(n10103), .ZN(
        P2_U3472) );
  INV_X1 U10923 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9606) );
  AOI22_X1 U10924 ( .A1(n10093), .A2(n9606), .B1(n9605), .B2(n10091), .ZN(
        P2_U3429) );
  INV_X1 U10925 ( .A(P1_WR_REG_SCAN_IN), .ZN(n10346) );
  XOR2_X1 U10926 ( .A(n10346), .B(P2_WR_REG_SCAN_IN), .Z(U123) );
  INV_X1 U10927 ( .A(P2_RD_REG_SCAN_IN), .ZN(n10485) );
  XOR2_X1 U10928 ( .A(n10485), .B(P1_RD_REG_SCAN_IN), .Z(U126) );
  INV_X1 U10929 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9624) );
  INV_X1 U10930 ( .A(n9607), .ZN(n9620) );
  NAND2_X1 U10931 ( .A1(n9609), .A2(n9608), .ZN(n9612) );
  NOR2_X1 U10932 ( .A1(n9665), .A2(n9610), .ZN(n9611) );
  NAND2_X1 U10933 ( .A1(n9612), .A2(n9611), .ZN(n9619) );
  NAND2_X1 U10934 ( .A1(n9614), .A2(n9613), .ZN(n9617) );
  NOR2_X1 U10935 ( .A1(n9649), .A2(n9615), .ZN(n9616) );
  NAND2_X1 U10936 ( .A1(n9617), .A2(n9616), .ZN(n9618) );
  OAI211_X1 U10937 ( .C1(n9704), .C2(n9620), .A(n9619), .B(n9618), .ZN(n9621)
         );
  INV_X1 U10938 ( .A(n9621), .ZN(n9623) );
  OAI211_X1 U10939 ( .C1(n9624), .C2(n9708), .A(n9623), .B(n9622), .ZN(
        P1_U3254) );
  INV_X1 U10940 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9636) );
  AOI211_X1 U10941 ( .C1(n9627), .C2(n9626), .A(n9625), .B(n9665), .ZN(n9632)
         );
  AOI211_X1 U10942 ( .C1(n9630), .C2(n9629), .A(n9628), .B(n9649), .ZN(n9631)
         );
  AOI211_X1 U10943 ( .C1(n9673), .C2(n9633), .A(n9632), .B(n9631), .ZN(n9635)
         );
  OAI211_X1 U10944 ( .C1(n9636), .C2(n9708), .A(n9635), .B(n9634), .ZN(
        P1_U3256) );
  INV_X1 U10945 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9648) );
  AOI211_X1 U10946 ( .C1(n9639), .C2(n9638), .A(n9637), .B(n9649), .ZN(n9644)
         );
  AOI211_X1 U10947 ( .C1(n9642), .C2(n9641), .A(n9640), .B(n9665), .ZN(n9643)
         );
  AOI211_X1 U10948 ( .C1(n9673), .C2(n9645), .A(n9644), .B(n9643), .ZN(n9647)
         );
  NAND2_X1 U10949 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9646) );
  OAI211_X1 U10950 ( .C1(n9648), .C2(n9708), .A(n9647), .B(n9646), .ZN(
        P1_U3257) );
  INV_X1 U10951 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9662) );
  AOI211_X1 U10952 ( .C1(n9652), .C2(n9651), .A(n9650), .B(n9649), .ZN(n9657)
         );
  AOI211_X1 U10953 ( .C1(n9655), .C2(n9654), .A(n9653), .B(n9665), .ZN(n9656)
         );
  AOI211_X1 U10954 ( .C1(n9673), .C2(n9658), .A(n9657), .B(n9656), .ZN(n9661)
         );
  NAND2_X1 U10955 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n9660) );
  OAI211_X1 U10956 ( .C1(n9662), .C2(n9708), .A(n9661), .B(n9660), .ZN(
        P1_U3258) );
  INV_X1 U10957 ( .A(n9663), .ZN(n9664) );
  AOI211_X1 U10958 ( .C1(n9667), .C2(n9666), .A(n9665), .B(n9664), .ZN(n9668)
         );
  AOI211_X1 U10959 ( .C1(P1_ADDR_REG_16__SCAN_IN), .C2(n9670), .A(n9669), .B(
        n9668), .ZN(n9677) );
  XNOR2_X1 U10960 ( .A(n9672), .B(n9671), .ZN(n9675) );
  AOI22_X1 U10961 ( .A1(n9675), .A2(n9699), .B1(n9674), .B2(n9673), .ZN(n9676)
         );
  NAND2_X1 U10962 ( .A1(n9677), .A2(n9676), .ZN(P1_U3259) );
  INV_X1 U10963 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9691) );
  OAI21_X1 U10964 ( .B1(n9680), .B2(n9679), .A(n9678), .ZN(n9681) );
  NAND2_X1 U10965 ( .A1(n9681), .A2(n9692), .ZN(n9686) );
  XNOR2_X1 U10966 ( .A(n9683), .B(n9682), .ZN(n9684) );
  NAND2_X1 U10967 ( .A1(n9684), .A2(n9699), .ZN(n9685) );
  OAI211_X1 U10968 ( .C1(n9704), .C2(n9687), .A(n9686), .B(n9685), .ZN(n9688)
         );
  INV_X1 U10969 ( .A(n9688), .ZN(n9690) );
  OAI211_X1 U10970 ( .C1(n9691), .C2(n9708), .A(n9690), .B(n9689), .ZN(
        P1_U3260) );
  OAI211_X1 U10971 ( .C1(n9695), .C2(n9694), .A(n9693), .B(n9692), .ZN(n9702)
         );
  NAND2_X1 U10972 ( .A1(n9697), .A2(n9696), .ZN(n9698) );
  NAND3_X1 U10973 ( .A1(n9700), .A2(n9699), .A3(n9698), .ZN(n9701) );
  OAI211_X1 U10974 ( .C1(n9704), .C2(n9703), .A(n9702), .B(n9701), .ZN(n9705)
         );
  INV_X1 U10975 ( .A(n9705), .ZN(n9707) );
  NAND2_X1 U10976 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9706) );
  OAI211_X1 U10977 ( .C1(n10419), .C2(n9708), .A(n9707), .B(n9706), .ZN(
        P1_U3261) );
  XNOR2_X1 U10978 ( .A(n9709), .B(n9712), .ZN(n9784) );
  NAND2_X1 U10979 ( .A1(n9711), .A2(n9710), .ZN(n9717) );
  AOI21_X1 U10980 ( .B1(n9714), .B2(n9713), .A(n9712), .ZN(n9716) );
  OAI21_X1 U10981 ( .B1(n9717), .B2(n9716), .A(n9715), .ZN(n9718) );
  AOI21_X1 U10982 ( .B1(n9784), .B2(n9719), .A(n9718), .ZN(n9781) );
  AOI222_X1 U10983 ( .A1(n9723), .A2(n9722), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n9721), .C1(n9733), .C2(n9720), .ZN(n9730) );
  INV_X1 U10984 ( .A(n9723), .ZN(n9780) );
  OAI211_X1 U10985 ( .C1(n9780), .C2(n9726), .A(n9725), .B(n9724), .ZN(n9778)
         );
  INV_X1 U10986 ( .A(n9778), .ZN(n9727) );
  AOI22_X1 U10987 ( .A1(n9784), .A2(n9728), .B1(n9731), .B2(n9727), .ZN(n9729)
         );
  OAI211_X1 U10988 ( .C1(n9744), .C2(n9781), .A(n9730), .B(n9729), .ZN(
        P1_U3282) );
  NAND2_X1 U10989 ( .A1(n9732), .A2(n9731), .ZN(n9736) );
  AOI22_X1 U10990 ( .A1(n9744), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n9734), .B2(
        n9733), .ZN(n9735) );
  OAI211_X1 U10991 ( .C1(n9738), .C2(n9737), .A(n9736), .B(n9735), .ZN(n9739)
         );
  AOI21_X1 U10992 ( .B1(n9741), .B2(n9740), .A(n9739), .ZN(n9742) );
  OAI21_X1 U10993 ( .B1(n9744), .B2(n9743), .A(n9742), .ZN(P1_U3289) );
  AND2_X1 U10994 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9746), .ZN(P1_U3294) );
  AND2_X1 U10995 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9746), .ZN(P1_U3295) );
  AND2_X1 U10996 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9746), .ZN(P1_U3296) );
  AND2_X1 U10997 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9746), .ZN(P1_U3297) );
  AND2_X1 U10998 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9746), .ZN(P1_U3298) );
  INV_X1 U10999 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10320) );
  NOR2_X1 U11000 ( .A1(n9745), .A2(n10320), .ZN(P1_U3299) );
  AND2_X1 U11001 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9746), .ZN(P1_U3300) );
  AND2_X1 U11002 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9746), .ZN(P1_U3301) );
  INV_X1 U11003 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10392) );
  NOR2_X1 U11004 ( .A1(n9745), .A2(n10392), .ZN(P1_U3302) );
  AND2_X1 U11005 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9746), .ZN(P1_U3303) );
  AND2_X1 U11006 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9746), .ZN(P1_U3304) );
  AND2_X1 U11007 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9746), .ZN(P1_U3305) );
  AND2_X1 U11008 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9746), .ZN(P1_U3306) );
  AND2_X1 U11009 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9746), .ZN(P1_U3307) );
  AND2_X1 U11010 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9746), .ZN(P1_U3308) );
  AND2_X1 U11011 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9746), .ZN(P1_U3309) );
  AND2_X1 U11012 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9746), .ZN(P1_U3310) );
  AND2_X1 U11013 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9746), .ZN(P1_U3311) );
  AND2_X1 U11014 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9746), .ZN(P1_U3312) );
  AND2_X1 U11015 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9746), .ZN(P1_U3313) );
  INV_X1 U11016 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10422) );
  NOR2_X1 U11017 ( .A1(n9745), .A2(n10422), .ZN(P1_U3314) );
  INV_X1 U11018 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10438) );
  NOR2_X1 U11019 ( .A1(n9745), .A2(n10438), .ZN(P1_U3315) );
  AND2_X1 U11020 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9746), .ZN(P1_U3316) );
  AND2_X1 U11021 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9746), .ZN(P1_U3317) );
  AND2_X1 U11022 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9746), .ZN(P1_U3318) );
  AND2_X1 U11023 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9746), .ZN(P1_U3319) );
  AND2_X1 U11024 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9746), .ZN(P1_U3320) );
  AND2_X1 U11025 ( .A1(n9746), .A2(P1_D_REG_4__SCAN_IN), .ZN(P1_U3321) );
  INV_X1 U11026 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10355) );
  NOR2_X1 U11027 ( .A1(n9745), .A2(n10355), .ZN(P1_U3322) );
  AND2_X1 U11028 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9746), .ZN(P1_U3323) );
  OAI21_X1 U11029 ( .B1(n9749), .B2(n9748), .A(n9747), .ZN(P1_U3439) );
  AOI21_X1 U11030 ( .B1(n9752), .B2(n9751), .A(n9750), .ZN(n9753) );
  AOI211_X1 U11031 ( .C1(n9756), .C2(n9755), .A(n9754), .B(n9753), .ZN(n9789)
         );
  INV_X1 U11032 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9757) );
  AOI22_X1 U11033 ( .A1(n9788), .A2(n9789), .B1(n9757), .B2(n9786), .ZN(
        P1_U3453) );
  INV_X1 U11034 ( .A(n9758), .ZN(n9759) );
  OAI21_X1 U11035 ( .B1(n5190), .B2(n9779), .A(n9759), .ZN(n9762) );
  INV_X1 U11036 ( .A(n9760), .ZN(n9761) );
  AOI211_X1 U11037 ( .C1(n9768), .C2(n9763), .A(n9762), .B(n9761), .ZN(n9790)
         );
  INV_X1 U11038 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10340) );
  AOI22_X1 U11039 ( .A1(n9788), .A2(n9790), .B1(n10340), .B2(n9786), .ZN(
        P1_U3456) );
  OAI211_X1 U11040 ( .C1(n9766), .C2(n9779), .A(n9765), .B(n9764), .ZN(n9767)
         );
  AOI21_X1 U11041 ( .B1(n9769), .B2(n9768), .A(n9767), .ZN(n9792) );
  INV_X1 U11042 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9770) );
  AOI22_X1 U11043 ( .A1(n9788), .A2(n9792), .B1(n9770), .B2(n9786), .ZN(
        P1_U3459) );
  OAI21_X1 U11044 ( .B1(n9772), .B2(n9779), .A(n9771), .ZN(n9773) );
  AOI21_X1 U11045 ( .B1(n9774), .B2(n9785), .A(n9773), .ZN(n9775) );
  AND2_X1 U11046 ( .A1(n9776), .A2(n9775), .ZN(n9794) );
  INV_X1 U11047 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9777) );
  AOI22_X1 U11048 ( .A1(n9788), .A2(n9794), .B1(n9777), .B2(n9786), .ZN(
        P1_U3474) );
  OAI21_X1 U11049 ( .B1(n9780), .B2(n9779), .A(n9778), .ZN(n9783) );
  INV_X1 U11050 ( .A(n9781), .ZN(n9782) );
  AOI211_X1 U11051 ( .C1(n9785), .C2(n9784), .A(n9783), .B(n9782), .ZN(n9796)
         );
  INV_X1 U11052 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9787) );
  AOI22_X1 U11053 ( .A1(n9788), .A2(n9796), .B1(n9787), .B2(n9786), .ZN(
        P1_U3486) );
  AOI22_X1 U11054 ( .A1(n9797), .A2(n9789), .B1(n6264), .B2(n9795), .ZN(
        P1_U3522) );
  AOI22_X1 U11055 ( .A1(n9797), .A2(n9790), .B1(n6687), .B2(n9795), .ZN(
        P1_U3523) );
  AOI22_X1 U11056 ( .A1(n9797), .A2(n9792), .B1(n9791), .B2(n9795), .ZN(
        P1_U3524) );
  AOI22_X1 U11057 ( .A1(n9797), .A2(n9794), .B1(n9793), .B2(n9795), .ZN(
        P1_U3529) );
  AOI22_X1 U11058 ( .A1(n9797), .A2(n9796), .B1(n6725), .B2(n9795), .ZN(
        P1_U3533) );
  OR2_X1 U11059 ( .A1(n10157), .A2(n9798), .ZN(n9808) );
  OAI21_X1 U11060 ( .B1(n9800), .B2(P2_REG1_REG_3__SCAN_IN), .A(n9799), .ZN(
        n9801) );
  NAND2_X1 U11061 ( .A1(n10153), .A2(n9801), .ZN(n9807) );
  INV_X1 U11062 ( .A(n9802), .ZN(n9806) );
  AOI21_X1 U11063 ( .B1(n9803), .B2(n7120), .A(n9815), .ZN(n9804) );
  OR2_X1 U11064 ( .A1(n10147), .A2(n9804), .ZN(n9805) );
  AND4_X1 U11065 ( .A1(n9808), .A2(n9807), .A3(n9806), .A4(n9805), .ZN(n9814)
         );
  OAI21_X1 U11066 ( .B1(n9811), .B2(n9810), .A(n9809), .ZN(n9812) );
  AOI22_X1 U11067 ( .A1(n9812), .A2(n10010), .B1(n10159), .B2(
        P2_ADDR_REG_3__SCAN_IN), .ZN(n9813) );
  NAND2_X1 U11068 ( .A1(n9814), .A2(n9813), .ZN(P2_U3185) );
  NOR2_X1 U11069 ( .A1(n9816), .A2(n9815), .ZN(n9817) );
  NAND2_X1 U11070 ( .A1(n9818), .A2(n9817), .ZN(n9819) );
  NAND2_X1 U11071 ( .A1(n9820), .A2(n9819), .ZN(n9822) );
  AOI21_X1 U11072 ( .B1(n9980), .B2(n9822), .A(n9821), .ZN(n9835) );
  INV_X1 U11073 ( .A(n9823), .ZN(n9824) );
  XNOR2_X1 U11074 ( .A(n9825), .B(n9824), .ZN(n9826) );
  NAND2_X1 U11075 ( .A1(n9826), .A2(n10010), .ZN(n9834) );
  OR2_X1 U11076 ( .A1(n10157), .A2(n9827), .ZN(n9833) );
  OAI21_X1 U11077 ( .B1(n9830), .B2(n9829), .A(n9828), .ZN(n9831) );
  NAND2_X1 U11078 ( .A1(n10153), .A2(n9831), .ZN(n9832) );
  AND4_X1 U11079 ( .A1(n9835), .A2(n9834), .A3(n9833), .A4(n9832), .ZN(n9836)
         );
  OAI21_X1 U11080 ( .B1(n9837), .B2(n10307), .A(n9836), .ZN(P2_U3186) );
  OAI21_X1 U11081 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(n9839), .A(n9838), .ZN(
        n9847) );
  AOI21_X1 U11082 ( .B1(n9841), .B2(n5848), .A(n9840), .ZN(n9845) );
  AOI21_X1 U11083 ( .B1(n10002), .B2(n9843), .A(n9842), .ZN(n9844) );
  OAI21_X1 U11084 ( .B1(n9845), .B2(n10147), .A(n9844), .ZN(n9846) );
  AOI21_X1 U11085 ( .B1(n9847), .B2(n10153), .A(n9846), .ZN(n9853) );
  OAI21_X1 U11086 ( .B1(n9850), .B2(n9849), .A(n9848), .ZN(n9851) );
  AOI22_X1 U11087 ( .A1(n9851), .A2(n10010), .B1(n10159), .B2(
        P2_ADDR_REG_7__SCAN_IN), .ZN(n9852) );
  NAND2_X1 U11088 ( .A1(n9853), .A2(n9852), .ZN(P2_U3189) );
  AOI21_X1 U11089 ( .B1(n10002), .B2(n9855), .A(n9854), .ZN(n9871) );
  OAI21_X1 U11090 ( .B1(n9858), .B2(n9857), .A(n9856), .ZN(n9859) );
  AOI22_X1 U11091 ( .A1(n10159), .A2(P2_ADDR_REG_8__SCAN_IN), .B1(n10010), 
        .B2(n9859), .ZN(n9870) );
  AOI21_X1 U11092 ( .B1(n9862), .B2(n9861), .A(n9860), .ZN(n9863) );
  OR2_X1 U11093 ( .A1(n9863), .A2(n10147), .ZN(n9869) );
  OAI21_X1 U11094 ( .B1(n9866), .B2(n9865), .A(n9864), .ZN(n9867) );
  NAND2_X1 U11095 ( .A1(n9867), .A2(n10153), .ZN(n9868) );
  NAND4_X1 U11096 ( .A1(n9871), .A2(n9870), .A3(n9869), .A4(n9868), .ZN(
        P2_U3190) );
  AOI22_X1 U11097 ( .A1(n9872), .A2(n10002), .B1(n10159), .B2(
        P2_ADDR_REG_9__SCAN_IN), .ZN(n9887) );
  OAI21_X1 U11098 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n9874), .A(n9873), .ZN(
        n9879) );
  OAI21_X1 U11099 ( .B1(n9877), .B2(n9876), .A(n9875), .ZN(n9878) );
  AOI22_X1 U11100 ( .A1(n9879), .A2(n10153), .B1(n10010), .B2(n9878), .ZN(
        n9886) );
  AOI21_X1 U11101 ( .B1(n9882), .B2(n9881), .A(n9880), .ZN(n9883) );
  OR2_X1 U11102 ( .A1(n10147), .A2(n9883), .ZN(n9884) );
  NAND4_X1 U11103 ( .A1(n9887), .A2(n9886), .A3(n9885), .A4(n9884), .ZN(
        P2_U3191) );
  AOI22_X1 U11104 ( .A1(n9888), .A2(n10002), .B1(n10159), .B2(
        P2_ADDR_REG_10__SCAN_IN), .ZN(n9903) );
  OAI21_X1 U11105 ( .B1(n9891), .B2(n9890), .A(n9889), .ZN(n9896) );
  OAI21_X1 U11106 ( .B1(n9894), .B2(n9893), .A(n9892), .ZN(n9895) );
  AOI22_X1 U11107 ( .A1(n9896), .A2(n10153), .B1(n10010), .B2(n9895), .ZN(
        n9902) );
  AOI21_X1 U11108 ( .B1(n4590), .B2(n9898), .A(n9897), .ZN(n9899) );
  OR2_X1 U11109 ( .A1(n9899), .A2(n10147), .ZN(n9900) );
  NAND4_X1 U11110 ( .A1(n9903), .A2(n9902), .A3(n9901), .A4(n9900), .ZN(
        P2_U3192) );
  AOI22_X1 U11111 ( .A1(n9904), .A2(n10002), .B1(n10159), .B2(
        P2_ADDR_REG_11__SCAN_IN), .ZN(n9918) );
  OAI21_X1 U11112 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n9906), .A(n9905), .ZN(
        n9911) );
  OAI21_X1 U11113 ( .B1(n9909), .B2(n9908), .A(n9907), .ZN(n9910) );
  AOI22_X1 U11114 ( .A1(n9911), .A2(n10153), .B1(n10010), .B2(n9910), .ZN(
        n9917) );
  AOI21_X1 U11115 ( .B1(n9913), .B2(n5897), .A(n9912), .ZN(n9914) );
  OR2_X1 U11116 ( .A1(n10147), .A2(n9914), .ZN(n9915) );
  NAND4_X1 U11117 ( .A1(n9918), .A2(n9917), .A3(n9916), .A4(n9915), .ZN(
        P2_U3193) );
  AOI22_X1 U11118 ( .A1(n9919), .A2(n10002), .B1(n10159), .B2(
        P2_ADDR_REG_12__SCAN_IN), .ZN(n9935) );
  OAI21_X1 U11119 ( .B1(n9922), .B2(n9921), .A(n9920), .ZN(n9927) );
  OAI21_X1 U11120 ( .B1(n9925), .B2(n9924), .A(n9923), .ZN(n9926) );
  AOI22_X1 U11121 ( .A1(n9927), .A2(n10153), .B1(n10010), .B2(n9926), .ZN(
        n9934) );
  AOI21_X1 U11122 ( .B1(n9930), .B2(n9929), .A(n9928), .ZN(n9931) );
  OR2_X1 U11123 ( .A1(n9931), .A2(n10147), .ZN(n9932) );
  NAND4_X1 U11124 ( .A1(n9935), .A2(n9934), .A3(n9933), .A4(n9932), .ZN(
        P2_U3194) );
  AOI22_X1 U11125 ( .A1(n9936), .A2(n10002), .B1(n10159), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n9951) );
  OAI21_X1 U11126 ( .B1(n9938), .B2(P2_REG1_REG_13__SCAN_IN), .A(n9937), .ZN(
        n9943) );
  OAI21_X1 U11127 ( .B1(n9941), .B2(n9940), .A(n9939), .ZN(n9942) );
  AOI22_X1 U11128 ( .A1(n9943), .A2(n10153), .B1(n10010), .B2(n9942), .ZN(
        n9950) );
  INV_X1 U11129 ( .A(n9944), .ZN(n9945) );
  NOR2_X1 U11130 ( .A1(n9945), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9946) );
  OAI21_X1 U11131 ( .B1(n9947), .B2(n9946), .A(n9980), .ZN(n9948) );
  NAND4_X1 U11132 ( .A1(n9951), .A2(n9950), .A3(n9949), .A4(n9948), .ZN(
        P2_U3195) );
  AOI22_X1 U11133 ( .A1(n9952), .A2(n10002), .B1(n10159), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n9968) );
  OAI21_X1 U11134 ( .B1(n9955), .B2(n9954), .A(n9953), .ZN(n9960) );
  OAI21_X1 U11135 ( .B1(n9958), .B2(n9957), .A(n9956), .ZN(n9959) );
  AOI22_X1 U11136 ( .A1(n9960), .A2(n10153), .B1(n10010), .B2(n9959), .ZN(
        n9967) );
  NAND2_X1 U11137 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n9966) );
  AOI21_X1 U11138 ( .B1(n9963), .B2(n9962), .A(n9961), .ZN(n9964) );
  OR2_X1 U11139 ( .A1(n10147), .A2(n9964), .ZN(n9965) );
  NAND4_X1 U11140 ( .A1(n9968), .A2(n9967), .A3(n9966), .A4(n9965), .ZN(
        P2_U3196) );
  AOI22_X1 U11141 ( .A1(n9969), .A2(n10002), .B1(n10159), .B2(
        P2_ADDR_REG_15__SCAN_IN), .ZN(n9984) );
  OAI21_X1 U11142 ( .B1(n9971), .B2(P2_REG1_REG_15__SCAN_IN), .A(n9970), .ZN(
        n9976) );
  OAI21_X1 U11143 ( .B1(n9974), .B2(n9973), .A(n9972), .ZN(n9975) );
  AOI22_X1 U11144 ( .A1(n9976), .A2(n10153), .B1(n10010), .B2(n9975), .ZN(
        n9983) );
  OAI21_X1 U11145 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n9978), .A(n9977), .ZN(
        n9979) );
  NAND2_X1 U11146 ( .A1(n9980), .A2(n9979), .ZN(n9981) );
  NAND4_X1 U11147 ( .A1(n9984), .A2(n9983), .A3(n9982), .A4(n9981), .ZN(
        P2_U3197) );
  AOI22_X1 U11148 ( .A1(n9985), .A2(n10002), .B1(n10159), .B2(
        P2_ADDR_REG_16__SCAN_IN), .ZN(n10001) );
  OAI21_X1 U11149 ( .B1(n9988), .B2(n9987), .A(n9986), .ZN(n9993) );
  OAI21_X1 U11150 ( .B1(n9991), .B2(n9990), .A(n9989), .ZN(n9992) );
  AOI22_X1 U11151 ( .A1(n9993), .A2(n10153), .B1(n10010), .B2(n9992), .ZN(
        n10000) );
  NAND2_X1 U11152 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3151), .ZN(n9999) );
  AOI21_X1 U11153 ( .B1(n9996), .B2(n9995), .A(n9994), .ZN(n9997) );
  OR2_X1 U11154 ( .A1(n10147), .A2(n9997), .ZN(n9998) );
  NAND4_X1 U11155 ( .A1(n10001), .A2(n10000), .A3(n9999), .A4(n9998), .ZN(
        P2_U3198) );
  AOI22_X1 U11156 ( .A1(n10003), .A2(n10002), .B1(n10159), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n10018) );
  OAI21_X1 U11157 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n10005), .A(n10004), 
        .ZN(n10011) );
  OAI21_X1 U11158 ( .B1(n10008), .B2(n10007), .A(n10006), .ZN(n10009) );
  AOI22_X1 U11159 ( .A1(n10011), .A2(n10153), .B1(n10010), .B2(n10009), .ZN(
        n10017) );
  NAND2_X1 U11160 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3151), .ZN(n10016)
         );
  NAND4_X1 U11161 ( .A1(n10018), .A2(n10017), .A3(n10016), .A4(n10015), .ZN(
        P2_U3199) );
  OAI21_X1 U11162 ( .B1(n10020), .B2(n10025), .A(n10019), .ZN(n10053) );
  OAI22_X1 U11163 ( .A1(n10050), .A2(n10023), .B1(n10022), .B2(n10021), .ZN(
        n10033) );
  NAND3_X1 U11164 ( .A1(n10026), .A2(n10025), .A3(n10024), .ZN(n10027) );
  AND2_X1 U11165 ( .A1(n10028), .A2(n10027), .ZN(n10029) );
  OAI222_X1 U11166 ( .A1(n10032), .A2(n4735), .B1(n10031), .B2(n10030), .C1(
        n10041), .C2(n10029), .ZN(n10051) );
  AOI211_X1 U11167 ( .C1(n10034), .C2(n10053), .A(n10033), .B(n10051), .ZN(
        n10036) );
  AOI22_X1 U11168 ( .A1(n10038), .A2(n10037), .B1(n10036), .B2(n10035), .ZN(
        P2_U3231) );
  INV_X1 U11169 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10045) );
  INV_X1 U11170 ( .A(n10039), .ZN(n10040) );
  AOI21_X1 U11171 ( .B1(n10041), .B2(n10084), .A(n10040), .ZN(n10042) );
  AOI211_X1 U11172 ( .C1(n10044), .C2(n10090), .A(n10043), .B(n10042), .ZN(
        n10094) );
  AOI22_X1 U11173 ( .A1(n10093), .A2(n10045), .B1(n10094), .B2(n10091), .ZN(
        P2_U3390) );
  INV_X1 U11174 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10363) );
  OAI21_X1 U11175 ( .B1(n10077), .B2(n10047), .A(n10046), .ZN(n10048) );
  AOI21_X1 U11176 ( .B1(n10082), .B2(n10049), .A(n10048), .ZN(n10096) );
  AOI22_X1 U11177 ( .A1(n10093), .A2(n10363), .B1(n10096), .B2(n10091), .ZN(
        P2_U3393) );
  NOR2_X1 U11178 ( .A1(n10050), .A2(n10077), .ZN(n10052) );
  AOI211_X1 U11179 ( .C1(n10082), .C2(n10053), .A(n10052), .B(n10051), .ZN(
        n10097) );
  AOI22_X1 U11180 ( .A1(n10093), .A2(n5781), .B1(n10097), .B2(n10091), .ZN(
        P2_U3396) );
  INV_X1 U11181 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10059) );
  INV_X1 U11182 ( .A(n10054), .ZN(n10058) );
  OAI22_X1 U11183 ( .A1(n10056), .A2(n10084), .B1(n10055), .B2(n10077), .ZN(
        n10057) );
  NOR2_X1 U11184 ( .A1(n10058), .A2(n10057), .ZN(n10098) );
  AOI22_X1 U11185 ( .A1(n10093), .A2(n10059), .B1(n10098), .B2(n10091), .ZN(
        P2_U3399) );
  INV_X1 U11186 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10065) );
  INV_X1 U11187 ( .A(n10060), .ZN(n10064) );
  OAI21_X1 U11188 ( .B1(n10062), .B2(n10077), .A(n10061), .ZN(n10063) );
  AOI21_X1 U11189 ( .B1(n10064), .B2(n10082), .A(n10063), .ZN(n10099) );
  AOI22_X1 U11190 ( .A1(n10093), .A2(n10065), .B1(n10099), .B2(n10091), .ZN(
        P2_U3408) );
  INV_X1 U11191 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10407) );
  OAI22_X1 U11192 ( .A1(n10068), .A2(n10067), .B1(n10066), .B2(n10077), .ZN(
        n10069) );
  NOR2_X1 U11193 ( .A1(n10070), .A2(n10069), .ZN(n10100) );
  AOI22_X1 U11194 ( .A1(n10093), .A2(n10407), .B1(n10100), .B2(n10091), .ZN(
        P2_U3411) );
  INV_X1 U11195 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10076) );
  INV_X1 U11196 ( .A(n10071), .ZN(n10075) );
  OAI22_X1 U11197 ( .A1(n10073), .A2(n10084), .B1(n10072), .B2(n10077), .ZN(
        n10074) );
  NOR2_X1 U11198 ( .A1(n10075), .A2(n10074), .ZN(n10101) );
  AOI22_X1 U11199 ( .A1(n10093), .A2(n10076), .B1(n10101), .B2(n10091), .ZN(
        P2_U3414) );
  INV_X1 U11200 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10083) );
  NOR2_X1 U11201 ( .A1(n10078), .A2(n10077), .ZN(n10080) );
  AOI211_X1 U11202 ( .C1(n10082), .C2(n10081), .A(n10080), .B(n10079), .ZN(
        n10102) );
  AOI22_X1 U11203 ( .A1(n10093), .A2(n10083), .B1(n10102), .B2(n10091), .ZN(
        P2_U3423) );
  INV_X1 U11204 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10092) );
  NOR2_X1 U11205 ( .A1(n10085), .A2(n10084), .ZN(n10088) );
  INV_X1 U11206 ( .A(n10086), .ZN(n10087) );
  AOI211_X1 U11207 ( .C1(n10090), .C2(n10089), .A(n10088), .B(n10087), .ZN(
        n10104) );
  AOI22_X1 U11208 ( .A1(n10093), .A2(n10092), .B1(n10104), .B2(n10091), .ZN(
        P2_U3426) );
  AOI22_X1 U11209 ( .A1(n10105), .A2(n10094), .B1(n5771), .B2(n10103), .ZN(
        P2_U3459) );
  INV_X1 U11210 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10095) );
  AOI22_X1 U11211 ( .A1(n10105), .A2(n10096), .B1(n10095), .B2(n10103), .ZN(
        P2_U3460) );
  AOI22_X1 U11212 ( .A1(n10105), .A2(n10097), .B1(n6843), .B2(n10103), .ZN(
        P2_U3461) );
  AOI22_X1 U11213 ( .A1(n10105), .A2(n10098), .B1(n6986), .B2(n10103), .ZN(
        P2_U3462) );
  AOI22_X1 U11214 ( .A1(n10105), .A2(n10099), .B1(n8308), .B2(n10103), .ZN(
        P2_U3465) );
  AOI22_X1 U11215 ( .A1(n10105), .A2(n10100), .B1(n5844), .B2(n10103), .ZN(
        P2_U3466) );
  AOI22_X1 U11216 ( .A1(n10105), .A2(n10101), .B1(n5834), .B2(n10103), .ZN(
        P2_U3467) );
  AOI22_X1 U11217 ( .A1(n10105), .A2(n10102), .B1(n5900), .B2(n10103), .ZN(
        P2_U3470) );
  AOI22_X1 U11218 ( .A1(n10105), .A2(n10104), .B1(n5916), .B2(n10103), .ZN(
        P2_U3471) );
  INV_X1 U11219 ( .A(n10106), .ZN(n10107) );
  NAND2_X1 U11220 ( .A1(n10108), .A2(n10107), .ZN(n10109) );
  XOR2_X1 U11221 ( .A(n10284), .B(n10109), .Z(ADD_1068_U5) );
  INV_X1 U11222 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10364) );
  INV_X1 U11223 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10110) );
  AOI22_X1 U11224 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n10364), .B2(n10110), .ZN(ADD_1068_U46) );
  AOI21_X1 U11225 ( .B1(n10419), .B2(n10112), .A(n10111), .ZN(n10113) );
  XOR2_X1 U11226 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10113), .Z(ADD_1068_U55)
         );
  OAI21_X1 U11227 ( .B1(n10116), .B2(n10115), .A(n10114), .ZN(ADD_1068_U56) );
  OAI21_X1 U11228 ( .B1(n10119), .B2(n10118), .A(n10117), .ZN(ADD_1068_U57) );
  OAI21_X1 U11229 ( .B1(n10122), .B2(n10121), .A(n10120), .ZN(ADD_1068_U58) );
  OAI21_X1 U11230 ( .B1(n10125), .B2(n10124), .A(n10123), .ZN(ADD_1068_U59) );
  OAI21_X1 U11231 ( .B1(n10128), .B2(n10127), .A(n10126), .ZN(ADD_1068_U60) );
  OAI21_X1 U11232 ( .B1(n10131), .B2(n10130), .A(n10129), .ZN(ADD_1068_U61) );
  AOI21_X1 U11233 ( .B1(n10134), .B2(n10133), .A(n10132), .ZN(ADD_1068_U62) );
  NAND2_X1 U11234 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10135) );
  NAND2_X1 U11235 ( .A1(n10136), .A2(n10135), .ZN(n10138) );
  XNOR2_X1 U11236 ( .A(n10138), .B(n10137), .ZN(ADD_1068_U63) );
  AOI211_X1 U11237 ( .C1(n10142), .C2(n10141), .A(n10140), .B(n10139), .ZN(
        n10143) );
  INV_X1 U11238 ( .A(n10143), .ZN(n10155) );
  OAI21_X1 U11239 ( .B1(n10145), .B2(P2_REG1_REG_5__SCAN_IN), .A(n10144), .ZN(
        n10152) );
  NAND2_X1 U11240 ( .A1(n10146), .A2(n6985), .ZN(n10148) );
  AOI21_X1 U11241 ( .B1(n10149), .B2(n10148), .A(n10147), .ZN(n10150) );
  AOI211_X1 U11242 ( .C1(n10153), .C2(n10152), .A(n10151), .B(n10150), .ZN(
        n10154) );
  OAI211_X1 U11243 ( .C1(n10157), .C2(n10156), .A(n10155), .B(n10154), .ZN(
        n10158) );
  AOI21_X1 U11244 ( .B1(n10159), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n10158), .ZN(
        n10546) );
  AOI22_X1 U11245 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(keyinput222), .B1(
        P2_IR_REG_26__SCAN_IN), .B2(keyinput207), .ZN(n10160) );
  OAI221_X1 U11246 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(keyinput222), .C1(
        P2_IR_REG_26__SCAN_IN), .C2(keyinput207), .A(n10160), .ZN(n10167) );
  AOI22_X1 U11247 ( .A1(P1_REG0_REG_24__SCAN_IN), .A2(keyinput166), .B1(
        P2_D_REG_21__SCAN_IN), .B2(keyinput223), .ZN(n10161) );
  OAI221_X1 U11248 ( .B1(P1_REG0_REG_24__SCAN_IN), .B2(keyinput166), .C1(
        P2_D_REG_21__SCAN_IN), .C2(keyinput223), .A(n10161), .ZN(n10166) );
  AOI22_X1 U11249 ( .A1(P1_REG0_REG_19__SCAN_IN), .A2(keyinput145), .B1(
        P2_D_REG_20__SCAN_IN), .B2(keyinput211), .ZN(n10162) );
  OAI221_X1 U11250 ( .B1(P1_REG0_REG_19__SCAN_IN), .B2(keyinput145), .C1(
        P2_D_REG_20__SCAN_IN), .C2(keyinput211), .A(n10162), .ZN(n10165) );
  AOI22_X1 U11251 ( .A1(P1_REG1_REG_13__SCAN_IN), .A2(keyinput172), .B1(
        P2_D_REG_30__SCAN_IN), .B2(keyinput205), .ZN(n10163) );
  OAI221_X1 U11252 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(keyinput172), .C1(
        P2_D_REG_30__SCAN_IN), .C2(keyinput205), .A(n10163), .ZN(n10164) );
  NOR4_X1 U11253 ( .A1(n10167), .A2(n10166), .A3(n10165), .A4(n10164), .ZN(
        n10195) );
  AOI22_X1 U11254 ( .A1(P1_REG0_REG_4__SCAN_IN), .A2(keyinput254), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(keyinput231), .ZN(n10168) );
  OAI221_X1 U11255 ( .B1(P1_REG0_REG_4__SCAN_IN), .B2(keyinput254), .C1(
        P2_DATAO_REG_24__SCAN_IN), .C2(keyinput231), .A(n10168), .ZN(n10175)
         );
  AOI22_X1 U11256 ( .A1(P1_REG1_REG_26__SCAN_IN), .A2(keyinput201), .B1(
        P2_IR_REG_9__SCAN_IN), .B2(keyinput180), .ZN(n10169) );
  OAI221_X1 U11257 ( .B1(P1_REG1_REG_26__SCAN_IN), .B2(keyinput201), .C1(
        P2_IR_REG_9__SCAN_IN), .C2(keyinput180), .A(n10169), .ZN(n10174) );
  AOI22_X1 U11258 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput225), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(keyinput226), .ZN(n10170) );
  OAI221_X1 U11259 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput225), .C1(
        P1_DATAO_REG_21__SCAN_IN), .C2(keyinput226), .A(n10170), .ZN(n10173)
         );
  AOI22_X1 U11260 ( .A1(P2_REG2_REG_5__SCAN_IN), .A2(keyinput218), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(keyinput255), .ZN(n10171) );
  OAI221_X1 U11261 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(keyinput218), .C1(
        P1_DATAO_REG_11__SCAN_IN), .C2(keyinput255), .A(n10171), .ZN(n10172)
         );
  NOR4_X1 U11262 ( .A1(n10175), .A2(n10174), .A3(n10173), .A4(n10172), .ZN(
        n10194) );
  AOI22_X1 U11263 ( .A1(P1_REG0_REG_15__SCAN_IN), .A2(keyinput139), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(keyinput193), .ZN(n10176) );
  OAI221_X1 U11264 ( .B1(P1_REG0_REG_15__SCAN_IN), .B2(keyinput139), .C1(
        P2_DATAO_REG_13__SCAN_IN), .C2(keyinput193), .A(n10176), .ZN(n10183)
         );
  AOI22_X1 U11265 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(keyinput246), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(keyinput169), .ZN(n10177) );
  OAI221_X1 U11266 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(keyinput246), .C1(
        P1_DATAO_REG_19__SCAN_IN), .C2(keyinput169), .A(n10177), .ZN(n10182)
         );
  AOI22_X1 U11267 ( .A1(P2_REG0_REG_19__SCAN_IN), .A2(keyinput204), .B1(
        P2_D_REG_26__SCAN_IN), .B2(keyinput138), .ZN(n10178) );
  OAI221_X1 U11268 ( .B1(P2_REG0_REG_19__SCAN_IN), .B2(keyinput204), .C1(
        P2_D_REG_26__SCAN_IN), .C2(keyinput138), .A(n10178), .ZN(n10181) );
  AOI22_X1 U11269 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(keyinput136), .B1(
        P2_IR_REG_22__SCAN_IN), .B2(keyinput141), .ZN(n10179) );
  OAI221_X1 U11270 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(keyinput136), .C1(
        P2_IR_REG_22__SCAN_IN), .C2(keyinput141), .A(n10179), .ZN(n10180) );
  NOR4_X1 U11271 ( .A1(n10183), .A2(n10182), .A3(n10181), .A4(n10180), .ZN(
        n10193) );
  AOI22_X1 U11272 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(keyinput212), .B1(
        P2_REG0_REG_18__SCAN_IN), .B2(keyinput196), .ZN(n10184) );
  OAI221_X1 U11273 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(keyinput212), .C1(
        P2_REG0_REG_18__SCAN_IN), .C2(keyinput196), .A(n10184), .ZN(n10191) );
  AOI22_X1 U11274 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput243), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput173), .ZN(n10185) );
  OAI221_X1 U11275 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput243), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput173), .A(n10185), .ZN(n10190) );
  AOI22_X1 U11276 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(keyinput182), .B1(
        P1_REG2_REG_26__SCAN_IN), .B2(keyinput185), .ZN(n10186) );
  OAI221_X1 U11277 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(keyinput182), .C1(
        P1_REG2_REG_26__SCAN_IN), .C2(keyinput185), .A(n10186), .ZN(n10189) );
  AOI22_X1 U11278 ( .A1(P1_REG1_REG_17__SCAN_IN), .A2(keyinput210), .B1(
        P2_REG1_REG_4__SCAN_IN), .B2(keyinput249), .ZN(n10187) );
  OAI221_X1 U11279 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(keyinput210), .C1(
        P2_REG1_REG_4__SCAN_IN), .C2(keyinput249), .A(n10187), .ZN(n10188) );
  NOR4_X1 U11280 ( .A1(n10191), .A2(n10190), .A3(n10189), .A4(n10188), .ZN(
        n10192) );
  NAND4_X1 U11281 ( .A1(n10195), .A2(n10194), .A3(n10193), .A4(n10192), .ZN(
        n10338) );
  AOI22_X1 U11282 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(keyinput213), .B1(
        P2_REG0_REG_2__SCAN_IN), .B2(keyinput168), .ZN(n10196) );
  OAI221_X1 U11283 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(keyinput213), .C1(
        P2_REG0_REG_2__SCAN_IN), .C2(keyinput168), .A(n10196), .ZN(n10203) );
  AOI22_X1 U11284 ( .A1(P1_WR_REG_SCAN_IN), .A2(keyinput203), .B1(
        P2_REG3_REG_25__SCAN_IN), .B2(keyinput132), .ZN(n10197) );
  OAI221_X1 U11285 ( .B1(P1_WR_REG_SCAN_IN), .B2(keyinput203), .C1(
        P2_REG3_REG_25__SCAN_IN), .C2(keyinput132), .A(n10197), .ZN(n10202) );
  AOI22_X1 U11286 ( .A1(P1_REG0_REG_14__SCAN_IN), .A2(keyinput235), .B1(
        P1_REG1_REG_24__SCAN_IN), .B2(keyinput189), .ZN(n10198) );
  OAI221_X1 U11287 ( .B1(P1_REG0_REG_14__SCAN_IN), .B2(keyinput235), .C1(
        P1_REG1_REG_24__SCAN_IN), .C2(keyinput189), .A(n10198), .ZN(n10201) );
  AOI22_X1 U11288 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput194), .B1(
        P2_REG3_REG_23__SCAN_IN), .B2(keyinput238), .ZN(n10199) );
  OAI221_X1 U11289 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput194), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput238), .A(n10199), .ZN(n10200) );
  NOR4_X1 U11290 ( .A1(n10203), .A2(n10202), .A3(n10201), .A4(n10200), .ZN(
        n10231) );
  AOI22_X1 U11291 ( .A1(P2_REG2_REG_3__SCAN_IN), .A2(keyinput167), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput140), .ZN(n10204) );
  OAI221_X1 U11292 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(keyinput167), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput140), .A(n10204), .ZN(n10211) );
  AOI22_X1 U11293 ( .A1(P1_REG1_REG_21__SCAN_IN), .A2(keyinput134), .B1(
        P2_REG0_REG_21__SCAN_IN), .B2(keyinput142), .ZN(n10205) );
  OAI221_X1 U11294 ( .B1(P1_REG1_REG_21__SCAN_IN), .B2(keyinput134), .C1(
        P2_REG0_REG_21__SCAN_IN), .C2(keyinput142), .A(n10205), .ZN(n10210) );
  AOI22_X1 U11295 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(keyinput241), .B1(
        P1_D_REG_4__SCAN_IN), .B2(keyinput252), .ZN(n10206) );
  OAI221_X1 U11296 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(keyinput241), .C1(
        P1_D_REG_4__SCAN_IN), .C2(keyinput252), .A(n10206), .ZN(n10209) );
  AOI22_X1 U11297 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(keyinput224), .B1(SI_25_), .B2(keyinput245), .ZN(n10207) );
  OAI221_X1 U11298 ( .B1(P2_DATAO_REG_6__SCAN_IN), .B2(keyinput224), .C1(
        SI_25_), .C2(keyinput245), .A(n10207), .ZN(n10208) );
  NOR4_X1 U11299 ( .A1(n10211), .A2(n10210), .A3(n10209), .A4(n10208), .ZN(
        n10230) );
  AOI22_X1 U11300 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(keyinput183), .B1(
        P2_IR_REG_20__SCAN_IN), .B2(keyinput155), .ZN(n10212) );
  OAI221_X1 U11301 ( .B1(P1_REG3_REG_8__SCAN_IN), .B2(keyinput183), .C1(
        P2_IR_REG_20__SCAN_IN), .C2(keyinput155), .A(n10212), .ZN(n10219) );
  AOI22_X1 U11302 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(keyinput187), .B1(
        P2_REG2_REG_4__SCAN_IN), .B2(keyinput230), .ZN(n10213) );
  OAI221_X1 U11303 ( .B1(P1_REG3_REG_9__SCAN_IN), .B2(keyinput187), .C1(
        P2_REG2_REG_4__SCAN_IN), .C2(keyinput230), .A(n10213), .ZN(n10218) );
  AOI22_X1 U11304 ( .A1(P1_REG1_REG_22__SCAN_IN), .A2(keyinput149), .B1(
        P1_REG1_REG_9__SCAN_IN), .B2(keyinput151), .ZN(n10214) );
  OAI221_X1 U11305 ( .B1(P1_REG1_REG_22__SCAN_IN), .B2(keyinput149), .C1(
        P1_REG1_REG_9__SCAN_IN), .C2(keyinput151), .A(n10214), .ZN(n10217) );
  AOI22_X1 U11306 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(keyinput164), .B1(
        P1_REG3_REG_28__SCAN_IN), .B2(keyinput165), .ZN(n10215) );
  OAI221_X1 U11307 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(keyinput164), .C1(
        P1_REG3_REG_28__SCAN_IN), .C2(keyinput165), .A(n10215), .ZN(n10216) );
  NOR4_X1 U11308 ( .A1(n10219), .A2(n10218), .A3(n10217), .A4(n10216), .ZN(
        n10229) );
  AOI22_X1 U11309 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(keyinput158), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(keyinput233), .ZN(n10220) );
  OAI221_X1 U11310 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(keyinput158), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput233), .A(n10220), .ZN(n10227) );
  INV_X1 U11311 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n10222) );
  AOI22_X1 U11312 ( .A1(P1_REG0_REG_1__SCAN_IN), .A2(keyinput236), .B1(n10222), 
        .B2(keyinput153), .ZN(n10221) );
  OAI221_X1 U11313 ( .B1(P1_REG0_REG_1__SCAN_IN), .B2(keyinput236), .C1(n10222), .C2(keyinput153), .A(n10221), .ZN(n10225) );
  AOI22_X1 U11314 ( .A1(n10418), .A2(keyinput156), .B1(keyinput152), .B2(
        n10370), .ZN(n10223) );
  OAI221_X1 U11315 ( .B1(n10418), .B2(keyinput156), .C1(n10370), .C2(
        keyinput152), .A(n10223), .ZN(n10224) );
  NOR4_X1 U11316 ( .A1(n10227), .A2(n10226), .A3(n10225), .A4(n10224), .ZN(
        n10228) );
  NAND4_X1 U11317 ( .A1(n10231), .A2(n10230), .A3(n10229), .A4(n10228), .ZN(
        n10337) );
  INV_X1 U11318 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10233) );
  AOI22_X1 U11319 ( .A1(n10234), .A2(keyinput154), .B1(keyinput188), .B2(
        n10233), .ZN(n10232) );
  OAI221_X1 U11320 ( .B1(n10234), .B2(keyinput154), .C1(n10233), .C2(
        keyinput188), .A(n10232), .ZN(n10243) );
  AOI22_X1 U11321 ( .A1(n10341), .A2(keyinput157), .B1(keyinput217), .B2(
        n10392), .ZN(n10235) );
  OAI221_X1 U11322 ( .B1(n10341), .B2(keyinput157), .C1(n10392), .C2(
        keyinput217), .A(n10235), .ZN(n10242) );
  INV_X1 U11323 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10237) );
  AOI22_X1 U11324 ( .A1(n10237), .A2(keyinput184), .B1(n10375), .B2(
        keyinput131), .ZN(n10236) );
  OAI221_X1 U11325 ( .B1(n10237), .B2(keyinput184), .C1(n10375), .C2(
        keyinput131), .A(n10236), .ZN(n10241) );
  INV_X1 U11326 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n10239) );
  AOI22_X1 U11327 ( .A1(n10239), .A2(keyinput176), .B1(n10454), .B2(
        keyinput146), .ZN(n10238) );
  OAI221_X1 U11328 ( .B1(n10239), .B2(keyinput176), .C1(n10454), .C2(
        keyinput146), .A(n10238), .ZN(n10240) );
  NOR4_X1 U11329 ( .A1(n10243), .A2(n10242), .A3(n10241), .A4(n10240), .ZN(
        n10282) );
  INV_X1 U11330 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10245) );
  AOI22_X1 U11331 ( .A1(n10246), .A2(keyinput133), .B1(keyinput253), .B2(
        n10245), .ZN(n10244) );
  OAI221_X1 U11332 ( .B1(n10246), .B2(keyinput133), .C1(n10245), .C2(
        keyinput253), .A(n10244), .ZN(n10255) );
  AOI22_X1 U11333 ( .A1(n6663), .A2(keyinput228), .B1(n10248), .B2(keyinput215), .ZN(n10247) );
  OAI221_X1 U11334 ( .B1(n6663), .B2(keyinput228), .C1(n10248), .C2(
        keyinput215), .A(n10247), .ZN(n10254) );
  AOI22_X1 U11335 ( .A1(n10404), .A2(keyinput170), .B1(keyinput220), .B2(
        n10409), .ZN(n10249) );
  OAI221_X1 U11336 ( .B1(n10404), .B2(keyinput170), .C1(n10409), .C2(
        keyinput220), .A(n10249), .ZN(n10253) );
  XOR2_X1 U11337 ( .A(n10360), .B(keyinput197), .Z(n10251) );
  XNOR2_X1 U11338 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(keyinput221), .ZN(n10250)
         );
  NAND2_X1 U11339 ( .A1(n10251), .A2(n10250), .ZN(n10252) );
  NOR4_X1 U11340 ( .A1(n10255), .A2(n10254), .A3(n10253), .A4(n10252), .ZN(
        n10281) );
  AOI22_X1 U11341 ( .A1(n10424), .A2(keyinput130), .B1(keyinput150), .B2(
        n10451), .ZN(n10256) );
  OAI221_X1 U11342 ( .B1(n10424), .B2(keyinput130), .C1(n10451), .C2(
        keyinput150), .A(n10256), .ZN(n10265) );
  XNOR2_X1 U11343 ( .A(P1_REG3_REG_1__SCAN_IN), .B(keyinput227), .ZN(n10260)
         );
  XNOR2_X1 U11344 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(keyinput232), .ZN(n10259)
         );
  XNOR2_X1 U11345 ( .A(P2_REG0_REG_22__SCAN_IN), .B(keyinput216), .ZN(n10258)
         );
  XNOR2_X1 U11346 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput242), .ZN(n10257) );
  NAND4_X1 U11347 ( .A1(n10260), .A2(n10259), .A3(n10258), .A4(n10257), .ZN(
        n10264) );
  XNOR2_X1 U11348 ( .A(keyinput202), .B(n5867), .ZN(n10263) );
  INV_X1 U11349 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10261) );
  XNOR2_X1 U11350 ( .A(keyinput174), .B(n10261), .ZN(n10262) );
  NOR4_X1 U11351 ( .A1(n10265), .A2(n10264), .A3(n10263), .A4(n10262), .ZN(
        n10280) );
  INV_X1 U11352 ( .A(SI_24_), .ZN(n10267) );
  AOI22_X1 U11353 ( .A1(n10439), .A2(keyinput250), .B1(n10267), .B2(
        keyinput178), .ZN(n10266) );
  OAI221_X1 U11354 ( .B1(n10439), .B2(keyinput250), .C1(n10267), .C2(
        keyinput178), .A(n10266), .ZN(n10274) );
  AOI22_X1 U11355 ( .A1(n10270), .A2(keyinput163), .B1(n10269), .B2(
        keyinput208), .ZN(n10268) );
  OAI221_X1 U11356 ( .B1(n10270), .B2(keyinput163), .C1(n10269), .C2(
        keyinput208), .A(n10268), .ZN(n10273) );
  XNOR2_X1 U11357 ( .A(n10271), .B(keyinput137), .ZN(n10272) );
  OR3_X1 U11358 ( .A1(n10274), .A2(n10273), .A3(n10272), .ZN(n10278) );
  INV_X1 U11359 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10448) );
  AOI22_X1 U11360 ( .A1(n5796), .A2(keyinput147), .B1(keyinput206), .B2(n10448), .ZN(n10275) );
  OAI221_X1 U11361 ( .B1(n5796), .B2(keyinput147), .C1(n10448), .C2(
        keyinput206), .A(n10275), .ZN(n10277) );
  XNOR2_X1 U11362 ( .A(n10419), .B(keyinput198), .ZN(n10276) );
  NOR3_X1 U11363 ( .A1(n10278), .A2(n10277), .A3(n10276), .ZN(n10279) );
  NAND4_X1 U11364 ( .A1(n10282), .A2(n10281), .A3(n10280), .A4(n10279), .ZN(
        n10336) );
  AOI22_X1 U11365 ( .A1(n10284), .A2(keyinput191), .B1(n7754), .B2(keyinput195), .ZN(n10283) );
  OAI221_X1 U11366 ( .B1(n10284), .B2(keyinput191), .C1(n7754), .C2(
        keyinput195), .A(n10283), .ZN(n10294) );
  AOI22_X1 U11367 ( .A1(n10484), .A2(keyinput143), .B1(keyinput200), .B2(
        n10438), .ZN(n10285) );
  OAI221_X1 U11368 ( .B1(n10484), .B2(keyinput143), .C1(n10438), .C2(
        keyinput200), .A(n10285), .ZN(n10293) );
  AOI22_X1 U11369 ( .A1(n10288), .A2(keyinput199), .B1(n10287), .B2(
        keyinput234), .ZN(n10286) );
  OAI221_X1 U11370 ( .B1(n10288), .B2(keyinput199), .C1(n10287), .C2(
        keyinput234), .A(n10286), .ZN(n10292) );
  XOR2_X1 U11371 ( .A(n7273), .B(keyinput160), .Z(n10290) );
  XNOR2_X1 U11372 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput177), .ZN(n10289) );
  NAND2_X1 U11373 ( .A1(n10290), .A2(n10289), .ZN(n10291) );
  NOR4_X1 U11374 ( .A1(n10294), .A2(n10293), .A3(n10292), .A4(n10291), .ZN(
        n10334) );
  AOI22_X1 U11375 ( .A1(n10297), .A2(keyinput239), .B1(keyinput162), .B2(
        n10296), .ZN(n10295) );
  OAI221_X1 U11376 ( .B1(n10297), .B2(keyinput239), .C1(n10296), .C2(
        keyinput162), .A(n10295), .ZN(n10305) );
  INV_X1 U11377 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U11378 ( .A1(n10355), .A2(keyinput190), .B1(keyinput192), .B2(
        n10432), .ZN(n10298) );
  OAI221_X1 U11379 ( .B1(n10355), .B2(keyinput190), .C1(n10432), .C2(
        keyinput192), .A(n10298), .ZN(n10304) );
  AOI22_X1 U11380 ( .A1(n5760), .A2(keyinput144), .B1(n10407), .B2(keyinput128), .ZN(n10299) );
  OAI221_X1 U11381 ( .B1(n5760), .B2(keyinput144), .C1(n10407), .C2(
        keyinput128), .A(n10299), .ZN(n10303) );
  XNOR2_X1 U11382 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(keyinput214), .ZN(n10301)
         );
  XNOR2_X1 U11383 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput237), .ZN(n10300) );
  NAND2_X1 U11384 ( .A1(n10301), .A2(n10300), .ZN(n10302) );
  NOR4_X1 U11385 ( .A1(n10305), .A2(n10304), .A3(n10303), .A4(n10302), .ZN(
        n10333) );
  AOI22_X1 U11386 ( .A1(n10363), .A2(keyinput251), .B1(keyinput181), .B2(
        n10307), .ZN(n10306) );
  OAI221_X1 U11387 ( .B1(n10363), .B2(keyinput251), .C1(n10307), .C2(
        keyinput181), .A(n10306), .ZN(n10317) );
  AOI22_X1 U11388 ( .A1(n10373), .A2(keyinput161), .B1(keyinput219), .B2(n6058), .ZN(n10308) );
  OAI221_X1 U11389 ( .B1(n10373), .B2(keyinput161), .C1(n6058), .C2(
        keyinput219), .A(n10308), .ZN(n10316) );
  AOI22_X1 U11390 ( .A1(n10311), .A2(keyinput186), .B1(n10310), .B2(
        keyinput175), .ZN(n10309) );
  OAI221_X1 U11391 ( .B1(n10311), .B2(keyinput186), .C1(n10310), .C2(
        keyinput175), .A(n10309), .ZN(n10315) );
  XOR2_X1 U11392 ( .A(n10485), .B(keyinput171), .Z(n10313) );
  XNOR2_X1 U11393 ( .A(P2_IR_REG_15__SCAN_IN), .B(keyinput248), .ZN(n10312) );
  NAND2_X1 U11394 ( .A1(n10313), .A2(n10312), .ZN(n10314) );
  NOR4_X1 U11395 ( .A1(n10317), .A2(n10316), .A3(n10315), .A4(n10314), .ZN(
        n10332) );
  AOI22_X1 U11396 ( .A1(n10320), .A2(keyinput129), .B1(keyinput148), .B2(
        n10319), .ZN(n10318) );
  OAI221_X1 U11397 ( .B1(n10320), .B2(keyinput129), .C1(n10319), .C2(
        keyinput148), .A(n10318), .ZN(n10330) );
  AOI22_X1 U11398 ( .A1(n10323), .A2(keyinput229), .B1(keyinput244), .B2(
        n10322), .ZN(n10321) );
  OAI221_X1 U11399 ( .B1(n10323), .B2(keyinput229), .C1(n10322), .C2(
        keyinput244), .A(n10321), .ZN(n10329) );
  AOI22_X1 U11400 ( .A1(n10422), .A2(keyinput159), .B1(n10325), .B2(
        keyinput135), .ZN(n10324) );
  OAI221_X1 U11401 ( .B1(n10422), .B2(keyinput159), .C1(n10325), .C2(
        keyinput135), .A(n10324), .ZN(n10328) );
  AOI22_X1 U11402 ( .A1(n10364), .A2(keyinput240), .B1(n5465), .B2(keyinput247), .ZN(n10326) );
  OAI221_X1 U11403 ( .B1(n10364), .B2(keyinput240), .C1(n5465), .C2(
        keyinput247), .A(n10326), .ZN(n10327) );
  NOR4_X1 U11404 ( .A1(n10330), .A2(n10329), .A3(n10328), .A4(n10327), .ZN(
        n10331) );
  NAND4_X1 U11405 ( .A1(n10334), .A2(n10333), .A3(n10332), .A4(n10331), .ZN(
        n10335) );
  NOR4_X1 U11406 ( .A1(n10338), .A2(n10337), .A3(n10336), .A4(n10335), .ZN(
        n10544) );
  AOI22_X1 U11407 ( .A1(n10341), .A2(keyinput29), .B1(keyinput108), .B2(n10340), .ZN(n10339) );
  OAI221_X1 U11408 ( .B1(n10341), .B2(keyinput29), .C1(n10340), .C2(
        keyinput108), .A(n10339), .ZN(n10352) );
  AOI22_X1 U11409 ( .A1(n10343), .A2(keyinput54), .B1(n7273), .B2(keyinput32), 
        .ZN(n10342) );
  OAI221_X1 U11410 ( .B1(n10343), .B2(keyinput54), .C1(n7273), .C2(keyinput32), 
        .A(n10342), .ZN(n10351) );
  INV_X1 U11411 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n10345) );
  AOI22_X1 U11412 ( .A1(n10346), .A2(keyinput75), .B1(n10345), .B2(keyinput57), 
        .ZN(n10344) );
  OAI221_X1 U11413 ( .B1(n10346), .B2(keyinput75), .C1(n10345), .C2(keyinput57), .A(n10344), .ZN(n10350) );
  XNOR2_X1 U11414 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput96), .ZN(n10348)
         );
  XNOR2_X1 U11415 ( .A(P2_REG1_REG_16__SCAN_IN), .B(keyinput101), .ZN(n10347)
         );
  NAND2_X1 U11416 ( .A1(n10348), .A2(n10347), .ZN(n10349) );
  NOR4_X1 U11417 ( .A1(n10352), .A2(n10351), .A3(n10350), .A4(n10349), .ZN(
        n10402) );
  AOI22_X1 U11418 ( .A1(n7754), .A2(keyinput67), .B1(n5781), .B2(keyinput40), 
        .ZN(n10353) );
  OAI221_X1 U11419 ( .B1(n7754), .B2(keyinput67), .C1(n5781), .C2(keyinput40), 
        .A(n10353), .ZN(n10358) );
  XNOR2_X1 U11420 ( .A(n10354), .B(keyinput109), .ZN(n10357) );
  XNOR2_X1 U11421 ( .A(n10355), .B(keyinput62), .ZN(n10356) );
  OR3_X1 U11422 ( .A1(n10358), .A2(n10357), .A3(n10356), .ZN(n10367) );
  AOI22_X1 U11423 ( .A1(n10361), .A2(keyinput37), .B1(keyinput69), .B2(n10360), 
        .ZN(n10359) );
  OAI221_X1 U11424 ( .B1(n10361), .B2(keyinput37), .C1(n10360), .C2(keyinput69), .A(n10359), .ZN(n10366) );
  AOI22_X1 U11425 ( .A1(n10364), .A2(keyinput112), .B1(n10363), .B2(
        keyinput123), .ZN(n10362) );
  OAI221_X1 U11426 ( .B1(n10364), .B2(keyinput112), .C1(n10363), .C2(
        keyinput123), .A(n10362), .ZN(n10365) );
  NOR3_X1 U11427 ( .A1(n10367), .A2(n10366), .A3(n10365), .ZN(n10401) );
  AOI22_X1 U11428 ( .A1(n10370), .A2(keyinput24), .B1(n10369), .B2(keyinput95), 
        .ZN(n10368) );
  OAI221_X1 U11429 ( .B1(n10370), .B2(keyinput24), .C1(n10369), .C2(keyinput95), .A(n10368), .ZN(n10383) );
  AOI22_X1 U11430 ( .A1(n10373), .A2(keyinput33), .B1(keyinput17), .B2(n10372), 
        .ZN(n10371) );
  OAI221_X1 U11431 ( .B1(n10373), .B2(keyinput33), .C1(n10372), .C2(keyinput17), .A(n10371), .ZN(n10382) );
  AOI22_X1 U11432 ( .A1(n10376), .A2(keyinput98), .B1(keyinput3), .B2(n10375), 
        .ZN(n10374) );
  OAI221_X1 U11433 ( .B1(n10376), .B2(keyinput98), .C1(n10375), .C2(keyinput3), 
        .A(n10374), .ZN(n10381) );
  INV_X1 U11434 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U11435 ( .A1(n10379), .A2(keyinput102), .B1(keyinput85), .B2(n10378), .ZN(n10377) );
  OAI221_X1 U11436 ( .B1(n10379), .B2(keyinput102), .C1(n10378), .C2(
        keyinput85), .A(n10377), .ZN(n10380) );
  NOR4_X1 U11437 ( .A1(n10383), .A2(n10382), .A3(n10381), .A4(n10380), .ZN(
        n10400) );
  INV_X1 U11438 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U11439 ( .A1(n10386), .A2(keyinput12), .B1(keyinput97), .B2(n10385), 
        .ZN(n10384) );
  OAI221_X1 U11440 ( .B1(n10386), .B2(keyinput12), .C1(n10385), .C2(keyinput97), .A(n10384), .ZN(n10398) );
  AOI22_X1 U11441 ( .A1(n10389), .A2(keyinput10), .B1(keyinput76), .B2(n10388), 
        .ZN(n10387) );
  OAI221_X1 U11442 ( .B1(n10389), .B2(keyinput10), .C1(n10388), .C2(keyinput76), .A(n10387), .ZN(n10397) );
  AOI22_X1 U11443 ( .A1(n10392), .A2(keyinput89), .B1(keyinput38), .B2(n10391), 
        .ZN(n10390) );
  OAI221_X1 U11444 ( .B1(n10392), .B2(keyinput89), .C1(n10391), .C2(keyinput38), .A(n10390), .ZN(n10396) );
  AOI22_X1 U11445 ( .A1(n10394), .A2(keyinput21), .B1(n5174), .B2(keyinput55), 
        .ZN(n10393) );
  OAI221_X1 U11446 ( .B1(n10394), .B2(keyinput21), .C1(n5174), .C2(keyinput55), 
        .A(n10393), .ZN(n10395) );
  NOR4_X1 U11447 ( .A1(n10398), .A2(n10397), .A3(n10396), .A4(n10395), .ZN(
        n10399) );
  NAND4_X1 U11448 ( .A1(n10402), .A2(n10401), .A3(n10400), .A4(n10399), .ZN(
        n10543) );
  INV_X1 U11449 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10405) );
  AOI22_X1 U11450 ( .A1(n10405), .A2(keyinput44), .B1(n10404), .B2(keyinput42), 
        .ZN(n10403) );
  OAI221_X1 U11451 ( .B1(n10405), .B2(keyinput44), .C1(n10404), .C2(keyinput42), .A(n10403), .ZN(n10416) );
  AOI22_X1 U11452 ( .A1(n6663), .A2(keyinput100), .B1(n10407), .B2(keyinput0), 
        .ZN(n10406) );
  OAI221_X1 U11453 ( .B1(n6663), .B2(keyinput100), .C1(n10407), .C2(keyinput0), 
        .A(n10406), .ZN(n10415) );
  AOI22_X1 U11454 ( .A1(n10410), .A2(keyinput14), .B1(keyinput92), .B2(n10409), 
        .ZN(n10408) );
  OAI221_X1 U11455 ( .B1(n10410), .B2(keyinput14), .C1(n10409), .C2(keyinput92), .A(n10408), .ZN(n10414) );
  XNOR2_X1 U11456 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput9), .ZN(n10412) );
  XNOR2_X1 U11457 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(keyinput93), .ZN(n10411)
         );
  NAND2_X1 U11458 ( .A1(n10412), .A2(n10411), .ZN(n10413) );
  NOR4_X1 U11459 ( .A1(n10416), .A2(n10415), .A3(n10414), .A4(n10413), .ZN(
        n10464) );
  AOI22_X1 U11460 ( .A1(n10419), .A2(keyinput70), .B1(n10418), .B2(keyinput28), 
        .ZN(n10417) );
  OAI221_X1 U11461 ( .B1(n10419), .B2(keyinput70), .C1(n10418), .C2(keyinput28), .A(n10417), .ZN(n10430) );
  AOI22_X1 U11462 ( .A1(n10422), .A2(keyinput31), .B1(keyinput84), .B2(n10421), 
        .ZN(n10420) );
  OAI221_X1 U11463 ( .B1(n10422), .B2(keyinput31), .C1(n10421), .C2(keyinput84), .A(n10420), .ZN(n10429) );
  AOI22_X1 U11464 ( .A1(P2_U3151), .A2(keyinput45), .B1(keyinput2), .B2(n10424), .ZN(n10423) );
  OAI221_X1 U11465 ( .B1(P2_U3151), .B2(keyinput45), .C1(n10424), .C2(
        keyinput2), .A(n10423), .ZN(n10428) );
  XNOR2_X1 U11466 ( .A(P2_REG0_REG_22__SCAN_IN), .B(keyinput88), .ZN(n10426)
         );
  XNOR2_X1 U11467 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput13), .ZN(n10425) );
  NAND2_X1 U11468 ( .A1(n10426), .A2(n10425), .ZN(n10427) );
  NOR4_X1 U11469 ( .A1(n10430), .A2(n10429), .A3(n10428), .A4(n10427), .ZN(
        n10463) );
  AOI22_X1 U11470 ( .A1(n10433), .A2(keyinput61), .B1(keyinput64), .B2(n10432), 
        .ZN(n10431) );
  OAI221_X1 U11471 ( .B1(n10433), .B2(keyinput61), .C1(n10432), .C2(keyinput64), .A(n10431), .ZN(n10445) );
  AOI22_X1 U11472 ( .A1(n10436), .A2(keyinput27), .B1(keyinput83), .B2(n10435), 
        .ZN(n10434) );
  OAI221_X1 U11473 ( .B1(n10436), .B2(keyinput27), .C1(n10435), .C2(keyinput83), .A(n10434), .ZN(n10444) );
  AOI22_X1 U11474 ( .A1(n10439), .A2(keyinput122), .B1(n10438), .B2(keyinput72), .ZN(n10437) );
  OAI221_X1 U11475 ( .B1(n10439), .B2(keyinput122), .C1(n10438), .C2(
        keyinput72), .A(n10437), .ZN(n10443) );
  XOR2_X1 U11476 ( .A(n5465), .B(keyinput119), .Z(n10441) );
  XNOR2_X1 U11477 ( .A(P2_IR_REG_15__SCAN_IN), .B(keyinput120), .ZN(n10440) );
  NAND2_X1 U11478 ( .A1(n10441), .A2(n10440), .ZN(n10442) );
  NOR4_X1 U11479 ( .A1(n10445), .A2(n10444), .A3(n10443), .A4(n10442), .ZN(
        n10462) );
  AOI22_X1 U11480 ( .A1(n10448), .A2(keyinput78), .B1(n10447), .B2(keyinput6), 
        .ZN(n10446) );
  OAI221_X1 U11481 ( .B1(n10448), .B2(keyinput78), .C1(n10447), .C2(keyinput6), 
        .A(n10446), .ZN(n10460) );
  INV_X1 U11482 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10450) );
  AOI22_X1 U11483 ( .A1(n10451), .A2(keyinput22), .B1(keyinput113), .B2(n10450), .ZN(n10449) );
  OAI221_X1 U11484 ( .B1(n10451), .B2(keyinput22), .C1(n10450), .C2(
        keyinput113), .A(n10449), .ZN(n10459) );
  AOI22_X1 U11485 ( .A1(n10454), .A2(keyinput18), .B1(keyinput127), .B2(n10453), .ZN(n10452) );
  OAI221_X1 U11486 ( .B1(n10454), .B2(keyinput18), .C1(n10453), .C2(
        keyinput127), .A(n10452), .ZN(n10458) );
  XNOR2_X1 U11487 ( .A(P1_REG3_REG_1__SCAN_IN), .B(keyinput99), .ZN(n10456) );
  XNOR2_X1 U11488 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(keyinput104), .ZN(n10455)
         );
  NAND2_X1 U11489 ( .A1(n10456), .A2(n10455), .ZN(n10457) );
  NOR4_X1 U11490 ( .A1(n10460), .A2(n10459), .A3(n10458), .A4(n10457), .ZN(
        n10461) );
  NAND4_X1 U11491 ( .A1(n10464), .A2(n10463), .A3(n10462), .A4(n10461), .ZN(
        n10542) );
  OAI22_X1 U11492 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(keyinput114), .B1(
        keyinput50), .B2(SI_24_), .ZN(n10465) );
  AOI221_X1 U11493 ( .B1(P2_IR_REG_13__SCAN_IN), .B2(keyinput114), .C1(SI_24_), 
        .C2(keyinput50), .A(n10465), .ZN(n10472) );
  OAI22_X1 U11494 ( .A1(P2_REG2_REG_24__SCAN_IN), .A2(keyinput91), .B1(
        P1_REG1_REG_26__SCAN_IN), .B2(keyinput73), .ZN(n10466) );
  AOI221_X1 U11495 ( .B1(P2_REG2_REG_24__SCAN_IN), .B2(keyinput91), .C1(
        keyinput73), .C2(P1_REG1_REG_26__SCAN_IN), .A(n10466), .ZN(n10471) );
  OAI22_X1 U11496 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(keyinput103), .B1(
        keyinput86), .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n10467) );
  AOI221_X1 U11497 ( .B1(P2_DATAO_REG_24__SCAN_IN), .B2(keyinput103), .C1(
        P1_DATAO_REG_15__SCAN_IN), .C2(keyinput86), .A(n10467), .ZN(n10470) );
  OAI22_X1 U11498 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput110), .B1(
        keyinput94), .B2(P1_REG2_REG_14__SCAN_IN), .ZN(n10468) );
  AOI221_X1 U11499 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput110), .C1(
        P1_REG2_REG_14__SCAN_IN), .C2(keyinput94), .A(n10468), .ZN(n10469) );
  NAND4_X1 U11500 ( .A1(n10472), .A2(n10471), .A3(n10470), .A4(n10469), .ZN(
        n10502) );
  OAI22_X1 U11501 ( .A1(P2_REG1_REG_21__SCAN_IN), .A2(keyinput47), .B1(
        P1_REG0_REG_10__SCAN_IN), .B2(keyinput125), .ZN(n10473) );
  AOI221_X1 U11502 ( .B1(P2_REG1_REG_21__SCAN_IN), .B2(keyinput47), .C1(
        keyinput125), .C2(P1_REG0_REG_10__SCAN_IN), .A(n10473), .ZN(n10480) );
  OAI22_X1 U11503 ( .A1(P2_REG2_REG_3__SCAN_IN), .A2(keyinput39), .B1(
        P1_REG3_REG_7__SCAN_IN), .B2(keyinput56), .ZN(n10474) );
  AOI221_X1 U11504 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(keyinput39), .C1(
        keyinput56), .C2(P1_REG3_REG_7__SCAN_IN), .A(n10474), .ZN(n10479) );
  OAI22_X1 U11505 ( .A1(P1_D_REG_26__SCAN_IN), .A2(keyinput1), .B1(keyinput34), 
        .B2(P1_REG3_REG_4__SCAN_IN), .ZN(n10475) );
  AOI221_X1 U11506 ( .B1(P1_D_REG_26__SCAN_IN), .B2(keyinput1), .C1(
        P1_REG3_REG_4__SCAN_IN), .C2(keyinput34), .A(n10475), .ZN(n10478) );
  OAI22_X1 U11507 ( .A1(P1_REG1_REG_29__SCAN_IN), .A2(keyinput35), .B1(
        keyinput87), .B2(P1_REG0_REG_26__SCAN_IN), .ZN(n10476) );
  AOI221_X1 U11508 ( .B1(P1_REG1_REG_29__SCAN_IN), .B2(keyinput35), .C1(
        P1_REG0_REG_26__SCAN_IN), .C2(keyinput87), .A(n10476), .ZN(n10477) );
  NAND4_X1 U11509 ( .A1(n10480), .A2(n10479), .A3(n10478), .A4(n10477), .ZN(
        n10501) );
  OAI22_X1 U11510 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(keyinput52), .B1(keyinput65), .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n10481) );
  AOI221_X1 U11511 ( .B1(P2_IR_REG_9__SCAN_IN), .B2(keyinput52), .C1(
        P2_DATAO_REG_13__SCAN_IN), .C2(keyinput65), .A(n10481), .ZN(n10491) );
  OAI22_X1 U11512 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput124), .B1(keyinput58), .B2(P1_ADDR_REG_5__SCAN_IN), .ZN(n10482) );
  AOI221_X1 U11513 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput124), .C1(
        P1_ADDR_REG_5__SCAN_IN), .C2(keyinput58), .A(n10482), .ZN(n10490) );
  OAI22_X1 U11514 ( .A1(n10485), .A2(keyinput43), .B1(n10484), .B2(keyinput15), 
        .ZN(n10483) );
  AOI221_X1 U11515 ( .B1(n10485), .B2(keyinput43), .C1(keyinput15), .C2(n10484), .A(n10483), .ZN(n10489) );
  OAI22_X1 U11516 ( .A1(n10487), .A2(keyinput68), .B1(keyinput107), .B2(
        P1_REG0_REG_14__SCAN_IN), .ZN(n10486) );
  AOI221_X1 U11517 ( .B1(n10487), .B2(keyinput68), .C1(P1_REG0_REG_14__SCAN_IN), .C2(keyinput107), .A(n10486), .ZN(n10488) );
  NAND4_X1 U11518 ( .A1(n10491), .A2(n10490), .A3(n10489), .A4(n10488), .ZN(
        n10500) );
  OAI22_X1 U11519 ( .A1(P2_D_REG_18__SCAN_IN), .A2(keyinput106), .B1(
        P1_REG0_REG_15__SCAN_IN), .B2(keyinput11), .ZN(n10492) );
  AOI221_X1 U11520 ( .B1(P2_D_REG_18__SCAN_IN), .B2(keyinput106), .C1(
        keyinput11), .C2(P1_REG0_REG_15__SCAN_IN), .A(n10492), .ZN(n10497) );
  OAI22_X1 U11521 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(keyinput79), .B1(
        keyinput82), .B2(P1_REG1_REG_17__SCAN_IN), .ZN(n10493) );
  AOI221_X1 U11522 ( .B1(P2_IR_REG_26__SCAN_IN), .B2(keyinput79), .C1(
        P1_REG1_REG_17__SCAN_IN), .C2(keyinput82), .A(n10493), .ZN(n10496) );
  OAI22_X1 U11523 ( .A1(P2_D_REG_30__SCAN_IN), .A2(keyinput77), .B1(
        P1_REG3_REG_9__SCAN_IN), .B2(keyinput59), .ZN(n10494) );
  AOI221_X1 U11524 ( .B1(P2_D_REG_30__SCAN_IN), .B2(keyinput77), .C1(
        keyinput59), .C2(P1_REG3_REG_9__SCAN_IN), .A(n10494), .ZN(n10495) );
  NAND4_X1 U11525 ( .A1(n10498), .A2(n10497), .A3(n10496), .A4(n10495), .ZN(
        n10499) );
  NOR4_X1 U11526 ( .A1(n10502), .A2(n10501), .A3(n10500), .A4(n10499), .ZN(
        n10540) );
  OAI22_X1 U11527 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(keyinput5), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(keyinput118), .ZN(n10503) );
  AOI221_X1 U11528 ( .B1(P1_DATAO_REG_26__SCAN_IN), .B2(keyinput5), .C1(
        keyinput118), .C2(P1_REG3_REG_0__SCAN_IN), .A(n10503), .ZN(n10510) );
  OAI22_X1 U11529 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(keyinput121), .B1(
        P1_REG0_REG_4__SCAN_IN), .B2(keyinput126), .ZN(n10504) );
  AOI221_X1 U11530 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(keyinput121), .C1(
        keyinput126), .C2(P1_REG0_REG_4__SCAN_IN), .A(n10504), .ZN(n10509) );
  OAI22_X1 U11531 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(keyinput71), .B1(
        keyinput74), .B2(P2_REG0_REG_9__SCAN_IN), .ZN(n10505) );
  AOI221_X1 U11532 ( .B1(P1_DATAO_REG_8__SCAN_IN), .B2(keyinput71), .C1(
        P2_REG0_REG_9__SCAN_IN), .C2(keyinput74), .A(n10505), .ZN(n10508) );
  OAI22_X1 U11533 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput66), .B1(
        keyinput81), .B2(P1_REG3_REG_20__SCAN_IN), .ZN(n10506) );
  AOI221_X1 U11534 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput66), .C1(
        P1_REG3_REG_20__SCAN_IN), .C2(keyinput81), .A(n10506), .ZN(n10507) );
  NAND4_X1 U11535 ( .A1(n10510), .A2(n10509), .A3(n10508), .A4(n10507), .ZN(
        n10538) );
  OAI22_X1 U11536 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(keyinput36), .B1(
        keyinput25), .B2(P1_REG2_REG_28__SCAN_IN), .ZN(n10511) );
  AOI221_X1 U11537 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(keyinput36), .C1(
        P1_REG2_REG_28__SCAN_IN), .C2(keyinput25), .A(n10511), .ZN(n10518) );
  OAI22_X1 U11538 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(keyinput41), .B1(
        P1_IR_REG_22__SCAN_IN), .B2(keyinput115), .ZN(n10512) );
  AOI221_X1 U11539 ( .B1(P1_DATAO_REG_19__SCAN_IN), .B2(keyinput41), .C1(
        keyinput115), .C2(P1_IR_REG_22__SCAN_IN), .A(n10512), .ZN(n10517) );
  OAI22_X1 U11540 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput4), .B1(
        keyinput26), .B2(P2_REG1_REG_20__SCAN_IN), .ZN(n10513) );
  AOI221_X1 U11541 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput4), .C1(
        P2_REG1_REG_20__SCAN_IN), .C2(keyinput26), .A(n10513), .ZN(n10516) );
  OAI22_X1 U11542 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(keyinput53), .B1(
        P2_ADDR_REG_1__SCAN_IN), .B2(keyinput63), .ZN(n10514) );
  AOI221_X1 U11543 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(keyinput53), .C1(
        keyinput63), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n10514), .ZN(n10515) );
  NAND4_X1 U11544 ( .A1(n10518), .A2(n10517), .A3(n10516), .A4(n10515), .ZN(
        n10537) );
  OAI22_X1 U11545 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput105), .B1(
        P2_REG2_REG_1__SCAN_IN), .B2(keyinput16), .ZN(n10519) );
  AOI221_X1 U11546 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput105), .C1(
        keyinput16), .C2(P2_REG2_REG_1__SCAN_IN), .A(n10519), .ZN(n10526) );
  OAI22_X1 U11547 ( .A1(P2_REG1_REG_30__SCAN_IN), .A2(keyinput80), .B1(
        P1_REG1_REG_9__SCAN_IN), .B2(keyinput23), .ZN(n10520) );
  AOI221_X1 U11548 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(keyinput80), .C1(
        keyinput23), .C2(P1_REG1_REG_9__SCAN_IN), .A(n10520), .ZN(n10525) );
  OAI22_X1 U11549 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(keyinput30), .B1(
        keyinput8), .B2(P2_REG1_REG_6__SCAN_IN), .ZN(n10521) );
  AOI221_X1 U11550 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(keyinput30), .C1(
        P2_REG1_REG_6__SCAN_IN), .C2(keyinput8), .A(n10521), .ZN(n10524) );
  OAI22_X1 U11551 ( .A1(SI_25_), .A2(keyinput117), .B1(keyinput90), .B2(
        P2_REG2_REG_5__SCAN_IN), .ZN(n10522) );
  AOI221_X1 U11552 ( .B1(SI_25_), .B2(keyinput117), .C1(P2_REG2_REG_5__SCAN_IN), .C2(keyinput90), .A(n10522), .ZN(n10523) );
  NAND4_X1 U11553 ( .A1(n10526), .A2(n10525), .A3(n10524), .A4(n10523), .ZN(
        n10536) );
  OAI22_X1 U11554 ( .A1(P1_REG2_REG_31__SCAN_IN), .A2(keyinput48), .B1(
        P2_ADDR_REG_10__SCAN_IN), .B2(keyinput116), .ZN(n10527) );
  AOI221_X1 U11555 ( .B1(P1_REG2_REG_31__SCAN_IN), .B2(keyinput48), .C1(
        keyinput116), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n10527), .ZN(n10534) );
  OAI22_X1 U11556 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(keyinput19), .B1(
        P1_IR_REG_31__SCAN_IN), .B2(keyinput49), .ZN(n10528) );
  AOI221_X1 U11557 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(keyinput19), .C1(
        keyinput49), .C2(P1_IR_REG_31__SCAN_IN), .A(n10528), .ZN(n10533) );
  OAI22_X1 U11558 ( .A1(SI_12_), .A2(keyinput7), .B1(keyinput60), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n10529) );
  AOI221_X1 U11559 ( .B1(SI_12_), .B2(keyinput7), .C1(P1_REG0_REG_17__SCAN_IN), 
        .C2(keyinput60), .A(n10529), .ZN(n10532) );
  OAI22_X1 U11560 ( .A1(P2_REG0_REG_25__SCAN_IN), .A2(keyinput111), .B1(
        P1_REG0_REG_12__SCAN_IN), .B2(keyinput46), .ZN(n10530) );
  AOI221_X1 U11561 ( .B1(P2_REG0_REG_25__SCAN_IN), .B2(keyinput111), .C1(
        keyinput46), .C2(P1_REG0_REG_12__SCAN_IN), .A(n10530), .ZN(n10531) );
  NAND4_X1 U11562 ( .A1(n10534), .A2(n10533), .A3(n10532), .A4(n10531), .ZN(
        n10535) );
  NOR4_X1 U11563 ( .A1(n10538), .A2(n10537), .A3(n10536), .A4(n10535), .ZN(
        n10539) );
  NAND2_X1 U11564 ( .A1(n10540), .A2(n10539), .ZN(n10541) );
  NOR4_X1 U11565 ( .A1(n10544), .A2(n10543), .A3(n10542), .A4(n10541), .ZN(
        n10545) );
  XNOR2_X1 U11566 ( .A(n10546), .B(n10545), .ZN(P2_U3187) );
  XOR2_X1 U11567 ( .A(n10547), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1068_U50) );
  NOR2_X1 U11568 ( .A1(n10549), .A2(n10548), .ZN(n10550) );
  XOR2_X1 U11569 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10550), .Z(ADD_1068_U51) );
  XOR2_X1 U11570 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10551), .Z(ADD_1068_U47) );
  XOR2_X1 U11571 ( .A(n10552), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1068_U49) );
  XOR2_X1 U11572 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10553), .Z(ADD_1068_U48) );
  XOR2_X1 U11573 ( .A(n10555), .B(n10554), .Z(ADD_1068_U54) );
  XOR2_X1 U11574 ( .A(n10557), .B(n10556), .Z(ADD_1068_U53) );
  XNOR2_X1 U11575 ( .A(n10559), .B(n10558), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U5015 ( .A(n6319), .Z(n4506) );
endmodule

