

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393;

  NAND2_X1 U4788 ( .A1(n5435), .A2(n5434), .ZN(n6484) );
  AND4_X1 U4789 ( .A1(n6446), .A2(n6445), .A3(n6444), .A4(n6443), .ZN(n9200)
         );
  NAND4_X1 U4790 ( .A1(n6434), .A2(n6433), .A3(n6432), .A4(n6431), .ZN(n9429)
         );
  CLKBUF_X1 U4791 ( .A(n6164), .Z(n4282) );
  INV_X1 U4792 ( .A(n6442), .ZN(n6563) );
  CLKBUF_X1 U4793 ( .A(n6164), .Z(n4283) );
  NAND2_X1 U4794 ( .A1(n5648), .A2(n5647), .ZN(n5854) );
  CLKBUF_X2 U4795 ( .A(n5347), .Z(n6990) );
  AOI21_X1 U4796 ( .B1(n4995), .B2(n4993), .A(n8178), .ZN(n4989) );
  INV_X1 U4797 ( .A(n8475), .ZN(n8499) );
  INV_X2 U4798 ( .A(n5754), .ZN(n5749) );
  AND2_X1 U4799 ( .A1(n9693), .A2(n4384), .ZN(n6710) );
  INV_X2 U4801 ( .A(n6164), .ZN(n8312) );
  INV_X2 U4802 ( .A(n5854), .ZN(n8311) );
  NAND2_X1 U4803 ( .A1(n6208), .A2(n7168), .ZN(n7173) );
  AND2_X1 U4804 ( .A1(n5600), .A2(n5599), .ZN(n5595) );
  CLKBUF_X2 U4805 ( .A(n6748), .Z(n6921) );
  INV_X1 U4806 ( .A(n6582), .ZN(n6589) );
  NAND2_X1 U4807 ( .A1(n6712), .A2(n6975), .ZN(n6970) );
  NAND2_X1 U4808 ( .A1(n8036), .A2(n9677), .ZN(n9352) );
  INV_X1 U4809 ( .A(n9429), .ZN(n7666) );
  INV_X1 U4810 ( .A(n7651), .ZN(n7425) );
  XNOR2_X1 U4811 ( .A(n4458), .B(n4713), .ZN(n7004) );
  INV_X2 U4812 ( .A(n9848), .ZN(n10077) );
  AND3_X2 U4813 ( .A1(n4702), .A2(n6031), .A3(n6030), .ZN(n6032) );
  INV_X1 U4814 ( .A(n5854), .ZN(n4281) );
  NAND2_X1 U4815 ( .A1(n5205), .A2(n5204), .ZN(n5365) );
  NOR2_X2 U4816 ( .A1(n6221), .A2(n6323), .ZN(n6222) );
  NOR2_X2 U4817 ( .A1(n5344), .A2(n5340), .ZN(n5582) );
  AOI21_X2 U4818 ( .B1(n6689), .B2(n6691), .A(n6690), .ZN(n6688) );
  INV_X2 U4819 ( .A(n7775), .ZN(n7880) );
  NAND2_X2 U4820 ( .A1(n6797), .A2(n6796), .ZN(n7775) );
  NAND2_X2 U4821 ( .A1(n9774), .A2(n4327), .ZN(n9775) );
  AOI21_X2 U4822 ( .B1(n9796), .B2(n9795), .A(n9388), .ZN(n9774) );
  NOR2_X1 U4823 ( .A1(n6739), .A2(n7425), .ZN(n7402) );
  OAI22_X2 U4824 ( .A1(n7682), .A2(n7681), .B1(n9925), .B2(n7685), .ZN(n9527)
         );
  NAND2_X1 U4825 ( .A1(n5648), .A2(n9055), .ZN(n6164) );
  AOI21_X2 U4826 ( .B1(n10043), .B2(n9549), .A(n10042), .ZN(n10204) );
  NOR2_X2 U4827 ( .A1(n8089), .A2(n8090), .ZN(n7961) );
  OAI21_X2 U4828 ( .B1(n4659), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n5212), .ZN(
        n5213) );
  INV_X4 U4829 ( .A(n6919), .ZN(n6727) );
  XNOR2_X2 U4830 ( .A(n5430), .B(n5429), .ZN(n7042) );
  NAND2_X2 U4831 ( .A1(n4594), .A2(n5243), .ZN(n5430) );
  NAND2_X1 U4832 ( .A1(n7875), .A2(n7997), .ZN(n9286) );
  OAI21_X1 U4833 ( .B1(n7436), .B2(n7437), .A(n6099), .ZN(n4495) );
  NAND2_X1 U4834 ( .A1(n4532), .A2(n5700), .ZN(n5760) );
  INV_X1 U4835 ( .A(n9430), .ZN(n7646) );
  NAND2_X1 U4836 ( .A1(n6057), .A2(n8500), .ZN(n8324) );
  CLKBUF_X3 U4837 ( .A(n6422), .Z(n6959) );
  AND2_X1 U4838 ( .A1(n5585), .A2(n4726), .ZN(n6422) );
  INV_X4 U4839 ( .A(n6911), .ZN(n4284) );
  NAND2_X1 U4840 ( .A1(n5372), .A2(n5366), .ZN(n5392) );
  INV_X4 U4841 ( .A(n5372), .ZN(n5052) );
  INV_X1 U4842 ( .A(n6301), .ZN(n4286) );
  NAND2_X1 U4843 ( .A1(n4465), .A2(n4316), .ZN(n7015) );
  INV_X1 U4844 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n10339) );
  INV_X2 U4845 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4520) );
  AOI21_X1 U4846 ( .B1(n6709), .B2(n9829), .A(n6708), .ZN(n9615) );
  INV_X1 U4847 ( .A(n8620), .ZN(n8650) );
  NAND2_X1 U4848 ( .A1(n4998), .A2(n5001), .ZN(n8620) );
  OAI22_X1 U4849 ( .A1(n6365), .A2(n6149), .B1(n8519), .B2(n8476), .ZN(n4497)
         );
  NAND2_X1 U4850 ( .A1(n4531), .A2(n8245), .ZN(n8610) );
  NAND2_X1 U4851 ( .A1(n9617), .A2(n6661), .ZN(n6663) );
  NAND2_X1 U4852 ( .A1(n4430), .A2(n6684), .ZN(n8839) );
  NAND2_X1 U4853 ( .A1(n8701), .A2(n8244), .ZN(n4531) );
  NAND2_X1 U4854 ( .A1(n8639), .A2(n8638), .ZN(n8701) );
  AND2_X1 U4855 ( .A1(n6972), .A2(n6971), .ZN(n8538) );
  OAI21_X2 U4856 ( .B1(n8888), .B2(n6182), .A(n8463), .ZN(n8878) );
  CLKBUF_X1 U4857 ( .A(n9073), .Z(n4673) );
  NAND2_X1 U4858 ( .A1(n4483), .A2(n5017), .ZN(n8630) );
  NAND2_X1 U4859 ( .A1(n8592), .A2(n4289), .ZN(n4483) );
  AOI22_X1 U4860 ( .A1(n9988), .A2(n8310), .B1(n8309), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n8999) );
  NAND2_X1 U4861 ( .A1(n4422), .A2(n4425), .ZN(n8823) );
  NAND2_X1 U4862 ( .A1(n8811), .A2(n4914), .ZN(n4912) );
  NAND2_X1 U4863 ( .A1(n5869), .A2(n8665), .ZN(n8592) );
  AOI21_X1 U4864 ( .B1(n8588), .B2(n8310), .A(n4408), .ZN(n9002) );
  CLKBUF_X1 U4865 ( .A(n6710), .Z(n9619) );
  NAND2_X1 U4866 ( .A1(n8666), .A2(n8664), .ZN(n5869) );
  NAND2_X1 U4867 ( .A1(n4468), .A2(n4521), .ZN(n8666) );
  OR2_X1 U4868 ( .A1(n9609), .A2(n10374), .ZN(n9312) );
  NAND2_X1 U4869 ( .A1(n9830), .A2(n6502), .ZN(n9811) );
  AND2_X1 U4870 ( .A1(n4522), .A2(n4985), .ZN(n4521) );
  AOI21_X1 U4871 ( .B1(n8798), .B2(n8796), .A(n8797), .ZN(n8795) );
  NAND2_X1 U4872 ( .A1(n4938), .A2(n6315), .ZN(n4943) );
  NAND2_X1 U4873 ( .A1(n4645), .A2(n8778), .ZN(n8796) );
  INV_X1 U4874 ( .A(n9721), .ZN(n9955) );
  NAND2_X1 U4875 ( .A1(n7930), .A2(n4637), .ZN(n8097) );
  NAND2_X1 U4876 ( .A1(n6577), .A2(n6576), .ZN(n9673) );
  OAI21_X1 U4877 ( .B1(n4598), .B2(n4597), .A(n5305), .ZN(n5543) );
  AND2_X1 U4878 ( .A1(n5512), .A2(n5511), .ZN(n9721) );
  NAND2_X1 U4879 ( .A1(n6485), .A2(n4564), .ZN(n7839) );
  AOI21_X1 U4880 ( .B1(n4289), .B2(n8591), .A(n4357), .ZN(n5017) );
  NAND2_X1 U4881 ( .A1(n7936), .A2(n8265), .ZN(n9840) );
  NAND2_X1 U4882 ( .A1(n4440), .A2(n7044), .ZN(n7966) );
  NAND2_X1 U4883 ( .A1(n7563), .A2(n6215), .ZN(n4440) );
  NOR2_X1 U4884 ( .A1(n9547), .A2(n9546), .ZN(n9565) );
  NAND2_X1 U4885 ( .A1(n5502), .A2(n5501), .ZN(n9734) );
  NAND2_X1 U4886 ( .A1(n5491), .A2(n5490), .ZN(n9900) );
  NAND2_X1 U4887 ( .A1(n4921), .A2(n7559), .ZN(n7563) );
  NAND2_X1 U4888 ( .A1(n5479), .A2(n5478), .ZN(n9911) );
  INV_X1 U4889 ( .A(n8403), .ZN(n8012) );
  AOI21_X1 U4890 ( .B1(n7822), .B2(n6637), .A(n5177), .ZN(n7748) );
  NAND2_X1 U4891 ( .A1(n6535), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6553) );
  NAND2_X1 U4892 ( .A1(n5456), .A2(n5455), .ZN(n9924) );
  NAND2_X1 U4893 ( .A1(n5447), .A2(n5446), .ZN(n9228) );
  AND2_X1 U4894 ( .A1(n4332), .A2(n4534), .ZN(n7697) );
  NAND2_X1 U4895 ( .A1(n7535), .A2(n6757), .ZN(n7592) );
  NAND2_X1 U4896 ( .A1(n4495), .A2(n7432), .ZN(n7505) );
  NAND2_X1 U4897 ( .A1(n7902), .A2(n7903), .ZN(n4977) );
  AND2_X1 U4898 ( .A1(n4665), .A2(n4664), .ZN(n7682) );
  AND2_X1 U4899 ( .A1(n6633), .A2(n6632), .ZN(n7895) );
  NAND2_X1 U4900 ( .A1(n4620), .A2(n4622), .ZN(n5449) );
  NAND2_X1 U4901 ( .A1(n6211), .A2(n7328), .ZN(n7372) );
  OAI22_X1 U4902 ( .A1(n7189), .A2(n7188), .B1(n7187), .B2(n7192), .ZN(n7190)
         );
  NAND2_X1 U4903 ( .A1(n4560), .A2(n4559), .ZN(n5415) );
  AND2_X1 U4904 ( .A1(n4445), .A2(n4444), .ZN(n7243) );
  CLKBUF_X1 U4905 ( .A(n6339), .Z(n4706) );
  INV_X1 U4906 ( .A(n5760), .ZN(n6339) );
  CLKBUF_X2 U4907 ( .A(n6740), .Z(n8544) );
  INV_X2 U4908 ( .A(n6740), .ZN(n6888) );
  NAND2_X1 U4909 ( .A1(n5220), .A2(n5219), .ZN(n5397) );
  INV_X2 U4910 ( .A(n6748), .ZN(n8547) );
  NOR2_X1 U4911 ( .A1(n7176), .A2(n4674), .ZN(n6303) );
  INV_X1 U4912 ( .A(n9279), .ZN(n4285) );
  NAND4_X1 U4913 ( .A1(n6427), .A2(n6426), .A3(n6425), .A4(n6424), .ZN(n9430)
         );
  NAND2_X1 U4914 ( .A1(n6159), .A2(n6158), .ZN(n10136) );
  NAND2_X1 U4915 ( .A1(n6666), .A2(n6665), .ZN(n6722) );
  AOI21_X1 U4916 ( .B1(n7100), .B2(n4290), .A(n7174), .ZN(n7176) );
  AND3_X1 U4917 ( .A1(n4535), .A2(n4479), .A3(n4478), .ZN(n8335) );
  BUF_X2 U4918 ( .A(n6911), .Z(n6918) );
  NAND2_X2 U4919 ( .A1(n8338), .A2(n8513), .ZN(n8475) );
  AND4_X1 U4920 ( .A1(n5733), .A2(n5732), .A3(n5731), .A4(n5730), .ZN(n7353)
         );
  AND3_X1 U4921 ( .A1(n5740), .A2(n5057), .A3(n5056), .ZN(n10156) );
  INV_X2 U4922 ( .A(n5773), .ZN(n8310) );
  OR2_X1 U4923 ( .A1(n5568), .A2(n5567), .ZN(n5569) );
  AND2_X1 U4924 ( .A1(n5682), .A2(n5681), .ZN(n8500) );
  XNOR2_X1 U4925 ( .A(n4547), .B(n5678), .ZN(n6057) );
  OAI21_X1 U4926 ( .B1(n5020), .B2(P2_IR_REG_20__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n4547) );
  NAND2_X1 U4927 ( .A1(n5583), .A2(n4727), .ZN(n9996) );
  XNOR2_X1 U4928 ( .A(n10339), .B(n5572), .ZN(n9414) );
  AND2_X1 U4929 ( .A1(n5581), .A2(n5580), .ZN(n4727) );
  NAND2_X1 U4930 ( .A1(n5583), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5584) );
  INV_X1 U4931 ( .A(n6070), .ZN(n6069) );
  NAND2_X2 U4932 ( .A1(n6990), .A2(P2_U3151), .ZN(n9063) );
  NAND2_X1 U4933 ( .A1(n4709), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U4934 ( .A1(n6052), .A2(n5643), .ZN(n6070) );
  INV_X1 U4935 ( .A(n5408), .ZN(n5142) );
  AND2_X1 U4936 ( .A1(n4967), .A2(n5182), .ZN(n4741) );
  NAND3_X1 U4937 ( .A1(n4844), .A2(n4429), .A3(n4628), .ZN(n5664) );
  AND4_X1 U4938 ( .A1(n4980), .A2(n4979), .A3(n4978), .A4(n4463), .ZN(n4811)
         );
  INV_X4 U4939 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U4940 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5597) );
  INV_X1 U4941 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5494) );
  INV_X1 U4942 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5870) );
  INV_X1 U4943 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5678) );
  INV_X4 U4944 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U4945 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4628) );
  NOR2_X1 U4946 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5896) );
  INV_X1 U4947 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5845) );
  NOR2_X1 U4948 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n4979) );
  INV_X1 U4949 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5673) );
  NOR2_X1 U4950 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4978) );
  NOR2_X1 U4951 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4980) );
  NAND2_X2 U4952 ( .A1(n8133), .A2(n8132), .ZN(n8131) );
  XNOR2_X2 U4953 ( .A(n5388), .B(P1_IR_REG_4__SCAN_IN), .ZN(n10055) );
  OAI21_X2 U4954 ( .B1(n9152), .B2(n6891), .A(n6890), .ZN(n9066) );
  BUF_X2 U4955 ( .A(n4375), .Z(n4287) );
  OAI21_X2 U4956 ( .B1(n5571), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5570) );
  OAI222_X1 U4957 ( .A1(n7143), .A2(P2_U3151), .B1(n9063), .B2(n4287), .C1(
        n5058), .C2(n9062), .ZN(P2_U3294) );
  INV_X2 U4958 ( .A(n9058), .ZN(n9062) );
  AND2_X1 U4959 ( .A1(n6052), .A2(n5654), .ZN(n6048) );
  INV_X1 U4960 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5654) );
  INV_X1 U4961 ( .A(n5859), .ZN(n5871) );
  NAND2_X1 U4962 ( .A1(n9051), .A2(n5647), .ZN(n5761) );
  NOR2_X1 U4963 ( .A1(n5266), .A2(n4618), .ZN(n4617) );
  INV_X1 U4964 ( .A(n5264), .ZN(n4618) );
  AND2_X1 U4965 ( .A1(n5844), .A2(n4996), .ZN(n4995) );
  AND2_X1 U4966 ( .A1(n4992), .A2(n8179), .ZN(n4991) );
  NAND2_X1 U4967 ( .A1(n4993), .A2(n5844), .ZN(n4992) );
  INV_X1 U4968 ( .A(n9051), .ZN(n5648) );
  NAND2_X1 U4969 ( .A1(n7364), .A2(n4643), .ZN(n6308) );
  OR2_X1 U4970 ( .A1(n7016), .A2(n7582), .ZN(n4643) );
  NOR2_X1 U4971 ( .A1(n8962), .A2(n8881), .ZN(n8280) );
  CLKBUF_X1 U4972 ( .A(n6043), .Z(n6044) );
  OR2_X1 U4973 ( .A1(n6113), .A2(n8192), .ZN(n4593) );
  NAND2_X1 U4974 ( .A1(n6113), .A2(n8192), .ZN(n5091) );
  AND4_X1 U4975 ( .A1(n5675), .A2(n5884), .A3(n10361), .A4(n5870), .ZN(n5676)
         );
  INV_X1 U4976 ( .A(n5817), .ZN(n5674) );
  NAND2_X1 U4977 ( .A1(n6722), .A2(n7636), .ZN(n6748) );
  INV_X1 U4978 ( .A(n9996), .ZN(n4726) );
  OR2_X1 U4979 ( .A1(n6586), .A2(n8275), .ZN(n6597) );
  INV_X1 U4980 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5336) );
  OAI21_X1 U4981 ( .B1(n5646), .B2(n4517), .A(n4516), .ZN(n4515) );
  NAND2_X1 U4982 ( .A1(n6070), .A2(n4480), .ZN(n4519) );
  NAND2_X1 U4983 ( .A1(n6069), .A2(n4339), .ZN(n4518) );
  AND2_X2 U4984 ( .A1(n5662), .A2(n5661), .ZN(n5754) );
  NAND2_X1 U4985 ( .A1(n8334), .A2(n6057), .ZN(n8336) );
  AND2_X1 U4986 ( .A1(n5091), .A2(n8499), .ZN(n8394) );
  INV_X1 U4987 ( .A(n8386), .ZN(n4827) );
  AND2_X1 U4988 ( .A1(n5469), .A2(n5457), .ZN(n4880) );
  NAND2_X1 U4989 ( .A1(n6092), .A2(n10156), .ZN(n8341) );
  OAI21_X1 U4990 ( .B1(n4591), .B2(n6115), .A(n4589), .ZN(n4511) );
  AND2_X1 U4991 ( .A1(n4796), .A2(n9352), .ZN(n4794) );
  NAND2_X1 U4992 ( .A1(n9411), .A2(n9342), .ZN(n4799) );
  INV_X1 U4993 ( .A(n5473), .ZN(n5259) );
  OAI21_X1 U4994 ( .B1(n4886), .B2(n5441), .A(n5253), .ZN(n4621) );
  AND2_X1 U4995 ( .A1(n5436), .A2(n5249), .ZN(n4892) );
  NAND2_X1 U4996 ( .A1(n8474), .A2(n4344), .ZN(n4842) );
  INV_X1 U4997 ( .A(n9002), .ZN(n8493) );
  NOR2_X1 U4998 ( .A1(n8757), .A2(n6301), .ZN(n4924) );
  NAND2_X1 U4999 ( .A1(n6300), .A2(n4286), .ZN(n4926) );
  NAND2_X1 U5000 ( .A1(n7243), .A2(n6210), .ZN(n6211) );
  OR2_X1 U5001 ( .A1(n8326), .A2(n6366), .ZN(n8487) );
  AOI21_X1 U5002 ( .B1(n4859), .B2(n4856), .A(n4855), .ZN(n4854) );
  NAND2_X1 U5003 ( .A1(n8908), .A2(n4859), .ZN(n4853) );
  INV_X1 U5004 ( .A(n4328), .ZN(n4856) );
  OR2_X1 U5005 ( .A1(n9031), .A2(n8948), .ZN(n8429) );
  NAND2_X1 U5006 ( .A1(n4507), .A2(n6129), .ZN(n8942) );
  OAI21_X1 U5007 ( .B1(n4533), .B2(n8415), .A(n4354), .ZN(n4507) );
  OR2_X1 U5008 ( .A1(n6101), .A2(n6100), .ZN(n6106) );
  AND2_X1 U5009 ( .A1(n8288), .A2(n6105), .ZN(n5190) );
  NAND2_X1 U5010 ( .A1(n5020), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5680) );
  NAND2_X1 U5011 ( .A1(n5668), .A2(n5667), .ZN(n5708) );
  NAND2_X1 U5012 ( .A1(n6869), .A2(n5125), .ZN(n5124) );
  INV_X1 U5013 ( .A(n9112), .ZN(n5125) );
  INV_X1 U5014 ( .A(n4965), .ZN(n4964) );
  OAI21_X1 U5015 ( .B1(n9626), .B2(n4966), .A(n5032), .ZN(n4965) );
  AND2_X1 U5016 ( .A1(n5043), .A2(n4740), .ZN(n9741) );
  NAND2_X1 U5017 ( .A1(n9783), .A2(n9801), .ZN(n4740) );
  OR2_X1 U5018 ( .A1(n7769), .A2(n7888), .ZN(n9377) );
  NAND2_X1 U5019 ( .A1(n9852), .A2(n10374), .ZN(n5035) );
  NAND2_X1 U5020 ( .A1(n8097), .A2(n4636), .ZN(n9806) );
  OR2_X1 U5021 ( .A1(n9228), .A2(n9835), .ZN(n4636) );
  XNOR2_X1 U5022 ( .A(n5319), .B(n5322), .ZN(n5550) );
  NAND2_X1 U5023 ( .A1(n5321), .A2(n5320), .ZN(n5319) );
  AND3_X1 U5024 ( .A1(n4291), .A2(n4358), .A3(n5182), .ZN(n4807) );
  AND2_X1 U5025 ( .A1(n5338), .A2(n5048), .ZN(n4967) );
  NAND2_X1 U5026 ( .A1(n5300), .A2(n5299), .ZN(n5538) );
  NAND2_X1 U5027 ( .A1(n4608), .A2(n4606), .ZN(n5300) );
  AOI21_X1 U5028 ( .B1(n4609), .B2(n4612), .A(n4607), .ZN(n4606) );
  AND2_X1 U5029 ( .A1(n5305), .A2(n5304), .ZN(n5537) );
  NAND2_X1 U5030 ( .A1(n4615), .A2(n4331), .ZN(n5273) );
  INV_X1 U5031 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U5032 ( .A1(n5458), .A2(n5457), .ZN(n5472) );
  INV_X1 U5033 ( .A(n4882), .ZN(n4560) );
  NAND2_X1 U5034 ( .A1(n5404), .A2(n5224), .ZN(n4583) );
  OR2_X1 U5035 ( .A1(n5843), .A2(n5842), .ZN(n5844) );
  AND2_X1 U5036 ( .A1(n5005), .A2(n5002), .ZN(n5001) );
  NAND2_X1 U5037 ( .A1(n6009), .A2(n5003), .ZN(n5002) );
  NAND2_X1 U5038 ( .A1(n4986), .A2(n4523), .ZN(n4522) );
  INV_X1 U5039 ( .A(n5816), .ZN(n4523) );
  NOR2_X1 U5040 ( .A1(n6045), .A2(n6044), .ZN(n6080) );
  NOR3_X1 U5041 ( .A1(n8501), .A2(n8500), .A3(n8499), .ZN(n8502) );
  AND2_X1 U5042 ( .A1(n4776), .A2(n5060), .ZN(n4558) );
  AND2_X1 U5043 ( .A1(n5910), .A2(n5909), .ZN(n8725) );
  OAI211_X1 U5044 ( .C1(n5691), .C2(n4760), .A(n4759), .B(
        P2_REG1_REG_1__SCAN_IN), .ZN(n4761) );
  OR2_X1 U5045 ( .A1(n4760), .A2(n4385), .ZN(n4759) );
  NAND2_X1 U5046 ( .A1(n4448), .A2(n6301), .ZN(n4908) );
  NAND3_X1 U5047 ( .A1(n4908), .A2(P2_REG2_REG_3__SCAN_IN), .A3(n7169), .ZN(
        n7171) );
  NOR2_X1 U5048 ( .A1(n7154), .A2(n4907), .ZN(n4899) );
  NAND2_X1 U5049 ( .A1(n6308), .A2(n7020), .ZN(n6309) );
  NAND2_X1 U5050 ( .A1(n4933), .A2(n7606), .ZN(n4932) );
  INV_X1 U5051 ( .A(n6216), .ZN(n4441) );
  NAND2_X1 U5052 ( .A1(n4920), .A2(n8796), .ZN(n8798) );
  AND2_X1 U5053 ( .A1(n6218), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4920) );
  NAND2_X1 U5054 ( .A1(n4744), .A2(n4746), .ZN(n4743) );
  NOR2_X1 U5055 ( .A1(n6695), .A2(n6696), .ZN(n6698) );
  NAND2_X1 U5056 ( .A1(n4577), .A2(n5062), .ZN(n8321) );
  AOI21_X1 U5057 ( .B1(n5064), .B2(n5068), .A(n4367), .ZN(n5062) );
  NAND2_X1 U5058 ( .A1(n8878), .A2(n5064), .ZN(n4577) );
  NAND2_X1 U5059 ( .A1(n8231), .A2(n8230), .ZN(n4510) );
  AND2_X1 U5060 ( .A1(n8441), .A2(n4295), .ZN(n8921) );
  INV_X1 U5061 ( .A(n4769), .ZN(n5974) );
  NAND2_X1 U5062 ( .A1(n8011), .A2(n8406), .ZN(n5074) );
  OAI211_X1 U5063 ( .C1(n5754), .C2(n7015), .A(n5759), .B(n5758), .ZN(n7339)
         );
  NAND2_X1 U5064 ( .A1(n6230), .A2(n7010), .ZN(n6081) );
  NAND2_X1 U5065 ( .A1(n5754), .A2(n5663), .ZN(n5757) );
  NAND2_X1 U5066 ( .A1(n5754), .A2(n6990), .ZN(n5773) );
  NAND2_X1 U5067 ( .A1(n4649), .A2(n4328), .ZN(n4857) );
  INV_X1 U5068 ( .A(n8908), .ZN(n4649) );
  OR2_X1 U5069 ( .A1(n8712), .A2(n8947), .ZN(n8422) );
  NAND2_X2 U5070 ( .A1(n5091), .A2(n4593), .ZN(n7721) );
  OR2_X1 U5071 ( .A1(n8475), .A2(n6184), .ZN(n6192) );
  AND2_X1 U5072 ( .A1(n6073), .A2(n10128), .ZN(n6190) );
  INV_X1 U5073 ( .A(n4760), .ZN(n4763) );
  NAND2_X1 U5074 ( .A1(n5691), .A2(n4385), .ZN(n4764) );
  NAND2_X1 U5075 ( .A1(n5871), .A2(n5023), .ZN(n5697) );
  NAND2_X1 U5076 ( .A1(n4292), .A2(n8060), .ZN(n5111) );
  OR2_X1 U5077 ( .A1(n6578), .A2(n9094), .ZN(n6586) );
  NOR2_X1 U5078 ( .A1(n5133), .A2(n5130), .ZN(n5129) );
  INV_X1 U5079 ( .A(n5136), .ZN(n5133) );
  INV_X1 U5080 ( .A(n5134), .ZN(n5130) );
  XNOR2_X1 U5081 ( .A(n6749), .B(n6748), .ZN(n6753) );
  AND2_X1 U5082 ( .A1(n6612), .A2(n6611), .ZN(n8550) );
  OR2_X1 U5083 ( .A1(n8579), .A2(n6615), .ZN(n6612) );
  AND2_X1 U5084 ( .A1(n6595), .A2(n6594), .ZN(n6909) );
  INV_X1 U5085 ( .A(n6588), .ZN(n6615) );
  INV_X1 U5086 ( .A(n10374), .ZN(n9628) );
  NAND2_X1 U5087 ( .A1(n5050), .A2(n5049), .ZN(n9617) );
  AND2_X1 U5088 ( .A1(n5168), .A2(n6659), .ZN(n5049) );
  AOI21_X1 U5089 ( .B1(n9667), .B2(n6657), .A(n6656), .ZN(n9663) );
  INV_X1 U5090 ( .A(n9877), .ZN(n9692) );
  NAND2_X1 U5091 ( .A1(n4631), .A2(n4629), .ZN(n6653) );
  INV_X1 U5092 ( .A(n4630), .ZN(n4629) );
  OR2_X1 U5093 ( .A1(n6484), .A2(n7981), .ZN(n9221) );
  AND2_X1 U5094 ( .A1(n7031), .A2(n8531), .ZN(n9834) );
  NAND2_X1 U5095 ( .A1(n5032), .A2(n5035), .ZN(n5031) );
  AND2_X1 U5096 ( .A1(n5029), .A2(n9306), .ZN(n5028) );
  NAND2_X1 U5097 ( .A1(n5031), .A2(n5034), .ZN(n5029) );
  INV_X1 U5098 ( .A(n5031), .ZN(n5030) );
  OR2_X1 U5099 ( .A1(n7652), .A2(n9349), .ZN(n9864) );
  AND2_X1 U5100 ( .A1(n5040), .A2(n4319), .ZN(n5039) );
  INV_X1 U5101 ( .A(n9795), .ZN(n5040) );
  OAI211_X1 U5102 ( .C1(n4736), .C2(n4732), .A(n4731), .B(n9295), .ZN(n7930)
         );
  INV_X1 U5103 ( .A(n4737), .ZN(n4732) );
  NAND2_X1 U5104 ( .A1(n4729), .A2(n4737), .ZN(n4731) );
  INV_X1 U5105 ( .A(n10107), .ZN(n9930) );
  NAND2_X1 U5106 ( .A1(n8036), .A2(n9366), .ZN(n7652) );
  INV_X1 U5107 ( .A(n9797), .ZN(n9829) );
  XNOR2_X1 U5108 ( .A(n5591), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U5109 ( .A1(n5590), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5591) );
  BUF_X4 U5110 ( .A(n5352), .Z(n5366) );
  AND4_X1 U5111 ( .A1(n5724), .A2(n5723), .A3(n5722), .A4(n5721), .ZN(n7440)
         );
  OR2_X1 U5112 ( .A1(n4283), .A2(n10193), .ZN(n5724) );
  INV_X1 U5113 ( .A(n8334), .ZN(n10154) );
  NAND2_X1 U5114 ( .A1(n6235), .A2(n6234), .ZN(n8846) );
  OR2_X1 U5115 ( .A1(P2_U3150), .A2(n6231), .ZN(n8088) );
  XNOR2_X1 U5116 ( .A(n5598), .B(n5597), .ZN(n8128) );
  AOI21_X1 U5117 ( .B1(n9350), .B2(n9276), .A(n4413), .ZN(n4436) );
  AND2_X2 U5118 ( .A1(n5620), .A2(n9986), .ZN(n10123) );
  NOR2_X1 U5119 ( .A1(n4827), .A2(n4824), .ZN(n4823) );
  INV_X1 U5120 ( .A(n8382), .ZN(n4824) );
  AND2_X1 U5121 ( .A1(n9221), .A2(n9377), .ZN(n4678) );
  INV_X1 U5122 ( .A(n8392), .ZN(n8387) );
  NOR2_X1 U5123 ( .A1(n4828), .A2(n4827), .ZN(n4826) );
  NOR2_X1 U5124 ( .A1(n4299), .A2(n8499), .ZN(n4837) );
  NAND2_X1 U5125 ( .A1(n4370), .A2(n4301), .ZN(n4835) );
  NOR2_X1 U5126 ( .A1(n8420), .A2(n8475), .ZN(n4838) );
  NAND2_X1 U5127 ( .A1(n4462), .A2(n4801), .ZN(n4461) );
  AOI21_X1 U5128 ( .B1(n9234), .B2(n9976), .A(n4802), .ZN(n4801) );
  INV_X1 U5129 ( .A(n4803), .ZN(n4462) );
  NAND2_X1 U5130 ( .A1(n9389), .A2(n9271), .ZN(n4802) );
  NAND2_X1 U5131 ( .A1(n4681), .A2(n4679), .ZN(n9229) );
  NOR2_X1 U5132 ( .A1(n9230), .A2(n4680), .ZN(n4679) );
  INV_X1 U5133 ( .A(n4837), .ZN(n4831) );
  NAND2_X1 U5134 ( .A1(n5188), .A2(n8414), .ZN(n8416) );
  AOI21_X1 U5135 ( .B1(n4561), .B2(n8413), .A(n8418), .ZN(n5188) );
  INV_X1 U5136 ( .A(n4835), .ZN(n4830) );
  INV_X1 U5137 ( .A(n8465), .ZN(n4541) );
  AND2_X1 U5138 ( .A1(n4976), .A2(n5187), .ZN(n9260) );
  AND2_X1 U5139 ( .A1(n7460), .A2(n8365), .ZN(n8355) );
  INV_X1 U5140 ( .A(n8347), .ZN(n6170) );
  INV_X1 U5141 ( .A(n8348), .ZN(n4694) );
  INV_X1 U5142 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n4775) );
  NAND2_X1 U5143 ( .A1(n6091), .A2(n6093), .ZN(n8340) );
  AOI21_X1 U5144 ( .B1(n4360), .B2(n5694), .A(n5179), .ZN(n6043) );
  NOR2_X1 U5145 ( .A1(n8887), .A2(n4860), .ZN(n4859) );
  INV_X1 U5146 ( .A(n4869), .ZN(n4800) );
  OAI211_X1 U5147 ( .C1(n9269), .C2(n9352), .A(n4871), .B(n4870), .ZN(n4869)
         );
  OR2_X1 U5148 ( .A1(n9420), .A2(n9271), .ZN(n4870) );
  NAND2_X1 U5149 ( .A1(n9269), .A2(n9420), .ZN(n4871) );
  AND2_X1 U5150 ( .A1(n9274), .A2(n9419), .ZN(n4798) );
  INV_X1 U5151 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5565) );
  OAI21_X1 U5152 ( .B1(n5366), .B2(n4699), .A(n4698), .ZN(n5225) );
  NAND2_X1 U5153 ( .A1(n5366), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n4698) );
  AND2_X1 U5154 ( .A1(n6006), .A2(n8624), .ZN(n6026) );
  INV_X2 U5155 ( .A(n6339), .ZN(n5903) );
  AND2_X1 U5156 ( .A1(n6334), .A2(n6025), .ZN(n4703) );
  NOR2_X1 U5157 ( .A1(n8493), .A2(n8279), .ZN(n8488) );
  AND3_X1 U5158 ( .A1(n8508), .A2(n4378), .A3(n4655), .ZN(n4654) );
  NAND2_X1 U5159 ( .A1(n8319), .A2(n8999), .ZN(n4655) );
  NOR2_X1 U5160 ( .A1(n7181), .A2(n10193), .ZN(n4674) );
  NAND2_X1 U5161 ( .A1(n6303), .A2(n6302), .ZN(n4948) );
  AND2_X1 U5162 ( .A1(n4906), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4903) );
  NAND3_X1 U5163 ( .A1(n4937), .A2(P2_REG1_REG_7__SCAN_IN), .A3(n6307), .ZN(
        n4936) );
  NAND2_X1 U5164 ( .A1(n4420), .A2(n4419), .ZN(n6316) );
  AOI21_X1 U5165 ( .B1(n7963), .B2(n7962), .A(n4397), .ZN(n4419) );
  NAND2_X1 U5166 ( .A1(n7961), .A2(n7962), .ZN(n4420) );
  OAI211_X1 U5167 ( .C1(n4942), .C2(n4941), .A(n4940), .B(n4406), .ZN(n6321)
         );
  AND2_X1 U5168 ( .A1(n4303), .A2(n4912), .ZN(n6221) );
  INV_X1 U5169 ( .A(n8280), .ZN(n8471) );
  AND2_X1 U5170 ( .A1(n5635), .A2(n4785), .ZN(n4784) );
  INV_X1 U5171 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n4785) );
  INV_X1 U5172 ( .A(n6014), .ZN(n5636) );
  INV_X1 U5173 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n4782) );
  INV_X1 U5174 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5632) );
  INV_X1 U5175 ( .A(n5915), .ZN(n5633) );
  INV_X1 U5176 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n4779) );
  INV_X1 U5177 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5630) );
  INV_X1 U5178 ( .A(n5861), .ZN(n5631) );
  NAND2_X1 U5179 ( .A1(n8369), .A2(n7696), .ZN(n6176) );
  NAND2_X1 U5180 ( .A1(n7383), .A2(n6097), .ZN(n7436) );
  NAND2_X1 U5181 ( .A1(n7353), .A2(n7484), .ZN(n8354) );
  INV_X1 U5182 ( .A(n10156), .ZN(n6093) );
  AND2_X1 U5183 ( .A1(n8429), .A2(n8428), .ZN(n8302) );
  NOR2_X1 U5184 ( .A1(n8221), .A2(n5076), .ZN(n5075) );
  INV_X1 U5185 ( .A(n8421), .ZN(n5076) );
  NAND2_X1 U5186 ( .A1(n8157), .A2(n6126), .ZN(n4533) );
  CLKBUF_X1 U5187 ( .A(n8021), .Z(n8022) );
  INV_X1 U5188 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5900) );
  INV_X1 U5189 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5884) );
  INV_X1 U5190 ( .A(n5708), .ZN(n5707) );
  NOR2_X1 U5191 ( .A1(n9306), .A2(n9305), .ZN(n4668) );
  INV_X1 U5192 ( .A(SI_18_), .ZN(n10300) );
  OR2_X1 U5193 ( .A1(n9855), .A2(n6909), .ZN(n9311) );
  NOR2_X1 U5194 ( .A1(n9947), .A2(n9660), .ZN(n5151) );
  OAI21_X1 U5195 ( .B1(n9721), .B2(n9729), .A(n9706), .ZN(n4630) );
  NAND2_X1 U5196 ( .A1(n9704), .A2(n5184), .ZN(n4631) );
  NAND2_X1 U5197 ( .A1(n4955), .A2(n9249), .ZN(n4954) );
  NAND2_X1 U5198 ( .A1(n4958), .A2(n9725), .ZN(n4955) );
  NAND2_X1 U5199 ( .A1(n4959), .A2(n4961), .ZN(n4958) );
  NOR2_X1 U5200 ( .A1(n4956), .A2(n4719), .ZN(n4718) );
  INV_X1 U5201 ( .A(n4720), .ZN(n4719) );
  NAND2_X1 U5202 ( .A1(n9249), .A2(n4959), .ZN(n4956) );
  AND2_X1 U5203 ( .A1(n9765), .A2(n9243), .ZN(n4720) );
  AND2_X1 U5204 ( .A1(n5158), .A2(n9783), .ZN(n5157) );
  NOR2_X1 U5205 ( .A1(n9911), .A2(n9820), .ZN(n5158) );
  NOR2_X2 U5206 ( .A1(n9840), .A2(n9924), .ZN(n9817) );
  NAND2_X1 U5207 ( .A1(n10101), .A2(n9428), .ZN(n9367) );
  NAND2_X1 U5208 ( .A1(n7647), .A2(n7900), .ZN(n9195) );
  INV_X1 U5209 ( .A(n9344), .ZN(n7031) );
  OR2_X1 U5210 ( .A1(n9269), .A2(n9270), .ZN(n9337) );
  NAND2_X1 U5211 ( .A1(n9625), .A2(n9626), .ZN(n9624) );
  OR2_X1 U5212 ( .A1(n9955), .A2(n9729), .ZN(n9250) );
  OR2_X1 U5213 ( .A1(n9911), .A2(n9180), .ZN(n9389) );
  NAND2_X1 U5214 ( .A1(n5543), .A2(n5314), .ZN(n5321) );
  INV_X1 U5215 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5345) );
  AND2_X1 U5216 ( .A1(n5299), .A2(n5298), .ZN(n5533) );
  AND4_X1 U5217 ( .A1(n5332), .A2(n5331), .A3(n10339), .A4(n5410), .ZN(n4291)
         );
  NOR2_X1 U5218 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5331) );
  AND2_X1 U5219 ( .A1(n5294), .A2(n5293), .ZN(n5529) );
  NOR2_X1 U5220 ( .A1(n5513), .A2(n4894), .ZN(n4893) );
  INV_X1 U5221 ( .A(n5279), .ZN(n4894) );
  INV_X1 U5222 ( .A(SI_20_), .ZN(n5504) );
  OAI21_X1 U5223 ( .B1(n5505), .B2(n5504), .A(n5503), .ZN(n5507) );
  INV_X1 U5224 ( .A(SI_19_), .ZN(n5267) );
  AOI21_X1 U5225 ( .B1(n4617), .B2(n5480), .A(n4359), .ZN(n4616) );
  NAND2_X1 U5226 ( .A1(n5261), .A2(n10264), .ZN(n5264) );
  AOI21_X1 U5227 ( .B1(n4878), .B2(n4879), .A(n4363), .ZN(n4876) );
  AOI21_X1 U5228 ( .B1(n4890), .B2(n4888), .A(n4887), .ZN(n4886) );
  INV_X1 U5229 ( .A(n5243), .ZN(n4888) );
  NAND2_X1 U5230 ( .A1(n4646), .A2(n4350), .ZN(n4887) );
  NAND2_X1 U5231 ( .A1(n5415), .A2(n4595), .ZN(n4594) );
  NOR2_X1 U5232 ( .A1(n5244), .A2(n4596), .ZN(n4595) );
  INV_X1 U5233 ( .A(n5239), .ZN(n4596) );
  NAND2_X1 U5234 ( .A1(n5415), .A2(n5239), .ZN(n5421) );
  INV_X1 U5235 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5410) );
  INV_X1 U5236 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4600) );
  OR2_X1 U5237 ( .A1(n9064), .A2(n6296), .ZN(n6072) );
  NAND2_X1 U5238 ( .A1(n8680), .A2(n4390), .ZN(n4476) );
  NAND2_X1 U5239 ( .A1(n7920), .A2(n7919), .ZN(n4470) );
  AOI22_X1 U5240 ( .A1(n4991), .A2(n4994), .B1(n4989), .B2(n4990), .ZN(n4985)
         );
  INV_X1 U5241 ( .A(n5844), .ZN(n4994) );
  INV_X1 U5242 ( .A(n4995), .ZN(n4990) );
  INV_X1 U5243 ( .A(n4989), .ZN(n4988) );
  INV_X1 U5244 ( .A(n4991), .ZN(n4987) );
  XNOR2_X1 U5245 ( .A(n5760), .B(n10156), .ZN(n5752) );
  OR2_X1 U5246 ( .A1(n8592), .A2(n8591), .ZN(n5019) );
  AND4_X1 U5247 ( .A1(n5642), .A2(n5641), .A3(n5683), .A4(n5640), .ZN(n5643)
         );
  INV_X1 U5248 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5640) );
  AND3_X1 U5249 ( .A1(n5893), .A2(n5892), .A3(n5891), .ZN(n8023) );
  AND3_X1 U5250 ( .A1(n5881), .A2(n5880), .A3(n5879), .ZN(n8669) );
  OR2_X1 U5251 ( .A1(n5742), .A2(n5741), .ZN(n5745) );
  NAND2_X1 U5252 ( .A1(n4281), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n4478) );
  AND2_X1 U5253 ( .A1(n5751), .A2(n5750), .ZN(n4535) );
  NAND2_X1 U5254 ( .A1(n8312), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4479) );
  OAI211_X1 U5255 ( .C1(n8755), .C2(n4923), .A(n4926), .B(n4925), .ZN(n4922)
         );
  INV_X1 U5256 ( .A(n6300), .ZN(n4927) );
  NAND2_X1 U5257 ( .A1(n8767), .A2(n4491), .ZN(n7096) );
  AND2_X1 U5258 ( .A1(n4492), .A2(n6240), .ZN(n4491) );
  NAND2_X1 U5259 ( .A1(n4464), .A2(n4463), .ZN(n5735) );
  NAND2_X1 U5260 ( .A1(n7171), .A2(n7169), .ZN(n6208) );
  NAND2_X1 U5261 ( .A1(n7184), .A2(n4489), .ZN(n4749) );
  NOR2_X1 U5262 ( .A1(n4752), .A2(n4490), .ZN(n4489) );
  INV_X1 U5263 ( .A(n7183), .ZN(n4490) );
  INV_X1 U5264 ( .A(n7164), .ZN(n4752) );
  NAND2_X1 U5265 ( .A1(n4749), .A2(n4747), .ZN(n7231) );
  NOR2_X1 U5266 ( .A1(n4748), .A2(n7234), .ZN(n4747) );
  INV_X1 U5267 ( .A(n4750), .ZN(n4748) );
  NAND2_X1 U5268 ( .A1(n4935), .A2(n7365), .ZN(n7364) );
  NAND2_X1 U5269 ( .A1(n4936), .A2(n6307), .ZN(n4935) );
  NAND2_X1 U5270 ( .A1(n4446), .A2(n7020), .ZN(n7560) );
  NAND2_X1 U5271 ( .A1(n7376), .A2(n6213), .ZN(n4446) );
  AND2_X1 U5272 ( .A1(n4308), .A2(n4932), .ZN(n7608) );
  INV_X1 U5273 ( .A(n6260), .ZN(n4485) );
  INV_X1 U5274 ( .A(n8774), .ZN(n4746) );
  NOR2_X1 U5275 ( .A1(n4708), .A2(n6220), .ZN(n8811) );
  AND2_X1 U5276 ( .A1(n6219), .A2(n6320), .ZN(n4708) );
  NAND2_X1 U5277 ( .A1(n4424), .A2(n6320), .ZN(n4423) );
  INV_X1 U5278 ( .A(n6321), .ZN(n4424) );
  NAND2_X1 U5279 ( .A1(n4423), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4422) );
  NAND2_X1 U5280 ( .A1(n6321), .A2(n8815), .ZN(n4425) );
  NAND2_X1 U5281 ( .A1(n8806), .A2(n8807), .ZN(n6280) );
  NAND2_X1 U5282 ( .A1(n8822), .A2(n4928), .ZN(n4432) );
  NAND2_X1 U5283 ( .A1(n4929), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4928) );
  NAND2_X1 U5284 ( .A1(n4432), .A2(n8845), .ZN(n6684) );
  NAND2_X1 U5285 ( .A1(n6151), .A2(n6150), .ZN(n8326) );
  AOI21_X1 U5286 ( .B1(n5067), .B2(n5066), .A(n5065), .ZN(n5064) );
  INV_X1 U5287 ( .A(n5070), .ZN(n5066) );
  NAND2_X1 U5288 ( .A1(n5072), .A2(n8468), .ZN(n5069) );
  NOR2_X1 U5289 ( .A1(n8280), .A2(n5071), .ZN(n5070) );
  INV_X1 U5290 ( .A(n8468), .ZN(n5071) );
  INV_X1 U5291 ( .A(n4318), .ZN(n5072) );
  AND2_X1 U5292 ( .A1(n8471), .A2(n8472), .ZN(n8870) );
  NAND2_X1 U5293 ( .A1(n8891), .A2(n10132), .ZN(n8866) );
  NAND2_X1 U5294 ( .A1(n5636), .A2(n4784), .ZN(n6062) );
  INV_X1 U5295 ( .A(n8438), .ZN(n5090) );
  OR2_X1 U5296 ( .A1(n5940), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5942) );
  NAND2_X1 U5297 ( .A1(n6181), .A2(n4345), .ZN(n5077) );
  AND2_X1 U5298 ( .A1(n5921), .A2(n5920), .ZN(n8708) );
  OR2_X1 U5299 ( .A1(n5904), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U5300 ( .A1(n8016), .A2(n8594), .ZN(n8405) );
  AND2_X1 U5301 ( .A1(n8407), .A2(n8405), .ZN(n5073) );
  NAND2_X1 U5302 ( .A1(n5628), .A2(n10238), .ZN(n5829) );
  INV_X1 U5303 ( .A(n5808), .ZN(n5628) );
  NAND2_X1 U5304 ( .A1(n4766), .A2(n4765), .ZN(n5808) );
  INV_X1 U5305 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n4765) );
  INV_X1 U5306 ( .A(n5797), .ZN(n4766) );
  AND4_X1 U5307 ( .A1(n5718), .A2(n5717), .A3(n5716), .A4(n5715), .ZN(n7474)
         );
  NOR2_X1 U5308 ( .A1(n8500), .A2(n7677), .ZN(n7304) );
  OR2_X1 U5309 ( .A1(n10172), .A2(n8338), .ZN(n6353) );
  AND2_X1 U5310 ( .A1(n8335), .A2(n10154), .ZN(n7299) );
  AND3_X1 U5311 ( .A1(n6360), .A2(n6359), .A3(n6358), .ZN(n7302) );
  NAND2_X1 U5312 ( .A1(n6033), .A2(n7008), .ZN(n7300) );
  AND2_X1 U5313 ( .A1(n4579), .A2(n8446), .ZN(n4578) );
  INV_X1 U5314 ( .A(n4313), .ZN(n5084) );
  AND2_X1 U5315 ( .A1(n8446), .A2(n8445), .ZN(n8903) );
  AND2_X1 U5316 ( .A1(n6022), .A2(n6021), .ZN(n8899) );
  INV_X1 U5317 ( .A(n4509), .ZN(n4508) );
  OAI21_X1 U5318 ( .B1(n4321), .B2(n8921), .A(n4677), .ZN(n4509) );
  OR2_X1 U5319 ( .A1(n8675), .A2(n8910), .ZN(n4677) );
  AOI21_X1 U5320 ( .B1(n5090), .B2(n4295), .A(n5089), .ZN(n5088) );
  AND2_X1 U5321 ( .A1(n4323), .A2(n8442), .ZN(n8909) );
  NAND2_X1 U5322 ( .A1(n4850), .A2(n4849), .ZN(n8231) );
  AOI21_X1 U5323 ( .B1(n4851), .B2(n8941), .A(n4362), .ZN(n4849) );
  NAND2_X1 U5324 ( .A1(n8930), .A2(n8429), .ZN(n8228) );
  AND2_X1 U5325 ( .A1(n8932), .A2(n4374), .ZN(n4851) );
  OR2_X1 U5326 ( .A1(n8942), .A2(n8941), .ZN(n4852) );
  OAI21_X1 U5327 ( .B1(n5077), .B2(n4573), .A(n4571), .ZN(n8930) );
  INV_X1 U5328 ( .A(n4572), .ZN(n4571) );
  OAI21_X1 U5329 ( .B1(n5075), .B2(n4573), .A(n8425), .ZN(n4572) );
  NAND2_X1 U5330 ( .A1(n8422), .A2(n4343), .ZN(n4573) );
  INV_X1 U5331 ( .A(n8302), .ZN(n8932) );
  AND2_X1 U5332 ( .A1(n5965), .A2(n5964), .ZN(n8947) );
  INV_X1 U5333 ( .A(n8608), .ZN(n8941) );
  NAND2_X1 U5334 ( .A1(n5077), .A2(n5075), .ZN(n8224) );
  OR2_X1 U5335 ( .A1(n8634), .A2(n8725), .ZN(n8419) );
  NAND2_X1 U5336 ( .A1(n8156), .A2(n8417), .ZN(n6181) );
  NAND2_X1 U5337 ( .A1(n4570), .A2(n8330), .ZN(n8156) );
  OAI21_X1 U5338 ( .B1(n5074), .B2(n4569), .A(n4567), .ZN(n4570) );
  AND2_X1 U5339 ( .A1(n4568), .A2(n8329), .ZN(n4567) );
  OR2_X1 U5340 ( .A1(n5073), .A2(n4569), .ZN(n4568) );
  OR2_X1 U5341 ( .A1(n8022), .A2(n8407), .ZN(n8025) );
  INV_X1 U5342 ( .A(n6114), .ZN(n4587) );
  OR2_X1 U5343 ( .A1(n8185), .A2(n8745), .ZN(n6116) );
  AOI21_X1 U5344 ( .B1(n7862), .B2(n8399), .A(n6180), .ZN(n8011) );
  AND2_X1 U5345 ( .A1(n7721), .A2(n6110), .ZN(n6111) );
  INV_X1 U5346 ( .A(n6109), .ZN(n6110) );
  INV_X1 U5347 ( .A(n8946), .ZN(n10132) );
  NAND2_X1 U5348 ( .A1(n7517), .A2(n5095), .ZN(n5094) );
  NOR2_X1 U5349 ( .A1(n8383), .A2(n5096), .ZN(n5095) );
  NAND2_X1 U5350 ( .A1(n6160), .A2(n8499), .ZN(n8946) );
  AND3_X1 U5351 ( .A1(n5778), .A2(n5777), .A3(n5776), .ZN(n10171) );
  XNOR2_X1 U5352 ( .A(n6051), .B(n6050), .ZN(n6229) );
  AND2_X1 U5353 ( .A1(n5645), .A2(n5646), .ZN(n5644) );
  NAND2_X1 U5354 ( .A1(n4843), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4504) );
  OAI22_X1 U5355 ( .A1(n5644), .A2(n4504), .B1(P2_IR_REG_31__SCAN_IN), .B2(
        n4843), .ZN(n4501) );
  INV_X1 U5356 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U5357 ( .A1(n5686), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5687) );
  NAND2_X1 U5358 ( .A1(n6048), .A2(n6050), .ZN(n5055) );
  NAND2_X1 U5359 ( .A1(n4526), .A2(n4524), .ZN(n5686) );
  INV_X1 U5360 ( .A(n4525), .ZN(n4524) );
  OR2_X1 U5361 ( .A1(n6048), .A2(n4520), .ZN(n4526) );
  OAI21_X1 U5362 ( .B1(n6050), .B2(n4520), .A(n5683), .ZN(n4525) );
  INV_X1 U5363 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5683) );
  AND2_X1 U5364 ( .A1(n5023), .A2(n5022), .ZN(n5021) );
  NAND2_X1 U5365 ( .A1(n4811), .A2(n4464), .ZN(n5825) );
  XNOR2_X1 U5366 ( .A(n5709), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6304) );
  NAND2_X1 U5367 ( .A1(n6390), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6478) );
  INV_X1 U5368 ( .A(n6472), .ZN(n6390) );
  NAND2_X1 U5369 ( .A1(n9162), .A2(n5127), .ZN(n5121) );
  AND2_X1 U5370 ( .A1(n6926), .A2(n6925), .ZN(n6928) );
  AND2_X1 U5371 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n6387) );
  NAND2_X1 U5372 ( .A1(n4687), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6487) );
  INV_X1 U5373 ( .A(n6478), .ZN(n4687) );
  NAND2_X1 U5374 ( .A1(n6569), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6578) );
  INV_X1 U5375 ( .A(n6571), .ZN(n6569) );
  XNOR2_X1 U5376 ( .A(n6760), .B(n8547), .ZN(n6761) );
  NAND2_X1 U5377 ( .A1(n6759), .A2(n6758), .ZN(n6760) );
  NAND2_X1 U5378 ( .A1(n4685), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n6472) );
  INV_X1 U5379 ( .A(n6463), .ZN(n4685) );
  AND2_X1 U5380 ( .A1(n6736), .A2(n6738), .ZN(n5097) );
  INV_X1 U5381 ( .A(n8042), .ZN(n5108) );
  AND2_X1 U5382 ( .A1(n8060), .A2(n6823), .ZN(n5110) );
  OR2_X1 U5383 ( .A1(n6829), .A2(n7978), .ZN(n6823) );
  NAND2_X1 U5384 ( .A1(n9074), .A2(n9075), .ZN(n9073) );
  NAND2_X1 U5385 ( .A1(n5138), .A2(n5137), .ZN(n5136) );
  INV_X1 U5386 ( .A(n5127), .ZN(n5117) );
  NAND2_X1 U5387 ( .A1(n5126), .A2(n5127), .ZN(n5116) );
  NAND2_X1 U5388 ( .A1(n5124), .A2(n5127), .ZN(n5115) );
  OR2_X1 U5389 ( .A1(n5126), .A2(n5124), .ZN(n5118) );
  OR2_X1 U5390 ( .A1(n7266), .A2(n8531), .ZN(n8264) );
  AND2_X1 U5391 ( .A1(n9985), .A2(n6940), .ZN(n6936) );
  OAI21_X1 U5392 ( .B1(n4792), .B2(n4872), .A(n4787), .ZN(n9350) );
  NAND2_X1 U5393 ( .A1(n9988), .A2(n5560), .ZN(n4625) );
  NAND2_X1 U5394 ( .A1(n6961), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6427) );
  NOR2_X2 U5395 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5024) );
  NOR2_X1 U5396 ( .A1(n5408), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5424) );
  AOI21_X1 U5397 ( .B1(n7132), .B2(n7131), .A(n7130), .ZN(n7134) );
  NOR2_X1 U5398 ( .A1(n7211), .A2(n4393), .ZN(n7189) );
  AND2_X1 U5399 ( .A1(n5452), .A2(n5451), .ZN(n5462) );
  XNOR2_X1 U5400 ( .A(n9534), .B(n4701), .ZN(n7686) );
  INV_X1 U5401 ( .A(n9533), .ZN(n4701) );
  NAND2_X1 U5402 ( .A1(n9550), .A2(n4394), .ZN(n9555) );
  NOR2_X1 U5403 ( .A1(n9555), .A2(n9554), .ZN(n9569) );
  AND2_X1 U5404 ( .A1(n5423), .A2(n5144), .ZN(n5143) );
  NOR2_X1 U5405 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5423) );
  NOR2_X1 U5406 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5333) );
  NOR2_X1 U5407 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5334) );
  AOI21_X1 U5408 ( .B1(n4962), .B2(n4297), .A(n4688), .ZN(n6958) );
  OAI21_X1 U5409 ( .B1(n4964), .B2(n4963), .A(n9336), .ZN(n4688) );
  INV_X1 U5410 ( .A(n9625), .ZN(n4962) );
  NAND2_X1 U5411 ( .A1(n9624), .A2(n9322), .ZN(n6705) );
  NAND2_X1 U5412 ( .A1(n9421), .A2(n9834), .ZN(n6707) );
  AND2_X1 U5413 ( .A1(n9311), .A2(n9322), .ZN(n9626) );
  AOI21_X1 U5414 ( .B1(n4974), .B2(n9669), .A(n4972), .ZN(n4971) );
  INV_X1 U5415 ( .A(n9316), .ZN(n4972) );
  INV_X1 U5416 ( .A(n4975), .ZN(n4974) );
  NAND2_X1 U5417 ( .A1(n9685), .A2(n4968), .ZN(n4970) );
  NOR2_X1 U5418 ( .A1(n4975), .A2(n4969), .ZN(n4968) );
  INV_X1 U5419 ( .A(n9670), .ZN(n4969) );
  NAND2_X1 U5420 ( .A1(n4970), .A2(n4574), .ZN(n9634) );
  AND2_X1 U5421 ( .A1(n4971), .A2(n9636), .ZN(n4574) );
  AND2_X1 U5422 ( .A1(n9301), .A2(n4973), .ZN(n9668) );
  NAND2_X1 U5423 ( .A1(n9685), .A2(n9670), .ZN(n4973) );
  AND2_X2 U5424 ( .A1(n9717), .A2(n9692), .ZN(n9693) );
  INV_X1 U5425 ( .A(n6537), .ZN(n6535) );
  AND2_X1 U5426 ( .A1(n6533), .A2(n6532), .ZN(n9728) );
  AND2_X1 U5427 ( .A1(n9395), .A2(n9401), .ZN(n9750) );
  NAND2_X1 U5428 ( .A1(n9775), .A2(n4720), .ZN(n9764) );
  AND2_X1 U5429 ( .A1(n9396), .A2(n9244), .ZN(n9765) );
  NAND2_X1 U5430 ( .A1(n6505), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6513) );
  INV_X1 U5431 ( .A(n6507), .ZN(n6505) );
  AND3_X1 U5432 ( .A1(n6517), .A2(n6516), .A3(n6515), .ZN(n9801) );
  AND4_X1 U5433 ( .A1(n6405), .A2(n6404), .A3(n6403), .A4(n6402), .ZN(n9807)
         );
  AND2_X1 U5434 ( .A1(n9387), .A2(n9232), .ZN(n9812) );
  NAND2_X1 U5435 ( .A1(n7111), .A2(n5560), .ZN(n5440) );
  AND2_X1 U5436 ( .A1(n9224), .A2(n9380), .ZN(n7934) );
  AND3_X1 U5437 ( .A1(n4565), .A2(n9293), .A3(n9220), .ZN(n4564) );
  NAND2_X1 U5438 ( .A1(n4733), .A2(n4736), .ZN(n7771) );
  NOR2_X1 U5439 ( .A1(n5178), .A2(n4734), .ZN(n4733) );
  INV_X1 U5440 ( .A(n6641), .ZN(n4734) );
  NAND2_X1 U5441 ( .A1(n7771), .A2(n9278), .ZN(n7770) );
  NAND2_X1 U5442 ( .A1(n7748), .A2(n6638), .ZN(n7988) );
  INV_X1 U5443 ( .A(n9281), .ZN(n7903) );
  NAND2_X1 U5444 ( .A1(n9367), .A2(n9195), .ZN(n9281) );
  INV_X1 U5445 ( .A(n9834), .ZN(n9802) );
  AND2_X1 U5446 ( .A1(n9275), .A2(n9353), .ZN(n9797) );
  AND2_X1 U5447 ( .A1(n9319), .A2(n9262), .ZN(n9636) );
  AOI21_X1 U5448 ( .B1(n9691), .B2(n6655), .A(n6654), .ZN(n9667) );
  NOR2_X1 U5449 ( .A1(n9877), .A2(n9714), .ZN(n6654) );
  OAI21_X1 U5450 ( .B1(n9806), .B2(n5038), .A(n5036), .ZN(n5043) );
  AOI21_X1 U5451 ( .B1(n5039), .B2(n5037), .A(n4369), .ZN(n5036) );
  INV_X1 U5452 ( .A(n5039), .ZN(n5038) );
  NAND2_X1 U5453 ( .A1(n4312), .A2(n9808), .ZN(n5042) );
  NAND2_X1 U5454 ( .A1(n9806), .A2(n4312), .ZN(n5041) );
  AND2_X1 U5455 ( .A1(n9389), .A2(n9233), .ZN(n9795) );
  NAND2_X1 U5456 ( .A1(n5045), .A2(n5047), .ZN(n4737) );
  INV_X1 U5457 ( .A(n7934), .ZN(n9295) );
  NAND2_X1 U5458 ( .A1(n4738), .A2(n4300), .ZN(n4729) );
  NOR2_X1 U5459 ( .A1(n7631), .A2(n5614), .ZN(n5620) );
  OR2_X1 U5460 ( .A1(n7635), .A2(n6934), .ZN(n5614) );
  NAND2_X1 U5461 ( .A1(n5345), .A2(n5339), .ZN(n5340) );
  INV_X1 U5462 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5339) );
  XNOR2_X1 U5463 ( .A(n5534), .B(n5533), .ZN(n8171) );
  NAND2_X1 U5464 ( .A1(n4605), .A2(n4609), .ZN(n5534) );
  OR2_X1 U5465 ( .A1(n5518), .A2(n4612), .ZN(n4605) );
  NAND2_X1 U5466 ( .A1(n4895), .A2(n5279), .ZN(n5514) );
  NAND2_X1 U5467 ( .A1(n5273), .A2(n5272), .ZN(n5505) );
  NAND2_X1 U5468 ( .A1(n5571), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5572) );
  XNOR2_X1 U5469 ( .A(n4725), .B(n5436), .ZN(n7111) );
  OAI21_X1 U5470 ( .B1(n5430), .B2(n5429), .A(n5249), .ZN(n4725) );
  NAND2_X1 U5471 ( .A1(n5142), .A2(n5143), .ZN(n5482) );
  OR2_X1 U5472 ( .A1(n5482), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5432) );
  AOI21_X1 U5473 ( .B1(n4583), .B2(n4885), .A(n4884), .ZN(n4883) );
  NAND2_X1 U5474 ( .A1(n6137), .A2(n6136), .ZN(n8962) );
  NAND2_X1 U5475 ( .A1(n5874), .A2(n5873), .ZN(n8597) );
  NOR2_X1 U5476 ( .A1(n8602), .A2(n8738), .ZN(n8649) );
  NAND2_X1 U5477 ( .A1(n4472), .A2(n4476), .ZN(n8602) );
  INV_X1 U5478 ( .A(n4473), .ZN(n4472) );
  AOI21_X1 U5479 ( .B1(n8680), .B2(n5986), .A(n8601), .ZN(n4473) );
  AND4_X1 U5480 ( .A1(n5824), .A2(n5823), .A3(n5822), .A4(n5821), .ZN(n8192)
         );
  OR2_X1 U5481 ( .A1(n5761), .A2(n10147), .ZN(n5764) );
  AND2_X1 U5482 ( .A1(n5980), .A2(n5979), .ZN(n8255) );
  NAND2_X1 U5483 ( .A1(n4529), .A2(n4528), .ZN(n4527) );
  INV_X1 U5484 ( .A(n8678), .ZN(n4528) );
  OAI21_X1 U5485 ( .B1(n8656), .B2(n4389), .A(n4530), .ZN(n4529) );
  NAND2_X1 U5486 ( .A1(n5772), .A2(n7440), .ZN(n5015) );
  OR2_X1 U5487 ( .A1(n7349), .A2(n7350), .ZN(n5016) );
  NAND2_X1 U5488 ( .A1(n4482), .A2(n4481), .ZN(n8639) );
  NAND2_X1 U5489 ( .A1(n8630), .A2(n8628), .ZN(n4481) );
  OAI21_X1 U5490 ( .B1(n8630), .B2(n8628), .A(n8741), .ZN(n4482) );
  AND2_X1 U5491 ( .A1(n5995), .A2(n5994), .ZN(n8920) );
  NAND2_X1 U5492 ( .A1(n4470), .A2(n4469), .ZN(n8051) );
  AND2_X1 U5493 ( .A1(n4320), .A2(n8052), .ZN(n4469) );
  INV_X1 U5494 ( .A(n8707), .ZN(n8722) );
  AND2_X1 U5495 ( .A1(n5929), .A2(n5928), .ZN(n8919) );
  NAND2_X1 U5496 ( .A1(n5957), .A2(n5956), .ZN(n8712) );
  OR3_X1 U5497 ( .A1(n6189), .A2(n6160), .A3(n6192), .ZN(n8724) );
  NAND2_X1 U5498 ( .A1(n6084), .A2(n6083), .ZN(n8727) );
  NAND2_X1 U5499 ( .A1(n8481), .A2(n4550), .ZN(n4549) );
  XNOR2_X1 U5500 ( .A(n6054), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8513) );
  INV_X1 U5501 ( .A(n8919), .ZN(n8934) );
  NAND2_X1 U5502 ( .A1(n5939), .A2(n5938), .ZN(n8933) );
  INV_X1 U5503 ( .A(n8725), .ZN(n8741) );
  INV_X1 U5504 ( .A(n8023), .ZN(n8743) );
  INV_X1 U5505 ( .A(n8669), .ZN(n8744) );
  INV_X1 U5506 ( .A(n8192), .ZN(n8746) );
  NAND2_X1 U5507 ( .A1(n7150), .A2(n6238), .ZN(n8769) );
  NAND2_X1 U5508 ( .A1(n8769), .A2(n8768), .ZN(n8767) );
  NAND2_X1 U5509 ( .A1(n4908), .A2(n7169), .ZN(n7105) );
  NAND2_X1 U5510 ( .A1(n7182), .A2(n6245), .ZN(n7165) );
  NAND2_X1 U5511 ( .A1(n8083), .A2(n8084), .ZN(n6267) );
  AND2_X1 U5512 ( .A1(n8796), .A2(n6218), .ZN(n8775) );
  NAND2_X1 U5513 ( .A1(n6324), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8837) );
  INV_X1 U5514 ( .A(n8839), .ZN(n6324) );
  INV_X1 U5515 ( .A(n8825), .ZN(n8856) );
  OR2_X1 U5516 ( .A1(n6699), .A2(n7497), .ZN(n4494) );
  OAI21_X1 U5517 ( .B1(n6698), .B2(n8850), .A(n7497), .ZN(n4493) );
  NAND2_X1 U5518 ( .A1(n4707), .A2(n8853), .ZN(n6703) );
  NAND2_X1 U5519 ( .A1(n6692), .A2(n6693), .ZN(n4707) );
  AND2_X1 U5520 ( .A1(n7253), .A2(n9064), .ZN(n8825) );
  XNOR2_X1 U5521 ( .A(n4758), .B(n4757), .ZN(n4756) );
  INV_X1 U5522 ( .A(n6295), .ZN(n4757) );
  AOI21_X1 U5523 ( .B1(n6694), .B2(n7497), .A(n6696), .ZN(n4758) );
  NAND2_X1 U5524 ( .A1(n4755), .A2(n4754), .ZN(n4753) );
  INV_X1 U5525 ( .A(n6297), .ZN(n4755) );
  NAND2_X1 U5526 ( .A1(n8848), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4754) );
  NAND2_X1 U5527 ( .A1(n6011), .A2(n6010), .ZN(n8884) );
  OR2_X1 U5528 ( .A1(n9014), .A2(n8958), .ZN(n4648) );
  NAND2_X1 U5529 ( .A1(n5074), .A2(n5073), .ZN(n8993) );
  OR2_X1 U5530 ( .A1(n10178), .A2(n7304), .ZN(n10128) );
  INV_X1 U5531 ( .A(n8925), .ZN(n8955) );
  INV_X1 U5532 ( .A(n9065), .ZN(n4814) );
  OR2_X1 U5533 ( .A1(n7314), .A2(n10128), .ZN(n8925) );
  OR2_X1 U5534 ( .A1(n6353), .A2(n6081), .ZN(n10129) );
  NAND2_X1 U5535 ( .A1(n10199), .A2(n10157), .ZN(n8991) );
  NAND2_X1 U5536 ( .A1(n8521), .A2(n6186), .ZN(n6371) );
  OAI21_X1 U5537 ( .B1(n4514), .B2(n10151), .A(n4512), .ZN(n9004) );
  AOI21_X1 U5538 ( .B1(n8736), .B2(n10131), .A(n4513), .ZN(n4512) );
  XNOR2_X1 U5539 ( .A(n8880), .B(n8879), .ZN(n4514) );
  NOR2_X1 U5540 ( .A1(n8899), .A2(n8946), .ZN(n4513) );
  AOI21_X1 U5541 ( .B1(n4653), .B2(n10136), .A(n4650), .ZN(n9009) );
  OAI21_X1 U5542 ( .B1(n8570), .B2(n4652), .A(n4651), .ZN(n4650) );
  XNOR2_X1 U5543 ( .A(n8890), .B(n8889), .ZN(n4653) );
  NAND2_X1 U5544 ( .A1(n8911), .A2(n10132), .ZN(n4651) );
  NAND2_X1 U5545 ( .A1(n5888), .A2(n5887), .ZN(n8716) );
  INV_X1 U5546 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7861) );
  OR2_X1 U5547 ( .A1(n5756), .A2(n4628), .ZN(n4465) );
  OAI21_X1 U5548 ( .B1(n9154), .B2(n6889), .A(n9151), .ZN(n6890) );
  AND3_X1 U5549 ( .A1(n5379), .A2(n5378), .A3(n5377), .ZN(n10089) );
  NAND2_X1 U5550 ( .A1(n7004), .A2(n5560), .ZN(n4457) );
  NAND2_X1 U5551 ( .A1(n9090), .A2(n6917), .ZN(n8273) );
  AND2_X1 U5552 ( .A1(n8271), .A2(n8272), .ZN(n6917) );
  NAND2_X1 U5553 ( .A1(n9091), .A2(n9092), .ZN(n9090) );
  OAI21_X1 U5554 ( .B1(n9621), .B2(n9186), .A(n8278), .ZN(n5146) );
  INV_X1 U5555 ( .A(n9417), .ZN(n4438) );
  NAND2_X1 U5556 ( .A1(n4625), .A2(n4623), .ZN(n9411) );
  NOR2_X1 U5557 ( .A1(n9273), .A2(n4624), .ZN(n4623) );
  INV_X1 U5558 ( .A(n5562), .ZN(n4624) );
  NAND2_X1 U5559 ( .A1(n6585), .A2(n6584), .ZN(n9627) );
  OR2_X1 U5560 ( .A1(n9642), .A2(n6615), .ZN(n6585) );
  INV_X1 U5561 ( .A(n7530), .ZN(n4580) );
  INV_X1 U5562 ( .A(n9200), .ZN(n9427) );
  AOI21_X1 U5563 ( .B1(n9499), .B2(n9498), .A(n9497), .ZN(n9496) );
  OR2_X1 U5564 ( .A1(n9519), .A2(n9520), .ZN(n4666) );
  NAND2_X1 U5565 ( .A1(n5164), .A2(n5160), .ZN(n9597) );
  NOR2_X1 U5566 ( .A1(n6970), .A2(n5165), .ZN(n6379) );
  NAND2_X1 U5567 ( .A1(n6623), .A2(n6622), .ZN(n6624) );
  XNOR2_X1 U5568 ( .A(n6614), .B(n6613), .ZN(n6625) );
  NAND2_X1 U5569 ( .A1(n7635), .A2(n9985), .ZN(n10072) );
  INV_X1 U5570 ( .A(n9884), .ZN(n9921) );
  INV_X1 U5571 ( .A(n10123), .ZN(n10120) );
  OAI21_X1 U5572 ( .B1(n6663), .B2(n5030), .A(n5028), .ZN(n6976) );
  NAND2_X1 U5573 ( .A1(n6663), .A2(n6662), .ZN(n4728) );
  INV_X1 U5574 ( .A(n5054), .ZN(n5053) );
  AND2_X1 U5575 ( .A1(n10115), .A2(n9930), .ZN(n9954) );
  INV_X1 U5576 ( .A(n9954), .ZN(n9975) );
  AND2_X1 U5577 ( .A1(n5616), .A2(n5615), .ZN(n9986) );
  INV_X1 U5578 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7787) );
  INV_X1 U5579 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U5580 ( .A1(n5496), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5498) );
  NOR2_X1 U5581 ( .A1(n10017), .A2(n10016), .ZN(n10387) );
  NOR2_X1 U5582 ( .A1(n10021), .A2(n10020), .ZN(n10222) );
  AOI21_X1 U5583 ( .B1(n10029), .B2(n10310), .A(n10028), .ZN(n10216) );
  NOR2_X1 U5584 ( .A1(n10218), .A2(n10217), .ZN(n10028) );
  NOR2_X1 U5585 ( .A1(n10034), .A2(n10033), .ZN(n10212) );
  NOR2_X1 U5586 ( .A1(n10214), .A2(n10213), .ZN(n10033) );
  NAND2_X1 U5587 ( .A1(n4553), .A2(n8339), .ZN(n8342) );
  AND2_X1 U5588 ( .A1(n8336), .A2(n8475), .ZN(n4554) );
  NAND2_X1 U5589 ( .A1(n8340), .A2(n8342), .ZN(n4818) );
  NAND2_X1 U5590 ( .A1(n4816), .A2(n4815), .ZN(n4539) );
  NAND2_X1 U5591 ( .A1(n8341), .A2(n8499), .ZN(n4815) );
  NAND2_X1 U5592 ( .A1(n4817), .A2(n8475), .ZN(n4816) );
  NAND2_X1 U5593 ( .A1(n4818), .A2(n8341), .ZN(n4817) );
  NOR2_X1 U5594 ( .A1(n4821), .A2(n4563), .ZN(n4820) );
  NAND2_X1 U5595 ( .A1(n8398), .A2(n8397), .ZN(n4821) );
  OAI21_X1 U5596 ( .B1(n4822), .B2(n4823), .A(n4364), .ZN(n4563) );
  NAND2_X1 U5597 ( .A1(n4466), .A2(n4683), .ZN(n9231) );
  NAND2_X1 U5598 ( .A1(n9226), .A2(n9352), .ZN(n4683) );
  NOR2_X1 U5599 ( .A1(n8418), .A2(n8499), .ZN(n4836) );
  INV_X1 U5600 ( .A(n9827), .ZN(n4680) );
  NAND2_X1 U5601 ( .A1(n9231), .A2(n4682), .ZN(n4681) );
  NAND2_X1 U5602 ( .A1(n4562), .A2(n5169), .ZN(n4561) );
  NAND2_X1 U5603 ( .A1(n4460), .A2(n4459), .ZN(n9238) );
  OR2_X1 U5604 ( .A1(n9236), .A2(n9237), .ZN(n4459) );
  NAND2_X1 U5605 ( .A1(n4805), .A2(n4461), .ZN(n4460) );
  NOR2_X1 U5606 ( .A1(n9649), .A2(n9352), .ZN(n9255) );
  OAI21_X1 U5607 ( .B1(n4556), .B2(n4555), .A(n8475), .ZN(n8426) );
  NAND2_X1 U5608 ( .A1(n8429), .A2(n4343), .ZN(n4555) );
  AOI21_X1 U5609 ( .B1(n4834), .B2(n4831), .A(n4340), .ZN(n4556) );
  AND2_X1 U5610 ( .A1(n4552), .A2(n8425), .ZN(n8427) );
  OAI21_X1 U5611 ( .B1(n8416), .B2(n4833), .A(n4829), .ZN(n4552) );
  AOI21_X1 U5612 ( .B1(n4830), .B2(n4832), .A(n4353), .ZN(n4829) );
  INV_X1 U5613 ( .A(n6116), .ZN(n4591) );
  OAI21_X1 U5614 ( .B1(n4592), .B2(n4591), .A(n8012), .ZN(n4590) );
  AND2_X1 U5615 ( .A1(n6635), .A2(n9211), .ZN(n9207) );
  OAI21_X1 U5616 ( .B1(n4543), .B2(n4542), .A(n4540), .ZN(n8467) );
  AOI21_X1 U5617 ( .B1(n4356), .B2(n8462), .A(n4541), .ZN(n4540) );
  INV_X1 U5618 ( .A(n8462), .ZN(n4542) );
  AOI21_X1 U5619 ( .B1(n8889), .B2(n4862), .A(n4348), .ZN(n4861) );
  INV_X1 U5620 ( .A(n4863), .ZN(n4862) );
  NAND2_X1 U5621 ( .A1(n8296), .A2(n4506), .ZN(n4505) );
  INV_X1 U5622 ( .A(n6127), .ZN(n4506) );
  NOR2_X1 U5623 ( .A1(n4352), .A2(n4846), .ZN(n4845) );
  INV_X1 U5624 ( .A(n6128), .ZN(n4846) );
  INV_X1 U5625 ( .A(n5533), .ZN(n4607) );
  NOR2_X1 U5626 ( .A1(n4711), .A2(n4614), .ZN(n4613) );
  INV_X1 U5627 ( .A(n5529), .ZN(n4614) );
  AOI21_X1 U5628 ( .B1(n5448), .B2(n4880), .A(n5258), .ZN(n4878) );
  INV_X1 U5629 ( .A(n4880), .ZN(n4879) );
  NAND2_X1 U5630 ( .A1(n4892), .A2(n5429), .ZN(n4646) );
  OAI21_X1 U5631 ( .B1(n5366), .B2(P1_DATAO_REG_11__SCAN_IN), .A(n4696), .ZN(
        n5246) );
  NAND2_X1 U5632 ( .A1(n5366), .A2(n7043), .ZN(n4696) );
  OAI21_X1 U5633 ( .B1(n5366), .B2(P1_DATAO_REG_8__SCAN_IN), .A(n4700), .ZN(
        n5229) );
  INV_X1 U5634 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4603) );
  INV_X1 U5635 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4602) );
  INV_X1 U5636 ( .A(n5986), .ZN(n5003) );
  NOR2_X1 U5637 ( .A1(n5000), .A2(n5004), .ZN(n4999) );
  INV_X1 U5638 ( .A(n6009), .ZN(n5004) );
  INV_X1 U5639 ( .A(n5982), .ZN(n5000) );
  INV_X1 U5640 ( .A(n8933), .ZN(n8247) );
  INV_X1 U5641 ( .A(n8610), .ZN(n8253) );
  NAND2_X1 U5642 ( .A1(n6043), .A2(n5696), .ZN(n4532) );
  NOR2_X1 U5643 ( .A1(n8480), .A2(n8323), .ZN(n8498) );
  NAND3_X1 U5644 ( .A1(n4293), .A2(n8325), .A3(n4675), .ZN(n8508) );
  INV_X1 U5645 ( .A(n8488), .ZN(n4675) );
  INV_X1 U5646 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U5647 ( .A1(n7563), .A2(n4439), .ZN(n6216) );
  AND2_X1 U5648 ( .A1(n8086), .A2(n6215), .ZN(n4439) );
  NOR2_X1 U5649 ( .A1(n5942), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n4769) );
  NOR2_X1 U5650 ( .A1(n6174), .A2(n6173), .ZN(n6175) );
  INV_X1 U5651 ( .A(n8366), .ZN(n6174) );
  INV_X1 U5652 ( .A(n8377), .ZN(n6173) );
  INV_X1 U5653 ( .A(n8369), .ZN(n8357) );
  AND2_X1 U5654 ( .A1(n5626), .A2(n5625), .ZN(n5701) );
  INV_X1 U5655 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U5656 ( .A1(n4366), .A2(n4692), .ZN(n6172) );
  OAI21_X1 U5657 ( .B1(n6170), .B2(n7382), .A(n6171), .ZN(n4581) );
  NAND2_X1 U5658 ( .A1(n8751), .A2(n10179), .ZN(n8369) );
  NAND2_X1 U5659 ( .A1(n4775), .A2(n7483), .ZN(n5779) );
  AND2_X1 U5660 ( .A1(n7298), .A2(n8341), .ZN(n10127) );
  INV_X1 U5661 ( .A(n6057), .ZN(n8338) );
  OR2_X1 U5662 ( .A1(n5083), .A2(n8281), .ZN(n5082) );
  AND2_X1 U5663 ( .A1(n8442), .A2(n5081), .ZN(n5080) );
  NOR2_X1 U5664 ( .A1(n8281), .A2(n5084), .ZN(n5081) );
  NAND2_X1 U5665 ( .A1(n8624), .A2(n4864), .ZN(n4863) );
  OR2_X1 U5666 ( .A1(n4867), .A2(n6133), .ZN(n4860) );
  AND2_X1 U5667 ( .A1(n8438), .A2(n8437), .ZN(n8304) );
  INV_X1 U5668 ( .A(n8410), .ZN(n4569) );
  AND2_X1 U5669 ( .A1(n8406), .A2(n8405), .ZN(n8403) );
  INV_X1 U5670 ( .A(n8395), .ZN(n8383) );
  INV_X1 U5671 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5645) );
  NOR2_X1 U5672 ( .A1(n5646), .A2(n4520), .ZN(n4480) );
  NOR2_X1 U5673 ( .A1(n5645), .A2(n4520), .ZN(n4517) );
  NAND2_X1 U5674 ( .A1(n5646), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4516) );
  AND2_X1 U5675 ( .A1(n5676), .A2(n5677), .ZN(n5023) );
  NAND2_X1 U5676 ( .A1(n5666), .A2(n5665), .ZN(n5774) );
  INV_X1 U5677 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5665) );
  NOR2_X1 U5678 ( .A1(n5113), .A2(n5124), .ZN(n5112) );
  NOR2_X1 U5679 ( .A1(n6875), .A2(n5123), .ZN(n5113) );
  NOR2_X1 U5680 ( .A1(n9162), .A2(n5127), .ZN(n5120) );
  AND2_X2 U5681 ( .A1(n6724), .A2(n6717), .ZN(n6740) );
  OR2_X1 U5682 ( .A1(n6721), .A2(n6720), .ZN(n6723) );
  NAND2_X1 U5683 ( .A1(n9336), .A2(n4875), .ZN(n4874) );
  NOR2_X1 U5684 ( .A1(n9332), .A2(n9352), .ZN(n4875) );
  AND2_X1 U5685 ( .A1(n9268), .A2(n9352), .ZN(n4868) );
  NOR2_X1 U5686 ( .A1(n4793), .A2(n9601), .ZN(n4670) );
  INV_X1 U5687 ( .A(n4794), .ZN(n4671) );
  OAI211_X1 U5688 ( .C1(n4799), .C2(n4791), .A(n9351), .B(n4789), .ZN(n4788)
         );
  OR2_X1 U5689 ( .A1(n4797), .A2(n4794), .ZN(n4791) );
  INV_X1 U5690 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10238) );
  OAI21_X1 U5691 ( .B1(n7283), .B2(n7685), .A(n7684), .ZN(n9534) );
  INV_X1 U5692 ( .A(n6717), .ZN(n7029) );
  NAND2_X1 U5693 ( .A1(n4976), .A2(n9313), .ZN(n4975) );
  AND2_X1 U5694 ( .A1(n5151), .A2(n5150), .ZN(n5149) );
  NOR2_X1 U5695 ( .A1(n6553), .A2(n6552), .ZN(n4689) );
  NAND2_X1 U5696 ( .A1(n9709), .A2(n4716), .ZN(n4715) );
  INV_X1 U5697 ( .A(n4954), .ZN(n4716) );
  NOR2_X1 U5698 ( .A1(n6513), .A2(n6512), .ZN(n4690) );
  NOR2_X1 U5699 ( .A1(n6496), .A2(n6399), .ZN(n6391) );
  NAND2_X1 U5700 ( .A1(n7761), .A2(n7848), .ZN(n7844) );
  AND2_X1 U5701 ( .A1(n7764), .A2(n9377), .ZN(n4566) );
  NAND2_X1 U5702 ( .A1(n4285), .A2(n6421), .ZN(n4952) );
  INV_X1 U5703 ( .A(n6421), .ZN(n4953) );
  AND2_X2 U5704 ( .A1(n6669), .A2(n9414), .ZN(n6720) );
  NAND2_X1 U5705 ( .A1(n9628), .A2(n9834), .ZN(n4723) );
  NAND2_X1 U5706 ( .A1(n9741), .A2(n9742), .ZN(n4739) );
  INV_X1 U5707 ( .A(n4312), .ZN(n5037) );
  AND2_X1 U5708 ( .A1(n6665), .A2(n9414), .ZN(n6721) );
  OR2_X1 U5709 ( .A1(n5318), .A2(n5317), .ZN(n5320) );
  AND2_X1 U5710 ( .A1(n5544), .A2(n5309), .ZN(n5542) );
  INV_X1 U5711 ( .A(n5537), .ZN(n4597) );
  INV_X1 U5712 ( .A(n5538), .ZN(n4598) );
  INV_X1 U5713 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U5714 ( .A1(n4351), .A2(n4710), .ZN(n4709) );
  AND2_X1 U5715 ( .A1(n4288), .A2(n5337), .ZN(n4710) );
  AOI21_X1 U5716 ( .B1(n4613), .B2(n4611), .A(n4610), .ZN(n4609) );
  INV_X1 U5717 ( .A(n5294), .ZN(n4610) );
  INV_X1 U5718 ( .A(n5287), .ZN(n4611) );
  INV_X1 U5719 ( .A(n4613), .ZN(n4612) );
  NAND2_X1 U5720 ( .A1(n5566), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5568) );
  INV_X1 U5721 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5567) );
  NOR2_X1 U5722 ( .A1(n5280), .A2(n4897), .ZN(n4896) );
  INV_X1 U5723 ( .A(n5272), .ZN(n4897) );
  NAND2_X1 U5724 ( .A1(n5564), .A2(n5563), .ZN(n5571) );
  NOR2_X1 U5725 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5563) );
  INV_X1 U5726 ( .A(n4443), .ZN(n5564) );
  NAND2_X1 U5727 ( .A1(n4442), .A2(n5142), .ZN(n4443) );
  AND2_X1 U5728 ( .A1(n5140), .A2(n4288), .ZN(n4442) );
  AND2_X1 U5729 ( .A1(n5143), .A2(n5488), .ZN(n5140) );
  INV_X1 U5730 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5488) );
  INV_X1 U5731 ( .A(n4621), .ZN(n4620) );
  NOR2_X1 U5732 ( .A1(n5432), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5444) );
  NOR2_X1 U5733 ( .A1(n4713), .A2(n4881), .ZN(n4885) );
  INV_X1 U5734 ( .A(n5226), .ZN(n4881) );
  NAND2_X1 U5735 ( .A1(n5352), .A2(n6986), .ZN(n5212) );
  CLKBUF_X1 U5736 ( .A(n5352), .Z(n4659) );
  NAND2_X1 U5737 ( .A1(n5347), .A2(n6992), .ZN(n4660) );
  INV_X1 U5738 ( .A(n8250), .ZN(n4530) );
  INV_X1 U5739 ( .A(n5786), .ZN(n5014) );
  INV_X1 U5740 ( .A(n5015), .ZN(n5012) );
  OR2_X1 U5741 ( .A1(n7349), .A2(n4477), .ZN(n4534) );
  INV_X1 U5742 ( .A(n5006), .ZN(n4477) );
  AOI21_X1 U5743 ( .B1(n7350), .B2(n5015), .A(n7471), .ZN(n5006) );
  NAND2_X1 U5744 ( .A1(n8650), .A2(n4703), .ZN(n4702) );
  INV_X1 U5745 ( .A(n5883), .ZN(n5018) );
  NAND2_X1 U5746 ( .A1(n8474), .A2(n8473), .ZN(n8485) );
  AND2_X1 U5747 ( .A1(n4842), .A2(n8325), .ZN(n8503) );
  NOR2_X1 U5748 ( .A1(n8507), .A2(n4551), .ZN(n4550) );
  NAND2_X1 U5749 ( .A1(n4842), .A2(n4840), .ZN(n8495) );
  OR2_X1 U5750 ( .A1(n8488), .A2(n8489), .ZN(n4712) );
  NOR2_X1 U5751 ( .A1(n8733), .A2(n8999), .ZN(n4841) );
  AND2_X1 U5752 ( .A1(n8318), .A2(n8317), .ZN(n8859) );
  OR2_X1 U5754 ( .A1(n7142), .A2(n7313), .ZN(n7140) );
  NAND2_X1 U5755 ( .A1(n6298), .A2(n4427), .ZN(n7146) );
  NAND2_X1 U5756 ( .A1(n4428), .A2(n4338), .ZN(n4427) );
  NOR2_X1 U5757 ( .A1(n7146), .A2(n10189), .ZN(n7145) );
  XNOR2_X1 U5758 ( .A(n7015), .B(n10147), .ZN(n8762) );
  XNOR2_X1 U5759 ( .A(n7015), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n8757) );
  NOR2_X1 U5760 ( .A1(n8757), .A2(n8756), .ZN(n8755) );
  AND2_X1 U5761 ( .A1(n7237), .A2(n4948), .ZN(n7157) );
  OR2_X1 U5762 ( .A1(n6302), .A2(n10195), .ZN(n4947) );
  OR2_X1 U5763 ( .A1(n7238), .A2(n4946), .ZN(n4945) );
  NOR2_X1 U5764 ( .A1(n7154), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4946) );
  NAND2_X1 U5765 ( .A1(n4944), .A2(n7154), .ZN(n7237) );
  INV_X1 U5766 ( .A(n6303), .ZN(n4944) );
  NAND2_X1 U5767 ( .A1(n4902), .A2(n7244), .ZN(n4444) );
  AOI21_X1 U5768 ( .B1(n4751), .B2(n7164), .A(n4355), .ZN(n4750) );
  INV_X1 U5769 ( .A(n6245), .ZN(n4751) );
  AND2_X1 U5770 ( .A1(n6213), .A2(n7606), .ZN(n4447) );
  INV_X1 U5771 ( .A(n6309), .ZN(n7555) );
  NAND2_X1 U5772 ( .A1(n4386), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8085) );
  INV_X1 U5773 ( .A(n6316), .ZN(n4938) );
  NAND2_X1 U5774 ( .A1(n7968), .A2(n4449), .ZN(n6218) );
  AND2_X1 U5775 ( .A1(n6217), .A2(n6315), .ZN(n4449) );
  INV_X1 U5776 ( .A(n4942), .ZN(n8791) );
  NAND2_X1 U5777 ( .A1(n7968), .A2(n6217), .ZN(n4645) );
  AND2_X1 U5778 ( .A1(n8811), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8809) );
  NAND2_X1 U5779 ( .A1(n6220), .A2(n4916), .ZN(n4913) );
  NOR2_X1 U5780 ( .A1(n8821), .A2(n4915), .ZN(n4914) );
  AND2_X1 U5781 ( .A1(n8487), .A2(n8322), .ZN(n8320) );
  INV_X1 U5782 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n4783) );
  OR2_X1 U5783 ( .A1(n6141), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8523) );
  AND2_X1 U5784 ( .A1(n8318), .A2(n6157), .ZN(n6366) );
  NAND2_X1 U5785 ( .A1(n4767), .A2(n5634), .ZN(n6014) );
  NAND2_X1 U5786 ( .A1(n4769), .A2(n4768), .ZN(n5989) );
  INV_X1 U5787 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n4768) );
  AND2_X1 U5788 ( .A1(n4305), .A2(n4781), .ZN(n4780) );
  INV_X1 U5789 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n4781) );
  NAND2_X1 U5790 ( .A1(n4847), .A2(n6128), .ZN(n8217) );
  NAND2_X1 U5791 ( .A1(n8205), .A2(n8296), .ZN(n4847) );
  NAND2_X1 U5792 ( .A1(n5633), .A2(n4305), .ZN(n5960) );
  NAND2_X1 U5793 ( .A1(n5633), .A2(n5632), .ZN(n5958) );
  AND2_X1 U5794 ( .A1(n4304), .A2(n4778), .ZN(n4777) );
  INV_X1 U5795 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n4778) );
  NAND2_X1 U5796 ( .A1(n5631), .A2(n4304), .ZN(n5889) );
  NAND2_X1 U5797 ( .A1(n5631), .A2(n5630), .ZN(n5875) );
  NAND2_X1 U5798 ( .A1(n4770), .A2(n5629), .ZN(n5861) );
  INV_X1 U5799 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5629) );
  INV_X1 U5800 ( .A(n5852), .ZN(n4770) );
  NAND2_X1 U5801 ( .A1(n4774), .A2(n4773), .ZN(n5831) );
  INV_X1 U5802 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n4773) );
  INV_X1 U5803 ( .A(n5829), .ZN(n4774) );
  NAND2_X1 U5804 ( .A1(n4772), .A2(n4771), .ZN(n5852) );
  INV_X1 U5805 ( .A(n5831), .ZN(n4772) );
  NAND2_X1 U5806 ( .A1(n5701), .A2(n5627), .ZN(n5797) );
  INV_X1 U5807 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U5808 ( .A1(n4865), .A2(n4863), .ZN(n8890) );
  NAND2_X1 U5809 ( .A1(n4857), .A2(n4858), .ZN(n4865) );
  INV_X1 U5810 ( .A(n4860), .ZN(n4858) );
  NAND2_X1 U5811 ( .A1(n5973), .A2(n5972), .ZN(n8675) );
  NAND2_X1 U5812 ( .A1(n4533), .A2(n6127), .ZN(n8205) );
  NAND2_X1 U5813 ( .A1(n4498), .A2(n6125), .ZN(n8157) );
  AND2_X1 U5814 ( .A1(n8419), .A2(n8417), .ZN(n8298) );
  NAND2_X1 U5815 ( .A1(n4584), .A2(n4593), .ZN(n7862) );
  NAND2_X1 U5816 ( .A1(n8384), .A2(n8382), .ZN(n8288) );
  NOR2_X1 U5817 ( .A1(n5656), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n4839) );
  OR2_X1 U5818 ( .A1(n5689), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U5819 ( .A1(n5680), .A2(n5679), .ZN(n5682) );
  NAND2_X1 U5820 ( .A1(n5871), .A2(n5676), .ZN(n5954) );
  XNOR2_X1 U5821 ( .A(n5794), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7016) );
  NAND2_X1 U5822 ( .A1(n5664), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5734) );
  NAND2_X1 U5823 ( .A1(n4628), .A2(n4520), .ZN(n4627) );
  NAND2_X1 U5824 ( .A1(n4844), .A2(n4429), .ZN(n5755) );
  NOR2_X1 U5825 ( .A1(n5100), .A2(n5103), .ZN(n5099) );
  OR2_X1 U5826 ( .A1(n6526), .A2(n6525), .ZN(n6537) );
  NOR2_X1 U5827 ( .A1(n9140), .A2(n5135), .ZN(n5134) );
  INV_X1 U5828 ( .A(n6879), .ZN(n5135) );
  INV_X1 U5829 ( .A(n6868), .ZN(n6869) );
  OAI21_X1 U5830 ( .B1(n6867), .B2(n9104), .A(n6866), .ZN(n6868) );
  NOR2_X1 U5831 ( .A1(n5189), .A2(n6863), .ZN(n6864) );
  NAND2_X1 U5832 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6436) );
  NAND2_X1 U5833 ( .A1(n6389), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U5834 ( .A1(n4686), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6494) );
  INV_X1 U5835 ( .A(n6487), .ZN(n4686) );
  INV_X1 U5836 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U5837 ( .A1(n6833), .A2(n6834), .ZN(n8061) );
  NAND2_X1 U5838 ( .A1(n4690), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6526) );
  NAND2_X1 U5839 ( .A1(n9131), .A2(n6771), .ZN(n7617) );
  NAND2_X1 U5840 ( .A1(n4669), .A2(n4667), .ZN(n9308) );
  AND2_X1 U5841 ( .A1(n4668), .A2(n4371), .ZN(n4667) );
  NAND2_X1 U5842 ( .A1(n6588), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6411) );
  NAND2_X1 U5843 ( .A1(n7050), .A2(n9445), .ZN(n9469) );
  AOI21_X1 U5844 ( .B1(n10049), .B2(n10048), .A(n10047), .ZN(n9480) );
  INV_X1 U5845 ( .A(n5337), .ZN(n5408) );
  NOR3_X1 U5846 ( .A1(n7204), .A2(n7203), .A3(n7207), .ZN(n7205) );
  NAND2_X1 U5847 ( .A1(n7686), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n9538) );
  NOR2_X1 U5848 ( .A1(n9569), .A2(n9570), .ZN(n9573) );
  NOR2_X1 U5849 ( .A1(n9565), .A2(n4663), .ZN(n9581) );
  OR2_X1 U5850 ( .A1(n9563), .A2(n9564), .ZN(n4663) );
  NAND2_X1 U5851 ( .A1(n9573), .A2(n9572), .ZN(n9585) );
  NOR2_X1 U5852 ( .A1(n5165), .A2(n8581), .ZN(n5163) );
  AND3_X1 U5853 ( .A1(n5159), .A2(n9274), .A3(n6975), .ZN(n5161) );
  INV_X1 U5854 ( .A(n5165), .ZN(n5159) );
  OR2_X1 U5855 ( .A1(n4796), .A2(n9269), .ZN(n5165) );
  INV_X1 U5856 ( .A(n9306), .ZN(n6613) );
  AND2_X1 U5857 ( .A1(n6597), .A2(n6587), .ZN(n9623) );
  NAND2_X1 U5858 ( .A1(n9693), .A2(n5151), .ZN(n9656) );
  AND2_X1 U5859 ( .A1(n6568), .A2(n6567), .ZN(n9652) );
  NAND2_X1 U5860 ( .A1(n4689), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6571) );
  INV_X1 U5861 ( .A(n4689), .ZN(n6561) );
  BUF_X1 U5862 ( .A(n9682), .Z(n9712) );
  NAND2_X1 U5863 ( .A1(n4714), .A2(n4954), .ZN(n9710) );
  NAND2_X1 U5864 ( .A1(n9775), .A2(n4718), .ZN(n4714) );
  NAND2_X1 U5865 ( .A1(n4957), .A2(n4959), .ZN(n9727) );
  NAND2_X1 U5866 ( .A1(n9764), .A2(n4960), .ZN(n4957) );
  AND2_X1 U5867 ( .A1(n9817), .A2(n5157), .ZN(n9779) );
  AND2_X1 U5868 ( .A1(n5157), .A2(n9763), .ZN(n5156) );
  OR2_X1 U5869 ( .A1(n9741), .A2(n9740), .ZN(n9758) );
  INV_X1 U5870 ( .A(n4690), .ZN(n6519) );
  NAND2_X1 U5871 ( .A1(n9817), .A2(n5158), .ZN(n9789) );
  AND2_X1 U5872 ( .A1(n9812), .A2(n9810), .ZN(n6502) );
  CLKBUF_X1 U5873 ( .A(n9817), .Z(n9839) );
  NAND2_X1 U5874 ( .A1(n8098), .A2(n9296), .ZN(n9828) );
  OR2_X1 U5875 ( .A1(n6494), .A2(n6493), .ZN(n6496) );
  NAND2_X1 U5876 ( .A1(n7933), .A2(n9380), .ZN(n8098) );
  AND4_X1 U5877 ( .A1(n6483), .A2(n6482), .A3(n6481), .A4(n6480), .ZN(n7981)
         );
  NOR2_X1 U5878 ( .A1(n5154), .A2(n7875), .ZN(n5152) );
  NAND2_X1 U5879 ( .A1(n5155), .A2(n4580), .ZN(n9211) );
  AND4_X1 U5880 ( .A1(n6461), .A2(n6460), .A3(n6459), .A4(n6458), .ZN(n7998)
         );
  AND4_X1 U5881 ( .A1(n6468), .A2(n6467), .A3(n6466), .A4(n6465), .ZN(n7997)
         );
  NAND2_X1 U5882 ( .A1(n7823), .A2(n5153), .ZN(n7989) );
  NAND2_X1 U5883 ( .A1(n6627), .A2(n7401), .ZN(n7400) );
  NOR2_X1 U5884 ( .A1(n9864), .A2(n6665), .ZN(n7635) );
  NAND2_X1 U5885 ( .A1(n8198), .A2(n5560), .ZN(n4898) );
  AOI21_X1 U5886 ( .B1(n4724), .B2(n9829), .A(n4721), .ZN(n9857) );
  NAND2_X1 U5887 ( .A1(n4723), .A2(n4722), .ZN(n4721) );
  OAI21_X1 U5888 ( .B1(n9625), .B2(n9626), .A(n9624), .ZN(n4724) );
  NAND2_X1 U5889 ( .A1(n9627), .A2(n9836), .ZN(n4722) );
  NAND2_X1 U5890 ( .A1(n5532), .A2(n5531), .ZN(n9660) );
  AND2_X1 U5891 ( .A1(n9249), .A2(n9246), .ZN(n9725) );
  NAND2_X1 U5892 ( .A1(n6837), .A2(n4638), .ZN(n4637) );
  INV_X1 U5893 ( .A(n8075), .ZN(n5155) );
  OR2_X1 U5894 ( .A1(n7652), .A2(n6721), .ZN(n10107) );
  NAND2_X1 U5895 ( .A1(n7416), .A2(n9279), .ZN(n4951) );
  NAND2_X1 U5896 ( .A1(n6990), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5051) );
  NAND2_X1 U5897 ( .A1(n7637), .A2(n9933), .ZN(n10112) );
  OAI211_X1 U5898 ( .C1(P1_B_REG_SCAN_IN), .C2(n8143), .A(n5612), .B(n5601), 
        .ZN(n9983) );
  XNOR2_X1 U5899 ( .A(n5555), .B(n5554), .ZN(n8588) );
  NOR2_X1 U5900 ( .A1(n5579), .A2(n5489), .ZN(n5576) );
  INV_X1 U5901 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5579) );
  INV_X1 U5902 ( .A(SI_29_), .ZN(n4691) );
  MUX2_X1 U5903 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5342), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5343) );
  XNOR2_X1 U5904 ( .A(n5547), .B(n5546), .ZN(n8530) );
  NAND2_X1 U5905 ( .A1(n5545), .A2(n5544), .ZN(n5547) );
  NAND2_X1 U5906 ( .A1(n5543), .A2(n5542), .ZN(n5545) );
  XNOR2_X1 U5907 ( .A(n5346), .B(n5345), .ZN(n5574) );
  XNOR2_X1 U5908 ( .A(n5543), .B(n5542), .ZN(n9061) );
  XNOR2_X1 U5909 ( .A(n5538), .B(n5537), .ZN(n8198) );
  XNOR2_X1 U5910 ( .A(n5510), .B(n5509), .ZN(n8039) );
  NAND2_X1 U5911 ( .A1(n4615), .A2(n4616), .ZN(n5493) );
  NAND2_X1 U5912 ( .A1(n4619), .A2(n5264), .ZN(n5487) );
  OR2_X1 U5913 ( .A1(n5481), .A2(n5480), .ZN(n4619) );
  XNOR2_X1 U5914 ( .A(n5472), .B(n5460), .ZN(n7345) );
  OAI21_X1 U5915 ( .B1(n5421), .B2(n4889), .A(n4886), .ZN(n5442) );
  NAND2_X1 U5916 ( .A1(n4583), .A2(n5226), .ZN(n4458) );
  XNOR2_X1 U5917 ( .A(n5209), .B(SI_3_), .ZN(n5371) );
  AND4_X1 U5918 ( .A1(n5802), .A2(n5801), .A3(n5800), .A4(n5799), .ZN(n7810)
         );
  INV_X1 U5919 ( .A(n6350), .ZN(n4981) );
  AND4_X1 U5920 ( .A1(n5814), .A2(n5813), .A3(n5812), .A4(n5811), .ZN(n7923)
         );
  NAND2_X1 U5921 ( .A1(n8687), .A2(n5192), .ZN(n4997) );
  NOR2_X1 U5922 ( .A1(n8649), .A2(n4474), .ZN(n8651) );
  INV_X1 U5923 ( .A(n8648), .ZN(n4475) );
  NAND2_X1 U5924 ( .A1(n4471), .A2(n4986), .ZN(n4468) );
  NAND2_X1 U5925 ( .A1(n6161), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5731) );
  OR2_X1 U5926 ( .A1(n4282), .A2(n5728), .ZN(n5733) );
  AND4_X1 U5927 ( .A1(n5706), .A2(n5705), .A3(n5704), .A4(n5703), .ZN(n7696)
         );
  NAND2_X1 U5928 ( .A1(n5019), .A2(n5883), .ZN(n8719) );
  NAND2_X1 U5929 ( .A1(n5019), .A2(n4289), .ZN(n8720) );
  INV_X1 U5930 ( .A(n8859), .ZN(n8733) );
  INV_X1 U5931 ( .A(n8899), .ZN(n8737) );
  INV_X1 U5932 ( .A(n8920), .ZN(n8738) );
  INV_X1 U5933 ( .A(n8255), .ZN(n8910) );
  INV_X1 U5934 ( .A(n8947), .ZN(n8740) );
  INV_X1 U5935 ( .A(n8708), .ZN(n8158) );
  OR2_X1 U5936 ( .A1(n6230), .A2(n6203), .ZN(n8742) );
  INV_X1 U5937 ( .A(n7923), .ZN(n8748) );
  INV_X1 U5938 ( .A(n7810), .ZN(n8749) );
  INV_X1 U5939 ( .A(n7696), .ZN(n8750) );
  INV_X1 U5940 ( .A(n7474), .ZN(n8751) );
  INV_X1 U5941 ( .A(n7440), .ZN(n8753) );
  NAND2_X1 U5942 ( .A1(n7184), .A2(n7183), .ZN(n7182) );
  NAND2_X1 U5943 ( .A1(n4749), .A2(n4750), .ZN(n7233) );
  NAND2_X1 U5944 ( .A1(n7231), .A2(n6249), .ZN(n7325) );
  NAND2_X1 U5945 ( .A1(n4909), .A2(n7372), .ZN(n7374) );
  INV_X1 U5946 ( .A(n4910), .ZN(n4909) );
  NAND2_X1 U5947 ( .A1(n6307), .A2(n4937), .ZN(n7327) );
  NAND2_X1 U5948 ( .A1(n4932), .A2(n6309), .ZN(n7609) );
  NAND2_X1 U5949 ( .A1(n6261), .A2(n6260), .ZN(n7552) );
  OAI21_X1 U5950 ( .B1(n6261), .B2(n4486), .A(n4484), .ZN(n8083) );
  AOI21_X1 U5951 ( .B1(n7553), .B2(n4485), .A(n4387), .ZN(n4484) );
  INV_X1 U5952 ( .A(n7553), .ZN(n4486) );
  OAI21_X1 U5953 ( .B1(n7961), .B2(n7963), .A(n7962), .ZN(n7960) );
  OAI21_X1 U5954 ( .B1(n6271), .B2(n4746), .A(n4744), .ZN(n8787) );
  NAND2_X1 U5955 ( .A1(n4421), .A2(n4425), .ZN(n8808) );
  INV_X1 U5956 ( .A(n4422), .ZN(n4421) );
  OAI21_X1 U5957 ( .B1(n6271), .B2(n4742), .A(n4487), .ZN(n8806) );
  AOI21_X1 U5958 ( .B1(n4488), .B2(n4745), .A(n4306), .ZN(n4487) );
  NAND2_X1 U5959 ( .A1(n4912), .A2(n4913), .ZN(n8820) );
  NAND2_X1 U5960 ( .A1(n4431), .A2(n6323), .ZN(n4430) );
  INV_X1 U5961 ( .A(n4432), .ZN(n4431) );
  INV_X1 U5962 ( .A(n8326), .ZN(n8524) );
  NAND2_X1 U5963 ( .A1(n5063), .A2(n5067), .ZN(n6370) );
  NAND2_X1 U5964 ( .A1(n8878), .A2(n5070), .ZN(n5063) );
  OAI21_X1 U5965 ( .B1(n8878), .B2(n5072), .A(n8468), .ZN(n8871) );
  AOI21_X1 U5966 ( .B1(n8869), .B2(n10136), .A(n8868), .ZN(n8964) );
  NAND2_X1 U5967 ( .A1(n8867), .A2(n8866), .ZN(n8868) );
  XNOR2_X1 U5968 ( .A(n8864), .B(n8870), .ZN(n8869) );
  AND2_X1 U5969 ( .A1(n4510), .A2(n4321), .ZN(n8917) );
  AOI21_X1 U5970 ( .B1(n8228), .B2(n8430), .A(n5090), .ZN(n8922) );
  NAND2_X1 U5971 ( .A1(n5077), .A2(n8421), .ZN(n8222) );
  NAND2_X1 U5972 ( .A1(n5074), .A2(n8405), .ZN(n8030) );
  NAND2_X1 U5973 ( .A1(n5828), .A2(n5827), .ZN(n5839) );
  NAND2_X1 U5974 ( .A1(n5712), .A2(n5711), .ZN(n7702) );
  INV_X1 U5975 ( .A(n7339), .ZN(n10161) );
  NAND2_X1 U5976 ( .A1(n5754), .A2(n4334), .ZN(n5057) );
  AND2_X1 U5977 ( .A1(n7258), .A2(n8343), .ZN(n10150) );
  AND2_X1 U5978 ( .A1(n6357), .A2(n6356), .ZN(n6361) );
  NAND2_X1 U5979 ( .A1(n8529), .A2(n6188), .ZN(n6362) );
  NAND2_X1 U5980 ( .A1(n6187), .A2(n6186), .ZN(n6188) );
  INV_X1 U5981 ( .A(n8884), .ZN(n9005) );
  NAND2_X1 U5982 ( .A1(n6013), .A2(n6012), .ZN(n9011) );
  OAI21_X1 U5983 ( .B1(n5086), .B2(n8228), .A(n5078), .ZN(n8902) );
  AOI21_X1 U5984 ( .B1(n5085), .B2(n5084), .A(n5083), .ZN(n5078) );
  NAND2_X1 U5985 ( .A1(n4857), .A2(n4866), .ZN(n8897) );
  NAND2_X1 U5986 ( .A1(n5988), .A2(n5987), .ZN(n9021) );
  NAND2_X1 U5987 ( .A1(n5087), .A2(n5088), .ZN(n8907) );
  NAND2_X1 U5988 ( .A1(n8228), .A2(n4313), .ZN(n5087) );
  NAND2_X1 U5989 ( .A1(n4852), .A2(n4851), .ZN(n8931) );
  AND2_X1 U5990 ( .A1(n8951), .A2(n8950), .ZN(n9036) );
  NAND2_X1 U5991 ( .A1(n8224), .A2(n8422), .ZN(n8940) );
  NAND2_X1 U5992 ( .A1(n5914), .A2(n5913), .ZN(n8644) );
  NAND2_X1 U5993 ( .A1(n6181), .A2(n8419), .ZN(n8204) );
  NAND2_X1 U5994 ( .A1(n5902), .A2(n5901), .ZN(n8634) );
  NAND2_X1 U5995 ( .A1(n8025), .A2(n6124), .ZN(n8145) );
  NAND2_X1 U5996 ( .A1(n8993), .A2(n8410), .ZN(n8144) );
  NAND2_X1 U5997 ( .A1(n5850), .A2(n5849), .ZN(n8185) );
  NAND2_X1 U5998 ( .A1(n6115), .A2(n6114), .ZN(n7863) );
  NAND2_X1 U5999 ( .A1(n7042), .A2(n8310), .ZN(n5819) );
  NAND2_X1 U6000 ( .A1(n4585), .A2(n5094), .ZN(n7717) );
  INV_X1 U6001 ( .A(n5839), .ZN(n8197) );
  NAND2_X1 U6002 ( .A1(n5807), .A2(n5806), .ZN(n7627) );
  AND2_X1 U6003 ( .A1(n6196), .A2(n6195), .ZN(n10186) );
  OR2_X1 U6004 ( .A1(n6190), .A2(n6189), .ZN(n6196) );
  AND2_X1 U6005 ( .A1(n6229), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7010) );
  NAND2_X1 U6006 ( .A1(n7007), .A2(n7006), .ZN(n7023) );
  NAND2_X1 U6007 ( .A1(n6069), .A2(n5644), .ZN(n9047) );
  INV_X1 U6008 ( .A(n4501), .ZN(n4500) );
  NAND2_X1 U6009 ( .A1(n6069), .A2(n4341), .ZN(n4502) );
  OR2_X1 U6010 ( .A1(n6069), .A2(n4504), .ZN(n4503) );
  INV_X1 U6011 ( .A(n5647), .ZN(n9055) );
  NAND2_X1 U6012 ( .A1(n5692), .A2(n5691), .ZN(n8203) );
  MUX2_X1 U6013 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5690), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5692) );
  OAI21_X1 U6014 ( .B1(n5055), .B2(n5689), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5690) );
  INV_X1 U6015 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8172) );
  INV_X1 U6016 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8140) );
  NAND2_X1 U6017 ( .A1(n5055), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5684) );
  INV_X1 U6018 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8035) );
  INV_X1 U6019 ( .A(n8513), .ZN(n8337) );
  INV_X1 U6020 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8575) );
  INV_X1 U6021 ( .A(n8500), .ZN(n8479) );
  INV_X1 U6022 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7678) );
  INV_X1 U6023 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7398) );
  INV_X1 U6024 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10323) );
  INV_X1 U6025 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7027) );
  INV_X1 U6026 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7022) );
  NAND2_X1 U6027 ( .A1(n5106), .A2(n4337), .ZN(n5105) );
  AND2_X1 U6028 ( .A1(n4294), .A2(n8261), .ZN(n5107) );
  AND2_X1 U6029 ( .A1(n8553), .A2(n9175), .ZN(n8554) );
  NOR2_X1 U6030 ( .A1(n6929), .A2(n6928), .ZN(n6927) );
  NAND2_X1 U6031 ( .A1(n6737), .A2(n6736), .ZN(n6744) );
  NAND2_X1 U6032 ( .A1(n5139), .A2(n9141), .ZN(n9084) );
  NAND2_X1 U6033 ( .A1(n4673), .A2(n5134), .ZN(n5139) );
  NAND2_X1 U6034 ( .A1(n5394), .A2(n5393), .ZN(n7900) );
  NAND2_X1 U6035 ( .A1(n6870), .A2(n6869), .ZN(n9113) );
  NAND2_X1 U6036 ( .A1(n9133), .A2(n9132), .ZN(n9131) );
  AND4_X1 U6037 ( .A1(n6477), .A2(n6476), .A3(n6475), .A4(n6474), .ZN(n7888)
         );
  AND2_X1 U6038 ( .A1(n6549), .A2(n6548), .ZN(n9729) );
  NAND2_X1 U6039 ( .A1(n4673), .A2(n6879), .ZN(n9144) );
  INV_X1 U6040 ( .A(n5104), .ZN(n8262) );
  AOI21_X1 U6041 ( .B1(n4294), .B2(n5109), .A(n4322), .ZN(n5104) );
  AOI21_X1 U6042 ( .B1(n5136), .B2(n5132), .A(n4326), .ZN(n5131) );
  INV_X1 U6043 ( .A(n9141), .ZN(n5132) );
  NAND2_X1 U6044 ( .A1(n5516), .A2(n5515), .ZN(n9877) );
  AND2_X1 U6045 ( .A1(n5118), .A2(n4401), .ZN(n9161) );
  INV_X1 U6046 ( .A(n9181), .ZN(n9155) );
  AND3_X1 U6047 ( .A1(n6511), .A2(n6510), .A3(n6509), .ZN(n9180) );
  NAND2_X1 U6048 ( .A1(n6946), .A2(n9834), .ZN(n9181) );
  OR2_X1 U6049 ( .A1(n9607), .A2(n6615), .ZN(n6603) );
  INV_X1 U6050 ( .A(n9652), .ZN(n9688) );
  INV_X1 U6051 ( .A(n9180), .ZN(n9815) );
  INV_X1 U6052 ( .A(n9807), .ZN(n9814) );
  INV_X1 U6053 ( .A(n7998), .ZN(n9426) );
  INV_X1 U6054 ( .A(n7647), .ZN(n9428) );
  NAND2_X1 U6055 ( .A1(n9472), .A2(n9473), .ZN(n10058) );
  OAI211_X1 U6056 ( .C1(n9486), .C2(n9502), .A(n7074), .B(n7073), .ZN(n9508)
         );
  OAI21_X1 U6057 ( .B1(n9496), .B2(n7120), .A(n7057), .ZN(n7132) );
  AOI22_X1 U6058 ( .A1(n7117), .A2(n7116), .B1(n7121), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7129) );
  AND2_X1 U6059 ( .A1(n5412), .A2(n5417), .ZN(n7137) );
  AND2_X1 U6060 ( .A1(n7088), .A2(n7087), .ZN(n7204) );
  AOI21_X1 U6061 ( .B1(n7286), .B2(n7285), .A(n7284), .ZN(n9514) );
  NAND2_X1 U6062 ( .A1(n9518), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4664) );
  NAND2_X1 U6063 ( .A1(n4662), .A2(n4661), .ZN(n9550) );
  INV_X1 U6064 ( .A(n9537), .ZN(n4661) );
  NAND2_X1 U6065 ( .A1(n9538), .A2(n9539), .ZN(n4662) );
  NAND2_X1 U6066 ( .A1(n7033), .A2(n7035), .ZN(n9596) );
  AOI21_X1 U6067 ( .B1(n9421), .B2(n9836), .A(n6966), .ZN(n6967) );
  NAND2_X1 U6068 ( .A1(n6707), .A2(n6706), .ZN(n6708) );
  OR3_X1 U6069 ( .A1(n6712), .A2(n6711), .A3(n9864), .ZN(n9611) );
  XNOR2_X1 U6070 ( .A(n4640), .B(n4639), .ZN(n9858) );
  INV_X1 U6071 ( .A(n9626), .ZN(n4639) );
  AND2_X1 U6072 ( .A1(n4970), .A2(n4971), .ZN(n9635) );
  NAND2_X1 U6073 ( .A1(n9764), .A2(n9244), .ZN(n9751) );
  AND2_X1 U6074 ( .A1(n6524), .A2(n6523), .ZN(n9749) );
  AND2_X1 U6075 ( .A1(n9775), .A2(n9243), .ZN(n9766) );
  INV_X1 U6076 ( .A(n9900), .ZN(n9763) );
  INV_X1 U6077 ( .A(n10072), .ZN(n9842) );
  INV_X1 U6078 ( .A(n9924), .ZN(n9846) );
  INV_X1 U6079 ( .A(n10075), .ZN(n9841) );
  NAND2_X1 U6080 ( .A1(n7770), .A2(n6642), .ZN(n7834) );
  AND2_X1 U6081 ( .A1(n4736), .A2(n4738), .ZN(n7792) );
  OR2_X1 U6082 ( .A1(n7641), .A2(n9677), .ZN(n10075) );
  XNOR2_X1 U6083 ( .A(n7902), .B(n7903), .ZN(n7904) );
  OR2_X1 U6084 ( .A1(n10077), .A2(n7640), .ZN(n10081) );
  INV_X1 U6085 ( .A(n10081), .ZN(n9819) );
  MUX2_X1 U6086 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9851), .S(n10123), .Z(n9854) );
  NOR2_X1 U6087 ( .A1(n9852), .A2(n9921), .ZN(n4634) );
  NAND2_X1 U6088 ( .A1(n5026), .A2(n5025), .ZN(n6977) );
  AOI21_X1 U6089 ( .B1(n5028), .B2(n5030), .A(n4349), .ZN(n5025) );
  NAND2_X1 U6090 ( .A1(n5050), .A2(n6659), .ZN(n9633) );
  INV_X1 U6091 ( .A(n5043), .ZN(n9773) );
  NAND2_X1 U6092 ( .A1(n5041), .A2(n4319), .ZN(n9786) );
  NAND2_X1 U6093 ( .A1(n4730), .A2(n4737), .ZN(n7931) );
  NAND2_X1 U6094 ( .A1(n4735), .A2(n4736), .ZN(n4730) );
  INV_X1 U6095 ( .A(n4729), .ZN(n4735) );
  AND2_X2 U6096 ( .A1(n5620), .A2(n5619), .ZN(n10115) );
  AND2_X1 U6097 ( .A1(n8128), .A2(n6932), .ZN(n9985) );
  INV_X1 U6098 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9989) );
  CLKBUF_X1 U6099 ( .A(n5573), .Z(n8531) );
  INV_X1 U6100 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8199) );
  INV_X1 U6101 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8174) );
  INV_X1 U6102 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8141) );
  INV_X1 U6103 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8130) );
  INV_X1 U6104 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8038) );
  INV_X1 U6105 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8040) );
  INV_X1 U6106 ( .A(n6669), .ZN(n9366) );
  XNOR2_X1 U6107 ( .A(n5505), .B(n5500), .ZN(n7859) );
  INV_X1 U6108 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7394) );
  AND2_X1 U6109 ( .A1(n5466), .A2(n5476), .ZN(n9533) );
  AND2_X1 U6110 ( .A1(n5426), .A2(n5432), .ZN(n7210) );
  INV_X1 U6111 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10359) );
  XNOR2_X1 U6112 ( .A(n5376), .B(n5375), .ZN(n9467) );
  OAI21_X1 U6113 ( .B1(n5366), .B2(n7013), .A(n4684), .ZN(n5367) );
  NAND2_X1 U6114 ( .A1(n5366), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4684) );
  XNOR2_X1 U6115 ( .A(n5356), .B(n5355), .ZN(n7064) );
  NAND2_X1 U6116 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5355) );
  AOI21_X1 U6117 ( .B1(n10019), .B2(n10294), .A(n10018), .ZN(n10383) );
  NOR2_X1 U6118 ( .A1(n10025), .A2(n10024), .ZN(n10220) );
  NOR2_X1 U6119 ( .A1(n10032), .A2(n10031), .ZN(n10214) );
  NOR2_X1 U6120 ( .A1(n10216), .A2(n10215), .ZN(n10031) );
  NOR2_X1 U6121 ( .A1(n10038), .A2(n10037), .ZN(n10210) );
  NAND2_X1 U6122 ( .A1(n4527), .A2(n8679), .ZN(n8259) );
  AND2_X1 U6123 ( .A1(n5016), .A2(n5015), .ZN(n7470) );
  OAI21_X1 U6124 ( .B1(n4557), .B2(n8515), .A(n8514), .ZN(P2_U3296) );
  XNOR2_X1 U6125 ( .A(n4548), .B(n7677), .ZN(n4557) );
  NAND2_X1 U6126 ( .A1(n8767), .A2(n6240), .ZN(n7098) );
  NAND2_X1 U6127 ( .A1(n7165), .A2(n7164), .ZN(n7163) );
  NAND2_X1 U6128 ( .A1(n6271), .A2(n6270), .ZN(n8773) );
  NAND2_X1 U6129 ( .A1(n4494), .A2(n4493), .ZN(n6702) );
  AOI21_X1 U6130 ( .B1(n4756), .B2(n8766), .A(n4753), .ZN(n6330) );
  OAI21_X1 U6131 ( .B1(n9004), .B2(n10148), .A(n4311), .ZN(n8886) );
  NAND2_X1 U6132 ( .A1(n8896), .A2(n4336), .ZN(P2_U3208) );
  AOI21_X1 U6133 ( .B1(n6373), .B2(n10199), .A(n4388), .ZN(n5186) );
  AOI21_X1 U6134 ( .B1(n6348), .B2(n6375), .A(n6374), .ZN(n6376) );
  INV_X1 U6135 ( .A(n5146), .ZN(n5145) );
  NOR2_X1 U6136 ( .A1(n4314), .A2(n4438), .ZN(n4437) );
  OR2_X1 U6137 ( .A1(n5166), .A2(n9921), .ZN(n5176) );
  AND2_X1 U6138 ( .A1(n4796), .A2(n9884), .ZN(n6381) );
  INV_X1 U6139 ( .A(n6673), .ZN(n6674) );
  OAI21_X1 U6140 ( .B1(n8576), .B2(n9927), .A(n6672), .ZN(n6673) );
  NAND2_X1 U6141 ( .A1(n4633), .A2(n4632), .ZN(P1_U3549) );
  AOI21_X1 U6142 ( .B1(n9613), .B2(n4635), .A(n4634), .ZN(n4633) );
  INV_X1 U6143 ( .A(n9854), .ZN(n4632) );
  INV_X1 U6144 ( .A(n9927), .ZN(n4635) );
  OR2_X1 U6145 ( .A1(n5166), .A2(n9975), .ZN(n5171) );
  AND2_X1 U6146 ( .A1(n4796), .A2(n9954), .ZN(n6384) );
  NAND2_X1 U6147 ( .A1(n6716), .A2(n6715), .ZN(P1_U3517) );
  NAND2_X1 U6148 ( .A1(n8260), .A2(n8934), .ZN(n8438) );
  AND4_X2 U6149 ( .A1(n5335), .A2(n5333), .A3(n5334), .A4(n5461), .ZN(n4288)
         );
  NAND2_X1 U6150 ( .A1(n6094), .A2(n10161), .ZN(n8347) );
  NOR2_X1 U6151 ( .A1(n8718), .A2(n5018), .ZN(n4289) );
  AND2_X1 U6152 ( .A1(n4925), .A2(n4926), .ZN(n4290) );
  NAND2_X1 U6153 ( .A1(n5997), .A2(n5996), .ZN(n8457) );
  INV_X1 U6154 ( .A(n8457), .ZN(n4864) );
  OR2_X1 U6155 ( .A1(n6832), .A2(n6831), .ZN(n4292) );
  AND3_X1 U6156 ( .A1(n8320), .A2(n4676), .A3(n4325), .ZN(n4293) );
  NAND2_X1 U6157 ( .A1(n5931), .A2(n5930), .ZN(n9031) );
  INV_X1 U6158 ( .A(n5068), .ZN(n5067) );
  OAI21_X1 U6159 ( .B1(n5069), .B2(n8280), .A(n8472), .ZN(n5068) );
  AND4_X1 U6160 ( .A1(n5858), .A2(n5857), .A3(n5856), .A4(n5855), .ZN(n8178)
         );
  AND2_X1 U6161 ( .A1(n5111), .A2(n5108), .ZN(n4294) );
  NAND2_X1 U6162 ( .A1(n6070), .A2(n4396), .ZN(n4760) );
  NAND2_X1 U6163 ( .A1(n8675), .A2(n8255), .ZN(n4295) );
  AND3_X1 U6164 ( .A1(n9395), .A2(n9396), .A3(n9352), .ZN(n4296) );
  INV_X1 U6165 ( .A(n5664), .ZN(n4464) );
  INV_X1 U6166 ( .A(n9303), .ZN(n4976) );
  AND2_X1 U6167 ( .A1(n9332), .A2(n9322), .ZN(n4297) );
  AND4_X1 U6168 ( .A1(n6452), .A2(n6451), .A3(n6450), .A4(n6449), .ZN(n7530)
         );
  AND2_X1 U6169 ( .A1(n5224), .A2(n5232), .ZN(n4298) );
  AND2_X1 U6170 ( .A1(n8422), .A2(n4324), .ZN(n4299) );
  AND2_X1 U6171 ( .A1(n4368), .A2(n6641), .ZN(n4300) );
  NAND2_X1 U6172 ( .A1(n8415), .A2(n4836), .ZN(n4301) );
  NAND2_X1 U6173 ( .A1(n7848), .A2(n7981), .ZN(n5047) );
  NAND2_X1 U6174 ( .A1(n6148), .A2(n6147), .ZN(n8865) );
  INV_X1 U6175 ( .A(n6837), .ZN(n8045) );
  NAND2_X1 U6176 ( .A1(n5440), .A2(n5439), .ZN(n6837) );
  AND3_X1 U6177 ( .A1(n5387), .A2(n5386), .A3(n5385), .ZN(n10095) );
  INV_X1 U6178 ( .A(n5519), .ZN(n4711) );
  AND2_X1 U6179 ( .A1(n8400), .A2(n8401), .ZN(n8399) );
  INV_X1 U6180 ( .A(n8399), .ZN(n4819) );
  AND2_X1 U6181 ( .A1(n5251), .A2(n5239), .ZN(n4302) );
  AND2_X1 U6182 ( .A1(n4913), .A2(n4405), .ZN(n4303) );
  AND2_X1 U6183 ( .A1(n5630), .A2(n4779), .ZN(n4304) );
  AND2_X1 U6184 ( .A1(n5632), .A2(n4782), .ZN(n4305) );
  AND2_X1 U6185 ( .A1(n6276), .A2(n6319), .ZN(n4306) );
  AND2_X1 U6186 ( .A1(n7554), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4307) );
  AND2_X1 U6187 ( .A1(n6309), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4308) );
  AND2_X1 U6188 ( .A1(n5010), .A2(n5013), .ZN(n4309) );
  AND3_X1 U6189 ( .A1(n4904), .A2(n4905), .A3(n4903), .ZN(n4310) );
  NAND2_X1 U6190 ( .A1(n4410), .A2(n7237), .ZN(n7156) );
  OR2_X1 U6191 ( .A1(n10145), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n4311) );
  NAND2_X1 U6192 ( .A1(n5796), .A2(n5795), .ZN(n7927) );
  INV_X1 U6193 ( .A(n6870), .ZN(n5126) );
  INV_X1 U6194 ( .A(n6416), .ZN(n6582) );
  AND2_X1 U6195 ( .A1(n6645), .A2(n6646), .ZN(n4312) );
  NAND2_X1 U6196 ( .A1(n5552), .A2(n5551), .ZN(n9269) );
  NAND2_X1 U6197 ( .A1(n8051), .A2(n5816), .ZN(n8687) );
  INV_X1 U6198 ( .A(n8307), .ZN(n5065) );
  NAND4_X1 U6199 ( .A1(n5785), .A2(n5784), .A3(n5783), .A4(n5782), .ZN(n8752)
         );
  NAND2_X1 U6200 ( .A1(n9693), .A2(n9675), .ZN(n9654) );
  INV_X1 U6201 ( .A(n8335), .ZN(n8754) );
  AND2_X1 U6202 ( .A1(n4295), .A2(n8430), .ZN(n4313) );
  AND3_X1 U6203 ( .A1(n9416), .A2(n9415), .A3(n9414), .ZN(n4314) );
  INV_X1 U6204 ( .A(n6887), .ZN(n5137) );
  NAND2_X1 U6205 ( .A1(n5549), .A2(n5548), .ZN(n8581) );
  AND2_X1 U6206 ( .A1(n9250), .A2(n9683), .ZN(n9709) );
  OR2_X1 U6207 ( .A1(n9734), .A2(n9078), .ZN(n9249) );
  INV_X1 U6208 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4843) );
  NAND2_X2 U6209 ( .A1(n5595), .A2(n5612), .ZN(n6717) );
  NAND2_X1 U6210 ( .A1(n5468), .A2(n5467), .ZN(n9820) );
  AND2_X1 U6211 ( .A1(n9693), .A2(n5149), .ZN(n4315) );
  AND2_X1 U6212 ( .A1(n5664), .A2(n4627), .ZN(n4316) );
  INV_X1 U6213 ( .A(n8887), .ZN(n8889) );
  AND2_X1 U6214 ( .A1(n8464), .A2(n8463), .ZN(n8887) );
  AND2_X1 U6215 ( .A1(n8478), .A2(n8486), .ZN(n4317) );
  NAND2_X1 U6216 ( .A1(n8884), .A2(n8570), .ZN(n4318) );
  INV_X1 U6217 ( .A(n8624), .ZN(n8911) );
  AND2_X1 U6218 ( .A1(n6005), .A2(n6004), .ZN(n8624) );
  AND2_X1 U6219 ( .A1(n5042), .A2(n5044), .ZN(n4319) );
  NAND2_X1 U6220 ( .A1(n5803), .A2(n7810), .ZN(n4320) );
  NAND2_X1 U6221 ( .A1(n8260), .A2(n8919), .ZN(n4321) );
  NOR2_X1 U6222 ( .A1(n6842), .A2(n6841), .ZN(n4322) );
  OR2_X1 U6223 ( .A1(n9021), .A2(n8920), .ZN(n4323) );
  OR2_X1 U6224 ( .A1(n8644), .A2(n8708), .ZN(n4324) );
  AND3_X1 U6225 ( .A1(n8307), .A2(n8870), .A3(n8306), .ZN(n4325) );
  INV_X1 U6226 ( .A(n9305), .ZN(n5032) );
  INV_X1 U6227 ( .A(n8179), .ZN(n4996) );
  NAND2_X1 U6228 ( .A1(n9839), .A2(n9976), .ZN(n9788) );
  AND2_X1 U6229 ( .A1(n9082), .A2(n6887), .ZN(n4326) );
  AND2_X1 U6230 ( .A1(n9243), .A2(n9239), .ZN(n4327) );
  INV_X1 U6231 ( .A(n9714), .ZN(n9253) );
  OR2_X1 U6232 ( .A1(n9021), .A2(n8738), .ZN(n4328) );
  NAND2_X1 U6233 ( .A1(n4625), .A2(n5562), .ZN(n9274) );
  INV_X1 U6234 ( .A(n8948), .ZN(n8739) );
  AND2_X1 U6235 ( .A1(n5947), .A2(n5946), .ZN(n8948) );
  AND2_X1 U6236 ( .A1(n8385), .A2(n8384), .ZN(n4329) );
  NOR2_X1 U6237 ( .A1(n9230), .A2(n9383), .ZN(n4330) );
  AND2_X1 U6238 ( .A1(n4616), .A2(n5271), .ZN(n4331) );
  NAND2_X1 U6239 ( .A1(n8363), .A2(n8354), .ZN(n4582) );
  XNOR2_X1 U6240 ( .A(n4728), .B(n5032), .ZN(n9853) );
  AND2_X1 U6241 ( .A1(n5010), .A2(n5009), .ZN(n4332) );
  NAND2_X1 U6242 ( .A1(n5349), .A2(n5348), .ZN(n4796) );
  AND2_X1 U6243 ( .A1(n5528), .A2(n5527), .ZN(n9675) );
  INV_X1 U6244 ( .A(n9675), .ZN(n9947) );
  NOR2_X1 U6245 ( .A1(n8809), .A2(n6220), .ZN(n4333) );
  AND2_X1 U6246 ( .A1(n5663), .A2(n5058), .ZN(n4334) );
  AND2_X1 U6247 ( .A1(n4425), .A2(n4423), .ZN(n4335) );
  AND2_X1 U6248 ( .A1(n4648), .A2(n8895), .ZN(n4336) );
  AND2_X1 U6249 ( .A1(n6621), .A2(n6620), .ZN(n9270) );
  INV_X1 U6250 ( .A(n9270), .ZN(n9420) );
  NAND2_X1 U6251 ( .A1(n6848), .A2(n6847), .ZN(n4337) );
  OR2_X1 U6252 ( .A1(n10187), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n4338) );
  NAND2_X1 U6253 ( .A1(n9947), .A2(n9652), .ZN(n9313) );
  AND2_X1 U6254 ( .A1(n5646), .A2(n5645), .ZN(n4339) );
  NAND2_X1 U6255 ( .A1(n8425), .A2(n8424), .ZN(n4340) );
  INV_X1 U6256 ( .A(n6642), .ZN(n5046) );
  AND2_X1 U6257 ( .A1(n5644), .A2(P2_IR_REG_30__SCAN_IN), .ZN(n4341) );
  INV_X1 U6258 ( .A(n5232), .ZN(n4884) );
  AND2_X1 U6259 ( .A1(n9190), .A2(n9195), .ZN(n4342) );
  NAND2_X1 U6260 ( .A1(n8613), .A2(n8933), .ZN(n4343) );
  AND2_X1 U6261 ( .A1(n4317), .A2(n8473), .ZN(n4344) );
  AND2_X1 U6262 ( .A1(n4324), .A2(n8419), .ZN(n4345) );
  INV_X1 U6263 ( .A(n9322), .ZN(n4966) );
  AND2_X1 U6264 ( .A1(n5933), .A2(n5932), .ZN(n8613) );
  AND2_X1 U6265 ( .A1(n6956), .A2(n6955), .ZN(n9332) );
  INV_X1 U6266 ( .A(n9332), .ZN(n4963) );
  INV_X1 U6267 ( .A(n4426), .ZN(n8756) );
  OR2_X1 U6268 ( .A1(n7145), .A2(n6299), .ZN(n4426) );
  AND2_X1 U6269 ( .A1(n5116), .A2(n5114), .ZN(n4346) );
  OR2_X1 U6270 ( .A1(n9750), .A2(n6534), .ZN(n4959) );
  AND2_X1 U6271 ( .A1(n5788), .A2(n8751), .ZN(n4347) );
  INV_X1 U6272 ( .A(n4961), .ZN(n4960) );
  NAND2_X1 U6273 ( .A1(n9401), .A2(n9244), .ZN(n4961) );
  AND2_X1 U6274 ( .A1(n8899), .A2(n8892), .ZN(n4348) );
  NOR2_X1 U6275 ( .A1(n6975), .A2(n8550), .ZN(n4349) );
  NAND2_X1 U6276 ( .A1(n5250), .A2(SI_12_), .ZN(n4350) );
  NAND2_X1 U6277 ( .A1(n4988), .A2(n4987), .ZN(n4986) );
  AND3_X1 U6278 ( .A1(n4291), .A2(n5182), .A3(n5048), .ZN(n4351) );
  INV_X1 U6279 ( .A(n5034), .ZN(n5033) );
  NAND2_X1 U6280 ( .A1(n5035), .A2(n6662), .ZN(n5034) );
  INV_X1 U6281 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6462) );
  INV_X1 U6282 ( .A(n5154), .ZN(n5153) );
  NAND2_X1 U6283 ( .A1(n7751), .A2(n5155), .ZN(n5154) );
  AND2_X1 U6284 ( .A1(n8712), .A2(n8740), .ZN(n4352) );
  INV_X1 U6285 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U6286 ( .A1(n4343), .A2(n8422), .ZN(n4353) );
  NAND2_X1 U6287 ( .A1(n9337), .A2(n9340), .ZN(n9307) );
  INV_X1 U6288 ( .A(n9307), .ZN(n4669) );
  AND2_X1 U6289 ( .A1(n4845), .A2(n4505), .ZN(n4354) );
  AND2_X1 U6290 ( .A1(n6246), .A2(n7154), .ZN(n4355) );
  NAND4_X1 U6291 ( .A1(n8447), .A2(n8446), .A3(n8445), .A4(n4323), .ZN(n4356)
         );
  INV_X1 U6292 ( .A(n6348), .ZN(n8519) );
  NAND2_X1 U6293 ( .A1(n6140), .A2(n6139), .ZN(n6348) );
  AND2_X1 U6294 ( .A1(n5895), .A2(n8743), .ZN(n4357) );
  AND4_X1 U6295 ( .A1(n5048), .A2(n5341), .A3(n5589), .A4(n5345), .ZN(n4358)
         );
  AND2_X1 U6296 ( .A1(n5265), .A2(SI_18_), .ZN(n4359) );
  AND2_X1 U6297 ( .A1(n5693), .A2(n7011), .ZN(n4360) );
  AND3_X1 U6298 ( .A1(n8366), .A2(n8364), .A3(n8363), .ZN(n4361) );
  AND2_X1 U6299 ( .A1(n6131), .A2(n8948), .ZN(n4362) );
  AND2_X1 U6300 ( .A1(n5259), .A2(SI_16_), .ZN(n4363) );
  OR2_X1 U6301 ( .A1(n4329), .A2(n4825), .ZN(n4364) );
  INV_X1 U6302 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7046) );
  AND2_X1 U6303 ( .A1(n9240), .A2(n9241), .ZN(n4365) );
  INV_X1 U6304 ( .A(n4833), .ZN(n4832) );
  OR2_X1 U6305 ( .A1(n4837), .A2(n8423), .ZN(n4833) );
  AND2_X1 U6306 ( .A1(n8355), .A2(n4581), .ZN(n4366) );
  INV_X1 U6307 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5227) );
  INV_X1 U6308 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5679) );
  INV_X1 U6309 ( .A(n5086), .ZN(n5085) );
  NAND2_X1 U6310 ( .A1(n5088), .A2(n4323), .ZN(n5086) );
  INV_X1 U6311 ( .A(n9855), .ZN(n9621) );
  NAND2_X1 U6312 ( .A1(n4898), .A2(n5539), .ZN(n9855) );
  AND2_X1 U6313 ( .A1(n6348), .A2(n8476), .ZN(n4367) );
  INV_X1 U6314 ( .A(n5583), .ZN(n9990) );
  INV_X1 U6315 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5048) );
  INV_X1 U6316 ( .A(n4767), .ZN(n5998) );
  NOR2_X1 U6317 ( .A1(n5989), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n4767) );
  AND2_X1 U6318 ( .A1(n5047), .A2(n6642), .ZN(n4368) );
  OR2_X1 U6319 ( .A1(n8581), .A2(n8550), .ZN(n9336) );
  OAI21_X1 U6320 ( .B1(n9278), .B2(n5046), .A(n7835), .ZN(n5045) );
  AND2_X1 U6321 ( .A1(n9911), .A2(n9815), .ZN(n4369) );
  INV_X1 U6322 ( .A(n7769), .ZN(n8010) );
  NAND2_X1 U6323 ( .A1(n8394), .A2(n4826), .ZN(n4825) );
  NAND2_X1 U6324 ( .A1(n4838), .A2(n8415), .ZN(n4370) );
  AND3_X1 U6325 ( .A1(n9626), .A2(n9636), .A3(n9304), .ZN(n4371) );
  AND3_X1 U6326 ( .A1(n9626), .A2(n9261), .A3(n9636), .ZN(n4372) );
  AND3_X1 U6327 ( .A1(n9332), .A2(n9336), .A3(n9312), .ZN(n4373) );
  NAND2_X1 U6328 ( .A1(n6130), .A2(n8933), .ZN(n4374) );
  AND4_X1 U6329 ( .A1(n5866), .A2(n5865), .A3(n5864), .A4(n5863), .ZN(n8594)
         );
  OR2_X1 U6330 ( .A1(n8675), .A2(n8255), .ZN(n8441) );
  INV_X1 U6331 ( .A(n8441), .ZN(n5089) );
  XOR2_X1 U6332 ( .A(n5059), .B(n5350), .Z(n4375) );
  AND2_X1 U6333 ( .A1(n9220), .A2(n9286), .ZN(n4376) );
  NOR2_X1 U6334 ( .A1(n8716), .A2(n8743), .ZN(n4377) );
  INV_X1 U6335 ( .A(n9783), .ZN(n9906) );
  AND2_X1 U6336 ( .A1(n5485), .A2(n5484), .ZN(n9783) );
  AND2_X1 U6337 ( .A1(n8498), .A2(n8500), .ZN(n4378) );
  OR2_X1 U6338 ( .A1(n5770), .A2(n7353), .ZN(n4379) );
  INV_X1 U6339 ( .A(n8442), .ZN(n5083) );
  AND2_X1 U6340 ( .A1(n8010), .A2(n5152), .ZN(n4380) );
  INV_X1 U6341 ( .A(n4867), .ZN(n4866) );
  NOR2_X1 U6342 ( .A1(n8920), .A2(n8456), .ZN(n4867) );
  AND2_X1 U6343 ( .A1(n4825), .A2(n4822), .ZN(n4381) );
  AND2_X1 U6344 ( .A1(n5736), .A2(n5735), .ZN(n6301) );
  AND2_X1 U6345 ( .A1(n7934), .A2(n9221), .ZN(n4382) );
  AND2_X1 U6346 ( .A1(n4852), .A2(n4374), .ZN(n4383) );
  AND2_X1 U6347 ( .A1(n9621), .A2(n5149), .ZN(n4384) );
  AND2_X1 U6348 ( .A1(n4892), .A2(n4891), .ZN(n4890) );
  INV_X1 U6349 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5646) );
  INV_X1 U6350 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4463) );
  INV_X1 U6351 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5672) );
  INV_X1 U6352 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5022) );
  INV_X1 U6353 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5677) );
  INV_X1 U6354 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5144) );
  NAND2_X1 U6355 ( .A1(n5536), .A2(n5535), .ZN(n9644) );
  INV_X1 U6356 ( .A(n9644), .ZN(n5150) );
  INV_X1 U6357 ( .A(n6132), .ZN(n8260) );
  NAND2_X1 U6358 ( .A1(n7573), .A2(n6107), .ZN(n7518) );
  NAND2_X1 U6359 ( .A1(n7823), .A2(n7751), .ZN(n7750) );
  AND2_X1 U6360 ( .A1(n7823), .A2(n4380), .ZN(n7761) );
  INV_X1 U6361 ( .A(n9383), .ZN(n4682) );
  AND2_X1 U6362 ( .A1(n5694), .A2(n5693), .ZN(n7005) );
  NAND2_X1 U6363 ( .A1(n5109), .A2(n5111), .ZN(n8041) );
  INV_X1 U6364 ( .A(n7606), .ZN(n7020) );
  AND2_X1 U6365 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4385) );
  NAND2_X1 U6366 ( .A1(n4443), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U6367 ( .A1(n4977), .A2(n9195), .ZN(n7815) );
  INV_X1 U6368 ( .A(n7143), .ZN(n4428) );
  AND2_X1 U6369 ( .A1(n7966), .A2(n6216), .ZN(n4386) );
  INV_X1 U6370 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n4919) );
  AND2_X1 U6371 ( .A1(n6263), .A2(n6310), .ZN(n4387) );
  AND2_X1 U6372 ( .A1(n6372), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n4388) );
  XNOR2_X1 U6373 ( .A(n5559), .B(n5558), .ZN(n9988) );
  AND2_X1 U6374 ( .A1(n8249), .A2(n8739), .ZN(n4389) );
  AND2_X1 U6375 ( .A1(n8601), .A2(n5986), .ZN(n4390) );
  XNOR2_X1 U6376 ( .A(n5687), .B(P2_IR_REG_25__SCAN_IN), .ZN(n6047) );
  AND2_X1 U6377 ( .A1(n6068), .A2(n6067), .ZN(n8881) );
  AND2_X1 U6378 ( .A1(n7839), .A2(n9221), .ZN(n7932) );
  AND2_X1 U6379 ( .A1(n4939), .A2(n8789), .ZN(n4391) );
  AND2_X1 U6380 ( .A1(n7823), .A2(n5152), .ZN(n4392) );
  AND2_X1 U6381 ( .A1(n5653), .A2(n5652), .ZN(n8570) );
  INV_X1 U6382 ( .A(n4745), .ZN(n4744) );
  OAI21_X1 U6383 ( .B1(n4746), .B2(n6270), .A(n6274), .ZN(n4745) );
  INV_X1 U6384 ( .A(n6317), .ZN(n8790) );
  NAND2_X1 U6385 ( .A1(n6316), .A2(n8778), .ZN(n6317) );
  INV_X1 U6386 ( .A(n5178), .ZN(n4738) );
  AND2_X1 U6387 ( .A1(n7210), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4393) );
  INV_X1 U6388 ( .A(n9609), .ZN(n9852) );
  NAND2_X1 U6389 ( .A1(n5541), .A2(n5540), .ZN(n9609) );
  OR2_X1 U6390 ( .A1(n9551), .A2(n9536), .ZN(n4394) );
  AND2_X1 U6391 ( .A1(n5041), .A2(n5039), .ZN(n4395) );
  NOR2_X2 U6392 ( .A1(n7844), .A2(n6837), .ZN(n7936) );
  OR2_X1 U6393 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4396) );
  AND2_X1 U6394 ( .A1(n6314), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4397) );
  INV_X1 U6395 ( .A(n4742), .ZN(n4488) );
  NAND2_X1 U6396 ( .A1(n4743), .A2(n8788), .ZN(n4742) );
  OR2_X1 U6397 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4398) );
  AND2_X1 U6398 ( .A1(n9817), .A2(n5156), .ZN(n9744) );
  AND2_X1 U6399 ( .A1(n6172), .A2(n8364), .ZN(n4399) );
  OR2_X1 U6400 ( .A1(n8524), .A2(n8991), .ZN(n4400) );
  NOR2_X1 U6401 ( .A1(n6875), .A2(n5117), .ZN(n4401) );
  OR2_X1 U6402 ( .A1(n9521), .A2(n4666), .ZN(n4665) );
  AND2_X1 U6403 ( .A1(n4470), .A2(n4320), .ZN(n4402) );
  NAND2_X1 U6404 ( .A1(n9660), .A2(n9673), .ZN(n4403) );
  NAND2_X1 U6405 ( .A1(n6341), .A2(n8679), .ZN(n4404) );
  INV_X1 U6406 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4429) );
  INV_X1 U6407 ( .A(n10145), .ZN(n10148) );
  AND2_X1 U6408 ( .A1(n6936), .A2(n6938), .ZN(n9175) );
  NAND2_X1 U6409 ( .A1(n6059), .A2(n6058), .ZN(n8679) );
  INV_X1 U6410 ( .A(n8835), .ZN(n8853) );
  NAND2_X2 U6411 ( .A1(n4457), .A2(n5413), .ZN(n8075) );
  XNOR2_X1 U6412 ( .A(n5421), .B(n5422), .ZN(n7025) );
  INV_X1 U6413 ( .A(n6302), .ZN(n7154) );
  NAND2_X1 U6414 ( .A1(n7306), .A2(n7307), .ZN(n7305) );
  OR2_X1 U6415 ( .A1(n6322), .A2(n8167), .ZN(n4405) );
  OR2_X1 U6416 ( .A1(n6319), .A2(n6318), .ZN(n4406) );
  NAND2_X1 U6417 ( .A1(n4951), .A2(n6421), .ZN(n7664) );
  INV_X1 U6418 ( .A(n7669), .ZN(n4658) );
  XNOR2_X1 U6419 ( .A(n10080), .B(n6725), .ZN(n6627) );
  AND2_X1 U6420 ( .A1(n4911), .A2(n7372), .ZN(n4407) );
  AND2_X1 U6421 ( .A1(n8309), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n4408) );
  OAI21_X1 U6422 ( .B1(n8383), .B2(n5093), .A(n8391), .ZN(n5092) );
  INV_X1 U6423 ( .A(n5092), .ZN(n4585) );
  NAND2_X1 U6424 ( .A1(n4931), .A2(n4930), .ZN(n4409) );
  NAND2_X1 U6425 ( .A1(n4658), .A2(n10095), .ZN(n7897) );
  INV_X1 U6426 ( .A(n7897), .ZN(n4657) );
  AND4_X1 U6427 ( .A1(n6492), .A2(n6491), .A3(n6490), .A4(n6489), .ZN(n9422)
         );
  INV_X1 U6428 ( .A(n9422), .ZN(n4638) );
  AND2_X1 U6429 ( .A1(n4948), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4410) );
  INV_X1 U6430 ( .A(n6307), .ZN(n7367) );
  NAND2_X1 U6431 ( .A1(n4934), .A2(n7328), .ZN(n6307) );
  AND2_X1 U6432 ( .A1(n4784), .A2(n4783), .ZN(n4411) );
  INV_X1 U6433 ( .A(n5013), .ZN(n5011) );
  NAND2_X1 U6434 ( .A1(n5014), .A2(n7352), .ZN(n5013) );
  INV_X1 U6435 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n4771) );
  XNOR2_X1 U6436 ( .A(n5698), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8509) );
  INV_X1 U6437 ( .A(n8509), .ZN(n7677) );
  XOR2_X1 U6438 ( .A(n7113), .B(P2_REG2_REG_12__SCAN_IN), .Z(n4412) );
  NAND2_X1 U6439 ( .A1(n7101), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7100) );
  AND2_X1 U6440 ( .A1(n9677), .A2(n9366), .ZN(n4413) );
  AND2_X1 U6441 ( .A1(n4901), .A2(n7154), .ZN(n4414) );
  AND2_X1 U6442 ( .A1(n9415), .A2(n9349), .ZN(n4415) );
  INV_X1 U6443 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7483) );
  INV_X1 U6444 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n4699) );
  INV_X1 U6445 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n4915) );
  INV_X1 U6446 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4604) );
  INV_X1 U6447 ( .A(n10131), .ZN(n4652) );
  NAND2_X1 U6448 ( .A1(n8865), .A2(n10131), .ZN(n8867) );
  OAI211_X1 U6449 ( .C1(n6331), .C2(n8835), .A(n6330), .B(n4416), .ZN(P2_U3201) );
  NAND2_X1 U6450 ( .A1(n4417), .A2(n8825), .ZN(n4416) );
  XNOR2_X1 U6451 ( .A(n4418), .B(n6329), .ZN(n4417) );
  OR2_X1 U6452 ( .A1(n6682), .A2(n6328), .ZN(n4418) );
  NAND2_X1 U6453 ( .A1(n4433), .A2(n5371), .ZN(n4697) );
  XNOR2_X1 U6454 ( .A(n4433), .B(n5371), .ZN(n6991) );
  NAND2_X1 U6455 ( .A1(n4647), .A2(n5208), .ZN(n4433) );
  NAND3_X1 U6456 ( .A1(n9418), .A2(n4437), .A3(n4434), .ZN(P1_U3242) );
  NAND2_X1 U6457 ( .A1(n4435), .A2(n4415), .ZN(n4434) );
  OAI21_X1 U6458 ( .B1(n4436), .B2(n9348), .A(n9347), .ZN(n4435) );
  NAND2_X1 U6459 ( .A1(n4441), .A2(n7966), .ZN(n4917) );
  NAND2_X1 U6460 ( .A1(n5495), .A2(n5494), .ZN(n5496) );
  NAND4_X1 U6461 ( .A1(n4904), .A2(n4905), .A3(n7244), .A4(n4903), .ZN(n4445)
         );
  NAND2_X1 U6462 ( .A1(n7376), .A2(n4447), .ZN(n6214) );
  NAND3_X1 U6463 ( .A1(n6214), .A2(P2_REG2_REG_9__SCAN_IN), .A3(n7560), .ZN(
        n7558) );
  NAND2_X1 U6464 ( .A1(n6207), .A2(n4286), .ZN(n7169) );
  INV_X1 U6465 ( .A(n6207), .ZN(n4448) );
  NAND2_X1 U6466 ( .A1(n4450), .A2(n4678), .ZN(n9223) );
  NAND2_X1 U6467 ( .A1(n4451), .A2(n4376), .ZN(n4450) );
  NAND2_X1 U6468 ( .A1(n9219), .A2(n9218), .ZN(n4451) );
  NAND2_X1 U6469 ( .A1(n9214), .A2(n9213), .ZN(n9219) );
  NAND2_X1 U6470 ( .A1(n4452), .A2(n4874), .ZN(n4873) );
  NAND2_X1 U6471 ( .A1(n4453), .A2(n4373), .ZN(n4452) );
  NAND2_X1 U6472 ( .A1(n4454), .A2(n9267), .ZN(n4453) );
  NAND2_X1 U6473 ( .A1(n4455), .A2(n4372), .ZN(n4454) );
  NAND2_X1 U6474 ( .A1(n4456), .A2(n9260), .ZN(n4455) );
  NAND3_X1 U6475 ( .A1(n9258), .A2(n9256), .A3(n9257), .ZN(n4456) );
  NAND2_X1 U6476 ( .A1(n9231), .A2(n9827), .ZN(n4804) );
  NAND2_X1 U6477 ( .A1(n4467), .A2(n9271), .ZN(n4466) );
  NAND2_X1 U6478 ( .A1(n9225), .A2(n9224), .ZN(n4467) );
  NOR2_X2 U6479 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5369) );
  NOR2_X2 U6480 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5382) );
  AND4_X2 U6481 ( .A1(n5382), .A2(n5369), .A3(n5024), .A4(n5336), .ZN(n5337)
         );
  INV_X1 U6482 ( .A(n8051), .ZN(n4471) );
  NAND2_X1 U6483 ( .A1(n4476), .A2(n4475), .ZN(n4474) );
  NOR2_X2 U6484 ( .A1(n7697), .A2(n4347), .ZN(n7802) );
  AND3_X2 U6485 ( .A1(n4810), .A2(n4811), .A3(n4808), .ZN(n6052) );
  INV_X1 U6486 ( .A(n7099), .ZN(n4492) );
  NAND2_X1 U6487 ( .A1(n10133), .A2(n6096), .ZN(n7383) );
  NAND2_X1 U6488 ( .A1(n8340), .A2(n8341), .ZN(n7306) );
  INV_X2 U6489 ( .A(n6092), .ZN(n6091) );
  AOI21_X1 U6490 ( .B1(n4496), .B2(n10136), .A(n6169), .ZN(n8529) );
  XNOR2_X1 U6491 ( .A(n4497), .B(n8320), .ZN(n4496) );
  NAND2_X1 U6492 ( .A1(n4499), .A2(n4848), .ZN(n4498) );
  NAND2_X1 U6493 ( .A1(n8021), .A2(n6124), .ZN(n4499) );
  NAND2_X1 U6494 ( .A1(n4511), .A2(n6122), .ZN(n8021) );
  NAND3_X1 U6495 ( .A1(n4503), .A2(n4502), .A3(n4500), .ZN(n9051) );
  OAI21_X2 U6496 ( .B1(n4510), .B2(n8921), .A(n4508), .ZN(n8908) );
  OAI21_X2 U6497 ( .B1(n7518), .B2(n6112), .A(n6111), .ZN(n6115) );
  NAND3_X1 U6498 ( .A1(n4519), .A2(n4518), .A3(n4515), .ZN(n5647) );
  NOR2_X1 U6499 ( .A1(n8657), .A2(n8658), .ZN(n8656) );
  OAI21_X2 U6500 ( .B1(n7505), .B2(n6106), .A(n5190), .ZN(n7573) );
  NAND2_X1 U6501 ( .A1(n4309), .A2(n4534), .ZN(n7698) );
  NAND2_X1 U6502 ( .A1(n8754), .A2(n10154), .ZN(n7307) );
  NAND2_X1 U6503 ( .A1(n4536), .A2(n8353), .ZN(n8361) );
  NAND2_X1 U6504 ( .A1(n8352), .A2(n4537), .ZN(n4536) );
  NAND2_X1 U6505 ( .A1(n4539), .A2(n4538), .ZN(n4537) );
  AND2_X1 U6506 ( .A1(n8346), .A2(n10135), .ZN(n4538) );
  NAND3_X1 U6507 ( .A1(n8440), .A2(n8439), .A3(n8921), .ZN(n4543) );
  NAND2_X1 U6508 ( .A1(n4626), .A2(n4544), .ZN(n8404) );
  NAND2_X1 U6509 ( .A1(n4545), .A2(n4820), .ZN(n4544) );
  NAND2_X1 U6510 ( .A1(n4546), .A2(n8381), .ZN(n4545) );
  NAND2_X1 U6511 ( .A1(n8376), .A2(n8375), .ZN(n4546) );
  NAND3_X1 U6512 ( .A1(n4811), .A2(n4464), .A3(n5672), .ZN(n5817) );
  NAND4_X1 U6513 ( .A1(n8505), .A2(n8506), .A3(n4558), .A4(n4549), .ZN(n4548)
         );
  NAND3_X1 U6514 ( .A1(n4676), .A2(n8490), .A3(n8519), .ZN(n4551) );
  NAND2_X1 U6515 ( .A1(n8335), .A2(n4554), .ZN(n4553) );
  NAND2_X1 U6516 ( .A1(n5404), .A2(n4298), .ZN(n4559) );
  NAND3_X1 U6517 ( .A1(n8404), .A2(n8402), .A3(n8403), .ZN(n4562) );
  NAND2_X1 U6518 ( .A1(n8197), .A2(n8747), .ZN(n8395) );
  NAND2_X1 U6519 ( .A1(n7763), .A2(n4566), .ZN(n4565) );
  NAND2_X2 U6520 ( .A1(n9634), .A2(n9262), .ZN(n9625) );
  NAND2_X2 U6521 ( .A1(n4575), .A2(n9690), .ZN(n9685) );
  NAND2_X1 U6522 ( .A1(n4576), .A2(n9683), .ZN(n4575) );
  INV_X1 U6523 ( .A(n9682), .ZN(n4576) );
  NAND2_X1 U6524 ( .A1(n5079), .A2(n4578), .ZN(n8888) );
  OR2_X1 U6525 ( .A1(n5085), .A2(n5082), .ZN(n4579) );
  NAND3_X1 U6526 ( .A1(n9218), .A2(n9197), .A3(n9207), .ZN(n9374) );
  INV_X1 U6527 ( .A(n4582), .ZN(n6171) );
  NAND2_X2 U6528 ( .A1(n9828), .A2(n6501), .ZN(n9830) );
  NAND3_X1 U6529 ( .A1(n5094), .A2(n4585), .A3(n5091), .ZN(n4584) );
  NAND2_X1 U6530 ( .A1(n4586), .A2(n5380), .ZN(n5216) );
  NAND2_X1 U6531 ( .A1(n4697), .A2(n5211), .ZN(n4586) );
  XNOR2_X1 U6532 ( .A(n5380), .B(n4586), .ZN(n6996) );
  NOR2_X1 U6533 ( .A1(n6117), .A2(n4587), .ZN(n4592) );
  NAND2_X1 U6534 ( .A1(n4588), .A2(n6116), .ZN(n8013) );
  NAND2_X1 U6535 ( .A1(n6115), .A2(n4592), .ZN(n4588) );
  INV_X1 U6536 ( .A(n4590), .ZN(n4589) );
  NAND2_X1 U6537 ( .A1(n4593), .A2(n8475), .ZN(n8392) );
  INV_X1 U6538 ( .A(n7721), .ZN(n8292) );
  AND2_X2 U6539 ( .A1(n4601), .A2(n4599), .ZN(n5347) );
  NAND3_X1 U6540 ( .A1(n4600), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4599) );
  NAND3_X1 U6541 ( .A1(n4604), .A2(n4603), .A3(n4602), .ZN(n4601) );
  NAND2_X1 U6542 ( .A1(n5518), .A2(n4609), .ZN(n4608) );
  AOI21_X1 U6543 ( .B1(n5518), .B2(n5287), .A(n4711), .ZN(n5530) );
  NAND2_X1 U6544 ( .A1(n5481), .A2(n4617), .ZN(n4615) );
  NAND3_X1 U6545 ( .A1(n4890), .A2(n5415), .A3(n4302), .ZN(n4622) );
  OAI21_X1 U6546 ( .B1(n5555), .B2(n5554), .A(n5553), .ZN(n5559) );
  NAND2_X1 U6547 ( .A1(n5325), .A2(n5324), .ZN(n5555) );
  NAND2_X1 U6548 ( .A1(n9272), .A2(n4795), .ZN(n4790) );
  NAND2_X1 U6549 ( .A1(n4895), .A2(n4893), .ZN(n5518) );
  INV_X4 U6550 ( .A(n5347), .ZN(n5352) );
  MUX2_X1 U6551 ( .A(n6985), .B(n6994), .S(n6990), .Z(n5217) );
  BUF_X4 U6552 ( .A(n5352), .Z(n5663) );
  NAND2_X1 U6553 ( .A1(n5244), .A2(n5243), .ZN(n4891) );
  AOI21_X1 U6554 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8794), .A(n8795), .ZN(
        n6219) );
  AOI21_X1 U6555 ( .B1(n4820), .B2(n4381), .A(n4819), .ZN(n4626) );
  NAND2_X2 U6556 ( .A1(n5223), .A2(n5222), .ZN(n5404) );
  NAND2_X1 U6557 ( .A1(n7140), .A2(n6205), .ZN(n8761) );
  NAND2_X1 U6558 ( .A1(n4911), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4910) );
  NAND2_X1 U6559 ( .A1(n4644), .A2(n6305), .ZN(n4911) );
  AOI21_X1 U6560 ( .B1(n7966), .B2(n4919), .A(n4412), .ZN(n4918) );
  NOR2_X1 U6561 ( .A1(n6219), .A2(n6320), .ZN(n6220) );
  NAND2_X1 U6562 ( .A1(n4877), .A2(n4876), .ZN(n5481) );
  OAI22_X1 U6563 ( .A1(n6135), .A2(n6134), .B1(n8570), .B2(n9005), .ZN(n8864)
         );
  OAI22_X2 U6564 ( .A1(n8864), .A2(n6138), .B1(n8736), .B2(n8962), .ZN(n6365)
         );
  OAI21_X1 U6565 ( .B1(n8253), .B2(n8933), .A(n8248), .ZN(n8657) );
  NAND2_X1 U6566 ( .A1(n7662), .A2(n6630), .ZN(n7639) );
  OR2_X2 U6567 ( .A1(n5392), .A2(n4287), .ZN(n5359) );
  NAND2_X1 U6568 ( .A1(n9617), .A2(n9616), .ZN(n4640) );
  XNOR2_X1 U6569 ( .A(n5354), .B(SI_1_), .ZN(n5059) );
  AOI22_X1 U6570 ( .A1(n7337), .A2(n7336), .B1(n7385), .B2(n5768), .ZN(n7221)
         );
  XNOR2_X1 U6571 ( .A(n5695), .B(P2_B_REG_SCAN_IN), .ZN(n5688) );
  NAND2_X1 U6572 ( .A1(n6313), .A2(n4641), .ZN(n8089) );
  NAND2_X1 U6573 ( .A1(n4642), .A2(n8086), .ZN(n4641) );
  INV_X1 U6574 ( .A(n6312), .ZN(n4642) );
  INV_X1 U6575 ( .A(n4890), .ZN(n4889) );
  INV_X1 U6576 ( .A(n8483), .ZN(n8478) );
  AOI21_X1 U6577 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n7235), .A(n7236), .ZN(
        n6306) );
  OAI21_X1 U6578 ( .B1(n6112), .B2(n7705), .A(n7719), .ZN(n6109) );
  INV_X1 U6579 ( .A(n6211), .ZN(n4644) );
  NAND2_X2 U6580 ( .A1(n9101), .A2(n6864), .ZN(n6870) );
  NAND2_X2 U6581 ( .A1(n8131), .A2(n5170), .ZN(n9101) );
  NAND2_X1 U6582 ( .A1(n4917), .A2(n4918), .ZN(n7968) );
  NOR2_X1 U6583 ( .A1(n6688), .A2(n6226), .ZN(n6227) );
  NAND2_X1 U6584 ( .A1(n5206), .A2(n5365), .ZN(n4647) );
  NAND2_X1 U6585 ( .A1(n4656), .A2(n4654), .ZN(n5060) );
  NAND2_X1 U6586 ( .A1(n8321), .A2(n8320), .ZN(n4656) );
  INV_X1 U6587 ( .A(n8526), .ZN(n6187) );
  NOR2_X1 U6588 ( .A1(n4582), .A2(n4694), .ZN(n4693) );
  NAND4_X1 U6589 ( .A1(n5672), .A2(n5677), .A3(n5022), .A4(n5638), .ZN(n4813)
         );
  NAND4_X1 U6590 ( .A1(n5870), .A2(n5900), .A3(n5673), .A4(n5845), .ZN(n4812)
         );
  NAND2_X1 U6591 ( .A1(n8228), .A2(n5080), .ZN(n5079) );
  NAND2_X1 U6592 ( .A1(n10127), .A2(n4693), .ZN(n4692) );
  NAND2_X2 U6593 ( .A1(n5573), .A2(n5574), .ZN(n5372) );
  NAND2_X2 U6594 ( .A1(n4657), .A2(n10101), .ZN(n7898) );
  NAND2_X1 U6595 ( .A1(n8477), .A2(n8478), .ZN(n8504) );
  OAI21_X1 U6596 ( .B1(n8436), .B2(n8435), .A(n8434), .ZN(n8440) );
  AOI21_X1 U6597 ( .B1(n8407), .B2(n6124), .A(n4377), .ZN(n4848) );
  OAI21_X1 U6598 ( .B1(n5347), .B2(P2_DATAO_REG_3__SCAN_IN), .A(n4660), .ZN(
        n5209) );
  INV_X1 U6599 ( .A(n6135), .ZN(n8880) );
  OAI21_X1 U6600 ( .B1(n9480), .B2(n9481), .A(n7055), .ZN(n9499) );
  NOR2_X1 U6601 ( .A1(n7205), .A2(n7061), .ZN(n7195) );
  MUX2_X1 U6602 ( .A(n7048), .B(P1_REG2_REG_1__SCAN_IN), .S(n7064), .Z(n9434)
         );
  OR2_X1 U6603 ( .A1(n5369), .A2(n5578), .ZN(n5384) );
  AOI21_X1 U6604 ( .B1(n4672), .B2(n4671), .A(n4670), .ZN(n4792) );
  NAND2_X2 U6605 ( .A1(n5128), .A2(n5131), .ZN(n9154) );
  NAND2_X1 U6606 ( .A1(n5122), .A2(n5119), .ZN(n9074) );
  NAND2_X1 U6607 ( .A1(n9120), .A2(n6905), .ZN(n9091) );
  NOR2_X1 U6608 ( .A1(n9066), .A2(n9067), .ZN(n9123) );
  INV_X1 U6609 ( .A(n6779), .ZN(n5103) );
  INV_X1 U6610 ( .A(n4799), .ZN(n4672) );
  INV_X1 U6611 ( .A(n4788), .ZN(n4787) );
  NAND2_X1 U6612 ( .A1(n6870), .A2(n5112), .ZN(n5122) );
  NAND2_X1 U6613 ( .A1(n7219), .A2(n4379), .ZN(n7349) );
  NAND2_X1 U6614 ( .A1(n4924), .A2(n4426), .ZN(n4925) );
  XNOR2_X2 U6615 ( .A(n5739), .B(n4844), .ZN(n7143) );
  NAND2_X1 U6616 ( .A1(n7839), .A2(n4382), .ZN(n7933) );
  NAND2_X1 U6617 ( .A1(n6301), .A2(n4927), .ZN(n4923) );
  INV_X1 U6618 ( .A(n4922), .ZN(n7101) );
  INV_X1 U6619 ( .A(n8480), .ZN(n4676) );
  NOR2_X1 U6620 ( .A1(n4712), .A2(n4841), .ZN(n4840) );
  AOI21_X1 U6621 ( .B1(n6368), .B2(n10136), .A(n6367), .ZN(n8516) );
  NAND2_X1 U6622 ( .A1(n5366), .A2(n10359), .ZN(n4700) );
  NAND2_X1 U6623 ( .A1(n4853), .A2(n4854), .ZN(n6135) );
  INV_X1 U6624 ( .A(n4861), .ZN(n4855) );
  NAND2_X1 U6625 ( .A1(n4739), .A2(n6651), .ZN(n9704) );
  NAND2_X1 U6626 ( .A1(n9235), .A2(n9352), .ZN(n4805) );
  NAND2_X1 U6627 ( .A1(n9242), .A2(n9394), .ZN(n4786) );
  INV_X1 U6628 ( .A(n6679), .ZN(n6680) );
  NAND2_X1 U6629 ( .A1(n7988), .A2(n6640), .ZN(n4736) );
  NAND2_X1 U6630 ( .A1(n7902), .A2(n9367), .ZN(n9193) );
  NAND2_X1 U6631 ( .A1(n7412), .A2(n4285), .ZN(n7411) );
  NAND2_X1 U6632 ( .A1(n9663), .A2(n4403), .ZN(n5050) );
  OAI21_X1 U6633 ( .B1(n4873), .B2(n4868), .A(n4669), .ZN(n4872) );
  NAND2_X1 U6634 ( .A1(n5027), .A2(n5031), .ZN(n6664) );
  AOI21_X1 U6635 ( .B1(n9247), .B2(n9251), .A(n9323), .ZN(n9248) );
  OAI22_X1 U6636 ( .A1(n5392), .A2(n7014), .B1(n5052), .B2(n5051), .ZN(n5054)
         );
  NAND2_X1 U6637 ( .A1(n6391), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6507) );
  XNOR2_X1 U6638 ( .A(n5550), .B(n4691), .ZN(n9054) );
  AOI21_X1 U6639 ( .B1(n8487), .B2(n8328), .A(n8327), .ZN(n8483) );
  NOR2_X1 U6640 ( .A1(n4809), .A2(n4813), .ZN(n4808) );
  NOR2_X1 U6641 ( .A1(n5664), .A2(n4812), .ZN(n4810) );
  NAND2_X1 U6642 ( .A1(n7299), .A2(n8345), .ZN(n7298) );
  INV_X1 U6643 ( .A(n4798), .ZN(n4793) );
  NAND2_X1 U6644 ( .A1(n4798), .A2(n4790), .ZN(n4789) );
  NAND2_X1 U6645 ( .A1(n4800), .A2(n4796), .ZN(n4795) );
  NAND2_X1 U6646 ( .A1(n5273), .A2(n4896), .ZN(n4895) );
  OR2_X1 U6647 ( .A1(n5061), .A2(n8324), .ZN(n4776) );
  NAND2_X1 U6648 ( .A1(n9054), .A2(n8310), .ZN(n6151) );
  OAI21_X2 U6649 ( .B1(n9625), .B2(n4966), .A(n4964), .ZN(n6957) );
  NAND2_X1 U6650 ( .A1(n4717), .A2(n4715), .ZN(n9682) );
  NAND2_X1 U6651 ( .A1(n9615), .A2(n9611), .ZN(n9851) );
  OAI21_X1 U6652 ( .B1(n4885), .B2(n4884), .A(n5238), .ZN(n4882) );
  OAI22_X1 U6653 ( .A1(n7274), .A2(n7275), .B1(n6091), .B2(n5753), .ZN(n7337)
         );
  NAND2_X1 U6654 ( .A1(n8173), .A2(n5688), .ZN(n5694) );
  OAI21_X1 U6655 ( .B1(n8573), .B2(n4704), .A(n8572), .ZN(P2_U3154) );
  NAND2_X1 U6656 ( .A1(n4705), .A2(n8679), .ZN(n4704) );
  NAND2_X1 U6657 ( .A1(n8567), .A2(n8566), .ZN(n4705) );
  NAND2_X1 U6658 ( .A1(n4899), .A2(n7173), .ZN(n4905) );
  INV_X2 U6659 ( .A(n5761), .ZN(n6161) );
  INV_X1 U6660 ( .A(n9132), .ZN(n5100) );
  NAND2_X1 U6661 ( .A1(n9133), .A2(n5099), .ZN(n5098) );
  NAND2_X1 U6662 ( .A1(n5231), .A2(n5232), .ZN(n4713) );
  NAND3_X1 U6663 ( .A1(n9775), .A2(n9709), .A3(n4718), .ZN(n4717) );
  AND2_X4 U6664 ( .A1(n4726), .A2(n6394), .ZN(n6588) );
  AND4_X2 U6665 ( .A1(n6441), .A2(n6440), .A3(n6438), .A4(n6439), .ZN(n7647)
         );
  NAND4_X1 U6666 ( .A1(n4288), .A2(n4741), .A3(n5337), .A4(n4291), .ZN(n5344)
         );
  AND4_X2 U6667 ( .A1(n5144), .A2(n5494), .A3(n5565), .A4(n5597), .ZN(n5182)
         );
  NAND2_X2 U6668 ( .A1(n4763), .A2(n4764), .ZN(n9064) );
  NAND2_X1 U6669 ( .A1(n4761), .A2(n4762), .ZN(n6237) );
  NAND3_X1 U6670 ( .A1(n4764), .A2(n4763), .A3(P2_REG2_REG_1__SCAN_IN), .ZN(
        n4762) );
  NAND3_X1 U6671 ( .A1(n7483), .A2(n4775), .A3(n5624), .ZN(n5781) );
  NAND2_X1 U6672 ( .A1(n5631), .A2(n4777), .ZN(n5904) );
  NAND2_X1 U6673 ( .A1(n5633), .A2(n4780), .ZN(n5940) );
  NAND2_X1 U6674 ( .A1(n5636), .A2(n4411), .ZN(n6141) );
  NAND2_X1 U6675 ( .A1(n5636), .A2(n5635), .ZN(n6016) );
  AOI21_X1 U6676 ( .B1(n4786), .B2(n4296), .A(n4365), .ZN(n9251) );
  NAND2_X1 U6677 ( .A1(n9238), .A2(n4327), .ZN(n9242) );
  NOR2_X1 U6678 ( .A1(n4800), .A2(n4796), .ZN(n4797) );
  AOI21_X1 U6679 ( .B1(n4804), .B2(n4330), .A(n9386), .ZN(n4803) );
  OR2_X1 U6680 ( .A1(n5561), .A2(n6989), .ZN(n5358) );
  NAND2_X2 U6681 ( .A1(n5372), .A2(n6990), .ZN(n5561) );
  NAND2_X1 U6682 ( .A1(n5343), .A2(n5577), .ZN(n5573) );
  NAND2_X1 U6683 ( .A1(n4806), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5342) );
  NAND3_X1 U6684 ( .A1(n5337), .A2(n4288), .A3(n4807), .ZN(n4806) );
  NAND4_X1 U6685 ( .A1(n4291), .A2(n4288), .A3(n5142), .A4(n5182), .ZN(n5593)
         );
  NAND2_X1 U6686 ( .A1(n5639), .A2(n5896), .ZN(n4809) );
  MUX2_X1 U6687 ( .A(n4429), .B(n4814), .S(n5754), .Z(n8334) );
  NAND3_X1 U6688 ( .A1(n8387), .A2(n8385), .A3(n8395), .ZN(n4822) );
  INV_X1 U6689 ( .A(n8391), .ZN(n4828) );
  NAND2_X1 U6690 ( .A1(n8416), .A2(n4835), .ZN(n4834) );
  NAND2_X1 U6691 ( .A1(n6048), .A2(n4839), .ZN(n5691) );
  INV_X1 U6692 ( .A(n5691), .ZN(n5658) );
  OAI21_X1 U6693 ( .B1(n8361), .B2(n7382), .A(n4361), .ZN(n8371) );
  INV_X2 U6694 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4844) );
  OR2_X1 U6695 ( .A1(n5755), .A2(n6236), .ZN(n6205) );
  OR2_X1 U6696 ( .A1(n5755), .A2(n10187), .ZN(n6298) );
  INV_X1 U6697 ( .A(n7306), .ZN(n8345) );
  NAND2_X1 U6698 ( .A1(n8942), .A2(n4851), .ZN(n4850) );
  INV_X1 U6699 ( .A(n4852), .ZN(n8945) );
  NAND2_X1 U6700 ( .A1(n5449), .A2(n4878), .ZN(n4877) );
  NAND2_X1 U6701 ( .A1(n5449), .A2(n5254), .ZN(n5458) );
  NAND2_X1 U6702 ( .A1(n7154), .A2(n4900), .ZN(n4904) );
  INV_X1 U6703 ( .A(n7173), .ZN(n4900) );
  NAND2_X1 U6704 ( .A1(n7173), .A2(n6209), .ZN(n4901) );
  AOI21_X1 U6705 ( .B1(n7173), .B2(n6209), .A(n6302), .ZN(n4902) );
  NAND3_X1 U6706 ( .A1(n4905), .A2(n4904), .A3(n4906), .ZN(n7155) );
  NAND2_X1 U6707 ( .A1(n7154), .A2(n4907), .ZN(n4906) );
  INV_X1 U6708 ( .A(n6209), .ZN(n4907) );
  NAND2_X1 U6709 ( .A1(n4910), .A2(n7372), .ZN(n6212) );
  INV_X1 U6710 ( .A(n8821), .ZN(n4916) );
  AND2_X1 U6711 ( .A1(n6214), .A2(n7560), .ZN(n7605) );
  NAND2_X1 U6712 ( .A1(n7558), .A2(n7560), .ZN(n4921) );
  INV_X1 U6713 ( .A(n6322), .ZN(n4929) );
  NAND2_X1 U6714 ( .A1(n8823), .A2(n8824), .ZN(n8822) );
  NAND2_X1 U6715 ( .A1(n7555), .A2(n7554), .ZN(n4930) );
  NAND3_X1 U6716 ( .A1(n4930), .A2(n6311), .A3(n4931), .ZN(n6312) );
  NAND3_X1 U6717 ( .A1(n4932), .A2(n6309), .A3(n4307), .ZN(n4931) );
  INV_X1 U6718 ( .A(n6308), .ZN(n4933) );
  NAND2_X1 U6719 ( .A1(n6306), .A2(n6305), .ZN(n4937) );
  INV_X1 U6720 ( .A(n6306), .ZN(n4934) );
  INV_X1 U6721 ( .A(n4936), .ZN(n7366) );
  NAND2_X1 U6722 ( .A1(n6317), .A2(n4942), .ZN(n4939) );
  NAND2_X1 U6723 ( .A1(n8790), .A2(n8789), .ZN(n4940) );
  INV_X1 U6724 ( .A(n8789), .ZN(n4941) );
  NAND2_X1 U6725 ( .A1(n4943), .A2(n6317), .ZN(n8779) );
  NAND3_X1 U6726 ( .A1(n4943), .A2(n6317), .A3(P2_REG1_REG_13__SCAN_IN), .ZN(
        n4942) );
  AOI21_X1 U6727 ( .B1(n6303), .B2(n4947), .A(n4945), .ZN(n7236) );
  NAND2_X1 U6728 ( .A1(n8347), .A2(n8348), .ZN(n10126) );
  INV_X1 U6729 ( .A(n8320), .ZN(n8308) );
  INV_X1 U6730 ( .A(n8508), .ZN(n5061) );
  NAND2_X2 U6731 ( .A1(n5819), .A2(n5818), .ZN(n6113) );
  NAND3_X1 U6732 ( .A1(n4950), .A2(n4949), .A3(n6428), .ZN(n7644) );
  NAND3_X1 U6733 ( .A1(n4952), .A2(n9369), .A3(n4953), .ZN(n4949) );
  NAND3_X1 U6734 ( .A1(n7416), .A2(n4952), .A3(n9369), .ZN(n4950) );
  NAND2_X2 U6735 ( .A1(n4977), .A2(n4342), .ZN(n9372) );
  NAND2_X1 U6736 ( .A1(n4982), .A2(n4981), .ZN(n4984) );
  NAND3_X1 U6737 ( .A1(n6337), .A2(n6336), .A3(n4983), .ZN(n4982) );
  INV_X1 U6738 ( .A(n4982), .ZN(n8573) );
  OAI211_X1 U6739 ( .C1(n4982), .C2(n4404), .A(n4984), .B(n6349), .ZN(P2_U3160) );
  NAND2_X1 U6740 ( .A1(n6336), .A2(n6337), .ZN(n8567) );
  INV_X1 U6741 ( .A(n8566), .ZN(n4983) );
  INV_X1 U6742 ( .A(n5192), .ZN(n4993) );
  NAND2_X1 U6743 ( .A1(n4997), .A2(n5844), .ZN(n8177) );
  NAND2_X1 U6744 ( .A1(n5983), .A2(n5982), .ZN(n8680) );
  NAND2_X1 U6745 ( .A1(n5983), .A2(n4999), .ZN(n4998) );
  INV_X1 U6746 ( .A(n6008), .ZN(n5005) );
  NAND3_X1 U6747 ( .A1(n5008), .A2(n5012), .A3(n5007), .ZN(n5010) );
  INV_X1 U6748 ( .A(n7471), .ZN(n5007) );
  NAND2_X1 U6749 ( .A1(n7350), .A2(n5015), .ZN(n5008) );
  NOR2_X1 U6750 ( .A1(n7699), .A2(n5011), .ZN(n5009) );
  INV_X1 U6751 ( .A(n5016), .ZN(n7348) );
  NAND2_X1 U6752 ( .A1(n5871), .A2(n5021), .ZN(n5020) );
  NAND3_X1 U6753 ( .A1(n5382), .A2(n5369), .A3(n5024), .ZN(n5398) );
  NAND2_X1 U6754 ( .A1(n6663), .A2(n5028), .ZN(n5026) );
  NAND2_X1 U6755 ( .A1(n6663), .A2(n5033), .ZN(n5027) );
  OR2_X1 U6756 ( .A1(n9820), .A2(n9833), .ZN(n5044) );
  INV_X1 U6757 ( .A(n9363), .ZN(n6750) );
  NAND2_X2 U6758 ( .A1(n5370), .A2(n5053), .ZN(n9363) );
  NAND3_X1 U6759 ( .A1(n6172), .A2(n8364), .A3(n6175), .ZN(n6178) );
  NAND3_X1 U6760 ( .A1(n4287), .A2(n6990), .A3(n5754), .ZN(n5056) );
  INV_X1 U6761 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5058) );
  NAND2_X1 U6762 ( .A1(n6161), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5721) );
  OAI21_X1 U6763 ( .B1(n8878), .B2(n5068), .A(n5064), .ZN(n6369) );
  NAND2_X1 U6764 ( .A1(n8289), .A2(n8385), .ZN(n5093) );
  OAI21_X1 U6765 ( .B1(n7517), .B2(n8289), .A(n8385), .ZN(n7704) );
  INV_X1 U6766 ( .A(n8385), .ZN(n5096) );
  NAND2_X1 U6767 ( .A1(n6737), .A2(n5097), .ZN(n7423) );
  NAND3_X1 U6768 ( .A1(n5098), .A2(n5101), .A3(n6786), .ZN(n7525) );
  NAND2_X1 U6769 ( .A1(n5102), .A2(n6779), .ZN(n5101) );
  INV_X1 U6770 ( .A(n6771), .ZN(n5102) );
  NAND2_X2 U6771 ( .A1(n6720), .A2(n6717), .ZN(n6911) );
  XNOR2_X1 U6772 ( .A(n5570), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U6773 ( .A1(n8261), .A2(n4322), .ZN(n5106) );
  AOI21_X2 U6774 ( .B1(n5109), .B2(n5107), .A(n5105), .ZN(n8133) );
  NAND2_X2 U6775 ( .A1(n7974), .A2(n5110), .ZN(n5109) );
  AND2_X1 U6776 ( .A1(n5115), .A2(n6875), .ZN(n5114) );
  AOI21_X1 U6777 ( .B1(n6875), .B2(n5121), .A(n5120), .ZN(n5119) );
  INV_X1 U6778 ( .A(n9162), .ZN(n5123) );
  OR2_X1 U6779 ( .A1(n6872), .A2(n6873), .ZN(n5127) );
  NAND2_X1 U6780 ( .A1(n9073), .A2(n5129), .ZN(n5128) );
  INV_X1 U6781 ( .A(n9082), .ZN(n5138) );
  NAND3_X1 U6782 ( .A1(n5142), .A2(n4288), .A3(n5143), .ZN(n5141) );
  OAI21_X1 U6783 ( .B1(n5148), .B2(n5147), .A(n5145), .ZN(P1_U3240) );
  AOI21_X1 U6784 ( .B1(n9090), .B2(n8272), .A(n8271), .ZN(n5147) );
  NAND2_X1 U6785 ( .A1(n8273), .A2(n9175), .ZN(n5148) );
  NAND2_X1 U6786 ( .A1(n5161), .A2(n6712), .ZN(n5160) );
  NAND2_X1 U6787 ( .A1(n5162), .A2(n5166), .ZN(n5164) );
  NAND2_X1 U6788 ( .A1(n6712), .A2(n5163), .ZN(n5162) );
  INV_X1 U6789 ( .A(n9274), .ZN(n5166) );
  OR2_X2 U6790 ( .A1(n6970), .A2(n9269), .ZN(n6971) );
  NAND2_X1 U6791 ( .A1(n6362), .A2(n10184), .ZN(n6199) );
  NAND2_X1 U6792 ( .A1(n6957), .A2(n6955), .ZN(n6614) );
  NAND2_X1 U6793 ( .A1(n8516), .A2(n6371), .ZN(n6373) );
  OR2_X1 U6794 ( .A1(n5684), .A2(n5683), .ZN(n5685) );
  INV_X1 U6795 ( .A(n7005), .ZN(n7006) );
  NAND2_X1 U6796 ( .A1(n5685), .A2(n5686), .ZN(n5695) );
  INV_X4 U6797 ( .A(n5392), .ZN(n5560) );
  NAND2_X1 U6798 ( .A1(n5674), .A2(n5183), .ZN(n5859) );
  NAND2_X1 U6799 ( .A1(n6047), .A2(n6046), .ZN(n6230) );
  OR2_X1 U6800 ( .A1(n8324), .A2(n6158), .ZN(n6191) );
  INV_X1 U6801 ( .A(n5585), .ZN(n6394) );
  OR2_X1 U6802 ( .A1(n8542), .A2(n9980), .ZN(n6982) );
  OR2_X1 U6803 ( .A1(n8542), .A2(n9927), .ZN(n6978) );
  NAND2_X1 U6804 ( .A1(n8565), .A2(n8554), .ZN(n8563) );
  NAND2_X1 U6805 ( .A1(n5596), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U6806 ( .A1(n9051), .A2(n9055), .ZN(n5742) );
  OR2_X1 U6807 ( .A1(n6382), .A2(n6381), .ZN(P1_U3552) );
  OR2_X1 U6808 ( .A1(n6385), .A2(n6384), .ZN(P1_U3520) );
  NAND2_X1 U6809 ( .A1(n5570), .A2(n5565), .ZN(n5566) );
  INV_X1 U6810 ( .A(n8581), .ZN(n6975) );
  INV_X1 U6811 ( .A(n6666), .ZN(n8036) );
  CLKBUF_X1 U6812 ( .A(n5574), .Z(n9999) );
  INV_X1 U6813 ( .A(n9414), .ZN(n9349) );
  OAI21_X1 U6814 ( .B1(n6968), .B2(n9797), .A(n6967), .ZN(n8539) );
  AND2_X2 U6815 ( .A1(n6361), .A2(n7302), .ZN(n10199) );
  INV_X1 U6816 ( .A(n10199), .ZN(n6372) );
  AND2_X1 U6817 ( .A1(n10141), .A2(n10172), .ZN(n10180) );
  AND2_X1 U6818 ( .A1(n4400), .A2(n6363), .ZN(n5167) );
  INV_X1 U6819 ( .A(n5742), .ZN(n5851) );
  INV_X1 U6820 ( .A(n8613), .ZN(n6130) );
  OR2_X1 U6821 ( .A1(n9644), .A2(n9627), .ZN(n5168) );
  AND2_X1 U6822 ( .A1(n8408), .A2(n8407), .ZN(n5169) );
  OR2_X1 U6823 ( .A1(n6853), .A2(n6852), .ZN(n5170) );
  INV_X1 U6824 ( .A(n8407), .ZN(n6123) );
  INV_X1 U6825 ( .A(n8550), .ZN(n9421) );
  AND2_X1 U6826 ( .A1(n8499), .A2(n6167), .ZN(n10131) );
  INV_X1 U6827 ( .A(n7113), .ZN(n6314) );
  AND2_X1 U6828 ( .A1(n8870), .A2(n8469), .ZN(n5172) );
  OR2_X1 U6829 ( .A1(n8519), .A2(n8991), .ZN(n5173) );
  AND2_X1 U6830 ( .A1(n5175), .A2(n6198), .ZN(n5174) );
  OR2_X1 U6831 ( .A1(n8524), .A2(n9044), .ZN(n5175) );
  NOR2_X1 U6832 ( .A1(n6636), .A2(n7747), .ZN(n5177) );
  NOR2_X1 U6833 ( .A1(n6639), .A2(n7791), .ZN(n5178) );
  AND2_X1 U6834 ( .A1(n8203), .A2(n5695), .ZN(n5179) );
  AND3_X1 U6835 ( .A1(n6023), .A2(n6333), .A3(n8618), .ZN(n5180) );
  NOR2_X1 U6836 ( .A1(n9619), .A2(n9618), .ZN(n5181) );
  AND2_X1 U6837 ( .A1(n5845), .A2(n5673), .ZN(n5183) );
  NAND2_X1 U6838 ( .A1(n5839), .A2(n8747), .ZN(n6108) );
  INV_X1 U6839 ( .A(n9031), .ZN(n6131) );
  AND2_X1 U6840 ( .A1(n9705), .A2(n9703), .ZN(n5184) );
  OR2_X2 U6841 ( .A1(n9732), .A2(n9734), .ZN(n5185) );
  NAND2_X1 U6842 ( .A1(n10184), .A2(n10157), .ZN(n9044) );
  INV_X1 U6843 ( .A(n9044), .ZN(n6375) );
  NAND2_X1 U6844 ( .A1(n6951), .A2(n9930), .ZN(n9186) );
  INV_X1 U6845 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5260) );
  INV_X1 U6846 ( .A(n9729), .ZN(n9687) );
  AND2_X2 U6847 ( .A1(n8128), .A2(n6984), .ZN(P1_U3973) );
  INV_X1 U6848 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5489) );
  NAND2_X2 U6849 ( .A1(n7641), .A2(n10072), .ZN(n9848) );
  OR2_X1 U6850 ( .A1(n9259), .A2(n9271), .ZN(n5187) );
  NAND2_X1 U6851 ( .A1(n5568), .A2(n5567), .ZN(n5596) );
  NAND2_X2 U6852 ( .A1(n7314), .A2(n10129), .ZN(n10145) );
  AND2_X1 U6853 ( .A1(n9104), .A2(n9103), .ZN(n5189) );
  NOR2_X1 U6854 ( .A1(n6816), .A2(n7881), .ZN(n5191) );
  AND2_X1 U6855 ( .A1(n8691), .A2(n5838), .ZN(n5192) );
  AND2_X1 U6856 ( .A1(n8369), .A2(n8368), .ZN(n8370) );
  NAND2_X1 U6857 ( .A1(n8360), .A2(n8499), .ZN(n8374) );
  AND2_X1 U6858 ( .A1(n8412), .A2(n8411), .ZN(n8413) );
  AND2_X1 U6859 ( .A1(n8460), .A2(n8459), .ZN(n8461) );
  AND2_X1 U6860 ( .A1(n8461), .A2(n8887), .ZN(n8462) );
  INV_X1 U6861 ( .A(n8747), .ZN(n5836) );
  AND2_X1 U6862 ( .A1(n7015), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6300) );
  OR2_X1 U6863 ( .A1(n5313), .A2(n5546), .ZN(n5315) );
  NAND2_X1 U6864 ( .A1(n5837), .A2(n5836), .ZN(n5838) );
  NAND2_X1 U6865 ( .A1(n6727), .A2(n6726), .ZN(n6728) );
  INV_X1 U6866 ( .A(n7385), .ZN(n6094) );
  NOR2_X1 U6867 ( .A1(n8884), .A2(n8891), .ZN(n6134) );
  INV_X1 U6868 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5624) );
  NOR2_X1 U6869 ( .A1(n9102), .A2(n9100), .ZN(n6863) );
  OR2_X1 U6870 ( .A1(n6919), .A2(n7425), .ZN(n6736) );
  INV_X1 U6871 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n10361) );
  INV_X1 U6872 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5578) );
  NOR2_X1 U6873 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5338) );
  AND2_X1 U6874 ( .A1(n5517), .A2(n5520), .ZN(n5287) );
  INV_X1 U6875 ( .A(n5508), .ZN(n5277) );
  INV_X1 U6876 ( .A(SI_17_), .ZN(n10264) );
  NAND2_X1 U6877 ( .A1(n7339), .A2(n7385), .ZN(n8348) );
  INV_X1 U6878 ( .A(n10180), .ZN(n6186) );
  INV_X1 U6879 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6399) );
  INV_X1 U6880 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6525) );
  INV_X1 U6881 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6512) );
  INV_X1 U6882 ( .A(n6959), .ZN(n6618) );
  NOR2_X1 U6883 ( .A1(n6965), .A2(n9277), .ZN(n6966) );
  NAND2_X1 U6884 ( .A1(n6669), .A2(n6666), .ZN(n9344) );
  INV_X1 U6885 ( .A(n7936), .ZN(n8102) );
  NAND2_X1 U6886 ( .A1(n5577), .A2(n5576), .ZN(n5581) );
  NAND2_X1 U6887 ( .A1(n5268), .A2(n5267), .ZN(n5272) );
  INV_X1 U6888 ( .A(SI_12_), .ZN(n10251) );
  XNOR2_X1 U6889 ( .A(n5903), .B(n7419), .ZN(n5769) );
  INV_X1 U6890 ( .A(n6026), .ZN(n8618) );
  AND2_X1 U6891 ( .A1(n8369), .A2(n8366), .ZN(n8285) );
  NOR2_X1 U6892 ( .A1(n8499), .A2(n6352), .ZN(n7303) );
  AND2_X1 U6893 ( .A1(n7007), .A2(n6074), .ZN(n6359) );
  OR2_X1 U6894 ( .A1(n7449), .A2(n6185), .ZN(n10141) );
  AND2_X1 U6895 ( .A1(n6192), .A2(n6191), .ZN(n6193) );
  OR2_X1 U6896 ( .A1(n6878), .A2(n6877), .ZN(n6879) );
  AND3_X1 U6897 ( .A1(n5588), .A2(n5587), .A3(n5586), .ZN(n9273) );
  INV_X1 U6898 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7079) );
  OR2_X1 U6899 ( .A1(n7035), .A2(n7034), .ZN(n9588) );
  INV_X1 U6900 ( .A(n9627), .ZN(n9653) );
  NAND2_X1 U6901 ( .A1(n6653), .A2(n6652), .ZN(n9691) );
  INV_X1 U6902 ( .A(n9864), .ZN(n9894) );
  NAND2_X1 U6903 ( .A1(n9221), .A2(n9222), .ZN(n7835) );
  NAND2_X1 U6904 ( .A1(n7031), .A2(n9455), .ZN(n9800) );
  OR2_X1 U6905 ( .A1(n6943), .A2(n5611), .ZN(n7631) );
  INV_X1 U6906 ( .A(n8724), .ZN(n8704) );
  OAI21_X1 U6907 ( .B1(n9005), .B2(n8731), .A(n6087), .ZN(n6088) );
  NAND2_X1 U6908 ( .A1(n6061), .A2(n10129), .ZN(n8711) );
  INV_X1 U6909 ( .A(n8846), .ZN(n8764) );
  INV_X1 U6910 ( .A(n8510), .ZN(n6296) );
  INV_X1 U6911 ( .A(n8088), .ZN(n8848) );
  INV_X1 U6912 ( .A(n8958), .ZN(n8927) );
  INV_X1 U6913 ( .A(n10129), .ZN(n8954) );
  INV_X1 U6914 ( .A(n8991), .ZN(n8983) );
  INV_X1 U6915 ( .A(n8304), .ZN(n8230) );
  NAND2_X1 U6916 ( .A1(n6057), .A2(n8337), .ZN(n10178) );
  INV_X1 U6917 ( .A(n10178), .ZN(n10157) );
  OR2_X1 U6918 ( .A1(n6194), .A2(n6193), .ZN(n6195) );
  INV_X1 U6919 ( .A(n6081), .ZN(n7007) );
  INV_X1 U6920 ( .A(n8264), .ZN(n9177) );
  INV_X1 U6921 ( .A(n9186), .ZN(n9168) );
  INV_X1 U6922 ( .A(n9164), .ZN(n9183) );
  AND3_X1 U6923 ( .A1(n6964), .A2(n6963), .A3(n6962), .ZN(n9277) );
  INV_X1 U6924 ( .A(n6665), .ZN(n9677) );
  INV_X1 U6925 ( .A(n9800), .ZN(n9836) );
  INV_X1 U6926 ( .A(n9850), .ZN(n9700) );
  AND2_X1 U6927 ( .A1(n10123), .A2(n9930), .ZN(n9884) );
  OAI21_X1 U6928 ( .B1(n8576), .B2(n9980), .A(n6678), .ZN(n6679) );
  INV_X1 U6929 ( .A(n10112), .ZN(n9916) );
  INV_X1 U6930 ( .A(n9230), .ZN(n9831) );
  OR2_X1 U6931 ( .A1(n9352), .A2(n9349), .ZN(n9933) );
  INV_X1 U6932 ( .A(n9986), .ZN(n5619) );
  XNOR2_X1 U6933 ( .A(n5594), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5599) );
  INV_X1 U6934 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10294) );
  NOR2_X1 U6935 ( .A1(n10222), .A2(n10221), .ZN(n10024) );
  INV_X1 U6936 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10310) );
  INV_X1 U6937 ( .A(n8679), .ZN(n8717) );
  INV_X1 U6938 ( .A(n8711), .ZN(n8731) );
  INV_X1 U6939 ( .A(n8570), .ZN(n8891) );
  INV_X1 U6940 ( .A(n8178), .ZN(n8745) );
  NAND2_X1 U6941 ( .A1(P2_U3893), .A2(n6296), .ZN(n8850) );
  NAND2_X1 U6942 ( .A1(n7253), .A2(n6228), .ZN(n8835) );
  NAND2_X1 U6943 ( .A1(n10145), .A2(n7459), .ZN(n8958) );
  NAND2_X1 U6944 ( .A1(n10199), .A2(n6186), .ZN(n8986) );
  INV_X1 U6945 ( .A(n8675), .ZN(n9028) );
  NAND2_X1 U6946 ( .A1(n10184), .A2(n6186), .ZN(n9039) );
  INV_X2 U6947 ( .A(n10186), .ZN(n10184) );
  INV_X1 U6948 ( .A(n7023), .ZN(n7024) );
  INV_X1 U6949 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n10375) );
  INV_X1 U6950 ( .A(n8086), .ZN(n7044) );
  NAND2_X1 U6951 ( .A1(n7265), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9164) );
  INV_X1 U6952 ( .A(n9175), .ZN(n9170) );
  INV_X1 U6953 ( .A(n6909), .ZN(n9637) );
  INV_X1 U6954 ( .A(n10061), .ZN(n9561) );
  OR2_X1 U6955 ( .A1(n10077), .A2(n7638), .ZN(n9850) );
  NAND2_X1 U6956 ( .A1(n10123), .A2(n10112), .ZN(n9927) );
  INV_X1 U6957 ( .A(n9660), .ZN(n9944) );
  INV_X1 U6958 ( .A(n9820), .ZN(n9976) );
  NAND2_X1 U6959 ( .A1(n10115), .A2(n10112), .ZN(n9980) );
  INV_X1 U6960 ( .A(n10115), .ZN(n10113) );
  INV_X1 U6961 ( .A(n10086), .ZN(n10087) );
  AND2_X1 U6962 ( .A1(n9985), .A2(n9983), .ZN(n10086) );
  INV_X1 U6963 ( .A(n5599), .ZN(n8143) );
  INV_X1 U6964 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7680) );
  INV_X1 U6965 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7043) );
  NOR2_X1 U6966 ( .A1(n10015), .A2(n10014), .ZN(n10385) );
  AOI21_X1 U6967 ( .B1(n10027), .B2(n10286), .A(n10026), .ZN(n10218) );
  INV_X2 U6968 ( .A(n8742), .ZN(P2_U3893) );
  INV_X1 U6969 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n5617) );
  INV_X1 U6970 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7013) );
  NAND2_X1 U6971 ( .A1(n5352), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5193) );
  INV_X1 U6972 ( .A(SI_2_), .ZN(n5364) );
  OAI211_X1 U6973 ( .C1(n5352), .C2(n7013), .A(n5193), .B(n5364), .ZN(n5206)
         );
  AND2_X1 U6974 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5351) );
  INV_X1 U6975 ( .A(n5351), .ZN(n5194) );
  INV_X1 U6976 ( .A(SI_1_), .ZN(n5199) );
  NAND2_X1 U6977 ( .A1(n5194), .A2(n5199), .ZN(n5195) );
  NAND2_X1 U6978 ( .A1(n5195), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U6979 ( .A1(n5351), .A2(SI_1_), .ZN(n5196) );
  NAND2_X1 U6980 ( .A1(n5197), .A2(n5196), .ZN(n5198) );
  NAND2_X1 U6981 ( .A1(n5352), .A2(n5198), .ZN(n5205) );
  NAND2_X1 U6982 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6983 ( .A1(n5353), .A2(n5199), .ZN(n5200) );
  NAND2_X1 U6984 ( .A1(n5200), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5202) );
  NAND3_X1 U6985 ( .A1(SI_1_), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n5201) );
  NAND2_X1 U6986 ( .A1(n5202), .A2(n5201), .ZN(n5203) );
  NAND2_X1 U6987 ( .A1(n5347), .A2(n5203), .ZN(n5204) );
  INV_X1 U6988 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6988) );
  NAND2_X1 U6989 ( .A1(n5352), .A2(n6988), .ZN(n5207) );
  OAI211_X1 U6990 ( .C1(n5352), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n5207), .B(
        SI_2_), .ZN(n5208) );
  INV_X1 U6991 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6987) );
  INV_X1 U6992 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6992) );
  INV_X1 U6993 ( .A(n5209), .ZN(n5210) );
  NAND2_X1 U6994 ( .A1(n5210), .A2(SI_3_), .ZN(n5211) );
  INV_X1 U6995 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6997) );
  INV_X1 U6996 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6986) );
  XNOR2_X1 U6997 ( .A(n5213), .B(SI_4_), .ZN(n5380) );
  INV_X1 U6998 ( .A(n5213), .ZN(n5214) );
  NAND2_X1 U6999 ( .A1(n5214), .A2(SI_4_), .ZN(n5215) );
  NAND2_X1 U7000 ( .A1(n5216), .A2(n5215), .ZN(n5390) );
  INV_X1 U7001 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6994) );
  INV_X1 U7002 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6985) );
  XNOR2_X1 U7003 ( .A(n5217), .B(SI_5_), .ZN(n5391) );
  NAND2_X1 U7004 ( .A1(n5390), .A2(n5391), .ZN(n5220) );
  INV_X1 U7005 ( .A(n5217), .ZN(n5218) );
  NAND2_X1 U7006 ( .A1(n5218), .A2(SI_5_), .ZN(n5219) );
  MUX2_X1 U7007 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5663), .Z(n5221) );
  INV_X1 U7008 ( .A(SI_6_), .ZN(n10340) );
  XNOR2_X1 U7009 ( .A(n5221), .B(n10340), .ZN(n5395) );
  NAND2_X1 U7010 ( .A1(n5397), .A2(n5395), .ZN(n5223) );
  NAND2_X1 U7011 ( .A1(n5221), .A2(SI_6_), .ZN(n5222) );
  XNOR2_X1 U7012 ( .A(n5225), .B(SI_7_), .ZN(n5403) );
  INV_X1 U7013 ( .A(n5403), .ZN(n5224) );
  NAND2_X1 U7014 ( .A1(n5225), .A2(SI_7_), .ZN(n5226) );
  INV_X1 U7015 ( .A(SI_8_), .ZN(n5228) );
  NAND2_X1 U7016 ( .A1(n5229), .A2(n5228), .ZN(n5232) );
  INV_X1 U7017 ( .A(n5229), .ZN(n5230) );
  NAND2_X1 U7018 ( .A1(n5230), .A2(SI_8_), .ZN(n5231) );
  INV_X1 U7019 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5233) );
  MUX2_X1 U7020 ( .A(n7022), .B(n5233), .S(n5366), .Z(n5235) );
  INV_X1 U7021 ( .A(SI_9_), .ZN(n5234) );
  NAND2_X1 U7022 ( .A1(n5235), .A2(n5234), .ZN(n5239) );
  INV_X1 U7023 ( .A(n5235), .ZN(n5236) );
  NAND2_X1 U7024 ( .A1(n5236), .A2(SI_9_), .ZN(n5237) );
  NAND2_X1 U7025 ( .A1(n5239), .A2(n5237), .ZN(n5414) );
  INV_X1 U7026 ( .A(n5414), .ZN(n5238) );
  INV_X1 U7027 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5240) );
  MUX2_X1 U7028 ( .A(n7027), .B(n5240), .S(n5663), .Z(n5241) );
  XNOR2_X1 U7029 ( .A(n5241), .B(SI_10_), .ZN(n5422) );
  INV_X1 U7030 ( .A(n5422), .ZN(n5244) );
  INV_X1 U7031 ( .A(n5241), .ZN(n5242) );
  NAND2_X1 U7032 ( .A1(n5242), .A2(SI_10_), .ZN(n5243) );
  INV_X1 U7033 ( .A(SI_11_), .ZN(n5245) );
  NAND2_X1 U7034 ( .A1(n5246), .A2(n5245), .ZN(n5249) );
  INV_X1 U7035 ( .A(n5246), .ZN(n5247) );
  NAND2_X1 U7036 ( .A1(n5247), .A2(SI_11_), .ZN(n5248) );
  NAND2_X1 U7037 ( .A1(n5249), .A2(n5248), .ZN(n5429) );
  MUX2_X1 U7038 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n5663), .Z(n5250) );
  XNOR2_X1 U7039 ( .A(n5250), .B(n10251), .ZN(n5436) );
  MUX2_X1 U7040 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5663), .Z(n5252) );
  XNOR2_X1 U7041 ( .A(n5252), .B(SI_13_), .ZN(n5441) );
  INV_X1 U7042 ( .A(n5441), .ZN(n5251) );
  NAND2_X1 U7043 ( .A1(n5252), .A2(SI_13_), .ZN(n5253) );
  MUX2_X1 U7044 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n5366), .Z(n5255) );
  XNOR2_X1 U7045 ( .A(n5255), .B(SI_14_), .ZN(n5448) );
  INV_X1 U7046 ( .A(n5448), .ZN(n5254) );
  NAND2_X1 U7047 ( .A1(n5255), .A2(SI_14_), .ZN(n5457) );
  MUX2_X1 U7048 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n5366), .Z(n5459) );
  NAND2_X1 U7049 ( .A1(n5459), .A2(SI_15_), .ZN(n5469) );
  MUX2_X1 U7050 ( .A(n10323), .B(n7394), .S(n5663), .Z(n5473) );
  INV_X1 U7051 ( .A(n5459), .ZN(n5257) );
  INV_X1 U7052 ( .A(SI_15_), .ZN(n5256) );
  NAND2_X1 U7053 ( .A1(n5257), .A2(n5256), .ZN(n5470) );
  OAI21_X1 U7054 ( .B1(SI_16_), .B2(n5259), .A(n5470), .ZN(n5258) );
  MUX2_X1 U7055 ( .A(n7398), .B(n5260), .S(n5366), .Z(n5261) );
  INV_X1 U7056 ( .A(n5261), .ZN(n5262) );
  NAND2_X1 U7057 ( .A1(n5262), .A2(SI_17_), .ZN(n5263) );
  NAND2_X1 U7058 ( .A1(n5264), .A2(n5263), .ZN(n5480) );
  MUX2_X1 U7059 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5366), .Z(n5265) );
  XNOR2_X1 U7060 ( .A(n5265), .B(n10300), .ZN(n5486) );
  INV_X1 U7061 ( .A(n5486), .ZN(n5266) );
  MUX2_X1 U7062 ( .A(n7678), .B(n7680), .S(n5663), .Z(n5268) );
  INV_X1 U7063 ( .A(n5268), .ZN(n5269) );
  NAND2_X1 U7064 ( .A1(n5269), .A2(SI_19_), .ZN(n5270) );
  NAND2_X1 U7065 ( .A1(n5272), .A2(n5270), .ZN(n5492) );
  INV_X1 U7066 ( .A(n5492), .ZN(n5271) );
  MUX2_X1 U7067 ( .A(n7861), .B(n7787), .S(n5366), .Z(n5503) );
  INV_X1 U7068 ( .A(n5503), .ZN(n5276) );
  MUX2_X1 U7069 ( .A(n8575), .B(n8040), .S(n5663), .Z(n5508) );
  OAI22_X1 U7070 ( .A1(SI_20_), .A2(n5276), .B1(n5277), .B2(SI_21_), .ZN(n5280) );
  INV_X1 U7071 ( .A(SI_21_), .ZN(n5274) );
  OAI21_X1 U7072 ( .B1(n5503), .B2(n5504), .A(n5274), .ZN(n5278) );
  AND2_X1 U7073 ( .A1(SI_21_), .A2(SI_20_), .ZN(n5275) );
  AOI22_X1 U7074 ( .A1(n5278), .A2(n5277), .B1(n5276), .B2(n5275), .ZN(n5279)
         );
  MUX2_X1 U7075 ( .A(n8035), .B(n8038), .S(n5663), .Z(n5282) );
  INV_X1 U7076 ( .A(SI_22_), .ZN(n5281) );
  NAND2_X1 U7077 ( .A1(n5282), .A2(n5281), .ZN(n5517) );
  INV_X1 U7078 ( .A(n5282), .ZN(n5283) );
  NAND2_X1 U7079 ( .A1(n5283), .A2(SI_22_), .ZN(n5284) );
  NAND2_X1 U7080 ( .A1(n5517), .A2(n5284), .ZN(n5513) );
  INV_X1 U7081 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5285) );
  MUX2_X1 U7082 ( .A(n5285), .B(n8130), .S(n5366), .Z(n5288) );
  INV_X1 U7083 ( .A(SI_23_), .ZN(n5286) );
  NAND2_X1 U7084 ( .A1(n5288), .A2(n5286), .ZN(n5520) );
  INV_X1 U7085 ( .A(n5288), .ZN(n5289) );
  NAND2_X1 U7086 ( .A1(n5289), .A2(SI_23_), .ZN(n5519) );
  MUX2_X1 U7087 ( .A(n8140), .B(n8141), .S(n5663), .Z(n5291) );
  INV_X1 U7088 ( .A(SI_24_), .ZN(n5290) );
  NAND2_X1 U7089 ( .A1(n5291), .A2(n5290), .ZN(n5294) );
  INV_X1 U7090 ( .A(n5291), .ZN(n5292) );
  NAND2_X1 U7091 ( .A1(n5292), .A2(SI_24_), .ZN(n5293) );
  MUX2_X1 U7092 ( .A(n8172), .B(n8174), .S(n5366), .Z(n5296) );
  INV_X1 U7093 ( .A(SI_25_), .ZN(n5295) );
  NAND2_X1 U7094 ( .A1(n5296), .A2(n5295), .ZN(n5299) );
  INV_X1 U7095 ( .A(n5296), .ZN(n5297) );
  NAND2_X1 U7096 ( .A1(n5297), .A2(SI_25_), .ZN(n5298) );
  INV_X1 U7097 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8201) );
  MUX2_X1 U7098 ( .A(n8201), .B(n8199), .S(n5663), .Z(n5302) );
  INV_X1 U7099 ( .A(SI_26_), .ZN(n5301) );
  NAND2_X1 U7100 ( .A1(n5302), .A2(n5301), .ZN(n5305) );
  INV_X1 U7101 ( .A(n5302), .ZN(n5303) );
  NAND2_X1 U7102 ( .A1(n5303), .A2(SI_26_), .ZN(n5304) );
  INV_X1 U7103 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10001) );
  MUX2_X1 U7104 ( .A(n10375), .B(n10001), .S(n5366), .Z(n5307) );
  INV_X1 U7105 ( .A(SI_27_), .ZN(n5306) );
  NAND2_X1 U7106 ( .A1(n5307), .A2(n5306), .ZN(n5544) );
  INV_X1 U7107 ( .A(n5307), .ZN(n5308) );
  NAND2_X1 U7108 ( .A1(n5308), .A2(SI_27_), .ZN(n5309) );
  INV_X1 U7109 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5310) );
  INV_X1 U7110 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8532) );
  MUX2_X1 U7111 ( .A(n5310), .B(n8532), .S(n5663), .Z(n5312) );
  INV_X1 U7112 ( .A(SI_28_), .ZN(n5311) );
  NAND2_X1 U7113 ( .A1(n5312), .A2(n5311), .ZN(n5316) );
  INV_X1 U7114 ( .A(n5316), .ZN(n5313) );
  XNOR2_X1 U7115 ( .A(n5312), .B(SI_28_), .ZN(n5546) );
  AND2_X1 U7116 ( .A1(n5542), .A2(n5315), .ZN(n5314) );
  INV_X1 U7117 ( .A(n5315), .ZN(n5318) );
  AND2_X1 U7118 ( .A1(n5544), .A2(n5316), .ZN(n5317) );
  MUX2_X1 U7119 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n5663), .Z(n5322) );
  NAND2_X1 U7120 ( .A1(n5550), .A2(SI_29_), .ZN(n5325) );
  AND2_X1 U7121 ( .A1(n5321), .A2(n5320), .ZN(n5323) );
  NAND2_X1 U7122 ( .A1(n5323), .A2(n5322), .ZN(n5324) );
  INV_X1 U7123 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n5326) );
  INV_X1 U7124 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8590) );
  MUX2_X1 U7125 ( .A(n5326), .B(n8590), .S(n5366), .Z(n5328) );
  INV_X1 U7126 ( .A(SI_30_), .ZN(n5327) );
  NAND2_X1 U7127 ( .A1(n5328), .A2(n5327), .ZN(n5553) );
  INV_X1 U7128 ( .A(n5328), .ZN(n5329) );
  NAND2_X1 U7129 ( .A1(n5329), .A2(SI_30_), .ZN(n5330) );
  NAND2_X1 U7130 ( .A1(n5553), .A2(n5330), .ZN(n5554) );
  NOR2_X1 U7131 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5332) );
  NOR2_X1 U7132 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5335) );
  INV_X1 U7133 ( .A(n5582), .ZN(n5577) );
  INV_X1 U7134 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U7135 ( .A1(n5344), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U7136 ( .A1(n8588), .A2(n5560), .ZN(n5349) );
  OR2_X1 U7137 ( .A1(n5561), .A2(n8590), .ZN(n5348) );
  MUX2_X1 U7138 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5663), .Z(n5350) );
  NAND2_X1 U7139 ( .A1(n5352), .A2(n5351), .ZN(n5362) );
  OAI21_X1 U7140 ( .B1(n5366), .B2(n5353), .A(n5362), .ZN(n5354) );
  INV_X1 U7141 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6989) );
  INV_X1 U7142 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5356) );
  OR2_X1 U7143 ( .A1(n5372), .A2(n7064), .ZN(n5357) );
  AND3_X4 U7144 ( .A1(n5358), .A2(n5359), .A3(n5357), .ZN(n10080) );
  INV_X1 U7145 ( .A(SI_0_), .ZN(n5361) );
  INV_X1 U7146 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5360) );
  OAI21_X1 U7147 ( .B1(n6990), .B2(n5361), .A(n5360), .ZN(n5363) );
  AND2_X1 U7148 ( .A1(n5363), .A2(n5362), .ZN(n10003) );
  MUX2_X1 U7149 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10003), .S(n5372), .Z(n7651)
         );
  NAND2_X1 U7150 ( .A1(n10080), .A2(n7425), .ZN(n7413) );
  XNOR2_X1 U7151 ( .A(n5365), .B(n5364), .ZN(n5368) );
  XNOR2_X1 U7152 ( .A(n5368), .B(n5367), .ZN(n7014) );
  INV_X1 U7153 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5373) );
  XNOR2_X1 U7154 ( .A(n5384), .B(n5373), .ZN(n9446) );
  OR2_X1 U7155 ( .A1(n5372), .A2(n9446), .ZN(n5370) );
  NOR2_X2 U7156 ( .A1(n7413), .A2(n9363), .ZN(n7670) );
  OR2_X1 U7157 ( .A1(n5392), .A2(n6991), .ZN(n5379) );
  OR2_X1 U7158 ( .A1(n5561), .A2(n6987), .ZN(n5378) );
  NAND2_X1 U7159 ( .A1(n5384), .A2(n5373), .ZN(n5374) );
  NAND2_X1 U7160 ( .A1(n5374), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5376) );
  INV_X1 U7161 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5375) );
  OR2_X1 U7162 ( .A1(n5372), .A2(n9467), .ZN(n5377) );
  NAND2_X1 U7163 ( .A1(n7670), .A2(n10089), .ZN(n7669) );
  INV_X1 U7164 ( .A(n6996), .ZN(n5381) );
  NAND2_X1 U7165 ( .A1(n5560), .A2(n5381), .ZN(n5387) );
  OR2_X1 U7166 ( .A1(n5382), .A2(n5489), .ZN(n5383) );
  NAND2_X1 U7167 ( .A1(n5384), .A2(n5383), .ZN(n5388) );
  OR2_X1 U7168 ( .A1(n5372), .A2(n10055), .ZN(n5386) );
  OR2_X1 U7169 ( .A1(n5561), .A2(n6986), .ZN(n5385) );
  INV_X1 U7170 ( .A(n10095), .ZN(n9134) );
  INV_X2 U7171 ( .A(n5561), .ZN(n5499) );
  OAI21_X1 U7172 ( .B1(n5388), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5389) );
  XNOR2_X1 U7173 ( .A(n5389), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9482) );
  AOI22_X1 U7174 ( .A1(n5499), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5052), .B2(
        n9482), .ZN(n5394) );
  XNOR2_X1 U7175 ( .A(n5390), .B(n5391), .ZN(n6993) );
  OR2_X1 U7176 ( .A1(n6993), .A2(n5392), .ZN(n5393) );
  INV_X1 U7177 ( .A(n5395), .ZN(n5396) );
  XNOR2_X1 U7178 ( .A(n5397), .B(n5396), .ZN(n6998) );
  NAND2_X1 U7179 ( .A1(n6998), .A2(n5560), .ZN(n5402) );
  NAND2_X1 U7180 ( .A1(n5398), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5399) );
  MUX2_X1 U7181 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5399), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5400) );
  AND2_X1 U7182 ( .A1(n5400), .A2(n5408), .ZN(n9503) );
  AOI22_X1 U7183 ( .A1(n5499), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5052), .B2(
        n9503), .ZN(n5401) );
  NAND2_X1 U7184 ( .A1(n5402), .A2(n5401), .ZN(n9199) );
  NOR2_X4 U7185 ( .A1(n7898), .A2(n9199), .ZN(n7823) );
  XNOR2_X1 U7186 ( .A(n5404), .B(n5403), .ZN(n7002) );
  NAND2_X1 U7187 ( .A1(n7002), .A2(n5560), .ZN(n5407) );
  NAND2_X1 U7188 ( .A1(n5408), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5405) );
  XNOR2_X1 U7189 ( .A(n5405), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7121) );
  AOI22_X1 U7190 ( .A1(n5499), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5052), .B2(
        n7121), .ZN(n5406) );
  NAND2_X1 U7191 ( .A1(n5407), .A2(n5406), .ZN(n7911) );
  INV_X1 U7192 ( .A(n7911), .ZN(n7751) );
  NOR2_X1 U7193 ( .A1(n5424), .A2(n5489), .ZN(n5409) );
  NAND2_X1 U7194 ( .A1(n5409), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5412) );
  INV_X1 U7195 ( .A(n5409), .ZN(n5411) );
  NAND2_X1 U7196 ( .A1(n5411), .A2(n5410), .ZN(n5417) );
  AOI22_X1 U7197 ( .A1(n5499), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5052), .B2(
        n7137), .ZN(n5413) );
  NAND2_X1 U7198 ( .A1(n4883), .A2(n5414), .ZN(n5416) );
  NAND2_X1 U7199 ( .A1(n5416), .A2(n5415), .ZN(n7018) );
  NAND2_X1 U7200 ( .A1(n7018), .A2(n5560), .ZN(n5420) );
  NAND2_X1 U7201 ( .A1(n5417), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5418) );
  XNOR2_X1 U7202 ( .A(n5418), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7092) );
  AOI22_X1 U7203 ( .A1(n5499), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5052), .B2(
        n7092), .ZN(n5419) );
  NAND2_X1 U7204 ( .A1(n5420), .A2(n5419), .ZN(n7875) );
  NAND2_X1 U7205 ( .A1(n7025), .A2(n5560), .ZN(n5428) );
  NAND2_X1 U7206 ( .A1(n5482), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5425) );
  MUX2_X1 U7207 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5425), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n5426) );
  AOI22_X1 U7208 ( .A1(n5499), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5052), .B2(
        n7210), .ZN(n5427) );
  NAND2_X1 U7209 ( .A1(n5428), .A2(n5427), .ZN(n7769) );
  NAND2_X1 U7210 ( .A1(n7042), .A2(n5560), .ZN(n5435) );
  NAND2_X1 U7211 ( .A1(n5432), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5431) );
  MUX2_X1 U7212 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5431), .S(
        P1_IR_REG_11__SCAN_IN), .Z(n5433) );
  INV_X1 U7213 ( .A(n5444), .ZN(n5437) );
  NAND2_X1 U7214 ( .A1(n5433), .A2(n5437), .ZN(n7192) );
  INV_X1 U7215 ( .A(n7192), .ZN(n7081) );
  AOI22_X1 U7216 ( .A1(n5499), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5052), .B2(
        n7081), .ZN(n5434) );
  INV_X1 U7217 ( .A(n6484), .ZN(n7848) );
  NAND2_X1 U7218 ( .A1(n5437), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5438) );
  XNOR2_X1 U7219 ( .A(n5438), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7280) );
  AOI22_X1 U7220 ( .A1(n5499), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5052), .B2(
        n7280), .ZN(n5439) );
  XNOR2_X1 U7221 ( .A(n5442), .B(n5441), .ZN(n7227) );
  NAND2_X1 U7222 ( .A1(n7227), .A2(n5560), .ZN(n5447) );
  INV_X1 U7223 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U7224 ( .A1(n5444), .A2(n5443), .ZN(n5450) );
  NAND2_X1 U7225 ( .A1(n5450), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5445) );
  XNOR2_X1 U7226 ( .A(n5445), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9518) );
  AOI22_X1 U7227 ( .A1(n5052), .A2(n9518), .B1(n5499), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n5446) );
  XNOR2_X1 U7228 ( .A(n5449), .B(n5448), .ZN(n7319) );
  NAND2_X1 U7229 ( .A1(n7319), .A2(n5560), .ZN(n5456) );
  INV_X1 U7230 ( .A(n5450), .ZN(n5452) );
  INV_X1 U7231 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5451) );
  INV_X1 U7232 ( .A(n5462), .ZN(n5453) );
  NAND2_X1 U7233 ( .A1(n5453), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5454) );
  XNOR2_X1 U7234 ( .A(n5454), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7320) );
  AOI22_X1 U7235 ( .A1(n7320), .A2(n5052), .B1(n5499), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n5455) );
  XNOR2_X1 U7236 ( .A(n5459), .B(SI_15_), .ZN(n5460) );
  NAND2_X1 U7237 ( .A1(n7345), .A2(n5560), .ZN(n5468) );
  AOI21_X1 U7238 ( .B1(n5462), .B2(n5461), .A(n5489), .ZN(n5463) );
  NAND2_X1 U7239 ( .A1(n5463), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n5466) );
  INV_X1 U7240 ( .A(n5463), .ZN(n5465) );
  INV_X1 U7241 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U7242 ( .A1(n5465), .A2(n5464), .ZN(n5476) );
  AOI22_X1 U7243 ( .A1(n9533), .A2(n5052), .B1(n5499), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n5467) );
  INV_X1 U7244 ( .A(n5469), .ZN(n5471) );
  OAI21_X1 U7245 ( .B1(n5472), .B2(n5471), .A(n5470), .ZN(n5475) );
  XNOR2_X1 U7246 ( .A(n5473), .B(SI_16_), .ZN(n5474) );
  XNOR2_X1 U7247 ( .A(n5475), .B(n5474), .ZN(n7393) );
  NAND2_X1 U7248 ( .A1(n7393), .A2(n5560), .ZN(n5479) );
  NAND2_X1 U7249 ( .A1(n5476), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5477) );
  XNOR2_X1 U7250 ( .A(n5477), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9535) );
  AOI22_X1 U7251 ( .A1(n9535), .A2(n5052), .B1(n5499), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n5478) );
  XNOR2_X1 U7252 ( .A(n5481), .B(n5480), .ZN(n7396) );
  NAND2_X1 U7253 ( .A1(n7396), .A2(n5560), .ZN(n5485) );
  NAND2_X1 U7254 ( .A1(n5141), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5483) );
  XNOR2_X1 U7255 ( .A(n5483), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9568) );
  AOI22_X1 U7256 ( .A1(n5499), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5052), .B2(
        n9568), .ZN(n5484) );
  XNOR2_X1 U7257 ( .A(n5487), .B(n5486), .ZN(n7495) );
  NAND2_X1 U7258 ( .A1(n7495), .A2(n5560), .ZN(n5491) );
  XNOR2_X1 U7259 ( .A(n5495), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9583) );
  AOI22_X1 U7260 ( .A1(n5499), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5052), .B2(
        n9583), .ZN(n5490) );
  XNOR2_X1 U7261 ( .A(n5493), .B(n5492), .ZN(n7676) );
  NAND2_X1 U7262 ( .A1(n7676), .A2(n5560), .ZN(n6524) );
  XNOR2_X2 U7263 ( .A(n5498), .B(n5497), .ZN(n6665) );
  AOI22_X1 U7264 ( .A1(n9677), .A2(n5052), .B1(n5499), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n6523) );
  NAND2_X1 U7265 ( .A1(n9744), .A2(n9749), .ZN(n9732) );
  XNOR2_X1 U7266 ( .A(n5503), .B(SI_20_), .ZN(n5500) );
  NAND2_X1 U7267 ( .A1(n7859), .A2(n5560), .ZN(n5502) );
  OR2_X1 U7268 ( .A1(n5561), .A2(n7787), .ZN(n5501) );
  NAND2_X1 U7269 ( .A1(n5505), .A2(n5504), .ZN(n5506) );
  NAND2_X1 U7270 ( .A1(n5507), .A2(n5506), .ZN(n5510) );
  XNOR2_X1 U7271 ( .A(n5508), .B(SI_21_), .ZN(n5509) );
  NAND2_X1 U7272 ( .A1(n8039), .A2(n5560), .ZN(n5512) );
  OR2_X1 U7273 ( .A1(n5561), .A2(n8040), .ZN(n5511) );
  NOR2_X2 U7274 ( .A1(n5185), .A2(n9955), .ZN(n9717) );
  XNOR2_X1 U7275 ( .A(n5514), .B(n5513), .ZN(n8034) );
  NAND2_X1 U7276 ( .A1(n8034), .A2(n5560), .ZN(n5516) );
  OR2_X1 U7277 ( .A1(n5561), .A2(n8038), .ZN(n5515) );
  AND2_X1 U7278 ( .A1(n5518), .A2(n5517), .ZN(n5521) );
  NAND2_X1 U7279 ( .A1(n5520), .A2(n5519), .ZN(n5522) );
  NAND2_X1 U7280 ( .A1(n5521), .A2(n5522), .ZN(n5526) );
  INV_X1 U7281 ( .A(n5521), .ZN(n5524) );
  INV_X1 U7282 ( .A(n5522), .ZN(n5523) );
  NAND2_X1 U7283 ( .A1(n5524), .A2(n5523), .ZN(n5525) );
  NAND2_X1 U7284 ( .A1(n5526), .A2(n5525), .ZN(n8127) );
  NAND2_X1 U7285 ( .A1(n8127), .A2(n5560), .ZN(n5528) );
  OR2_X1 U7286 ( .A1(n5561), .A2(n8130), .ZN(n5527) );
  XNOR2_X1 U7287 ( .A(n5530), .B(n5529), .ZN(n8139) );
  NAND2_X1 U7288 ( .A1(n8139), .A2(n5560), .ZN(n5532) );
  OR2_X1 U7289 ( .A1(n5561), .A2(n8141), .ZN(n5531) );
  NAND2_X1 U7290 ( .A1(n8171), .A2(n5560), .ZN(n5536) );
  OR2_X1 U7291 ( .A1(n5561), .A2(n8174), .ZN(n5535) );
  OR2_X1 U7292 ( .A1(n5561), .A2(n8199), .ZN(n5539) );
  NAND2_X1 U7293 ( .A1(n9061), .A2(n5560), .ZN(n5541) );
  OR2_X1 U7294 ( .A1(n5561), .A2(n10001), .ZN(n5540) );
  AND2_X2 U7295 ( .A1(n6710), .A2(n9852), .ZN(n6712) );
  NAND2_X1 U7296 ( .A1(n8530), .A2(n5560), .ZN(n5549) );
  OR2_X1 U7297 ( .A1(n5561), .A2(n8532), .ZN(n5548) );
  NAND2_X1 U7298 ( .A1(n9054), .A2(n5560), .ZN(n5552) );
  INV_X1 U7299 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9997) );
  OR2_X1 U7300 ( .A1(n5561), .A2(n9997), .ZN(n5551) );
  INV_X1 U7301 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5556) );
  INV_X1 U7302 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9994) );
  MUX2_X1 U7303 ( .A(n5556), .B(n9994), .S(n5663), .Z(n5557) );
  XNOR2_X1 U7304 ( .A(n5557), .B(SI_31_), .ZN(n5558) );
  OR2_X1 U7305 ( .A1(n5561), .A2(n9994), .ZN(n5562) );
  AND2_X2 U7306 ( .A1(n5569), .A2(n5596), .ZN(n6666) );
  INV_X1 U7307 ( .A(n9999), .ZN(n9452) );
  NAND2_X1 U7308 ( .A1(n9452), .A2(P1_B_REG_SCAN_IN), .ZN(n5575) );
  NAND2_X1 U7309 ( .A1(n9834), .A2(n5575), .ZN(n6965) );
  NAND2_X1 U7310 ( .A1(n5579), .A2(n5578), .ZN(n5580) );
  NAND2_X1 U7311 ( .A1(n5582), .A2(n5579), .ZN(n5583) );
  XNOR2_X2 U7312 ( .A(n5584), .B(n9989), .ZN(n5585) );
  NAND2_X1 U7313 ( .A1(n6959), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5588) );
  AND2_X2 U7314 ( .A1(n9996), .A2(n6394), .ZN(n6423) );
  INV_X2 U7315 ( .A(n6423), .ZN(n6442) );
  INV_X2 U7316 ( .A(n6442), .ZN(n6960) );
  NAND2_X1 U7317 ( .A1(n6960), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5587) );
  AND2_X2 U7318 ( .A1(n9996), .A2(n5585), .ZN(n6416) );
  NAND2_X1 U7319 ( .A1(n6589), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5586) );
  NOR2_X1 U7320 ( .A1(n6965), .A2(n9273), .ZN(n6380) );
  AOI21_X1 U7321 ( .B1(n9597), .B2(n9894), .A(n6380), .ZN(n5621) );
  NAND2_X1 U7322 ( .A1(n5592), .A2(n5589), .ZN(n5590) );
  XNOR2_X1 U7323 ( .A(n5592), .B(P1_IR_REG_25__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U7324 ( .A1(n5593), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5594) );
  OAI211_X1 U7325 ( .C1(n9344), .C2(n6721), .A(n6717), .B(n8128), .ZN(n6943)
         );
  INV_X1 U7326 ( .A(n5600), .ZN(n8176) );
  NAND3_X1 U7327 ( .A1(n8176), .A2(P1_B_REG_SCAN_IN), .A3(n8143), .ZN(n5601)
         );
  INV_X1 U7328 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10248) );
  INV_X1 U7329 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10267) );
  INV_X1 U7330 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10260) );
  INV_X1 U7331 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10297) );
  NAND4_X1 U7332 ( .A1(n10248), .A2(n10267), .A3(n10260), .A4(n10297), .ZN(
        n5602) );
  NOR3_X1 U7333 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        n5602), .ZN(n10227) );
  NOR4_X1 U7334 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n5609) );
  NOR4_X1 U7335 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n5608) );
  NOR4_X1 U7336 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5606) );
  NOR4_X1 U7337 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5605) );
  NOR4_X1 U7338 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5604) );
  NOR4_X1 U7339 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n5603) );
  AND4_X1 U7340 ( .A1(n5606), .A2(n5605), .A3(n5604), .A4(n5603), .ZN(n5607)
         );
  AND4_X1 U7341 ( .A1(n10227), .A2(n5609), .A3(n5608), .A4(n5607), .ZN(n5610)
         );
  OR2_X1 U7342 ( .A1(n9983), .A2(n5610), .ZN(n6933) );
  NAND2_X1 U7343 ( .A1(n6933), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5611) );
  OR2_X1 U7344 ( .A1(n9983), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5613) );
  INV_X1 U7345 ( .A(n5612), .ZN(n8200) );
  NAND2_X1 U7346 ( .A1(n8200), .A2(n8176), .ZN(n9984) );
  NAND2_X1 U7347 ( .A1(n5613), .A2(n9984), .ZN(n7632) );
  INV_X1 U7348 ( .A(n7632), .ZN(n6934) );
  OR2_X1 U7349 ( .A1(n9983), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U7350 ( .A1(n8200), .A2(n8143), .ZN(n5615) );
  MUX2_X1 U7351 ( .A(n5617), .B(n5621), .S(n10123), .Z(n5618) );
  NAND2_X1 U7352 ( .A1(n5618), .A2(n5176), .ZN(P1_U3553) );
  INV_X1 U7353 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n5622) );
  MUX2_X1 U7354 ( .A(n5622), .B(n5621), .S(n10115), .Z(n5623) );
  NAND2_X1 U7355 ( .A1(n5623), .A2(n5171), .ZN(P1_U3521) );
  INV_X1 U7356 ( .A(n5781), .ZN(n5626) );
  INV_X1 U7357 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5634) );
  INV_X1 U7358 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U7359 ( .A1(n6016), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5637) );
  NAND2_X1 U7360 ( .A1(n6062), .A2(n5637), .ZN(n8883) );
  NOR2_X1 U7361 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5639) );
  NOR2_X1 U7362 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5642) );
  NOR2_X1 U7363 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n5641) );
  NAND2_X1 U7364 ( .A1(n8883), .A2(n6143), .ZN(n5653) );
  INV_X1 U7365 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8882) );
  NAND2_X1 U7366 ( .A1(n8312), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U7367 ( .A1(n8311), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5649) );
  OAI211_X1 U7368 ( .C1(n8882), .C2(n4695), .A(n5650), .B(n5649), .ZN(n5651)
         );
  INV_X1 U7369 ( .A(n5651), .ZN(n5652) );
  NAND2_X1 U7370 ( .A1(n5683), .A2(n5655), .ZN(n5689) );
  NOR2_X1 U7371 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n5657) );
  OAI21_X1 U7372 ( .B1(n5658), .B2(n4520), .A(n5657), .ZN(n5662) );
  NAND2_X1 U7373 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n5659) );
  NOR2_X1 U7374 ( .A1(n4520), .A2(n5659), .ZN(n5660) );
  NAND2_X1 U7375 ( .A1(n5691), .A2(n5660), .ZN(n5661) );
  NAND2_X1 U7376 ( .A1(n7002), .A2(n8310), .ZN(n5671) );
  INV_X1 U7378 ( .A(n5735), .ZN(n5666) );
  INV_X1 U7379 ( .A(n5774), .ZN(n5668) );
  INV_X1 U7380 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5667) );
  INV_X1 U7381 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U7382 ( .A1(n5707), .A2(n5669), .ZN(n5804) );
  NAND2_X1 U7383 ( .A1(n5804), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5792) );
  XNOR2_X1 U7384 ( .A(n5792), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6305) );
  AOI22_X1 U7385 ( .A1(n8309), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6305), .B2(
        n5749), .ZN(n5670) );
  NAND2_X1 U7386 ( .A1(n5671), .A2(n5670), .ZN(n7572) );
  NOR2_X1 U7387 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5675) );
  OR2_X1 U7388 ( .A1(n5680), .A2(n5679), .ZN(n5681) );
  INV_X1 U7389 ( .A(n8324), .ZN(n5696) );
  INV_X1 U7390 ( .A(P2_B_REG_SCAN_IN), .ZN(n6168) );
  INV_X1 U7391 ( .A(n8203), .ZN(n5693) );
  INV_X1 U7392 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7011) );
  NAND2_X1 U7393 ( .A1(n5697), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5698) );
  NAND2_X1 U7394 ( .A1(n6057), .A2(n8509), .ZN(n5699) );
  NAND2_X1 U7395 ( .A1(n5699), .A2(n8479), .ZN(n5700) );
  XNOR2_X1 U7396 ( .A(n7572), .B(n5903), .ZN(n5789) );
  INV_X1 U7397 ( .A(n5789), .ZN(n5790) );
  NAND2_X1 U7398 ( .A1(n6161), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5706) );
  INV_X1 U7399 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10266) );
  OR2_X1 U7400 ( .A1(n4283), .A2(n10266), .ZN(n5705) );
  INV_X1 U7401 ( .A(n5701), .ZN(n5714) );
  NAND2_X1 U7402 ( .A1(n5714), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5702) );
  AND2_X1 U7403 ( .A1(n5797), .A2(n5702), .ZN(n7804) );
  OR2_X1 U7404 ( .A1(n5742), .A2(n7804), .ZN(n5704) );
  INV_X1 U7405 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10311) );
  OR2_X1 U7406 ( .A1(n5854), .A2(n10311), .ZN(n5703) );
  NAND2_X1 U7407 ( .A1(n5708), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5709) );
  AND2_X1 U7408 ( .A1(n5749), .A2(n6304), .ZN(n5710) );
  AOI21_X1 U7409 ( .B1(n8309), .B2(P1_DATAO_REG_6__SCAN_IN), .A(n5710), .ZN(
        n5712) );
  NAND2_X1 U7410 ( .A1(n6998), .A2(n8310), .ZN(n5711) );
  XNOR2_X1 U7411 ( .A(n5903), .B(n7702), .ZN(n5787) );
  INV_X1 U7412 ( .A(n5787), .ZN(n5788) );
  NAND2_X1 U7413 ( .A1(n8311), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5718) );
  INV_X1 U7414 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10197) );
  OR2_X1 U7415 ( .A1(n4282), .A2(n10197), .ZN(n5717) );
  NAND2_X1 U7416 ( .A1(n5781), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5713) );
  AND2_X1 U7417 ( .A1(n5714), .A2(n5713), .ZN(n7492) );
  OR2_X1 U7418 ( .A1(n5742), .A2(n7492), .ZN(n5716) );
  INV_X1 U7419 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7491) );
  OR2_X1 U7420 ( .A1(n5761), .A2(n7491), .ZN(n5715) );
  INV_X1 U7421 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5719) );
  OR2_X1 U7422 ( .A1(n5854), .A2(n5719), .ZN(n5723) );
  NAND2_X1 U7423 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5720) );
  AND2_X1 U7424 ( .A1(n5779), .A2(n5720), .ZN(n7356) );
  OR2_X1 U7425 ( .A1(n5742), .A2(n7356), .ZN(n5722) );
  INV_X1 U7426 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7464) );
  OR2_X1 U7427 ( .A1(n5773), .A2(n6996), .ZN(n5727) );
  NAND2_X1 U7428 ( .A1(n5735), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5725) );
  XNOR2_X1 U7429 ( .A(n5725), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7181) );
  NAND2_X1 U7430 ( .A1(n5749), .A2(n7181), .ZN(n5726) );
  OAI211_X1 U7431 ( .C1(n5757), .C2(n6997), .A(n5727), .B(n5726), .ZN(n7466)
         );
  INV_X1 U7432 ( .A(n7466), .ZN(n10167) );
  XNOR2_X1 U7433 ( .A(n5903), .B(n10167), .ZN(n5771) );
  INV_X1 U7434 ( .A(n5771), .ZN(n5772) );
  INV_X1 U7435 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5728) );
  OR2_X1 U7436 ( .A1(n5742), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5732) );
  INV_X1 U7437 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7482) );
  INV_X1 U7438 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5729) );
  OR2_X1 U7439 ( .A1(n5854), .A2(n5729), .ZN(n5730) );
  OR2_X1 U7440 ( .A1(n5773), .A2(n6991), .ZN(n5738) );
  MUX2_X1 U7441 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5734), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5736) );
  NAND2_X1 U7442 ( .A1(n5749), .A2(n6301), .ZN(n5737) );
  OAI211_X1 U7443 ( .C1(n5757), .C2(n6992), .A(n5738), .B(n5737), .ZN(n7484)
         );
  INV_X1 U7444 ( .A(n7484), .ZN(n7419) );
  INV_X1 U7445 ( .A(n5769), .ZN(n5770) );
  NAND2_X1 U7446 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5739) );
  NAND2_X1 U7447 ( .A1(n5749), .A2(n7143), .ZN(n5740) );
  NAND2_X1 U7448 ( .A1(n6161), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5747) );
  INV_X1 U7449 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10189) );
  OR2_X1 U7450 ( .A1(n6164), .A2(n10189), .ZN(n5746) );
  INV_X1 U7451 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n5741) );
  INV_X1 U7452 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5743) );
  OR2_X1 U7453 ( .A1(n5854), .A2(n5743), .ZN(n5744) );
  AND4_X2 U7454 ( .A1(n5747), .A2(n5746), .A3(n5745), .A4(n5744), .ZN(n6092)
         );
  XNOR2_X1 U7455 ( .A(n5752), .B(n6092), .ZN(n7274) );
  NAND2_X1 U7456 ( .A1(n6990), .A2(SI_0_), .ZN(n5748) );
  XNOR2_X1 U7457 ( .A(n5748), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9065) );
  INV_X1 U7458 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7451) );
  OR2_X1 U7459 ( .A1(n5742), .A2(n7451), .ZN(n5751) );
  INV_X1 U7460 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10187) );
  INV_X1 U7461 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6236) );
  OR2_X1 U7462 ( .A1(n5761), .A2(n6236), .ZN(n5750) );
  AOI21_X1 U7463 ( .B1(n6339), .B2(n8334), .A(n7299), .ZN(n7275) );
  INV_X1 U7464 ( .A(n5752), .ZN(n5753) );
  NAND2_X1 U7465 ( .A1(n5755), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5756) );
  OR2_X1 U7466 ( .A1(n5757), .A2(n7013), .ZN(n5759) );
  OR2_X1 U7467 ( .A1(n5773), .A2(n7014), .ZN(n5758) );
  XNOR2_X1 U7468 ( .A(n5760), .B(n10161), .ZN(n5767) );
  NAND2_X1 U7469 ( .A1(n5851), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5766) );
  INV_X1 U7470 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10191) );
  OR2_X1 U7471 ( .A1(n4283), .A2(n10191), .ZN(n5765) );
  INV_X1 U7472 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10147) );
  INV_X1 U7473 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5762) );
  OR2_X1 U7474 ( .A1(n5854), .A2(n5762), .ZN(n5763) );
  AND4_X2 U7475 ( .A1(n5766), .A2(n5765), .A3(n5764), .A4(n5763), .ZN(n7385)
         );
  XNOR2_X1 U7476 ( .A(n5767), .B(n7385), .ZN(n7336) );
  INV_X1 U7477 ( .A(n5767), .ZN(n5768) );
  XNOR2_X1 U7478 ( .A(n5769), .B(n7353), .ZN(n7220) );
  NAND2_X1 U7479 ( .A1(n7221), .A2(n7220), .ZN(n7219) );
  XNOR2_X1 U7480 ( .A(n5771), .B(n8753), .ZN(n7350) );
  NAND2_X1 U7481 ( .A1(n8309), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5778) );
  OR2_X1 U7482 ( .A1(n5773), .A2(n6993), .ZN(n5777) );
  NAND2_X1 U7483 ( .A1(n5774), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5775) );
  XNOR2_X1 U7484 ( .A(n5775), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U7485 ( .A1(n5749), .A2(n6302), .ZN(n5776) );
  XNOR2_X1 U7486 ( .A(n5903), .B(n10171), .ZN(n5786) );
  INV_X1 U7487 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10195) );
  OR2_X1 U7488 ( .A1(n4282), .A2(n10195), .ZN(n5785) );
  NAND2_X1 U7489 ( .A1(n6161), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5784) );
  NAND2_X1 U7490 ( .A1(n8311), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U7491 ( .A1(n5779), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5780) );
  AND2_X1 U7492 ( .A1(n5781), .A2(n5780), .ZN(n7445) );
  OR2_X1 U7493 ( .A1(n5742), .A2(n7445), .ZN(n5782) );
  XNOR2_X1 U7494 ( .A(n5786), .B(n8752), .ZN(n7471) );
  XNOR2_X1 U7495 ( .A(n5787), .B(n7474), .ZN(n7699) );
  XNOR2_X1 U7496 ( .A(n5789), .B(n8750), .ZN(n7801) );
  NAND2_X1 U7497 ( .A1(n7802), .A2(n7801), .ZN(n7800) );
  OAI21_X1 U7498 ( .B1(n5790), .B2(n8750), .A(n7800), .ZN(n7920) );
  NAND2_X1 U7499 ( .A1(n7004), .A2(n8310), .ZN(n5796) );
  INV_X1 U7500 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5791) );
  NAND2_X1 U7501 ( .A1(n5792), .A2(n5791), .ZN(n5793) );
  NAND2_X1 U7502 ( .A1(n5793), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5794) );
  AOI22_X1 U7503 ( .A1(n8309), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7016), .B2(
        n5749), .ZN(n5795) );
  XNOR2_X1 U7504 ( .A(n7927), .B(n6338), .ZN(n5803) );
  NAND2_X1 U7505 ( .A1(n8311), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5802) );
  INV_X1 U7506 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7582) );
  OR2_X1 U7507 ( .A1(n4283), .A2(n7582), .ZN(n5801) );
  NAND2_X1 U7508 ( .A1(n5797), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5798) );
  AND2_X1 U7509 ( .A1(n5808), .A2(n5798), .ZN(n7924) );
  OR2_X1 U7510 ( .A1(n5742), .A2(n7924), .ZN(n5800) );
  INV_X1 U7511 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7586) );
  OR2_X1 U7512 ( .A1(n5761), .A2(n7586), .ZN(n5799) );
  XNOR2_X1 U7513 ( .A(n5803), .B(n8749), .ZN(n7919) );
  NAND2_X1 U7514 ( .A1(n7018), .A2(n8310), .ZN(n5807) );
  OAI21_X1 U7515 ( .B1(n5804), .B2(n4398), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5805) );
  XNOR2_X1 U7516 ( .A(n5805), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7606) );
  AOI22_X1 U7517 ( .A1(n8309), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7606), .B2(
        n5749), .ZN(n5806) );
  INV_X2 U7518 ( .A(n4706), .ZN(n6338) );
  XNOR2_X1 U7519 ( .A(n7627), .B(n6338), .ZN(n5815) );
  NAND2_X1 U7520 ( .A1(n8311), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5814) );
  INV_X1 U7521 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7629) );
  OR2_X1 U7522 ( .A1(n4282), .A2(n7629), .ZN(n5813) );
  NAND2_X1 U7523 ( .A1(n5808), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5809) );
  AND2_X1 U7524 ( .A1(n5829), .A2(n5809), .ZN(n8054) );
  OR2_X1 U7525 ( .A1(n5742), .A2(n8054), .ZN(n5812) );
  INV_X1 U7526 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5810) );
  OR2_X1 U7527 ( .A1(n5761), .A2(n5810), .ZN(n5811) );
  XNOR2_X1 U7528 ( .A(n5815), .B(n8748), .ZN(n8052) );
  OR2_X1 U7529 ( .A1(n5815), .A2(n7923), .ZN(n5816) );
  NAND2_X1 U7530 ( .A1(n5817), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5846) );
  XNOR2_X1 U7531 ( .A(n5846), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8086) );
  AOI22_X1 U7532 ( .A1(n8309), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8086), .B2(
        n5749), .ZN(n5818) );
  NAND2_X1 U7533 ( .A1(n8312), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U7534 ( .A1(n5831), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U7535 ( .A1(n5852), .A2(n5820), .ZN(n7730) );
  INV_X1 U7536 ( .A(n7730), .ZN(n8695) );
  OR2_X1 U7537 ( .A1(n8695), .A2(n5742), .ZN(n5823) );
  OR2_X1 U7538 ( .A1(n4695), .A2(n4919), .ZN(n5822) );
  INV_X1 U7539 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7724) );
  OR2_X1 U7540 ( .A1(n5854), .A2(n7724), .ZN(n5821) );
  XNOR2_X1 U7541 ( .A(n8292), .B(n6338), .ZN(n8691) );
  NAND2_X1 U7542 ( .A1(n7025), .A2(n8310), .ZN(n5828) );
  NAND2_X1 U7543 ( .A1(n5825), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5826) );
  XNOR2_X1 U7544 ( .A(n5826), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6310) );
  AOI22_X1 U7545 ( .A1(n8309), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6310), .B2(
        n5749), .ZN(n5827) );
  XNOR2_X1 U7546 ( .A(n8197), .B(n5903), .ZN(n8688) );
  INV_X1 U7547 ( .A(n8688), .ZN(n5837) );
  NAND2_X1 U7548 ( .A1(n8312), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5835) );
  NAND2_X1 U7549 ( .A1(n6161), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U7550 ( .A1(n8311), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U7551 ( .A1(n5829), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5830) );
  AND2_X1 U7552 ( .A1(n5831), .A2(n5830), .ZN(n7742) );
  OR2_X1 U7553 ( .A1(n5742), .A2(n7742), .ZN(n5832) );
  NAND4_X1 U7554 ( .A1(n5835), .A2(n5834), .A3(n5833), .A4(n5832), .ZN(n8747)
         );
  NOR2_X1 U7555 ( .A1(n6108), .A2(n6338), .ZN(n5840) );
  AOI211_X1 U7556 ( .C1(n8746), .C2(n6338), .A(n5840), .B(n8292), .ZN(n5843)
         );
  NOR2_X1 U7557 ( .A1(n6338), .A2(n8192), .ZN(n5841) );
  AOI211_X1 U7558 ( .C1(n8383), .C2(n6338), .A(n5841), .B(n7721), .ZN(n5842)
         );
  NAND2_X1 U7559 ( .A1(n7111), .A2(n8310), .ZN(n5850) );
  NAND2_X1 U7560 ( .A1(n5846), .A2(n5845), .ZN(n5847) );
  NAND2_X1 U7561 ( .A1(n5847), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5848) );
  XNOR2_X1 U7562 ( .A(n5848), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7113) );
  AOI22_X1 U7563 ( .A1(n8309), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7113), .B2(
        n5749), .ZN(n5849) );
  XOR2_X1 U7564 ( .A(n6338), .B(n8185), .Z(n8179) );
  NAND2_X1 U7565 ( .A1(n5852), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5853) );
  NAND2_X1 U7566 ( .A1(n5861), .A2(n5853), .ZN(n8184) );
  NAND2_X1 U7567 ( .A1(n6143), .A2(n8184), .ZN(n5858) );
  INV_X1 U7568 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7865) );
  OR2_X1 U7569 ( .A1(n5854), .A2(n7865), .ZN(n5857) );
  INV_X1 U7570 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7868) );
  OR2_X1 U7571 ( .A1(n4283), .A2(n7868), .ZN(n5856) );
  INV_X1 U7572 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10223) );
  OR2_X1 U7573 ( .A1(n4695), .A2(n10223), .ZN(n5855) );
  NAND2_X1 U7574 ( .A1(n7227), .A2(n8310), .ZN(n6121) );
  NAND2_X1 U7575 ( .A1(n5859), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5860) );
  XNOR2_X1 U7576 ( .A(n5860), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6315) );
  AOI22_X1 U7577 ( .A1(n8309), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6315), .B2(
        n5749), .ZN(n6119) );
  NAND2_X1 U7578 ( .A1(n6121), .A2(n6119), .ZN(n8016) );
  XNOR2_X1 U7579 ( .A(n8016), .B(n6338), .ZN(n5867) );
  NAND2_X1 U7580 ( .A1(n5861), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U7581 ( .A1(n5875), .A2(n5862), .ZN(n8671) );
  NAND2_X1 U7582 ( .A1(n8671), .A2(n6143), .ZN(n5866) );
  NAND2_X1 U7583 ( .A1(n8311), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5865) );
  NAND2_X1 U7584 ( .A1(n8312), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U7585 ( .A1(n6161), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U7586 ( .A1(n5867), .A2(n8594), .ZN(n8664) );
  INV_X1 U7587 ( .A(n5867), .ZN(n5868) );
  NAND2_X1 U7588 ( .A1(n5868), .A2(n6118), .ZN(n8665) );
  NAND2_X1 U7589 ( .A1(n7319), .A2(n8310), .ZN(n5874) );
  NAND2_X1 U7590 ( .A1(n5871), .A2(n5870), .ZN(n5872) );
  NAND2_X1 U7591 ( .A1(n5872), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5899) );
  XNOR2_X1 U7592 ( .A(n5899), .B(P2_IR_REG_14__SCAN_IN), .ZN(n6319) );
  AOI22_X1 U7593 ( .A1(n8309), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6319), .B2(
        n5749), .ZN(n5873) );
  XNOR2_X1 U7594 ( .A(n8597), .B(n6338), .ZN(n5882) );
  NAND2_X1 U7595 ( .A1(n5875), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5876) );
  NAND2_X1 U7596 ( .A1(n5889), .A2(n5876), .ZN(n8596) );
  NAND2_X1 U7597 ( .A1(n8596), .A2(n6143), .ZN(n5881) );
  NAND2_X1 U7598 ( .A1(n8311), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U7599 ( .A1(n8312), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5877) );
  AND2_X1 U7600 ( .A1(n5878), .A2(n5877), .ZN(n5880) );
  NAND2_X1 U7601 ( .A1(n6161), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5879) );
  XNOR2_X1 U7602 ( .A(n5882), .B(n8669), .ZN(n8591) );
  NAND2_X1 U7603 ( .A1(n5882), .A2(n8669), .ZN(n5883) );
  NAND2_X1 U7604 ( .A1(n7345), .A2(n8310), .ZN(n5888) );
  NAND2_X1 U7605 ( .A1(n5899), .A2(n5884), .ZN(n5885) );
  NAND2_X1 U7606 ( .A1(n5885), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5886) );
  XNOR2_X1 U7607 ( .A(n5886), .B(P2_IR_REG_15__SCAN_IN), .ZN(n6320) );
  AOI22_X1 U7608 ( .A1(n8309), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6320), .B2(
        n5749), .ZN(n5887) );
  XNOR2_X1 U7609 ( .A(n8716), .B(n6338), .ZN(n5894) );
  NAND2_X1 U7610 ( .A1(n5889), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U7611 ( .A1(n5904), .A2(n5890), .ZN(n8728) );
  NAND2_X1 U7612 ( .A1(n8728), .A2(n6143), .ZN(n5893) );
  AOI22_X1 U7613 ( .A1(n8311), .A2(P2_REG0_REG_15__SCAN_IN), .B1(n8312), .B2(
        P2_REG1_REG_15__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7614 ( .A1(n6161), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5891) );
  XNOR2_X1 U7615 ( .A(n5894), .B(n8023), .ZN(n8718) );
  INV_X1 U7616 ( .A(n5894), .ZN(n5895) );
  NAND2_X1 U7617 ( .A1(n7393), .A2(n8310), .ZN(n5902) );
  INV_X1 U7618 ( .A(n5896), .ZN(n5897) );
  NAND2_X1 U7619 ( .A1(n5897), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U7620 ( .A1(n5899), .A2(n5898), .ZN(n5911) );
  XNOR2_X1 U7621 ( .A(n5911), .B(n5900), .ZN(n6322) );
  AOI22_X1 U7622 ( .A1(n8309), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5749), .B2(
        n6322), .ZN(n5901) );
  XOR2_X1 U7623 ( .A(n5903), .B(n8634), .Z(n8628) );
  NAND2_X1 U7624 ( .A1(n5904), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5905) );
  NAND2_X1 U7625 ( .A1(n5915), .A2(n5905), .ZN(n8633) );
  NAND2_X1 U7626 ( .A1(n8633), .A2(n6143), .ZN(n5910) );
  INV_X1 U7627 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8167) );
  NAND2_X1 U7628 ( .A1(n8312), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U7629 ( .A1(n8311), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5906) );
  OAI211_X1 U7630 ( .C1(n4695), .C2(n8167), .A(n5907), .B(n5906), .ZN(n5908)
         );
  INV_X1 U7631 ( .A(n5908), .ZN(n5909) );
  NAND2_X1 U7632 ( .A1(n7396), .A2(n8310), .ZN(n5914) );
  OAI21_X1 U7633 ( .B1(n5911), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5912) );
  XNOR2_X1 U7634 ( .A(n5912), .B(P2_IR_REG_17__SCAN_IN), .ZN(n6323) );
  AOI22_X1 U7635 ( .A1(n8309), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6323), .B2(
        n5749), .ZN(n5913) );
  XNOR2_X1 U7636 ( .A(n8644), .B(n6338), .ZN(n5952) );
  NAND2_X1 U7637 ( .A1(n5915), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5916) );
  NAND2_X1 U7638 ( .A1(n5958), .A2(n5916), .ZN(n8643) );
  NAND2_X1 U7639 ( .A1(n8643), .A2(n6143), .ZN(n5921) );
  INV_X1 U7640 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8213) );
  NAND2_X1 U7641 ( .A1(n8311), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5918) );
  NAND2_X1 U7642 ( .A1(n8312), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5917) );
  OAI211_X1 U7643 ( .C1(n8213), .C2(n4695), .A(n5918), .B(n5917), .ZN(n5919)
         );
  INV_X1 U7644 ( .A(n5919), .ZN(n5920) );
  NAND2_X1 U7645 ( .A1(n5952), .A2(n8708), .ZN(n8638) );
  NAND2_X1 U7646 ( .A1(n8039), .A2(n8310), .ZN(n5923) );
  NAND2_X1 U7647 ( .A1(n8309), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5922) );
  NAND2_X1 U7648 ( .A1(n5923), .A2(n5922), .ZN(n6132) );
  XNOR2_X1 U7649 ( .A(n6132), .B(n6338), .ZN(n5971) );
  NAND2_X1 U7650 ( .A1(n5942), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7651 ( .A1(n5974), .A2(n5924), .ZN(n8257) );
  NAND2_X1 U7652 ( .A1(n8257), .A2(n6143), .ZN(n5929) );
  INV_X1 U7653 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8240) );
  NAND2_X1 U7654 ( .A1(n8312), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U7655 ( .A1(n8311), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5925) );
  OAI211_X1 U7656 ( .C1(n8240), .C2(n4695), .A(n5926), .B(n5925), .ZN(n5927)
         );
  INV_X1 U7657 ( .A(n5927), .ZN(n5928) );
  XNOR2_X1 U7658 ( .A(n5971), .B(n8934), .ZN(n8250) );
  NAND2_X1 U7659 ( .A1(n7859), .A2(n8310), .ZN(n5931) );
  NAND2_X1 U7660 ( .A1(n8309), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5930) );
  XNOR2_X1 U7661 ( .A(n9031), .B(n4706), .ZN(n8249) );
  NAND2_X1 U7662 ( .A1(n7676), .A2(n8310), .ZN(n5933) );
  AOI22_X1 U7663 ( .A1(n8309), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8509), .B2(
        n5749), .ZN(n5932) );
  XNOR2_X1 U7664 ( .A(n8613), .B(n4706), .ZN(n8246) );
  NAND2_X1 U7665 ( .A1(n5960), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5934) );
  NAND2_X1 U7666 ( .A1(n5940), .A2(n5934), .ZN(n8953) );
  NAND2_X1 U7667 ( .A1(n8953), .A2(n6143), .ZN(n5939) );
  INV_X1 U7668 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8952) );
  NAND2_X1 U7669 ( .A1(n8311), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U7670 ( .A1(n8312), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5935) );
  OAI211_X1 U7671 ( .C1(n8952), .C2(n4695), .A(n5936), .B(n5935), .ZN(n5937)
         );
  INV_X1 U7672 ( .A(n5937), .ZN(n5938) );
  NAND2_X1 U7673 ( .A1(n5940), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U7674 ( .A1(n5942), .A2(n5941), .ZN(n8937) );
  NAND2_X1 U7675 ( .A1(n8937), .A2(n6143), .ZN(n5947) );
  INV_X1 U7676 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8936) );
  NAND2_X1 U7677 ( .A1(n8311), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U7678 ( .A1(n8312), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5943) );
  OAI211_X1 U7679 ( .C1(n8936), .C2(n4695), .A(n5944), .B(n5943), .ZN(n5945)
         );
  INV_X1 U7680 ( .A(n5945), .ZN(n5946) );
  OAI21_X1 U7681 ( .B1(n8246), .B2(n8247), .A(n8948), .ZN(n5950) );
  INV_X1 U7682 ( .A(n8246), .ZN(n5949) );
  NOR2_X1 U7683 ( .A1(n8948), .A2(n8247), .ZN(n5948) );
  AOI22_X1 U7684 ( .A1(n8249), .A2(n5950), .B1(n5949), .B2(n5948), .ZN(n5951)
         );
  NAND2_X1 U7685 ( .A1(n8250), .A2(n5951), .ZN(n8251) );
  INV_X1 U7686 ( .A(n8251), .ZN(n5967) );
  INV_X1 U7687 ( .A(n5952), .ZN(n5953) );
  NAND2_X1 U7688 ( .A1(n5953), .A2(n8158), .ZN(n8700) );
  NAND2_X1 U7689 ( .A1(n7495), .A2(n8310), .ZN(n5957) );
  NAND2_X1 U7690 ( .A1(n5954), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5955) );
  XNOR2_X1 U7691 ( .A(n5955), .B(P2_IR_REG_18__SCAN_IN), .ZN(n6325) );
  AOI22_X1 U7692 ( .A1(n8309), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6325), .B2(
        n5749), .ZN(n5956) );
  XNOR2_X1 U7693 ( .A(n8712), .B(n6338), .ZN(n5970) );
  NAND2_X1 U7694 ( .A1(n5958), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U7695 ( .A1(n5960), .A2(n5959), .ZN(n8710) );
  NAND2_X1 U7696 ( .A1(n8710), .A2(n6143), .ZN(n5965) );
  INV_X1 U7697 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n10275) );
  NAND2_X1 U7698 ( .A1(n8311), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7699 ( .A1(n6161), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5961) );
  OAI211_X1 U7700 ( .C1(n4282), .C2(n10275), .A(n5962), .B(n5961), .ZN(n5963)
         );
  INV_X1 U7701 ( .A(n5963), .ZN(n5964) );
  XNOR2_X1 U7702 ( .A(n5970), .B(n8947), .ZN(n8703) );
  INV_X1 U7703 ( .A(n8703), .ZN(n5966) );
  AND2_X1 U7704 ( .A1(n8700), .A2(n5966), .ZN(n8244) );
  AND2_X1 U7705 ( .A1(n5967), .A2(n8244), .ZN(n5968) );
  NAND2_X1 U7706 ( .A1(n8701), .A2(n5968), .ZN(n5983) );
  INV_X1 U7707 ( .A(n8249), .ZN(n5969) );
  AOI22_X1 U7708 ( .A1(n5969), .A2(n8948), .B1(n8247), .B2(n8246), .ZN(n8252)
         );
  NAND2_X1 U7709 ( .A1(n5970), .A2(n8947), .ZN(n8245) );
  AOI21_X1 U7710 ( .B1(n8252), .B2(n8245), .A(n8251), .ZN(n5981) );
  AND2_X1 U7711 ( .A1(n5971), .A2(n8919), .ZN(n8677) );
  NAND2_X1 U7712 ( .A1(n8034), .A2(n8310), .ZN(n5973) );
  NAND2_X1 U7713 ( .A1(n8309), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5972) );
  XNOR2_X1 U7714 ( .A(n8675), .B(n6338), .ZN(n5984) );
  NAND2_X1 U7715 ( .A1(n5974), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U7716 ( .A1(n5989), .A2(n5975), .ZN(n8923) );
  NAND2_X1 U7717 ( .A1(n8923), .A2(n6143), .ZN(n5980) );
  INV_X1 U7718 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n10279) );
  NAND2_X1 U7719 ( .A1(n8311), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U7720 ( .A1(n6161), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5976) );
  OAI211_X1 U7721 ( .C1(n4283), .C2(n10279), .A(n5977), .B(n5976), .ZN(n5978)
         );
  INV_X1 U7722 ( .A(n5978), .ZN(n5979) );
  XNOR2_X1 U7723 ( .A(n5984), .B(n8255), .ZN(n8676) );
  NOR3_X1 U7724 ( .A1(n5981), .A2(n8677), .A3(n8676), .ZN(n5982) );
  INV_X1 U7725 ( .A(n5984), .ZN(n5985) );
  NAND2_X1 U7726 ( .A1(n5985), .A2(n8910), .ZN(n5986) );
  NAND2_X1 U7727 ( .A1(n8127), .A2(n8310), .ZN(n5988) );
  NAND2_X1 U7728 ( .A1(n8309), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5987) );
  XNOR2_X1 U7729 ( .A(n9021), .B(n6338), .ZN(n8601) );
  NAND2_X1 U7730 ( .A1(n5989), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7731 ( .A1(n5998), .A2(n5990), .ZN(n8914) );
  NAND2_X1 U7732 ( .A1(n8914), .A2(n6143), .ZN(n5995) );
  INV_X1 U7733 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8913) );
  NAND2_X1 U7734 ( .A1(n8311), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U7735 ( .A1(n8312), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5991) );
  OAI211_X1 U7736 ( .C1(n8913), .C2(n4695), .A(n5992), .B(n5991), .ZN(n5993)
         );
  INV_X1 U7737 ( .A(n5993), .ZN(n5994) );
  NAND2_X1 U7738 ( .A1(n8601), .A2(n8920), .ZN(n6009) );
  NAND2_X1 U7739 ( .A1(n8139), .A2(n8310), .ZN(n5997) );
  NAND2_X1 U7740 ( .A1(n8309), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5996) );
  XNOR2_X1 U7741 ( .A(n8457), .B(n6338), .ZN(n6006) );
  INV_X1 U7742 ( .A(n6006), .ZN(n6007) );
  NAND2_X1 U7743 ( .A1(n5998), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U7744 ( .A1(n6014), .A2(n5999), .ZN(n8901) );
  NAND2_X1 U7745 ( .A1(n8901), .A2(n6143), .ZN(n6005) );
  INV_X1 U7746 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7747 ( .A1(n8311), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6001) );
  NAND2_X1 U7748 ( .A1(n8312), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6000) );
  OAI211_X1 U7749 ( .C1(n6002), .C2(n4695), .A(n6001), .B(n6000), .ZN(n6003)
         );
  INV_X1 U7750 ( .A(n6003), .ZN(n6004) );
  AOI21_X1 U7751 ( .B1(n6007), .B2(n8911), .A(n6026), .ZN(n8648) );
  OAI21_X1 U7752 ( .B1(n8920), .B2(n8601), .A(n8648), .ZN(n6008) );
  NAND2_X1 U7753 ( .A1(n8198), .A2(n8310), .ZN(n6011) );
  NAND2_X1 U7754 ( .A1(n8309), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6010) );
  XNOR2_X1 U7755 ( .A(n8884), .B(n6338), .ZN(n6334) );
  INV_X1 U7756 ( .A(n6334), .ZN(n6023) );
  NAND2_X1 U7757 ( .A1(n8171), .A2(n8310), .ZN(n6013) );
  NAND2_X1 U7758 ( .A1(n8309), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6012) );
  XNOR2_X1 U7759 ( .A(n9011), .B(n4706), .ZN(n6024) );
  INV_X1 U7760 ( .A(n6024), .ZN(n6332) );
  NAND2_X1 U7761 ( .A1(n6014), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7762 ( .A1(n6016), .A2(n6015), .ZN(n8894) );
  NAND2_X1 U7763 ( .A1(n8894), .A2(n6143), .ZN(n6022) );
  INV_X1 U7764 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U7765 ( .A1(n8311), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7766 ( .A1(n8312), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6017) );
  OAI211_X1 U7767 ( .C1(n6019), .C2(n4695), .A(n6018), .B(n6017), .ZN(n6020)
         );
  INV_X1 U7768 ( .A(n6020), .ZN(n6021) );
  NAND2_X1 U7769 ( .A1(n6332), .A2(n8899), .ZN(n6333) );
  NAND2_X1 U7770 ( .A1(n8620), .A2(n5180), .ZN(n6031) );
  NAND2_X1 U7771 ( .A1(n6024), .A2(n8737), .ZN(n6025) );
  INV_X1 U7772 ( .A(n6025), .ZN(n6029) );
  OAI21_X1 U7773 ( .B1(n6026), .B2(n8899), .A(n6332), .ZN(n6027) );
  OAI211_X1 U7774 ( .C1(n8618), .C2(n8737), .A(n6334), .B(n6027), .ZN(n6028)
         );
  OAI21_X1 U7775 ( .B1(n6029), .B2(n6334), .A(n6028), .ZN(n6030) );
  NAND2_X1 U7776 ( .A1(n6032), .A2(n8570), .ZN(n6337) );
  OAI21_X1 U7777 ( .B1(n8570), .B2(n6032), .A(n6337), .ZN(n6060) );
  INV_X1 U7778 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10237) );
  NAND2_X1 U7779 ( .A1(n7005), .A2(n10237), .ZN(n6033) );
  INV_X1 U7780 ( .A(n6047), .ZN(n8173) );
  NAND2_X1 U7781 ( .A1(n8173), .A2(n8203), .ZN(n7008) );
  NOR4_X1 U7782 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n10236) );
  NOR2_X1 U7783 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .ZN(
        n6036) );
  NOR4_X1 U7784 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6035) );
  NOR4_X1 U7785 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n6034) );
  NAND4_X1 U7786 ( .A1(n10236), .A2(n6036), .A3(n6035), .A4(n6034), .ZN(n6042)
         );
  NOR4_X1 U7787 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6040) );
  NOR4_X1 U7788 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6039) );
  NOR4_X1 U7789 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6038) );
  NOR4_X1 U7790 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6037) );
  NAND4_X1 U7791 ( .A1(n6040), .A2(n6039), .A3(n6038), .A4(n6037), .ZN(n6041)
         );
  OAI21_X1 U7792 ( .B1(n6042), .B2(n6041), .A(n7005), .ZN(n6074) );
  NAND2_X1 U7793 ( .A1(n7300), .A2(n6074), .ZN(n6045) );
  NOR2_X1 U7794 ( .A1(n8203), .A2(n5695), .ZN(n6046) );
  INV_X1 U7795 ( .A(n6048), .ZN(n6049) );
  NAND2_X1 U7796 ( .A1(n6049), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7797 ( .A1(n6080), .A2(n7007), .ZN(n6189) );
  INV_X1 U7798 ( .A(n6052), .ZN(n6053) );
  NAND2_X1 U7799 ( .A1(n6053), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U7800 ( .A1(n8509), .A2(n8513), .ZN(n6158) );
  OR2_X1 U7801 ( .A1(n6189), .A2(n6191), .ZN(n6059) );
  INV_X1 U7802 ( .A(n7300), .ZN(n6055) );
  NAND2_X1 U7803 ( .A1(n6055), .A2(n6044), .ZN(n6360) );
  INV_X1 U7804 ( .A(n6360), .ZN(n6056) );
  NAND2_X1 U7805 ( .A1(n6056), .A2(n6359), .ZN(n6194) );
  NAND3_X1 U7806 ( .A1(n8475), .A2(n6191), .A3(n10178), .ZN(n6073) );
  OR2_X1 U7807 ( .A1(n6194), .A2(n6073), .ZN(n6058) );
  NAND2_X1 U7808 ( .A1(n6060), .A2(n8679), .ZN(n6090) );
  OR2_X1 U7809 ( .A1(n6194), .A2(n10178), .ZN(n6061) );
  NAND2_X1 U7810 ( .A1(n7304), .A2(n8337), .ZN(n10172) );
  NAND2_X1 U7811 ( .A1(n6062), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7812 ( .A1(n6141), .A2(n6063), .ZN(n8872) );
  NAND2_X1 U7813 ( .A1(n8872), .A2(n6143), .ZN(n6068) );
  INV_X1 U7814 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n10276) );
  NAND2_X1 U7815 ( .A1(n6161), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7816 ( .A1(n8312), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6064) );
  OAI211_X1 U7817 ( .C1(n5854), .C2(n10276), .A(n6065), .B(n6064), .ZN(n6066)
         );
  INV_X1 U7818 ( .A(n6066), .ZN(n6067) );
  INV_X1 U7819 ( .A(n8881), .ZN(n8736) );
  NAND2_X1 U7820 ( .A1(n6070), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6071) );
  XNOR2_X1 U7821 ( .A(n6071), .B(P2_IR_REG_28__SCAN_IN), .ZN(n8510) );
  NAND2_X1 U7822 ( .A1(n6072), .A2(n5754), .ZN(n6167) );
  INV_X1 U7823 ( .A(n6167), .ZN(n6160) );
  NAND2_X1 U7824 ( .A1(n8479), .A2(n7677), .ZN(n6184) );
  OR3_X1 U7825 ( .A1(n6189), .A2(n6192), .A3(n6167), .ZN(n8707) );
  INV_X1 U7826 ( .A(n6074), .ZN(n6075) );
  NOR2_X1 U7827 ( .A1(n6360), .A2(n6075), .ZN(n6078) );
  NAND2_X1 U7828 ( .A1(n8499), .A2(n6184), .ZN(n6358) );
  AND3_X1 U7829 ( .A1(n6358), .A2(n6230), .A3(n6229), .ZN(n6077) );
  OR2_X1 U7830 ( .A1(n6080), .A2(n6191), .ZN(n6076) );
  OAI211_X1 U7831 ( .C1(n6190), .C2(n6078), .A(n6077), .B(n6076), .ZN(n6079)
         );
  NAND2_X1 U7832 ( .A1(n6079), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6084) );
  INV_X1 U7833 ( .A(n6080), .ZN(n6082) );
  NOR2_X1 U7834 ( .A1(n6192), .A2(n6081), .ZN(n8511) );
  NAND2_X1 U7835 ( .A1(n6082), .A2(n8511), .ZN(n6083) );
  AOI22_X1 U7836 ( .A1(n8883), .A2(n8727), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n6085) );
  OAI21_X1 U7837 ( .B1(n8899), .B2(n8707), .A(n6085), .ZN(n6086) );
  AOI21_X1 U7838 ( .B1(n8736), .B2(n8704), .A(n6086), .ZN(n6087) );
  INV_X1 U7839 ( .A(n6088), .ZN(n6089) );
  NAND2_X1 U7840 ( .A1(n6090), .A2(n6089), .ZN(P2_U3180) );
  NAND2_X1 U7841 ( .A1(n6093), .A2(n6092), .ZN(n10134) );
  NAND2_X1 U7842 ( .A1(n7305), .A2(n10134), .ZN(n6095) );
  NAND2_X1 U7843 ( .A1(n6095), .A2(n10126), .ZN(n10133) );
  NAND2_X1 U7844 ( .A1(n10161), .A2(n7385), .ZN(n6096) );
  INV_X1 U7845 ( .A(n7353), .ZN(n10130) );
  NAND2_X1 U7846 ( .A1(n10130), .A2(n7484), .ZN(n6097) );
  AND2_X1 U7847 ( .A1(n8753), .A2(n7466), .ZN(n7437) );
  NAND2_X1 U7848 ( .A1(n7419), .A2(n7353), .ZN(n7435) );
  NAND2_X1 U7849 ( .A1(n10167), .A2(n7440), .ZN(n7438) );
  INV_X1 U7850 ( .A(n8752), .ZN(n7352) );
  NAND2_X1 U7851 ( .A1(n10171), .A2(n7352), .ZN(n7433) );
  OAI211_X1 U7852 ( .C1(n7435), .C2(n7437), .A(n7438), .B(n7433), .ZN(n6098)
         );
  INV_X1 U7853 ( .A(n6098), .ZN(n6099) );
  INV_X1 U7854 ( .A(n10171), .ZN(n7446) );
  NAND2_X1 U7855 ( .A1(n7446), .A2(n8752), .ZN(n7432) );
  AND2_X1 U7856 ( .A1(n7702), .A2(n8751), .ZN(n6101) );
  AND2_X1 U7857 ( .A1(n7572), .A2(n8750), .ZN(n6100) );
  OR2_X1 U7858 ( .A1(n7927), .A2(n7810), .ZN(n8384) );
  NAND2_X1 U7859 ( .A1(n7927), .A2(n7810), .ZN(n8382) );
  INV_X1 U7860 ( .A(n7572), .ZN(n7803) );
  OAI21_X1 U7861 ( .B1(n7702), .B2(n8751), .A(n8750), .ZN(n6104) );
  NAND2_X1 U7862 ( .A1(n7696), .A2(n7474), .ZN(n6102) );
  NOR2_X1 U7863 ( .A1(n7702), .A2(n6102), .ZN(n6103) );
  AOI21_X1 U7864 ( .B1(n7803), .B2(n6104), .A(n6103), .ZN(n6105) );
  NAND2_X1 U7865 ( .A1(n7927), .A2(n8749), .ZN(n6107) );
  NAND2_X1 U7866 ( .A1(n7627), .A2(n8748), .ZN(n7706) );
  NAND2_X1 U7867 ( .A1(n6108), .A2(n7706), .ZN(n6112) );
  OR2_X1 U7868 ( .A1(n7627), .A2(n8748), .ZN(n7705) );
  NAND2_X1 U7869 ( .A1(n8197), .A2(n5836), .ZN(n7719) );
  NAND2_X1 U7870 ( .A1(n6113), .A2(n8746), .ZN(n6114) );
  AND2_X1 U7871 ( .A1(n8185), .A2(n8745), .ZN(n6117) );
  INV_X1 U7872 ( .A(n8594), .ZN(n6118) );
  AND2_X1 U7873 ( .A1(n6119), .A2(n6118), .ZN(n6120) );
  NAND2_X1 U7874 ( .A1(n6121), .A2(n6120), .ZN(n8406) );
  OR2_X1 U7875 ( .A1(n8016), .A2(n6118), .ZN(n6122) );
  XNOR2_X1 U7876 ( .A(n8597), .B(n8744), .ZN(n8407) );
  NAND2_X1 U7877 ( .A1(n8597), .A2(n8744), .ZN(n6124) );
  NAND2_X1 U7878 ( .A1(n8716), .A2(n8743), .ZN(n6125) );
  NAND2_X1 U7879 ( .A1(n8634), .A2(n8725), .ZN(n8417) );
  INV_X1 U7880 ( .A(n8298), .ZN(n6126) );
  NAND2_X1 U7881 ( .A1(n8634), .A2(n8741), .ZN(n6127) );
  NAND2_X1 U7882 ( .A1(n8644), .A2(n8708), .ZN(n8421) );
  NAND2_X1 U7883 ( .A1(n4324), .A2(n8421), .ZN(n8296) );
  NAND2_X1 U7884 ( .A1(n8644), .A2(n8158), .ZN(n6128) );
  OR2_X1 U7885 ( .A1(n8712), .A2(n8740), .ZN(n6129) );
  NAND2_X1 U7886 ( .A1(n6130), .A2(n8247), .ZN(n8425) );
  NAND2_X1 U7887 ( .A1(n4343), .A2(n8425), .ZN(n8608) );
  NAND2_X1 U7888 ( .A1(n9031), .A2(n8948), .ZN(n8428) );
  NAND2_X1 U7889 ( .A1(n6132), .A2(n8919), .ZN(n8437) );
  INV_X1 U7890 ( .A(n9021), .ZN(n8456) );
  NOR2_X1 U7891 ( .A1(n4864), .A2(n8624), .ZN(n6133) );
  NOR2_X1 U7892 ( .A1(n9011), .A2(n8899), .ZN(n6182) );
  INV_X1 U7893 ( .A(n6182), .ZN(n8464) );
  NAND2_X1 U7894 ( .A1(n9011), .A2(n8899), .ZN(n8463) );
  INV_X1 U7895 ( .A(n9011), .ZN(n8892) );
  NAND2_X1 U7896 ( .A1(n9061), .A2(n8310), .ZN(n6137) );
  NAND2_X1 U7897 ( .A1(n8309), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6136) );
  INV_X1 U7898 ( .A(n8962), .ZN(n8874) );
  NOR2_X1 U7899 ( .A1(n8874), .A2(n8881), .ZN(n6138) );
  NAND2_X1 U7900 ( .A1(n8530), .A2(n8310), .ZN(n6140) );
  NAND2_X1 U7901 ( .A1(n8309), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7902 ( .A1(n6141), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U7903 ( .A1(n8523), .A2(n6142), .ZN(n8517) );
  NAND2_X1 U7904 ( .A1(n8517), .A2(n6143), .ZN(n6148) );
  INV_X1 U7905 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10325) );
  NAND2_X1 U7906 ( .A1(n6161), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6145) );
  INV_X1 U7907 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n10299) );
  OR2_X1 U7908 ( .A1(n4282), .A2(n10299), .ZN(n6144) );
  OAI211_X1 U7909 ( .C1(n5854), .C2(n10325), .A(n6145), .B(n6144), .ZN(n6146)
         );
  INV_X1 U7910 ( .A(n6146), .ZN(n6147) );
  NOR2_X1 U7911 ( .A1(n6348), .A2(n8865), .ZN(n6149) );
  INV_X1 U7912 ( .A(n8865), .ZN(n8476) );
  NAND2_X1 U7913 ( .A1(n8309), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6150) );
  INV_X1 U7914 ( .A(n8523), .ZN(n6152) );
  NAND2_X1 U7915 ( .A1(n6152), .A2(n6143), .ZN(n8318) );
  INV_X1 U7916 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7917 ( .A1(n8311), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U7918 ( .A1(n6161), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6153) );
  OAI211_X1 U7919 ( .C1(n6155), .C2(n4283), .A(n6154), .B(n6153), .ZN(n6156)
         );
  INV_X1 U7920 ( .A(n6156), .ZN(n6157) );
  NAND2_X1 U7921 ( .A1(n8326), .A2(n6366), .ZN(n8322) );
  OR2_X1 U7922 ( .A1(n8479), .A2(n6057), .ZN(n6159) );
  INV_X1 U7923 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n10326) );
  NAND2_X1 U7924 ( .A1(n8311), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7925 ( .A1(n6161), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6162) );
  OAI211_X1 U7926 ( .C1(n4282), .C2(n10326), .A(n6163), .B(n6162), .ZN(n6165)
         );
  INV_X1 U7927 ( .A(n6165), .ZN(n6166) );
  NAND2_X1 U7928 ( .A1(n8318), .A2(n6166), .ZN(n8734) );
  INV_X1 U7929 ( .A(n8734), .ZN(n8279) );
  OAI21_X1 U7930 ( .B1(n5749), .B2(n6168), .A(n10131), .ZN(n8858) );
  OAI22_X1 U7931 ( .A1(n8476), .A2(n8946), .B1(n8279), .B2(n8858), .ZN(n6169)
         );
  NAND2_X1 U7932 ( .A1(n7466), .A2(n7440), .ZN(n8363) );
  NAND2_X1 U7933 ( .A1(n10167), .A2(n8753), .ZN(n7460) );
  NAND2_X1 U7934 ( .A1(n10171), .A2(n8752), .ZN(n8365) );
  NOR2_X1 U7935 ( .A1(n7484), .A2(n7353), .ZN(n7382) );
  NAND2_X1 U7936 ( .A1(n7446), .A2(n7352), .ZN(n8364) );
  NAND2_X1 U7937 ( .A1(n7702), .A2(n7474), .ZN(n8366) );
  NAND2_X1 U7938 ( .A1(n7572), .A2(n7696), .ZN(n8377) );
  INV_X1 U7939 ( .A(n7702), .ZN(n10179) );
  AOI22_X1 U7940 ( .A1(n7803), .A2(n6176), .B1(n8357), .B2(n8750), .ZN(n6177)
         );
  NAND3_X1 U7941 ( .A1(n6178), .A2(n8384), .A3(n6177), .ZN(n6179) );
  NAND2_X1 U7942 ( .A1(n6179), .A2(n8382), .ZN(n7517) );
  OR2_X1 U7943 ( .A1(n7627), .A2(n7923), .ZN(n8385) );
  NAND2_X1 U7944 ( .A1(n7627), .A2(n7923), .ZN(n8386) );
  NAND2_X1 U7945 ( .A1(n8385), .A2(n8386), .ZN(n8289) );
  NAND2_X1 U7946 ( .A1(n5839), .A2(n5836), .ZN(n8391) );
  OR2_X1 U7947 ( .A1(n8185), .A2(n8178), .ZN(n8400) );
  NAND2_X1 U7948 ( .A1(n8185), .A2(n8178), .ZN(n8401) );
  INV_X1 U7949 ( .A(n8400), .ZN(n6180) );
  OR2_X1 U7950 ( .A1(n8597), .A2(n8669), .ZN(n8410) );
  NAND2_X1 U7951 ( .A1(n8716), .A2(n8023), .ZN(n8329) );
  OR2_X1 U7952 ( .A1(n8716), .A2(n8023), .ZN(n8330) );
  NAND2_X1 U7953 ( .A1(n8712), .A2(n8947), .ZN(n8424) );
  NAND2_X1 U7954 ( .A1(n8422), .A2(n8424), .ZN(n8221) );
  AND2_X1 U7955 ( .A1(n8437), .A2(n8428), .ZN(n8430) );
  NAND2_X1 U7956 ( .A1(n9021), .A2(n8920), .ZN(n8442) );
  AND2_X1 U7957 ( .A1(n8457), .A2(n8624), .ZN(n8281) );
  OR2_X1 U7958 ( .A1(n8457), .A2(n8624), .ZN(n8446) );
  OR2_X1 U7959 ( .A1(n8884), .A2(n8570), .ZN(n8468) );
  NAND2_X1 U7960 ( .A1(n8962), .A2(n8881), .ZN(n8472) );
  XNOR2_X1 U7961 ( .A(n6348), .B(n8865), .ZN(n8307) );
  XNOR2_X1 U7962 ( .A(n8321), .B(n8308), .ZN(n8526) );
  NAND2_X1 U7963 ( .A1(n6192), .A2(n10178), .ZN(n7449) );
  NOR2_X1 U7964 ( .A1(n8509), .A2(n8337), .ZN(n6351) );
  INV_X1 U7965 ( .A(n6351), .ZN(n6183) );
  AND2_X1 U7966 ( .A1(n6184), .A2(n6183), .ZN(n6185) );
  INV_X1 U7967 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6197) );
  OR2_X1 U7968 ( .A1(n10184), .A2(n6197), .ZN(n6198) );
  NAND2_X1 U7969 ( .A1(n6199), .A2(n5174), .ZN(P2_U3456) );
  INV_X1 U7970 ( .A(n6230), .ZN(n6200) );
  OR2_X1 U7971 ( .A1(n8499), .A2(n6200), .ZN(n6201) );
  NAND2_X1 U7972 ( .A1(n6201), .A2(n6229), .ZN(n6232) );
  NAND2_X1 U7973 ( .A1(n6232), .A2(n5754), .ZN(n6202) );
  NAND2_X1 U7974 ( .A1(n6202), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U7975 ( .A(n7010), .ZN(n6203) );
  INV_X1 U7976 ( .A(n6319), .ZN(n8794) );
  NOR2_X1 U7977 ( .A1(n6236), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6204) );
  OAI21_X1 U7978 ( .B1(n7143), .B2(n6204), .A(n6205), .ZN(n7142) );
  INV_X1 U7979 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7313) );
  NAND2_X1 U7980 ( .A1(n8762), .A2(n8761), .ZN(n8760) );
  NAND2_X1 U7981 ( .A1(n7015), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7982 ( .A1(n8760), .A2(n6206), .ZN(n6207) );
  XNOR2_X1 U7983 ( .A(n7181), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n7168) );
  OR2_X1 U7984 ( .A1(n7181), .A2(n7464), .ZN(n6209) );
  INV_X1 U7985 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7444) );
  XNOR2_X1 U7986 ( .A(n6304), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n7244) );
  OR2_X1 U7987 ( .A1(n6304), .A2(n7491), .ZN(n6210) );
  INV_X1 U7988 ( .A(n6305), .ZN(n7328) );
  XNOR2_X1 U7989 ( .A(n7016), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n7371) );
  NAND2_X1 U7990 ( .A1(n6212), .A2(n7371), .ZN(n7376) );
  OR2_X1 U7991 ( .A1(n7016), .A2(n7586), .ZN(n6213) );
  XNOR2_X1 U7992 ( .A(n6310), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n7559) );
  INV_X1 U7993 ( .A(n6310), .ZN(n7557) );
  NAND2_X1 U7994 ( .A1(n7557), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6215) );
  OR2_X1 U7995 ( .A1(n7113), .A2(n10223), .ZN(n6217) );
  INV_X1 U7996 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8033) );
  XNOR2_X1 U7997 ( .A(n6319), .B(n8033), .ZN(n8797) );
  XOR2_X1 U7998 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n6322), .Z(n8821) );
  AOI21_X1 U7999 ( .B1(n6221), .B2(n6323), .A(n6222), .ZN(n8841) );
  NAND2_X1 U8000 ( .A1(n8841), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6689) );
  INV_X1 U8001 ( .A(n6222), .ZN(n6691) );
  INV_X1 U8002 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6223) );
  OR2_X1 U8003 ( .A1(n6325), .A2(n6223), .ZN(n6225) );
  NAND2_X1 U8004 ( .A1(n6325), .A2(n6223), .ZN(n6224) );
  NAND2_X1 U8005 ( .A1(n6225), .A2(n6224), .ZN(n6690) );
  INV_X1 U8006 ( .A(n6225), .ZN(n6226) );
  XNOR2_X1 U8007 ( .A(n8509), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n6292) );
  XNOR2_X1 U8008 ( .A(n6227), .B(n6292), .ZN(n6331) );
  AND2_X1 U8009 ( .A1(n8510), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9057) );
  AND2_X1 U8010 ( .A1(n6232), .A2(n9057), .ZN(n7253) );
  INV_X1 U8011 ( .A(n9064), .ZN(n6228) );
  INV_X1 U8012 ( .A(n6229), .ZN(n8116) );
  NOR2_X1 U8013 ( .A1(n6230), .A2(n8116), .ZN(n6231) );
  NAND2_X1 U8014 ( .A1(n6232), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6233) );
  NAND2_X1 U8015 ( .A1(n6233), .A2(n6296), .ZN(n6235) );
  AOI21_X1 U8016 ( .B1(n8742), .B2(n8510), .A(n5749), .ZN(n6234) );
  NAND2_X1 U8017 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8611) );
  OAI21_X1 U8018 ( .B1(n8846), .B2(n7677), .A(n8611), .ZN(n6297) );
  INV_X1 U8019 ( .A(n6325), .ZN(n7497) );
  XNOR2_X1 U8020 ( .A(n6237), .B(n4428), .ZN(n7151) );
  MUX2_X1 U8021 ( .A(n6236), .B(n10187), .S(n9064), .Z(n7251) );
  NAND2_X1 U8022 ( .A1(n7251), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7250) );
  NAND2_X1 U8023 ( .A1(n7151), .A2(n7250), .ZN(n7150) );
  NAND2_X1 U8024 ( .A1(n6237), .A2(n7143), .ZN(n6238) );
  MUX2_X1 U8025 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n9064), .Z(n6239) );
  INV_X1 U8026 ( .A(n7015), .ZN(n8763) );
  XNOR2_X1 U8027 ( .A(n6239), .B(n8763), .ZN(n8768) );
  NAND2_X1 U8028 ( .A1(n6239), .A2(n7015), .ZN(n6240) );
  MUX2_X1 U8029 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n9064), .Z(n6241) );
  XNOR2_X1 U8030 ( .A(n6241), .B(n4286), .ZN(n7099) );
  INV_X1 U8031 ( .A(n6241), .ZN(n6242) );
  NAND2_X1 U8032 ( .A1(n6242), .A2(n6301), .ZN(n6243) );
  AND2_X1 U8033 ( .A1(n7096), .A2(n6243), .ZN(n7184) );
  MUX2_X1 U8034 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n9064), .Z(n6244) );
  XNOR2_X1 U8035 ( .A(n6244), .B(n7181), .ZN(n7183) );
  INV_X1 U8036 ( .A(n7181), .ZN(n6995) );
  NAND2_X1 U8037 ( .A1(n6244), .A2(n6995), .ZN(n6245) );
  MUX2_X1 U8038 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n9064), .Z(n6246) );
  XNOR2_X1 U8039 ( .A(n6246), .B(n6302), .ZN(n7164) );
  MUX2_X1 U8040 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n9064), .Z(n6247) );
  INV_X1 U8041 ( .A(n6304), .ZN(n7235) );
  XNOR2_X1 U8042 ( .A(n6247), .B(n7235), .ZN(n7234) );
  INV_X1 U8043 ( .A(n6247), .ZN(n6248) );
  NAND2_X1 U8044 ( .A1(n6248), .A2(n6304), .ZN(n6249) );
  MUX2_X1 U8045 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n9064), .Z(n6250) );
  XNOR2_X1 U8046 ( .A(n6250), .B(n6305), .ZN(n7326) );
  NAND2_X1 U8047 ( .A1(n7325), .A2(n7326), .ZN(n6253) );
  INV_X1 U8048 ( .A(n6250), .ZN(n6251) );
  NAND2_X1 U8049 ( .A1(n6251), .A2(n6305), .ZN(n6252) );
  NAND2_X1 U8050 ( .A1(n6253), .A2(n6252), .ZN(n7362) );
  MUX2_X1 U8051 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n9064), .Z(n6254) );
  XNOR2_X1 U8052 ( .A(n6254), .B(n7016), .ZN(n7363) );
  NAND2_X1 U8053 ( .A1(n7362), .A2(n7363), .ZN(n6257) );
  INV_X1 U8054 ( .A(n6254), .ZN(n6255) );
  NAND2_X1 U8055 ( .A1(n6255), .A2(n7016), .ZN(n6256) );
  NAND2_X1 U8056 ( .A1(n6257), .A2(n6256), .ZN(n7603) );
  MUX2_X1 U8057 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n9064), .Z(n6258) );
  XNOR2_X1 U8058 ( .A(n6258), .B(n7606), .ZN(n7604) );
  NAND2_X1 U8059 ( .A1(n7603), .A2(n7604), .ZN(n6261) );
  INV_X1 U8060 ( .A(n6258), .ZN(n6259) );
  NAND2_X1 U8061 ( .A1(n6259), .A2(n7606), .ZN(n6260) );
  MUX2_X1 U8062 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n9064), .Z(n6262) );
  XNOR2_X1 U8063 ( .A(n6262), .B(n6310), .ZN(n7553) );
  INV_X1 U8064 ( .A(n6262), .ZN(n6263) );
  MUX2_X1 U8065 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n9064), .Z(n6264) );
  XNOR2_X1 U8066 ( .A(n6264), .B(n8086), .ZN(n8084) );
  INV_X1 U8067 ( .A(n6264), .ZN(n6265) );
  NAND2_X1 U8068 ( .A1(n6265), .A2(n8086), .ZN(n6266) );
  NAND2_X1 U8069 ( .A1(n6267), .A2(n6266), .ZN(n7958) );
  MUX2_X1 U8070 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n9064), .Z(n6268) );
  XNOR2_X1 U8071 ( .A(n6268), .B(n7113), .ZN(n7959) );
  NAND2_X1 U8072 ( .A1(n7958), .A2(n7959), .ZN(n6271) );
  INV_X1 U8073 ( .A(n6268), .ZN(n6269) );
  NAND2_X1 U8074 ( .A1(n6269), .A2(n7113), .ZN(n6270) );
  MUX2_X1 U8075 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n9064), .Z(n6272) );
  XNOR2_X1 U8076 ( .A(n6272), .B(n6315), .ZN(n8774) );
  INV_X1 U8077 ( .A(n6272), .ZN(n6273) );
  NAND2_X1 U8078 ( .A1(n6273), .A2(n6315), .ZN(n6274) );
  MUX2_X1 U8079 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n9064), .Z(n6275) );
  XNOR2_X1 U8080 ( .A(n6275), .B(n6319), .ZN(n8788) );
  INV_X1 U8081 ( .A(n6275), .ZN(n6276) );
  MUX2_X1 U8082 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n9064), .Z(n6277) );
  XNOR2_X1 U8083 ( .A(n6277), .B(n6320), .ZN(n8807) );
  INV_X1 U8084 ( .A(n6277), .ZN(n6278) );
  NAND2_X1 U8085 ( .A1(n6278), .A2(n6320), .ZN(n6279) );
  NAND2_X1 U8086 ( .A1(n6280), .A2(n6279), .ZN(n8828) );
  MUX2_X1 U8087 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n9064), .Z(n6281) );
  XNOR2_X1 U8088 ( .A(n6281), .B(n6322), .ZN(n8829) );
  NAND2_X1 U8089 ( .A1(n8828), .A2(n8829), .ZN(n6284) );
  INV_X1 U8090 ( .A(n6281), .ZN(n6282) );
  NAND2_X1 U8091 ( .A1(n6282), .A2(n6322), .ZN(n6283) );
  NAND2_X1 U8092 ( .A1(n6284), .A2(n6283), .ZN(n8842) );
  MUX2_X1 U8093 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n9064), .Z(n6285) );
  XNOR2_X1 U8094 ( .A(n6285), .B(n6323), .ZN(n8843) );
  INV_X1 U8095 ( .A(n6285), .ZN(n6286) );
  AND2_X1 U8096 ( .A1(n6286), .A2(n6323), .ZN(n6287) );
  AOI21_X1 U8097 ( .B1(n8842), .B2(n8843), .A(n6287), .ZN(n6291) );
  INV_X1 U8098 ( .A(n6291), .ZN(n6289) );
  MUX2_X1 U8099 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n9064), .Z(n6290) );
  INV_X1 U8100 ( .A(n6290), .ZN(n6288) );
  NAND2_X1 U8101 ( .A1(n6289), .A2(n6288), .ZN(n6694) );
  AND2_X1 U8102 ( .A1(n6291), .A2(n6290), .ZN(n6696) );
  INV_X1 U8103 ( .A(n6292), .ZN(n6294) );
  XNOR2_X1 U8104 ( .A(n8509), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n6329) );
  INV_X1 U8105 ( .A(n6329), .ZN(n6293) );
  MUX2_X1 U8106 ( .A(n6294), .B(n6293), .S(n9064), .Z(n6295) );
  INV_X1 U8107 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8163) );
  INV_X1 U8108 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6318) );
  INV_X1 U8109 ( .A(n6298), .ZN(n6299) );
  XNOR2_X1 U8110 ( .A(n7181), .B(n10193), .ZN(n7174) );
  XNOR2_X1 U8111 ( .A(n6304), .B(n10197), .ZN(n7238) );
  XNOR2_X1 U8112 ( .A(n7016), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n7365) );
  XNOR2_X1 U8113 ( .A(n6310), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n7554) );
  INV_X1 U8114 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7715) );
  NAND2_X1 U8115 ( .A1(n7557), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U8116 ( .A1(n6312), .A2(n7044), .ZN(n6313) );
  INV_X1 U8117 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8090) );
  INV_X1 U8118 ( .A(n6313), .ZN(n7963) );
  XNOR2_X1 U8119 ( .A(n7113), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n7962) );
  INV_X1 U8120 ( .A(n6315), .ZN(n8778) );
  INV_X1 U8121 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8780) );
  XNOR2_X1 U8122 ( .A(n6319), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n8789) );
  INV_X1 U8123 ( .A(n6320), .ZN(n8815) );
  INV_X1 U8124 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8149) );
  XNOR2_X1 U8125 ( .A(n6322), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8824) );
  INV_X1 U8126 ( .A(n6323), .ZN(n8845) );
  INV_X1 U8127 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8840) );
  OR2_X1 U8128 ( .A1(n6325), .A2(n10275), .ZN(n6327) );
  NAND2_X1 U8129 ( .A1(n6325), .A2(n10275), .ZN(n6326) );
  NAND2_X1 U8130 ( .A1(n6327), .A2(n6326), .ZN(n6683) );
  AOI21_X1 U8131 ( .B1(n8837), .B2(n6684), .A(n6683), .ZN(n6682) );
  INV_X1 U8132 ( .A(n6327), .ZN(n6328) );
  XNOR2_X1 U8133 ( .A(n6332), .B(n8899), .ZN(n8619) );
  AOI21_X1 U8134 ( .B1(n8620), .B2(n8618), .A(n8619), .ZN(n8621) );
  INV_X1 U8135 ( .A(n6333), .ZN(n6335) );
  OAI21_X1 U8136 ( .B1(n8621), .B2(n6335), .A(n6334), .ZN(n6336) );
  XNOR2_X1 U8137 ( .A(n8962), .B(n6338), .ZN(n6344) );
  XNOR2_X1 U8138 ( .A(n6344), .B(n8881), .ZN(n8566) );
  XNOR2_X1 U8139 ( .A(n8865), .B(n4706), .ZN(n6340) );
  XNOR2_X1 U8140 ( .A(n6348), .B(n6340), .ZN(n6341) );
  INV_X1 U8141 ( .A(n6341), .ZN(n6345) );
  OAI211_X1 U8142 ( .C1(n8881), .C2(n6344), .A(n6345), .B(n8679), .ZN(n6350)
         );
  INV_X1 U8143 ( .A(n6366), .ZN(n8735) );
  NAND2_X1 U8144 ( .A1(n8735), .A2(n8704), .ZN(n6343) );
  AOI22_X1 U8145 ( .A1(n8517), .A2(n8727), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n6342) );
  OAI211_X1 U8146 ( .C1(n8881), .C2(n8707), .A(n6343), .B(n6342), .ZN(n6347)
         );
  NOR4_X1 U8147 ( .A1(n6345), .A2(n6344), .A3(n8881), .A4(n8717), .ZN(n6346)
         );
  AOI211_X1 U8148 ( .C1(n6348), .C2(n8711), .A(n6347), .B(n6346), .ZN(n6349)
         );
  AND2_X1 U8149 ( .A1(n6351), .A2(n8500), .ZN(n6352) );
  NAND2_X1 U8150 ( .A1(n6353), .A2(n6044), .ZN(n6354) );
  NAND2_X1 U8151 ( .A1(n7303), .A2(n6354), .ZN(n6357) );
  INV_X1 U8152 ( .A(n7303), .ZN(n6355) );
  NAND2_X1 U8153 ( .A1(n6355), .A2(n7300), .ZN(n6356) );
  NAND2_X1 U8154 ( .A1(n6362), .A2(n10199), .ZN(n6364) );
  NAND2_X1 U8155 ( .A1(n6372), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6363) );
  NAND2_X1 U8156 ( .A1(n6364), .A2(n5167), .ZN(P2_U3488) );
  XNOR2_X1 U8157 ( .A(n6365), .B(n5065), .ZN(n6368) );
  OAI22_X1 U8158 ( .A1(n6366), .A2(n4652), .B1(n8881), .B2(n8946), .ZN(n6367)
         );
  OAI21_X1 U8159 ( .B1(n6370), .B2(n8307), .A(n6369), .ZN(n8521) );
  NAND2_X1 U8160 ( .A1(n5186), .A2(n5173), .ZN(P2_U3487) );
  NAND2_X1 U8161 ( .A1(n6373), .A2(n10184), .ZN(n6377) );
  NOR2_X1 U8162 ( .A1(n10184), .A2(n10325), .ZN(n6374) );
  NAND2_X1 U8163 ( .A1(n6377), .A2(n6376), .ZN(P2_U3455) );
  AND2_X1 U8164 ( .A1(n6971), .A2(n4796), .ZN(n6378) );
  OR3_X2 U8165 ( .A1(n6379), .A2(n6378), .A3(n9864), .ZN(n9605) );
  INV_X1 U8166 ( .A(n6380), .ZN(n9598) );
  NAND2_X1 U8167 ( .A1(n9605), .A2(n9598), .ZN(n6383) );
  MUX2_X1 U8168 ( .A(n6383), .B(P1_REG1_REG_30__SCAN_IN), .S(n10120), .Z(n6382) );
  MUX2_X1 U8169 ( .A(n6383), .B(P1_REG0_REG_30__SCAN_IN), .S(n10113), .Z(n6385) );
  INV_X1 U8170 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6626) );
  NAND2_X1 U8171 ( .A1(n6589), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6398) );
  INV_X1 U8172 ( .A(n6436), .ZN(n6386) );
  NAND2_X1 U8173 ( .A1(n6386), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6455) );
  INV_X1 U8174 ( .A(n6455), .ZN(n6388) );
  NAND2_X1 U8175 ( .A1(n6388), .A2(n6387), .ZN(n6457) );
  INV_X1 U8176 ( .A(n6457), .ZN(n6389) );
  INV_X1 U8177 ( .A(n6391), .ZN(n6401) );
  INV_X1 U8178 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6392) );
  NAND2_X1 U8179 ( .A1(n6401), .A2(n6392), .ZN(n6393) );
  AND2_X1 U8180 ( .A1(n6507), .A2(n6393), .ZN(n9818) );
  NAND2_X1 U8181 ( .A1(n9818), .A2(n6588), .ZN(n6397) );
  NAND2_X1 U8182 ( .A1(n6959), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6396) );
  NAND2_X1 U8183 ( .A1(n6563), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6395) );
  NAND4_X1 U8184 ( .A1(n6398), .A2(n6397), .A3(n6396), .A4(n6395), .ZN(n9833)
         );
  INV_X1 U8185 ( .A(n9833), .ZN(n9799) );
  OR2_X1 U8186 ( .A1(n9820), .A2(n9799), .ZN(n9387) );
  NAND2_X1 U8187 ( .A1(n9820), .A2(n9799), .ZN(n9232) );
  NAND2_X1 U8188 ( .A1(n6959), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U8189 ( .A1(n6589), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6404) );
  NAND2_X1 U8190 ( .A1(n6496), .A2(n6399), .ZN(n6400) );
  AND2_X1 U8191 ( .A1(n6401), .A2(n6400), .ZN(n9843) );
  NAND2_X1 U8192 ( .A1(n6588), .A2(n9843), .ZN(n6403) );
  NAND2_X1 U8193 ( .A1(n6563), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6402) );
  OR2_X1 U8194 ( .A1(n9924), .A2(n9807), .ZN(n9810) );
  NAND2_X1 U8195 ( .A1(n6588), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6409) );
  NAND2_X1 U8196 ( .A1(n6416), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6408) );
  NAND2_X1 U8197 ( .A1(n6422), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U8198 ( .A1(n6423), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6406) );
  NAND4_X2 U8199 ( .A1(n6409), .A2(n6408), .A3(n6407), .A4(n6406), .ZN(n6725)
         );
  INV_X1 U8200 ( .A(n6627), .ZN(n7399) );
  NAND2_X1 U8201 ( .A1(n6423), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U8202 ( .A1(n6416), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6412) );
  NAND2_X1 U8203 ( .A1(n6422), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6410) );
  NAND4_X2 U8204 ( .A1(n6413), .A2(n6412), .A3(n6411), .A4(n6410), .ZN(n6739)
         );
  NAND2_X1 U8205 ( .A1(n7399), .A2(n7402), .ZN(n6415) );
  INV_X1 U8206 ( .A(n6725), .ZN(n7539) );
  NAND2_X1 U8207 ( .A1(n7539), .A2(n6726), .ZN(n6414) );
  NAND2_X1 U8208 ( .A1(n6415), .A2(n6414), .ZN(n7416) );
  NAND2_X1 U8209 ( .A1(n6588), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U8210 ( .A1(n6416), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6419) );
  NAND2_X1 U8211 ( .A1(n6422), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6418) );
  NAND2_X1 U8212 ( .A1(n6423), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6417) );
  NAND4_X2 U8213 ( .A1(n6420), .A2(n6419), .A3(n6418), .A4(n6417), .ZN(n9431)
         );
  XNOR2_X1 U8214 ( .A(n9431), .B(n9363), .ZN(n9279) );
  INV_X1 U8215 ( .A(n9431), .ZN(n9364) );
  NAND2_X1 U8216 ( .A1(n9364), .A2(n9363), .ZN(n6421) );
  NAND2_X1 U8217 ( .A1(n6422), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6426) );
  INV_X1 U8218 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7595) );
  NAND2_X1 U8219 ( .A1(n6588), .A2(n7595), .ZN(n6425) );
  NAND2_X1 U8220 ( .A1(n6423), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6424) );
  NAND2_X1 U8221 ( .A1(n9430), .A2(n10089), .ZN(n9369) );
  INV_X1 U8222 ( .A(n10089), .ZN(n7672) );
  NAND2_X1 U8223 ( .A1(n7646), .A2(n7672), .ZN(n6428) );
  NAND2_X1 U8224 ( .A1(n6959), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6434) );
  NAND2_X1 U8225 ( .A1(n6416), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6433) );
  INV_X1 U8226 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6429) );
  NAND2_X1 U8227 ( .A1(n7595), .A2(n6429), .ZN(n6430) );
  AND2_X1 U8228 ( .A1(n6430), .A2(n6436), .ZN(n9135) );
  NAND2_X1 U8229 ( .A1(n6588), .A2(n9135), .ZN(n6432) );
  NAND2_X1 U8230 ( .A1(n6960), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6431) );
  NAND2_X1 U8231 ( .A1(n9429), .A2(n10095), .ZN(n9368) );
  NAND2_X1 U8232 ( .A1(n7644), .A2(n9368), .ZN(n9196) );
  NAND2_X1 U8233 ( .A1(n7666), .A2(n9134), .ZN(n9194) );
  NAND2_X1 U8234 ( .A1(n9196), .A2(n9194), .ZN(n7902) );
  NAND2_X1 U8235 ( .A1(n6959), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6441) );
  NAND2_X1 U8236 ( .A1(n6416), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6440) );
  INV_X1 U8237 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6435) );
  NAND2_X1 U8238 ( .A1(n6436), .A2(n6435), .ZN(n6437) );
  AND2_X1 U8239 ( .A1(n6455), .A2(n6437), .ZN(n7899) );
  NAND2_X1 U8240 ( .A1(n6588), .A2(n7899), .ZN(n6439) );
  NAND2_X1 U8241 ( .A1(n6563), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6438) );
  INV_X1 U8242 ( .A(n7900), .ZN(n10101) );
  NAND2_X1 U8243 ( .A1(n6416), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6446) );
  XNOR2_X1 U8244 ( .A(n6455), .B(P1_REG3_REG_6__SCAN_IN), .ZN(n7826) );
  NAND2_X1 U8245 ( .A1(n6588), .A2(n7826), .ZN(n6445) );
  NAND2_X1 U8246 ( .A1(n6959), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6444) );
  NAND2_X1 U8247 ( .A1(n6960), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6443) );
  NAND2_X1 U8248 ( .A1(n9200), .A2(n9199), .ZN(n9190) );
  INV_X1 U8249 ( .A(n9190), .ZN(n9285) );
  NAND2_X1 U8250 ( .A1(n6959), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6452) );
  INV_X2 U8251 ( .A(n6582), .ZN(n6961) );
  NAND2_X1 U8252 ( .A1(n6961), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6451) );
  INV_X1 U8253 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U8254 ( .A1(n6457), .A2(n6447), .ZN(n6448) );
  AND2_X1 U8255 ( .A1(n6463), .A2(n6448), .ZN(n8074) );
  NAND2_X1 U8256 ( .A1(n6588), .A2(n8074), .ZN(n6450) );
  NAND2_X1 U8257 ( .A1(n6563), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6449) );
  NAND2_X1 U8258 ( .A1(n8075), .A2(n7530), .ZN(n9212) );
  NAND2_X1 U8259 ( .A1(n6589), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6461) );
  INV_X1 U8260 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6454) );
  INV_X1 U8261 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6453) );
  OAI21_X1 U8262 ( .B1(n6455), .B2(n6454), .A(n6453), .ZN(n6456) );
  AND2_X1 U8263 ( .A1(n6457), .A2(n6456), .ZN(n7910) );
  NAND2_X1 U8264 ( .A1(n6588), .A2(n7910), .ZN(n6460) );
  NAND2_X1 U8265 ( .A1(n6959), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6459) );
  NAND2_X1 U8266 ( .A1(n6960), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U8267 ( .A1(n7911), .A2(n7998), .ZN(n7992) );
  NAND2_X1 U8268 ( .A1(n9212), .A2(n7992), .ZN(n7788) );
  NAND2_X1 U8269 ( .A1(n7788), .A2(n9211), .ZN(n6469) );
  NAND2_X1 U8270 ( .A1(n6959), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U8271 ( .A1(n6961), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U8272 ( .A1(n6463), .A2(n6462), .ZN(n6464) );
  AND2_X1 U8273 ( .A1(n6472), .A2(n6464), .ZN(n7890) );
  NAND2_X1 U8274 ( .A1(n6588), .A2(n7890), .ZN(n6466) );
  NAND2_X1 U8275 ( .A1(n6960), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6465) );
  NAND2_X1 U8276 ( .A1(n6469), .A2(n9286), .ZN(n6470) );
  OR2_X1 U8277 ( .A1(n7875), .A2(n7997), .ZN(n9218) );
  NAND2_X1 U8278 ( .A1(n6470), .A2(n9218), .ZN(n9373) );
  OR2_X1 U8279 ( .A1(n7998), .A2(n7911), .ZN(n6635) );
  INV_X1 U8280 ( .A(n9199), .ZN(n10108) );
  NAND2_X1 U8281 ( .A1(n10108), .A2(n9427), .ZN(n9197) );
  NAND2_X1 U8282 ( .A1(n9373), .A2(n9374), .ZN(n7763) );
  NAND2_X1 U8283 ( .A1(n6959), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U8284 ( .A1(n6961), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6476) );
  INV_X1 U8285 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U8286 ( .A1(n6472), .A2(n6471), .ZN(n6473) );
  AND2_X1 U8287 ( .A1(n6478), .A2(n6473), .ZN(n7984) );
  NAND2_X1 U8288 ( .A1(n6588), .A2(n7984), .ZN(n6475) );
  NAND2_X1 U8289 ( .A1(n6960), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6474) );
  NAND3_X1 U8290 ( .A1(n9372), .A2(n7763), .A3(n9377), .ZN(n6485) );
  NAND2_X1 U8291 ( .A1(n6589), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U8292 ( .A1(n6478), .A2(n7079), .ZN(n6479) );
  AND2_X1 U8293 ( .A1(n6487), .A2(n6479), .ZN(n8067) );
  NAND2_X1 U8294 ( .A1(n6588), .A2(n8067), .ZN(n6482) );
  NAND2_X1 U8295 ( .A1(n6959), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6481) );
  NAND2_X1 U8296 ( .A1(n6960), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U8297 ( .A1(n6484), .A2(n7981), .ZN(n9222) );
  INV_X1 U8298 ( .A(n7835), .ZN(n9293) );
  NAND2_X1 U8299 ( .A1(n7769), .A2(n7888), .ZN(n9220) );
  INV_X1 U8300 ( .A(n7788), .ZN(n9288) );
  NAND2_X1 U8301 ( .A1(n9286), .A2(n9288), .ZN(n7764) );
  NAND2_X1 U8302 ( .A1(n6961), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6492) );
  NAND2_X1 U8303 ( .A1(n6959), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6491) );
  INV_X1 U8304 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U8305 ( .A1(n6487), .A2(n6486), .ZN(n6488) );
  AND2_X1 U8306 ( .A1(n6494), .A2(n6488), .ZN(n8048) );
  NAND2_X1 U8307 ( .A1(n6588), .A2(n8048), .ZN(n6490) );
  NAND2_X1 U8308 ( .A1(n6563), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6489) );
  OR2_X1 U8309 ( .A1(n6837), .A2(n9422), .ZN(n9224) );
  NAND2_X1 U8310 ( .A1(n6837), .A2(n9422), .ZN(n9380) );
  NAND2_X1 U8311 ( .A1(n6959), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6500) );
  NAND2_X1 U8312 ( .A1(n6961), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6499) );
  NAND2_X1 U8313 ( .A1(n6494), .A2(n6493), .ZN(n6495) );
  AND2_X1 U8314 ( .A1(n6496), .A2(n6495), .ZN(n8268) );
  NAND2_X1 U8315 ( .A1(n6588), .A2(n8268), .ZN(n6498) );
  NAND2_X1 U8316 ( .A1(n6563), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6497) );
  NAND4_X1 U8317 ( .A1(n6500), .A2(n6499), .A3(n6498), .A4(n6497), .ZN(n9835)
         );
  XNOR2_X1 U8318 ( .A(n9228), .B(n9835), .ZN(n9296) );
  INV_X1 U8319 ( .A(n9835), .ZN(n9227) );
  NAND2_X1 U8320 ( .A1(n9228), .A2(n9227), .ZN(n9827) );
  XNOR2_X1 U8321 ( .A(n9924), .B(n9807), .ZN(n9230) );
  AND2_X1 U8322 ( .A1(n9827), .A2(n9831), .ZN(n6501) );
  NAND2_X1 U8323 ( .A1(n9811), .A2(n9232), .ZN(n9796) );
  NAND2_X1 U8324 ( .A1(n6959), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U8325 ( .A1(n6589), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6503) );
  AND2_X1 U8326 ( .A1(n6504), .A2(n6503), .ZN(n6511) );
  INV_X1 U8327 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U8328 ( .A1(n6507), .A2(n6506), .ZN(n6508) );
  NAND2_X1 U8329 ( .A1(n6513), .A2(n6508), .ZN(n9792) );
  OR2_X1 U8330 ( .A1(n6615), .A2(n9792), .ZN(n6510) );
  NAND2_X1 U8331 ( .A1(n6563), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U8332 ( .A1(n9911), .A2(n9180), .ZN(n9233) );
  NAND2_X1 U8333 ( .A1(n6513), .A2(n6512), .ZN(n6514) );
  AND2_X1 U8334 ( .A1(n6519), .A2(n6514), .ZN(n9780) );
  NAND2_X1 U8335 ( .A1(n9780), .A2(n6588), .ZN(n6517) );
  AOI22_X1 U8336 ( .A1(n6959), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n6589), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n6516) );
  NAND2_X1 U8337 ( .A1(n6563), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6515) );
  OR2_X1 U8338 ( .A1(n9906), .A2(n9801), .ZN(n9243) );
  NAND2_X1 U8339 ( .A1(n9906), .A2(n9801), .ZN(n9239) );
  INV_X1 U8340 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9571) );
  INV_X1 U8341 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6518) );
  NAND2_X1 U8342 ( .A1(n6519), .A2(n6518), .ZN(n6520) );
  NAND2_X1 U8343 ( .A1(n6526), .A2(n6520), .ZN(n9760) );
  OR2_X1 U8344 ( .A1(n9760), .A2(n6615), .ZN(n6522) );
  AOI22_X1 U8345 ( .A1(n6959), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n6961), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n6521) );
  OAI211_X1 U8346 ( .C1(n6442), .C2(n9571), .A(n6522), .B(n6521), .ZN(n9776)
         );
  INV_X1 U8347 ( .A(n9776), .ZN(n9115) );
  OR2_X1 U8348 ( .A1(n9900), .A2(n9115), .ZN(n9396) );
  NAND2_X1 U8349 ( .A1(n9900), .A2(n9115), .ZN(n9244) );
  NAND2_X1 U8350 ( .A1(n6524), .A2(n6523), .ZN(n9893) );
  NAND2_X1 U8351 ( .A1(n6526), .A2(n6525), .ZN(n6527) );
  AND2_X1 U8352 ( .A1(n6537), .A2(n6527), .ZN(n9747) );
  NAND2_X1 U8353 ( .A1(n9747), .A2(n6588), .ZN(n6533) );
  INV_X1 U8354 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n6530) );
  NAND2_X1 U8355 ( .A1(n6959), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6529) );
  NAND2_X1 U8356 ( .A1(n6961), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6528) );
  OAI211_X1 U8357 ( .C1(n6530), .C2(n6442), .A(n6529), .B(n6528), .ZN(n6531)
         );
  INV_X1 U8358 ( .A(n6531), .ZN(n6532) );
  OR2_X1 U8359 ( .A1(n9893), .A2(n9728), .ZN(n9395) );
  NAND2_X1 U8360 ( .A1(n9893), .A2(n9728), .ZN(n9401) );
  INV_X1 U8361 ( .A(n9401), .ZN(n6534) );
  INV_X1 U8362 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6536) );
  NAND2_X1 U8363 ( .A1(n6537), .A2(n6536), .ZN(n6538) );
  NAND2_X1 U8364 ( .A1(n6553), .A2(n6538), .ZN(n9145) );
  OR2_X1 U8365 ( .A1(n9145), .A2(n6615), .ZN(n6543) );
  INV_X1 U8366 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9891) );
  NAND2_X1 U8367 ( .A1(n6563), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6540) );
  NAND2_X1 U8368 ( .A1(n6589), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6539) );
  OAI211_X1 U8369 ( .C1(n6618), .C2(n9891), .A(n6540), .B(n6539), .ZN(n6541)
         );
  INV_X1 U8370 ( .A(n6541), .ZN(n6542) );
  NAND2_X1 U8371 ( .A1(n6543), .A2(n6542), .ZN(n9752) );
  INV_X1 U8372 ( .A(n9752), .ZN(n9078) );
  NAND2_X1 U8373 ( .A1(n9734), .A2(n9078), .ZN(n9246) );
  XNOR2_X1 U8374 ( .A(n6553), .B(P1_REG3_REG_21__SCAN_IN), .ZN(n9718) );
  NAND2_X1 U8375 ( .A1(n9718), .A2(n6588), .ZN(n6549) );
  INV_X1 U8376 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U8377 ( .A1(n6959), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6545) );
  NAND2_X1 U8378 ( .A1(n6961), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6544) );
  OAI211_X1 U8379 ( .C1(n6546), .C2(n6442), .A(n6545), .B(n6544), .ZN(n6547)
         );
  INV_X1 U8380 ( .A(n6547), .ZN(n6548) );
  NAND2_X1 U8381 ( .A1(n9955), .A2(n9729), .ZN(n9683) );
  INV_X1 U8382 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6551) );
  INV_X1 U8383 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6550) );
  OAI21_X1 U8384 ( .B1(n6553), .B2(n6551), .A(n6550), .ZN(n6554) );
  NAND2_X1 U8385 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .ZN(n6552) );
  NAND2_X1 U8386 ( .A1(n6554), .A2(n6561), .ZN(n9695) );
  OR2_X1 U8387 ( .A1(n9695), .A2(n6615), .ZN(n6559) );
  INV_X1 U8388 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10291) );
  NAND2_X1 U8389 ( .A1(n6563), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U8390 ( .A1(n6589), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6555) );
  OAI211_X1 U8391 ( .C1(n6618), .C2(n10291), .A(n6556), .B(n6555), .ZN(n6557)
         );
  INV_X1 U8392 ( .A(n6557), .ZN(n6558) );
  NAND2_X1 U8393 ( .A1(n6559), .A2(n6558), .ZN(n9714) );
  XNOR2_X1 U8394 ( .A(n9877), .B(n9714), .ZN(n9690) );
  NAND2_X1 U8395 ( .A1(n9877), .A2(n9253), .ZN(n9670) );
  INV_X1 U8396 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6560) );
  NAND2_X1 U8397 ( .A1(n6561), .A2(n6560), .ZN(n6562) );
  NAND2_X1 U8398 ( .A1(n6571), .A2(n6562), .ZN(n9676) );
  OR2_X1 U8399 ( .A1(n9676), .A2(n6615), .ZN(n6568) );
  INV_X1 U8400 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9872) );
  NAND2_X1 U8401 ( .A1(n6589), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6565) );
  NAND2_X1 U8402 ( .A1(n6563), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6564) );
  OAI211_X1 U8403 ( .C1(n6618), .C2(n9872), .A(n6565), .B(n6564), .ZN(n6566)
         );
  INV_X1 U8404 ( .A(n6566), .ZN(n6567) );
  OR2_X1 U8405 ( .A1(n9947), .A2(n9652), .ZN(n9259) );
  NAND2_X1 U8406 ( .A1(n9259), .A2(n9313), .ZN(n9669) );
  INV_X1 U8407 ( .A(n9313), .ZN(n9649) );
  INV_X1 U8408 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6570) );
  NAND2_X1 U8409 ( .A1(n6571), .A2(n6570), .ZN(n6572) );
  NAND2_X1 U8410 ( .A1(n6578), .A2(n6572), .ZN(n9658) );
  OR2_X1 U8411 ( .A1(n9658), .A2(n6615), .ZN(n6577) );
  INV_X1 U8412 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9868) );
  NAND2_X1 U8413 ( .A1(n6589), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6574) );
  NAND2_X1 U8414 ( .A1(n6960), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6573) );
  OAI211_X1 U8415 ( .C1(n6618), .C2(n9868), .A(n6574), .B(n6573), .ZN(n6575)
         );
  INV_X1 U8416 ( .A(n6575), .ZN(n6576) );
  INV_X1 U8417 ( .A(n9673), .ZN(n6658) );
  OR2_X1 U8418 ( .A1(n9660), .A2(n6658), .ZN(n9316) );
  NAND2_X1 U8419 ( .A1(n9660), .A2(n6658), .ZN(n9325) );
  NAND2_X1 U8420 ( .A1(n9316), .A2(n9325), .ZN(n9303) );
  INV_X1 U8421 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U8422 ( .A1(n6578), .A2(n9094), .ZN(n6579) );
  NAND2_X1 U8423 ( .A1(n6586), .A2(n6579), .ZN(n9642) );
  INV_X1 U8424 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10356) );
  NAND2_X1 U8425 ( .A1(n6959), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6581) );
  NAND2_X1 U8426 ( .A1(n6960), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6580) );
  OAI211_X1 U8427 ( .C1(n6582), .C2(n10356), .A(n6581), .B(n6580), .ZN(n6583)
         );
  INV_X1 U8428 ( .A(n6583), .ZN(n6584) );
  OR2_X1 U8429 ( .A1(n9644), .A2(n9653), .ZN(n9319) );
  NAND2_X1 U8430 ( .A1(n9644), .A2(n9653), .ZN(n9262) );
  INV_X1 U8431 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8275) );
  NAND2_X1 U8432 ( .A1(n6586), .A2(n8275), .ZN(n6587) );
  NAND2_X1 U8433 ( .A1(n9623), .A2(n6588), .ZN(n6595) );
  INV_X1 U8434 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n6592) );
  NAND2_X1 U8435 ( .A1(n6589), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6591) );
  NAND2_X1 U8436 ( .A1(n6960), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6590) );
  OAI211_X1 U8437 ( .C1(n6618), .C2(n6592), .A(n6591), .B(n6590), .ZN(n6593)
         );
  INV_X1 U8438 ( .A(n6593), .ZN(n6594) );
  NAND2_X1 U8439 ( .A1(n9855), .A2(n6909), .ZN(n9322) );
  INV_X1 U8440 ( .A(n6597), .ZN(n6596) );
  NAND2_X1 U8441 ( .A1(n6596), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6606) );
  INV_X1 U8442 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n10278) );
  NAND2_X1 U8443 ( .A1(n6597), .A2(n10278), .ZN(n6598) );
  NAND2_X1 U8444 ( .A1(n6606), .A2(n6598), .ZN(n9607) );
  INV_X1 U8445 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n10293) );
  NAND2_X1 U8446 ( .A1(n6961), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6600) );
  NAND2_X1 U8447 ( .A1(n6960), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6599) );
  OAI211_X1 U8448 ( .C1(n6618), .C2(n10293), .A(n6600), .B(n6599), .ZN(n6601)
         );
  INV_X1 U8449 ( .A(n6601), .ZN(n6602) );
  AND2_X2 U8450 ( .A1(n6603), .A2(n6602), .ZN(n10374) );
  NAND2_X1 U8451 ( .A1(n9609), .A2(n10374), .ZN(n6955) );
  NAND2_X1 U8452 ( .A1(n9312), .A2(n6955), .ZN(n9305) );
  INV_X1 U8453 ( .A(n6606), .ZN(n6604) );
  NAND2_X1 U8454 ( .A1(n6604), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8533) );
  INV_X1 U8455 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6605) );
  NAND2_X1 U8456 ( .A1(n6606), .A2(n6605), .ZN(n6607) );
  NAND2_X1 U8457 ( .A1(n8533), .A2(n6607), .ZN(n8579) );
  NAND2_X1 U8458 ( .A1(n6961), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6609) );
  NAND2_X1 U8459 ( .A1(n6960), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6608) );
  OAI211_X1 U8460 ( .C1(n6618), .C2(n6626), .A(n6609), .B(n6608), .ZN(n6610)
         );
  INV_X1 U8461 ( .A(n6610), .ZN(n6611) );
  NAND2_X1 U8462 ( .A1(n8581), .A2(n8550), .ZN(n6956) );
  NAND2_X1 U8463 ( .A1(n9336), .A2(n6956), .ZN(n9306) );
  NAND2_X1 U8464 ( .A1(n6666), .A2(n9677), .ZN(n9275) );
  NAND2_X1 U8465 ( .A1(n6669), .A2(n9349), .ZN(n9353) );
  OR2_X1 U8466 ( .A1(n8533), .A2(n6615), .ZN(n6621) );
  INV_X1 U8467 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6974) );
  NAND2_X1 U8468 ( .A1(n6960), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6617) );
  NAND2_X1 U8469 ( .A1(n6961), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6616) );
  OAI211_X1 U8470 ( .C1(n6618), .C2(n6974), .A(n6617), .B(n6616), .ZN(n6619)
         );
  INV_X1 U8471 ( .A(n6619), .ZN(n6620) );
  NAND2_X1 U8472 ( .A1(n9420), .A2(n9834), .ZN(n6623) );
  INV_X1 U8473 ( .A(n8531), .ZN(n9455) );
  NAND2_X1 U8474 ( .A1(n9628), .A2(n9836), .ZN(n6622) );
  AOI21_X1 U8475 ( .B1(n6625), .B2(n9829), .A(n6624), .ZN(n8587) );
  OAI211_X1 U8476 ( .C1(n6975), .C2(n6712), .A(n9894), .B(n6970), .ZN(n8583)
         );
  AND2_X1 U8477 ( .A1(n8587), .A2(n8583), .ZN(n6676) );
  MUX2_X1 U8478 ( .A(n6626), .B(n6676), .S(n10123), .Z(n6675) );
  NAND2_X1 U8479 ( .A1(n6739), .A2(n7651), .ZN(n7401) );
  NAND2_X1 U8480 ( .A1(n7539), .A2(n10080), .ZN(n6628) );
  NAND2_X1 U8481 ( .A1(n7400), .A2(n6628), .ZN(n7412) );
  NAND2_X1 U8482 ( .A1(n9364), .A2(n6750), .ZN(n6629) );
  NAND2_X1 U8483 ( .A1(n7411), .A2(n6629), .ZN(n7663) );
  XNOR2_X1 U8484 ( .A(n9430), .B(n10089), .ZN(n9282) );
  NAND2_X1 U8485 ( .A1(n7663), .A2(n9282), .ZN(n7662) );
  NAND2_X1 U8486 ( .A1(n7646), .A2(n10089), .ZN(n6630) );
  XNOR2_X1 U8487 ( .A(n9429), .B(n10095), .ZN(n9284) );
  AND2_X1 U8488 ( .A1(n9284), .A2(n9281), .ZN(n6631) );
  NAND2_X1 U8489 ( .A1(n7639), .A2(n6631), .ZN(n6633) );
  NAND2_X1 U8490 ( .A1(n7666), .A2(n10095), .ZN(n7893) );
  OR2_X1 U8491 ( .A1(n7903), .A2(n7893), .ZN(n6632) );
  NAND2_X1 U8492 ( .A1(n7647), .A2(n10101), .ZN(n6634) );
  NAND2_X1 U8493 ( .A1(n7895), .A2(n6634), .ZN(n7822) );
  NAND2_X1 U8494 ( .A1(n9190), .A2(n9197), .ZN(n7821) );
  NAND2_X1 U8495 ( .A1(n6635), .A2(n7992), .ZN(n9201) );
  AND2_X1 U8496 ( .A1(n7821), .A2(n9201), .ZN(n6637) );
  INV_X1 U8497 ( .A(n9201), .ZN(n6636) );
  NAND2_X1 U8498 ( .A1(n9200), .A2(n10108), .ZN(n7747) );
  OR2_X1 U8499 ( .A1(n9426), .A2(n7911), .ZN(n6638) );
  NAND2_X1 U8500 ( .A1(n9211), .A2(n9212), .ZN(n7994) );
  NAND2_X1 U8501 ( .A1(n9218), .A2(n9286), .ZN(n7793) );
  AND2_X1 U8502 ( .A1(n7994), .A2(n7793), .ZN(n6640) );
  INV_X1 U8503 ( .A(n7793), .ZN(n6639) );
  OR2_X1 U8504 ( .A1(n8075), .A2(n4580), .ZN(n7791) );
  INV_X1 U8505 ( .A(n7997), .ZN(n9425) );
  OR2_X1 U8506 ( .A1(n7875), .A2(n9425), .ZN(n6641) );
  NAND2_X1 U8507 ( .A1(n9377), .A2(n9220), .ZN(n9278) );
  INV_X1 U8508 ( .A(n7888), .ZN(n9424) );
  OR2_X1 U8509 ( .A1(n7769), .A2(n9424), .ZN(n6642) );
  NOR2_X1 U8510 ( .A1(n9924), .A2(n9814), .ZN(n9808) );
  NAND2_X1 U8511 ( .A1(n9228), .A2(n9835), .ZN(n9805) );
  NAND2_X1 U8512 ( .A1(n9805), .A2(n9807), .ZN(n6644) );
  INV_X1 U8513 ( .A(n9805), .ZN(n6643) );
  AOI22_X1 U8514 ( .A1(n9924), .A2(n6644), .B1(n6643), .B2(n9814), .ZN(n6646)
         );
  NAND2_X1 U8515 ( .A1(n9820), .A2(n9833), .ZN(n6645) );
  OR2_X1 U8516 ( .A1(n9900), .A2(n9776), .ZN(n9742) );
  INV_X1 U8517 ( .A(n9801), .ZN(n9767) );
  NAND2_X1 U8518 ( .A1(n9906), .A2(n9767), .ZN(n6647) );
  NAND2_X1 U8519 ( .A1(n6647), .A2(n9115), .ZN(n6648) );
  INV_X1 U8520 ( .A(n6647), .ZN(n9740) );
  AOI22_X1 U8521 ( .A1(n9900), .A2(n6648), .B1(n9740), .B2(n9776), .ZN(n6649)
         );
  OAI21_X1 U8522 ( .B1(n9728), .B2(n9749), .A(n6649), .ZN(n6650) );
  INV_X1 U8523 ( .A(n6650), .ZN(n6651) );
  OR2_X1 U8524 ( .A1(n9734), .A2(n9752), .ZN(n9705) );
  NAND2_X1 U8525 ( .A1(n9749), .A2(n9728), .ZN(n9703) );
  NAND2_X1 U8526 ( .A1(n9734), .A2(n9752), .ZN(n9706) );
  NAND2_X1 U8527 ( .A1(n9721), .A2(n9729), .ZN(n6652) );
  NAND2_X1 U8528 ( .A1(n9877), .A2(n9714), .ZN(n6655) );
  NAND2_X1 U8529 ( .A1(n9675), .A2(n9652), .ZN(n6657) );
  NOR2_X1 U8530 ( .A1(n9675), .A2(n9652), .ZN(n6656) );
  NAND2_X1 U8531 ( .A1(n9944), .A2(n6658), .ZN(n6659) );
  OR2_X1 U8532 ( .A1(n9621), .A2(n6909), .ZN(n6660) );
  NAND2_X1 U8533 ( .A1(n9644), .A2(n9627), .ZN(n9616) );
  AND2_X1 U8534 ( .A1(n6660), .A2(n9616), .ZN(n6661) );
  NAND2_X1 U8535 ( .A1(n9621), .A2(n6909), .ZN(n6662) );
  OAI21_X1 U8536 ( .B1(n6664), .B2(n9306), .A(n6976), .ZN(n8576) );
  INV_X1 U8537 ( .A(n6721), .ZN(n6667) );
  NAND2_X1 U8538 ( .A1(n6722), .A2(n6667), .ZN(n6668) );
  AND2_X1 U8539 ( .A1(n6668), .A2(n7652), .ZN(n6671) );
  INV_X1 U8540 ( .A(n6722), .ZN(n6670) );
  NAND2_X1 U8541 ( .A1(n6670), .A2(n6720), .ZN(n7653) );
  NAND2_X1 U8542 ( .A1(n6671), .A2(n7653), .ZN(n7637) );
  NAND2_X1 U8543 ( .A1(n8581), .A2(n9884), .ZN(n6672) );
  NAND2_X1 U8544 ( .A1(n6675), .A2(n6674), .ZN(P1_U3550) );
  INV_X1 U8545 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6677) );
  MUX2_X1 U8546 ( .A(n6677), .B(n6676), .S(n10115), .Z(n6681) );
  NAND2_X1 U8547 ( .A1(n8581), .A2(n9954), .ZN(n6678) );
  NAND2_X1 U8548 ( .A1(n6681), .A2(n6680), .ZN(P1_U3518) );
  INV_X1 U8549 ( .A(n6682), .ZN(n6686) );
  NAND3_X1 U8550 ( .A1(n8837), .A2(n6684), .A3(n6683), .ZN(n6685) );
  AOI21_X1 U8551 ( .B1(n6686), .B2(n6685), .A(n8856), .ZN(n6687) );
  INV_X1 U8552 ( .A(n6687), .ZN(n6704) );
  INV_X1 U8553 ( .A(n6688), .ZN(n6693) );
  NAND3_X1 U8554 ( .A1(n6689), .A2(n6691), .A3(n6690), .ZN(n6692) );
  INV_X1 U8555 ( .A(n6694), .ZN(n6695) );
  INV_X1 U8556 ( .A(n6698), .ZN(n6697) );
  OAI21_X1 U8557 ( .B1(n6697), .B2(n8742), .A(n8846), .ZN(n6699) );
  INV_X1 U8558 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10205) );
  NAND2_X1 U8559 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8705) );
  OAI21_X1 U8560 ( .B1(n8088), .B2(n10205), .A(n8705), .ZN(n6700) );
  INV_X1 U8561 ( .A(n6700), .ZN(n6701) );
  NAND4_X1 U8562 ( .A1(n6704), .A2(n6703), .A3(n6702), .A4(n6701), .ZN(
        P2_U3200) );
  OAI21_X1 U8563 ( .B1(n5032), .B2(n6705), .A(n6957), .ZN(n6709) );
  NAND2_X1 U8564 ( .A1(n9637), .A2(n9836), .ZN(n6706) );
  NOR2_X1 U8565 ( .A1(n9852), .A2(n9619), .ZN(n6711) );
  MUX2_X1 U8566 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9851), .S(n10115), .Z(n6713) );
  INV_X1 U8567 ( .A(n6713), .ZN(n6716) );
  OAI22_X1 U8568 ( .A1(n9853), .A2(n9980), .B1(n9852), .B2(n9975), .ZN(n6714)
         );
  INV_X1 U8569 ( .A(n6714), .ZN(n6715) );
  OR2_X4 U8570 ( .A1(n6720), .A2(n7029), .ZN(n6919) );
  OAI22_X1 U8571 ( .A1(n9692), .A2(n6919), .B1(n9253), .B2(n6918), .ZN(n6718)
         );
  INV_X1 U8572 ( .A(n6720), .ZN(n7636) );
  XNOR2_X1 U8573 ( .A(n6718), .B(n6921), .ZN(n6889) );
  INV_X1 U8574 ( .A(n6889), .ZN(n9152) );
  OAI22_X1 U8575 ( .A1(n9721), .A2(n6919), .B1(n9729), .B2(n6918), .ZN(n6719)
         );
  XNOR2_X1 U8576 ( .A(n6719), .B(n6921), .ZN(n9082) );
  NAND2_X1 U8577 ( .A1(n6723), .A2(n6722), .ZN(n6724) );
  OAI22_X1 U8578 ( .A1(n9721), .A2(n6918), .B1(n9729), .B2(n6888), .ZN(n6887)
         );
  NAND2_X1 U8579 ( .A1(n6725), .A2(n4284), .ZN(n6729) );
  INV_X1 U8580 ( .A(n10080), .ZN(n6726) );
  NAND2_X1 U8581 ( .A1(n6729), .A2(n6728), .ZN(n6730) );
  XNOR2_X1 U8582 ( .A(n8547), .B(n6730), .ZN(n6735) );
  INV_X1 U8583 ( .A(n6735), .ZN(n6733) );
  NOR2_X1 U8584 ( .A1(n6911), .A2(n10080), .ZN(n6731) );
  AOI21_X1 U8585 ( .B1(n8544), .B2(n6725), .A(n6731), .ZN(n6734) );
  INV_X1 U8586 ( .A(n6734), .ZN(n6732) );
  NAND2_X1 U8587 ( .A1(n6733), .A2(n6732), .ZN(n7262) );
  NAND2_X1 U8588 ( .A1(n6735), .A2(n6734), .ZN(n7261) );
  NAND2_X1 U8589 ( .A1(n6739), .A2(n4284), .ZN(n6737) );
  NAND2_X1 U8590 ( .A1(n7029), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6738) );
  AOI22_X1 U8591 ( .A1(n4284), .A2(n7651), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n7029), .ZN(n6742) );
  NAND2_X1 U8592 ( .A1(n6740), .A2(n6739), .ZN(n6741) );
  NAND2_X1 U8593 ( .A1(n6742), .A2(n6741), .ZN(n7424) );
  NAND2_X1 U8594 ( .A1(n7423), .A2(n7424), .ZN(n6743) );
  OAI21_X1 U8595 ( .B1(n6744), .B2(n6921), .A(n6743), .ZN(n7264) );
  NAND2_X1 U8596 ( .A1(n7261), .A2(n7264), .ZN(n6745) );
  NAND2_X1 U8597 ( .A1(n7262), .A2(n6745), .ZN(n7534) );
  INV_X1 U8598 ( .A(n7534), .ZN(n6752) );
  NAND2_X1 U8599 ( .A1(n6727), .A2(n9363), .ZN(n6747) );
  NAND2_X1 U8600 ( .A1(n9431), .A2(n4284), .ZN(n6746) );
  NAND2_X1 U8601 ( .A1(n6747), .A2(n6746), .ZN(n6749) );
  OAI22_X1 U8602 ( .A1(n9364), .A2(n6888), .B1(n6750), .B2(n6911), .ZN(n6754)
         );
  XNOR2_X1 U8603 ( .A(n6753), .B(n6754), .ZN(n7537) );
  INV_X1 U8604 ( .A(n7537), .ZN(n6751) );
  NAND2_X1 U8605 ( .A1(n6752), .A2(n6751), .ZN(n7535) );
  INV_X1 U8606 ( .A(n6753), .ZN(n6756) );
  INV_X1 U8607 ( .A(n6754), .ZN(n6755) );
  NAND2_X1 U8608 ( .A1(n6756), .A2(n6755), .ZN(n6757) );
  NAND2_X1 U8609 ( .A1(n9430), .A2(n4284), .ZN(n6759) );
  NAND2_X1 U8610 ( .A1(n6727), .A2(n7672), .ZN(n6758) );
  OAI22_X1 U8611 ( .A1(n7646), .A2(n6888), .B1(n10089), .B2(n6918), .ZN(n6762)
         );
  XNOR2_X1 U8612 ( .A(n6761), .B(n6762), .ZN(n7591) );
  INV_X1 U8613 ( .A(n6761), .ZN(n6763) );
  NOR2_X1 U8614 ( .A1(n6763), .A2(n6762), .ZN(n6764) );
  AOI21_X2 U8615 ( .B1(n7592), .B2(n7591), .A(n6764), .ZN(n9133) );
  NAND2_X1 U8616 ( .A1(n6727), .A2(n9134), .ZN(n6766) );
  NAND2_X1 U8617 ( .A1(n9429), .A2(n4284), .ZN(n6765) );
  NAND2_X1 U8618 ( .A1(n6766), .A2(n6765), .ZN(n6767) );
  XNOR2_X1 U8619 ( .A(n6767), .B(n8547), .ZN(n6768) );
  OAI22_X1 U8620 ( .A1(n7666), .A2(n6888), .B1(n10095), .B2(n6918), .ZN(n6769)
         );
  XNOR2_X1 U8621 ( .A(n6768), .B(n6769), .ZN(n9132) );
  INV_X1 U8622 ( .A(n6768), .ZN(n6770) );
  NAND2_X1 U8623 ( .A1(n6770), .A2(n6769), .ZN(n6771) );
  OAI22_X1 U8624 ( .A1(n7647), .A2(n6911), .B1(n10101), .B2(n6919), .ZN(n6772)
         );
  XNOR2_X1 U8625 ( .A(n6772), .B(n8547), .ZN(n7544) );
  OR2_X1 U8626 ( .A1(n7647), .A2(n6888), .ZN(n6774) );
  NAND2_X1 U8627 ( .A1(n4284), .A2(n7900), .ZN(n6773) );
  NAND2_X1 U8628 ( .A1(n6774), .A2(n6773), .ZN(n6782) );
  INV_X1 U8629 ( .A(n6782), .ZN(n7546) );
  NAND2_X1 U8630 ( .A1(n6727), .A2(n9199), .ZN(n6775) );
  OAI21_X1 U8631 ( .B1(n9200), .B2(n6918), .A(n6775), .ZN(n6776) );
  XNOR2_X1 U8632 ( .A(n6776), .B(n8547), .ZN(n7620) );
  OR2_X1 U8633 ( .A1(n9200), .A2(n6888), .ZN(n6778) );
  NAND2_X1 U8634 ( .A1(n9199), .A2(n4284), .ZN(n6777) );
  NAND2_X1 U8635 ( .A1(n6778), .A2(n6777), .ZN(n6781) );
  INV_X1 U8636 ( .A(n6781), .ZN(n7619) );
  AOI22_X1 U8637 ( .A1(n7544), .A2(n7546), .B1(n7620), .B2(n7619), .ZN(n6779)
         );
  INV_X1 U8638 ( .A(n7544), .ZN(n7618) );
  NAND2_X1 U8639 ( .A1(n7618), .A2(n6782), .ZN(n6780) );
  NAND2_X1 U8640 ( .A1(n6780), .A2(n7619), .ZN(n6785) );
  INV_X1 U8641 ( .A(n7620), .ZN(n6784) );
  AND2_X1 U8642 ( .A1(n6782), .A2(n6781), .ZN(n6783) );
  AOI22_X1 U8643 ( .A1(n6785), .A2(n6784), .B1(n6783), .B2(n7618), .ZN(n6786)
         );
  INV_X1 U8644 ( .A(n7525), .ZN(n6797) );
  NAND2_X1 U8645 ( .A1(n7911), .A2(n6727), .ZN(n6787) );
  OAI21_X1 U8646 ( .B1(n7998), .B2(n6911), .A(n6787), .ZN(n6788) );
  XNOR2_X1 U8647 ( .A(n6788), .B(n8547), .ZN(n6791) );
  OR2_X1 U8648 ( .A1(n7998), .A2(n6888), .ZN(n6790) );
  NAND2_X1 U8649 ( .A1(n7911), .A2(n8543), .ZN(n6789) );
  AND2_X1 U8650 ( .A1(n6790), .A2(n6789), .ZN(n6792) );
  NAND2_X1 U8651 ( .A1(n6791), .A2(n6792), .ZN(n7776) );
  INV_X1 U8652 ( .A(n6791), .ZN(n6794) );
  INV_X1 U8653 ( .A(n6792), .ZN(n6793) );
  NAND2_X1 U8654 ( .A1(n6794), .A2(n6793), .ZN(n6795) );
  NAND2_X1 U8655 ( .A1(n7776), .A2(n6795), .ZN(n7526) );
  INV_X1 U8656 ( .A(n7526), .ZN(n6796) );
  NAND2_X1 U8657 ( .A1(n8075), .A2(n6727), .ZN(n6799) );
  OR2_X1 U8658 ( .A1(n7530), .A2(n6918), .ZN(n6798) );
  NAND2_X1 U8659 ( .A1(n6799), .A2(n6798), .ZN(n6800) );
  XNOR2_X1 U8660 ( .A(n6800), .B(n6921), .ZN(n6811) );
  NAND2_X1 U8661 ( .A1(n8075), .A2(n8543), .ZN(n6802) );
  OR2_X1 U8662 ( .A1(n7530), .A2(n6888), .ZN(n6801) );
  NAND2_X1 U8663 ( .A1(n6802), .A2(n6801), .ZN(n7777) );
  NAND2_X1 U8664 ( .A1(n6811), .A2(n7777), .ZN(n7879) );
  NAND2_X1 U8665 ( .A1(n7875), .A2(n6727), .ZN(n6804) );
  OR2_X1 U8666 ( .A1(n7997), .A2(n6918), .ZN(n6803) );
  NAND2_X1 U8667 ( .A1(n6804), .A2(n6803), .ZN(n6805) );
  XNOR2_X1 U8668 ( .A(n6805), .B(n6921), .ZN(n6810) );
  INV_X1 U8669 ( .A(n6810), .ZN(n6807) );
  NOR2_X1 U8670 ( .A1(n7997), .A2(n6888), .ZN(n6806) );
  AOI21_X1 U8671 ( .B1(n7875), .B2(n8543), .A(n6806), .ZN(n6809) );
  OR2_X1 U8672 ( .A1(n6807), .A2(n6809), .ZN(n6808) );
  AND2_X1 U8673 ( .A1(n7879), .A2(n6808), .ZN(n6817) );
  INV_X1 U8674 ( .A(n6808), .ZN(n6816) );
  XNOR2_X1 U8675 ( .A(n6810), .B(n6809), .ZN(n7884) );
  INV_X1 U8676 ( .A(n6811), .ZN(n7878) );
  NAND2_X1 U8677 ( .A1(n7776), .A2(n7777), .ZN(n6814) );
  INV_X1 U8678 ( .A(n7776), .ZN(n6813) );
  INV_X1 U8679 ( .A(n7777), .ZN(n6812) );
  AOI22_X1 U8680 ( .A1(n7878), .A2(n6814), .B1(n6813), .B2(n6812), .ZN(n6815)
         );
  AND2_X1 U8681 ( .A1(n7884), .A2(n6815), .ZN(n7881) );
  AOI21_X2 U8682 ( .B1(n7880), .B2(n6817), .A(n5191), .ZN(n7974) );
  NAND2_X1 U8683 ( .A1(n7769), .A2(n6727), .ZN(n6819) );
  OR2_X1 U8684 ( .A1(n7888), .A2(n6918), .ZN(n6818) );
  NAND2_X1 U8685 ( .A1(n6819), .A2(n6818), .ZN(n6820) );
  XNOR2_X1 U8686 ( .A(n6820), .B(n6921), .ZN(n6829) );
  NAND2_X1 U8687 ( .A1(n7769), .A2(n8543), .ZN(n6822) );
  OR2_X1 U8688 ( .A1(n7888), .A2(n6888), .ZN(n6821) );
  NAND2_X1 U8689 ( .A1(n6822), .A2(n6821), .ZN(n7978) );
  NAND2_X1 U8690 ( .A1(n6484), .A2(n6727), .ZN(n6825) );
  OR2_X1 U8691 ( .A1(n7981), .A2(n6911), .ZN(n6824) );
  NAND2_X1 U8692 ( .A1(n6825), .A2(n6824), .ZN(n6826) );
  XNOR2_X1 U8693 ( .A(n6826), .B(n6921), .ZN(n6833) );
  NAND2_X1 U8694 ( .A1(n6484), .A2(n8543), .ZN(n6828) );
  OR2_X1 U8695 ( .A1(n7981), .A2(n6888), .ZN(n6827) );
  NAND2_X1 U8696 ( .A1(n6828), .A2(n6827), .ZN(n6834) );
  INV_X1 U8697 ( .A(n8061), .ZN(n6832) );
  INV_X1 U8698 ( .A(n6829), .ZN(n7975) );
  INV_X1 U8699 ( .A(n7978), .ZN(n6830) );
  NOR2_X1 U8700 ( .A1(n7975), .A2(n6830), .ZN(n6831) );
  INV_X1 U8701 ( .A(n6833), .ZN(n6836) );
  INV_X1 U8702 ( .A(n6834), .ZN(n6835) );
  NAND2_X1 U8703 ( .A1(n6836), .A2(n6835), .ZN(n8060) );
  NAND2_X1 U8704 ( .A1(n6837), .A2(n6727), .ZN(n6839) );
  OR2_X1 U8705 ( .A1(n9422), .A2(n6918), .ZN(n6838) );
  NAND2_X1 U8706 ( .A1(n6839), .A2(n6838), .ZN(n6840) );
  XNOR2_X1 U8707 ( .A(n6840), .B(n6921), .ZN(n6842) );
  OAI22_X1 U8708 ( .A1(n8045), .A2(n6918), .B1(n9422), .B2(n6888), .ZN(n6841)
         );
  XNOR2_X1 U8709 ( .A(n6842), .B(n6841), .ZN(n8042) );
  NAND2_X1 U8710 ( .A1(n9228), .A2(n6727), .ZN(n6844) );
  NAND2_X1 U8711 ( .A1(n9835), .A2(n4284), .ZN(n6843) );
  NAND2_X1 U8712 ( .A1(n6844), .A2(n6843), .ZN(n6845) );
  XNOR2_X1 U8713 ( .A(n6845), .B(n6921), .ZN(n6846) );
  AOI22_X1 U8714 ( .A1(n9228), .A2(n8543), .B1(n8544), .B2(n9835), .ZN(n6847)
         );
  XNOR2_X1 U8715 ( .A(n6846), .B(n6847), .ZN(n8261) );
  INV_X1 U8716 ( .A(n6846), .ZN(n6848) );
  NOR2_X1 U8717 ( .A1(n9807), .A2(n6911), .ZN(n6849) );
  AOI21_X1 U8718 ( .B1(n9924), .B2(n6727), .A(n6849), .ZN(n6850) );
  XNOR2_X1 U8719 ( .A(n6850), .B(n6921), .ZN(n6852) );
  OAI22_X1 U8720 ( .A1(n9846), .A2(n6918), .B1(n9807), .B2(n6888), .ZN(n6851)
         );
  XNOR2_X1 U8721 ( .A(n6852), .B(n6851), .ZN(n8132) );
  INV_X1 U8722 ( .A(n6851), .ZN(n6853) );
  NAND2_X1 U8723 ( .A1(n9911), .A2(n6727), .ZN(n6855) );
  NAND2_X1 U8724 ( .A1(n9815), .A2(n8543), .ZN(n6854) );
  NAND2_X1 U8725 ( .A1(n6855), .A2(n6854), .ZN(n6856) );
  XNOR2_X1 U8726 ( .A(n6856), .B(n8547), .ZN(n9104) );
  NOR2_X1 U8727 ( .A1(n9180), .A2(n6888), .ZN(n6857) );
  AOI21_X1 U8728 ( .B1(n9911), .B2(n8543), .A(n6857), .ZN(n9103) );
  NAND2_X1 U8729 ( .A1(n9820), .A2(n6727), .ZN(n6859) );
  NAND2_X1 U8730 ( .A1(n9833), .A2(n4284), .ZN(n6858) );
  NAND2_X1 U8731 ( .A1(n6859), .A2(n6858), .ZN(n6860) );
  XNOR2_X1 U8732 ( .A(n6860), .B(n6921), .ZN(n9102) );
  NAND2_X1 U8733 ( .A1(n9820), .A2(n8543), .ZN(n6862) );
  NAND2_X1 U8734 ( .A1(n8544), .A2(n9833), .ZN(n6861) );
  NAND2_X1 U8735 ( .A1(n6862), .A2(n6861), .ZN(n9100) );
  INV_X1 U8736 ( .A(n9103), .ZN(n6865) );
  AOI21_X1 U8737 ( .B1(n9102), .B2(n9100), .A(n6865), .ZN(n6867) );
  NAND3_X1 U8738 ( .A1(n9102), .A2(n9100), .A3(n6865), .ZN(n6866) );
  OAI22_X1 U8739 ( .A1(n9783), .A2(n6919), .B1(n9801), .B2(n6918), .ZN(n6871)
         );
  XNOR2_X1 U8740 ( .A(n6871), .B(n6921), .ZN(n6872) );
  OAI22_X1 U8741 ( .A1(n9783), .A2(n6918), .B1(n9801), .B2(n6888), .ZN(n6873)
         );
  XNOR2_X1 U8742 ( .A(n6872), .B(n6873), .ZN(n9112) );
  OAI22_X1 U8743 ( .A1(n9763), .A2(n6919), .B1(n9115), .B2(n6918), .ZN(n6874)
         );
  XOR2_X1 U8744 ( .A(n6921), .B(n6874), .Z(n6875) );
  OAI22_X1 U8745 ( .A1(n9763), .A2(n6918), .B1(n9115), .B2(n6888), .ZN(n9162)
         );
  OAI22_X1 U8746 ( .A1(n9749), .A2(n6911), .B1(n9728), .B2(n6888), .ZN(n6877)
         );
  OAI22_X1 U8747 ( .A1(n9749), .A2(n6919), .B1(n9728), .B2(n6918), .ZN(n6876)
         );
  XNOR2_X1 U8748 ( .A(n6876), .B(n6921), .ZN(n6878) );
  XOR2_X1 U8749 ( .A(n6877), .B(n6878), .Z(n9075) );
  NAND2_X1 U8750 ( .A1(n9734), .A2(n6727), .ZN(n6881) );
  NAND2_X1 U8751 ( .A1(n9752), .A2(n8543), .ZN(n6880) );
  NAND2_X1 U8752 ( .A1(n6881), .A2(n6880), .ZN(n6882) );
  XNOR2_X1 U8753 ( .A(n6882), .B(n6921), .ZN(n6886) );
  NAND2_X1 U8754 ( .A1(n9734), .A2(n4284), .ZN(n6884) );
  NAND2_X1 U8755 ( .A1(n9752), .A2(n8544), .ZN(n6883) );
  NAND2_X1 U8756 ( .A1(n6884), .A2(n6883), .ZN(n6885) );
  NOR2_X1 U8757 ( .A1(n6886), .A2(n6885), .ZN(n9140) );
  NAND2_X1 U8758 ( .A1(n6886), .A2(n6885), .ZN(n9141) );
  INV_X1 U8759 ( .A(n9154), .ZN(n6891) );
  OAI22_X1 U8760 ( .A1(n9692), .A2(n6911), .B1(n9253), .B2(n6888), .ZN(n9151)
         );
  OAI22_X1 U8761 ( .A1(n9675), .A2(n6919), .B1(n9652), .B2(n6911), .ZN(n6892)
         );
  XOR2_X1 U8762 ( .A(n6921), .B(n6892), .Z(n6894) );
  AOI22_X1 U8763 ( .A1(n9947), .A2(n8543), .B1(n8544), .B2(n9688), .ZN(n6893)
         );
  NAND2_X1 U8764 ( .A1(n6894), .A2(n6893), .ZN(n6895) );
  OAI21_X1 U8765 ( .B1(n6894), .B2(n6893), .A(n6895), .ZN(n9067) );
  INV_X1 U8766 ( .A(n6895), .ZN(n9122) );
  NAND2_X1 U8767 ( .A1(n9660), .A2(n6727), .ZN(n6897) );
  NAND2_X1 U8768 ( .A1(n9673), .A2(n8543), .ZN(n6896) );
  NAND2_X1 U8769 ( .A1(n6897), .A2(n6896), .ZN(n6898) );
  XNOR2_X1 U8770 ( .A(n6898), .B(n8547), .ZN(n6900) );
  AND2_X1 U8771 ( .A1(n9673), .A2(n8544), .ZN(n6899) );
  AOI21_X1 U8772 ( .B1(n9660), .B2(n4284), .A(n6899), .ZN(n6901) );
  NAND2_X1 U8773 ( .A1(n6900), .A2(n6901), .ZN(n6905) );
  INV_X1 U8774 ( .A(n6900), .ZN(n6903) );
  INV_X1 U8775 ( .A(n6901), .ZN(n6902) );
  NAND2_X1 U8776 ( .A1(n6903), .A2(n6902), .ZN(n6904) );
  AND2_X1 U8777 ( .A1(n6905), .A2(n6904), .ZN(n9121) );
  OAI21_X2 U8778 ( .B1(n9123), .B2(n9122), .A(n9121), .ZN(n9120) );
  NAND2_X1 U8779 ( .A1(n9644), .A2(n6727), .ZN(n6907) );
  NAND2_X1 U8780 ( .A1(n9627), .A2(n8543), .ZN(n6906) );
  NAND2_X1 U8781 ( .A1(n6907), .A2(n6906), .ZN(n6908) );
  XNOR2_X1 U8782 ( .A(n6908), .B(n6921), .ZN(n6914) );
  AOI22_X1 U8783 ( .A1(n9644), .A2(n8543), .B1(n8544), .B2(n9627), .ZN(n6915)
         );
  XNOR2_X1 U8784 ( .A(n6914), .B(n6915), .ZN(n9092) );
  OAI22_X1 U8785 ( .A1(n9621), .A2(n6919), .B1(n6909), .B2(n6918), .ZN(n6910)
         );
  XNOR2_X1 U8786 ( .A(n6910), .B(n8547), .ZN(n6924) );
  OR2_X1 U8787 ( .A1(n9621), .A2(n6911), .ZN(n6913) );
  NAND2_X1 U8788 ( .A1(n9637), .A2(n8544), .ZN(n6912) );
  NAND2_X1 U8789 ( .A1(n6913), .A2(n6912), .ZN(n6925) );
  XNOR2_X1 U8790 ( .A(n6924), .B(n6925), .ZN(n8271) );
  INV_X1 U8791 ( .A(n6914), .ZN(n6916) );
  NAND2_X1 U8792 ( .A1(n6916), .A2(n6915), .ZN(n8272) );
  OAI22_X1 U8793 ( .A1(n9852), .A2(n6919), .B1(n10374), .B2(n6918), .ZN(n6920)
         );
  XOR2_X1 U8794 ( .A(n6921), .B(n6920), .Z(n6923) );
  AOI22_X1 U8795 ( .A1(n9609), .A2(n8543), .B1(n8544), .B2(n9628), .ZN(n6922)
         );
  NAND2_X1 U8796 ( .A1(n6923), .A2(n6922), .ZN(n8559) );
  OAI21_X1 U8797 ( .B1(n6923), .B2(n6922), .A(n8559), .ZN(n6929) );
  INV_X1 U8798 ( .A(n6924), .ZN(n6926) );
  AND2_X2 U8799 ( .A1(n8273), .A2(n6927), .ZN(n8565) );
  INV_X1 U8800 ( .A(n6928), .ZN(n6931) );
  INV_X1 U8801 ( .A(n6929), .ZN(n6930) );
  AOI21_X1 U8802 ( .B1(n8273), .B2(n6931), .A(n6930), .ZN(n6935) );
  AND2_X1 U8803 ( .A1(n6717), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6932) );
  AND3_X1 U8804 ( .A1(n6934), .A2(n9986), .A3(n6933), .ZN(n6940) );
  AND2_X1 U8805 ( .A1(n10107), .A2(n9344), .ZN(n6938) );
  OAI21_X1 U8806 ( .B1(n8565), .B2(n6935), .A(n9175), .ZN(n6954) );
  INV_X1 U8807 ( .A(n6936), .ZN(n6950) );
  NOR2_X1 U8808 ( .A1(n6950), .A2(n7653), .ZN(n6946) );
  INV_X1 U8809 ( .A(n6946), .ZN(n7266) );
  INV_X1 U8810 ( .A(n7653), .ZN(n6937) );
  AND2_X1 U8811 ( .A1(n6937), .A2(n9985), .ZN(n9357) );
  INV_X1 U8812 ( .A(n6938), .ZN(n6939) );
  OR2_X1 U8813 ( .A1(n9414), .A2(P1_U3086), .ZN(n7785) );
  NAND2_X1 U8814 ( .A1(n6939), .A2(n7785), .ZN(n6942) );
  INV_X1 U8815 ( .A(n6940), .ZN(n6941) );
  OAI21_X1 U8816 ( .B1(n9357), .B2(n6942), .A(n6941), .ZN(n6945) );
  INV_X1 U8817 ( .A(n6943), .ZN(n6944) );
  NAND2_X1 U8818 ( .A1(n6945), .A2(n6944), .ZN(n7265) );
  OAI22_X1 U8819 ( .A1(n9607), .A2(n9164), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10278), .ZN(n6948) );
  NOR2_X1 U8820 ( .A1(n8550), .A2(n9181), .ZN(n6947) );
  AOI211_X1 U8821 ( .C1(n9177), .C2(n9637), .A(n6948), .B(n6947), .ZN(n6953)
         );
  NAND2_X1 U8822 ( .A1(n9985), .A2(n9414), .ZN(n6949) );
  NAND2_X1 U8823 ( .A1(n6950), .A2(n6949), .ZN(n6951) );
  NAND2_X1 U8824 ( .A1(n9609), .A2(n9168), .ZN(n6952) );
  NAND3_X1 U8825 ( .A1(n6954), .A2(n6953), .A3(n6952), .ZN(P1_U3214) );
  NAND2_X1 U8826 ( .A1(n9269), .A2(n9270), .ZN(n9340) );
  XNOR2_X1 U8827 ( .A(n6958), .B(n9307), .ZN(n6968) );
  NAND2_X1 U8828 ( .A1(n6959), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6964) );
  NAND2_X1 U8829 ( .A1(n6960), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6963) );
  NAND2_X1 U8830 ( .A1(n6961), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6962) );
  INV_X1 U8831 ( .A(n9269), .ZN(n6969) );
  NOR2_X1 U8832 ( .A1(n6969), .A2(n10107), .ZN(n6973) );
  AOI21_X1 U8833 ( .B1(n9269), .B2(n6970), .A(n9864), .ZN(n6972) );
  NOR3_X1 U8834 ( .A1(n8539), .A2(n6973), .A3(n8538), .ZN(n6980) );
  MUX2_X1 U8835 ( .A(n6974), .B(n6980), .S(n10123), .Z(n6979) );
  XNOR2_X1 U8836 ( .A(n6977), .B(n9307), .ZN(n8542) );
  NAND2_X1 U8837 ( .A1(n6979), .A2(n6978), .ZN(P1_U3551) );
  INV_X1 U8838 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6981) );
  MUX2_X1 U8839 ( .A(n6981), .B(n6980), .S(n10115), .Z(n6983) );
  NAND2_X1 U8840 ( .A1(n6983), .A2(n6982), .ZN(P1_U3519) );
  NOR2_X1 U8841 ( .A1(n6717), .A2(P1_U3086), .ZN(n6984) );
  NAND2_X1 U8842 ( .A1(n6990), .A2(P1_U3086), .ZN(n9993) );
  INV_X1 U8843 ( .A(n9993), .ZN(n7346) );
  INV_X1 U8844 ( .A(n7346), .ZN(n10002) );
  NOR2_X1 U8845 ( .A1(n6990), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9987) );
  INV_X2 U8846 ( .A(n9987), .ZN(n8589) );
  INV_X1 U8847 ( .A(n9482), .ZN(n9477) );
  OAI222_X1 U8848 ( .A1(n10002), .A2(n6985), .B1(n8589), .B2(n6993), .C1(
        P1_U3086), .C2(n9477), .ZN(P1_U3350) );
  OAI222_X1 U8849 ( .A1(n6986), .A2(n9993), .B1(P1_U3086), .B2(n10055), .C1(
        n8589), .C2(n6996), .ZN(P1_U3351) );
  OAI222_X1 U8850 ( .A1(n10002), .A2(n6987), .B1(n8589), .B2(n6991), .C1(
        P1_U3086), .C2(n9467), .ZN(P1_U3352) );
  OAI222_X1 U8851 ( .A1(P1_U3086), .A2(n9446), .B1(n8589), .B2(n7014), .C1(
        n6988), .C2(n10002), .ZN(P1_U3353) );
  OAI222_X1 U8852 ( .A1(n7064), .A2(P1_U3086), .B1(n8589), .B2(n4287), .C1(
        n6989), .C2(n10002), .ZN(P1_U3354) );
  NOR2_X1 U8853 ( .A1(n6990), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9058) );
  OAI222_X1 U8854 ( .A1(n9062), .A2(n6992), .B1(n9063), .B2(n6991), .C1(
        P2_U3151), .C2(n4286), .ZN(P2_U3292) );
  OAI222_X1 U8855 ( .A1(n9062), .A2(n6994), .B1(n9063), .B2(n6993), .C1(
        P2_U3151), .C2(n7154), .ZN(P2_U3290) );
  OAI222_X1 U8856 ( .A1(n9062), .A2(n6997), .B1(n9063), .B2(n6996), .C1(
        P2_U3151), .C2(n6995), .ZN(P2_U3291) );
  INV_X1 U8857 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6999) );
  INV_X1 U8858 ( .A(n6998), .ZN(n7000) );
  INV_X1 U8859 ( .A(n9503), .ZN(n7072) );
  OAI222_X1 U8860 ( .A1(n10002), .A2(n6999), .B1(n8589), .B2(n7000), .C1(
        P1_U3086), .C2(n7072), .ZN(P1_U3349) );
  INV_X1 U8861 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7001) );
  OAI222_X1 U8862 ( .A1(n9062), .A2(n7001), .B1(n9063), .B2(n7000), .C1(
        P2_U3151), .C2(n7235), .ZN(P2_U3289) );
  INV_X1 U8863 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7003) );
  INV_X1 U8864 ( .A(n7002), .ZN(n7012) );
  INV_X1 U8865 ( .A(n7121), .ZN(n7118) );
  OAI222_X1 U8866 ( .A1(n10002), .A2(n7003), .B1(n8589), .B2(n7012), .C1(
        P1_U3086), .C2(n7118), .ZN(P1_U3348) );
  INV_X1 U8867 ( .A(n7004), .ZN(n7017) );
  INV_X1 U8868 ( .A(n7137), .ZN(n7077) );
  OAI222_X1 U8869 ( .A1(n10002), .A2(n10359), .B1(n8589), .B2(n7017), .C1(
        P1_U3086), .C2(n7077), .ZN(P1_U3347) );
  INV_X1 U8870 ( .A(n7008), .ZN(n7009) );
  AOI22_X1 U8871 ( .A1(n7023), .A2(n10237), .B1(n7009), .B2(n7010), .ZN(
        P2_U3377) );
  AOI22_X1 U8872 ( .A1(n7023), .A2(n7011), .B1(n5179), .B2(n7010), .ZN(
        P2_U3376) );
  OAI222_X1 U8873 ( .A1(n9062), .A2(n4699), .B1(n9063), .B2(n7012), .C1(
        P2_U3151), .C2(n7328), .ZN(P2_U3288) );
  OAI222_X1 U8874 ( .A1(n7015), .A2(P2_U3151), .B1(n9063), .B2(n7014), .C1(
        n7013), .C2(n9062), .ZN(P2_U3293) );
  INV_X1 U8875 ( .A(n7016), .ZN(n7370) );
  OAI222_X1 U8876 ( .A1(P2_U3151), .A2(n7370), .B1(n9063), .B2(n7017), .C1(
        n9062), .C2(n5227), .ZN(P2_U3287) );
  AND2_X1 U8877 ( .A1(n7023), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8878 ( .A1(n7023), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8879 ( .A1(n7023), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8880 ( .A1(n7023), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8881 ( .A1(n7023), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8882 ( .A1(n7023), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8883 ( .A1(n7023), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8884 ( .A1(n7023), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8885 ( .A1(n7023), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8886 ( .A1(n7023), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8887 ( .A1(n7023), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8888 ( .A1(n7023), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8889 ( .A1(n7023), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8890 ( .A1(n7023), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8891 ( .A1(n7023), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8892 ( .A1(n7023), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8893 ( .A1(n7023), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8894 ( .A1(n7023), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8895 ( .A1(n7023), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8896 ( .A1(n7023), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8897 ( .A1(n7023), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8898 ( .A1(n7023), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8899 ( .A1(n7023), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U8900 ( .A(n7018), .ZN(n7021) );
  AOI22_X1 U8901 ( .A1(n7092), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n7346), .ZN(n7019) );
  OAI21_X1 U8902 ( .B1(n7021), .B2(n8589), .A(n7019), .ZN(P1_U3346) );
  OAI222_X1 U8903 ( .A1(n9062), .A2(n7022), .B1(n9063), .B2(n7021), .C1(
        P2_U3151), .C2(n7020), .ZN(P2_U3286) );
  INV_X1 U8904 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10247) );
  NOR2_X1 U8905 ( .A1(n7024), .A2(n10247), .ZN(P2_U3239) );
  INV_X1 U8906 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10338) );
  NOR2_X1 U8907 ( .A1(n7024), .A2(n10338), .ZN(P2_U3256) );
  INV_X1 U8908 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10327) );
  NOR2_X1 U8909 ( .A1(n7024), .A2(n10327), .ZN(P2_U3252) );
  INV_X1 U8910 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10347) );
  NOR2_X1 U8911 ( .A1(n7024), .A2(n10347), .ZN(P2_U3262) );
  INV_X1 U8912 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10263) );
  NOR2_X1 U8913 ( .A1(n7024), .A2(n10263), .ZN(P2_U3260) );
  INV_X1 U8914 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n10250) );
  NOR2_X1 U8915 ( .A1(n7024), .A2(n10250), .ZN(P2_U3257) );
  INV_X1 U8916 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10284) );
  NOR2_X1 U8917 ( .A1(n7024), .A2(n10284), .ZN(P2_U3258) );
  INV_X1 U8918 ( .A(n7025), .ZN(n7028) );
  AOI22_X1 U8919 ( .A1(n7210), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n7346), .ZN(n7026) );
  OAI21_X1 U8920 ( .B1(n7028), .B2(n8589), .A(n7026), .ZN(P1_U3345) );
  OAI222_X1 U8921 ( .A1(P2_U3151), .A2(n7557), .B1(n9063), .B2(n7028), .C1(
        n7027), .C2(n9062), .ZN(P2_U3285) );
  NAND2_X1 U8922 ( .A1(n8128), .A2(n7029), .ZN(n7030) );
  NAND2_X1 U8923 ( .A1(n7030), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7034) );
  INV_X1 U8924 ( .A(n7034), .ZN(n7033) );
  NAND2_X1 U8925 ( .A1(n7031), .A2(n8128), .ZN(n7032) );
  NAND2_X1 U8926 ( .A1(n7032), .A2(n5372), .ZN(n7035) );
  INV_X1 U8927 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7040) );
  INV_X1 U8928 ( .A(n9588), .ZN(n7038) );
  INV_X1 U8929 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7661) );
  AOI21_X1 U8930 ( .B1(n9452), .B2(n7661), .A(n8531), .ZN(n9458) );
  OAI21_X1 U8931 ( .B1(n9452), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9458), .ZN(
        n7036) );
  XNOR2_X1 U8932 ( .A(n7036), .B(P1_IR_REG_0__SCAN_IN), .ZN(n7037) );
  AOI22_X1 U8933 ( .A1(n7038), .A2(n7037), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n7039) );
  OAI21_X1 U8934 ( .B1(n9596), .B2(n7040), .A(n7039), .ZN(P1_U3243) );
  NAND2_X1 U8935 ( .A1(n8158), .A2(P2_U3893), .ZN(n7041) );
  OAI21_X1 U8936 ( .B1(P2_U3893), .B2(n5260), .A(n7041), .ZN(P2_U3508) );
  INV_X1 U8937 ( .A(n7042), .ZN(n7045) );
  OAI222_X1 U8938 ( .A1(n10002), .A2(n7043), .B1(n8589), .B2(n7045), .C1(
        P1_U3086), .C2(n7192), .ZN(P1_U3344) );
  OAI222_X1 U8939 ( .A1(n9062), .A2(n7046), .B1(n9063), .B2(n7045), .C1(
        P2_U3151), .C2(n7044), .ZN(P2_U3284) );
  INV_X1 U8940 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7047) );
  MUX2_X1 U8941 ( .A(n7047), .B(P1_REG2_REG_2__SCAN_IN), .S(n9446), .Z(n7050)
         );
  INV_X1 U8942 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n7048) );
  AND2_X1 U8943 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9453) );
  NAND2_X1 U8944 ( .A1(n9434), .A2(n9453), .ZN(n9433) );
  INV_X1 U8945 ( .A(n7064), .ZN(n9438) );
  NAND2_X1 U8946 ( .A1(n9438), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7049) );
  NAND2_X1 U8947 ( .A1(n9433), .A2(n7049), .ZN(n9445) );
  INV_X1 U8948 ( .A(n9446), .ZN(n9459) );
  NAND2_X1 U8949 ( .A1(n9459), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9468) );
  NAND2_X1 U8950 ( .A1(n9469), .A2(n9468), .ZN(n7052) );
  INV_X1 U8951 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7668) );
  MUX2_X1 U8952 ( .A(n7668), .B(P1_REG2_REG_3__SCAN_IN), .S(n9467), .Z(n7051)
         );
  NAND2_X1 U8953 ( .A1(n7052), .A2(n7051), .ZN(n10049) );
  INV_X1 U8954 ( .A(n9467), .ZN(n9466) );
  NAND2_X1 U8955 ( .A1(n9466), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n10048) );
  INV_X1 U8956 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7053) );
  MUX2_X1 U8957 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7053), .S(n10055), .Z(n10047) );
  NOR2_X1 U8958 ( .A1(n10055), .A2(n7053), .ZN(n9481) );
  INV_X1 U8959 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7054) );
  MUX2_X1 U8960 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7054), .S(n9482), .Z(n7055)
         );
  NAND2_X1 U8961 ( .A1(n9482), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9498) );
  INV_X1 U8962 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7828) );
  MUX2_X1 U8963 ( .A(n7828), .B(P1_REG2_REG_6__SCAN_IN), .S(n9503), .Z(n9497)
         );
  NOR2_X1 U8964 ( .A1(n7072), .A2(n7828), .ZN(n7120) );
  INV_X1 U8965 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7056) );
  MUX2_X1 U8966 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7056), .S(n7121), .Z(n7057)
         );
  NAND2_X1 U8967 ( .A1(n7121), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7131) );
  INV_X1 U8968 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7058) );
  MUX2_X1 U8969 ( .A(n7058), .B(P1_REG2_REG_8__SCAN_IN), .S(n7137), .Z(n7130)
         );
  AOI21_X1 U8970 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n7137), .A(n7134), .ZN(
        n7088) );
  INV_X1 U8971 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7059) );
  MUX2_X1 U8972 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n7059), .S(n7092), .Z(n7087)
         );
  NOR2_X1 U8973 ( .A1(n7092), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7203) );
  INV_X1 U8974 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7060) );
  MUX2_X1 U8975 ( .A(n7060), .B(P1_REG2_REG_10__SCAN_IN), .S(n7210), .Z(n7207)
         );
  AND2_X1 U8976 ( .A1(n7210), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7061) );
  INV_X1 U8977 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7193) );
  XNOR2_X1 U8978 ( .A(n7192), .B(n7193), .ZN(n7194) );
  XNOR2_X1 U8979 ( .A(n7195), .B(n7194), .ZN(n7084) );
  NOR2_X1 U8980 ( .A1(n9999), .A2(n8531), .ZN(n9356) );
  INV_X1 U8981 ( .A(n9356), .ZN(n7062) );
  NOR2_X2 U8982 ( .A1(n9588), .A2(n7062), .ZN(n10052) );
  INV_X1 U8983 ( .A(n10052), .ZN(n9556) );
  INV_X1 U8984 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7187) );
  XNOR2_X1 U8985 ( .A(n7192), .B(n7187), .ZN(n7188) );
  XNOR2_X1 U8986 ( .A(n9446), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9443) );
  INV_X1 U8987 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7063) );
  MUX2_X1 U8988 ( .A(n7063), .B(P1_REG1_REG_1__SCAN_IN), .S(n7064), .Z(n9436)
         );
  AND2_X1 U8989 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9437) );
  NAND2_X1 U8990 ( .A1(n9436), .A2(n9437), .ZN(n9435) );
  OR2_X1 U8991 ( .A1(n7064), .A2(n7063), .ZN(n7065) );
  NAND2_X1 U8992 ( .A1(n9435), .A2(n7065), .ZN(n9444) );
  NAND2_X1 U8993 ( .A1(n9443), .A2(n9444), .ZN(n7067) );
  NAND2_X1 U8994 ( .A1(n9459), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7066) );
  NAND2_X1 U8995 ( .A1(n7067), .A2(n7066), .ZN(n9472) );
  INV_X1 U8996 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7068) );
  MUX2_X1 U8997 ( .A(n7068), .B(P1_REG1_REG_3__SCAN_IN), .S(n9467), .Z(n9473)
         );
  NAND2_X1 U8998 ( .A1(n9466), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10057) );
  NAND2_X1 U8999 ( .A1(n10058), .A2(n10057), .ZN(n7071) );
  INV_X1 U9000 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7069) );
  MUX2_X1 U9001 ( .A(n7069), .B(P1_REG1_REG_4__SCAN_IN), .S(n10055), .Z(n7070)
         );
  NAND2_X1 U9002 ( .A1(n7071), .A2(n7070), .ZN(n10060) );
  INV_X1 U9003 ( .A(n10055), .ZN(n10053) );
  NAND2_X1 U9004 ( .A1(n10053), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9488) );
  INV_X1 U9005 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10118) );
  MUX2_X1 U9006 ( .A(n10118), .B(P1_REG1_REG_5__SCAN_IN), .S(n9482), .Z(n9487)
         );
  AOI21_X1 U9007 ( .B1(n10060), .B2(n9488), .A(n9487), .ZN(n9486) );
  NOR2_X1 U9008 ( .A1(n9477), .A2(n10118), .ZN(n9502) );
  NAND2_X1 U9009 ( .A1(n9503), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7074) );
  INV_X1 U9010 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10121) );
  NAND2_X1 U9011 ( .A1(n7072), .A2(n10121), .ZN(n7073) );
  NAND2_X1 U9012 ( .A1(n9508), .A2(n7074), .ZN(n7117) );
  INV_X1 U9013 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7075) );
  XNOR2_X1 U9014 ( .A(n7121), .B(n7075), .ZN(n7116) );
  XNOR2_X1 U9015 ( .A(n7137), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n7128) );
  INV_X1 U9016 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7076) );
  OAI22_X1 U9017 ( .A1(n7129), .A2(n7128), .B1(n7077), .B2(n7076), .ZN(n7085)
         );
  XNOR2_X1 U9018 ( .A(n7092), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n7086) );
  NOR2_X1 U9019 ( .A1(n7085), .A2(n7086), .ZN(n7214) );
  NOR2_X1 U9020 ( .A1(n7092), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7213) );
  XNOR2_X1 U9021 ( .A(n7210), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n7212) );
  NOR3_X1 U9022 ( .A1(n7214), .A2(n7213), .A3(n7212), .ZN(n7211) );
  XOR2_X1 U9023 ( .A(n7188), .B(n7189), .Z(n7078) );
  NOR2_X2 U9024 ( .A1(n9588), .A2(n9452), .ZN(n10061) );
  NAND2_X1 U9025 ( .A1(n7078), .A2(n10061), .ZN(n7083) );
  NOR2_X2 U9026 ( .A1(n9588), .A2(n9455), .ZN(n10054) );
  NOR2_X1 U9027 ( .A1(n7079), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8068) );
  INV_X1 U9028 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10286) );
  NOR2_X1 U9029 ( .A1(n9596), .A2(n10286), .ZN(n7080) );
  AOI211_X1 U9030 ( .C1(n10054), .C2(n7081), .A(n8068), .B(n7080), .ZN(n7082)
         );
  OAI211_X1 U9031 ( .C1(n7084), .C2(n9556), .A(n7083), .B(n7082), .ZN(P1_U3254) );
  AOI21_X1 U9032 ( .B1(n7086), .B2(n7085), .A(n7214), .ZN(n7095) );
  NOR2_X1 U9033 ( .A1(n7088), .A2(n7087), .ZN(n7089) );
  OAI21_X1 U9034 ( .B1(n7089), .B2(n7204), .A(n10052), .ZN(n7094) );
  INV_X1 U9035 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7090) );
  NAND2_X1 U9036 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7886) );
  OAI21_X1 U9037 ( .B1(n9596), .B2(n7090), .A(n7886), .ZN(n7091) );
  AOI21_X1 U9038 ( .B1(n7092), .B2(n10054), .A(n7091), .ZN(n7093) );
  OAI211_X1 U9039 ( .C1(n7095), .C2(n9561), .A(n7094), .B(n7093), .ZN(P1_U3252) );
  INV_X1 U9040 ( .A(n7096), .ZN(n7097) );
  AOI21_X1 U9041 ( .B1(n7099), .B2(n7098), .A(n7097), .ZN(n7110) );
  OAI21_X1 U9042 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n7101), .A(n7100), .ZN(
        n7102) );
  NAND2_X1 U9043 ( .A1(n8825), .A2(n7102), .ZN(n7103) );
  NAND2_X1 U9044 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3151), .ZN(n7222) );
  NAND2_X1 U9045 ( .A1(n7103), .A2(n7222), .ZN(n7108) );
  INV_X1 U9046 ( .A(n7171), .ZN(n7104) );
  AOI21_X1 U9047 ( .B1(n7482), .B2(n7105), .A(n7104), .ZN(n7106) );
  OAI22_X1 U9048 ( .A1(n7106), .A2(n8835), .B1(n8846), .B2(n4286), .ZN(n7107)
         );
  AOI211_X1 U9049 ( .C1(n8848), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n7108), .B(
        n7107), .ZN(n7109) );
  OAI21_X1 U9050 ( .B1(n7110), .B2(n8850), .A(n7109), .ZN(P2_U3185) );
  INV_X1 U9051 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7112) );
  INV_X1 U9052 ( .A(n7111), .ZN(n7115) );
  INV_X1 U9053 ( .A(n7280), .ZN(n7286) );
  OAI222_X1 U9054 ( .A1(n10002), .A2(n7112), .B1(n8589), .B2(n7115), .C1(n7286), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U9055 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7114) );
  OAI222_X1 U9056 ( .A1(P2_U3151), .A2(n6314), .B1(n9063), .B2(n7115), .C1(
        n7114), .C2(n9062), .ZN(P2_U3283) );
  XNOR2_X1 U9057 ( .A(n7117), .B(n7116), .ZN(n7127) );
  INV_X1 U9058 ( .A(n9596), .ZN(n10063) );
  AND2_X1 U9059 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7527) );
  INV_X1 U9060 ( .A(n10054), .ZN(n9580) );
  NOR2_X1 U9061 ( .A1(n9580), .A2(n7118), .ZN(n7119) );
  AOI211_X1 U9062 ( .C1(n10063), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n7527), .B(
        n7119), .ZN(n7126) );
  INV_X1 U9063 ( .A(n7120), .ZN(n7123) );
  MUX2_X1 U9064 ( .A(n7056), .B(P1_REG2_REG_7__SCAN_IN), .S(n7121), .Z(n7122)
         );
  NAND2_X1 U9065 ( .A1(n7123), .A2(n7122), .ZN(n7124) );
  OAI211_X1 U9066 ( .C1(n9496), .C2(n7124), .A(n10052), .B(n7132), .ZN(n7125)
         );
  OAI211_X1 U9067 ( .C1(n7127), .C2(n9561), .A(n7126), .B(n7125), .ZN(P1_U3250) );
  XNOR2_X1 U9068 ( .A(n7129), .B(n7128), .ZN(n7139) );
  NAND2_X1 U9069 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7779) );
  OAI21_X1 U9070 ( .B1(n9596), .B2(n10294), .A(n7779), .ZN(n7136) );
  AND3_X1 U9071 ( .A1(n7132), .A2(n7131), .A3(n7130), .ZN(n7133) );
  NOR3_X1 U9072 ( .A1(n9556), .A2(n7134), .A3(n7133), .ZN(n7135) );
  AOI211_X1 U9073 ( .C1(n10054), .C2(n7137), .A(n7136), .B(n7135), .ZN(n7138)
         );
  OAI21_X1 U9074 ( .B1(n7139), .B2(n9561), .A(n7138), .ZN(P1_U3251) );
  INV_X1 U9075 ( .A(n7140), .ZN(n7141) );
  AOI21_X1 U9076 ( .B1(n7313), .B2(n7142), .A(n7141), .ZN(n7144) );
  OAI22_X1 U9077 ( .A1(n7144), .A2(n8835), .B1(n8846), .B2(n7143), .ZN(n7149)
         );
  AOI21_X1 U9078 ( .B1(n10189), .B2(n7146), .A(n7145), .ZN(n7147) );
  OAI22_X1 U9079 ( .A1(n8856), .A2(n7147), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5741), .ZN(n7148) );
  AOI211_X1 U9080 ( .C1(n8848), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n7149), .B(
        n7148), .ZN(n7153) );
  INV_X1 U9081 ( .A(n8850), .ZN(n8766) );
  OAI211_X1 U9082 ( .C1(n7151), .C2(n7250), .A(n7150), .B(n8766), .ZN(n7152)
         );
  NAND2_X1 U9083 ( .A1(n7153), .A2(n7152), .ZN(P2_U3183) );
  NAND2_X1 U9084 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3151), .ZN(n7472) );
  OAI21_X1 U9085 ( .B1(n8846), .B2(n7154), .A(n7472), .ZN(n7162) );
  AOI21_X1 U9086 ( .B1(n7444), .B2(n7155), .A(n4310), .ZN(n7160) );
  OAI21_X1 U9087 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n7157), .A(n7156), .ZN(
        n7158) );
  NAND2_X1 U9088 ( .A1(n7158), .A2(n8825), .ZN(n7159) );
  OAI21_X1 U9089 ( .B1(n7160), .B2(n8835), .A(n7159), .ZN(n7161) );
  AOI211_X1 U9090 ( .C1(n8848), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n7162), .B(
        n7161), .ZN(n7167) );
  OAI211_X1 U9091 ( .C1(n7165), .C2(n7164), .A(n7163), .B(n8766), .ZN(n7166)
         );
  NAND2_X1 U9092 ( .A1(n7167), .A2(n7166), .ZN(P2_U3187) );
  INV_X1 U9093 ( .A(n7168), .ZN(n7170) );
  NAND3_X1 U9094 ( .A1(n7171), .A2(n7170), .A3(n7169), .ZN(n7172) );
  AOI21_X1 U9095 ( .B1(n7173), .B2(n7172), .A(n8835), .ZN(n7180) );
  INV_X1 U9096 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7178) );
  AND3_X1 U9097 ( .A1(n7100), .A2(n7174), .A3(n4290), .ZN(n7175) );
  OAI21_X1 U9098 ( .B1(n7176), .B2(n7175), .A(n8825), .ZN(n7177) );
  NAND2_X1 U9099 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7351) );
  OAI211_X1 U9100 ( .C1(n7178), .C2(n8088), .A(n7177), .B(n7351), .ZN(n7179)
         );
  AOI211_X1 U9101 ( .C1(n8764), .C2(n7181), .A(n7180), .B(n7179), .ZN(n7186)
         );
  OAI211_X1 U9102 ( .C1(n7184), .C2(n7183), .A(n7182), .B(n8766), .ZN(n7185)
         );
  NAND2_X1 U9103 ( .A1(n7186), .A2(n7185), .ZN(P2_U3186) );
  XNOR2_X1 U9104 ( .A(n7280), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n7191) );
  NOR2_X1 U9105 ( .A1(n7190), .A2(n7191), .ZN(n9521) );
  AOI21_X1 U9106 ( .B1(n7191), .B2(n7190), .A(n9521), .ZN(n7202) );
  NAND2_X1 U9107 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8043) );
  OAI21_X1 U9108 ( .B1(n9596), .B2(n10310), .A(n8043), .ZN(n7200) );
  XNOR2_X1 U9109 ( .A(n7280), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n7197) );
  OAI22_X1 U9110 ( .A1(n7195), .A2(n7194), .B1(n7193), .B2(n7192), .ZN(n7196)
         );
  NOR2_X1 U9111 ( .A1(n7196), .A2(n7197), .ZN(n7284) );
  AOI21_X1 U9112 ( .B1(n7197), .B2(n7196), .A(n7284), .ZN(n7198) );
  NOR2_X1 U9113 ( .A1(n7198), .A2(n9556), .ZN(n7199) );
  AOI211_X1 U9114 ( .C1(n10054), .C2(n7280), .A(n7200), .B(n7199), .ZN(n7201)
         );
  OAI21_X1 U9115 ( .B1(n7202), .B2(n9561), .A(n7201), .ZN(P1_U3255) );
  INV_X1 U9116 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10023) );
  NAND2_X1 U9117 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7979) );
  OAI21_X1 U9118 ( .B1(n9596), .B2(n10023), .A(n7979), .ZN(n7209) );
  OR2_X1 U9119 ( .A1(n7204), .A2(n7203), .ZN(n7206) );
  AOI211_X1 U9120 ( .C1(n7207), .C2(n7206), .A(n9556), .B(n7205), .ZN(n7208)
         );
  AOI211_X1 U9121 ( .C1(n10054), .C2(n7210), .A(n7209), .B(n7208), .ZN(n7218)
         );
  INV_X1 U9122 ( .A(n7211), .ZN(n7216) );
  OAI21_X1 U9123 ( .B1(n7214), .B2(n7213), .A(n7212), .ZN(n7215) );
  NAND3_X1 U9124 ( .A1(n7216), .A2(n10061), .A3(n7215), .ZN(n7217) );
  NAND2_X1 U9125 ( .A1(n7218), .A2(n7217), .ZN(P1_U3253) );
  NOR2_X1 U9126 ( .A1(n10063), .A2(P1_U3973), .ZN(P1_U3085) );
  OAI211_X1 U9127 ( .C1(n7221), .C2(n7220), .A(n7219), .B(n8679), .ZN(n7226)
         );
  OAI22_X1 U9128 ( .A1(n7385), .A2(n8707), .B1(n8724), .B2(n7440), .ZN(n7224)
         );
  OAI21_X1 U9129 ( .B1(n8731), .B2(n7419), .A(n7222), .ZN(n7223) );
  AOI211_X1 U9130 ( .C1(n7483), .C2(n8727), .A(n7224), .B(n7223), .ZN(n7225)
         );
  NAND2_X1 U9131 ( .A1(n7226), .A2(n7225), .ZN(P2_U3158) );
  INV_X1 U9132 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7228) );
  INV_X1 U9133 ( .A(n7227), .ZN(n7229) );
  INV_X1 U9134 ( .A(n9518), .ZN(n7287) );
  OAI222_X1 U9135 ( .A1(n10002), .A2(n7228), .B1(n8589), .B2(n7229), .C1(
        P1_U3086), .C2(n7287), .ZN(P1_U3342) );
  INV_X1 U9136 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7230) );
  OAI222_X1 U9137 ( .A1(n9062), .A2(n7230), .B1(n9063), .B2(n7229), .C1(
        P2_U3151), .C2(n8778), .ZN(P2_U3282) );
  INV_X1 U9138 ( .A(n7231), .ZN(n7232) );
  AOI21_X1 U9139 ( .B1(n7234), .B2(n7233), .A(n7232), .ZN(n7249) );
  NAND2_X1 U9140 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7692) );
  OAI21_X1 U9141 ( .B1(n8846), .B2(n7235), .A(n7692), .ZN(n7242) );
  INV_X1 U9142 ( .A(n7236), .ZN(n7240) );
  NAND3_X1 U9143 ( .A1(n7156), .A2(n7238), .A3(n7237), .ZN(n7239) );
  AOI21_X1 U9144 ( .B1(n7240), .B2(n7239), .A(n8856), .ZN(n7241) );
  AOI211_X1 U9145 ( .C1(n8848), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n7242), .B(
        n7241), .ZN(n7248) );
  INV_X1 U9146 ( .A(n7243), .ZN(n7246) );
  NOR3_X1 U9147 ( .A1(n4310), .A2(n4414), .A3(n7244), .ZN(n7245) );
  OAI21_X1 U9148 ( .B1(n7246), .B2(n7245), .A(n8853), .ZN(n7247) );
  OAI211_X1 U9149 ( .C1(n7249), .C2(n8850), .A(n7248), .B(n7247), .ZN(P2_U3188) );
  INV_X1 U9150 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n7257) );
  OAI21_X1 U9151 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n7251), .A(n7250), .ZN(n7252) );
  OAI21_X1 U9152 ( .B1(n7253), .B2(n8766), .A(n7252), .ZN(n7254) );
  OAI21_X1 U9153 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7451), .A(n7254), .ZN(n7255) );
  AOI21_X1 U9154 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n8764), .A(n7255), .ZN(n7256) );
  OAI21_X1 U9155 ( .B1(n8088), .B2(n7257), .A(n7256), .ZN(P2_U3182) );
  INV_X1 U9156 ( .A(n7299), .ZN(n7258) );
  NAND2_X1 U9157 ( .A1(n8334), .A2(n8754), .ZN(n8343) );
  OR2_X1 U9158 ( .A1(n8727), .A2(P2_U3151), .ZN(n7338) );
  NAND2_X1 U9159 ( .A1(n7338), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7260) );
  AOI22_X1 U9160 ( .A1(n8704), .A2(n6091), .B1(n8711), .B2(n10154), .ZN(n7259)
         );
  OAI211_X1 U9161 ( .C1(n10150), .C2(n8717), .A(n7260), .B(n7259), .ZN(
        P2_U3172) );
  NAND2_X1 U9162 ( .A1(n7261), .A2(n7262), .ZN(n7263) );
  XOR2_X1 U9163 ( .A(n7264), .B(n7263), .Z(n7270) );
  OR2_X1 U9164 ( .A1(n7265), .A2(P1_U3086), .ZN(n7541) );
  NAND2_X1 U9165 ( .A1(n9834), .A2(n9431), .ZN(n7403) );
  OAI22_X1 U9166 ( .A1(n7266), .A2(n7403), .B1(n10080), .B2(n9186), .ZN(n7268)
         );
  INV_X1 U9167 ( .A(n6739), .ZN(n7405) );
  NOR2_X1 U9168 ( .A1(n8264), .A2(n7405), .ZN(n7267) );
  AOI211_X1 U9169 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n7541), .A(n7268), .B(
        n7267), .ZN(n7269) );
  OAI21_X1 U9170 ( .B1(n7270), .B2(n9170), .A(n7269), .ZN(P1_U3222) );
  INV_X1 U9171 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7273) );
  AND2_X1 U9172 ( .A1(n6739), .A2(n7425), .ZN(n9361) );
  NOR2_X1 U9173 ( .A1(n7402), .A2(n9361), .ZN(n9280) );
  INV_X1 U9174 ( .A(n9280), .ZN(n7654) );
  OAI21_X1 U9175 ( .B1(n9829), .B2(n10112), .A(n7654), .ZN(n7271) );
  NAND2_X1 U9176 ( .A1(n9834), .A2(n6725), .ZN(n7655) );
  OAI211_X1 U9177 ( .C1(n7652), .C2(n7425), .A(n7271), .B(n7655), .ZN(n9935)
         );
  NAND2_X1 U9178 ( .A1(n9935), .A2(n10115), .ZN(n7272) );
  OAI21_X1 U9179 ( .B1(n10115), .B2(n7273), .A(n7272), .ZN(P1_U3453) );
  XOR2_X1 U9180 ( .A(n7275), .B(n7274), .Z(n7279) );
  AOI22_X1 U9181 ( .A1(n8722), .A2(n8754), .B1(n8711), .B2(n10156), .ZN(n7276)
         );
  OAI21_X1 U9182 ( .B1(n7385), .B2(n8724), .A(n7276), .ZN(n7277) );
  AOI21_X1 U9183 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7338), .A(n7277), .ZN(
        n7278) );
  OAI21_X1 U9184 ( .B1(n8717), .B2(n7279), .A(n7278), .ZN(P2_U3162) );
  NOR2_X1 U9185 ( .A1(n7280), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9520) );
  XNOR2_X1 U9186 ( .A(n9518), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9519) );
  XNOR2_X1 U9187 ( .A(n7320), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n7681) );
  XNOR2_X1 U9188 ( .A(n7682), .B(n7681), .ZN(n7296) );
  INV_X1 U9189 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7281) );
  NAND2_X1 U9190 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8134) );
  OAI21_X1 U9191 ( .B1(n9596), .B2(n7281), .A(n8134), .ZN(n7282) );
  AOI21_X1 U9192 ( .B1(n7320), .B2(n10054), .A(n7282), .ZN(n7295) );
  INV_X1 U9193 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7283) );
  MUX2_X1 U9194 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n7283), .S(n7320), .Z(n7289)
         );
  INV_X1 U9195 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7288) );
  AOI22_X1 U9196 ( .A1(n9518), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7288), .B2(
        n7287), .ZN(n9513) );
  INV_X1 U9197 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7285) );
  NAND2_X1 U9198 ( .A1(n9513), .A2(n9514), .ZN(n9512) );
  OAI21_X1 U9199 ( .B1(n7288), .B2(n7287), .A(n9512), .ZN(n7290) );
  NAND2_X1 U9200 ( .A1(n7289), .A2(n7290), .ZN(n7684) );
  MUX2_X1 U9201 ( .A(n7283), .B(P1_REG2_REG_14__SCAN_IN), .S(n7320), .Z(n7292)
         );
  INV_X1 U9202 ( .A(n7290), .ZN(n7291) );
  NAND2_X1 U9203 ( .A1(n7292), .A2(n7291), .ZN(n7293) );
  NAND3_X1 U9204 ( .A1(n10052), .A2(n7684), .A3(n7293), .ZN(n7294) );
  OAI211_X1 U9205 ( .C1(n7296), .C2(n9561), .A(n7295), .B(n7294), .ZN(P1_U3257) );
  INV_X1 U9206 ( .A(n9273), .ZN(n9338) );
  NAND2_X1 U9207 ( .A1(P1_U3973), .A2(n9338), .ZN(n7297) );
  OAI21_X1 U9208 ( .B1(P1_U3973), .B2(n5556), .A(n7297), .ZN(P1_U3585) );
  OAI21_X1 U9209 ( .B1(n8345), .B2(n7299), .A(n7298), .ZN(n10158) );
  INV_X1 U9210 ( .A(n10158), .ZN(n7317) );
  NAND2_X1 U9211 ( .A1(n7303), .A2(n7300), .ZN(n7301) );
  OAI211_X1 U9212 ( .C1(n6044), .C2(n7303), .A(n7302), .B(n7301), .ZN(n7314)
         );
  NAND2_X1 U9213 ( .A1(n8338), .A2(n7304), .ZN(n7458) );
  INV_X1 U9214 ( .A(n7458), .ZN(n10144) );
  NAND2_X1 U9215 ( .A1(n10145), .A2(n10144), .ZN(n7745) );
  OAI21_X1 U9216 ( .B1(n7307), .B2(n7306), .A(n7305), .ZN(n7308) );
  NAND2_X1 U9217 ( .A1(n7308), .A2(n10136), .ZN(n7312) );
  AOI22_X1 U9218 ( .A1(n10132), .A2(n8754), .B1(n10131), .B2(n6094), .ZN(n7311) );
  INV_X1 U9219 ( .A(n10141), .ZN(n7309) );
  NAND2_X1 U9220 ( .A1(n10158), .A2(n7309), .ZN(n7310) );
  AND3_X1 U9221 ( .A1(n7312), .A2(n7311), .A3(n7310), .ZN(n10160) );
  MUX2_X1 U9222 ( .A(n7313), .B(n10160), .S(n10145), .Z(n7316) );
  AOI22_X1 U9223 ( .A1(n8955), .A2(n10156), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8954), .ZN(n7315) );
  OAI211_X1 U9224 ( .C1(n7317), .C2(n7745), .A(n7316), .B(n7315), .ZN(P2_U3232) );
  NAND2_X1 U9225 ( .A1(n4580), .A2(P1_U3973), .ZN(n7318) );
  OAI21_X1 U9226 ( .B1(P1_U3973), .B2(n5227), .A(n7318), .ZN(P1_U3562) );
  INV_X1 U9227 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7321) );
  INV_X1 U9228 ( .A(n7319), .ZN(n7322) );
  INV_X1 U9229 ( .A(n7320), .ZN(n7685) );
  OAI222_X1 U9230 ( .A1(n10002), .A2(n7321), .B1(n8589), .B2(n7322), .C1(
        P1_U3086), .C2(n7685), .ZN(P1_U3341) );
  INV_X1 U9231 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7323) );
  OAI222_X1 U9232 ( .A1(n9062), .A2(n7323), .B1(n9063), .B2(n7322), .C1(
        P2_U3151), .C2(n8794), .ZN(P2_U3281) );
  INV_X1 U9233 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n10313) );
  NAND2_X1 U9234 ( .A1(P1_U3973), .A2(n6739), .ZN(n7324) );
  OAI21_X1 U9235 ( .B1(P1_U3973), .B2(n10313), .A(n7324), .ZN(P1_U3554) );
  XOR2_X1 U9236 ( .A(n7326), .B(n7325), .Z(n7335) );
  OAI21_X1 U9237 ( .B1(n4407), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7374), .ZN(
        n7333) );
  AOI21_X1 U9238 ( .B1(n10266), .B2(n7327), .A(n7366), .ZN(n7331) );
  NAND2_X1 U9239 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7806) );
  OAI21_X1 U9240 ( .B1(n8846), .B2(n7328), .A(n7806), .ZN(n7329) );
  AOI21_X1 U9241 ( .B1(n8848), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7329), .ZN(
        n7330) );
  OAI21_X1 U9242 ( .B1(n7331), .B2(n8856), .A(n7330), .ZN(n7332) );
  AOI21_X1 U9243 ( .B1(n8853), .B2(n7333), .A(n7332), .ZN(n7334) );
  OAI21_X1 U9244 ( .B1(n7335), .B2(n8850), .A(n7334), .ZN(P2_U3189) );
  XNOR2_X1 U9245 ( .A(n7337), .B(n7336), .ZN(n7343) );
  NAND2_X1 U9246 ( .A1(n7338), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7341) );
  AOI22_X1 U9247 ( .A1(n8722), .A2(n6091), .B1(n8711), .B2(n7339), .ZN(n7340)
         );
  OAI211_X1 U9248 ( .C1(n7353), .C2(n8724), .A(n7341), .B(n7340), .ZN(n7342)
         );
  AOI21_X1 U9249 ( .B1(n7343), .B2(n8679), .A(n7342), .ZN(n7344) );
  INV_X1 U9250 ( .A(n7344), .ZN(P2_U3177) );
  INV_X1 U9251 ( .A(n7345), .ZN(n7360) );
  AOI22_X1 U9252 ( .A1(n9533), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n7346), .ZN(n7347) );
  OAI21_X1 U9253 ( .B1(n7360), .B2(n8589), .A(n7347), .ZN(P1_U3340) );
  AOI21_X1 U9254 ( .B1(n7350), .B2(n7349), .A(n7348), .ZN(n7359) );
  INV_X1 U9255 ( .A(n7351), .ZN(n7355) );
  OAI22_X1 U9256 ( .A1(n7353), .A2(n8707), .B1(n8724), .B2(n7352), .ZN(n7354)
         );
  AOI211_X1 U9257 ( .C1(n7466), .C2(n8711), .A(n7355), .B(n7354), .ZN(n7358)
         );
  INV_X1 U9258 ( .A(n7356), .ZN(n7465) );
  NAND2_X1 U9259 ( .A1(n8727), .A2(n7465), .ZN(n7357) );
  OAI211_X1 U9260 ( .C1(n7359), .C2(n8717), .A(n7358), .B(n7357), .ZN(P2_U3170) );
  INV_X1 U9261 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7361) );
  OAI222_X1 U9262 ( .A1(n9062), .A2(n7361), .B1(n9063), .B2(n7360), .C1(
        P2_U3151), .C2(n8815), .ZN(P2_U3280) );
  XOR2_X1 U9263 ( .A(n7363), .B(n7362), .Z(n7381) );
  INV_X1 U9264 ( .A(n7364), .ZN(n7369) );
  NOR3_X1 U9265 ( .A1(n7367), .A2(n7366), .A3(n7365), .ZN(n7368) );
  OAI21_X1 U9266 ( .B1(n7369), .B2(n7368), .A(n8825), .ZN(n7380) );
  NAND2_X1 U9267 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7921) );
  OAI21_X1 U9268 ( .B1(n8846), .B2(n7370), .A(n7921), .ZN(n7378) );
  INV_X1 U9269 ( .A(n7371), .ZN(n7373) );
  NAND3_X1 U9270 ( .A1(n7374), .A2(n7373), .A3(n7372), .ZN(n7375) );
  AOI21_X1 U9271 ( .B1(n7376), .B2(n7375), .A(n8835), .ZN(n7377) );
  AOI211_X1 U9272 ( .C1(n8848), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7378), .B(
        n7377), .ZN(n7379) );
  OAI211_X1 U9273 ( .C1(n7381), .C2(n8850), .A(n7380), .B(n7379), .ZN(P2_U3190) );
  INV_X1 U9274 ( .A(n7382), .ZN(n8362) );
  NAND2_X1 U9275 ( .A1(n8362), .A2(n8354), .ZN(n8282) );
  XNOR2_X1 U9276 ( .A(n7383), .B(n8282), .ZN(n7387) );
  NAND2_X1 U9277 ( .A1(n10131), .A2(n8753), .ZN(n7384) );
  OAI21_X1 U9278 ( .B1(n8946), .B2(n7385), .A(n7384), .ZN(n7386) );
  AOI21_X1 U9279 ( .B1(n7387), .B2(n10136), .A(n7386), .ZN(n7481) );
  OR2_X1 U9280 ( .A1(n10127), .A2(n10126), .ZN(n10124) );
  NAND2_X1 U9281 ( .A1(n10124), .A2(n8348), .ZN(n7389) );
  INV_X1 U9282 ( .A(n8282), .ZN(n7388) );
  NAND2_X1 U9283 ( .A1(n7389), .A2(n7388), .ZN(n7430) );
  OAI21_X1 U9284 ( .B1(n7389), .B2(n7388), .A(n7430), .ZN(n7480) );
  NAND2_X1 U9285 ( .A1(n7480), .A2(n6186), .ZN(n7390) );
  NAND2_X1 U9286 ( .A1(n7481), .A2(n7390), .ZN(n7421) );
  MUX2_X1 U9287 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n7421), .S(n10199), .Z(n7391)
         );
  AOI21_X1 U9288 ( .B1(n8983), .B2(n7484), .A(n7391), .ZN(n7392) );
  INV_X1 U9289 ( .A(n7392), .ZN(P2_U3462) );
  INV_X1 U9290 ( .A(n7393), .ZN(n7395) );
  INV_X1 U9291 ( .A(n9535), .ZN(n9551) );
  OAI222_X1 U9292 ( .A1(n10002), .A2(n7394), .B1(n8589), .B2(n7395), .C1(n9551), .C2(P1_U3086), .ZN(P1_U3339) );
  OAI222_X1 U9293 ( .A1(n9062), .A2(n10323), .B1(P2_U3151), .B2(n4929), .C1(
        n7395), .C2(n9063), .ZN(P2_U3279) );
  INV_X1 U9294 ( .A(n9568), .ZN(n9553) );
  INV_X1 U9295 ( .A(n7396), .ZN(n7397) );
  OAI222_X1 U9296 ( .A1(P1_U3086), .A2(n9553), .B1(n8589), .B2(n7397), .C1(
        n10002), .C2(n5260), .ZN(P1_U3338) );
  OAI222_X1 U9297 ( .A1(n9062), .A2(n7398), .B1(n9063), .B2(n7397), .C1(
        P2_U3151), .C2(n8845), .ZN(P2_U3278) );
  INV_X1 U9298 ( .A(n9933), .ZN(n7757) );
  OAI21_X1 U9299 ( .B1(n6627), .B2(n7401), .A(n7400), .ZN(n10070) );
  OAI211_X1 U9300 ( .C1(n10080), .C2(n7425), .A(n9894), .B(n7413), .ZN(n10074)
         );
  INV_X1 U9301 ( .A(n10074), .ZN(n7409) );
  XNOR2_X1 U9302 ( .A(n7399), .B(n7402), .ZN(n7407) );
  INV_X1 U9303 ( .A(n7637), .ZN(n7842) );
  NAND2_X1 U9304 ( .A1(n10070), .A2(n7842), .ZN(n7404) );
  OAI211_X1 U9305 ( .C1(n7405), .C2(n9800), .A(n7404), .B(n7403), .ZN(n7406)
         );
  AOI21_X1 U9306 ( .B1(n7407), .B2(n9829), .A(n7406), .ZN(n10085) );
  INV_X1 U9307 ( .A(n10085), .ZN(n7408) );
  AOI211_X1 U9308 ( .C1(n7757), .C2(n10070), .A(n7409), .B(n7408), .ZN(n7457)
         );
  AOI22_X1 U9309 ( .A1(n9884), .A2(n6726), .B1(n10120), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n7410) );
  OAI21_X1 U9310 ( .B1(n7457), .B2(n10120), .A(n7410), .ZN(P1_U3523) );
  OAI21_X1 U9311 ( .B1(n7412), .B2(n4285), .A(n7411), .ZN(n7856) );
  NAND2_X1 U9312 ( .A1(n7413), .A2(n9363), .ZN(n7414) );
  NAND2_X1 U9313 ( .A1(n9894), .A2(n7414), .ZN(n7415) );
  NOR2_X1 U9314 ( .A1(n7415), .A2(n7670), .ZN(n7852) );
  XNOR2_X1 U9315 ( .A(n7416), .B(n4285), .ZN(n7417) );
  OAI222_X1 U9316 ( .A1(n9800), .A2(n7539), .B1(n9802), .B2(n7646), .C1(n9797), 
        .C2(n7417), .ZN(n7851) );
  AOI211_X1 U9317 ( .C1(n10112), .C2(n7856), .A(n7852), .B(n7851), .ZN(n7429)
         );
  AOI22_X1 U9318 ( .A1(n9884), .A2(n9363), .B1(n10120), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n7418) );
  OAI21_X1 U9319 ( .B1(n7429), .B2(n10120), .A(n7418), .ZN(P1_U3524) );
  OAI22_X1 U9320 ( .A1(n9044), .A2(n7419), .B1(n5729), .B2(n10184), .ZN(n7420)
         );
  AOI21_X1 U9321 ( .B1(n7421), .B2(n10184), .A(n7420), .ZN(n7422) );
  INV_X1 U9322 ( .A(n7422), .ZN(P2_U3399) );
  XNOR2_X1 U9323 ( .A(n7423), .B(n7424), .ZN(n9454) );
  OAI22_X1 U9324 ( .A1(n9181), .A2(n7539), .B1(n9186), .B2(n7425), .ZN(n7426)
         );
  AOI21_X1 U9325 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n7541), .A(n7426), .ZN(
        n7427) );
  OAI21_X1 U9326 ( .B1(n9170), .B2(n9454), .A(n7427), .ZN(P1_U3232) );
  AOI22_X1 U9327 ( .A1(n9954), .A2(n9363), .B1(n10113), .B2(
        P1_REG0_REG_2__SCAN_IN), .ZN(n7428) );
  OAI21_X1 U9328 ( .B1(n7429), .B2(n10113), .A(n7428), .ZN(P1_U3459) );
  NAND2_X1 U9329 ( .A1(n7430), .A2(n8354), .ZN(n7461) );
  INV_X1 U9330 ( .A(n8363), .ZN(n7431) );
  OAI21_X1 U9331 ( .B1(n7461), .B2(n7431), .A(n7460), .ZN(n7434) );
  NAND2_X1 U9332 ( .A1(n7433), .A2(n7432), .ZN(n8284) );
  XNOR2_X1 U9333 ( .A(n7434), .B(n8284), .ZN(n10173) );
  AND2_X1 U9334 ( .A1(n7436), .A2(n7435), .ZN(n7462) );
  AOI21_X1 U9335 ( .B1(n7462), .B2(n7438), .A(n7437), .ZN(n7439) );
  XOR2_X1 U9336 ( .A(n8284), .B(n7439), .Z(n7443) );
  OAI22_X1 U9337 ( .A1(n4652), .A2(n7474), .B1(n7440), .B2(n8946), .ZN(n7442)
         );
  NOR2_X1 U9338 ( .A1(n10173), .A2(n10141), .ZN(n7441) );
  AOI211_X1 U9339 ( .C1(n10136), .C2(n7443), .A(n7442), .B(n7441), .ZN(n10170)
         );
  MUX2_X1 U9340 ( .A(n7444), .B(n10170), .S(n10145), .Z(n7448) );
  INV_X1 U9341 ( .A(n7445), .ZN(n7477) );
  AOI22_X1 U9342 ( .A1(n8955), .A2(n7446), .B1(n8954), .B2(n7477), .ZN(n7447)
         );
  OAI211_X1 U9343 ( .C1(n10173), .C2(n7745), .A(n7448), .B(n7447), .ZN(
        P2_U3228) );
  NAND2_X1 U9344 ( .A1(n10131), .A2(n6091), .ZN(n10149) );
  OAI21_X1 U9345 ( .B1(n10150), .B2(n7449), .A(n10149), .ZN(n7450) );
  MUX2_X1 U9346 ( .A(P2_REG2_REG_0__SCAN_IN), .B(n7450), .S(n10145), .Z(n7453)
         );
  OAI22_X1 U9347 ( .A1(n8925), .A2(n8334), .B1(n7451), .B2(n10129), .ZN(n7452)
         );
  OR2_X1 U9348 ( .A1(n7453), .A2(n7452), .ZN(P2_U3233) );
  INV_X1 U9349 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7454) );
  OAI22_X1 U9350 ( .A1(n9975), .A2(n10080), .B1(n10115), .B2(n7454), .ZN(n7455) );
  INV_X1 U9351 ( .A(n7455), .ZN(n7456) );
  OAI21_X1 U9352 ( .B1(n7457), .B2(n10113), .A(n7456), .ZN(P1_U3456) );
  NAND2_X1 U9353 ( .A1(n10141), .A2(n7458), .ZN(n7459) );
  AND2_X1 U9354 ( .A1(n7460), .A2(n8363), .ZN(n8353) );
  XNOR2_X1 U9355 ( .A(n7461), .B(n8353), .ZN(n10169) );
  INV_X1 U9356 ( .A(n10169), .ZN(n7469) );
  XNOR2_X1 U9357 ( .A(n7462), .B(n8353), .ZN(n7463) );
  AOI222_X1 U9358 ( .A1(n10136), .A2(n7463), .B1(n8752), .B2(n10131), .C1(
        n10130), .C2(n10132), .ZN(n10166) );
  MUX2_X1 U9359 ( .A(n7464), .B(n10166), .S(n10145), .Z(n7468) );
  AOI22_X1 U9360 ( .A1(n8955), .A2(n7466), .B1(n8954), .B2(n7465), .ZN(n7467)
         );
  OAI211_X1 U9361 ( .C1(n8958), .C2(n7469), .A(n7468), .B(n7467), .ZN(P2_U3229) );
  XOR2_X1 U9362 ( .A(n7471), .B(n7470), .Z(n7479) );
  NAND2_X1 U9363 ( .A1(n8722), .A2(n8753), .ZN(n7473) );
  OAI211_X1 U9364 ( .C1(n7474), .C2(n8724), .A(n7473), .B(n7472), .ZN(n7476)
         );
  NOR2_X1 U9365 ( .A1(n8731), .A2(n10171), .ZN(n7475) );
  AOI211_X1 U9366 ( .C1(n7477), .C2(n8727), .A(n7476), .B(n7475), .ZN(n7478)
         );
  OAI21_X1 U9367 ( .B1(n7479), .B2(n8717), .A(n7478), .ZN(P2_U3167) );
  INV_X1 U9368 ( .A(n7480), .ZN(n7487) );
  MUX2_X1 U9369 ( .A(n7482), .B(n7481), .S(n10145), .Z(n7486) );
  AOI22_X1 U9370 ( .A1(n8955), .A2(n7484), .B1(n8954), .B2(n7483), .ZN(n7485)
         );
  OAI211_X1 U9371 ( .C1(n7487), .C2(n8958), .A(n7486), .B(n7485), .ZN(P2_U3230) );
  INV_X1 U9372 ( .A(n8285), .ZN(n7489) );
  OR2_X1 U9373 ( .A1(n4399), .A2(n7489), .ZN(n7500) );
  INV_X1 U9374 ( .A(n7500), .ZN(n7488) );
  AOI21_X1 U9375 ( .B1(n4399), .B2(n7489), .A(n7488), .ZN(n10181) );
  XNOR2_X1 U9376 ( .A(n7505), .B(n8285), .ZN(n7490) );
  AOI222_X1 U9377 ( .A1(n10136), .A2(n7490), .B1(n8750), .B2(n10131), .C1(
        n8752), .C2(n10132), .ZN(n10177) );
  MUX2_X1 U9378 ( .A(n7491), .B(n10177), .S(n10145), .Z(n7494) );
  INV_X1 U9379 ( .A(n7492), .ZN(n7691) );
  AOI22_X1 U9380 ( .A1(n8955), .A2(n7702), .B1(n8954), .B2(n7691), .ZN(n7493)
         );
  OAI211_X1 U9381 ( .C1(n10181), .C2(n8958), .A(n7494), .B(n7493), .ZN(
        P2_U3227) );
  INV_X1 U9382 ( .A(n7495), .ZN(n7498) );
  INV_X1 U9383 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7496) );
  OAI222_X1 U9384 ( .A1(P2_U3151), .A2(n7497), .B1(n9063), .B2(n7498), .C1(
        n7496), .C2(n9062), .ZN(P2_U3277) );
  INV_X1 U9385 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7499) );
  INV_X1 U9386 ( .A(n9583), .ZN(n9579) );
  OAI222_X1 U9387 ( .A1(n10002), .A2(n7499), .B1(n8589), .B2(n7498), .C1(n9579), .C2(P1_U3086), .ZN(P1_U3337) );
  INV_X1 U9388 ( .A(n10172), .ZN(n10165) );
  NAND2_X1 U9389 ( .A1(n7500), .A2(n8366), .ZN(n7503) );
  INV_X1 U9390 ( .A(n7503), .ZN(n7501) );
  XNOR2_X1 U9391 ( .A(n7572), .B(n8750), .ZN(n8375) );
  NAND2_X1 U9392 ( .A1(n7501), .A2(n8375), .ZN(n7569) );
  INV_X1 U9393 ( .A(n8375), .ZN(n7502) );
  NAND2_X1 U9394 ( .A1(n7503), .A2(n7502), .ZN(n7504) );
  NAND2_X1 U9395 ( .A1(n7569), .A2(n7504), .ZN(n7513) );
  INV_X1 U9396 ( .A(n7513), .ZN(n7601) );
  OAI21_X1 U9397 ( .B1(n7505), .B2(n8751), .A(n7702), .ZN(n7507) );
  NAND2_X1 U9398 ( .A1(n7505), .A2(n8751), .ZN(n7506) );
  NAND2_X1 U9399 ( .A1(n7507), .A2(n7506), .ZN(n7508) );
  OR2_X1 U9400 ( .A1(n7508), .A2(n8375), .ZN(n7571) );
  NAND2_X1 U9401 ( .A1(n7508), .A2(n8375), .ZN(n7509) );
  NAND2_X1 U9402 ( .A1(n7571), .A2(n7509), .ZN(n7510) );
  NAND2_X1 U9403 ( .A1(n7510), .A2(n10136), .ZN(n7512) );
  AOI22_X1 U9404 ( .A1(n10132), .A2(n8751), .B1(n10131), .B2(n8749), .ZN(n7511) );
  OAI211_X1 U9405 ( .C1(n7513), .C2(n10141), .A(n7512), .B(n7511), .ZN(n7598)
         );
  AOI21_X1 U9406 ( .B1(n10165), .B2(n7601), .A(n7598), .ZN(n7515) );
  MUX2_X1 U9407 ( .A(n10311), .B(n7515), .S(n10184), .Z(n7514) );
  OAI21_X1 U9408 ( .B1(n7803), .B2(n9044), .A(n7514), .ZN(P2_U3411) );
  MUX2_X1 U9409 ( .A(n10266), .B(n7515), .S(n10199), .Z(n7516) );
  OAI21_X1 U9410 ( .B1(n7803), .B2(n8991), .A(n7516), .ZN(P2_U3466) );
  XNOR2_X1 U9411 ( .A(n7517), .B(n8289), .ZN(n7523) );
  INV_X1 U9412 ( .A(n7523), .ZN(n7738) );
  INV_X1 U9413 ( .A(n8289), .ZN(n7519) );
  XNOR2_X1 U9414 ( .A(n7518), .B(n7519), .ZN(n7520) );
  NAND2_X1 U9415 ( .A1(n7520), .A2(n10136), .ZN(n7522) );
  AOI22_X1 U9416 ( .A1(n10132), .A2(n8749), .B1(n10131), .B2(n8747), .ZN(n7521) );
  OAI211_X1 U9417 ( .C1(n7523), .C2(n10141), .A(n7522), .B(n7521), .ZN(n7734)
         );
  AOI21_X1 U9418 ( .B1(n10165), .B2(n7738), .A(n7734), .ZN(n7628) );
  AOI22_X1 U9419 ( .A1(n6375), .A2(n7627), .B1(n10186), .B2(
        P2_REG0_REG_9__SCAN_IN), .ZN(n7524) );
  OAI21_X1 U9420 ( .B1(n7628), .B2(n10186), .A(n7524), .ZN(P2_U3417) );
  AOI21_X1 U9421 ( .B1(n7526), .B2(n7525), .A(n7880), .ZN(n7533) );
  NAND2_X1 U9422 ( .A1(n9183), .A2(n7910), .ZN(n7529) );
  AOI21_X1 U9423 ( .B1(n9177), .B2(n9427), .A(n7527), .ZN(n7528) );
  OAI211_X1 U9424 ( .C1(n7530), .C2(n9181), .A(n7529), .B(n7528), .ZN(n7531)
         );
  AOI21_X1 U9425 ( .B1(n9168), .B2(n7911), .A(n7531), .ZN(n7532) );
  OAI21_X1 U9426 ( .B1(n7533), .B2(n9170), .A(n7532), .ZN(P1_U3213) );
  INV_X1 U9427 ( .A(n7535), .ZN(n7536) );
  AOI21_X1 U9428 ( .B1(n7537), .B2(n7534), .A(n7536), .ZN(n7543) );
  AOI22_X1 U9429 ( .A1(n9155), .A2(n9430), .B1(n9168), .B2(n9363), .ZN(n7538)
         );
  OAI21_X1 U9430 ( .B1(n7539), .B2(n8264), .A(n7538), .ZN(n7540) );
  AOI21_X1 U9431 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n7541), .A(n7540), .ZN(
        n7542) );
  OAI21_X1 U9432 ( .B1(n7543), .B2(n9170), .A(n7542), .ZN(P1_U3237) );
  INV_X1 U9433 ( .A(n7899), .ZN(n7551) );
  XNOR2_X1 U9434 ( .A(n7617), .B(n7544), .ZN(n7545) );
  NAND2_X1 U9435 ( .A1(n7545), .A2(n7546), .ZN(n7616) );
  OAI21_X1 U9436 ( .B1(n7546), .B2(n7545), .A(n7616), .ZN(n7547) );
  NAND2_X1 U9437 ( .A1(n7547), .A2(n9175), .ZN(n7550) );
  AND2_X1 U9438 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9479) );
  OAI22_X1 U9439 ( .A1(n8264), .A2(n7666), .B1(n9200), .B2(n9181), .ZN(n7548)
         );
  AOI211_X1 U9440 ( .C1(n9168), .C2(n7900), .A(n9479), .B(n7548), .ZN(n7549)
         );
  OAI211_X1 U9441 ( .C1(n9164), .C2(n7551), .A(n7550), .B(n7549), .ZN(P1_U3227) );
  XOR2_X1 U9442 ( .A(n7553), .B(n7552), .Z(n7568) );
  NOR3_X1 U9443 ( .A1(n7608), .A2(n7555), .A3(n7554), .ZN(n7556) );
  OAI21_X1 U9444 ( .B1(n4409), .B2(n7556), .A(n8825), .ZN(n7567) );
  NAND2_X1 U9445 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8190) );
  OAI21_X1 U9446 ( .B1(n8846), .B2(n7557), .A(n8190), .ZN(n7565) );
  INV_X1 U9447 ( .A(n7559), .ZN(n7561) );
  NAND3_X1 U9448 ( .A1(n7558), .A2(n7561), .A3(n7560), .ZN(n7562) );
  AOI21_X1 U9449 ( .B1(n7563), .B2(n7562), .A(n8835), .ZN(n7564) );
  AOI211_X1 U9450 ( .C1(n8848), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n7565), .B(
        n7564), .ZN(n7566) );
  OAI211_X1 U9451 ( .C1(n7568), .C2(n8850), .A(n7567), .B(n7566), .ZN(P2_U3192) );
  OR2_X1 U9452 ( .A1(n7572), .A2(n7696), .ZN(n8378) );
  NAND2_X1 U9453 ( .A1(n7569), .A2(n8378), .ZN(n7570) );
  XOR2_X1 U9454 ( .A(n8288), .B(n7570), .Z(n7590) );
  INV_X1 U9455 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7579) );
  OAI21_X1 U9456 ( .B1(n8750), .B2(n7572), .A(n7571), .ZN(n7576) );
  INV_X1 U9457 ( .A(n8288), .ZN(n7575) );
  INV_X1 U9458 ( .A(n10136), .ZN(n10151) );
  INV_X1 U9459 ( .A(n7573), .ZN(n7574) );
  AOI211_X1 U9460 ( .C1(n7576), .C2(n7575), .A(n10151), .B(n7574), .ZN(n7578)
         );
  OAI22_X1 U9461 ( .A1(n4652), .A2(n7923), .B1(n7696), .B2(n8946), .ZN(n7577)
         );
  NOR2_X1 U9462 ( .A1(n7578), .A2(n7577), .ZN(n7585) );
  MUX2_X1 U9463 ( .A(n7579), .B(n7585), .S(n10184), .Z(n7581) );
  NAND2_X1 U9464 ( .A1(n6375), .A2(n7927), .ZN(n7580) );
  OAI211_X1 U9465 ( .C1(n7590), .C2(n9039), .A(n7581), .B(n7580), .ZN(P2_U3414) );
  MUX2_X1 U9466 ( .A(n7582), .B(n7585), .S(n10199), .Z(n7584) );
  NAND2_X1 U9467 ( .A1(n8983), .A2(n7927), .ZN(n7583) );
  OAI211_X1 U9468 ( .C1(n7590), .C2(n8986), .A(n7584), .B(n7583), .ZN(P2_U3467) );
  MUX2_X1 U9469 ( .A(n7586), .B(n7585), .S(n10145), .Z(n7589) );
  INV_X1 U9470 ( .A(n7924), .ZN(n7587) );
  AOI22_X1 U9471 ( .A1(n8955), .A2(n7927), .B1(n8954), .B2(n7587), .ZN(n7588)
         );
  OAI211_X1 U9472 ( .C1(n7590), .C2(n8958), .A(n7589), .B(n7588), .ZN(P2_U3225) );
  XOR2_X1 U9473 ( .A(n7592), .B(n7591), .Z(n7597) );
  AOI22_X1 U9474 ( .A1(n9155), .A2(n9429), .B1(n9177), .B2(n9431), .ZN(n7593)
         );
  NAND2_X1 U9475 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9463) );
  OAI211_X1 U9476 ( .C1(n10089), .C2(n9186), .A(n7593), .B(n9463), .ZN(n7594)
         );
  AOI21_X1 U9477 ( .B1(n9183), .B2(n7595), .A(n7594), .ZN(n7596) );
  OAI21_X1 U9478 ( .B1(n7597), .B2(n9170), .A(n7596), .ZN(P1_U3218) );
  INV_X1 U9479 ( .A(n7745), .ZN(n7737) );
  OAI22_X1 U9480 ( .A1(n8925), .A2(n7803), .B1(n7804), .B2(n10129), .ZN(n7600)
         );
  MUX2_X1 U9481 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7598), .S(n10145), .Z(n7599)
         );
  AOI211_X1 U9482 ( .C1(n7601), .C2(n7737), .A(n7600), .B(n7599), .ZN(n7602)
         );
  INV_X1 U9483 ( .A(n7602), .ZN(P2_U3226) );
  XOR2_X1 U9484 ( .A(n7604), .B(n7603), .Z(n7615) );
  OAI21_X1 U9485 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n7605), .A(n7558), .ZN(
        n7613) );
  INV_X1 U9486 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10337) );
  NAND2_X1 U9487 ( .A1(n8764), .A2(n7606), .ZN(n7607) );
  NAND2_X1 U9488 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8053) );
  OAI211_X1 U9489 ( .C1(n10337), .C2(n8088), .A(n7607), .B(n8053), .ZN(n7612)
         );
  AOI21_X1 U9490 ( .B1(n7629), .B2(n7609), .A(n7608), .ZN(n7610) );
  NOR2_X1 U9491 ( .A1(n7610), .A2(n8856), .ZN(n7611) );
  AOI211_X1 U9492 ( .C1(n8853), .C2(n7613), .A(n7612), .B(n7611), .ZN(n7614)
         );
  OAI21_X1 U9493 ( .B1(n7615), .B2(n8850), .A(n7614), .ZN(P2_U3191) );
  OAI21_X1 U9494 ( .B1(n7618), .B2(n7617), .A(n7616), .ZN(n7622) );
  XNOR2_X1 U9495 ( .A(n7620), .B(n7619), .ZN(n7621) );
  XNOR2_X1 U9496 ( .A(n7622), .B(n7621), .ZN(n7626) );
  NAND2_X1 U9497 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9493) );
  OAI21_X1 U9498 ( .B1(n8264), .B2(n7647), .A(n9493), .ZN(n7623) );
  AOI21_X1 U9499 ( .B1(n9155), .B2(n9426), .A(n7623), .ZN(n7625) );
  AOI22_X1 U9500 ( .A1(n9183), .A2(n7826), .B1(n9168), .B2(n9199), .ZN(n7624)
         );
  OAI211_X1 U9501 ( .C1(n7626), .C2(n9170), .A(n7625), .B(n7624), .ZN(P1_U3239) );
  INV_X1 U9502 ( .A(n7627), .ZN(n8059) );
  MUX2_X1 U9503 ( .A(n7629), .B(n7628), .S(n10199), .Z(n7630) );
  OAI21_X1 U9504 ( .B1(n8059), .B2(n8991), .A(n7630), .ZN(P2_U3468) );
  INV_X1 U9505 ( .A(n7631), .ZN(n7634) );
  NOR2_X1 U9506 ( .A1(n9986), .A2(n7632), .ZN(n7633) );
  NAND2_X1 U9507 ( .A1(n7634), .A2(n7633), .ZN(n7641) );
  OR2_X1 U9508 ( .A1(n7636), .A2(n6665), .ZN(n7843) );
  AND2_X1 U9509 ( .A1(n7637), .A2(n7843), .ZN(n7638) );
  NAND2_X1 U9510 ( .A1(n7639), .A2(n9284), .ZN(n7894) );
  OAI21_X1 U9511 ( .B1(n7639), .B2(n9284), .A(n7894), .ZN(n10098) );
  OR2_X1 U9512 ( .A1(n7652), .A2(n9414), .ZN(n7640) );
  OAI211_X1 U9513 ( .C1(n4658), .C2(n10095), .A(n9894), .B(n7897), .ZN(n10094)
         );
  INV_X1 U9514 ( .A(n10094), .ZN(n7642) );
  AOI22_X1 U9515 ( .A1(n9841), .A2(n7642), .B1(n9135), .B2(n9842), .ZN(n7643)
         );
  OAI21_X1 U9516 ( .B1(n10095), .B2(n10081), .A(n7643), .ZN(n7649) );
  XNOR2_X1 U9517 ( .A(n7644), .B(n9284), .ZN(n7645) );
  OAI222_X1 U9518 ( .A1(n9802), .A2(n7647), .B1(n9800), .B2(n7646), .C1(n9797), 
        .C2(n7645), .ZN(n10096) );
  MUX2_X1 U9519 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10096), .S(n9848), .Z(n7648)
         );
  AOI211_X1 U9520 ( .C1(n9700), .C2(n10098), .A(n7649), .B(n7648), .ZN(n7650)
         );
  INV_X1 U9521 ( .A(n7650), .ZN(P1_U3289) );
  NOR2_X1 U9522 ( .A1(n10075), .A2(n9864), .ZN(n9756) );
  OAI21_X1 U9523 ( .B1(n9819), .B2(n9756), .A(n7651), .ZN(n7660) );
  INV_X1 U9524 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7657) );
  NAND3_X1 U9525 ( .A1(n7654), .A2(n7653), .A3(n7652), .ZN(n7656) );
  OAI211_X1 U9526 ( .C1(n10072), .C2(n7657), .A(n7656), .B(n7655), .ZN(n7658)
         );
  NAND2_X1 U9527 ( .A1(n9848), .A2(n7658), .ZN(n7659) );
  OAI211_X1 U9528 ( .C1(n7661), .C2(n9848), .A(n7660), .B(n7659), .ZN(P1_U3293) );
  OAI21_X1 U9529 ( .B1(n7663), .B2(n9282), .A(n7662), .ZN(n10092) );
  INV_X1 U9530 ( .A(n10092), .ZN(n7675) );
  XNOR2_X1 U9531 ( .A(n7664), .B(n9282), .ZN(n7665) );
  OAI222_X1 U9532 ( .A1(n9800), .A2(n9364), .B1(n9802), .B2(n7666), .C1(n9797), 
        .C2(n7665), .ZN(n10090) );
  INV_X1 U9533 ( .A(n10090), .ZN(n7667) );
  MUX2_X1 U9534 ( .A(n7668), .B(n7667), .S(n9848), .Z(n7674) );
  OAI211_X1 U9535 ( .C1(n7670), .C2(n10089), .A(n9894), .B(n7669), .ZN(n10088)
         );
  OAI22_X1 U9536 ( .A1(n10075), .A2(n10088), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10072), .ZN(n7671) );
  AOI21_X1 U9537 ( .B1(n9819), .B2(n7672), .A(n7671), .ZN(n7673) );
  OAI211_X1 U9538 ( .C1(n7675), .C2(n9850), .A(n7674), .B(n7673), .ZN(P1_U3290) );
  INV_X1 U9539 ( .A(n7676), .ZN(n7679) );
  OAI222_X1 U9540 ( .A1(n9062), .A2(n7678), .B1(n9063), .B2(n7679), .C1(
        P2_U3151), .C2(n7677), .ZN(P2_U3276) );
  OAI222_X1 U9541 ( .A1(n10002), .A2(n7680), .B1(n8589), .B2(n7679), .C1(n6665), .C2(P1_U3086), .ZN(P1_U3336) );
  INV_X1 U9542 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9925) );
  INV_X1 U9543 ( .A(n9527), .ZN(n7683) );
  XNOR2_X1 U9544 ( .A(n7683), .B(n9533), .ZN(n9526) );
  XNOR2_X1 U9545 ( .A(n9526), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n7690) );
  INV_X1 U9546 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10036) );
  OAI211_X1 U9547 ( .C1(P1_REG2_REG_15__SCAN_IN), .C2(n7686), .A(n10052), .B(
        n9538), .ZN(n7687) );
  NAND2_X1 U9548 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9178) );
  OAI211_X1 U9549 ( .C1(n9596), .C2(n10036), .A(n7687), .B(n9178), .ZN(n7688)
         );
  AOI21_X1 U9550 ( .B1(n9533), .B2(n10054), .A(n7688), .ZN(n7689) );
  OAI21_X1 U9551 ( .B1(n7690), .B2(n9561), .A(n7689), .ZN(P1_U3258) );
  NAND2_X1 U9552 ( .A1(n8727), .A2(n7691), .ZN(n7695) );
  INV_X1 U9553 ( .A(n7692), .ZN(n7693) );
  AOI21_X1 U9554 ( .B1(n8722), .B2(n8752), .A(n7693), .ZN(n7694) );
  OAI211_X1 U9555 ( .C1(n7696), .C2(n8724), .A(n7695), .B(n7694), .ZN(n7701)
         );
  AOI211_X1 U9556 ( .C1(n7699), .C2(n7698), .A(n8717), .B(n7697), .ZN(n7700)
         );
  AOI211_X1 U9557 ( .C1(n7702), .C2(n8711), .A(n7701), .B(n7700), .ZN(n7703)
         );
  INV_X1 U9558 ( .A(n7703), .ZN(P2_U3179) );
  INV_X1 U9559 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7712) );
  XNOR2_X1 U9560 ( .A(n5839), .B(n8747), .ZN(n8290) );
  XNOR2_X1 U9561 ( .A(n7704), .B(n8290), .ZN(n7746) );
  INV_X1 U9562 ( .A(n7746), .ZN(n7711) );
  NAND2_X1 U9563 ( .A1(n7518), .A2(n7705), .ZN(n7707) );
  NAND2_X1 U9564 ( .A1(n7707), .A2(n7706), .ZN(n7720) );
  XNOR2_X1 U9565 ( .A(n7720), .B(n8290), .ZN(n7708) );
  NAND2_X1 U9566 ( .A1(n7708), .A2(n10136), .ZN(n7710) );
  AOI22_X1 U9567 ( .A1(n10132), .A2(n8748), .B1(n10131), .B2(n8746), .ZN(n7709) );
  OAI211_X1 U9568 ( .C1(n7746), .C2(n10141), .A(n7710), .B(n7709), .ZN(n7740)
         );
  AOI21_X1 U9569 ( .B1(n10165), .B2(n7711), .A(n7740), .ZN(n7714) );
  MUX2_X1 U9570 ( .A(n7712), .B(n7714), .S(n10184), .Z(n7713) );
  OAI21_X1 U9571 ( .B1(n8197), .B2(n9044), .A(n7713), .ZN(P2_U3420) );
  MUX2_X1 U9572 ( .A(n7715), .B(n7714), .S(n10199), .Z(n7716) );
  OAI21_X1 U9573 ( .B1(n8197), .B2(n8991), .A(n7716), .ZN(P2_U3469) );
  XNOR2_X1 U9574 ( .A(n7717), .B(n7721), .ZN(n7733) );
  INV_X1 U9575 ( .A(n6108), .ZN(n7718) );
  AOI21_X1 U9576 ( .B1(n7720), .B2(n7719), .A(n7718), .ZN(n7722) );
  XNOR2_X1 U9577 ( .A(n7722), .B(n7721), .ZN(n7723) );
  AOI222_X1 U9578 ( .A1(n10136), .A2(n7723), .B1(n8745), .B2(n10131), .C1(
        n8747), .C2(n10132), .ZN(n7729) );
  MUX2_X1 U9579 ( .A(n7724), .B(n7729), .S(n10184), .Z(n7726) );
  NAND2_X1 U9580 ( .A1(n6113), .A2(n6375), .ZN(n7725) );
  OAI211_X1 U9581 ( .C1(n7733), .C2(n9039), .A(n7726), .B(n7725), .ZN(P2_U3423) );
  MUX2_X1 U9582 ( .A(n8090), .B(n7729), .S(n10199), .Z(n7728) );
  NAND2_X1 U9583 ( .A1(n6113), .A2(n8983), .ZN(n7727) );
  OAI211_X1 U9584 ( .C1(n8986), .C2(n7733), .A(n7728), .B(n7727), .ZN(P2_U3470) );
  MUX2_X1 U9585 ( .A(n4919), .B(n7729), .S(n10145), .Z(n7732) );
  AOI22_X1 U9586 ( .A1(n6113), .A2(n8955), .B1(n8954), .B2(n7730), .ZN(n7731)
         );
  OAI211_X1 U9587 ( .C1(n7733), .C2(n8958), .A(n7732), .B(n7731), .ZN(P2_U3222) );
  OAI22_X1 U9588 ( .A1(n8059), .A2(n8925), .B1(n8054), .B2(n10129), .ZN(n7736)
         );
  MUX2_X1 U9589 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7734), .S(n10145), .Z(n7735)
         );
  AOI211_X1 U9590 ( .C1(n7738), .C2(n7737), .A(n7736), .B(n7735), .ZN(n7739)
         );
  INV_X1 U9591 ( .A(n7739), .ZN(P2_U3224) );
  MUX2_X1 U9592 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n7740), .S(n10145), .Z(n7741) );
  INV_X1 U9593 ( .A(n7741), .ZN(n7744) );
  INV_X1 U9594 ( .A(n7742), .ZN(n8194) );
  AOI22_X1 U9595 ( .A1(n5839), .A2(n8955), .B1(n8954), .B2(n8194), .ZN(n7743)
         );
  OAI211_X1 U9596 ( .C1(n7746), .C2(n7745), .A(n7744), .B(n7743), .ZN(P2_U3223) );
  NAND2_X1 U9597 ( .A1(n7822), .A2(n7821), .ZN(n7820) );
  NAND2_X1 U9598 ( .A1(n7820), .A2(n7747), .ZN(n7749) );
  OAI21_X1 U9599 ( .B1(n7749), .B2(n9201), .A(n7748), .ZN(n7917) );
  OAI211_X1 U9600 ( .C1(n7823), .C2(n7751), .A(n9894), .B(n7750), .ZN(n7913)
         );
  INV_X1 U9601 ( .A(n7913), .ZN(n7756) );
  NAND2_X1 U9602 ( .A1(n9372), .A2(n9197), .ZN(n7752) );
  NOR2_X1 U9603 ( .A1(n7752), .A2(n9201), .ZN(n7991) );
  AOI21_X1 U9604 ( .B1(n9201), .B2(n7752), .A(n7991), .ZN(n7755) );
  AOI22_X1 U9605 ( .A1(n9836), .A2(n9427), .B1(n4580), .B2(n9834), .ZN(n7754)
         );
  NAND2_X1 U9606 ( .A1(n7917), .A2(n7842), .ZN(n7753) );
  OAI211_X1 U9607 ( .C1(n7755), .C2(n9797), .A(n7754), .B(n7753), .ZN(n7914)
         );
  AOI211_X1 U9608 ( .C1(n7757), .C2(n7917), .A(n7756), .B(n7914), .ZN(n7760)
         );
  AOI22_X1 U9609 ( .A1(n9884), .A2(n7911), .B1(n10120), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7758) );
  OAI21_X1 U9610 ( .B1(n7760), .B2(n10120), .A(n7758), .ZN(P1_U3529) );
  AOI22_X1 U9611 ( .A1(n9954), .A2(n7911), .B1(n10113), .B2(
        P1_REG0_REG_7__SCAN_IN), .ZN(n7759) );
  OAI21_X1 U9612 ( .B1(n7760), .B2(n10113), .A(n7759), .ZN(P1_U3474) );
  OAI21_X1 U9613 ( .B1(n4392), .B2(n8010), .A(n9894), .ZN(n7762) );
  NOR2_X1 U9614 ( .A1(n7762), .A2(n7761), .ZN(n8004) );
  OAI21_X1 U9615 ( .B1(n9372), .B2(n7764), .A(n7763), .ZN(n7765) );
  NOR2_X1 U9616 ( .A1(n7765), .A2(n9278), .ZN(n7837) );
  AOI21_X1 U9617 ( .B1(n9278), .B2(n7765), .A(n7837), .ZN(n7766) );
  OAI222_X1 U9618 ( .A1(n9802), .A2(n7981), .B1(n9800), .B2(n7997), .C1(n9797), 
        .C2(n7766), .ZN(n8003) );
  AOI21_X1 U9619 ( .B1(n8004), .B2(n6665), .A(n8003), .ZN(n7774) );
  INV_X1 U9620 ( .A(n7984), .ZN(n7767) );
  OAI22_X1 U9621 ( .A1(n9848), .A2(n7060), .B1(n7767), .B2(n10072), .ZN(n7768)
         );
  AOI21_X1 U9622 ( .B1(n9819), .B2(n7769), .A(n7768), .ZN(n7773) );
  OAI21_X1 U9623 ( .B1(n7771), .B2(n9278), .A(n7770), .ZN(n8005) );
  NAND2_X1 U9624 ( .A1(n8005), .A2(n9700), .ZN(n7772) );
  OAI211_X1 U9625 ( .C1(n7774), .C2(n10077), .A(n7773), .B(n7772), .ZN(
        P1_U3283) );
  NAND2_X1 U9626 ( .A1(n7775), .A2(n7776), .ZN(n7877) );
  XNOR2_X1 U9627 ( .A(n7877), .B(n7878), .ZN(n7778) );
  NOR2_X1 U9628 ( .A1(n7778), .A2(n7777), .ZN(n7876) );
  AOI21_X1 U9629 ( .B1(n7778), .B2(n7777), .A(n7876), .ZN(n7784) );
  NAND2_X1 U9630 ( .A1(n9177), .A2(n9426), .ZN(n7780) );
  OAI211_X1 U9631 ( .C1(n9181), .C2(n7997), .A(n7780), .B(n7779), .ZN(n7781)
         );
  AOI21_X1 U9632 ( .B1(n8074), .B2(n9183), .A(n7781), .ZN(n7783) );
  NAND2_X1 U9633 ( .A1(n9168), .A2(n8075), .ZN(n7782) );
  OAI211_X1 U9634 ( .C1(n7784), .C2(n9170), .A(n7783), .B(n7782), .ZN(P1_U3221) );
  NAND2_X1 U9635 ( .A1(n7859), .A2(n9987), .ZN(n7786) );
  OAI211_X1 U9636 ( .C1(n7787), .C2(n9993), .A(n7786), .B(n7785), .ZN(P1_U3335) );
  OAI21_X1 U9637 ( .B1(n7991), .B2(n7788), .A(n9211), .ZN(n7789) );
  XNOR2_X1 U9638 ( .A(n7789), .B(n7793), .ZN(n7790) );
  AOI22_X1 U9639 ( .A1(n7790), .A2(n9829), .B1(n9836), .B2(n4580), .ZN(n7951)
         );
  MUX2_X1 U9640 ( .A(n7059), .B(n7951), .S(n9848), .Z(n7799) );
  NAND2_X1 U9641 ( .A1(n7988), .A2(n7994), .ZN(n7987) );
  NAND2_X1 U9642 ( .A1(n7987), .A2(n7791), .ZN(n7794) );
  OAI21_X1 U9643 ( .B1(n7794), .B2(n7793), .A(n7792), .ZN(n7954) );
  XOR2_X1 U9644 ( .A(n7875), .B(n7989), .Z(n7795) );
  AOI22_X1 U9645 ( .A1(n7795), .A2(n9894), .B1(n9834), .B2(n9424), .ZN(n7950)
         );
  AOI22_X1 U9646 ( .A1(n9819), .A2(n7875), .B1(n9842), .B2(n7890), .ZN(n7796)
         );
  OAI21_X1 U9647 ( .B1(n7950), .B2(n10075), .A(n7796), .ZN(n7797) );
  AOI21_X1 U9648 ( .B1(n7954), .B2(n9700), .A(n7797), .ZN(n7798) );
  NAND2_X1 U9649 ( .A1(n7799), .A2(n7798), .ZN(P1_U3284) );
  OAI21_X1 U9650 ( .B1(n7802), .B2(n7801), .A(n7800), .ZN(n7813) );
  NOR2_X1 U9651 ( .A1(n8731), .A2(n7803), .ZN(n7812) );
  INV_X1 U9652 ( .A(n7804), .ZN(n7805) );
  NAND2_X1 U9653 ( .A1(n8727), .A2(n7805), .ZN(n7809) );
  INV_X1 U9654 ( .A(n7806), .ZN(n7807) );
  AOI21_X1 U9655 ( .B1(n8722), .B2(n8751), .A(n7807), .ZN(n7808) );
  OAI211_X1 U9656 ( .C1(n7810), .C2(n8724), .A(n7809), .B(n7808), .ZN(n7811)
         );
  AOI211_X1 U9657 ( .C1(n7813), .C2(n8679), .A(n7812), .B(n7811), .ZN(n7814)
         );
  INV_X1 U9658 ( .A(n7814), .ZN(P2_U3153) );
  INV_X1 U9659 ( .A(n7821), .ZN(n7816) );
  XNOR2_X1 U9660 ( .A(n7815), .B(n7816), .ZN(n7817) );
  NAND2_X1 U9661 ( .A1(n7817), .A2(n9829), .ZN(n7819) );
  AOI22_X1 U9662 ( .A1(n9836), .A2(n9428), .B1(n9426), .B2(n9834), .ZN(n7818)
         );
  NAND2_X1 U9663 ( .A1(n7819), .A2(n7818), .ZN(n10109) );
  INV_X1 U9664 ( .A(n10109), .ZN(n7833) );
  OAI21_X1 U9665 ( .B1(n7822), .B2(n7821), .A(n7820), .ZN(n10111) );
  INV_X1 U9666 ( .A(n7898), .ZN(n7825) );
  INV_X1 U9667 ( .A(n7823), .ZN(n7824) );
  OAI211_X1 U9668 ( .C1(n10108), .C2(n7825), .A(n7824), .B(n9894), .ZN(n10106)
         );
  INV_X1 U9669 ( .A(n7826), .ZN(n7827) );
  OAI22_X1 U9670 ( .A1(n9848), .A2(n7828), .B1(n7827), .B2(n10072), .ZN(n7829)
         );
  AOI21_X1 U9671 ( .B1(n9819), .B2(n9199), .A(n7829), .ZN(n7830) );
  OAI21_X1 U9672 ( .B1(n10075), .B2(n10106), .A(n7830), .ZN(n7831) );
  AOI21_X1 U9673 ( .B1(n10111), .B2(n9700), .A(n7831), .ZN(n7832) );
  OAI21_X1 U9674 ( .B1(n7833), .B2(n10077), .A(n7832), .ZN(P1_U3287) );
  XNOR2_X1 U9675 ( .A(n7834), .B(n7835), .ZN(n9928) );
  INV_X1 U9676 ( .A(n9220), .ZN(n7836) );
  OAI21_X1 U9677 ( .B1(n7837), .B2(n7836), .A(n7835), .ZN(n7838) );
  AND3_X1 U9678 ( .A1(n7839), .A2(n7838), .A3(n9829), .ZN(n7841) );
  OAI22_X1 U9679 ( .A1(n9802), .A2(n9422), .B1(n7888), .B2(n9800), .ZN(n7840)
         );
  AOI211_X1 U9680 ( .C1(n9928), .C2(n7842), .A(n7841), .B(n7840), .ZN(n9932)
         );
  NOR2_X1 U9681 ( .A1(n10077), .A2(n7843), .ZN(n10071) );
  INV_X1 U9682 ( .A(n7761), .ZN(n7845) );
  INV_X1 U9683 ( .A(n7844), .ZN(n7937) );
  AOI211_X1 U9684 ( .C1(n6484), .C2(n7845), .A(n9864), .B(n7937), .ZN(n9929)
         );
  NAND2_X1 U9685 ( .A1(n9929), .A2(n9841), .ZN(n7847) );
  AOI22_X1 U9686 ( .A1(n10077), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8067), .B2(
        n9842), .ZN(n7846) );
  OAI211_X1 U9687 ( .C1(n7848), .C2(n10081), .A(n7847), .B(n7846), .ZN(n7849)
         );
  AOI21_X1 U9688 ( .B1(n9928), .B2(n10071), .A(n7849), .ZN(n7850) );
  OAI21_X1 U9689 ( .B1(n9932), .B2(n10077), .A(n7850), .ZN(P1_U3282) );
  INV_X1 U9690 ( .A(n7851), .ZN(n7858) );
  NAND2_X1 U9691 ( .A1(n9819), .A2(n9363), .ZN(n7854) );
  AOI22_X1 U9692 ( .A1(n9841), .A2(n7852), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9842), .ZN(n7853) );
  OAI211_X1 U9693 ( .C1(n7047), .C2(n9848), .A(n7854), .B(n7853), .ZN(n7855)
         );
  AOI21_X1 U9694 ( .B1(n9700), .B2(n7856), .A(n7855), .ZN(n7857) );
  OAI21_X1 U9695 ( .B1(n10077), .B2(n7858), .A(n7857), .ZN(P1_U3291) );
  INV_X1 U9696 ( .A(n7859), .ZN(n7860) );
  OAI222_X1 U9697 ( .A1(n9062), .A2(n7861), .B1(n9063), .B2(n7860), .C1(n8479), 
        .C2(P2_U3151), .ZN(P2_U3275) );
  XNOR2_X1 U9698 ( .A(n7862), .B(n8399), .ZN(n7874) );
  XNOR2_X1 U9699 ( .A(n7863), .B(n8399), .ZN(n7864) );
  AOI222_X1 U9700 ( .A1(n10136), .A2(n7864), .B1(n6118), .B2(n10131), .C1(
        n8746), .C2(n10132), .ZN(n7871) );
  MUX2_X1 U9701 ( .A(n7865), .B(n7871), .S(n10184), .Z(n7867) );
  NAND2_X1 U9702 ( .A1(n8185), .A2(n6375), .ZN(n7866) );
  OAI211_X1 U9703 ( .C1(n7874), .C2(n9039), .A(n7867), .B(n7866), .ZN(P2_U3426) );
  MUX2_X1 U9704 ( .A(n7868), .B(n7871), .S(n10199), .Z(n7870) );
  NAND2_X1 U9705 ( .A1(n8185), .A2(n8983), .ZN(n7869) );
  OAI211_X1 U9706 ( .C1(n7874), .C2(n8986), .A(n7870), .B(n7869), .ZN(P2_U3471) );
  MUX2_X1 U9707 ( .A(n10223), .B(n7871), .S(n10145), .Z(n7873) );
  AOI22_X1 U9708 ( .A1(n8185), .A2(n8955), .B1(n8954), .B2(n8184), .ZN(n7872)
         );
  OAI211_X1 U9709 ( .C1(n7874), .C2(n8958), .A(n7873), .B(n7872), .ZN(P2_U3221) );
  INV_X1 U9710 ( .A(n7875), .ZN(n7952) );
  AOI21_X1 U9711 ( .B1(n7878), .B2(n7877), .A(n7876), .ZN(n7885) );
  NAND2_X1 U9712 ( .A1(n7880), .A2(n7879), .ZN(n7882) );
  NAND2_X1 U9713 ( .A1(n7882), .A2(n7881), .ZN(n7883) );
  OAI211_X1 U9714 ( .C1(n7885), .C2(n7884), .A(n9175), .B(n7883), .ZN(n7892)
         );
  NAND2_X1 U9715 ( .A1(n9177), .A2(n4580), .ZN(n7887) );
  OAI211_X1 U9716 ( .C1(n9181), .C2(n7888), .A(n7887), .B(n7886), .ZN(n7889)
         );
  AOI21_X1 U9717 ( .B1(n7890), .B2(n9183), .A(n7889), .ZN(n7891) );
  OAI211_X1 U9718 ( .C1(n7952), .C2(n9186), .A(n7892), .B(n7891), .ZN(P1_U3231) );
  NAND2_X1 U9719 ( .A1(n7894), .A2(n7893), .ZN(n7896) );
  OAI21_X1 U9720 ( .B1(n7896), .B2(n9281), .A(n7895), .ZN(n10104) );
  OAI211_X1 U9721 ( .C1(n4657), .C2(n10101), .A(n9894), .B(n7898), .ZN(n10100)
         );
  AOI22_X1 U9722 ( .A1(n9819), .A2(n7900), .B1(n9842), .B2(n7899), .ZN(n7901)
         );
  OAI21_X1 U9723 ( .B1(n10075), .B2(n10100), .A(n7901), .ZN(n7908) );
  NAND2_X1 U9724 ( .A1(n7904), .A2(n9829), .ZN(n7906) );
  AOI22_X1 U9725 ( .A1(n9834), .A2(n9427), .B1(n9836), .B2(n9429), .ZN(n7905)
         );
  NAND2_X1 U9726 ( .A1(n7906), .A2(n7905), .ZN(n10102) );
  MUX2_X1 U9727 ( .A(n10102), .B(P1_REG2_REG_5__SCAN_IN), .S(n10077), .Z(n7907) );
  AOI211_X1 U9728 ( .C1(n9700), .C2(n10104), .A(n7908), .B(n7907), .ZN(n7909)
         );
  INV_X1 U9729 ( .A(n7909), .ZN(P1_U3288) );
  AOI22_X1 U9730 ( .A1(n9819), .A2(n7911), .B1(n9842), .B2(n7910), .ZN(n7912)
         );
  OAI21_X1 U9731 ( .B1(n10075), .B2(n7913), .A(n7912), .ZN(n7916) );
  MUX2_X1 U9732 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7914), .S(n9848), .Z(n7915)
         );
  AOI211_X1 U9733 ( .C1(n10071), .C2(n7917), .A(n7916), .B(n7915), .ZN(n7918)
         );
  INV_X1 U9734 ( .A(n7918), .ZN(P1_U3286) );
  XOR2_X1 U9735 ( .A(n7920), .B(n7919), .Z(n7929) );
  NAND2_X1 U9736 ( .A1(n8722), .A2(n8750), .ZN(n7922) );
  OAI211_X1 U9737 ( .C1(n7923), .C2(n8724), .A(n7922), .B(n7921), .ZN(n7926)
         );
  INV_X1 U9738 ( .A(n8727), .ZN(n8696) );
  NOR2_X1 U9739 ( .A1(n8696), .A2(n7924), .ZN(n7925) );
  AOI211_X1 U9740 ( .C1(n7927), .C2(n8711), .A(n7926), .B(n7925), .ZN(n7928)
         );
  OAI21_X1 U9741 ( .B1(n7929), .B2(n8717), .A(n7928), .ZN(P2_U3161) );
  OAI21_X1 U9742 ( .B1(n7931), .B2(n9295), .A(n7930), .ZN(n7949) );
  OAI21_X1 U9743 ( .B1(n7932), .B2(n7934), .A(n7933), .ZN(n7935) );
  INV_X1 U9744 ( .A(n7981), .ZN(n9423) );
  AOI222_X1 U9745 ( .A1(n9829), .A2(n7935), .B1(n9423), .B2(n9836), .C1(n9835), 
        .C2(n9834), .ZN(n7943) );
  OAI211_X1 U9746 ( .C1(n7937), .C2(n8045), .A(n9894), .B(n8102), .ZN(n7944)
         );
  OAI211_X1 U9747 ( .C1(n8045), .C2(n10107), .A(n7943), .B(n7944), .ZN(n7940)
         );
  NAND2_X1 U9748 ( .A1(n7940), .A2(n10123), .ZN(n7939) );
  NAND2_X1 U9749 ( .A1(n10120), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7938) );
  OAI211_X1 U9750 ( .C1(n7949), .C2(n9927), .A(n7939), .B(n7938), .ZN(P1_U3534) );
  NAND2_X1 U9751 ( .A1(n7940), .A2(n10115), .ZN(n7942) );
  NAND2_X1 U9752 ( .A1(n10113), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7941) );
  OAI211_X1 U9753 ( .C1(n7949), .C2(n9980), .A(n7942), .B(n7941), .ZN(P1_U3489) );
  OAI21_X1 U9754 ( .B1(n9677), .B2(n7944), .A(n7943), .ZN(n7947) );
  AOI22_X1 U9755 ( .A1(n10077), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8048), .B2(
        n9842), .ZN(n7945) );
  OAI21_X1 U9756 ( .B1(n8045), .B2(n10081), .A(n7945), .ZN(n7946) );
  AOI21_X1 U9757 ( .B1(n7947), .B2(n9848), .A(n7946), .ZN(n7948) );
  OAI21_X1 U9758 ( .B1(n7949), .B2(n9850), .A(n7948), .ZN(P1_U3281) );
  OAI211_X1 U9759 ( .C1(n7952), .C2(n10107), .A(n7951), .B(n7950), .ZN(n7953)
         );
  AOI21_X1 U9760 ( .B1(n10112), .B2(n7954), .A(n7953), .ZN(n7957) );
  NAND2_X1 U9761 ( .A1(n10120), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7955) );
  OAI21_X1 U9762 ( .B1(n7957), .B2(n10120), .A(n7955), .ZN(P1_U3531) );
  NAND2_X1 U9763 ( .A1(n10113), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7956) );
  OAI21_X1 U9764 ( .B1(n7957), .B2(n10113), .A(n7956), .ZN(P1_U3480) );
  XOR2_X1 U9765 ( .A(n7959), .B(n7958), .Z(n7973) );
  INV_X1 U9766 ( .A(n7960), .ZN(n7965) );
  NOR3_X1 U9767 ( .A1(n7961), .A2(n7963), .A3(n7962), .ZN(n7964) );
  OAI21_X1 U9768 ( .B1(n7965), .B2(n7964), .A(n8825), .ZN(n7972) );
  NAND2_X1 U9769 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8181) );
  OAI21_X1 U9770 ( .B1(n8846), .B2(n6314), .A(n8181), .ZN(n7970) );
  NAND3_X1 U9771 ( .A1(n8085), .A2(n4412), .A3(n7966), .ZN(n7967) );
  AOI21_X1 U9772 ( .B1(n7968), .B2(n7967), .A(n8835), .ZN(n7969) );
  AOI211_X1 U9773 ( .C1(n8848), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n7970), .B(
        n7969), .ZN(n7971) );
  OAI211_X1 U9774 ( .C1(n7973), .C2(n8850), .A(n7972), .B(n7971), .ZN(P2_U3194) );
  INV_X1 U9775 ( .A(n7974), .ZN(n7976) );
  NAND2_X1 U9776 ( .A1(n7976), .A2(n7975), .ZN(n8062) );
  OAI21_X1 U9777 ( .B1(n7976), .B2(n7975), .A(n8062), .ZN(n7977) );
  NOR2_X1 U9778 ( .A1(n7977), .A2(n7978), .ZN(n8064) );
  AOI21_X1 U9779 ( .B1(n7978), .B2(n7977), .A(n8064), .ZN(n7986) );
  NAND2_X1 U9780 ( .A1(n9177), .A2(n9425), .ZN(n7980) );
  OAI211_X1 U9781 ( .C1(n9181), .C2(n7981), .A(n7980), .B(n7979), .ZN(n7983)
         );
  NOR2_X1 U9782 ( .A1(n8010), .A2(n9186), .ZN(n7982) );
  AOI211_X1 U9783 ( .C1(n9183), .C2(n7984), .A(n7983), .B(n7982), .ZN(n7985)
         );
  OAI21_X1 U9784 ( .B1(n7986), .B2(n9170), .A(n7985), .ZN(P1_U3217) );
  OAI21_X1 U9785 ( .B1(n7988), .B2(n7994), .A(n7987), .ZN(n8081) );
  INV_X1 U9786 ( .A(n7750), .ZN(n7990) );
  OAI211_X1 U9787 ( .C1(n7990), .C2(n5155), .A(n9894), .B(n7989), .ZN(n8077)
         );
  OAI21_X1 U9788 ( .B1(n5155), .B2(n10107), .A(n8077), .ZN(n7999) );
  INV_X1 U9789 ( .A(n7991), .ZN(n7993) );
  NAND2_X1 U9790 ( .A1(n7993), .A2(n7992), .ZN(n7995) );
  XNOR2_X1 U9791 ( .A(n7995), .B(n7994), .ZN(n7996) );
  OAI222_X1 U9792 ( .A1(n9800), .A2(n7998), .B1(n9802), .B2(n7997), .C1(n7996), 
        .C2(n9797), .ZN(n8078) );
  AOI211_X1 U9793 ( .C1(n10112), .C2(n8081), .A(n7999), .B(n8078), .ZN(n8002)
         );
  NAND2_X1 U9794 ( .A1(n10113), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8000) );
  OAI21_X1 U9795 ( .B1(n8002), .B2(n10113), .A(n8000), .ZN(P1_U3477) );
  NAND2_X1 U9796 ( .A1(n10120), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8001) );
  OAI21_X1 U9797 ( .B1(n8002), .B2(n10120), .A(n8001), .ZN(P1_U3530) );
  INV_X1 U9798 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10336) );
  AOI211_X1 U9799 ( .C1(n10112), .C2(n8005), .A(n8004), .B(n8003), .ZN(n8007)
         );
  MUX2_X1 U9800 ( .A(n10336), .B(n8007), .S(n10123), .Z(n8006) );
  OAI21_X1 U9801 ( .B1(n8010), .B2(n9921), .A(n8006), .ZN(P1_U3532) );
  INV_X1 U9802 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n8008) );
  MUX2_X1 U9803 ( .A(n8008), .B(n8007), .S(n10115), .Z(n8009) );
  OAI21_X1 U9804 ( .B1(n8010), .B2(n9975), .A(n8009), .ZN(P1_U3483) );
  XNOR2_X1 U9805 ( .A(n8011), .B(n8012), .ZN(n8112) );
  INV_X1 U9806 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8015) );
  XNOR2_X1 U9807 ( .A(n8013), .B(n8012), .ZN(n8014) );
  AOI222_X1 U9808 ( .A1(n10136), .A2(n8014), .B1(n8744), .B2(n10131), .C1(
        n8745), .C2(n10132), .ZN(n8109) );
  MUX2_X1 U9809 ( .A(n8015), .B(n8109), .S(n10184), .Z(n8018) );
  INV_X1 U9810 ( .A(n8016), .ZN(n8108) );
  NAND2_X1 U9811 ( .A1(n8016), .A2(n6375), .ZN(n8017) );
  OAI211_X1 U9812 ( .C1(n8112), .C2(n9039), .A(n8018), .B(n8017), .ZN(P2_U3429) );
  MUX2_X1 U9813 ( .A(n8780), .B(n8109), .S(n10199), .Z(n8020) );
  NAND2_X1 U9814 ( .A1(n8016), .A2(n8983), .ZN(n8019) );
  OAI211_X1 U9815 ( .C1(n8112), .C2(n8986), .A(n8020), .B(n8019), .ZN(P2_U3472) );
  AOI21_X1 U9816 ( .B1(n8022), .B2(n8407), .A(n10151), .ZN(n8026) );
  OAI22_X1 U9817 ( .A1(n8023), .A2(n4652), .B1(n8594), .B2(n8946), .ZN(n8024)
         );
  AOI21_X1 U9818 ( .B1(n8026), .B2(n8025), .A(n8024), .ZN(n8995) );
  INV_X1 U9819 ( .A(n8995), .ZN(n8029) );
  INV_X1 U9820 ( .A(n8597), .ZN(n8996) );
  INV_X1 U9821 ( .A(n8596), .ZN(n8027) );
  OAI22_X1 U9822 ( .A1(n8996), .A2(n10128), .B1(n8027), .B2(n10129), .ZN(n8028) );
  OAI21_X1 U9823 ( .B1(n8029), .B2(n8028), .A(n10145), .ZN(n8032) );
  NAND2_X1 U9824 ( .A1(n8030), .A2(n6123), .ZN(n8992) );
  NAND3_X1 U9825 ( .A1(n8993), .A2(n8992), .A3(n8927), .ZN(n8031) );
  OAI211_X1 U9826 ( .C1(n10145), .C2(n8033), .A(n8032), .B(n8031), .ZN(
        P2_U3219) );
  INV_X1 U9827 ( .A(n8034), .ZN(n8037) );
  OAI222_X1 U9828 ( .A1(n9062), .A2(n8035), .B1(n9063), .B2(n8037), .C1(
        P2_U3151), .C2(n8337), .ZN(P2_U3273) );
  OAI222_X1 U9829 ( .A1(n10002), .A2(n8038), .B1(n8589), .B2(n8037), .C1(
        P1_U3086), .C2(n8036), .ZN(P1_U3333) );
  INV_X1 U9830 ( .A(n8039), .ZN(n8574) );
  OAI222_X1 U9831 ( .A1(P1_U3086), .A2(n9366), .B1(n8589), .B2(n8574), .C1(
        n8040), .C2(n10002), .ZN(P1_U3334) );
  XOR2_X1 U9832 ( .A(n8042), .B(n8041), .Z(n8050) );
  NAND2_X1 U9833 ( .A1(n9177), .A2(n9423), .ZN(n8044) );
  OAI211_X1 U9834 ( .C1(n9181), .C2(n9227), .A(n8044), .B(n8043), .ZN(n8047)
         );
  NOR2_X1 U9835 ( .A1(n8045), .A2(n9186), .ZN(n8046) );
  AOI211_X1 U9836 ( .C1(n9183), .C2(n8048), .A(n8047), .B(n8046), .ZN(n8049)
         );
  OAI21_X1 U9837 ( .B1(n8050), .B2(n9170), .A(n8049), .ZN(P1_U3224) );
  OAI211_X1 U9838 ( .C1(n4402), .C2(n8052), .A(n8051), .B(n8679), .ZN(n8058)
         );
  OAI21_X1 U9839 ( .B1(n8724), .B2(n5836), .A(n8053), .ZN(n8056) );
  NOR2_X1 U9840 ( .A1(n8696), .A2(n8054), .ZN(n8055) );
  AOI211_X1 U9841 ( .C1(n8722), .C2(n8749), .A(n8056), .B(n8055), .ZN(n8057)
         );
  OAI211_X1 U9842 ( .C1(n8059), .C2(n8731), .A(n8058), .B(n8057), .ZN(P2_U3171) );
  NAND2_X1 U9843 ( .A1(n8061), .A2(n8060), .ZN(n8066) );
  INV_X1 U9844 ( .A(n8062), .ZN(n8063) );
  NOR2_X1 U9845 ( .A1(n8064), .A2(n8063), .ZN(n8065) );
  XOR2_X1 U9846 ( .A(n8066), .B(n8065), .Z(n8073) );
  NAND2_X1 U9847 ( .A1(n9183), .A2(n8067), .ZN(n8070) );
  AOI21_X1 U9848 ( .B1(n9177), .B2(n9424), .A(n8068), .ZN(n8069) );
  OAI211_X1 U9849 ( .C1(n9422), .C2(n9181), .A(n8070), .B(n8069), .ZN(n8071)
         );
  AOI21_X1 U9850 ( .B1(n9168), .B2(n6484), .A(n8071), .ZN(n8072) );
  OAI21_X1 U9851 ( .B1(n8073), .B2(n9170), .A(n8072), .ZN(P1_U3236) );
  AOI22_X1 U9852 ( .A1(n9819), .A2(n8075), .B1(n9842), .B2(n8074), .ZN(n8076)
         );
  OAI21_X1 U9853 ( .B1(n8077), .B2(n10075), .A(n8076), .ZN(n8080) );
  MUX2_X1 U9854 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n8078), .S(n9848), .Z(n8079)
         );
  AOI211_X1 U9855 ( .C1(n9700), .C2(n8081), .A(n8080), .B(n8079), .ZN(n8082)
         );
  INV_X1 U9856 ( .A(n8082), .ZN(P1_U3285) );
  XOR2_X1 U9857 ( .A(n8084), .B(n8083), .Z(n8096) );
  OAI21_X1 U9858 ( .B1(P2_REG2_REG_11__SCAN_IN), .B2(n4386), .A(n8085), .ZN(
        n8094) );
  INV_X1 U9859 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10027) );
  NAND2_X1 U9860 ( .A1(n8764), .A2(n8086), .ZN(n8087) );
  NAND2_X1 U9861 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8692) );
  OAI211_X1 U9862 ( .C1(n10027), .C2(n8088), .A(n8087), .B(n8692), .ZN(n8093)
         );
  AOI21_X1 U9863 ( .B1(n8090), .B2(n8089), .A(n7961), .ZN(n8091) );
  NOR2_X1 U9864 ( .A1(n8091), .A2(n8856), .ZN(n8092) );
  AOI211_X1 U9865 ( .C1(n8853), .C2(n8094), .A(n8093), .B(n8092), .ZN(n8095)
         );
  OAI21_X1 U9866 ( .B1(n8096), .B2(n8850), .A(n8095), .ZN(P2_U3193) );
  XOR2_X1 U9867 ( .A(n9296), .B(n8097), .Z(n8126) );
  XNOR2_X1 U9868 ( .A(n8098), .B(n9296), .ZN(n8101) );
  NAND2_X1 U9869 ( .A1(n9814), .A2(n9834), .ZN(n8099) );
  OAI21_X1 U9870 ( .B1(n9422), .B2(n9800), .A(n8099), .ZN(n8100) );
  AOI21_X1 U9871 ( .B1(n8101), .B2(n9829), .A(n8100), .ZN(n8120) );
  INV_X1 U9872 ( .A(n8120), .ZN(n8106) );
  INV_X1 U9873 ( .A(n9228), .ZN(n8265) );
  OAI211_X1 U9874 ( .C1(n7936), .C2(n8265), .A(n9894), .B(n9840), .ZN(n8119)
         );
  AOI22_X1 U9875 ( .A1(n10077), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8268), .B2(
        n9842), .ZN(n8104) );
  NAND2_X1 U9876 ( .A1(n9228), .A2(n9819), .ZN(n8103) );
  OAI211_X1 U9877 ( .C1(n8119), .C2(n10075), .A(n8104), .B(n8103), .ZN(n8105)
         );
  AOI21_X1 U9878 ( .B1(n8106), .B2(n9848), .A(n8105), .ZN(n8107) );
  OAI21_X1 U9879 ( .B1(n8126), .B2(n9850), .A(n8107), .ZN(P1_U3280) );
  NOR2_X1 U9880 ( .A1(n8108), .A2(n10128), .ZN(n8111) );
  INV_X1 U9881 ( .A(n8109), .ZN(n8110) );
  AOI211_X1 U9882 ( .C1(n8954), .C2(n8671), .A(n8111), .B(n8110), .ZN(n8115)
         );
  INV_X1 U9883 ( .A(n8112), .ZN(n8113) );
  AOI22_X1 U9884 ( .A1(n8113), .A2(n8927), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n10148), .ZN(n8114) );
  OAI21_X1 U9885 ( .B1(n8115), .B2(n10148), .A(n8114), .ZN(P2_U3220) );
  INV_X1 U9886 ( .A(n8127), .ZN(n8118) );
  NAND2_X1 U9887 ( .A1(n9058), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8117) );
  NAND2_X1 U9888 ( .A1(n8116), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8515) );
  OAI211_X1 U9889 ( .C1(n8118), .C2(n9063), .A(n8117), .B(n8515), .ZN(P2_U3272) );
  AOI22_X1 U9890 ( .A1(n9228), .A2(n9884), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n10120), .ZN(n8122) );
  NAND2_X1 U9891 ( .A1(n8120), .A2(n8119), .ZN(n8123) );
  NAND2_X1 U9892 ( .A1(n8123), .A2(n10123), .ZN(n8121) );
  OAI211_X1 U9893 ( .C1(n8126), .C2(n9927), .A(n8122), .B(n8121), .ZN(P1_U3535) );
  AOI22_X1 U9894 ( .A1(n9228), .A2(n9954), .B1(P1_REG0_REG_13__SCAN_IN), .B2(
        n10113), .ZN(n8125) );
  NAND2_X1 U9895 ( .A1(n8123), .A2(n10115), .ZN(n8124) );
  OAI211_X1 U9896 ( .C1(n8126), .C2(n9980), .A(n8125), .B(n8124), .ZN(P1_U3492) );
  NAND2_X1 U9897 ( .A1(n8127), .A2(n9987), .ZN(n8129) );
  OR2_X1 U9898 ( .A1(n8128), .A2(P1_U3086), .ZN(n9359) );
  OAI211_X1 U9899 ( .C1(n8130), .C2(n9993), .A(n8129), .B(n9359), .ZN(P1_U3332) );
  OAI211_X1 U9900 ( .C1(n8133), .C2(n8132), .A(n8131), .B(n9175), .ZN(n8138)
         );
  NAND2_X1 U9901 ( .A1(n9177), .A2(n9835), .ZN(n8135) );
  OAI211_X1 U9902 ( .C1(n9181), .C2(n9799), .A(n8135), .B(n8134), .ZN(n8136)
         );
  AOI21_X1 U9903 ( .B1(n9843), .B2(n9183), .A(n8136), .ZN(n8137) );
  OAI211_X1 U9904 ( .C1(n9846), .C2(n9186), .A(n8138), .B(n8137), .ZN(P1_U3215) );
  INV_X1 U9905 ( .A(n8139), .ZN(n8142) );
  OAI222_X1 U9906 ( .A1(P2_U3151), .A2(n5695), .B1(n9063), .B2(n8142), .C1(
        n8140), .C2(n9062), .ZN(P2_U3271) );
  OAI222_X1 U9907 ( .A1(n8143), .A2(P1_U3086), .B1(n8589), .B2(n8142), .C1(
        n8141), .C2(n10002), .ZN(P1_U3331) );
  XNOR2_X1 U9908 ( .A(n8716), .B(n8743), .ZN(n8412) );
  XNOR2_X1 U9909 ( .A(n8144), .B(n8412), .ZN(n8155) );
  INV_X1 U9910 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n10353) );
  XNOR2_X1 U9911 ( .A(n8145), .B(n8412), .ZN(n8146) );
  AOI222_X1 U9912 ( .A1(n10136), .A2(n8146), .B1(n8741), .B2(n10131), .C1(
        n8744), .C2(n10132), .ZN(n8152) );
  MUX2_X1 U9913 ( .A(n10353), .B(n8152), .S(n10184), .Z(n8148) );
  NAND2_X1 U9914 ( .A1(n8716), .A2(n6375), .ZN(n8147) );
  OAI211_X1 U9915 ( .C1(n8155), .C2(n9039), .A(n8148), .B(n8147), .ZN(P2_U3435) );
  MUX2_X1 U9916 ( .A(n8149), .B(n8152), .S(n10199), .Z(n8151) );
  NAND2_X1 U9917 ( .A1(n8716), .A2(n8983), .ZN(n8150) );
  OAI211_X1 U9918 ( .C1(n8986), .C2(n8155), .A(n8151), .B(n8150), .ZN(P2_U3474) );
  MUX2_X1 U9919 ( .A(n4915), .B(n8152), .S(n10145), .Z(n8154) );
  AOI22_X1 U9920 ( .A1(n8716), .A2(n8955), .B1(n8954), .B2(n8728), .ZN(n8153)
         );
  OAI211_X1 U9921 ( .C1(n8155), .C2(n8958), .A(n8154), .B(n8153), .ZN(P2_U3218) );
  XNOR2_X1 U9922 ( .A(n8156), .B(n8298), .ZN(n8170) );
  INV_X1 U9923 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8160) );
  XNOR2_X1 U9924 ( .A(n8157), .B(n8298), .ZN(n8159) );
  AOI222_X1 U9925 ( .A1(n10136), .A2(n8159), .B1(n8158), .B2(n10131), .C1(
        n8743), .C2(n10132), .ZN(n8166) );
  MUX2_X1 U9926 ( .A(n8160), .B(n8166), .S(n10184), .Z(n8162) );
  NAND2_X1 U9927 ( .A1(n8634), .A2(n6375), .ZN(n8161) );
  OAI211_X1 U9928 ( .C1(n8170), .C2(n9039), .A(n8162), .B(n8161), .ZN(P2_U3438) );
  MUX2_X1 U9929 ( .A(n8163), .B(n8166), .S(n10199), .Z(n8165) );
  NAND2_X1 U9930 ( .A1(n8634), .A2(n8983), .ZN(n8164) );
  OAI211_X1 U9931 ( .C1(n8170), .C2(n8986), .A(n8165), .B(n8164), .ZN(P2_U3475) );
  MUX2_X1 U9932 ( .A(n8167), .B(n8166), .S(n10145), .Z(n8169) );
  AOI22_X1 U9933 ( .A1(n8634), .A2(n8955), .B1(n8954), .B2(n8633), .ZN(n8168)
         );
  OAI211_X1 U9934 ( .C1(n8170), .C2(n8958), .A(n8169), .B(n8168), .ZN(P2_U3217) );
  INV_X1 U9935 ( .A(n8171), .ZN(n8175) );
  OAI222_X1 U9936 ( .A1(P2_U3151), .A2(n8173), .B1(n9063), .B2(n8175), .C1(
        n8172), .C2(n9062), .ZN(P2_U3270) );
  OAI222_X1 U9937 ( .A1(n8176), .A2(P1_U3086), .B1(n8589), .B2(n8175), .C1(
        n8174), .C2(n10002), .ZN(P1_U3330) );
  XNOR2_X1 U9938 ( .A(n8179), .B(n8178), .ZN(n8180) );
  XNOR2_X1 U9939 ( .A(n8177), .B(n8180), .ZN(n8188) );
  NAND2_X1 U9940 ( .A1(n8722), .A2(n8746), .ZN(n8182) );
  OAI211_X1 U9941 ( .C1(n8594), .C2(n8724), .A(n8182), .B(n8181), .ZN(n8183)
         );
  AOI21_X1 U9942 ( .B1(n8184), .B2(n8727), .A(n8183), .ZN(n8187) );
  NAND2_X1 U9943 ( .A1(n8185), .A2(n8711), .ZN(n8186) );
  OAI211_X1 U9944 ( .C1(n8188), .C2(n8717), .A(n8187), .B(n8186), .ZN(P2_U3164) );
  XNOR2_X1 U9945 ( .A(n8687), .B(n8747), .ZN(n8689) );
  XNOR2_X1 U9946 ( .A(n8689), .B(n8688), .ZN(n8189) );
  NAND2_X1 U9947 ( .A1(n8189), .A2(n8679), .ZN(n8196) );
  NAND2_X1 U9948 ( .A1(n8722), .A2(n8748), .ZN(n8191) );
  OAI211_X1 U9949 ( .C1(n8192), .C2(n8724), .A(n8191), .B(n8190), .ZN(n8193)
         );
  AOI21_X1 U9950 ( .B1(n8194), .B2(n8727), .A(n8193), .ZN(n8195) );
  OAI211_X1 U9951 ( .C1(n8197), .C2(n8731), .A(n8196), .B(n8195), .ZN(P2_U3157) );
  INV_X1 U9952 ( .A(n8198), .ZN(n8202) );
  OAI222_X1 U9953 ( .A1(n8200), .A2(P1_U3086), .B1(n8589), .B2(n8202), .C1(
        n8199), .C2(n10002), .ZN(P1_U3329) );
  OAI222_X1 U9954 ( .A1(P2_U3151), .A2(n8203), .B1(n9063), .B2(n8202), .C1(
        n8201), .C2(n9062), .ZN(P2_U3269) );
  INV_X1 U9955 ( .A(n8296), .ZN(n8415) );
  XNOR2_X1 U9956 ( .A(n8204), .B(n8415), .ZN(n8216) );
  INV_X1 U9957 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8207) );
  XNOR2_X1 U9958 ( .A(n8205), .B(n8415), .ZN(n8206) );
  AOI222_X1 U9959 ( .A1(n10136), .A2(n8206), .B1(n8740), .B2(n10131), .C1(
        n8741), .C2(n10132), .ZN(n8212) );
  MUX2_X1 U9960 ( .A(n8207), .B(n8212), .S(n10184), .Z(n8209) );
  NAND2_X1 U9961 ( .A1(n8644), .A2(n6375), .ZN(n8208) );
  OAI211_X1 U9962 ( .C1(n8216), .C2(n9039), .A(n8209), .B(n8208), .ZN(P2_U3441) );
  MUX2_X1 U9963 ( .A(n8840), .B(n8212), .S(n10199), .Z(n8211) );
  NAND2_X1 U9964 ( .A1(n8644), .A2(n8983), .ZN(n8210) );
  OAI211_X1 U9965 ( .C1(n8216), .C2(n8986), .A(n8211), .B(n8210), .ZN(P2_U3476) );
  MUX2_X1 U9966 ( .A(n8213), .B(n8212), .S(n10145), .Z(n8215) );
  AOI22_X1 U9967 ( .A1(n8644), .A2(n8955), .B1(n8954), .B2(n8643), .ZN(n8214)
         );
  OAI211_X1 U9968 ( .C1(n8216), .C2(n8958), .A(n8215), .B(n8214), .ZN(P2_U3216) );
  INV_X1 U9969 ( .A(n8221), .ZN(n8299) );
  XNOR2_X1 U9970 ( .A(n8217), .B(n8299), .ZN(n8220) );
  NAND2_X1 U9971 ( .A1(n8933), .A2(n10131), .ZN(n8218) );
  OAI21_X1 U9972 ( .B1(n8708), .B2(n8946), .A(n8218), .ZN(n8219) );
  AOI21_X1 U9973 ( .B1(n8220), .B2(n10136), .A(n8219), .ZN(n8989) );
  NAND2_X1 U9974 ( .A1(n8222), .A2(n8221), .ZN(n8223) );
  AND2_X1 U9975 ( .A1(n8224), .A2(n8223), .ZN(n8987) );
  INV_X1 U9976 ( .A(n8712), .ZN(n9045) );
  AOI22_X1 U9977 ( .A1(n10148), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8954), .B2(
        n8710), .ZN(n8225) );
  OAI21_X1 U9978 ( .B1(n9045), .B2(n8925), .A(n8225), .ZN(n8226) );
  AOI21_X1 U9979 ( .B1(n8987), .B2(n8927), .A(n8226), .ZN(n8227) );
  OAI21_X1 U9980 ( .B1(n8989), .B2(n10148), .A(n8227), .ZN(P2_U3215) );
  NAND2_X1 U9981 ( .A1(n8228), .A2(n8428), .ZN(n8229) );
  XNOR2_X1 U9982 ( .A(n8229), .B(n8230), .ZN(n8243) );
  INV_X1 U9983 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8233) );
  XNOR2_X1 U9984 ( .A(n8231), .B(n8230), .ZN(n8232) );
  AOI222_X1 U9985 ( .A1(n10136), .A2(n8232), .B1(n8910), .B2(n10131), .C1(
        n8739), .C2(n10132), .ZN(n8239) );
  MUX2_X1 U9986 ( .A(n8233), .B(n8239), .S(n10184), .Z(n8235) );
  NAND2_X1 U9987 ( .A1(n6132), .A2(n6375), .ZN(n8234) );
  OAI211_X1 U9988 ( .C1(n8243), .C2(n9039), .A(n8235), .B(n8234), .ZN(P2_U3448) );
  INV_X1 U9989 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8236) );
  MUX2_X1 U9990 ( .A(n8236), .B(n8239), .S(n10199), .Z(n8238) );
  NAND2_X1 U9991 ( .A1(n6132), .A2(n8983), .ZN(n8237) );
  OAI211_X1 U9992 ( .C1(n8986), .C2(n8243), .A(n8238), .B(n8237), .ZN(P2_U3480) );
  MUX2_X1 U9993 ( .A(n8240), .B(n8239), .S(n10145), .Z(n8242) );
  AOI22_X1 U9994 ( .A1(n6132), .A2(n8955), .B1(n8954), .B2(n8257), .ZN(n8241)
         );
  OAI211_X1 U9995 ( .C1(n8243), .C2(n8958), .A(n8242), .B(n8241), .ZN(P2_U3212) );
  OAI21_X1 U9996 ( .B1(n8610), .B2(n8247), .A(n8246), .ZN(n8248) );
  XNOR2_X1 U9997 ( .A(n8249), .B(n8739), .ZN(n8658) );
  AOI21_X1 U9998 ( .B1(n8253), .B2(n8252), .A(n8251), .ZN(n8678) );
  AOI22_X1 U9999 ( .A1(n8739), .A2(n8722), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8254) );
  OAI21_X1 U10000 ( .B1(n8255), .B2(n8724), .A(n8254), .ZN(n8256) );
  AOI21_X1 U10001 ( .B1(n8257), .B2(n8727), .A(n8256), .ZN(n8258) );
  OAI211_X1 U10002 ( .C1(n8260), .C2(n8731), .A(n8259), .B(n8258), .ZN(
        P2_U3163) );
  XOR2_X1 U10003 ( .A(n8262), .B(n8261), .Z(n8270) );
  NAND2_X1 U10004 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9515) );
  NAND2_X1 U10005 ( .A1(n9155), .A2(n9814), .ZN(n8263) );
  OAI211_X1 U10006 ( .C1(n8264), .C2(n9422), .A(n9515), .B(n8263), .ZN(n8267)
         );
  NOR2_X1 U10007 ( .A1(n8265), .A2(n9186), .ZN(n8266) );
  AOI211_X1 U10008 ( .C1(n9183), .C2(n8268), .A(n8267), .B(n8266), .ZN(n8269)
         );
  OAI21_X1 U10009 ( .B1(n8270), .B2(n9170), .A(n8269), .ZN(P1_U3234) );
  NAND2_X1 U10010 ( .A1(n9627), .A2(n9177), .ZN(n8274) );
  OAI21_X1 U10011 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n8275), .A(n8274), .ZN(
        n8277) );
  NOR2_X1 U10012 ( .A1(n10374), .A2(n9181), .ZN(n8276) );
  AOI211_X1 U10013 ( .C1(n9183), .C2(n9623), .A(n8277), .B(n8276), .ZN(n8278)
         );
  NOR2_X1 U10014 ( .A1(n9002), .A2(n8734), .ZN(n8480) );
  NAND2_X1 U10015 ( .A1(n8468), .A2(n4318), .ZN(n8879) );
  INV_X1 U10016 ( .A(n8281), .ZN(n8445) );
  INV_X1 U10017 ( .A(n10126), .ZN(n10135) );
  NAND4_X1 U10018 ( .A1(n8345), .A2(n10135), .A3(n10150), .A4(n6057), .ZN(
        n8283) );
  NOR2_X1 U10019 ( .A1(n8283), .A2(n8282), .ZN(n8286) );
  NAND4_X1 U10020 ( .A1(n8286), .A2(n8285), .A3(n8353), .A4(n8284), .ZN(n8287)
         );
  NOR3_X1 U10021 ( .A1(n8289), .A2(n8288), .A3(n8287), .ZN(n8291) );
  NAND4_X1 U10022 ( .A1(n8292), .A2(n8291), .A3(n8375), .A4(n8290), .ZN(n8293)
         );
  NOR2_X1 U10023 ( .A1(n4819), .A2(n8293), .ZN(n8294) );
  NAND3_X1 U10024 ( .A1(n8407), .A2(n8403), .A3(n8294), .ZN(n8295) );
  NOR2_X1 U10025 ( .A1(n8296), .A2(n8295), .ZN(n8297) );
  NAND4_X1 U10026 ( .A1(n8299), .A2(n8298), .A3(n8297), .A4(n8412), .ZN(n8300)
         );
  NOR2_X1 U10027 ( .A1(n8608), .A2(n8300), .ZN(n8301) );
  AND4_X1 U10028 ( .A1(n8302), .A2(n8921), .A3(n8909), .A4(n8301), .ZN(n8303)
         );
  NAND4_X1 U10029 ( .A1(n8887), .A2(n8304), .A3(n8903), .A4(n8303), .ZN(n8305)
         );
  NOR2_X1 U10030 ( .A1(n8879), .A2(n8305), .ZN(n8306) );
  INV_X1 U10031 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8315) );
  NAND2_X1 U10032 ( .A1(n8311), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8314) );
  NAND2_X1 U10033 ( .A1(n8312), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8313) );
  OAI211_X1 U10034 ( .C1(n8315), .C2(n4695), .A(n8314), .B(n8313), .ZN(n8316)
         );
  INV_X1 U10035 ( .A(n8316), .ZN(n8317) );
  NAND2_X1 U10036 ( .A1(n8999), .A2(n8733), .ZN(n8325) );
  NAND2_X1 U10037 ( .A1(n9002), .A2(n8859), .ZN(n8319) );
  INV_X1 U10038 ( .A(n8322), .ZN(n8323) );
  INV_X1 U10039 ( .A(n8325), .ZN(n8507) );
  NAND2_X1 U10040 ( .A1(n8326), .A2(n8499), .ZN(n8328) );
  AND2_X1 U10041 ( .A1(n8735), .A2(n8499), .ZN(n8327) );
  INV_X1 U10042 ( .A(n8329), .ZN(n8332) );
  NAND2_X1 U10043 ( .A1(n8419), .A2(n8330), .ZN(n8331) );
  MUX2_X1 U10044 ( .A(n8332), .B(n8331), .S(n8475), .Z(n8333) );
  INV_X1 U10045 ( .A(n8333), .ZN(n8414) );
  NAND3_X1 U10046 ( .A1(n10154), .A2(n8338), .A3(n8337), .ZN(n8339) );
  INV_X1 U10047 ( .A(n8342), .ZN(n8344) );
  NAND3_X1 U10048 ( .A1(n8345), .A2(n8344), .A3(n8343), .ZN(n8346) );
  NAND2_X1 U10049 ( .A1(n8362), .A2(n8347), .ZN(n8350) );
  NAND2_X1 U10050 ( .A1(n8354), .A2(n8348), .ZN(n8349) );
  MUX2_X1 U10051 ( .A(n8350), .B(n8349), .S(n8475), .Z(n8351) );
  INV_X1 U10052 ( .A(n8351), .ZN(n8352) );
  INV_X1 U10053 ( .A(n8354), .ZN(n8356) );
  OAI21_X1 U10054 ( .B1(n8361), .B2(n8356), .A(n8355), .ZN(n8359) );
  AND2_X1 U10055 ( .A1(n8366), .A2(n8364), .ZN(n8358) );
  AOI21_X1 U10056 ( .B1(n8359), .B2(n8358), .A(n8357), .ZN(n8360) );
  INV_X1 U10057 ( .A(n8365), .ZN(n8367) );
  NAND2_X1 U10058 ( .A1(n8367), .A2(n8366), .ZN(n8368) );
  AOI21_X1 U10059 ( .B1(n8371), .B2(n8370), .A(n8499), .ZN(n8372) );
  INV_X1 U10060 ( .A(n8372), .ZN(n8373) );
  NAND2_X1 U10061 ( .A1(n8374), .A2(n8373), .ZN(n8376) );
  AND2_X1 U10062 ( .A1(n8382), .A2(n8377), .ZN(n8380) );
  AND2_X1 U10063 ( .A1(n8384), .A2(n8378), .ZN(n8379) );
  MUX2_X1 U10064 ( .A(n8380), .B(n8379), .S(n8475), .Z(n8381) );
  AND2_X1 U10065 ( .A1(n8499), .A2(n8746), .ZN(n8389) );
  OAI21_X1 U10066 ( .B1(n8499), .B2(n8746), .A(n6113), .ZN(n8388) );
  OAI21_X1 U10067 ( .B1(n8389), .B2(n6113), .A(n8388), .ZN(n8390) );
  OAI21_X1 U10068 ( .B1(n8392), .B2(n8391), .A(n8390), .ZN(n8393) );
  INV_X1 U10069 ( .A(n8393), .ZN(n8398) );
  INV_X1 U10070 ( .A(n8394), .ZN(n8396) );
  OR2_X1 U10071 ( .A1(n8396), .A2(n8395), .ZN(n8397) );
  MUX2_X1 U10072 ( .A(n8401), .B(n8400), .S(n8499), .Z(n8402) );
  MUX2_X1 U10073 ( .A(n8406), .B(n8405), .S(n8499), .Z(n8408) );
  NAND2_X1 U10074 ( .A1(n8597), .A2(n8669), .ZN(n8409) );
  MUX2_X1 U10075 ( .A(n8410), .B(n8409), .S(n8475), .Z(n8411) );
  INV_X1 U10076 ( .A(n8417), .ZN(n8418) );
  INV_X1 U10077 ( .A(n8419), .ZN(n8420) );
  NAND2_X1 U10078 ( .A1(n8424), .A2(n8421), .ZN(n8423) );
  OAI21_X1 U10079 ( .B1(n8427), .B2(n8475), .A(n8426), .ZN(n8436) );
  INV_X1 U10080 ( .A(n8428), .ZN(n8435) );
  NAND2_X1 U10081 ( .A1(n8438), .A2(n8429), .ZN(n8432) );
  INV_X1 U10082 ( .A(n8430), .ZN(n8431) );
  MUX2_X1 U10083 ( .A(n8432), .B(n8431), .S(n8475), .Z(n8433) );
  INV_X1 U10084 ( .A(n8433), .ZN(n8434) );
  MUX2_X1 U10085 ( .A(n8438), .B(n8437), .S(n8499), .Z(n8439) );
  NAND2_X1 U10086 ( .A1(n8442), .A2(n4295), .ZN(n8443) );
  MUX2_X1 U10087 ( .A(n5089), .B(n8443), .S(n8475), .Z(n8444) );
  INV_X1 U10088 ( .A(n8444), .ZN(n8447) );
  NOR2_X1 U10089 ( .A1(n8738), .A2(n8475), .ZN(n8449) );
  NAND2_X1 U10090 ( .A1(n9021), .A2(n8449), .ZN(n8448) );
  OAI21_X1 U10091 ( .B1(n8911), .B2(n8475), .A(n8448), .ZN(n8453) );
  NAND2_X1 U10092 ( .A1(n8738), .A2(n8475), .ZN(n8454) );
  OAI21_X1 U10093 ( .B1(n8624), .B2(n8454), .A(n8456), .ZN(n8452) );
  INV_X1 U10094 ( .A(n8449), .ZN(n8450) );
  OAI21_X1 U10095 ( .B1(n8911), .B2(n8450), .A(n9021), .ZN(n8451) );
  AOI22_X1 U10096 ( .A1(n8457), .A2(n8453), .B1(n8452), .B2(n8451), .ZN(n8460)
         );
  INV_X1 U10097 ( .A(n8454), .ZN(n8455) );
  AOI22_X1 U10098 ( .A1(n8456), .A2(n8455), .B1(n8475), .B2(n8911), .ZN(n8458)
         );
  OR2_X1 U10099 ( .A1(n8458), .A2(n8457), .ZN(n8459) );
  MUX2_X1 U10100 ( .A(n8464), .B(n8463), .S(n8475), .Z(n8465) );
  INV_X1 U10101 ( .A(n8879), .ZN(n8466) );
  NAND2_X1 U10102 ( .A1(n8467), .A2(n8466), .ZN(n8470) );
  MUX2_X1 U10103 ( .A(n4318), .B(n8468), .S(n8499), .Z(n8469) );
  NAND2_X1 U10104 ( .A1(n8470), .A2(n5172), .ZN(n8474) );
  MUX2_X1 U10105 ( .A(n8472), .B(n8471), .S(n8475), .Z(n8473) );
  MUX2_X1 U10106 ( .A(n8476), .B(n8519), .S(n8475), .Z(n8484) );
  NAND2_X1 U10107 ( .A1(n8485), .A2(n8484), .ZN(n8477) );
  INV_X1 U10108 ( .A(n8504), .ZN(n8481) );
  AND2_X1 U10109 ( .A1(n8499), .A2(n8479), .ZN(n8490) );
  AOI21_X1 U10110 ( .B1(n8499), .B2(n8734), .A(n9002), .ZN(n8482) );
  NOR2_X1 U10111 ( .A1(n8734), .A2(n8499), .ZN(n8492) );
  NOR4_X1 U10112 ( .A1(n8482), .A2(n8500), .A3(n8492), .A4(n8733), .ZN(n8497)
         );
  INV_X1 U10113 ( .A(n8999), .ZN(n8496) );
  INV_X1 U10114 ( .A(n8484), .ZN(n8486) );
  INV_X1 U10115 ( .A(n8487), .ZN(n8489) );
  NAND2_X1 U10116 ( .A1(n8734), .A2(n8490), .ZN(n8491) );
  OAI211_X1 U10117 ( .C1(n8493), .C2(n8492), .A(n8733), .B(n8491), .ZN(n8494)
         );
  OAI211_X1 U10118 ( .C1(n8497), .C2(n8496), .A(n8495), .B(n8494), .ZN(n8506)
         );
  INV_X1 U10119 ( .A(n8498), .ZN(n8501) );
  OAI211_X1 U10120 ( .C1(n8865), .C2(n8504), .A(n8503), .B(n8502), .ZN(n8505)
         );
  NAND3_X1 U10121 ( .A1(n8511), .A2(n8510), .A3(n9064), .ZN(n8512) );
  OAI211_X1 U10122 ( .C1(n8513), .C2(n8515), .A(n8512), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8514) );
  AOI22_X1 U10123 ( .A1(n8517), .A2(n8954), .B1(n10148), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8518) );
  OAI21_X1 U10124 ( .B1(n8519), .B2(n8925), .A(n8518), .ZN(n8520) );
  AOI21_X1 U10125 ( .B1(n8521), .B2(n8927), .A(n8520), .ZN(n8522) );
  OAI21_X1 U10126 ( .B1(n8516), .B2(n10148), .A(n8522), .ZN(P2_U3205) );
  NOR2_X1 U10127 ( .A1(n8523), .A2(n10129), .ZN(n8860) );
  NOR2_X1 U10128 ( .A1(n8524), .A2(n8925), .ZN(n8525) );
  AOI211_X1 U10129 ( .C1(n10148), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8860), .B(
        n8525), .ZN(n8528) );
  OR2_X1 U10130 ( .A1(n8526), .A2(n8958), .ZN(n8527) );
  OAI211_X1 U10131 ( .C1(n8529), .C2(n10148), .A(n8528), .B(n8527), .ZN(
        P2_U3204) );
  INV_X1 U10132 ( .A(n8530), .ZN(n9060) );
  OAI222_X1 U10133 ( .A1(n10002), .A2(n8532), .B1(P1_U3086), .B2(n8531), .C1(
        n8589), .C2(n9060), .ZN(P1_U3327) );
  NAND2_X1 U10134 ( .A1(n9269), .A2(n9819), .ZN(n8536) );
  INV_X1 U10135 ( .A(n8533), .ZN(n8534) );
  AOI22_X1 U10136 ( .A1(n8534), .A2(n9842), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n10077), .ZN(n8535) );
  NAND2_X1 U10137 ( .A1(n8536), .A2(n8535), .ZN(n8537) );
  AOI21_X1 U10138 ( .B1(n8538), .B2(n9841), .A(n8537), .ZN(n8541) );
  NAND2_X1 U10139 ( .A1(n8539), .A2(n9848), .ZN(n8540) );
  OAI211_X1 U10140 ( .C1(n8542), .C2(n9850), .A(n8541), .B(n8540), .ZN(
        P1_U3356) );
  NAND2_X1 U10141 ( .A1(n8581), .A2(n8543), .ZN(n8546) );
  NAND2_X1 U10142 ( .A1(n9421), .A2(n8544), .ZN(n8545) );
  NAND2_X1 U10143 ( .A1(n8546), .A2(n8545), .ZN(n8548) );
  XNOR2_X1 U10144 ( .A(n8548), .B(n8547), .ZN(n8552) );
  NAND2_X1 U10145 ( .A1(n8581), .A2(n6727), .ZN(n8549) );
  OAI21_X1 U10146 ( .B1(n8550), .B2(n6918), .A(n8549), .ZN(n8551) );
  XNOR2_X1 U10147 ( .A(n8552), .B(n8551), .ZN(n8553) );
  INV_X1 U10148 ( .A(n8553), .ZN(n8558) );
  NAND3_X1 U10149 ( .A1(n8559), .A2(n9175), .A3(n8558), .ZN(n8564) );
  NAND2_X1 U10150 ( .A1(n9628), .A2(n9177), .ZN(n8557) );
  INV_X1 U10151 ( .A(n8579), .ZN(n8555) );
  AOI22_X1 U10152 ( .A1(n8555), .A2(n9183), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n8556) );
  OAI211_X1 U10153 ( .C1(n9270), .C2(n9181), .A(n8557), .B(n8556), .ZN(n8561)
         );
  NOR3_X1 U10154 ( .A1(n8559), .A2(n8558), .A3(n9170), .ZN(n8560) );
  AOI211_X1 U10155 ( .C1(n9168), .C2(n8581), .A(n8561), .B(n8560), .ZN(n8562)
         );
  OAI211_X1 U10156 ( .C1(n8565), .C2(n8564), .A(n8563), .B(n8562), .ZN(
        P1_U3220) );
  NAND2_X1 U10157 ( .A1(n8865), .A2(n8704), .ZN(n8569) );
  AOI22_X1 U10158 ( .A1(n8872), .A2(n8727), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8568) );
  OAI211_X1 U10159 ( .C1(n8570), .C2(n8707), .A(n8569), .B(n8568), .ZN(n8571)
         );
  AOI21_X1 U10160 ( .B1(n8962), .B2(n8711), .A(n8571), .ZN(n8572) );
  OAI222_X1 U10161 ( .A1(n9062), .A2(n8575), .B1(n9063), .B2(n8574), .C1(n6057), .C2(P2_U3151), .ZN(P2_U3274) );
  INV_X1 U10162 ( .A(n8576), .ZN(n8577) );
  NAND2_X1 U10163 ( .A1(n8577), .A2(n9700), .ZN(n8586) );
  INV_X1 U10164 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n8578) );
  OAI22_X1 U10165 ( .A1(n8579), .A2(n10072), .B1(n8578), .B2(n9848), .ZN(n8580) );
  AOI21_X1 U10166 ( .B1(n8581), .B2(n9819), .A(n8580), .ZN(n8582) );
  OAI21_X1 U10167 ( .B1(n8583), .B2(n10075), .A(n8582), .ZN(n8584) );
  INV_X1 U10168 ( .A(n8584), .ZN(n8585) );
  OAI211_X1 U10169 ( .C1(n8587), .C2(n10077), .A(n8586), .B(n8585), .ZN(
        P1_U3265) );
  INV_X1 U10170 ( .A(n8588), .ZN(n9053) );
  OAI222_X1 U10171 ( .A1(n10002), .A2(n8590), .B1(n8589), .B2(n9053), .C1(
        n5585), .C2(P1_U3086), .ZN(P1_U3325) );
  XOR2_X1 U10172 ( .A(n8592), .B(n8591), .Z(n8600) );
  NAND2_X1 U10173 ( .A1(n8704), .A2(n8743), .ZN(n8593) );
  NAND2_X1 U10174 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8793) );
  OAI211_X1 U10175 ( .C1(n8594), .C2(n8707), .A(n8593), .B(n8793), .ZN(n8595)
         );
  AOI21_X1 U10176 ( .B1(n8596), .B2(n8727), .A(n8595), .ZN(n8599) );
  NAND2_X1 U10177 ( .A1(n8597), .A2(n8711), .ZN(n8598) );
  OAI211_X1 U10178 ( .C1(n8600), .C2(n8717), .A(n8599), .B(n8598), .ZN(
        P2_U3155) );
  AOI21_X1 U10179 ( .B1(n8738), .B2(n8602), .A(n8649), .ZN(n8607) );
  AOI22_X1 U10180 ( .A1(n8910), .A2(n8722), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8604) );
  NAND2_X1 U10181 ( .A1(n8914), .A2(n8727), .ZN(n8603) );
  OAI211_X1 U10182 ( .C1(n8624), .C2(n8724), .A(n8604), .B(n8603), .ZN(n8605)
         );
  AOI21_X1 U10183 ( .B1(n9021), .B2(n8711), .A(n8605), .ZN(n8606) );
  OAI21_X1 U10184 ( .B1(n8607), .B2(n8717), .A(n8606), .ZN(P2_U3156) );
  XNOR2_X1 U10185 ( .A(n8608), .B(n6338), .ZN(n8609) );
  XNOR2_X1 U10186 ( .A(n8610), .B(n8609), .ZN(n8617) );
  NAND2_X1 U10187 ( .A1(n8740), .A2(n8722), .ZN(n8612) );
  OAI211_X1 U10188 ( .C1(n8948), .C2(n8724), .A(n8612), .B(n8611), .ZN(n8615)
         );
  NOR2_X1 U10189 ( .A1(n8613), .A2(n8731), .ZN(n8614) );
  AOI211_X1 U10190 ( .C1(n8953), .C2(n8727), .A(n8615), .B(n8614), .ZN(n8616)
         );
  OAI21_X1 U10191 ( .B1(n8617), .B2(n8717), .A(n8616), .ZN(P2_U3159) );
  AND3_X1 U10192 ( .A1(n8620), .A2(n8619), .A3(n8618), .ZN(n8622) );
  OAI21_X1 U10193 ( .B1(n8622), .B2(n8621), .A(n8679), .ZN(n8627) );
  AOI22_X1 U10194 ( .A1(n8894), .A2(n8727), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8623) );
  OAI21_X1 U10195 ( .B1(n8624), .B2(n8707), .A(n8623), .ZN(n8625) );
  AOI21_X1 U10196 ( .B1(n8891), .B2(n8704), .A(n8625), .ZN(n8626) );
  OAI211_X1 U10197 ( .C1(n8892), .C2(n8731), .A(n8627), .B(n8626), .ZN(
        P2_U3165) );
  XNOR2_X1 U10198 ( .A(n8628), .B(n8725), .ZN(n8629) );
  XNOR2_X1 U10199 ( .A(n8630), .B(n8629), .ZN(n8637) );
  NAND2_X1 U10200 ( .A1(n8722), .A2(n8743), .ZN(n8631) );
  NAND2_X1 U10201 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8827) );
  OAI211_X1 U10202 ( .C1(n8708), .C2(n8724), .A(n8631), .B(n8827), .ZN(n8632)
         );
  AOI21_X1 U10203 ( .B1(n8633), .B2(n8727), .A(n8632), .ZN(n8636) );
  NAND2_X1 U10204 ( .A1(n8634), .A2(n8711), .ZN(n8635) );
  OAI211_X1 U10205 ( .C1(n8637), .C2(n8717), .A(n8636), .B(n8635), .ZN(
        P2_U3166) );
  NAND2_X1 U10206 ( .A1(n8700), .A2(n8638), .ZN(n8640) );
  XOR2_X1 U10207 ( .A(n8640), .B(n8639), .Z(n8647) );
  NAND2_X1 U10208 ( .A1(n8722), .A2(n8741), .ZN(n8641) );
  NAND2_X1 U10209 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8844) );
  OAI211_X1 U10210 ( .C1(n8947), .C2(n8724), .A(n8641), .B(n8844), .ZN(n8642)
         );
  AOI21_X1 U10211 ( .B1(n8643), .B2(n8727), .A(n8642), .ZN(n8646) );
  NAND2_X1 U10212 ( .A1(n8644), .A2(n8711), .ZN(n8645) );
  OAI211_X1 U10213 ( .C1(n8647), .C2(n8717), .A(n8646), .B(n8645), .ZN(
        P2_U3168) );
  OAI21_X1 U10214 ( .B1(n8651), .B2(n8650), .A(n8679), .ZN(n8655) );
  AOI22_X1 U10215 ( .A1(n8901), .A2(n8727), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8652) );
  OAI21_X1 U10216 ( .B1(n8920), .B2(n8707), .A(n8652), .ZN(n8653) );
  AOI21_X1 U10217 ( .B1(n8737), .B2(n8704), .A(n8653), .ZN(n8654) );
  OAI211_X1 U10218 ( .C1(n4864), .C2(n8731), .A(n8655), .B(n8654), .ZN(
        P2_U3169) );
  AOI211_X1 U10219 ( .C1(n8658), .C2(n8657), .A(n8717), .B(n8656), .ZN(n8659)
         );
  INV_X1 U10220 ( .A(n8659), .ZN(n8663) );
  AOI22_X1 U10221 ( .A1(n8933), .A2(n8722), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8660) );
  OAI21_X1 U10222 ( .B1(n8919), .B2(n8724), .A(n8660), .ZN(n8661) );
  AOI21_X1 U10223 ( .B1(n8937), .B2(n8727), .A(n8661), .ZN(n8662) );
  OAI211_X1 U10224 ( .C1(n6131), .C2(n8731), .A(n8663), .B(n8662), .ZN(
        P2_U3173) );
  NAND2_X1 U10225 ( .A1(n8665), .A2(n8664), .ZN(n8667) );
  XOR2_X1 U10226 ( .A(n8667), .B(n8666), .Z(n8674) );
  NAND2_X1 U10227 ( .A1(n8722), .A2(n8745), .ZN(n8668) );
  NAND2_X1 U10228 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8776) );
  OAI211_X1 U10229 ( .C1(n8669), .C2(n8724), .A(n8668), .B(n8776), .ZN(n8670)
         );
  AOI21_X1 U10230 ( .B1(n8671), .B2(n8727), .A(n8670), .ZN(n8673) );
  NAND2_X1 U10231 ( .A1(n8016), .A2(n8711), .ZN(n8672) );
  OAI211_X1 U10232 ( .C1(n8674), .C2(n8717), .A(n8673), .B(n8672), .ZN(
        P2_U3174) );
  OAI21_X1 U10233 ( .B1(n8678), .B2(n8677), .A(n8676), .ZN(n8681) );
  NAND3_X1 U10234 ( .A1(n8681), .A2(n8680), .A3(n8679), .ZN(n8686) );
  INV_X1 U10235 ( .A(n8923), .ZN(n8683) );
  AOI22_X1 U10236 ( .A1(n8934), .A2(n8722), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8682) );
  OAI21_X1 U10237 ( .B1(n8683), .B2(n8696), .A(n8682), .ZN(n8684) );
  AOI21_X1 U10238 ( .B1(n8704), .B2(n8738), .A(n8684), .ZN(n8685) );
  OAI211_X1 U10239 ( .C1(n9028), .C2(n8731), .A(n8686), .B(n8685), .ZN(
        P2_U3175) );
  OAI22_X1 U10240 ( .A1(n8689), .A2(n8688), .B1(n8747), .B2(n8687), .ZN(n8690)
         );
  XOR2_X1 U10241 ( .A(n8691), .B(n8690), .Z(n8699) );
  OAI21_X1 U10242 ( .B1(n8707), .B2(n5836), .A(n8692), .ZN(n8693) );
  AOI21_X1 U10243 ( .B1(n8704), .B2(n8745), .A(n8693), .ZN(n8694) );
  OAI21_X1 U10244 ( .B1(n8696), .B2(n8695), .A(n8694), .ZN(n8697) );
  AOI21_X1 U10245 ( .B1(n6113), .B2(n8711), .A(n8697), .ZN(n8698) );
  OAI21_X1 U10246 ( .B1(n8699), .B2(n8717), .A(n8698), .ZN(P2_U3176) );
  NAND2_X1 U10247 ( .A1(n8701), .A2(n8700), .ZN(n8702) );
  XOR2_X1 U10248 ( .A(n8703), .B(n8702), .Z(n8715) );
  NAND2_X1 U10249 ( .A1(n8933), .A2(n8704), .ZN(n8706) );
  OAI211_X1 U10250 ( .C1(n8708), .C2(n8707), .A(n8706), .B(n8705), .ZN(n8709)
         );
  AOI21_X1 U10251 ( .B1(n8710), .B2(n8727), .A(n8709), .ZN(n8714) );
  NAND2_X1 U10252 ( .A1(n8712), .A2(n8711), .ZN(n8713) );
  OAI211_X1 U10253 ( .C1(n8715), .C2(n8717), .A(n8714), .B(n8713), .ZN(
        P2_U3178) );
  INV_X1 U10254 ( .A(n8716), .ZN(n8732) );
  AOI21_X1 U10255 ( .B1(n8719), .B2(n8718), .A(n8717), .ZN(n8721) );
  NAND2_X1 U10256 ( .A1(n8721), .A2(n8720), .ZN(n8730) );
  NAND2_X1 U10257 ( .A1(n8722), .A2(n8744), .ZN(n8723) );
  NAND2_X1 U10258 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8814) );
  OAI211_X1 U10259 ( .C1(n8725), .C2(n8724), .A(n8723), .B(n8814), .ZN(n8726)
         );
  AOI21_X1 U10260 ( .B1(n8728), .B2(n8727), .A(n8726), .ZN(n8729) );
  OAI211_X1 U10261 ( .C1(n8732), .C2(n8731), .A(n8730), .B(n8729), .ZN(
        P2_U3181) );
  MUX2_X1 U10262 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8733), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10263 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8734), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10264 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8735), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10265 ( .A(n8865), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8742), .Z(
        P2_U3519) );
  MUX2_X1 U10266 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8736), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10267 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8891), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10268 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8737), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10269 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8911), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10270 ( .A(n8738), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8742), .Z(
        P2_U3514) );
  MUX2_X1 U10271 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8910), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10272 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8934), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10273 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8739), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10274 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8933), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10275 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8740), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10276 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8741), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10277 ( .A(n8743), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8742), .Z(
        P2_U3506) );
  MUX2_X1 U10278 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8744), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10279 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n6118), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10280 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8745), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U10281 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8746), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10282 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8747), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10283 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8748), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10284 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8749), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U10285 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8750), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U10286 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8751), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U10287 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8752), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U10288 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8753), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U10289 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n10130), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U10290 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n6094), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U10291 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6091), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U10292 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8754), .S(P2_U3893), .Z(
        P2_U3491) );
  AOI21_X1 U10293 ( .B1(n8757), .B2(n8756), .A(n8755), .ZN(n8758) );
  INV_X1 U10294 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10358) );
  OAI22_X1 U10295 ( .A1(n8856), .A2(n8758), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10358), .ZN(n8759) );
  AOI21_X1 U10296 ( .B1(n8848), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n8759), .ZN(
        n8772) );
  OAI21_X1 U10297 ( .B1(n8762), .B2(n8761), .A(n8760), .ZN(n8765) );
  AOI22_X1 U10298 ( .A1(n8853), .A2(n8765), .B1(n8764), .B2(n8763), .ZN(n8771)
         );
  OAI211_X1 U10299 ( .C1(n8769), .C2(n8768), .A(n8767), .B(n8766), .ZN(n8770)
         );
  NAND3_X1 U10300 ( .A1(n8772), .A2(n8771), .A3(n8770), .ZN(P2_U3184) );
  XOR2_X1 U10301 ( .A(n8774), .B(n8773), .Z(n8786) );
  OAI21_X1 U10302 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n8775), .A(n8798), .ZN(
        n8784) );
  NAND2_X1 U10303 ( .A1(n8848), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n8777) );
  OAI211_X1 U10304 ( .C1(n8846), .C2(n8778), .A(n8777), .B(n8776), .ZN(n8783)
         );
  AOI21_X1 U10305 ( .B1(n8780), .B2(n8779), .A(n8791), .ZN(n8781) );
  NOR2_X1 U10306 ( .A1(n8781), .A2(n8856), .ZN(n8782) );
  AOI211_X1 U10307 ( .C1(n8853), .C2(n8784), .A(n8783), .B(n8782), .ZN(n8785)
         );
  OAI21_X1 U10308 ( .B1(n8786), .B2(n8850), .A(n8785), .ZN(P2_U3195) );
  XOR2_X1 U10309 ( .A(n8788), .B(n8787), .Z(n8805) );
  NOR3_X1 U10310 ( .A1(n8791), .A2(n8790), .A3(n8789), .ZN(n8792) );
  OAI21_X1 U10311 ( .B1(n4391), .B2(n8792), .A(n8825), .ZN(n8804) );
  OAI21_X1 U10312 ( .B1(n8846), .B2(n8794), .A(n8793), .ZN(n8802) );
  INV_X1 U10313 ( .A(n8795), .ZN(n8800) );
  NAND3_X1 U10314 ( .A1(n8798), .A2(n8797), .A3(n8796), .ZN(n8799) );
  AOI21_X1 U10315 ( .B1(n8800), .B2(n8799), .A(n8835), .ZN(n8801) );
  AOI211_X1 U10316 ( .C1(n8848), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n8802), .B(
        n8801), .ZN(n8803) );
  OAI211_X1 U10317 ( .C1(n8805), .C2(n8850), .A(n8804), .B(n8803), .ZN(
        P2_U3196) );
  XOR2_X1 U10318 ( .A(n8807), .B(n8806), .Z(n8819) );
  OAI21_X1 U10319 ( .B1(n4335), .B2(P2_REG1_REG_15__SCAN_IN), .A(n8808), .ZN(
        n8813) );
  INV_X1 U10320 ( .A(n8809), .ZN(n8810) );
  OAI21_X1 U10321 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n8811), .A(n8810), .ZN(
        n8812) );
  AOI22_X1 U10322 ( .A1(n8813), .A2(n8825), .B1(n8853), .B2(n8812), .ZN(n8818)
         );
  OAI21_X1 U10323 ( .B1(n8846), .B2(n8815), .A(n8814), .ZN(n8816) );
  AOI21_X1 U10324 ( .B1(n8848), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8816), .ZN(
        n8817) );
  OAI211_X1 U10325 ( .C1(n8819), .C2(n8850), .A(n8818), .B(n8817), .ZN(
        P2_U3197) );
  AOI21_X1 U10326 ( .B1(n4333), .B2(n8821), .A(n8820), .ZN(n8836) );
  OAI21_X1 U10327 ( .B1(n8824), .B2(n8823), .A(n8822), .ZN(n8826) );
  NAND2_X1 U10328 ( .A1(n8826), .A2(n8825), .ZN(n8834) );
  OAI21_X1 U10329 ( .B1(n8846), .B2(n4929), .A(n8827), .ZN(n8832) );
  XOR2_X1 U10330 ( .A(n8829), .B(n8828), .Z(n8830) );
  NOR2_X1 U10331 ( .A1(n8830), .A2(n8850), .ZN(n8831) );
  AOI211_X1 U10332 ( .C1(n8848), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n8832), .B(
        n8831), .ZN(n8833) );
  OAI211_X1 U10333 ( .C1(n8836), .C2(n8835), .A(n8834), .B(n8833), .ZN(
        P2_U3198) );
  INV_X1 U10334 ( .A(n8837), .ZN(n8838) );
  AOI21_X1 U10335 ( .B1(n8840), .B2(n8839), .A(n8838), .ZN(n8857) );
  OAI21_X1 U10336 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n8841), .A(n6689), .ZN(
        n8854) );
  XOR2_X1 U10337 ( .A(n8843), .B(n8842), .Z(n8851) );
  OAI21_X1 U10338 ( .B1(n8846), .B2(n8845), .A(n8844), .ZN(n8847) );
  AOI21_X1 U10339 ( .B1(n8848), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8847), .ZN(
        n8849) );
  OAI21_X1 U10340 ( .B1(n8851), .B2(n8850), .A(n8849), .ZN(n8852) );
  AOI21_X1 U10341 ( .B1(n8854), .B2(n8853), .A(n8852), .ZN(n8855) );
  OAI21_X1 U10342 ( .B1(n8857), .B2(n8856), .A(n8855), .ZN(P2_U3199) );
  NOR2_X1 U10343 ( .A1(n8859), .A2(n8858), .ZN(n8997) );
  AOI21_X1 U10344 ( .B1(n8997), .B2(n10145), .A(n8860), .ZN(n8863) );
  NAND2_X1 U10345 ( .A1(n10148), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8861) );
  OAI211_X1 U10346 ( .C1(n8999), .C2(n8925), .A(n8863), .B(n8861), .ZN(
        P2_U3202) );
  NAND2_X1 U10347 ( .A1(n10148), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8862) );
  OAI211_X1 U10348 ( .C1(n9002), .C2(n8925), .A(n8863), .B(n8862), .ZN(
        P2_U3203) );
  XNOR2_X1 U10349 ( .A(n8871), .B(n8870), .ZN(n8965) );
  INV_X1 U10350 ( .A(n8965), .ZN(n8876) );
  AOI22_X1 U10351 ( .A1(n8872), .A2(n8954), .B1(n10148), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8873) );
  OAI21_X1 U10352 ( .B1(n8874), .B2(n8925), .A(n8873), .ZN(n8875) );
  AOI21_X1 U10353 ( .B1(n8876), .B2(n8927), .A(n8875), .ZN(n8877) );
  OAI21_X1 U10354 ( .B1(n8964), .B2(n10148), .A(n8877), .ZN(P2_U3206) );
  XNOR2_X1 U10355 ( .A(n8878), .B(n8879), .ZN(n9006) );
  AOI22_X1 U10356 ( .A1(n8884), .A2(n8955), .B1(n8954), .B2(n8883), .ZN(n8885)
         );
  OAI211_X1 U10357 ( .C1(n9006), .C2(n8958), .A(n8886), .B(n8885), .ZN(
        P2_U3207) );
  XNOR2_X1 U10358 ( .A(n8888), .B(n8887), .ZN(n9014) );
  OAI21_X1 U10359 ( .B1(n8892), .B2(n10128), .A(n9009), .ZN(n8893) );
  NAND2_X1 U10360 ( .A1(n8893), .A2(n10145), .ZN(n8896) );
  AOI22_X1 U10361 ( .A1(n8894), .A2(n8954), .B1(n10148), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8895) );
  NOR2_X1 U10362 ( .A1(n4864), .A2(n10128), .ZN(n8900) );
  XOR2_X1 U10363 ( .A(n8903), .B(n8897), .Z(n8898) );
  OAI222_X1 U10364 ( .A1(n4652), .A2(n8899), .B1(n8946), .B2(n8920), .C1(n8898), .C2(n10151), .ZN(n9015) );
  AOI211_X1 U10365 ( .C1(n8954), .C2(n8901), .A(n8900), .B(n9015), .ZN(n8906)
         );
  XOR2_X1 U10366 ( .A(n8903), .B(n8902), .Z(n9016) );
  INV_X1 U10367 ( .A(n9016), .ZN(n8904) );
  AOI22_X1 U10368 ( .A1(n8904), .A2(n8927), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n10148), .ZN(n8905) );
  OAI21_X1 U10369 ( .B1(n8906), .B2(n10148), .A(n8905), .ZN(P2_U3209) );
  XNOR2_X1 U10370 ( .A(n8907), .B(n8909), .ZN(n9024) );
  XOR2_X1 U10371 ( .A(n8908), .B(n8909), .Z(n8912) );
  AOI222_X1 U10372 ( .A1(n10136), .A2(n8912), .B1(n8911), .B2(n10131), .C1(
        n8910), .C2(n10132), .ZN(n9019) );
  MUX2_X1 U10373 ( .A(n8913), .B(n9019), .S(n10145), .Z(n8916) );
  AOI22_X1 U10374 ( .A1(n9021), .A2(n8955), .B1(n8954), .B2(n8914), .ZN(n8915)
         );
  OAI211_X1 U10375 ( .C1(n9024), .C2(n8958), .A(n8916), .B(n8915), .ZN(
        P2_U3210) );
  XOR2_X1 U10376 ( .A(n8917), .B(n8921), .Z(n8918) );
  OAI222_X1 U10377 ( .A1(n4652), .A2(n8920), .B1(n8946), .B2(n8919), .C1(
        n10151), .C2(n8918), .ZN(n8976) );
  INV_X1 U10378 ( .A(n8976), .ZN(n8929) );
  XNOR2_X1 U10379 ( .A(n8922), .B(n8921), .ZN(n8977) );
  AOI22_X1 U10380 ( .A1(n8923), .A2(n8954), .B1(n10148), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n8924) );
  OAI21_X1 U10381 ( .B1(n9028), .B2(n8925), .A(n8924), .ZN(n8926) );
  AOI21_X1 U10382 ( .B1(n8977), .B2(n8927), .A(n8926), .ZN(n8928) );
  OAI21_X1 U10383 ( .B1(n8929), .B2(n10148), .A(n8928), .ZN(P2_U3211) );
  XNOR2_X1 U10384 ( .A(n8932), .B(n8930), .ZN(n9034) );
  OAI21_X1 U10385 ( .B1(n4383), .B2(n8932), .A(n8931), .ZN(n8935) );
  AOI222_X1 U10386 ( .A1(n10136), .A2(n8935), .B1(n8934), .B2(n10131), .C1(
        n8933), .C2(n10132), .ZN(n9029) );
  MUX2_X1 U10387 ( .A(n8936), .B(n9029), .S(n10145), .Z(n8939) );
  AOI22_X1 U10388 ( .A1(n9031), .A2(n8955), .B1(n8954), .B2(n8937), .ZN(n8938)
         );
  OAI211_X1 U10389 ( .C1(n9034), .C2(n8958), .A(n8939), .B(n8938), .ZN(
        P2_U3213) );
  XNOR2_X1 U10390 ( .A(n8940), .B(n8941), .ZN(n9040) );
  NAND2_X1 U10391 ( .A1(n8942), .A2(n8941), .ZN(n8943) );
  NAND2_X1 U10392 ( .A1(n8943), .A2(n10136), .ZN(n8944) );
  OR2_X1 U10393 ( .A1(n8945), .A2(n8944), .ZN(n8951) );
  OAI22_X1 U10394 ( .A1(n8948), .A2(n4652), .B1(n8947), .B2(n8946), .ZN(n8949)
         );
  INV_X1 U10395 ( .A(n8949), .ZN(n8950) );
  MUX2_X1 U10396 ( .A(n9036), .B(n8952), .S(n10148), .Z(n8957) );
  AOI22_X1 U10397 ( .A1(n6130), .A2(n8955), .B1(n8954), .B2(n8953), .ZN(n8956)
         );
  OAI211_X1 U10398 ( .C1(n9040), .C2(n8958), .A(n8957), .B(n8956), .ZN(
        P2_U3214) );
  NAND2_X1 U10399 ( .A1(n6372), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8959) );
  NAND2_X1 U10400 ( .A1(n8997), .A2(n10199), .ZN(n8961) );
  OAI211_X1 U10401 ( .C1(n8999), .C2(n8991), .A(n8959), .B(n8961), .ZN(
        P2_U3490) );
  NAND2_X1 U10402 ( .A1(n6372), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8960) );
  OAI211_X1 U10403 ( .C1(n9002), .C2(n8991), .A(n8961), .B(n8960), .ZN(
        P2_U3489) );
  NAND2_X1 U10404 ( .A1(n8962), .A2(n10157), .ZN(n8963) );
  OAI211_X1 U10405 ( .C1(n10180), .C2(n8965), .A(n8964), .B(n8963), .ZN(n9003)
         );
  MUX2_X1 U10406 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9003), .S(n10199), .Z(
        P2_U3486) );
  MUX2_X1 U10407 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9004), .S(n10199), .Z(
        n8967) );
  OAI22_X1 U10408 ( .A1(n9006), .A2(n8986), .B1(n9005), .B2(n8991), .ZN(n8966)
         );
  OR2_X1 U10409 ( .A1(n8967), .A2(n8966), .ZN(P2_U3485) );
  INV_X1 U10410 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8968) );
  MUX2_X1 U10411 ( .A(n8968), .B(n9009), .S(n10199), .Z(n8970) );
  NAND2_X1 U10412 ( .A1(n9011), .A2(n8983), .ZN(n8969) );
  OAI211_X1 U10413 ( .C1(n9014), .C2(n8986), .A(n8970), .B(n8969), .ZN(
        P2_U3484) );
  MUX2_X1 U10414 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9015), .S(n10199), .Z(
        n8972) );
  OAI22_X1 U10415 ( .A1(n9016), .A2(n8986), .B1(n4864), .B2(n8991), .ZN(n8971)
         );
  OR2_X1 U10416 ( .A1(n8972), .A2(n8971), .ZN(P2_U3483) );
  INV_X1 U10417 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8973) );
  MUX2_X1 U10418 ( .A(n8973), .B(n9019), .S(n10199), .Z(n8975) );
  NAND2_X1 U10419 ( .A1(n9021), .A2(n8983), .ZN(n8974) );
  OAI211_X1 U10420 ( .C1(n9024), .C2(n8986), .A(n8975), .B(n8974), .ZN(
        P2_U3482) );
  AOI21_X1 U10421 ( .B1(n6186), .B2(n8977), .A(n8976), .ZN(n9025) );
  MUX2_X1 U10422 ( .A(n10279), .B(n9025), .S(n10199), .Z(n8978) );
  OAI21_X1 U10423 ( .B1(n9028), .B2(n8991), .A(n8978), .ZN(P2_U3481) );
  INV_X1 U10424 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8979) );
  MUX2_X1 U10425 ( .A(n8979), .B(n9029), .S(n10199), .Z(n8981) );
  NAND2_X1 U10426 ( .A1(n9031), .A2(n8983), .ZN(n8980) );
  OAI211_X1 U10427 ( .C1(n8986), .C2(n9034), .A(n8981), .B(n8980), .ZN(
        P2_U3479) );
  INV_X1 U10428 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8982) );
  MUX2_X1 U10429 ( .A(n8982), .B(n9036), .S(n10199), .Z(n8985) );
  NAND2_X1 U10430 ( .A1(n6130), .A2(n8983), .ZN(n8984) );
  OAI211_X1 U10431 ( .C1(n9040), .C2(n8986), .A(n8985), .B(n8984), .ZN(
        P2_U3478) );
  NAND2_X1 U10432 ( .A1(n8987), .A2(n6186), .ZN(n8988) );
  AND2_X1 U10433 ( .A1(n8989), .A2(n8988), .ZN(n9042) );
  MUX2_X1 U10434 ( .A(n9042), .B(n10275), .S(n6372), .Z(n8990) );
  OAI21_X1 U10435 ( .B1(n9045), .B2(n8991), .A(n8990), .ZN(P2_U3477) );
  NAND3_X1 U10436 ( .A1(n8993), .A2(n6186), .A3(n8992), .ZN(n8994) );
  OAI211_X1 U10437 ( .C1(n8996), .C2(n10178), .A(n8995), .B(n8994), .ZN(n9046)
         );
  MUX2_X1 U10438 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9046), .S(n10199), .Z(
        P2_U3473) );
  NAND2_X1 U10439 ( .A1(n10186), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8998) );
  NAND2_X1 U10440 ( .A1(n8997), .A2(n10184), .ZN(n9001) );
  OAI211_X1 U10441 ( .C1(n8999), .C2(n9044), .A(n8998), .B(n9001), .ZN(
        P2_U3458) );
  NAND2_X1 U10442 ( .A1(n10186), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9000) );
  OAI211_X1 U10443 ( .C1(n9002), .C2(n9044), .A(n9001), .B(n9000), .ZN(
        P2_U3457) );
  MUX2_X1 U10444 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9003), .S(n10184), .Z(
        P2_U3454) );
  MUX2_X1 U10445 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9004), .S(n10184), .Z(
        n9008) );
  OAI22_X1 U10446 ( .A1(n9006), .A2(n9039), .B1(n9005), .B2(n9044), .ZN(n9007)
         );
  OR2_X1 U10447 ( .A1(n9008), .A2(n9007), .ZN(P2_U3453) );
  INV_X1 U10448 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9010) );
  MUX2_X1 U10449 ( .A(n9010), .B(n9009), .S(n10184), .Z(n9013) );
  NAND2_X1 U10450 ( .A1(n9011), .A2(n6375), .ZN(n9012) );
  OAI211_X1 U10451 ( .C1(n9014), .C2(n9039), .A(n9013), .B(n9012), .ZN(
        P2_U3452) );
  MUX2_X1 U10452 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9015), .S(n10184), .Z(
        n9018) );
  OAI22_X1 U10453 ( .A1(n9016), .A2(n9039), .B1(n4864), .B2(n9044), .ZN(n9017)
         );
  OR2_X1 U10454 ( .A1(n9018), .A2(n9017), .ZN(P2_U3451) );
  INV_X1 U10455 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9020) );
  MUX2_X1 U10456 ( .A(n9020), .B(n9019), .S(n10184), .Z(n9023) );
  NAND2_X1 U10457 ( .A1(n9021), .A2(n6375), .ZN(n9022) );
  OAI211_X1 U10458 ( .C1(n9024), .C2(n9039), .A(n9023), .B(n9022), .ZN(
        P2_U3450) );
  INV_X1 U10459 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9026) );
  MUX2_X1 U10460 ( .A(n9026), .B(n9025), .S(n10184), .Z(n9027) );
  OAI21_X1 U10461 ( .B1(n9028), .B2(n9044), .A(n9027), .ZN(P2_U3449) );
  INV_X1 U10462 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9030) );
  MUX2_X1 U10463 ( .A(n9030), .B(n9029), .S(n10184), .Z(n9033) );
  NAND2_X1 U10464 ( .A1(n9031), .A2(n6375), .ZN(n9032) );
  OAI211_X1 U10465 ( .C1(n9034), .C2(n9039), .A(n9033), .B(n9032), .ZN(
        P2_U3447) );
  INV_X1 U10466 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9035) );
  MUX2_X1 U10467 ( .A(n9036), .B(n9035), .S(n10186), .Z(n9038) );
  NAND2_X1 U10468 ( .A1(n6130), .A2(n6375), .ZN(n9037) );
  OAI211_X1 U10469 ( .C1(n9040), .C2(n9039), .A(n9038), .B(n9037), .ZN(
        P2_U3446) );
  INV_X1 U10470 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9041) );
  MUX2_X1 U10471 ( .A(n9042), .B(n9041), .S(n10186), .Z(n9043) );
  OAI21_X1 U10472 ( .B1(n9045), .B2(n9044), .A(n9043), .ZN(P2_U3444) );
  MUX2_X1 U10473 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n9046), .S(n10184), .Z(
        P2_U3432) );
  INV_X1 U10474 ( .A(n9988), .ZN(n9050) );
  NOR4_X1 U10475 ( .A1(n9047), .A2(P2_IR_REG_30__SCAN_IN), .A3(n4520), .A4(
        P2_U3151), .ZN(n9048) );
  AOI21_X1 U10476 ( .B1(n9058), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9048), .ZN(
        n9049) );
  OAI21_X1 U10477 ( .B1(n9050), .B2(n9063), .A(n9049), .ZN(P2_U3264) );
  AOI22_X1 U10478 ( .A1(n9051), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9058), .ZN(n9052) );
  OAI21_X1 U10479 ( .B1(n9053), .B2(n9063), .A(n9052), .ZN(P2_U3265) );
  INV_X1 U10480 ( .A(n9054), .ZN(n9995) );
  AOI22_X1 U10481 ( .A1(n9055), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9058), .ZN(n9056) );
  OAI21_X1 U10482 ( .B1(n9995), .B2(n9063), .A(n9056), .ZN(P2_U3266) );
  AOI21_X1 U10483 ( .B1(n9058), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n9057), .ZN(
        n9059) );
  OAI21_X1 U10484 ( .B1(n9060), .B2(n9063), .A(n9059), .ZN(P2_U3267) );
  INV_X1 U10485 ( .A(n9061), .ZN(n9998) );
  OAI222_X1 U10486 ( .A1(P2_U3151), .A2(n9064), .B1(n9063), .B2(n9998), .C1(
        n10375), .C2(n9062), .ZN(P2_U3268) );
  MUX2_X1 U10487 ( .A(n9065), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AOI21_X1 U10488 ( .B1(n9067), .B2(n9066), .A(n9123), .ZN(n9072) );
  NAND2_X1 U10489 ( .A1(n9673), .A2(n9155), .ZN(n9069) );
  AOI22_X1 U10490 ( .A1(n9714), .A2(n9177), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9068) );
  OAI211_X1 U10491 ( .C1(n9164), .C2(n9676), .A(n9069), .B(n9068), .ZN(n9070)
         );
  AOI21_X1 U10492 ( .B1(n9947), .B2(n9168), .A(n9070), .ZN(n9071) );
  OAI21_X1 U10493 ( .B1(n9072), .B2(n9170), .A(n9071), .ZN(P1_U3216) );
  OAI21_X1 U10494 ( .B1(n9075), .B2(n9074), .A(n4673), .ZN(n9076) );
  NAND2_X1 U10495 ( .A1(n9076), .A2(n9175), .ZN(n9081) );
  NAND2_X1 U10496 ( .A1(n9177), .A2(n9776), .ZN(n9077) );
  NAND2_X1 U10497 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9594) );
  OAI211_X1 U10498 ( .C1(n9078), .C2(n9181), .A(n9077), .B(n9594), .ZN(n9079)
         );
  AOI21_X1 U10499 ( .B1(n9747), .B2(n9183), .A(n9079), .ZN(n9080) );
  OAI211_X1 U10500 ( .C1(n9749), .C2(n9186), .A(n9081), .B(n9080), .ZN(
        P1_U3219) );
  XNOR2_X1 U10501 ( .A(n9082), .B(n5137), .ZN(n9083) );
  XNOR2_X1 U10502 ( .A(n9084), .B(n9083), .ZN(n9089) );
  AOI22_X1 U10503 ( .A1(n9752), .A2(n9177), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9086) );
  NAND2_X1 U10504 ( .A1(n9183), .A2(n9718), .ZN(n9085) );
  OAI211_X1 U10505 ( .C1(n9253), .C2(n9181), .A(n9086), .B(n9085), .ZN(n9087)
         );
  AOI21_X1 U10506 ( .B1(n9955), .B2(n9168), .A(n9087), .ZN(n9088) );
  OAI21_X1 U10507 ( .B1(n9089), .B2(n9170), .A(n9088), .ZN(P1_U3223) );
  OAI21_X1 U10508 ( .B1(n9092), .B2(n9091), .A(n9090), .ZN(n9093) );
  NAND2_X1 U10509 ( .A1(n9093), .A2(n9175), .ZN(n9099) );
  NOR2_X1 U10510 ( .A1(n9094), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9095) );
  AOI21_X1 U10511 ( .B1(n9673), .B2(n9177), .A(n9095), .ZN(n9096) );
  OAI21_X1 U10512 ( .B1(n9642), .B2(n9164), .A(n9096), .ZN(n9097) );
  AOI21_X1 U10513 ( .B1(n9637), .B2(n9155), .A(n9097), .ZN(n9098) );
  OAI211_X1 U10514 ( .C1(n5150), .C2(n9186), .A(n9099), .B(n9098), .ZN(
        P1_U3225) );
  XOR2_X1 U10515 ( .A(n9101), .B(n9102), .Z(n9174) );
  INV_X1 U10516 ( .A(n9100), .ZN(n9173) );
  NAND2_X1 U10517 ( .A1(n9174), .A2(n9173), .ZN(n9172) );
  OAI21_X1 U10518 ( .B1(n9102), .B2(n9101), .A(n9172), .ZN(n9106) );
  XNOR2_X1 U10519 ( .A(n9104), .B(n9103), .ZN(n9105) );
  XNOR2_X1 U10520 ( .A(n9106), .B(n9105), .ZN(n9111) );
  NOR2_X1 U10521 ( .A1(n9164), .A2(n9792), .ZN(n9109) );
  NAND2_X1 U10522 ( .A1(n9177), .A2(n9833), .ZN(n9107) );
  NAND2_X1 U10523 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9531) );
  OAI211_X1 U10524 ( .C1(n9181), .C2(n9801), .A(n9107), .B(n9531), .ZN(n9108)
         );
  AOI211_X1 U10525 ( .C1(n9911), .C2(n9168), .A(n9109), .B(n9108), .ZN(n9110)
         );
  OAI21_X1 U10526 ( .B1(n9111), .B2(n9170), .A(n9110), .ZN(P1_U3226) );
  XOR2_X1 U10527 ( .A(n9113), .B(n9112), .Z(n9119) );
  NAND2_X1 U10528 ( .A1(n9177), .A2(n9815), .ZN(n9114) );
  NAND2_X1 U10529 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9548) );
  OAI211_X1 U10530 ( .C1(n9181), .C2(n9115), .A(n9114), .B(n9548), .ZN(n9117)
         );
  NOR2_X1 U10531 ( .A1(n9783), .A2(n9186), .ZN(n9116) );
  AOI211_X1 U10532 ( .C1(n9183), .C2(n9780), .A(n9117), .B(n9116), .ZN(n9118)
         );
  OAI21_X1 U10533 ( .B1(n9119), .B2(n9170), .A(n9118), .ZN(P1_U3228) );
  INV_X1 U10534 ( .A(n9120), .ZN(n9125) );
  NOR3_X1 U10535 ( .A1(n9123), .A2(n9122), .A3(n9121), .ZN(n9124) );
  OAI21_X1 U10536 ( .B1(n9125), .B2(n9124), .A(n9175), .ZN(n9130) );
  INV_X1 U10537 ( .A(n9658), .ZN(n9128) );
  AOI22_X1 U10538 ( .A1(n9688), .A2(n9177), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9126) );
  OAI21_X1 U10539 ( .B1(n9653), .B2(n9181), .A(n9126), .ZN(n9127) );
  AOI21_X1 U10540 ( .B1(n9128), .B2(n9183), .A(n9127), .ZN(n9129) );
  OAI211_X1 U10541 ( .C1(n9944), .C2(n9186), .A(n9130), .B(n9129), .ZN(
        P1_U3229) );
  OAI211_X1 U10542 ( .C1(n9133), .C2(n9132), .A(n9131), .B(n9175), .ZN(n9139)
         );
  AOI22_X1 U10543 ( .A1(n9168), .A2(n9134), .B1(P1_REG3_REG_4__SCAN_IN), .B2(
        P1_U3086), .ZN(n9138) );
  AOI22_X1 U10544 ( .A1(n9155), .A2(n9428), .B1(n9177), .B2(n9430), .ZN(n9137)
         );
  NAND2_X1 U10545 ( .A1(n9183), .A2(n9135), .ZN(n9136) );
  NAND4_X1 U10546 ( .A1(n9139), .A2(n9138), .A3(n9137), .A4(n9136), .ZN(
        P1_U3230) );
  INV_X1 U10547 ( .A(n9140), .ZN(n9142) );
  NAND2_X1 U10548 ( .A1(n9142), .A2(n9141), .ZN(n9143) );
  XNOR2_X1 U10549 ( .A(n9144), .B(n9143), .ZN(n9150) );
  INV_X1 U10550 ( .A(n9145), .ZN(n9733) );
  NAND2_X1 U10551 ( .A1(n9183), .A2(n9733), .ZN(n9147) );
  INV_X1 U10552 ( .A(n9728), .ZN(n9768) );
  AOI22_X1 U10553 ( .A1(n9768), .A2(n9177), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9146) );
  OAI211_X1 U10554 ( .C1(n9729), .C2(n9181), .A(n9147), .B(n9146), .ZN(n9148)
         );
  AOI21_X1 U10555 ( .B1(n9734), .B2(n9168), .A(n9148), .ZN(n9149) );
  OAI21_X1 U10556 ( .B1(n9150), .B2(n9170), .A(n9149), .ZN(P1_U3233) );
  XNOR2_X1 U10557 ( .A(n9152), .B(n9151), .ZN(n9153) );
  XNOR2_X1 U10558 ( .A(n9154), .B(n9153), .ZN(n9160) );
  AOI22_X1 U10559 ( .A1(n9688), .A2(n9155), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9157) );
  NAND2_X1 U10560 ( .A1(n9687), .A2(n9177), .ZN(n9156) );
  OAI211_X1 U10561 ( .C1(n9164), .C2(n9695), .A(n9157), .B(n9156), .ZN(n9158)
         );
  AOI21_X1 U10562 ( .B1(n9877), .B2(n9168), .A(n9158), .ZN(n9159) );
  OAI21_X1 U10563 ( .B1(n9160), .B2(n9170), .A(n9159), .ZN(P1_U3235) );
  NOR2_X1 U10564 ( .A1(n9161), .A2(n4346), .ZN(n9163) );
  XNOR2_X1 U10565 ( .A(n9163), .B(n9162), .ZN(n9171) );
  NOR2_X1 U10566 ( .A1(n9164), .A2(n9760), .ZN(n9167) );
  NAND2_X1 U10567 ( .A1(n9177), .A2(n9767), .ZN(n9165) );
  NAND2_X1 U10568 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9575) );
  OAI211_X1 U10569 ( .C1(n9181), .C2(n9728), .A(n9165), .B(n9575), .ZN(n9166)
         );
  AOI211_X1 U10570 ( .C1(n9900), .C2(n9168), .A(n9167), .B(n9166), .ZN(n9169)
         );
  OAI21_X1 U10571 ( .B1(n9171), .B2(n9170), .A(n9169), .ZN(P1_U3238) );
  OAI21_X1 U10572 ( .B1(n9174), .B2(n9173), .A(n9172), .ZN(n9176) );
  NAND2_X1 U10573 ( .A1(n9176), .A2(n9175), .ZN(n9185) );
  NAND2_X1 U10574 ( .A1(n9177), .A2(n9814), .ZN(n9179) );
  OAI211_X1 U10575 ( .C1(n9181), .C2(n9180), .A(n9179), .B(n9178), .ZN(n9182)
         );
  AOI21_X1 U10576 ( .B1(n9818), .B2(n9183), .A(n9182), .ZN(n9184) );
  OAI211_X1 U10577 ( .C1(n9976), .C2(n9186), .A(n9185), .B(n9184), .ZN(
        P1_U3241) );
  OAI21_X1 U10578 ( .B1(n4963), .B2(n9312), .A(n9336), .ZN(n9268) );
  INV_X1 U10579 ( .A(n9352), .ZN(n9271) );
  NAND3_X1 U10580 ( .A1(n9249), .A2(n9271), .A3(n9395), .ZN(n9241) );
  NAND3_X1 U10581 ( .A1(n9249), .A2(n9749), .A3(n9395), .ZN(n9187) );
  OAI21_X1 U10582 ( .B1(n9728), .B2(n9271), .A(n9187), .ZN(n9188) );
  NAND2_X1 U10583 ( .A1(n9188), .A2(n9246), .ZN(n9240) );
  INV_X1 U10584 ( .A(n9233), .ZN(n9388) );
  OAI21_X1 U10585 ( .B1(n9388), .B2(n9799), .A(n9271), .ZN(n9234) );
  INV_X1 U10586 ( .A(n9234), .ZN(n9237) );
  AND2_X1 U10587 ( .A1(n9820), .A2(n9799), .ZN(n9189) );
  AOI21_X1 U10588 ( .B1(n9189), .B2(n9389), .A(n9388), .ZN(n9236) );
  NAND3_X1 U10589 ( .A1(n9190), .A2(n9195), .A3(n9271), .ZN(n9191) );
  NOR2_X1 U10590 ( .A1(n9201), .A2(n9191), .ZN(n9192) );
  NAND2_X1 U10591 ( .A1(n9193), .A2(n9192), .ZN(n9210) );
  NAND3_X1 U10592 ( .A1(n9196), .A2(n9195), .A3(n9194), .ZN(n9206) );
  NAND3_X1 U10593 ( .A1(n9197), .A2(n9367), .A3(n9352), .ZN(n9198) );
  NOR2_X1 U10594 ( .A1(n9201), .A2(n9198), .ZN(n9205) );
  NAND3_X1 U10595 ( .A1(n9200), .A2(n9199), .A3(n9352), .ZN(n9203) );
  NAND3_X1 U10596 ( .A1(n9427), .A2(n10108), .A3(n9271), .ZN(n9202) );
  AOI21_X1 U10597 ( .B1(n9203), .B2(n9202), .A(n9201), .ZN(n9204) );
  AOI21_X1 U10598 ( .B1(n9206), .B2(n9205), .A(n9204), .ZN(n9209) );
  MUX2_X1 U10599 ( .A(n9207), .B(n9288), .S(n9352), .Z(n9208) );
  NAND3_X1 U10600 ( .A1(n9210), .A2(n9209), .A3(n9208), .ZN(n9214) );
  MUX2_X1 U10601 ( .A(n9212), .B(n9211), .S(n9352), .Z(n9213) );
  NAND2_X1 U10602 ( .A1(n9377), .A2(n9218), .ZN(n9215) );
  AOI21_X1 U10603 ( .B1(n9219), .B2(n9286), .A(n9215), .ZN(n9216) );
  NAND2_X1 U10604 ( .A1(n9222), .A2(n9220), .ZN(n9376) );
  AND2_X1 U10605 ( .A1(n9224), .A2(n9221), .ZN(n9379) );
  OAI21_X1 U10606 ( .B1(n9216), .B2(n9376), .A(n9379), .ZN(n9217) );
  NAND2_X1 U10607 ( .A1(n9217), .A2(n9380), .ZN(n9226) );
  NAND3_X1 U10608 ( .A1(n9223), .A2(n9380), .A3(n9222), .ZN(n9225) );
  NOR2_X1 U10609 ( .A1(n9228), .A2(n9227), .ZN(n9383) );
  AND2_X1 U10610 ( .A1(n9387), .A2(n9810), .ZN(n9385) );
  NAND3_X1 U10611 ( .A1(n9229), .A2(n9385), .A3(n9389), .ZN(n9235) );
  OAI211_X1 U10612 ( .C1(n9846), .C2(n9814), .A(n9233), .B(n9232), .ZN(n9386)
         );
  AND2_X1 U10613 ( .A1(n9244), .A2(n9239), .ZN(n9394) );
  INV_X1 U10614 ( .A(n9242), .ZN(n9245) );
  NAND2_X1 U10615 ( .A1(n9396), .A2(n9243), .ZN(n9390) );
  OAI211_X1 U10616 ( .C1(n9245), .C2(n9390), .A(n9401), .B(n9244), .ZN(n9247)
         );
  NAND2_X1 U10617 ( .A1(n9683), .A2(n9246), .ZN(n9323) );
  INV_X1 U10618 ( .A(n9250), .ZN(n9327) );
  OAI211_X1 U10619 ( .C1(n9248), .C2(n9327), .A(n9255), .B(n9690), .ZN(n9258)
         );
  NAND2_X1 U10620 ( .A1(n9250), .A2(n9249), .ZN(n9320) );
  OAI21_X1 U10621 ( .B1(n9251), .B2(n9320), .A(n9683), .ZN(n9252) );
  NAND3_X1 U10622 ( .A1(n9252), .A2(n9690), .A3(n9352), .ZN(n9257) );
  OR2_X1 U10623 ( .A1(n9877), .A2(n9253), .ZN(n9254) );
  NAND2_X1 U10624 ( .A1(n9259), .A2(n9254), .ZN(n9314) );
  NAND2_X1 U10625 ( .A1(n9313), .A2(n9670), .ZN(n9324) );
  AOI22_X1 U10626 ( .A1(n9255), .A2(n9314), .B1(n9324), .B2(n9352), .ZN(n9256)
         );
  MUX2_X1 U10627 ( .A(n9316), .B(n9325), .S(n9352), .Z(n9261) );
  INV_X1 U10628 ( .A(n9262), .ZN(n9329) );
  OAI21_X1 U10629 ( .B1(n4966), .B2(n9329), .A(n9311), .ZN(n9266) );
  INV_X1 U10630 ( .A(n9311), .ZN(n9264) );
  INV_X1 U10631 ( .A(n9319), .ZN(n9263) );
  OAI21_X1 U10632 ( .B1(n9264), .B2(n9263), .A(n9322), .ZN(n9265) );
  MUX2_X1 U10633 ( .A(n9266), .B(n9265), .S(n9352), .Z(n9267) );
  INV_X1 U10634 ( .A(n9277), .ZN(n9419) );
  NAND2_X1 U10635 ( .A1(n9419), .A2(n9338), .ZN(n9342) );
  INV_X1 U10636 ( .A(n4796), .ZN(n9601) );
  NAND2_X1 U10637 ( .A1(n9352), .A2(n9601), .ZN(n9272) );
  NAND2_X1 U10638 ( .A1(n9274), .A2(n9273), .ZN(n9351) );
  INV_X1 U10639 ( .A(n9275), .ZN(n9276) );
  OR2_X1 U10640 ( .A1(n4796), .A2(n9277), .ZN(n9407) );
  NAND2_X1 U10641 ( .A1(n4796), .A2(n9277), .ZN(n9341) );
  NAND2_X1 U10642 ( .A1(n9407), .A2(n9341), .ZN(n9309) );
  INV_X1 U10643 ( .A(n9669), .ZN(n9301) );
  INV_X1 U10644 ( .A(n9278), .ZN(n9292) );
  NAND4_X1 U10645 ( .A1(n9280), .A2(n7399), .A3(n9279), .A4(n9366), .ZN(n9283)
         );
  NOR3_X1 U10646 ( .A1(n9283), .A2(n9282), .A3(n9281), .ZN(n9289) );
  NOR2_X1 U10647 ( .A1(n9285), .A2(n9284), .ZN(n9287) );
  NAND4_X1 U10648 ( .A1(n9289), .A2(n9288), .A3(n9287), .A4(n9286), .ZN(n9290)
         );
  NOR2_X1 U10649 ( .A1(n9290), .A2(n9374), .ZN(n9291) );
  NAND3_X1 U10650 ( .A1(n9293), .A2(n9292), .A3(n9291), .ZN(n9294) );
  NOR2_X1 U10651 ( .A1(n9295), .A2(n9294), .ZN(n9297) );
  AND4_X1 U10652 ( .A1(n9812), .A2(n9297), .A3(n9831), .A4(n9296), .ZN(n9298)
         );
  AND4_X1 U10653 ( .A1(n9765), .A2(n9795), .A3(n4327), .A4(n9298), .ZN(n9299)
         );
  AND3_X1 U10654 ( .A1(n9725), .A2(n9750), .A3(n9299), .ZN(n9300) );
  NAND4_X1 U10655 ( .A1(n9301), .A2(n9709), .A3(n9300), .A4(n9690), .ZN(n9302)
         );
  NOR2_X1 U10656 ( .A1(n9303), .A2(n9302), .ZN(n9304) );
  NOR2_X1 U10657 ( .A1(n9309), .A2(n9308), .ZN(n9310) );
  AND3_X1 U10658 ( .A1(n9310), .A2(n9411), .A3(n9351), .ZN(n9348) );
  NAND2_X1 U10659 ( .A1(n9312), .A2(n9311), .ZN(n9334) );
  INV_X1 U10660 ( .A(n9334), .ZN(n9402) );
  NAND2_X1 U10661 ( .A1(n9314), .A2(n9313), .ZN(n9315) );
  NAND2_X1 U10662 ( .A1(n9316), .A2(n9315), .ZN(n9317) );
  NAND2_X1 U10663 ( .A1(n9317), .A2(n9325), .ZN(n9318) );
  AND2_X1 U10664 ( .A1(n9319), .A2(n9318), .ZN(n9331) );
  INV_X1 U10665 ( .A(n9331), .ZN(n9321) );
  OR2_X1 U10666 ( .A1(n9321), .A2(n9320), .ZN(n9399) );
  OAI21_X1 U10667 ( .B1(n9399), .B2(n9727), .A(n9322), .ZN(n9335) );
  INV_X1 U10668 ( .A(n9323), .ZN(n9328) );
  INV_X1 U10669 ( .A(n9324), .ZN(n9326) );
  OAI211_X1 U10670 ( .C1(n9328), .C2(n9327), .A(n9326), .B(n9325), .ZN(n9330)
         );
  AOI21_X1 U10671 ( .B1(n9331), .B2(n9330), .A(n9329), .ZN(n9333) );
  OAI21_X1 U10672 ( .B1(n9334), .B2(n9333), .A(n9332), .ZN(n9360) );
  AOI21_X1 U10673 ( .B1(n9402), .B2(n9335), .A(n9360), .ZN(n9339) );
  NAND2_X1 U10674 ( .A1(n9337), .A2(n9336), .ZN(n9404) );
  OAI22_X1 U10675 ( .A1(n9339), .A2(n9404), .B1(n9601), .B2(n9338), .ZN(n9343)
         );
  NAND2_X1 U10676 ( .A1(n9341), .A2(n9340), .ZN(n9408) );
  OAI22_X1 U10677 ( .A1(n9343), .A2(n9408), .B1(n4796), .B2(n9342), .ZN(n9345)
         );
  INV_X1 U10678 ( .A(n9351), .ZN(n9410) );
  AOI211_X1 U10679 ( .C1(n9345), .C2(n9411), .A(n9344), .B(n9410), .ZN(n9346)
         );
  OAI21_X1 U10680 ( .B1(n9346), .B2(n9348), .A(n6665), .ZN(n9347) );
  INV_X1 U10681 ( .A(n9359), .ZN(n9415) );
  OAI21_X1 U10682 ( .B1(n9352), .B2(n9351), .A(n9350), .ZN(n9355) );
  NOR3_X1 U10683 ( .A1(n9359), .A2(n6666), .A3(n9353), .ZN(n9354) );
  OAI211_X1 U10684 ( .C1(n9411), .C2(n6665), .A(n9355), .B(n9354), .ZN(n9418)
         );
  NAND2_X1 U10685 ( .A1(n9357), .A2(n9356), .ZN(n9358) );
  OAI211_X1 U10686 ( .C1(n6666), .C2(n9359), .A(n9358), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9417) );
  INV_X1 U10687 ( .A(n9360), .ZN(n9406) );
  INV_X1 U10688 ( .A(n9361), .ZN(n9362) );
  OAI21_X1 U10689 ( .B1(n9364), .B2(n9363), .A(n9362), .ZN(n9365) );
  AOI211_X1 U10690 ( .C1(n10080), .C2(n6725), .A(n9366), .B(n9365), .ZN(n9370)
         );
  AND4_X1 U10691 ( .A1(n9370), .A2(n9369), .A3(n9368), .A4(n9367), .ZN(n9371)
         );
  NOR2_X1 U10692 ( .A1(n9372), .A2(n9371), .ZN(n9375) );
  OAI21_X1 U10693 ( .B1(n9375), .B2(n9374), .A(n9373), .ZN(n9378) );
  AOI21_X1 U10694 ( .B1(n9378), .B2(n9377), .A(n9376), .ZN(n9382) );
  INV_X1 U10695 ( .A(n9379), .ZN(n9381) );
  OAI211_X1 U10696 ( .C1(n9382), .C2(n9381), .A(n9380), .B(n9827), .ZN(n9384)
         );
  NAND3_X1 U10697 ( .A1(n9385), .A2(n9384), .A3(n4682), .ZN(n9393) );
  OAI21_X1 U10698 ( .B1(n9388), .B2(n9387), .A(n9386), .ZN(n9392) );
  INV_X1 U10699 ( .A(n9389), .ZN(n9391) );
  AOI211_X1 U10700 ( .C1(n9393), .C2(n9392), .A(n9391), .B(n9390), .ZN(n9398)
         );
  INV_X1 U10701 ( .A(n9394), .ZN(n9397) );
  OAI211_X1 U10702 ( .C1(n9398), .C2(n9397), .A(n9396), .B(n9395), .ZN(n9400)
         );
  AOI21_X1 U10703 ( .B1(n9401), .B2(n9400), .A(n9399), .ZN(n9403) );
  OAI21_X1 U10704 ( .B1(n9403), .B2(n4966), .A(n9402), .ZN(n9405) );
  AOI21_X1 U10705 ( .B1(n9406), .B2(n9405), .A(n9404), .ZN(n9409) );
  OAI21_X1 U10706 ( .B1(n9409), .B2(n9408), .A(n9407), .ZN(n9412) );
  AOI21_X1 U10707 ( .B1(n9412), .B2(n9411), .A(n9410), .ZN(n9413) );
  XNOR2_X1 U10708 ( .A(n9413), .B(n6665), .ZN(n9416) );
  MUX2_X1 U10709 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9419), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10710 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9420), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10711 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9421), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10712 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9637), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10713 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9627), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10714 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9673), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10715 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9688), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10716 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9714), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10717 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9687), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10718 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9752), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10719 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9768), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10720 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9776), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10721 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9767), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10722 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9815), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10723 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9833), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10724 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9814), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10725 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9835), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10726 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n4638), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10727 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9423), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10728 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9424), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10729 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9425), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10730 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9426), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10731 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9427), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10732 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9428), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10733 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9429), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10734 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9430), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10735 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9431), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10736 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6725), .S(P1_U3973), .Z(
        P1_U3555) );
  OAI211_X1 U10737 ( .C1(n9453), .C2(n9434), .A(n10052), .B(n9433), .ZN(n9442)
         );
  OAI211_X1 U10738 ( .C1(n9437), .C2(n9436), .A(n10061), .B(n9435), .ZN(n9441)
         );
  AOI22_X1 U10739 ( .A1(n10063), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9440) );
  NAND2_X1 U10740 ( .A1(n10054), .A2(n9438), .ZN(n9439) );
  NAND4_X1 U10741 ( .A1(n9442), .A2(n9441), .A3(n9440), .A4(n9439), .ZN(
        P1_U3244) );
  XOR2_X1 U10742 ( .A(n9444), .B(n9443), .Z(n9451) );
  INV_X1 U10743 ( .A(n9445), .ZN(n9449) );
  MUX2_X1 U10744 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n7047), .S(n9446), .Z(n9448)
         );
  INV_X1 U10745 ( .A(n9469), .ZN(n9447) );
  AOI211_X1 U10746 ( .C1(n9449), .C2(n9448), .A(n9447), .B(n9556), .ZN(n9450)
         );
  AOI21_X1 U10747 ( .B1(n10061), .B2(n9451), .A(n9450), .ZN(n9462) );
  AOI22_X1 U10748 ( .A1(n10063), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n9461) );
  MUX2_X1 U10749 ( .A(n9454), .B(n9453), .S(n9452), .Z(n9456) );
  NAND2_X1 U10750 ( .A1(n9456), .A2(n9455), .ZN(n9457) );
  OAI211_X1 U10751 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9458), .A(n9457), .B(
        P1_U3973), .ZN(n10068) );
  NAND2_X1 U10752 ( .A1(n10054), .A2(n9459), .ZN(n9460) );
  NAND4_X1 U10753 ( .A1(n9462), .A2(n9461), .A3(n10068), .A4(n9460), .ZN(
        P1_U3245) );
  INV_X1 U10754 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9464) );
  OAI21_X1 U10755 ( .B1(n9596), .B2(n9464), .A(n9463), .ZN(n9465) );
  AOI21_X1 U10756 ( .B1(n9466), .B2(n10054), .A(n9465), .ZN(n9476) );
  MUX2_X1 U10757 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n7668), .S(n9467), .Z(n9470)
         );
  NAND3_X1 U10758 ( .A1(n9470), .A2(n9469), .A3(n9468), .ZN(n9471) );
  NAND3_X1 U10759 ( .A1(n10052), .A2(n10049), .A3(n9471), .ZN(n9475) );
  OAI211_X1 U10760 ( .C1(n9473), .C2(n9472), .A(n10061), .B(n10058), .ZN(n9474) );
  NAND3_X1 U10761 ( .A1(n9476), .A2(n9475), .A3(n9474), .ZN(P1_U3246) );
  NOR2_X1 U10762 ( .A1(n9580), .A2(n9477), .ZN(n9478) );
  AOI211_X1 U10763 ( .C1(n10063), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n9479), .B(
        n9478), .ZN(n9492) );
  INV_X1 U10764 ( .A(n9480), .ZN(n10051) );
  INV_X1 U10765 ( .A(n9481), .ZN(n9484) );
  MUX2_X1 U10766 ( .A(n7054), .B(P1_REG2_REG_5__SCAN_IN), .S(n9482), .Z(n9483)
         );
  NAND3_X1 U10767 ( .A1(n10051), .A2(n9484), .A3(n9483), .ZN(n9485) );
  NAND3_X1 U10768 ( .A1(n10052), .A2(n9499), .A3(n9485), .ZN(n9491) );
  INV_X1 U10769 ( .A(n9486), .ZN(n9506) );
  NAND3_X1 U10770 ( .A1(n10060), .A2(n9488), .A3(n9487), .ZN(n9489) );
  NAND3_X1 U10771 ( .A1(n10061), .A2(n9506), .A3(n9489), .ZN(n9490) );
  NAND3_X1 U10772 ( .A1(n9492), .A2(n9491), .A3(n9490), .ZN(P1_U3248) );
  INV_X1 U10773 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9494) );
  OAI21_X1 U10774 ( .B1(n9596), .B2(n9494), .A(n9493), .ZN(n9495) );
  AOI21_X1 U10775 ( .B1(n9503), .B2(n10054), .A(n9495), .ZN(n9511) );
  INV_X1 U10776 ( .A(n9496), .ZN(n9501) );
  NAND3_X1 U10777 ( .A1(n9499), .A2(n9498), .A3(n9497), .ZN(n9500) );
  NAND3_X1 U10778 ( .A1(n10052), .A2(n9501), .A3(n9500), .ZN(n9510) );
  INV_X1 U10779 ( .A(n9502), .ZN(n9505) );
  MUX2_X1 U10780 ( .A(n10121), .B(P1_REG1_REG_6__SCAN_IN), .S(n9503), .Z(n9504) );
  NAND3_X1 U10781 ( .A1(n9506), .A2(n9505), .A3(n9504), .ZN(n9507) );
  NAND3_X1 U10782 ( .A1(n10061), .A2(n9508), .A3(n9507), .ZN(n9509) );
  NAND3_X1 U10783 ( .A1(n9511), .A2(n9510), .A3(n9509), .ZN(P1_U3249) );
  OAI211_X1 U10784 ( .C1(n9514), .C2(n9513), .A(n10052), .B(n9512), .ZN(n9525)
         );
  INV_X1 U10785 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9516) );
  OAI21_X1 U10786 ( .B1(n9596), .B2(n9516), .A(n9515), .ZN(n9517) );
  AOI21_X1 U10787 ( .B1(n9518), .B2(n10054), .A(n9517), .ZN(n9524) );
  OAI21_X1 U10788 ( .B1(n9521), .B2(n9520), .A(n9519), .ZN(n9522) );
  NAND3_X1 U10789 ( .A1(n4665), .A2(n10061), .A3(n9522), .ZN(n9523) );
  NAND3_X1 U10790 ( .A1(n9525), .A2(n9524), .A3(n9523), .ZN(P1_U3256) );
  AOI22_X1 U10791 ( .A1(n9527), .A2(n9533), .B1(P1_REG1_REG_15__SCAN_IN), .B2(
        n9526), .ZN(n9529) );
  NOR2_X1 U10792 ( .A1(n9535), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9544) );
  AOI21_X1 U10793 ( .B1(n9535), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9544), .ZN(
        n9528) );
  NOR2_X1 U10794 ( .A1(n9529), .A2(n9528), .ZN(n9530) );
  AND2_X1 U10795 ( .A1(n9529), .A2(n9528), .ZN(n9545) );
  OAI21_X1 U10796 ( .B1(n9530), .B2(n9545), .A(n10061), .ZN(n9543) );
  INV_X1 U10797 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10040) );
  OAI21_X1 U10798 ( .B1(n9596), .B2(n10040), .A(n9531), .ZN(n9532) );
  AOI21_X1 U10799 ( .B1(n9535), .B2(n10054), .A(n9532), .ZN(n9542) );
  NAND2_X1 U10800 ( .A1(n9534), .A2(n9533), .ZN(n9539) );
  INV_X1 U10801 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9536) );
  MUX2_X1 U10802 ( .A(n9536), .B(P1_REG2_REG_16__SCAN_IN), .S(n9535), .Z(n9537) );
  NAND3_X1 U10803 ( .A1(n9539), .A2(n9538), .A3(n9537), .ZN(n9540) );
  NAND3_X1 U10804 ( .A1(n9550), .A2(n10052), .A3(n9540), .ZN(n9541) );
  NAND3_X1 U10805 ( .A1(n9543), .A2(n9542), .A3(n9541), .ZN(P1_U3259) );
  NOR2_X1 U10806 ( .A1(n9545), .A2(n9544), .ZN(n9547) );
  XNOR2_X1 U10807 ( .A(n9568), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9546) );
  AOI21_X1 U10808 ( .B1(n9547), .B2(n9546), .A(n9565), .ZN(n9562) );
  INV_X1 U10809 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9549) );
  OAI21_X1 U10810 ( .B1(n9596), .B2(n9549), .A(n9548), .ZN(n9559) );
  INV_X1 U10811 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9552) );
  AOI22_X1 U10812 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9553), .B1(n9568), .B2(
        n9552), .ZN(n9554) );
  AOI21_X1 U10813 ( .B1(n9555), .B2(n9554), .A(n9569), .ZN(n9557) );
  NOR2_X1 U10814 ( .A1(n9557), .A2(n9556), .ZN(n9558) );
  AOI211_X1 U10815 ( .C1(n10054), .C2(n9568), .A(n9559), .B(n9558), .ZN(n9560)
         );
  OAI21_X1 U10816 ( .B1(n9562), .B2(n9561), .A(n9560), .ZN(P1_U3260) );
  NOR2_X1 U10817 ( .A1(n9568), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9564) );
  XNOR2_X1 U10818 ( .A(n9583), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9563) );
  INV_X1 U10819 ( .A(n9581), .ZN(n9567) );
  OAI21_X1 U10820 ( .B1(n9565), .B2(n9564), .A(n9563), .ZN(n9566) );
  NAND3_X1 U10821 ( .A1(n9567), .A2(n10061), .A3(n9566), .ZN(n9578) );
  NOR2_X1 U10822 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9568), .ZN(n9570) );
  XNOR2_X1 U10823 ( .A(n9583), .B(n9571), .ZN(n9572) );
  OAI211_X1 U10824 ( .C1(n9573), .C2(n9572), .A(n10052), .B(n9585), .ZN(n9574)
         );
  NAND2_X1 U10825 ( .A1(n9575), .A2(n9574), .ZN(n9576) );
  AOI21_X1 U10826 ( .B1(n10063), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n9576), .ZN(
        n9577) );
  OAI211_X1 U10827 ( .C1(n9580), .C2(n9579), .A(n9578), .B(n9577), .ZN(
        P1_U3261) );
  AOI21_X1 U10828 ( .B1(n9583), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9581), .ZN(
        n9582) );
  XOR2_X1 U10829 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9582), .Z(n9591) );
  INV_X1 U10830 ( .A(n9591), .ZN(n9587) );
  NAND2_X1 U10831 ( .A1(n9583), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9584) );
  NAND2_X1 U10832 ( .A1(n9585), .A2(n9584), .ZN(n9586) );
  XNOR2_X1 U10833 ( .A(n9586), .B(n6530), .ZN(n9589) );
  AOI22_X1 U10834 ( .A1(n9587), .A2(n10061), .B1(n10052), .B2(n9589), .ZN(
        n9593) );
  NOR3_X1 U10835 ( .A1(n9589), .A2(n9588), .A3(n9999), .ZN(n9590) );
  AOI211_X1 U10836 ( .C1(n9591), .C2(n10061), .A(n9590), .B(n10054), .ZN(n9592) );
  MUX2_X1 U10837 ( .A(n9593), .B(n9592), .S(n9677), .Z(n9595) );
  OAI211_X1 U10838 ( .C1(n4604), .C2(n9596), .A(n9595), .B(n9594), .ZN(
        P1_U3262) );
  NAND2_X1 U10839 ( .A1(n9597), .A2(n9756), .ZN(n9600) );
  NOR2_X1 U10840 ( .A1(n10077), .A2(n9598), .ZN(n9603) );
  AOI21_X1 U10841 ( .B1(n10077), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9603), .ZN(
        n9599) );
  OAI211_X1 U10842 ( .C1(n5166), .C2(n10081), .A(n9600), .B(n9599), .ZN(
        P1_U3263) );
  NOR2_X1 U10843 ( .A1(n9601), .A2(n10081), .ZN(n9602) );
  AOI211_X1 U10844 ( .C1(n10077), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9603), .B(
        n9602), .ZN(n9604) );
  OAI21_X1 U10845 ( .B1(n10075), .B2(n9605), .A(n9604), .ZN(P1_U3264) );
  INV_X1 U10846 ( .A(n9853), .ZN(n9613) );
  INV_X1 U10847 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9606) );
  OAI22_X1 U10848 ( .A1(n9607), .A2(n10072), .B1(n9606), .B2(n9848), .ZN(n9608) );
  AOI21_X1 U10849 ( .B1(n9609), .B2(n9819), .A(n9608), .ZN(n9610) );
  OAI21_X1 U10850 ( .B1(n9611), .B2(n10075), .A(n9610), .ZN(n9612) );
  AOI21_X1 U10851 ( .B1(n9613), .B2(n9700), .A(n9612), .ZN(n9614) );
  OAI21_X1 U10852 ( .B1(n10077), .B2(n9615), .A(n9614), .ZN(P1_U3266) );
  NOR2_X1 U10853 ( .A1(n4315), .A2(n9621), .ZN(n9618) );
  INV_X1 U10854 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9620) );
  OAI22_X1 U10855 ( .A1(n9621), .A2(n10081), .B1(n9620), .B2(n9848), .ZN(n9622) );
  AOI21_X1 U10856 ( .B1(n5181), .B2(n9756), .A(n9622), .ZN(n9632) );
  INV_X1 U10857 ( .A(n9623), .ZN(n9629) );
  OAI21_X1 U10858 ( .B1(n9629), .B2(n10072), .A(n9857), .ZN(n9630) );
  NAND2_X1 U10859 ( .A1(n9630), .A2(n9848), .ZN(n9631) );
  OAI211_X1 U10860 ( .C1(n9858), .C2(n9850), .A(n9632), .B(n9631), .ZN(
        P1_U3267) );
  XNOR2_X1 U10861 ( .A(n9633), .B(n9636), .ZN(n9938) );
  OAI21_X1 U10862 ( .B1(n9636), .B2(n9635), .A(n9634), .ZN(n9638) );
  AOI222_X1 U10863 ( .A1(n9829), .A2(n9638), .B1(n9637), .B2(n9834), .C1(n9673), .C2(n9836), .ZN(n9860) );
  INV_X1 U10864 ( .A(n9860), .ZN(n9647) );
  NAND2_X1 U10865 ( .A1(n9656), .A2(n9644), .ZN(n9639) );
  NAND2_X1 U10866 ( .A1(n9639), .A2(n9894), .ZN(n9640) );
  OR2_X1 U10867 ( .A1(n4315), .A2(n9640), .ZN(n9859) );
  INV_X1 U10868 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9641) );
  OAI22_X1 U10869 ( .A1(n9642), .A2(n10072), .B1(n9641), .B2(n9848), .ZN(n9643) );
  AOI21_X1 U10870 ( .B1(n9644), .B2(n9819), .A(n9643), .ZN(n9645) );
  OAI21_X1 U10871 ( .B1(n9859), .B2(n10075), .A(n9645), .ZN(n9646) );
  AOI21_X1 U10872 ( .B1(n9647), .B2(n9848), .A(n9646), .ZN(n9648) );
  OAI21_X1 U10873 ( .B1(n9938), .B2(n9850), .A(n9648), .ZN(P1_U3268) );
  NOR2_X1 U10874 ( .A1(n9668), .A2(n9649), .ZN(n9650) );
  XNOR2_X1 U10875 ( .A(n9650), .B(n4976), .ZN(n9651) );
  OAI222_X1 U10876 ( .A1(n9802), .A2(n9653), .B1(n9800), .B2(n9652), .C1(n9651), .C2(n9797), .ZN(n9866) );
  NAND2_X1 U10877 ( .A1(n9654), .A2(n9660), .ZN(n9655) );
  NAND2_X1 U10878 ( .A1(n9656), .A2(n9655), .ZN(n9863) );
  INV_X1 U10879 ( .A(n9756), .ZN(n9662) );
  INV_X1 U10880 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9657) );
  OAI22_X1 U10881 ( .A1(n9658), .A2(n10072), .B1(n9848), .B2(n9657), .ZN(n9659) );
  AOI21_X1 U10882 ( .B1(n9660), .B2(n9819), .A(n9659), .ZN(n9661) );
  OAI21_X1 U10883 ( .B1(n9863), .B2(n9662), .A(n9661), .ZN(n9665) );
  XNOR2_X1 U10884 ( .A(n9663), .B(n4976), .ZN(n9865) );
  NOR2_X1 U10885 ( .A1(n9865), .A2(n9850), .ZN(n9664) );
  AOI211_X1 U10886 ( .C1(n9848), .C2(n9866), .A(n9665), .B(n9664), .ZN(n9666)
         );
  INV_X1 U10887 ( .A(n9666), .ZN(P1_U3269) );
  XNOR2_X1 U10888 ( .A(n9667), .B(n9669), .ZN(n9950) );
  INV_X1 U10889 ( .A(n9668), .ZN(n9672) );
  NAND3_X1 U10890 ( .A1(n9685), .A2(n9670), .A3(n9669), .ZN(n9671) );
  NAND2_X1 U10891 ( .A1(n9672), .A2(n9671), .ZN(n9674) );
  AOI222_X1 U10892 ( .A1(n9829), .A2(n9674), .B1(n9673), .B2(n9834), .C1(n9714), .C2(n9836), .ZN(n9871) );
  INV_X1 U10893 ( .A(n9871), .ZN(n9679) );
  OAI211_X1 U10894 ( .C1(n9693), .C2(n9675), .A(n9894), .B(n9654), .ZN(n9870)
         );
  OAI22_X1 U10895 ( .A1(n9870), .A2(n9677), .B1(n10072), .B2(n9676), .ZN(n9678) );
  OAI21_X1 U10896 ( .B1(n9679), .B2(n9678), .A(n9848), .ZN(n9681) );
  AOI22_X1 U10897 ( .A1(n9947), .A2(n9819), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n10077), .ZN(n9680) );
  OAI211_X1 U10898 ( .C1(n9950), .C2(n9850), .A(n9681), .B(n9680), .ZN(
        P1_U3270) );
  INV_X1 U10899 ( .A(n9690), .ZN(n9684) );
  NAND2_X1 U10900 ( .A1(n9684), .A2(n9683), .ZN(n9686) );
  OAI21_X1 U10901 ( .B1(n9712), .B2(n9686), .A(n9685), .ZN(n9689) );
  AOI222_X1 U10902 ( .A1(n9829), .A2(n9689), .B1(n9688), .B2(n9834), .C1(n9687), .C2(n9836), .ZN(n9879) );
  XNOR2_X1 U10903 ( .A(n9691), .B(n9690), .ZN(n9880) );
  INV_X1 U10904 ( .A(n9880), .ZN(n9701) );
  OAI21_X1 U10905 ( .B1(n9717), .B2(n9692), .A(n9894), .ZN(n9694) );
  OR2_X1 U10906 ( .A1(n9694), .A2(n9693), .ZN(n9875) );
  INV_X1 U10907 ( .A(n9695), .ZN(n9696) );
  AOI22_X1 U10908 ( .A1(n9696), .A2(n9842), .B1(n10077), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9698) );
  NAND2_X1 U10909 ( .A1(n9877), .A2(n9819), .ZN(n9697) );
  OAI211_X1 U10910 ( .C1(n9875), .C2(n10075), .A(n9698), .B(n9697), .ZN(n9699)
         );
  AOI21_X1 U10911 ( .B1(n9701), .B2(n9700), .A(n9699), .ZN(n9702) );
  OAI21_X1 U10912 ( .B1(n10077), .B2(n9879), .A(n9702), .ZN(P1_U3271) );
  NAND2_X1 U10913 ( .A1(n9704), .A2(n9703), .ZN(n9724) );
  INV_X1 U10914 ( .A(n9705), .ZN(n9707) );
  OAI21_X1 U10915 ( .B1(n9724), .B2(n9707), .A(n9706), .ZN(n9708) );
  XOR2_X1 U10916 ( .A(n9709), .B(n9708), .Z(n9958) );
  NOR2_X1 U10917 ( .A1(n9710), .A2(n9709), .ZN(n9711) );
  OR2_X1 U10918 ( .A1(n9712), .A2(n9711), .ZN(n9713) );
  NAND2_X1 U10919 ( .A1(n9713), .A2(n9829), .ZN(n9716) );
  AOI22_X1 U10920 ( .A1(n9714), .A2(n9834), .B1(n9836), .B2(n9752), .ZN(n9715)
         );
  NAND2_X1 U10921 ( .A1(n9716), .A2(n9715), .ZN(n9882) );
  AOI211_X1 U10922 ( .C1(n9955), .C2(n5185), .A(n9864), .B(n9717), .ZN(n9881)
         );
  NAND2_X1 U10923 ( .A1(n9881), .A2(n9841), .ZN(n9720) );
  AOI22_X1 U10924 ( .A1(n10077), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9718), 
        .B2(n9842), .ZN(n9719) );
  OAI211_X1 U10925 ( .C1(n9721), .C2(n10081), .A(n9720), .B(n9719), .ZN(n9722)
         );
  AOI21_X1 U10926 ( .B1(n9882), .B2(n9848), .A(n9722), .ZN(n9723) );
  OAI21_X1 U10927 ( .B1(n9958), .B2(n9850), .A(n9723), .ZN(P1_U3272) );
  XNOR2_X1 U10928 ( .A(n9724), .B(n9725), .ZN(n9962) );
  INV_X1 U10929 ( .A(n9725), .ZN(n9726) );
  XNOR2_X1 U10930 ( .A(n9727), .B(n9726), .ZN(n9731) );
  OAI22_X1 U10931 ( .A1(n9729), .A2(n9802), .B1(n9728), .B2(n9800), .ZN(n9730)
         );
  AOI21_X1 U10932 ( .B1(n9731), .B2(n9829), .A(n9730), .ZN(n9888) );
  INV_X1 U10933 ( .A(n9888), .ZN(n9738) );
  INV_X1 U10934 ( .A(n9732), .ZN(n9745) );
  INV_X1 U10935 ( .A(n9734), .ZN(n9889) );
  OAI211_X1 U10936 ( .C1(n9745), .C2(n9889), .A(n5185), .B(n9894), .ZN(n9887)
         );
  AOI22_X1 U10937 ( .A1(n10077), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9733), 
        .B2(n9842), .ZN(n9736) );
  NAND2_X1 U10938 ( .A1(n9734), .A2(n9819), .ZN(n9735) );
  OAI211_X1 U10939 ( .C1(n9887), .C2(n10075), .A(n9736), .B(n9735), .ZN(n9737)
         );
  AOI21_X1 U10940 ( .B1(n9738), .B2(n9848), .A(n9737), .ZN(n9739) );
  OAI21_X1 U10941 ( .B1(n9962), .B2(n9850), .A(n9739), .ZN(P1_U3273) );
  AOI22_X1 U10942 ( .A1(n9758), .A2(n9742), .B1(n9776), .B2(n9900), .ZN(n9743)
         );
  XNOR2_X1 U10943 ( .A(n9743), .B(n9750), .ZN(n9898) );
  INV_X1 U10944 ( .A(n9744), .ZN(n9746) );
  AOI21_X1 U10945 ( .B1(n9893), .B2(n9746), .A(n9745), .ZN(n9895) );
  AOI22_X1 U10946 ( .A1(n10077), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9747), 
        .B2(n9842), .ZN(n9748) );
  OAI21_X1 U10947 ( .B1(n9749), .B2(n10081), .A(n9748), .ZN(n9755) );
  XNOR2_X1 U10948 ( .A(n9751), .B(n9750), .ZN(n9753) );
  AOI222_X1 U10949 ( .A1(n9829), .A2(n9753), .B1(n9752), .B2(n9834), .C1(n9776), .C2(n9836), .ZN(n9897) );
  NOR2_X1 U10950 ( .A1(n9897), .A2(n10077), .ZN(n9754) );
  AOI211_X1 U10951 ( .C1(n9895), .C2(n9756), .A(n9755), .B(n9754), .ZN(n9757)
         );
  OAI21_X1 U10952 ( .B1(n9898), .B2(n9850), .A(n9757), .ZN(P1_U3274) );
  XOR2_X1 U10953 ( .A(n9765), .B(n9758), .Z(n9903) );
  INV_X1 U10954 ( .A(n9779), .ZN(n9759) );
  AOI211_X1 U10955 ( .C1(n9900), .C2(n9759), .A(n9864), .B(n9744), .ZN(n9899)
         );
  INV_X1 U10956 ( .A(n9760), .ZN(n9761) );
  AOI22_X1 U10957 ( .A1(n10077), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9761), 
        .B2(n9842), .ZN(n9762) );
  OAI21_X1 U10958 ( .B1(n9763), .B2(n10081), .A(n9762), .ZN(n9771) );
  OAI21_X1 U10959 ( .B1(n9766), .B2(n9765), .A(n9764), .ZN(n9769) );
  AOI222_X1 U10960 ( .A1(n9829), .A2(n9769), .B1(n9768), .B2(n9834), .C1(n9767), .C2(n9836), .ZN(n9902) );
  NOR2_X1 U10961 ( .A1(n9902), .A2(n10077), .ZN(n9770) );
  AOI211_X1 U10962 ( .C1(n9899), .C2(n9841), .A(n9771), .B(n9770), .ZN(n9772)
         );
  OAI21_X1 U10963 ( .B1(n9903), .B2(n9850), .A(n9772), .ZN(P1_U3275) );
  XNOR2_X1 U10964 ( .A(n9773), .B(n4327), .ZN(n9967) );
  OAI211_X1 U10965 ( .C1(n9774), .C2(n4327), .A(n9829), .B(n9775), .ZN(n9778)
         );
  AOI22_X1 U10966 ( .A1(n9776), .A2(n9834), .B1(n9836), .B2(n9815), .ZN(n9777)
         );
  NAND2_X1 U10967 ( .A1(n9778), .A2(n9777), .ZN(n9904) );
  AOI211_X1 U10968 ( .C1(n9906), .C2(n9789), .A(n9864), .B(n9779), .ZN(n9905)
         );
  NAND2_X1 U10969 ( .A1(n9905), .A2(n9841), .ZN(n9782) );
  AOI22_X1 U10970 ( .A1(n10077), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9780), 
        .B2(n9842), .ZN(n9781) );
  OAI211_X1 U10971 ( .C1(n9783), .C2(n10081), .A(n9782), .B(n9781), .ZN(n9784)
         );
  AOI21_X1 U10972 ( .B1(n9904), .B2(n9848), .A(n9784), .ZN(n9785) );
  OAI21_X1 U10973 ( .B1(n9967), .B2(n9850), .A(n9785), .ZN(P1_U3276) );
  AOI21_X1 U10974 ( .B1(n9795), .B2(n9786), .A(n4395), .ZN(n9787) );
  INV_X1 U10975 ( .A(n9787), .ZN(n9971) );
  INV_X1 U10976 ( .A(n9789), .ZN(n9790) );
  AOI211_X1 U10977 ( .C1(n9911), .C2(n9788), .A(n9864), .B(n9790), .ZN(n9910)
         );
  INV_X1 U10978 ( .A(n9911), .ZN(n9791) );
  NOR2_X1 U10979 ( .A1(n9791), .A2(n10081), .ZN(n9794) );
  OAI22_X1 U10980 ( .A1(n9848), .A2(n9536), .B1(n9792), .B2(n10072), .ZN(n9793) );
  AOI211_X1 U10981 ( .C1(n9910), .C2(n9841), .A(n9794), .B(n9793), .ZN(n9804)
         );
  XOR2_X1 U10982 ( .A(n9796), .B(n9795), .Z(n9798) );
  OAI222_X1 U10983 ( .A1(n9802), .A2(n9801), .B1(n9800), .B2(n9799), .C1(n9798), .C2(n9797), .ZN(n9909) );
  NAND2_X1 U10984 ( .A1(n9909), .A2(n9848), .ZN(n9803) );
  OAI211_X1 U10985 ( .C1(n9971), .C2(n9850), .A(n9804), .B(n9803), .ZN(
        P1_U3277) );
  AND2_X1 U10986 ( .A1(n9806), .A2(n9805), .ZN(n9826) );
  OAI22_X1 U10987 ( .A1(n9826), .A2(n9808), .B1(n9807), .B2(n9846), .ZN(n9809)
         );
  XOR2_X1 U10988 ( .A(n9812), .B(n9809), .Z(n9917) );
  AND2_X1 U10989 ( .A1(n9830), .A2(n9810), .ZN(n9813) );
  OAI21_X1 U10990 ( .B1(n9813), .B2(n9812), .A(n9811), .ZN(n9816) );
  AOI222_X1 U10991 ( .A1(n9829), .A2(n9816), .B1(n9815), .B2(n9834), .C1(n9814), .C2(n9836), .ZN(n9915) );
  INV_X1 U10992 ( .A(n9915), .ZN(n9824) );
  OAI211_X1 U10993 ( .C1(n9839), .C2(n9976), .A(n9894), .B(n9788), .ZN(n9914)
         );
  AOI22_X1 U10994 ( .A1(n10077), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9818), 
        .B2(n9842), .ZN(n9822) );
  NAND2_X1 U10995 ( .A1(n9820), .A2(n9819), .ZN(n9821) );
  OAI211_X1 U10996 ( .C1(n9914), .C2(n10075), .A(n9822), .B(n9821), .ZN(n9823)
         );
  AOI21_X1 U10997 ( .B1(n9824), .B2(n9848), .A(n9823), .ZN(n9825) );
  OAI21_X1 U10998 ( .B1(n9917), .B2(n9850), .A(n9825), .ZN(P1_U3278) );
  XNOR2_X1 U10999 ( .A(n9826), .B(n9831), .ZN(n9981) );
  AND2_X1 U11000 ( .A1(n9828), .A2(n9827), .ZN(n9832) );
  OAI211_X1 U11001 ( .C1(n9832), .C2(n9831), .A(n9830), .B(n9829), .ZN(n9838)
         );
  AOI22_X1 U11002 ( .A1(n9836), .A2(n9835), .B1(n9834), .B2(n9833), .ZN(n9837)
         );
  NAND2_X1 U11003 ( .A1(n9838), .A2(n9837), .ZN(n9922) );
  AOI211_X1 U11004 ( .C1(n9924), .C2(n9840), .A(n9864), .B(n9839), .ZN(n9923)
         );
  NAND2_X1 U11005 ( .A1(n9923), .A2(n9841), .ZN(n9845) );
  AOI22_X1 U11006 ( .A1(n10077), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9843), 
        .B2(n9842), .ZN(n9844) );
  OAI211_X1 U11007 ( .C1(n9846), .C2(n10081), .A(n9845), .B(n9844), .ZN(n9847)
         );
  AOI21_X1 U11008 ( .B1(n9848), .B2(n9922), .A(n9847), .ZN(n9849) );
  OAI21_X1 U11009 ( .B1(n9981), .B2(n9850), .A(n9849), .ZN(P1_U3279) );
  AOI22_X1 U11010 ( .A1(n5181), .A2(n9894), .B1(n9930), .B2(n9855), .ZN(n9856)
         );
  OAI211_X1 U11011 ( .C1(n9858), .C2(n9916), .A(n9857), .B(n9856), .ZN(n9936)
         );
  MUX2_X1 U11012 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9936), .S(n10123), .Z(
        P1_U3548) );
  NAND2_X1 U11013 ( .A1(n9860), .A2(n9859), .ZN(n9937) );
  MUX2_X1 U11014 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9937), .S(n10123), .Z(
        n9862) );
  OAI22_X1 U11015 ( .A1(n9938), .A2(n9927), .B1(n5150), .B2(n9921), .ZN(n9861)
         );
  OR2_X1 U11016 ( .A1(n9862), .A2(n9861), .ZN(P1_U3547) );
  OAI22_X1 U11017 ( .A1(n9865), .A2(n9916), .B1(n9864), .B2(n9863), .ZN(n9867)
         );
  NOR2_X1 U11018 ( .A1(n9867), .A2(n9866), .ZN(n9941) );
  MUX2_X1 U11019 ( .A(n9868), .B(n9941), .S(n10123), .Z(n9869) );
  OAI21_X1 U11020 ( .B1(n9944), .B2(n9921), .A(n9869), .ZN(P1_U3546) );
  AND2_X1 U11021 ( .A1(n9871), .A2(n9870), .ZN(n9945) );
  MUX2_X1 U11022 ( .A(n9872), .B(n9945), .S(n10123), .Z(n9874) );
  NAND2_X1 U11023 ( .A1(n9947), .A2(n9884), .ZN(n9873) );
  OAI211_X1 U11024 ( .C1(n9950), .C2(n9927), .A(n9874), .B(n9873), .ZN(
        P1_U3545) );
  INV_X1 U11025 ( .A(n9875), .ZN(n9876) );
  AOI21_X1 U11026 ( .B1(n9930), .B2(n9877), .A(n9876), .ZN(n9878) );
  OAI211_X1 U11027 ( .C1(n9880), .C2(n9916), .A(n9879), .B(n9878), .ZN(n9951)
         );
  MUX2_X1 U11028 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9951), .S(n10123), .Z(
        P1_U3544) );
  INV_X1 U11029 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9883) );
  NOR2_X1 U11030 ( .A1(n9882), .A2(n9881), .ZN(n9952) );
  MUX2_X1 U11031 ( .A(n9883), .B(n9952), .S(n10123), .Z(n9886) );
  NAND2_X1 U11032 ( .A1(n9955), .A2(n9884), .ZN(n9885) );
  OAI211_X1 U11033 ( .C1(n9958), .C2(n9927), .A(n9886), .B(n9885), .ZN(
        P1_U3543) );
  OAI211_X1 U11034 ( .C1(n9889), .C2(n10107), .A(n9888), .B(n9887), .ZN(n9890)
         );
  INV_X1 U11035 ( .A(n9890), .ZN(n9959) );
  MUX2_X1 U11036 ( .A(n9891), .B(n9959), .S(n10123), .Z(n9892) );
  OAI21_X1 U11037 ( .B1(n9962), .B2(n9927), .A(n9892), .ZN(P1_U3542) );
  AOI22_X1 U11038 ( .A1(n9895), .A2(n9894), .B1(n9930), .B2(n9893), .ZN(n9896)
         );
  OAI211_X1 U11039 ( .C1(n9898), .C2(n9916), .A(n9897), .B(n9896), .ZN(n9963)
         );
  MUX2_X1 U11040 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9963), .S(n10123), .Z(
        P1_U3541) );
  AOI21_X1 U11041 ( .B1(n9930), .B2(n9900), .A(n9899), .ZN(n9901) );
  OAI211_X1 U11042 ( .C1(n9903), .C2(n9916), .A(n9902), .B(n9901), .ZN(n9964)
         );
  MUX2_X1 U11043 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9964), .S(n10123), .Z(
        P1_U3540) );
  INV_X1 U11044 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9907) );
  AOI211_X1 U11045 ( .C1(n9930), .C2(n9906), .A(n9905), .B(n9904), .ZN(n9965)
         );
  MUX2_X1 U11046 ( .A(n9907), .B(n9965), .S(n10123), .Z(n9908) );
  OAI21_X1 U11047 ( .B1(n9967), .B2(n9927), .A(n9908), .ZN(P1_U3539) );
  INV_X1 U11048 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9912) );
  AOI211_X1 U11049 ( .C1(n9930), .C2(n9911), .A(n9910), .B(n9909), .ZN(n9968)
         );
  MUX2_X1 U11050 ( .A(n9912), .B(n9968), .S(n10123), .Z(n9913) );
  OAI21_X1 U11051 ( .B1(n9971), .B2(n9927), .A(n9913), .ZN(P1_U3538) );
  INV_X1 U11052 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9919) );
  OAI211_X1 U11053 ( .C1(n9917), .C2(n9916), .A(n9915), .B(n9914), .ZN(n9918)
         );
  INV_X1 U11054 ( .A(n9918), .ZN(n9972) );
  MUX2_X1 U11055 ( .A(n9919), .B(n9972), .S(n10123), .Z(n9920) );
  OAI21_X1 U11056 ( .B1(n9976), .B2(n9921), .A(n9920), .ZN(P1_U3537) );
  AOI211_X1 U11057 ( .C1(n9930), .C2(n9924), .A(n9923), .B(n9922), .ZN(n9977)
         );
  MUX2_X1 U11058 ( .A(n9925), .B(n9977), .S(n10123), .Z(n9926) );
  OAI21_X1 U11059 ( .B1(n9981), .B2(n9927), .A(n9926), .ZN(P1_U3536) );
  INV_X1 U11060 ( .A(n9928), .ZN(n9934) );
  AOI21_X1 U11061 ( .B1(n9930), .B2(n6484), .A(n9929), .ZN(n9931) );
  OAI211_X1 U11062 ( .C1(n9934), .C2(n9933), .A(n9932), .B(n9931), .ZN(n9982)
         );
  MUX2_X1 U11063 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9982), .S(n10123), .Z(
        P1_U3533) );
  MUX2_X1 U11064 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9935), .S(n10123), .Z(
        P1_U3522) );
  MUX2_X1 U11065 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9936), .S(n10115), .Z(
        P1_U3516) );
  MUX2_X1 U11066 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9937), .S(n10115), .Z(
        n9940) );
  OAI22_X1 U11067 ( .A1(n9938), .A2(n9980), .B1(n5150), .B2(n9975), .ZN(n9939)
         );
  OR2_X1 U11068 ( .A1(n9940), .A2(n9939), .ZN(P1_U3515) );
  INV_X1 U11069 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9942) );
  MUX2_X1 U11070 ( .A(n9942), .B(n9941), .S(n10115), .Z(n9943) );
  OAI21_X1 U11071 ( .B1(n9944), .B2(n9975), .A(n9943), .ZN(P1_U3514) );
  INV_X1 U11072 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9946) );
  MUX2_X1 U11073 ( .A(n9946), .B(n9945), .S(n10115), .Z(n9949) );
  NAND2_X1 U11074 ( .A1(n9947), .A2(n9954), .ZN(n9948) );
  OAI211_X1 U11075 ( .C1(n9950), .C2(n9980), .A(n9949), .B(n9948), .ZN(
        P1_U3513) );
  MUX2_X1 U11076 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9951), .S(n10115), .Z(
        P1_U3512) );
  INV_X1 U11077 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9953) );
  MUX2_X1 U11078 ( .A(n9953), .B(n9952), .S(n10115), .Z(n9957) );
  NAND2_X1 U11079 ( .A1(n9955), .A2(n9954), .ZN(n9956) );
  OAI211_X1 U11080 ( .C1(n9958), .C2(n9980), .A(n9957), .B(n9956), .ZN(
        P1_U3511) );
  INV_X1 U11081 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9960) );
  MUX2_X1 U11082 ( .A(n9960), .B(n9959), .S(n10115), .Z(n9961) );
  OAI21_X1 U11083 ( .B1(n9962), .B2(n9980), .A(n9961), .ZN(P1_U3510) );
  MUX2_X1 U11084 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9963), .S(n10115), .Z(
        P1_U3509) );
  MUX2_X1 U11085 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9964), .S(n10115), .Z(
        P1_U3507) );
  INV_X1 U11086 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10261) );
  MUX2_X1 U11087 ( .A(n10261), .B(n9965), .S(n10115), .Z(n9966) );
  OAI21_X1 U11088 ( .B1(n9967), .B2(n9980), .A(n9966), .ZN(P1_U3504) );
  INV_X1 U11089 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9969) );
  MUX2_X1 U11090 ( .A(n9969), .B(n9968), .S(n10115), .Z(n9970) );
  OAI21_X1 U11091 ( .B1(n9971), .B2(n9980), .A(n9970), .ZN(P1_U3501) );
  INV_X1 U11092 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9973) );
  MUX2_X1 U11093 ( .A(n9973), .B(n9972), .S(n10115), .Z(n9974) );
  OAI21_X1 U11094 ( .B1(n9976), .B2(n9975), .A(n9974), .ZN(P1_U3498) );
  INV_X1 U11095 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9978) );
  MUX2_X1 U11096 ( .A(n9978), .B(n9977), .S(n10115), .Z(n9979) );
  OAI21_X1 U11097 ( .B1(n9981), .B2(n9980), .A(n9979), .ZN(P1_U3495) );
  MUX2_X1 U11098 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n9982), .S(n10115), .Z(
        P1_U3486) );
  MUX2_X1 U11099 ( .A(P1_D_REG_1__SCAN_IN), .B(n9984), .S(n10086), .Z(P1_U3440) );
  MUX2_X1 U11100 ( .A(P1_D_REG_0__SCAN_IN), .B(n9986), .S(n9985), .Z(P1_U3439)
         );
  NAND2_X1 U11101 ( .A1(n9988), .A2(n9987), .ZN(n9992) );
  NAND4_X1 U11102 ( .A1(n9990), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .A4(n9989), .ZN(n9991) );
  OAI211_X1 U11103 ( .C1(n9994), .C2(n9993), .A(n9992), .B(n9991), .ZN(
        P1_U3324) );
  OAI222_X1 U11104 ( .A1(n10002), .A2(n9997), .B1(P1_U3086), .B2(n9996), .C1(
        n8589), .C2(n9995), .ZN(P1_U3326) );
  OAI222_X1 U11105 ( .A1(n10002), .A2(n10001), .B1(P1_U3086), .B2(n9999), .C1(
        n8589), .C2(n9998), .ZN(P1_U3328) );
  MUX2_X1 U11106 ( .A(n10003), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U11107 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10043) );
  INV_X1 U11108 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10041) );
  NOR2_X1 U11109 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10038) );
  NOR2_X1 U11110 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10034) );
  NOR2_X1 U11111 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10032) );
  INV_X1 U11112 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10029) );
  NOR2_X1 U11113 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10025) );
  NOR2_X1 U11114 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10021) );
  INV_X1 U11115 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10019) );
  NOR2_X1 U11116 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10017) );
  NOR2_X1 U11117 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10015) );
  NOR2_X1 U11118 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10013) );
  NOR2_X1 U11119 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10011) );
  NAND2_X1 U11120 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10009) );
  XOR2_X1 U11121 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10391) );
  NAND2_X1 U11122 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n10007) );
  AOI21_X1 U11123 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10201) );
  INV_X1 U11124 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10296) );
  NAND2_X1 U11125 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n10004) );
  NOR2_X1 U11126 ( .A1(n10296), .A2(n10004), .ZN(n10200) );
  NOR2_X1 U11127 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10200), .ZN(n10005) );
  NOR2_X1 U11128 ( .A1(n10201), .A2(n10005), .ZN(n10389) );
  XOR2_X1 U11129 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10388) );
  NAND2_X1 U11130 ( .A1(n10389), .A2(n10388), .ZN(n10006) );
  NAND2_X1 U11131 ( .A1(n10007), .A2(n10006), .ZN(n10390) );
  NAND2_X1 U11132 ( .A1(n10391), .A2(n10390), .ZN(n10008) );
  NAND2_X1 U11133 ( .A1(n10009), .A2(n10008), .ZN(n10393) );
  XNOR2_X1 U11134 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10392) );
  NOR2_X1 U11135 ( .A1(n10393), .A2(n10392), .ZN(n10010) );
  NOR2_X1 U11136 ( .A1(n10011), .A2(n10010), .ZN(n10381) );
  XNOR2_X1 U11137 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10380) );
  NOR2_X1 U11138 ( .A1(n10381), .A2(n10380), .ZN(n10012) );
  NOR2_X1 U11139 ( .A1(n10013), .A2(n10012), .ZN(n10379) );
  XNOR2_X1 U11140 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10378) );
  NOR2_X1 U11141 ( .A1(n10379), .A2(n10378), .ZN(n10014) );
  XNOR2_X1 U11142 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10384) );
  NOR2_X1 U11143 ( .A1(n10385), .A2(n10384), .ZN(n10016) );
  AOI22_X1 U11144 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10294), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n10019), .ZN(n10386) );
  NOR2_X1 U11145 ( .A1(n10387), .A2(n10386), .ZN(n10018) );
  AOI22_X1 U11146 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7090), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n10337), .ZN(n10382) );
  NOR2_X1 U11147 ( .A1(n10383), .A2(n10382), .ZN(n10020) );
  INV_X1 U11148 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10022) );
  AOI22_X1 U11149 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n10023), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n10022), .ZN(n10221) );
  AOI22_X1 U11150 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n10286), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n10027), .ZN(n10219) );
  NOR2_X1 U11151 ( .A1(n10220), .A2(n10219), .ZN(n10026) );
  AOI22_X1 U11152 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n10310), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n10029), .ZN(n10217) );
  INV_X1 U11153 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10030) );
  AOI22_X1 U11154 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n9516), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n10030), .ZN(n10215) );
  XNOR2_X1 U11155 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10213) );
  INV_X1 U11156 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10035) );
  AOI22_X1 U11157 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n10036), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n10035), .ZN(n10211) );
  NOR2_X1 U11158 ( .A1(n10212), .A2(n10211), .ZN(n10037) );
  AOI22_X1 U11159 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n10040), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n10041), .ZN(n10209) );
  NOR2_X1 U11160 ( .A1(n10210), .A2(n10209), .ZN(n10039) );
  AOI21_X1 U11161 ( .B1(n10041), .B2(n10040), .A(n10039), .ZN(n10208) );
  AOI22_X1 U11162 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n9549), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n10043), .ZN(n10207) );
  NOR2_X1 U11163 ( .A1(n10208), .A2(n10207), .ZN(n10042) );
  NOR2_X1 U11164 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10204), .ZN(n10044) );
  NAND2_X1 U11165 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10204), .ZN(n10203) );
  OAI21_X1 U11166 ( .B1(n10205), .B2(n10044), .A(n10203), .ZN(n10046) );
  XNOR2_X1 U11167 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n10045) );
  XNOR2_X1 U11168 ( .A(n10046), .B(n10045), .ZN(ADD_1068_U4) );
  INV_X1 U11169 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10355) );
  XOR2_X1 U11170 ( .A(n10355), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  XNOR2_X1 U11171 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  NAND3_X1 U11172 ( .A1(n10049), .A2(n10048), .A3(n10047), .ZN(n10050) );
  NAND3_X1 U11173 ( .A1(n10052), .A2(n10051), .A3(n10050), .ZN(n10067) );
  NAND2_X1 U11174 ( .A1(n10054), .A2(n10053), .ZN(n10066) );
  MUX2_X1 U11175 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n7069), .S(n10055), .Z(
        n10056) );
  NAND3_X1 U11176 ( .A1(n10058), .A2(n10057), .A3(n10056), .ZN(n10059) );
  NAND3_X1 U11177 ( .A1(n10061), .A2(n10060), .A3(n10059), .ZN(n10065) );
  AND2_X1 U11178 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10062) );
  AOI21_X1 U11179 ( .B1(n10063), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n10062), .ZN(
        n10064) );
  AND4_X1 U11180 ( .A1(n10067), .A2(n10066), .A3(n10065), .A4(n10064), .ZN(
        n10069) );
  NAND2_X1 U11181 ( .A1(n10069), .A2(n10068), .ZN(P1_U3247) );
  AND2_X1 U11182 ( .A1(n10071), .A2(n10070), .ZN(n10083) );
  INV_X1 U11183 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10073) );
  OAI22_X1 U11184 ( .A1(n10075), .A2(n10074), .B1(n10073), .B2(n10072), .ZN(
        n10076) );
  INV_X1 U11185 ( .A(n10076), .ZN(n10079) );
  NAND2_X1 U11186 ( .A1(n10077), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10078) );
  OAI211_X1 U11187 ( .C1(n10081), .C2(n10080), .A(n10079), .B(n10078), .ZN(
        n10082) );
  NOR2_X1 U11188 ( .A1(n10083), .A2(n10082), .ZN(n10084) );
  OAI21_X1 U11189 ( .B1(n10077), .B2(n10085), .A(n10084), .ZN(P1_U3292) );
  AND2_X1 U11190 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10087), .ZN(P1_U3294) );
  NOR2_X1 U11191 ( .A1(n10086), .A2(n10260), .ZN(P1_U3295) );
  NOR2_X1 U11192 ( .A1(n10086), .A2(n10297), .ZN(P1_U3296) );
  AND2_X1 U11193 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10087), .ZN(P1_U3297) );
  AND2_X1 U11194 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10087), .ZN(P1_U3298) );
  NOR2_X1 U11195 ( .A1(n10086), .A2(n10267), .ZN(P1_U3299) );
  INV_X1 U11196 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10314) );
  NOR2_X1 U11197 ( .A1(n10086), .A2(n10314), .ZN(P1_U3300) );
  AND2_X1 U11198 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10087), .ZN(P1_U3301) );
  NOR2_X1 U11199 ( .A1(n10086), .A2(n10248), .ZN(P1_U3302) );
  AND2_X1 U11200 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10087), .ZN(P1_U3303) );
  AND2_X1 U11201 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10087), .ZN(P1_U3304) );
  AND2_X1 U11202 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10087), .ZN(P1_U3305) );
  AND2_X1 U11203 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10087), .ZN(P1_U3306) );
  AND2_X1 U11204 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10087), .ZN(P1_U3307) );
  AND2_X1 U11205 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10087), .ZN(P1_U3308) );
  AND2_X1 U11206 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10087), .ZN(P1_U3309) );
  AND2_X1 U11207 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10087), .ZN(P1_U3310) );
  AND2_X1 U11208 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10087), .ZN(P1_U3311) );
  AND2_X1 U11209 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10087), .ZN(P1_U3312) );
  AND2_X1 U11210 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10087), .ZN(P1_U3313) );
  AND2_X1 U11211 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10087), .ZN(P1_U3314) );
  AND2_X1 U11212 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10087), .ZN(P1_U3315) );
  AND2_X1 U11213 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10087), .ZN(P1_U3316) );
  AND2_X1 U11214 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10087), .ZN(P1_U3317) );
  AND2_X1 U11215 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10087), .ZN(P1_U3318) );
  AND2_X1 U11216 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10087), .ZN(P1_U3319) );
  AND2_X1 U11217 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10087), .ZN(P1_U3320) );
  INV_X1 U11218 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10346) );
  NOR2_X1 U11219 ( .A1(n10086), .A2(n10346), .ZN(P1_U3321) );
  AND2_X1 U11220 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10087), .ZN(P1_U3322) );
  AND2_X1 U11221 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10087), .ZN(P1_U3323) );
  OAI21_X1 U11222 ( .B1(n10089), .B2(n10107), .A(n10088), .ZN(n10091) );
  AOI211_X1 U11223 ( .C1(n10112), .C2(n10092), .A(n10091), .B(n10090), .ZN(
        n10116) );
  INV_X1 U11224 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10093) );
  AOI22_X1 U11225 ( .A1(n10115), .A2(n10116), .B1(n10093), .B2(n10113), .ZN(
        P1_U3462) );
  OAI21_X1 U11226 ( .B1(n10095), .B2(n10107), .A(n10094), .ZN(n10097) );
  AOI211_X1 U11227 ( .C1(n10112), .C2(n10098), .A(n10097), .B(n10096), .ZN(
        n10117) );
  INV_X1 U11228 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10099) );
  AOI22_X1 U11229 ( .A1(n10115), .A2(n10117), .B1(n10099), .B2(n10113), .ZN(
        P1_U3465) );
  OAI21_X1 U11230 ( .B1(n10101), .B2(n10107), .A(n10100), .ZN(n10103) );
  AOI211_X1 U11231 ( .C1(n10112), .C2(n10104), .A(n10103), .B(n10102), .ZN(
        n10119) );
  INV_X1 U11232 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10105) );
  AOI22_X1 U11233 ( .A1(n10115), .A2(n10119), .B1(n10105), .B2(n10113), .ZN(
        P1_U3468) );
  OAI21_X1 U11234 ( .B1(n10108), .B2(n10107), .A(n10106), .ZN(n10110) );
  AOI211_X1 U11235 ( .C1(n10112), .C2(n10111), .A(n10110), .B(n10109), .ZN(
        n10122) );
  INV_X1 U11236 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10114) );
  AOI22_X1 U11237 ( .A1(n10115), .A2(n10122), .B1(n10114), .B2(n10113), .ZN(
        P1_U3471) );
  AOI22_X1 U11238 ( .A1(n10123), .A2(n10116), .B1(n7068), .B2(n10120), .ZN(
        P1_U3525) );
  AOI22_X1 U11239 ( .A1(n10123), .A2(n10117), .B1(n7069), .B2(n10120), .ZN(
        P1_U3526) );
  AOI22_X1 U11240 ( .A1(n10123), .A2(n10119), .B1(n10118), .B2(n10120), .ZN(
        P1_U3527) );
  AOI22_X1 U11241 ( .A1(n10123), .A2(n10122), .B1(n10121), .B2(n10120), .ZN(
        P1_U3528) );
  INV_X1 U11242 ( .A(n10124), .ZN(n10125) );
  AOI21_X1 U11243 ( .B1(n10127), .B2(n10126), .A(n10125), .ZN(n10142) );
  INV_X1 U11244 ( .A(n10142), .ZN(n10164) );
  OAI22_X1 U11245 ( .A1(n10129), .A2(n10358), .B1(n10161), .B2(n10128), .ZN(
        n10143) );
  AOI22_X1 U11246 ( .A1(n10132), .A2(n6091), .B1(n10131), .B2(n10130), .ZN(
        n10140) );
  INV_X1 U11247 ( .A(n10133), .ZN(n10138) );
  AND3_X1 U11248 ( .A1(n7305), .A2(n10135), .A3(n10134), .ZN(n10137) );
  OAI21_X1 U11249 ( .B1(n10138), .B2(n10137), .A(n10136), .ZN(n10139) );
  OAI211_X1 U11250 ( .C1(n10142), .C2(n10141), .A(n10140), .B(n10139), .ZN(
        n10162) );
  AOI211_X1 U11251 ( .C1(n10144), .C2(n10164), .A(n10143), .B(n10162), .ZN(
        n10146) );
  AOI22_X1 U11252 ( .A1(n10148), .A2(n10147), .B1(n10146), .B2(n10145), .ZN(
        P2_U3231) );
  INV_X1 U11253 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10155) );
  INV_X1 U11254 ( .A(n10149), .ZN(n10153) );
  AOI21_X1 U11255 ( .B1(n10180), .B2(n10151), .A(n10150), .ZN(n10152) );
  AOI211_X1 U11256 ( .C1(n10154), .C2(n10157), .A(n10153), .B(n10152), .ZN(
        n10188) );
  AOI22_X1 U11257 ( .A1(n10186), .A2(n10155), .B1(n10188), .B2(n10184), .ZN(
        P2_U3390) );
  AOI22_X1 U11258 ( .A1(n10158), .A2(n10165), .B1(n10157), .B2(n10156), .ZN(
        n10159) );
  AND2_X1 U11259 ( .A1(n10160), .A2(n10159), .ZN(n10190) );
  AOI22_X1 U11260 ( .A1(n10186), .A2(n5743), .B1(n10190), .B2(n10184), .ZN(
        P2_U3393) );
  NOR2_X1 U11261 ( .A1(n10161), .A2(n10178), .ZN(n10163) );
  AOI211_X1 U11262 ( .C1(n10165), .C2(n10164), .A(n10163), .B(n10162), .ZN(
        n10192) );
  AOI22_X1 U11263 ( .A1(n10186), .A2(n5762), .B1(n10192), .B2(n10184), .ZN(
        P2_U3396) );
  OAI21_X1 U11264 ( .B1(n10167), .B2(n10178), .A(n10166), .ZN(n10168) );
  AOI21_X1 U11265 ( .B1(n10169), .B2(n6186), .A(n10168), .ZN(n10194) );
  AOI22_X1 U11266 ( .A1(n10186), .A2(n5719), .B1(n10194), .B2(n10184), .ZN(
        P2_U3402) );
  INV_X1 U11267 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10176) );
  INV_X1 U11268 ( .A(n10170), .ZN(n10175) );
  OAI22_X1 U11269 ( .A1(n10173), .A2(n10172), .B1(n10171), .B2(n10178), .ZN(
        n10174) );
  NOR2_X1 U11270 ( .A1(n10175), .A2(n10174), .ZN(n10196) );
  AOI22_X1 U11271 ( .A1(n10186), .A2(n10176), .B1(n10196), .B2(n10184), .ZN(
        P2_U3405) );
  INV_X1 U11272 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10185) );
  INV_X1 U11273 ( .A(n10177), .ZN(n10183) );
  OAI22_X1 U11274 ( .A1(n10181), .A2(n10180), .B1(n10179), .B2(n10178), .ZN(
        n10182) );
  NOR2_X1 U11275 ( .A1(n10183), .A2(n10182), .ZN(n10198) );
  AOI22_X1 U11276 ( .A1(n10186), .A2(n10185), .B1(n10198), .B2(n10184), .ZN(
        P2_U3408) );
  AOI22_X1 U11277 ( .A1(n10199), .A2(n10188), .B1(n10187), .B2(n6372), .ZN(
        P2_U3459) );
  AOI22_X1 U11278 ( .A1(n10199), .A2(n10190), .B1(n10189), .B2(n6372), .ZN(
        P2_U3460) );
  AOI22_X1 U11279 ( .A1(n10199), .A2(n10192), .B1(n10191), .B2(n6372), .ZN(
        P2_U3461) );
  INV_X1 U11280 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10193) );
  AOI22_X1 U11281 ( .A1(n10199), .A2(n10194), .B1(n10193), .B2(n6372), .ZN(
        P2_U3463) );
  AOI22_X1 U11282 ( .A1(n10199), .A2(n10196), .B1(n10195), .B2(n6372), .ZN(
        P2_U3464) );
  AOI22_X1 U11283 ( .A1(n10199), .A2(n10198), .B1(n10197), .B2(n6372), .ZN(
        P2_U3465) );
  NOR2_X1 U11284 ( .A1(n10201), .A2(n10200), .ZN(n10202) );
  XOR2_X1 U11285 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10202), .Z(ADD_1068_U5) );
  XOR2_X1 U11286 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI21_X1 U11287 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10204), .A(n10203), 
        .ZN(n10206) );
  XOR2_X1 U11288 ( .A(n10206), .B(n10205), .Z(ADD_1068_U55) );
  XNOR2_X1 U11289 ( .A(n10208), .B(n10207), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11290 ( .A(n10210), .B(n10209), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11291 ( .A(n10212), .B(n10211), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11292 ( .A(n10214), .B(n10213), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11293 ( .A(n10216), .B(n10215), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11294 ( .A(n10218), .B(n10217), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11295 ( .A(n10220), .B(n10219), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11296 ( .A(n10222), .B(n10221), .ZN(ADD_1068_U63) );
  NAND4_X1 U11297 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .A3(n10223), .A4(n10310), .ZN(n10234) );
  NOR4_X1 U11298 ( .A1(SI_18_), .A2(P2_REG1_REG_30__SCAN_IN), .A3(n10293), 
        .A4(n10299), .ZN(n10226) );
  NOR4_X1 U11299 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(P1_DATAO_REG_10__SCAN_IN), .A3(P2_REG0_REG_28__SCAN_IN), .A4(P2_REG2_REG_21__SCAN_IN), .ZN(n10225) );
  NOR3_X1 U11300 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .A3(P2_REG0_REG_7__SCAN_IN), .ZN(n10224) );
  NAND4_X1 U11301 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(n10226), .A3(n10225), 
        .A4(n10224), .ZN(n10233) );
  NAND4_X1 U11302 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(P1_REG2_REG_19__SCAN_IN), 
        .A3(P1_REG0_REG_2__SCAN_IN), .A4(P2_IR_REG_15__SCAN_IN), .ZN(n10232)
         );
  INV_X1 U11303 ( .A(n10227), .ZN(n10230) );
  NOR3_X1 U11304 ( .A1(SI_8_), .A2(P2_REG0_REG_15__SCAN_IN), .A3(n10356), .ZN(
        n10228) );
  NAND4_X1 U11305 ( .A1(n10358), .A2(P2_WR_REG_SCAN_IN), .A3(n10228), .A4(
        P1_ADDR_REG_17__SCAN_IN), .ZN(n10229) );
  OR4_X1 U11306 ( .A1(n10230), .A2(n10339), .A3(n10336), .A4(n10229), .ZN(
        n10231) );
  NOR4_X1 U11307 ( .A1(n10234), .A2(n10233), .A3(n10232), .A4(n10231), .ZN(
        n10373) );
  NAND3_X1 U11308 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        n4771), .ZN(n10245) );
  NOR4_X1 U11309 ( .A1(P2_REG0_REG_4__SCAN_IN), .A2(P2_ADDR_REG_9__SCAN_IN), 
        .A3(P1_ADDR_REG_8__SCAN_IN), .A4(n10296), .ZN(n10235) );
  NAND4_X1 U11310 ( .A1(SI_6_), .A2(n10236), .A3(P2_D_REG_9__SCAN_IN), .A4(
        n10235), .ZN(n10244) );
  NAND4_X1 U11311 ( .A1(n10237), .A2(n10278), .A3(P2_DATAO_REG_7__SCAN_IN), 
        .A4(P1_REG1_REG_2__SCAN_IN), .ZN(n10242) );
  NOR4_X1 U11312 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(P2_REG0_REG_2__SCAN_IN), 
        .A3(n10276), .A4(n10291), .ZN(n10240) );
  NOR4_X1 U11313 ( .A1(SI_17_), .A2(n10261), .A3(n10238), .A4(n10266), .ZN(
        n10239) );
  NAND4_X1 U11314 ( .A1(n10279), .A2(P1_REG0_REG_13__SCAN_IN), .A3(n10240), 
        .A4(n10239), .ZN(n10241) );
  OR4_X1 U11315 ( .A1(n10286), .A2(n10284), .A3(n10242), .A4(n10241), .ZN(
        n10243) );
  NOR4_X1 U11316 ( .A1(SI_12_), .A2(n10245), .A3(n10244), .A4(n10243), .ZN(
        n10372) );
  AOI22_X1 U11317 ( .A1(n10248), .A2(keyinput54), .B1(keyinput62), .B2(n10247), 
        .ZN(n10246) );
  OAI221_X1 U11318 ( .B1(n10248), .B2(keyinput54), .C1(n10247), .C2(keyinput62), .A(n10246), .ZN(n10258) );
  AOI22_X1 U11319 ( .A1(n10251), .A2(keyinput45), .B1(keyinput63), .B2(n10250), 
        .ZN(n10249) );
  OAI221_X1 U11320 ( .B1(n10251), .B2(keyinput45), .C1(n10250), .C2(keyinput63), .A(n10249), .ZN(n10257) );
  AOI22_X1 U11321 ( .A1(n5719), .A2(keyinput51), .B1(n4771), .B2(keyinput46), 
        .ZN(n10252) );
  OAI221_X1 U11322 ( .B1(n5719), .B2(keyinput51), .C1(n4771), .C2(keyinput46), 
        .A(n10252), .ZN(n10256) );
  XNOR2_X1 U11323 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput40), .ZN(n10254) );
  XNOR2_X1 U11324 ( .A(P2_REG3_REG_9__SCAN_IN), .B(keyinput24), .ZN(n10253) );
  NAND2_X1 U11325 ( .A1(n10254), .A2(n10253), .ZN(n10255) );
  NOR4_X1 U11326 ( .A1(n10258), .A2(n10257), .A3(n10256), .A4(n10255), .ZN(
        n10308) );
  AOI22_X1 U11327 ( .A1(n10261), .A2(keyinput11), .B1(n10260), .B2(keyinput23), 
        .ZN(n10259) );
  OAI221_X1 U11328 ( .B1(n10261), .B2(keyinput11), .C1(n10260), .C2(keyinput23), .A(n10259), .ZN(n10273) );
  AOI22_X1 U11329 ( .A1(n10264), .A2(keyinput44), .B1(keyinput49), .B2(n10263), 
        .ZN(n10262) );
  OAI221_X1 U11330 ( .B1(n10264), .B2(keyinput44), .C1(n10263), .C2(keyinput49), .A(n10262), .ZN(n10272) );
  AOI22_X1 U11331 ( .A1(n10267), .A2(keyinput8), .B1(keyinput56), .B2(n10266), 
        .ZN(n10265) );
  OAI221_X1 U11332 ( .B1(n10267), .B2(keyinput8), .C1(n10266), .C2(keyinput56), 
        .A(n10265), .ZN(n10271) );
  XNOR2_X1 U11333 ( .A(P2_D_REG_1__SCAN_IN), .B(keyinput43), .ZN(n10269) );
  XNOR2_X1 U11334 ( .A(P1_REG1_REG_2__SCAN_IN), .B(keyinput37), .ZN(n10268) );
  NAND2_X1 U11335 ( .A1(n10269), .A2(n10268), .ZN(n10270) );
  NOR4_X1 U11336 ( .A1(n10273), .A2(n10272), .A3(n10271), .A4(n10270), .ZN(
        n10307) );
  AOI22_X1 U11337 ( .A1(n10276), .A2(keyinput38), .B1(keyinput42), .B2(n10275), 
        .ZN(n10274) );
  OAI221_X1 U11338 ( .B1(n10276), .B2(keyinput38), .C1(n10275), .C2(keyinput42), .A(n10274), .ZN(n10282) );
  AOI22_X1 U11339 ( .A1(n10279), .A2(keyinput29), .B1(n10278), .B2(keyinput13), 
        .ZN(n10277) );
  OAI221_X1 U11340 ( .B1(n10279), .B2(keyinput29), .C1(n10278), .C2(keyinput13), .A(n10277), .ZN(n10281) );
  XOR2_X1 U11341 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput31), .Z(n10280) );
  OR3_X1 U11342 ( .A1(n10282), .A2(n10281), .A3(n10280), .ZN(n10289) );
  INV_X1 U11343 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10285) );
  AOI22_X1 U11344 ( .A1(n10285), .A2(keyinput55), .B1(keyinput57), .B2(n10284), 
        .ZN(n10283) );
  OAI221_X1 U11345 ( .B1(n10285), .B2(keyinput55), .C1(n10284), .C2(keyinput57), .A(n10283), .ZN(n10288) );
  XNOR2_X1 U11346 ( .A(n10286), .B(keyinput33), .ZN(n10287) );
  NOR3_X1 U11347 ( .A1(n10289), .A2(n10288), .A3(n10287), .ZN(n10306) );
  AOI22_X1 U11348 ( .A1(n10291), .A2(keyinput3), .B1(keyinput15), .B2(n5762), 
        .ZN(n10290) );
  OAI221_X1 U11349 ( .B1(n10291), .B2(keyinput3), .C1(n5762), .C2(keyinput15), 
        .A(n10290), .ZN(n10304) );
  AOI22_X1 U11350 ( .A1(n10294), .A2(keyinput21), .B1(n10293), .B2(keyinput9), 
        .ZN(n10292) );
  OAI221_X1 U11351 ( .B1(n10294), .B2(keyinput21), .C1(n10293), .C2(keyinput9), 
        .A(n10292), .ZN(n10303) );
  AOI22_X1 U11352 ( .A1(n10297), .A2(keyinput1), .B1(keyinput17), .B2(n10296), 
        .ZN(n10295) );
  OAI221_X1 U11353 ( .B1(n10297), .B2(keyinput1), .C1(n10296), .C2(keyinput17), 
        .A(n10295), .ZN(n10302) );
  AOI22_X1 U11354 ( .A1(n10300), .A2(keyinput10), .B1(keyinput32), .B2(n10299), 
        .ZN(n10298) );
  OAI221_X1 U11355 ( .B1(n10300), .B2(keyinput10), .C1(n10299), .C2(keyinput32), .A(n10298), .ZN(n10301) );
  NOR4_X1 U11356 ( .A1(n10304), .A2(n10303), .A3(n10302), .A4(n10301), .ZN(
        n10305) );
  NAND4_X1 U11357 ( .A1(n10308), .A2(n10307), .A3(n10306), .A4(n10305), .ZN(
        n10371) );
  AOI22_X1 U11358 ( .A1(n10311), .A2(keyinput20), .B1(keyinput52), .B2(n10310), 
        .ZN(n10309) );
  OAI221_X1 U11359 ( .B1(n10311), .B2(keyinput20), .C1(n10310), .C2(keyinput52), .A(n10309), .ZN(n10321) );
  AOI22_X1 U11360 ( .A1(n10314), .A2(keyinput2), .B1(keyinput22), .B2(n10313), 
        .ZN(n10312) );
  OAI221_X1 U11361 ( .B1(n10314), .B2(keyinput2), .C1(n10313), .C2(keyinput22), 
        .A(n10312), .ZN(n10320) );
  XNOR2_X1 U11362 ( .A(SI_8_), .B(keyinput5), .ZN(n10318) );
  XNOR2_X1 U11363 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput18), .ZN(n10317) );
  XNOR2_X1 U11364 ( .A(P2_REG2_REG_12__SCAN_IN), .B(keyinput28), .ZN(n10316)
         );
  XNOR2_X1 U11365 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput14), .ZN(n10315) );
  NAND4_X1 U11366 ( .A1(n10318), .A2(n10317), .A3(n10316), .A4(n10315), .ZN(
        n10319) );
  NOR3_X1 U11367 ( .A1(n10321), .A2(n10320), .A3(n10319), .ZN(n10369) );
  AOI22_X1 U11368 ( .A1(n10323), .A2(keyinput59), .B1(keyinput19), .B2(n8240), 
        .ZN(n10322) );
  OAI221_X1 U11369 ( .B1(n10323), .B2(keyinput59), .C1(n8240), .C2(keyinput19), 
        .A(n10322), .ZN(n10334) );
  AOI22_X1 U11370 ( .A1(n10326), .A2(keyinput4), .B1(keyinput53), .B2(n10325), 
        .ZN(n10324) );
  OAI221_X1 U11371 ( .B1(n10326), .B2(keyinput4), .C1(n10325), .C2(keyinput53), 
        .A(n10324), .ZN(n10333) );
  XNOR2_X1 U11372 ( .A(n10327), .B(keyinput26), .ZN(n10332) );
  XOR2_X1 U11373 ( .A(n6546), .B(keyinput16), .Z(n10330) );
  XNOR2_X1 U11374 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(keyinput48), .ZN(n10329)
         );
  XNOR2_X1 U11375 ( .A(P1_REG3_REG_8__SCAN_IN), .B(keyinput58), .ZN(n10328) );
  NAND3_X1 U11376 ( .A1(n10330), .A2(n10329), .A3(n10328), .ZN(n10331) );
  NOR4_X1 U11377 ( .A1(n10334), .A2(n10333), .A3(n10332), .A4(n10331), .ZN(
        n10368) );
  AOI22_X1 U11378 ( .A1(n10337), .A2(keyinput12), .B1(n10336), .B2(keyinput47), 
        .ZN(n10335) );
  OAI221_X1 U11379 ( .B1(n10337), .B2(keyinput12), .C1(n10336), .C2(keyinput47), .A(n10335), .ZN(n10344) );
  XNOR2_X1 U11380 ( .A(n10338), .B(keyinput36), .ZN(n10343) );
  XNOR2_X1 U11381 ( .A(n10339), .B(keyinput30), .ZN(n10342) );
  XNOR2_X1 U11382 ( .A(n10340), .B(keyinput7), .ZN(n10341) );
  OR4_X1 U11383 ( .A1(n10344), .A2(n10343), .A3(n10342), .A4(n10341), .ZN(
        n10350) );
  AOI22_X1 U11384 ( .A1(n9549), .A2(keyinput39), .B1(n10346), .B2(keyinput0), 
        .ZN(n10345) );
  OAI221_X1 U11385 ( .B1(n9549), .B2(keyinput39), .C1(n10346), .C2(keyinput0), 
        .A(n10345), .ZN(n10349) );
  XNOR2_X1 U11386 ( .A(n10347), .B(keyinput27), .ZN(n10348) );
  NOR3_X1 U11387 ( .A1(n10350), .A2(n10349), .A3(n10348), .ZN(n10367) );
  INV_X1 U11388 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10352) );
  AOI22_X1 U11389 ( .A1(n10353), .A2(keyinput35), .B1(n10352), .B2(keyinput6), 
        .ZN(n10351) );
  OAI221_X1 U11390 ( .B1(n10353), .B2(keyinput35), .C1(n10352), .C2(keyinput6), 
        .A(n10351), .ZN(n10365) );
  AOI22_X1 U11391 ( .A1(n10356), .A2(keyinput50), .B1(keyinput60), .B2(n10355), 
        .ZN(n10354) );
  OAI221_X1 U11392 ( .B1(n10356), .B2(keyinput50), .C1(n10355), .C2(keyinput60), .A(n10354), .ZN(n10364) );
  AOI22_X1 U11393 ( .A1(n10359), .A2(keyinput41), .B1(keyinput34), .B2(n10358), 
        .ZN(n10357) );
  OAI221_X1 U11394 ( .B1(n10359), .B2(keyinput41), .C1(n10358), .C2(keyinput34), .A(n10357), .ZN(n10363) );
  AOI22_X1 U11395 ( .A1(n10361), .A2(keyinput61), .B1(n6530), .B2(keyinput25), 
        .ZN(n10360) );
  OAI221_X1 U11396 ( .B1(n10361), .B2(keyinput61), .C1(n6530), .C2(keyinput25), 
        .A(n10360), .ZN(n10362) );
  NOR4_X1 U11397 ( .A1(n10365), .A2(n10364), .A3(n10363), .A4(n10362), .ZN(
        n10366) );
  NAND4_X1 U11398 ( .A1(n10369), .A2(n10368), .A3(n10367), .A4(n10366), .ZN(
        n10370) );
  AOI211_X1 U11399 ( .C1(n10373), .C2(n10372), .A(n10371), .B(n10370), .ZN(
        n10377) );
  MUX2_X1 U11400 ( .A(n10375), .B(n10374), .S(P1_U3973), .Z(n10376) );
  XNOR2_X1 U11401 ( .A(n10377), .B(n10376), .ZN(P1_U3581) );
  XNOR2_X1 U11402 ( .A(n10379), .B(n10378), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11403 ( .A(n10381), .B(n10380), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11404 ( .A(n10383), .B(n10382), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11405 ( .A(n10385), .B(n10384), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11406 ( .A(n10387), .B(n10386), .ZN(ADD_1068_U48) );
  XOR2_X1 U11407 ( .A(n10389), .B(n10388), .Z(ADD_1068_U54) );
  XOR2_X1 U11408 ( .A(n10391), .B(n10390), .Z(ADD_1068_U53) );
  XNOR2_X1 U11409 ( .A(n10393), .B(n10392), .ZN(ADD_1068_U52) );
  INV_X1 U4787 ( .A(n6918), .ZN(n8543) );
  CLKBUF_X1 U4800 ( .A(n5761), .Z(n4695) );
  CLKBUF_X1 U5753 ( .A(n5851), .Z(n6143) );
  INV_X2 U7377 ( .A(n5757), .ZN(n8309) );
endmodule

