

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347;

  CLKBUF_X2 U2527 ( .A(n3107), .Z(n3794) );
  OAI21_X1 U2528 ( .B1(n3107), .B2(n2574), .A(n2573), .ZN(n3116) );
  NAND2_X1 U2529 ( .A1(n2823), .A2(IR_REG_31__SCAN_IN), .ZN(n2824) );
  NOR2_X4 U2530 ( .A1(n2768), .A2(n2634), .ZN(n2765) );
  AND2_X4 U2531 ( .A1(n3000), .A2(n2958), .ZN(n4050) );
  XNOR2_X2 U2532 ( .A(n2824), .B(n4800), .ZN(n2908) );
  NAND2_X1 U2533 ( .A1(n4072), .A2(n4071), .ZN(n4200) );
  AND2_X1 U2534 ( .A1(n2568), .A2(n2535), .ZN(n5281) );
  OR2_X1 U2535 ( .A1(n3765), .A2(n2715), .ZN(n2570) );
  NAND2_X2 U2536 ( .A1(n3856), .A2(n3859), .ZN(n3080) );
  INV_X4 U2537 ( .A(n3024), .ZN(n3490) );
  INV_X8 U2538 ( .A(n4112), .ZN(n3492) );
  CLKBUF_X3 U2539 ( .A(n3240), .Z(n2494) );
  AND2_X1 U2540 ( .A1(n5066), .A2(n2924), .ZN(n3240) );
  NOR2_X1 U2542 ( .A1(n4089), .A2(n4099), .ZN(n4179) );
  OAI21_X1 U2543 ( .B1(n4108), .B2(n4107), .A(n4106), .ZN(n4213) );
  NAND2_X1 U2544 ( .A1(n4898), .A2(n2513), .ZN(n4880) );
  AND2_X1 U2545 ( .A1(n4484), .A2(n4467), .ZN(n4465) );
  NAND2_X1 U2546 ( .A1(n4921), .A2(n2585), .ZN(n4890) );
  OR2_X1 U2547 ( .A1(n4987), .A2(n4956), .ZN(n4963) );
  NAND2_X1 U2548 ( .A1(n3523), .A2(n3522), .ZN(n3620) );
  AND2_X1 U2549 ( .A1(n3320), .A2(n3319), .ZN(n3343) );
  OAI22_X1 U2550 ( .A1(n3257), .A2(n3256), .B1(n3334), .B2(n4232), .ZN(n3260)
         );
  OAI21_X1 U2551 ( .B1(n3157), .B2(n3156), .A(n3870), .ZN(n3223) );
  CLKBUF_X1 U2552 ( .A(n4219), .Z(n5276) );
  NOR2_X1 U2553 ( .A1(n3054), .A2(n5068), .ZN(n4219) );
  NOR2_X1 U2554 ( .A1(n3230), .A2(n3334), .ZN(n3251) );
  AND2_X1 U2555 ( .A1(n3860), .A2(n3863), .ZN(n3837) );
  NAND2_X4 U2556 ( .A1(n4999), .A2(n3000), .ZN(n3024) );
  NAND4_X1 U2557 ( .A1(n2994), .A2(n2993), .A3(n2992), .A4(n2991), .ZN(n4234)
         );
  NAND4_X1 U2558 ( .A1(n2955), .A2(n2954), .A3(n2953), .A4(n2952), .ZN(n4236)
         );
  NAND4_X1 U2559 ( .A1(n3061), .A2(n3060), .A3(n3059), .A4(n3058), .ZN(n3108)
         );
  NAND2_X1 U2560 ( .A1(n2999), .A2(n2998), .ZN(n4999) );
  OAI21_X1 U2561 ( .B1(n3107), .B2(n2572), .A(n2571), .ZN(n3079) );
  INV_X1 U2562 ( .A(n3099), .ZN(n3000) );
  INV_X1 U2563 ( .A(n3208), .ZN(n3215) );
  AND2_X2 U2564 ( .A1(n2925), .A2(n2924), .ZN(n3057) );
  AND2_X2 U2565 ( .A1(n5067), .A2(n5066), .ZN(n3109) );
  AND2_X1 U2566 ( .A1(n2997), .A2(n3858), .ZN(n3099) );
  AND2_X2 U2567 ( .A1(n5067), .A2(n2925), .ZN(n3056) );
  INV_X1 U2568 ( .A(n2924), .ZN(n5067) );
  XNOR2_X1 U2569 ( .A(n2956), .B(n4789), .ZN(n2961) );
  OR3_X1 U2570 ( .A1(n2956), .A2(n2957), .A3(n5064), .ZN(n2640) );
  XNOR2_X1 U2571 ( .A(n2827), .B(n4801), .ZN(n3043) );
  XNOR2_X1 U2572 ( .A(n2922), .B(IR_REG_30__SCAN_IN), .ZN(n5066) );
  OAI211_X1 U2573 ( .C1(IR_REG_29__SCAN_IN), .C2(IR_REG_31__SCAN_IN), .A(n2920), .B(n2921), .ZN(n2924) );
  NAND2_X1 U2574 ( .A1(n2836), .A2(IR_REG_31__SCAN_IN), .ZN(n2837) );
  NAND2_X1 U2575 ( .A1(n2813), .A2(IR_REG_31__SCAN_IN), .ZN(n2956) );
  NAND2_X1 U2576 ( .A1(n2915), .A2(n2741), .ZN(n2920) );
  OAI21_X1 U2577 ( .B1(n2566), .B2(n2565), .A(IR_REG_31__SCAN_IN), .ZN(n2841)
         );
  AND2_X1 U2578 ( .A1(n2821), .A2(n2666), .ZN(n2812) );
  NOR2_X1 U2579 ( .A1(n2566), .A2(IR_REG_22__SCAN_IN), .ZN(n2825) );
  AND2_X1 U2580 ( .A1(n2498), .A2(n2511), .ZN(n2666) );
  INV_X1 U2581 ( .A(n2913), .ZN(n2565) );
  AND2_X1 U2582 ( .A1(n2913), .A2(n2840), .ZN(n2918) );
  AND2_X1 U2583 ( .A1(n2504), .A2(n4776), .ZN(n2497) );
  AND2_X1 U2584 ( .A1(n2839), .A2(n2838), .ZN(n2913) );
  AND2_X1 U2585 ( .A1(n2829), .A2(n2828), .ZN(n2839) );
  AND2_X1 U2586 ( .A1(n4806), .A2(n4613), .ZN(n2838) );
  AND2_X1 U2587 ( .A1(n2747), .A2(n4766), .ZN(n2632) );
  NOR2_X1 U2588 ( .A1(IR_REG_25__SCAN_IN), .A2(IR_REG_22__SCAN_IN), .ZN(n2829)
         );
  NOR2_X1 U2589 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2828)
         );
  INV_X1 U2590 ( .A(IR_REG_4__SCAN_IN), .ZN(n2747) );
  NOR2_X2 U2591 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2783)
         );
  INV_X1 U2592 ( .A(IR_REG_3__SCAN_IN), .ZN(n4571) );
  INV_X1 U2593 ( .A(IR_REG_2__SCAN_IN), .ZN(n4766) );
  INV_X1 U2594 ( .A(IR_REG_12__SCAN_IN), .ZN(n4587) );
  INV_X1 U2595 ( .A(IR_REG_11__SCAN_IN), .ZN(n4781) );
  INV_X1 U2596 ( .A(IR_REG_10__SCAN_IN), .ZN(n4775) );
  NOR2_X1 U2597 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2633)
         );
  BUF_X1 U2598 ( .A(n5013), .Z(n2492) );
  INV_X1 U2599 ( .A(n2961), .ZN(n5130) );
  AND2_X1 U2600 ( .A1(n2925), .A2(n2924), .ZN(n2493) );
  NAND2_X2 U2601 ( .A1(n3099), .A2(n2958), .ZN(n4112) );
  OR2_X2 U2602 ( .A1(n4449), .A2(n4431), .ZN(n4432) );
  NOR2_X4 U2603 ( .A1(n4432), .A2(n4386), .ZN(n5330) );
  AND2_X4 U2604 ( .A1(n4050), .A2(n3188), .ZN(n3026) );
  XNOR2_X2 U2605 ( .A(n2837), .B(n4613), .ZN(n2846) );
  NOR2_X1 U2606 ( .A1(n4443), .A2(n2550), .ZN(n2549) );
  INV_X1 U2607 ( .A(n4406), .ZN(n2550) );
  AOI21_X1 U2608 ( .B1(n3930), .B2(n2618), .A(n2617), .ZN(n2616) );
  INV_X1 U2609 ( .A(n3965), .ZN(n2617) );
  INV_X1 U2610 ( .A(n3930), .ZN(n2619) );
  NOR2_X1 U2611 ( .A1(REG2_REG_16__SCAN_IN), .A2(n4335), .ZN(n4334) );
  NAND2_X1 U2612 ( .A1(n4456), .A2(n4378), .ZN(n4440) );
  AND2_X1 U2613 ( .A1(n4425), .A2(n2691), .ZN(n2690) );
  NAND2_X1 U2614 ( .A1(n4379), .A2(n4382), .ZN(n2691) );
  AND2_X1 U2615 ( .A1(n3965), .A2(n3927), .ZN(n3930) );
  AND2_X1 U2616 ( .A1(n4096), .A2(n4097), .ZN(n2631) );
  INV_X1 U2617 ( .A(n5270), .ZN(n3991) );
  OR2_X1 U2618 ( .A1(n3731), .A2(n3730), .ZN(n3733) );
  AND2_X1 U2619 ( .A1(n3928), .A2(n3640), .ZN(n3644) );
  NAND2_X1 U2620 ( .A1(n3691), .A2(REG3_REG_26__SCAN_IN), .ZN(n3779) );
  NAND2_X1 U2621 ( .A1(n2945), .A2(n2944), .ZN(n2943) );
  NOR2_X1 U2622 ( .A1(n4263), .A2(n5187), .ZN(n4262) );
  XNOR2_X1 U2623 ( .A(n2795), .B(n2794), .ZN(n4273) );
  INV_X1 U2624 ( .A(n5074), .ZN(n2794) );
  NAND2_X1 U2625 ( .A1(n4273), .A2(REG2_REG_8__SCAN_IN), .ZN(n4272) );
  XNOR2_X1 U2626 ( .A(n3463), .B(n2872), .ZN(n4304) );
  NAND2_X1 U2627 ( .A1(n3943), .A2(n3942), .ZN(n3941) );
  OAI21_X1 U2628 ( .B1(n2606), .B2(n4334), .A(n2537), .ZN(n4356) );
  NAND2_X1 U2629 ( .A1(n2610), .A2(n2607), .ZN(n2606) );
  INV_X1 U2630 ( .A(n4358), .ZN(n2607) );
  NAND2_X1 U2631 ( .A1(n2688), .A2(n2686), .ZN(n2685) );
  OR2_X1 U2632 ( .A1(n2690), .A2(n2693), .ZN(n2686) );
  NAND2_X1 U2633 ( .A1(n2554), .A2(n4406), .ZN(n4444) );
  INV_X1 U2634 ( .A(n2553), .ZN(n4442) );
  NAND2_X1 U2635 ( .A1(n2676), .A2(n2674), .ZN(n4456) );
  AOI21_X1 U2636 ( .B1(n2677), .B2(n2679), .A(n2675), .ZN(n2674) );
  AOI21_X1 U2637 ( .B1(n2697), .B2(n3817), .A(n4374), .ZN(n2695) );
  OR2_X1 U2638 ( .A1(n4935), .A2(n2696), .ZN(n2694) );
  INV_X1 U2639 ( .A(n2697), .ZN(n2696) );
  OR2_X1 U2640 ( .A1(n3751), .A2(n4195), .ZN(n3745) );
  AOI21_X1 U2641 ( .B1(n2712), .B2(n2709), .A(n2519), .ZN(n2708) );
  NOR2_X1 U2642 ( .A1(n2713), .A2(n3655), .ZN(n2709) );
  NAND2_X1 U2643 ( .A1(n2712), .A2(n2711), .ZN(n2710) );
  INV_X1 U2644 ( .A(n3655), .ZN(n2711) );
  INV_X1 U2645 ( .A(n2714), .ZN(n2713) );
  OAI21_X1 U2646 ( .B1(n2496), .B2(n3541), .A(n2715), .ZN(n2714) );
  NAND2_X1 U2647 ( .A1(n3581), .A2(n3626), .ZN(n3538) );
  AND2_X1 U2648 ( .A1(n4236), .A2(n3079), .ZN(n3081) );
  INV_X1 U2649 ( .A(IR_REG_19__SCAN_IN), .ZN(n4789) );
  NAND2_X1 U2650 ( .A1(n4093), .A2(n4098), .ZN(n2630) );
  AND2_X1 U2651 ( .A1(n4458), .A2(n4485), .ZN(n3809) );
  INV_X1 U2652 ( .A(n3080), .ZN(n3839) );
  OAI21_X1 U2653 ( .B1(n3500), .B2(n3501), .A(n3505), .ZN(n2645) );
  AND2_X1 U2654 ( .A1(n3415), .A2(n3413), .ZN(n3500) );
  INV_X1 U2655 ( .A(n3823), .ZN(n3858) );
  AND2_X1 U2656 ( .A1(n3355), .A2(REG1_REG_9__SCAN_IN), .ZN(n2867) );
  OAI21_X1 U2657 ( .B1(n4313), .B2(n2725), .A(n2724), .ZN(n2882) );
  NAND2_X1 U2658 ( .A1(n4320), .A2(n2726), .ZN(n2724) );
  INV_X1 U2659 ( .A(n4341), .ZN(n2611) );
  AND2_X1 U2660 ( .A1(n2553), .A2(n2552), .ZN(n4426) );
  NAND2_X1 U2661 ( .A1(n2554), .A2(n2549), .ZN(n2553) );
  OR2_X1 U2662 ( .A1(n4222), .A2(n4944), .ZN(n4902) );
  NOR2_X1 U2663 ( .A1(n5281), .A2(n5290), .ZN(n4395) );
  NOR2_X1 U2664 ( .A1(n2672), .A2(n2669), .ZN(n2668) );
  NOR2_X1 U2665 ( .A1(n3657), .A2(n2705), .ZN(n2704) );
  INV_X1 U2666 ( .A(n2708), .ZN(n2705) );
  NAND2_X1 U2667 ( .A1(n3515), .A2(n2581), .ZN(n2580) );
  INV_X1 U2668 ( .A(n3353), .ZN(n2699) );
  OAI21_X1 U2669 ( .B1(n3840), .B2(n2560), .A(n3816), .ZN(n2559) );
  INV_X1 U2670 ( .A(n3874), .ZN(n2560) );
  AND2_X1 U2671 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n3110) );
  NOR2_X1 U2672 ( .A1(n3586), .A2(n3634), .ZN(n3585) );
  INV_X1 U2673 ( .A(IR_REG_28__SCAN_IN), .ZN(n2840) );
  AND3_X1 U2674 ( .A1(n4587), .A2(n4775), .A3(n4781), .ZN(n2748) );
  INV_X1 U2675 ( .A(IR_REG_9__SCAN_IN), .ZN(n4776) );
  NOR2_X1 U2676 ( .A1(n2768), .A2(IR_REG_3__SCAN_IN), .ZN(n2776) );
  NAND2_X1 U2677 ( .A1(n2650), .A2(n2503), .ZN(n2649) );
  AND2_X1 U2678 ( .A1(n2503), .A2(n3330), .ZN(n2651) );
  INV_X1 U2679 ( .A(n4154), .ZN(n4080) );
  NAND2_X1 U2680 ( .A1(n4007), .A2(n2657), .ZN(n2656) );
  INV_X1 U2681 ( .A(n2628), .ZN(n2626) );
  NAND2_X1 U2682 ( .A1(n3619), .A2(n3618), .ZN(n2664) );
  NAND2_X1 U2683 ( .A1(n3620), .A2(n2665), .ZN(n2663) );
  OR2_X1 U2684 ( .A1(n3619), .A2(n3618), .ZN(n2665) );
  INV_X1 U2685 ( .A(n3659), .ZN(n3658) );
  INV_X1 U2686 ( .A(n4104), .ZN(n4105) );
  NAND2_X1 U2687 ( .A1(n3970), .A2(n2514), .ZN(n3985) );
  NOR2_X1 U2688 ( .A1(n3542), .A2(n4726), .ZN(n3560) );
  NAND2_X1 U2689 ( .A1(n2739), .A2(REG1_REG_3__SCAN_IN), .ZN(n2737) );
  OR2_X1 U2690 ( .A1(n2853), .A2(n4248), .ZN(n2739) );
  AND2_X1 U2691 ( .A1(n2853), .A2(n4248), .ZN(n2854) );
  NAND2_X1 U2692 ( .A1(n4254), .A2(n2788), .ZN(n2789) );
  NAND2_X1 U2693 ( .A1(n4259), .A2(n2793), .ZN(n2945) );
  OAI21_X1 U2694 ( .B1(n4262), .B2(n2734), .A(n2733), .ZN(n2863) );
  NAND2_X1 U2695 ( .A1(n2941), .A2(n2735), .ZN(n2733) );
  OR2_X1 U2696 ( .A1(n2860), .A2(n2862), .ZN(n2734) );
  NOR2_X1 U2697 ( .A1(n4282), .A2(n4281), .ZN(n4280) );
  INV_X1 U2698 ( .A(n2602), .ZN(n2596) );
  NOR2_X1 U2699 ( .A1(n3373), .A2(n2603), .ZN(n2602) );
  NAND2_X1 U2700 ( .A1(n2601), .A2(n2600), .ZN(n2599) );
  NAND2_X1 U2701 ( .A1(n2604), .A2(n2603), .ZN(n2598) );
  INV_X1 U2702 ( .A(n2743), .ZN(n2600) );
  NAND2_X1 U2703 ( .A1(n2800), .A2(n3481), .ZN(n2801) );
  NAND2_X1 U2704 ( .A1(n2871), .A2(n2870), .ZN(n2872) );
  NOR2_X1 U2705 ( .A1(n5236), .A2(n4304), .ZN(n4303) );
  NAND2_X1 U2706 ( .A1(n3941), .A2(n2803), .ZN(n2804) );
  XNOR2_X1 U2707 ( .A(n2807), .B(n3654), .ZN(n4335) );
  XNOR2_X1 U2708 ( .A(n2882), .B(n3654), .ZN(n4332) );
  AND2_X1 U2709 ( .A1(n2690), .A2(n2693), .ZN(n2683) );
  AOI21_X1 U2710 ( .B1(n2690), .B2(n2692), .A(n2525), .ZN(n2688) );
  INV_X1 U2711 ( .A(n4382), .ZN(n2692) );
  NOR2_X1 U2712 ( .A1(n4424), .A2(n2551), .ZN(n4427) );
  NAND2_X1 U2713 ( .A1(n2546), .A2(n2544), .ZN(n2551) );
  NAND2_X1 U2714 ( .A1(n2548), .A2(n2545), .ZN(n2544) );
  OR2_X1 U2715 ( .A1(n4460), .A2(n2547), .ZN(n2546) );
  NOR2_X2 U2716 ( .A1(n4890), .A2(n4485), .ZN(n4484) );
  AOI21_X1 U2717 ( .B1(n2680), .B2(n2678), .A(n2520), .ZN(n2677) );
  INV_X1 U2718 ( .A(n4376), .ZN(n2678) );
  INV_X1 U2719 ( .A(n2680), .ZN(n2679) );
  AND2_X1 U2720 ( .A1(n2506), .A2(n4477), .ZN(n2680) );
  NAND2_X1 U2721 ( .A1(n2694), .A2(n2516), .ZN(n4898) );
  NAND2_X1 U2722 ( .A1(n3690), .A2(n3689), .ZN(n3731) );
  AND2_X1 U2723 ( .A1(n2500), .A2(n4919), .ZN(n2697) );
  NAND2_X1 U2724 ( .A1(n3666), .A2(n3667), .ZN(n3949) );
  OR2_X1 U2725 ( .A1(n3672), .A2(n3894), .ZN(n5290) );
  INV_X1 U2726 ( .A(n3966), .ZN(n3974) );
  AOI21_X1 U2727 ( .B1(n2713), .B2(n2496), .A(n2524), .ZN(n2712) );
  INV_X1 U2728 ( .A(n3634), .ZN(n3649) );
  NAND2_X1 U2729 ( .A1(n2577), .A2(n3626), .ZN(n3586) );
  NAND2_X1 U2730 ( .A1(n3424), .A2(n3532), .ZN(n3471) );
  NOR2_X1 U2731 ( .A1(n3820), .A2(n3468), .ZN(n3469) );
  AND2_X1 U2732 ( .A1(n3880), .A2(n3876), .ZN(n3838) );
  AND2_X1 U2733 ( .A1(n3077), .A2(n3076), .ZN(n5288) );
  NAND2_X1 U2734 ( .A1(n3223), .A2(n3841), .ZN(n3158) );
  NOR2_X1 U2735 ( .A1(n5296), .A2(n5130), .ZN(n2962) );
  NAND2_X1 U2736 ( .A1(n2575), .A2(n3349), .ZN(n3230) );
  OR2_X1 U2737 ( .A1(n3099), .A2(n4997), .ZN(n2999) );
  AOI21_X1 U2738 ( .B1(n2997), .B2(n3082), .A(n5130), .ZN(n2998) );
  INV_X1 U2739 ( .A(n2850), .ZN(n2574) );
  INV_X1 U2740 ( .A(n5288), .ZN(n5124) );
  INV_X1 U2741 ( .A(IR_REG_29__SCAN_IN), .ZN(n4811) );
  AND2_X1 U2742 ( .A1(n2957), .A2(n4789), .ZN(n2639) );
  OAI21_X1 U2743 ( .B1(n2957), .B2(n4789), .A(IR_REG_31__SCAN_IN), .ZN(n2637)
         );
  INV_X1 U2744 ( .A(IR_REG_8__SCAN_IN), .ZN(n2635) );
  NAND2_X1 U2745 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2721)
         );
  NOR2_X1 U2746 ( .A1(n2626), .A2(n4093), .ZN(n2625) );
  NAND2_X1 U2747 ( .A1(n2631), .A2(n5271), .ZN(n2628) );
  INV_X1 U2748 ( .A(n2631), .ZN(n2622) );
  NAND2_X1 U2749 ( .A1(n3107), .A2(DATAI_0_), .ZN(n2571) );
  NAND2_X1 U2750 ( .A1(n3787), .A2(n3786), .ZN(n4464) );
  OR2_X1 U2751 ( .A1(n4468), .A2(n3790), .ZN(n3698) );
  NAND2_X1 U2752 ( .A1(n3716), .A2(n3715), .ZN(n4909) );
  NAND4_X1 U2753 ( .A1(n3300), .A2(n3299), .A3(n3298), .A4(n3297), .ZN(n4229)
         );
  XNOR2_X1 U2754 ( .A(n2850), .B(n2849), .ZN(n4239) );
  NAND2_X1 U2755 ( .A1(n2796), .A2(n4272), .ZN(n4286) );
  XNOR2_X1 U2756 ( .A(n2719), .B(n2541), .ZN(n2718) );
  NAND2_X1 U2757 ( .A1(n4361), .A2(n2886), .ZN(n2719) );
  NOR2_X1 U2758 ( .A1(n4356), .A2(n2540), .ZN(n2816) );
  OAI21_X1 U2759 ( .B1(n3080), .B2(n3081), .A(n3118), .ZN(n5140) );
  NAND2_X1 U2760 ( .A1(n2933), .A2(n2791), .ZN(n2792) );
  NAND2_X1 U2761 ( .A1(n2717), .A2(n2857), .ZN(n2858) );
  NAND2_X1 U2762 ( .A1(n2876), .A2(n2875), .ZN(n2877) );
  NAND2_X1 U2763 ( .A1(n4322), .A2(n2539), .ZN(n2807) );
  NAND2_X1 U2764 ( .A1(n5072), .A2(REG2_REG_17__SCAN_IN), .ZN(n2612) );
  NAND2_X1 U2765 ( .A1(n2548), .A2(n2675), .ZN(n2547) );
  AND2_X1 U2766 ( .A1(n4425), .A2(n2552), .ZN(n2548) );
  INV_X1 U2767 ( .A(n2549), .ZN(n2545) );
  NAND2_X1 U2768 ( .A1(n3210), .A2(n3266), .ZN(n3866) );
  NAND2_X1 U2769 ( .A1(n3281), .A2(n3108), .ZN(n3870) );
  NAND2_X1 U2770 ( .A1(n3866), .A2(n3870), .ZN(n3134) );
  NAND2_X1 U2771 ( .A1(n3839), .A2(n2567), .ZN(n3104) );
  INV_X1 U2772 ( .A(IR_REG_18__SCAN_IN), .ZN(n2811) );
  INV_X1 U2773 ( .A(IR_REG_15__SCAN_IN), .ZN(n4597) );
  INV_X1 U2774 ( .A(IR_REG_14__SCAN_IN), .ZN(n2749) );
  NAND3_X1 U2775 ( .A1(n2644), .A2(n2642), .A3(n2641), .ZN(n2647) );
  NAND2_X1 U2776 ( .A1(n2643), .A2(n3506), .ZN(n2642) );
  INV_X1 U2777 ( .A(n2645), .ZN(n2644) );
  INV_X1 U2778 ( .A(n4050), .ZN(n4123) );
  NOR2_X1 U2779 ( .A1(n3161), .A2(n3160), .ZN(n3241) );
  OR2_X1 U2780 ( .A1(n3295), .A2(n4561), .ZN(n3358) );
  NAND2_X1 U2781 ( .A1(n3241), .A2(REG3_REG_8__SCAN_IN), .ZN(n3295) );
  INV_X1 U2782 ( .A(n4006), .ZN(n2659) );
  INV_X1 U2783 ( .A(n4160), .ZN(n2660) );
  NAND2_X1 U2784 ( .A1(n2647), .A2(n2646), .ZN(n3523) );
  INV_X1 U2785 ( .A(n3510), .ZN(n2646) );
  NAND2_X1 U2786 ( .A1(n3110), .A2(REG3_REG_5__SCAN_IN), .ZN(n3161) );
  NAND2_X1 U2787 ( .A1(n2614), .A2(n2613), .ZN(n3984) );
  AOI21_X1 U2788 ( .B1(n2616), .B2(n2619), .A(n2514), .ZN(n2613) );
  AND2_X1 U2789 ( .A1(n3053), .A2(n3913), .ZN(n3069) );
  NAND2_X1 U2790 ( .A1(n2590), .A2(n2589), .ZN(n2983) );
  NAND2_X1 U2791 ( .A1(n2848), .A2(REG2_REG_2__SCAN_IN), .ZN(n2589) );
  OR2_X1 U2792 ( .A1(n2848), .A2(REG2_REG_2__SCAN_IN), .ZN(n2590) );
  OAI21_X1 U2793 ( .B1(n3184), .B2(n2987), .A(n2981), .ZN(n2787) );
  NAND2_X1 U2794 ( .A1(n5115), .A2(n2790), .ZN(n2935) );
  NAND2_X1 U2795 ( .A1(n2935), .A2(n2934), .ZN(n2933) );
  AND2_X1 U2796 ( .A1(n2737), .A2(n2736), .ZN(n2855) );
  XNOR2_X1 U2797 ( .A(n2792), .B(n5183), .ZN(n4260) );
  AND2_X1 U2798 ( .A1(n4269), .A2(n2865), .ZN(n4282) );
  NAND2_X1 U2799 ( .A1(n2864), .A2(n5074), .ZN(n2865) );
  NAND2_X1 U2800 ( .A1(n2943), .A2(n2517), .ZN(n2795) );
  INV_X1 U2801 ( .A(REG3_REG_9__SCAN_IN), .ZN(n4561) );
  INV_X1 U2802 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3512) );
  XNOR2_X1 U2803 ( .A(n2732), .B(n3373), .ZN(n4294) );
  NOR2_X1 U2804 ( .A1(n4294), .A2(n5218), .ZN(n4293) );
  NAND2_X1 U2805 ( .A1(n4300), .A2(n2802), .ZN(n3943) );
  INV_X1 U2806 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4726) );
  NOR2_X1 U2807 ( .A1(n4314), .A2(n5252), .ZN(n4313) );
  NAND2_X1 U2808 ( .A1(n4310), .A2(n2805), .ZN(n4324) );
  NAND2_X1 U2809 ( .A1(n4324), .A2(n4323), .ZN(n4322) );
  NOR2_X1 U2810 ( .A1(n4334), .A2(n2808), .ZN(n4342) );
  NAND2_X1 U2811 ( .A1(n4331), .A2(n2508), .ZN(n2727) );
  INV_X1 U2812 ( .A(n2608), .ZN(n4357) );
  OAI21_X1 U2813 ( .B1(n4334), .B2(n2609), .A(n2612), .ZN(n2608) );
  NAND2_X1 U2814 ( .A1(n4465), .A2(n4450), .ZN(n4449) );
  AND2_X1 U2815 ( .A1(n3781), .A2(n3780), .ZN(n4451) );
  OR2_X1 U2816 ( .A1(n4407), .A2(n3850), .ZN(n4443) );
  AND2_X1 U2817 ( .A1(n3707), .A2(n3706), .ZN(n4458) );
  OR2_X1 U2818 ( .A1(n4094), .A2(n3790), .ZN(n3707) );
  AND2_X1 U2819 ( .A1(n2502), .A2(n4891), .ZN(n2585) );
  NAND2_X1 U2820 ( .A1(n4921), .A2(n2502), .ZN(n4911) );
  NAND2_X1 U2821 ( .A1(n4989), .A2(n4988), .ZN(n4987) );
  AOI21_X1 U2822 ( .B1(n4984), .B2(n2671), .A(n2523), .ZN(n2670) );
  INV_X1 U2823 ( .A(n2512), .ZN(n2671) );
  OR2_X1 U2824 ( .A1(n3813), .A2(n4396), .ZN(n4955) );
  NOR2_X1 U2825 ( .A1(n4370), .A2(n3956), .ZN(n4989) );
  NAND2_X1 U2826 ( .A1(n2703), .A2(n2702), .ZN(n3668) );
  AOI21_X1 U2827 ( .B1(n2704), .B2(n2710), .A(n2501), .ZN(n2702) );
  NAND2_X1 U2828 ( .A1(n2586), .A2(n3667), .ZN(n3956) );
  INV_X1 U2829 ( .A(n3594), .ZN(n3593) );
  NAND2_X1 U2830 ( .A1(n3560), .A2(REG3_REG_15__SCAN_IN), .ZN(n3594) );
  NAND2_X1 U2831 ( .A1(n2570), .A2(n2569), .ZN(n2568) );
  NOR2_X1 U2832 ( .A1(n3828), .A2(n3670), .ZN(n2569) );
  AND2_X1 U2833 ( .A1(n3585), .A2(n3933), .ZN(n3603) );
  NAND2_X1 U2834 ( .A1(n3603), .A2(n3974), .ZN(n5292) );
  INV_X1 U2835 ( .A(n2570), .ZN(n3671) );
  INV_X1 U2836 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4759) );
  NAND2_X1 U2837 ( .A1(n2579), .A2(n3532), .ZN(n2578) );
  INV_X1 U2838 ( .A(n2580), .ZN(n2579) );
  NOR2_X1 U2839 ( .A1(n3368), .A2(n2580), .ZN(n3436) );
  INV_X1 U2840 ( .A(n4228), .ZN(n3467) );
  NAND2_X1 U2841 ( .A1(n3443), .A2(n4229), .ZN(n2701) );
  AND2_X1 U2842 ( .A1(n3884), .A2(n3550), .ZN(n3819) );
  OR2_X1 U2843 ( .A1(n3289), .A2(n3398), .ZN(n3368) );
  NOR2_X1 U2844 ( .A1(n3368), .A2(n3443), .ZN(n3388) );
  INV_X1 U2845 ( .A(n4229), .ZN(n3386) );
  AOI21_X1 U2846 ( .B1(n2558), .B2(n2560), .A(n2533), .ZN(n2556) );
  INV_X1 U2847 ( .A(n2559), .ZN(n2558) );
  NAND2_X1 U2848 ( .A1(n3251), .A2(n4138), .ZN(n3289) );
  NAND2_X1 U2849 ( .A1(n2557), .A2(n3874), .ZN(n3301) );
  NAND2_X1 U2850 ( .A1(n3238), .A2(n3840), .ZN(n2557) );
  NAND2_X1 U2851 ( .A1(n3907), .A2(n5121), .ZN(n5315) );
  AND2_X1 U2852 ( .A1(n3872), .A2(n3874), .ZN(n3840) );
  NAND2_X1 U2853 ( .A1(n3106), .A2(n3865), .ZN(n3157) );
  INV_X1 U2854 ( .A(n5315), .ZN(n5325) );
  INV_X1 U2855 ( .A(n3214), .ZN(n2576) );
  NAND2_X1 U2856 ( .A1(n2543), .A2(n3860), .ZN(n3207) );
  INV_X1 U2857 ( .A(n3108), .ZN(n3210) );
  MUX2_X1 U2858 ( .A(n2848), .B(DATAI_2_), .S(n3107), .Z(n3187) );
  AND2_X1 U2859 ( .A1(n3198), .A2(n3185), .ZN(n3216) );
  OR2_X1 U2860 ( .A1(n5296), .A2(n2961), .ZN(n5005) );
  NOR2_X1 U2861 ( .A1(n3116), .A2(n3079), .ZN(n3185) );
  INV_X1 U2862 ( .A(n5286), .ZN(n5127) );
  NAND2_X1 U2863 ( .A1(n4999), .A2(n5156), .ZN(n5258) );
  INV_X1 U2864 ( .A(IR_REG_27__SCAN_IN), .ZN(n4613) );
  INV_X1 U2865 ( .A(IR_REG_26__SCAN_IN), .ZN(n4806) );
  NOR2_X1 U2866 ( .A1(n2820), .A2(n2831), .ZN(n2583) );
  NAND2_X1 U2867 ( .A1(n2839), .A2(n2830), .ZN(n2831) );
  NAND2_X1 U2868 ( .A1(n2821), .A2(n2748), .ZN(n2756) );
  INV_X1 U2869 ( .A(IR_REG_7__SCAN_IN), .ZN(n4579) );
  OR2_X1 U2870 ( .A1(n2774), .A2(IR_REG_6__SCAN_IN), .ZN(n2770) );
  NAND2_X1 U2871 ( .A1(n3342), .A2(n2651), .ZN(n2648) );
  NAND2_X1 U2872 ( .A1(n3929), .A2(n3928), .ZN(n2615) );
  NAND2_X1 U2873 ( .A1(n4200), .A2(n4075), .ZN(n4153) );
  INV_X1 U2874 ( .A(n2647), .ZN(n3509) );
  INV_X1 U2875 ( .A(n3493), .ZN(n3515) );
  NAND2_X1 U2876 ( .A1(n2656), .A2(n4037), .ZN(n4159) );
  NAND2_X1 U2877 ( .A1(n2663), .A2(n2664), .ZN(n3622) );
  NAND2_X1 U2878 ( .A1(n5273), .A2(n3994), .ZN(n4002) );
  OAI21_X1 U2879 ( .B1(n4007), .B2(n2655), .A(n2652), .ZN(n4193) );
  AOI21_X1 U2880 ( .B1(n2658), .B2(n2654), .A(n2653), .ZN(n2652) );
  INV_X1 U2881 ( .A(n4049), .ZN(n2653) );
  INV_X1 U2882 ( .A(n4964), .ZN(n4956) );
  NOR2_X1 U2883 ( .A1(n3623), .A2(n2662), .ZN(n2661) );
  INV_X1 U2884 ( .A(n2664), .ZN(n2662) );
  INV_X1 U2885 ( .A(n5268), .ZN(n4216) );
  INV_X1 U2886 ( .A(n3187), .ZN(n3198) );
  NAND2_X1 U2887 ( .A1(n3342), .A2(n3330), .ZN(n3404) );
  INV_X1 U2888 ( .A(n5266), .ZN(n4214) );
  NOR2_X1 U2889 ( .A1(n2746), .A2(n4105), .ZN(n4106) );
  AND2_X1 U2890 ( .A1(n3069), .A2(n5068), .ZN(n5268) );
  INV_X1 U2891 ( .A(n5280), .ZN(n4183) );
  NAND2_X1 U2892 ( .A1(n3739), .A2(n3738), .ZN(n4930) );
  OR2_X1 U2893 ( .A1(n4913), .A2(n3790), .ZN(n3739) );
  NAND2_X1 U2894 ( .A1(n3729), .A2(n3728), .ZN(n4373) );
  OR2_X1 U2895 ( .A1(n4922), .A2(n3790), .ZN(n3729) );
  OR2_X1 U2896 ( .A1(n3747), .A2(n3746), .ZN(n4982) );
  OR2_X1 U2897 ( .A1(n2888), .A2(n2889), .ZN(n5104) );
  NAND2_X1 U2898 ( .A1(n4239), .A2(n4238), .ZN(n4237) );
  XNOR2_X1 U2899 ( .A(n2787), .B(n2588), .ZN(n4255) );
  NAND2_X1 U2900 ( .A1(n4255), .A2(REG2_REG_3__SCAN_IN), .ZN(n4254) );
  NOR2_X1 U2901 ( .A1(n2737), .A2(n2854), .ZN(n4251) );
  OR2_X1 U2902 ( .A1(n2738), .A2(n2854), .ZN(n4252) );
  INV_X1 U2903 ( .A(n2739), .ZN(n2738) );
  XNOR2_X1 U2904 ( .A(n2789), .B(n5164), .ZN(n5117) );
  OR2_X1 U2905 ( .A1(n2932), .A2(n2931), .ZN(n2717) );
  NOR2_X1 U2906 ( .A1(n4262), .A2(n2860), .ZN(n2942) );
  XNOR2_X1 U2907 ( .A(n2863), .B(n5074), .ZN(n4270) );
  NAND2_X1 U2908 ( .A1(n4270), .A2(REG1_REG_8__SCAN_IN), .ZN(n4269) );
  OAI211_X1 U2909 ( .C1(n4286), .C2(n2597), .A(REG2_REG_10__SCAN_IN), .B(n2594), .ZN(n4290) );
  NAND2_X1 U2910 ( .A1(n2499), .A2(n2605), .ZN(n2597) );
  AND2_X1 U2911 ( .A1(n2596), .A2(n2499), .ZN(n2595) );
  OAI211_X1 U2912 ( .C1(n4286), .C2(n2605), .A(n2499), .B(n2593), .ZN(n4291)
         );
  NAND2_X1 U2913 ( .A1(n4286), .A2(n2602), .ZN(n2593) );
  OAI21_X1 U2914 ( .B1(n4294), .B2(n2730), .A(n2729), .ZN(n3479) );
  NAND2_X1 U2915 ( .A1(n2731), .A2(REG1_REG_10__SCAN_IN), .ZN(n2730) );
  NAND2_X1 U2916 ( .A1(n2869), .A2(n2731), .ZN(n2729) );
  INV_X1 U2917 ( .A(n3480), .ZN(n2731) );
  NAND2_X1 U2918 ( .A1(n4301), .A2(REG2_REG_12__SCAN_IN), .ZN(n4300) );
  NOR2_X1 U2919 ( .A1(n4303), .A2(n2874), .ZN(n3940) );
  INV_X1 U2920 ( .A(n2872), .ZN(n2873) );
  NOR2_X1 U2921 ( .A1(n3940), .A2(n3939), .ZN(n3938) );
  XNOR2_X1 U2922 ( .A(n2804), .B(n2587), .ZN(n4311) );
  NOR2_X1 U2923 ( .A1(n4313), .A2(n2879), .ZN(n4321) );
  NAND2_X1 U2924 ( .A1(n2688), .A2(n4409), .ZN(n2687) );
  OAI21_X1 U2925 ( .B1(n2693), .B2(n2688), .A(n2685), .ZN(n2684) );
  NAND2_X1 U2926 ( .A1(n2689), .A2(n4382), .ZN(n4421) );
  OR2_X1 U2927 ( .A1(n4428), .A2(n2526), .ZN(n4438) );
  AND2_X1 U2928 ( .A1(n4430), .A2(n5286), .ZN(n2564) );
  OAI21_X1 U2929 ( .B1(n4880), .B2(n2679), .A(n2677), .ZN(n4457) );
  NAND2_X1 U2930 ( .A1(n2681), .A2(n2680), .ZN(n4475) );
  AND2_X1 U2931 ( .A1(n2681), .A2(n2506), .ZN(n4474) );
  NAND2_X1 U2932 ( .A1(n4880), .A2(n4376), .ZN(n2681) );
  AND2_X1 U2933 ( .A1(n2694), .A2(n2695), .ZN(n4899) );
  AND2_X1 U2934 ( .A1(n2698), .A2(n2500), .ZN(n4920) );
  NAND2_X1 U2935 ( .A1(n4935), .A2(n4936), .ZN(n2698) );
  NAND2_X1 U2936 ( .A1(n4985), .A2(n4984), .ZN(n4983) );
  NAND2_X1 U2937 ( .A1(n2673), .A2(n2512), .ZN(n4985) );
  NAND2_X1 U2938 ( .A1(n4369), .A2(n4368), .ZN(n2673) );
  NAND2_X1 U2939 ( .A1(n2706), .A2(n2708), .ZN(n5291) );
  OR2_X1 U2940 ( .A1(n3576), .A2(n2710), .ZN(n2706) );
  NAND2_X1 U2941 ( .A1(n2707), .A2(n2712), .ZN(n3656) );
  NAND2_X1 U2942 ( .A1(n3576), .A2(n2713), .ZN(n2707) );
  AOI21_X1 U2943 ( .B1(n3576), .B2(n3541), .A(n2496), .ZN(n3591) );
  NAND2_X1 U2944 ( .A1(n3354), .A2(n3353), .ZN(n3385) );
  INV_X1 U2945 ( .A(n3288), .ZN(n3354) );
  OR2_X1 U2946 ( .A1(n5005), .A2(n3090), .ZN(n4991) );
  XNOR2_X1 U2947 ( .A(n3080), .B(n3855), .ZN(n3087) );
  INV_X1 U2948 ( .A(n4991), .ZN(n5303) );
  NAND2_X1 U2949 ( .A1(n2563), .A2(n2561), .ZN(n5052) );
  INV_X1 U2950 ( .A(n4438), .ZN(n2563) );
  INV_X1 U2951 ( .A(n2562), .ZN(n2561) );
  OAI21_X1 U2952 ( .B1(n5011), .B2(n5297), .A(n5010), .ZN(n2562) );
  AND2_X2 U2953 ( .A1(n5050), .A2(n5049), .ZN(n5347) );
  AND2_X1 U2954 ( .A1(n2830), .A2(n4811), .ZN(n2917) );
  XNOR2_X1 U2955 ( .A(n2835), .B(IR_REG_26__SCAN_IN), .ZN(n5069) );
  XNOR2_X1 U2956 ( .A(n2843), .B(n2830), .ZN(n3823) );
  OAI21_X1 U2957 ( .B1(n2957), .B2(IR_REG_31__SCAN_IN), .A(n2637), .ZN(n2636)
         );
  NAND2_X1 U2958 ( .A1(n2956), .A2(n2639), .ZN(n2638) );
  XNOR2_X1 U2959 ( .A(n2591), .B(IR_REG_2__SCAN_IN), .ZN(n2848) );
  NAND2_X1 U2960 ( .A1(n2592), .A2(IR_REG_31__SCAN_IN), .ZN(n2591) );
  INV_X1 U2961 ( .A(n2783), .ZN(n2592) );
  NAND2_X1 U2962 ( .A1(n2722), .A2(n2720), .ZN(n2850) );
  NAND2_X1 U2963 ( .A1(n2721), .A2(IR_REG_1__SCAN_IN), .ZN(n2720) );
  NAND2_X1 U2964 ( .A1(n2628), .A2(n2622), .ZN(n2621) );
  NAND2_X1 U2965 ( .A1(n2718), .A2(n4362), .ZN(n2894) );
  INV_X1 U2966 ( .A(n3056), .ZN(n2923) );
  AND2_X1 U2967 ( .A1(n3566), .A2(n3649), .ZN(n2496) );
  NOR2_X1 U2968 ( .A1(n4108), .A2(n4100), .ZN(n4178) );
  AND2_X1 U2969 ( .A1(n2505), .A2(n2749), .ZN(n2498) );
  INV_X1 U2970 ( .A(n4984), .ZN(n2672) );
  INV_X1 U2971 ( .A(n4285), .ZN(n2603) );
  AND2_X1 U2972 ( .A1(n2598), .A2(n2599), .ZN(n2499) );
  INV_X1 U2973 ( .A(n3855), .ZN(n2567) );
  OR2_X1 U2974 ( .A1(n4222), .A2(n4938), .ZN(n2500) );
  AND2_X1 U2975 ( .A1(n2716), .A2(n5294), .ZN(n2501) );
  INV_X1 U2976 ( .A(n3373), .ZN(n2601) );
  AND2_X1 U2977 ( .A1(n4384), .A2(n4912), .ZN(n2502) );
  NAND2_X1 U2978 ( .A1(n3402), .A2(n3401), .ZN(n2503) );
  INV_X1 U2979 ( .A(n2566), .ZN(n2914) );
  NAND4_X1 U2980 ( .A1(n2582), .A2(n2497), .A3(n2765), .A4(n2830), .ZN(n2566)
         );
  NAND2_X1 U2981 ( .A1(n2832), .A2(n5069), .ZN(n2958) );
  AND4_X1 U2982 ( .A1(n4591), .A2(n4587), .A3(n4775), .A4(n4781), .ZN(n2504)
         );
  AND2_X1 U2983 ( .A1(n2748), .A2(n4591), .ZN(n2505) );
  MUX2_X1 U2984 ( .A(n5113), .B(DATAI_4_), .S(n3107), .Z(n3266) );
  INV_X1 U2985 ( .A(n3266), .ZN(n3281) );
  NAND2_X1 U2986 ( .A1(n4479), .A2(n4891), .ZN(n2506) );
  NOR2_X1 U2987 ( .A1(n4179), .A2(n4181), .ZN(n2507) );
  NAND2_X1 U2988 ( .A1(n2783), .A2(n4766), .ZN(n2779) );
  AND2_X1 U2989 ( .A1(n2883), .A2(n2728), .ZN(n2508) );
  NAND2_X1 U2990 ( .A1(n2584), .A2(IR_REG_31__SCAN_IN), .ZN(n2835) );
  NOR2_X1 U2991 ( .A1(n4321), .A2(n4320), .ZN(n2509) );
  XOR2_X1 U2992 ( .A(n2816), .B(n2815), .Z(n2510) );
  INV_X1 U2993 ( .A(n2610), .ZN(n2609) );
  NOR2_X1 U2994 ( .A1(n2808), .A2(n2611), .ZN(n2610) );
  AND2_X1 U2995 ( .A1(n2819), .A2(n4597), .ZN(n2511) );
  INV_X1 U2996 ( .A(n3443), .ZN(n2581) );
  INV_X1 U2997 ( .A(n4459), .ZN(n2675) );
  AOI21_X1 U2998 ( .B1(n4193), .B2(n4190), .A(n4189), .ZN(n4166) );
  INV_X1 U2999 ( .A(n3843), .ZN(n2715) );
  OR2_X1 U3000 ( .A1(n4371), .A2(n4370), .ZN(n2512) );
  OR2_X1 U3001 ( .A1(n4930), .A2(n4375), .ZN(n2513) );
  INV_X1 U3002 ( .A(n2605), .ZN(n2604) );
  NAND2_X1 U3003 ( .A1(n4007), .A2(n4006), .ZN(n4039) );
  XOR2_X1 U3004 ( .A(n3969), .B(n3490), .Z(n2514) );
  INV_X1 U3005 ( .A(n3526), .ZN(n3532) );
  INV_X1 U3006 ( .A(n4093), .ZN(n2629) );
  INV_X1 U3007 ( .A(n4409), .ZN(n2693) );
  INV_X1 U3008 ( .A(n4368), .ZN(n2669) );
  AND2_X1 U3009 ( .A1(n2581), .A2(n3386), .ZN(n2515) );
  NAND2_X1 U3010 ( .A1(n3986), .A2(n3985), .ZN(n5269) );
  NAND2_X1 U3011 ( .A1(n2821), .A2(n2498), .ZN(n2752) );
  AND2_X1 U3012 ( .A1(n2695), .A2(n4904), .ZN(n2516) );
  INV_X1 U3013 ( .A(n4222), .ZN(n4960) );
  NAND2_X1 U3014 ( .A1(n3722), .A2(n3721), .ZN(n4222) );
  OR2_X1 U3015 ( .A1(n5191), .A2(n3253), .ZN(n2517) );
  NAND2_X1 U3016 ( .A1(n2698), .A2(n2697), .ZN(n2518) );
  NOR2_X1 U3017 ( .A1(n5283), .A2(n3974), .ZN(n2519) );
  NOR2_X1 U3018 ( .A1(n4458), .A2(n4478), .ZN(n2520) );
  AND2_X1 U3019 ( .A1(n2615), .A2(n3930), .ZN(n2521) );
  AND2_X1 U3020 ( .A1(n2656), .A2(n2654), .ZN(n2522) );
  AND2_X1 U3021 ( .A1(n4194), .A2(n4988), .ZN(n2523) );
  NOR2_X1 U3022 ( .A1(n3921), .A2(n4224), .ZN(n2524) );
  INV_X1 U3023 ( .A(n2655), .ZN(n2654) );
  NAND2_X1 U3024 ( .A1(n2660), .A2(n4037), .ZN(n2655) );
  NOR2_X1 U3025 ( .A1(n4383), .A2(n4422), .ZN(n2525) );
  INV_X1 U3026 ( .A(n2658), .ZN(n2657) );
  OR2_X1 U3027 ( .A1(n4038), .A2(n2659), .ZN(n2658) );
  INV_X1 U3028 ( .A(n4379), .ZN(n4380) );
  NOR2_X1 U3029 ( .A1(n4464), .A2(n4381), .ZN(n4379) );
  AND2_X1 U3030 ( .A1(n4921), .A2(n4384), .ZN(n4910) );
  OR2_X1 U3031 ( .A1(n4429), .A2(n2564), .ZN(n2526) );
  OR2_X1 U3032 ( .A1(n4982), .A2(n4956), .ZN(n2527) );
  INV_X1 U3033 ( .A(IR_REG_31__SCAN_IN), .ZN(n5064) );
  NOR2_X1 U3034 ( .A1(n4093), .A2(n4098), .ZN(n2528) );
  AND2_X1 U3035 ( .A1(n4080), .A2(n4075), .ZN(n2529) );
  NAND2_X1 U3036 ( .A1(n2821), .A2(n2505), .ZN(n2530) );
  INV_X1 U3037 ( .A(n2862), .ZN(n2735) );
  AND2_X1 U3038 ( .A1(n3239), .A2(REG1_REG_7__SCAN_IN), .ZN(n2862) );
  OR2_X1 U3039 ( .A1(n2515), .A2(n2699), .ZN(n2531) );
  OR2_X1 U3040 ( .A1(n2630), .A2(n2626), .ZN(n2532) );
  NAND3_X1 U3041 ( .A1(n2640), .A2(n2638), .A3(n2636), .ZN(n2997) );
  INV_X1 U3042 ( .A(n4223), .ZN(n2716) );
  NAND2_X1 U3043 ( .A1(n2663), .A2(n2661), .ZN(n3643) );
  INV_X1 U3044 ( .A(n4372), .ZN(n4988) );
  NAND2_X1 U3045 ( .A1(n2648), .A2(n2649), .ZN(n3507) );
  INV_X1 U3046 ( .A(n3134), .ZN(n3138) );
  AND2_X1 U3047 ( .A1(n4231), .A2(n4138), .ZN(n2533) );
  NAND2_X1 U3048 ( .A1(n2822), .A2(IR_REG_31__SCAN_IN), .ZN(n2833) );
  INV_X1 U3049 ( .A(n3928), .ZN(n2618) );
  NOR2_X1 U3050 ( .A1(n3276), .A2(n3316), .ZN(n2534) );
  NAND2_X1 U3051 ( .A1(n5267), .A2(n3974), .ZN(n2535) );
  NOR2_X1 U3052 ( .A1(n4293), .A2(n2869), .ZN(n2536) );
  INV_X1 U3053 ( .A(n2586), .ZN(n5293) );
  NOR2_X1 U3054 ( .A1(n5292), .A2(n5265), .ZN(n2586) );
  INV_X1 U3055 ( .A(n2577), .ZN(n3474) );
  NOR2_X1 U3056 ( .A1(n3368), .A2(n2578), .ZN(n2577) );
  XNOR2_X1 U3057 ( .A(n2841), .B(n2840), .ZN(n2845) );
  INV_X1 U3058 ( .A(n3547), .ZN(n2587) );
  OR2_X1 U3059 ( .A1(n2612), .A2(n4358), .ZN(n2537) );
  NAND2_X1 U3060 ( .A1(n2576), .A2(n3281), .ZN(n3229) );
  INV_X1 U3061 ( .A(n3229), .ZN(n2575) );
  NOR2_X1 U3062 ( .A1(n2942), .A2(n2941), .ZN(n2538) );
  OR2_X1 U3063 ( .A1(n4328), .A2(n2806), .ZN(n2539) );
  INV_X1 U3064 ( .A(n2881), .ZN(n2726) );
  AND2_X1 U3065 ( .A1(n5073), .A2(REG1_REG_15__SCAN_IN), .ZN(n2881) );
  INV_X1 U3066 ( .A(IR_REG_0__SCAN_IN), .ZN(n2572) );
  XNOR2_X1 U3067 ( .A(n2782), .B(IR_REG_3__SCAN_IN), .ZN(n4248) );
  INV_X1 U3068 ( .A(n4248), .ZN(n2588) );
  AND2_X1 U3069 ( .A1(n5071), .A2(REG2_REG_18__SCAN_IN), .ZN(n2540) );
  XOR2_X1 U3070 ( .A(n2961), .B(REG1_REG_19__SCAN_IN), .Z(n2541) );
  NAND2_X1 U3071 ( .A1(n2543), .A2(n2542), .ZN(n3183) );
  OR2_X1 U3072 ( .A1(n3179), .A2(n3837), .ZN(n2542) );
  NAND2_X1 U3073 ( .A1(n3179), .A2(n3837), .ZN(n2543) );
  OR2_X2 U3074 ( .A1(n4460), .A2(n4459), .ZN(n2554) );
  INV_X1 U3075 ( .A(n4407), .ZN(n2552) );
  NAND2_X1 U3076 ( .A1(n3238), .A2(n2558), .ZN(n2555) );
  NAND2_X1 U3077 ( .A1(n2555), .A2(n2556), .ZN(n3356) );
  NAND3_X1 U3078 ( .A1(n2582), .A2(n2497), .A3(n2765), .ZN(n2916) );
  NAND2_X1 U3079 ( .A1(n3107), .A2(DATAI_1_), .ZN(n2573) );
  INV_X1 U3080 ( .A(n2820), .ZN(n2582) );
  NAND3_X1 U3081 ( .A1(n2497), .A2(n2583), .A3(n2765), .ZN(n2584) );
  AND2_X1 U3082 ( .A1(n2765), .A2(n4776), .ZN(n2821) );
  NAND2_X1 U3083 ( .A1(n2835), .A2(n4806), .ZN(n2836) );
  NAND2_X1 U3084 ( .A1(n4286), .A2(n2595), .ZN(n2594) );
  NAND2_X1 U3085 ( .A1(n4286), .A2(n4285), .ZN(n4284) );
  NAND2_X1 U3086 ( .A1(n4284), .A2(n2743), .ZN(n2798) );
  NAND2_X1 U3087 ( .A1(n3373), .A2(n2743), .ZN(n2605) );
  NAND2_X1 U3088 ( .A1(n2921), .A2(IR_REG_31__SCAN_IN), .ZN(n2922) );
  OAI21_X2 U3089 ( .B1(n4883), .B2(n4403), .A(n4402), .ZN(n4476) );
  NAND2_X1 U3090 ( .A1(n2786), .A2(n2785), .ZN(n2981) );
  OAI21_X1 U3091 ( .B1(n3929), .B2(n2619), .A(n2616), .ZN(n3971) );
  NAND2_X1 U3092 ( .A1(n3929), .A2(n2616), .ZN(n2614) );
  OR2_X1 U3093 ( .A1(n4179), .A2(n2532), .ZN(n2623) );
  NAND2_X1 U3094 ( .A1(n4178), .A2(n2629), .ZN(n2620) );
  OAI211_X1 U3095 ( .C1(n4178), .C2(n2528), .A(n2620), .B(n2628), .ZN(n2627)
         );
  NAND4_X1 U3096 ( .A1(n2627), .A2(n2624), .A3(n2623), .A4(n2621), .ZN(U3222)
         );
  NAND3_X1 U3097 ( .A1(n4179), .A2(n4182), .A3(n2625), .ZN(n2624) );
  NAND2_X1 U3098 ( .A1(n2632), .A2(n2783), .ZN(n2768) );
  NAND4_X1 U3099 ( .A1(n2633), .A2(n4571), .A3(n2635), .A4(n2769), .ZN(n2634)
         );
  NAND2_X2 U3100 ( .A1(n2997), .A2(n5121), .ZN(n5296) );
  NAND3_X1 U3101 ( .A1(n3342), .A2(n2651), .A3(n3506), .ZN(n2641) );
  INV_X1 U3102 ( .A(n3403), .ZN(n2650) );
  INV_X1 U3103 ( .A(n2649), .ZN(n2643) );
  NAND3_X1 U3104 ( .A1(n3986), .A2(n3991), .A3(n3985), .ZN(n5273) );
  NAND2_X1 U3105 ( .A1(n4200), .A2(n2529), .ZN(n4151) );
  NAND2_X1 U3106 ( .A1(n4369), .A2(n2668), .ZN(n2667) );
  NAND2_X1 U3107 ( .A1(n2667), .A2(n2670), .ZN(n4952) );
  NAND2_X1 U3108 ( .A1(n4880), .A2(n2677), .ZN(n2676) );
  NAND2_X1 U3109 ( .A1(n4440), .A2(n2683), .ZN(n2682) );
  OAI211_X1 U3110 ( .C1(n4440), .C2(n2687), .A(n2684), .B(n2682), .ZN(n5000)
         );
  NAND2_X1 U3111 ( .A1(n4440), .A2(n4380), .ZN(n2689) );
  OAI21_X1 U3112 ( .B1(n3288), .B2(n2531), .A(n2701), .ZN(n2700) );
  INV_X1 U3113 ( .A(n2700), .ZN(n3470) );
  NAND2_X1 U3114 ( .A1(n3576), .A2(n2704), .ZN(n2703) );
  INV_X1 U3115 ( .A(n2717), .ZN(n2930) );
  NOR2_X1 U3116 ( .A1(n5109), .A2(n2856), .ZN(n2932) );
  INV_X1 U3117 ( .A(IR_REG_1__SCAN_IN), .ZN(n2723) );
  NAND3_X1 U3118 ( .A1(n2723), .A2(IR_REG_31__SCAN_IN), .A3(IR_REG_0__SCAN_IN), 
        .ZN(n2722) );
  OR2_X1 U3119 ( .A1(n2879), .A2(n2881), .ZN(n2725) );
  NAND2_X1 U3120 ( .A1(n2727), .A2(n2884), .ZN(n4363) );
  NAND2_X1 U3121 ( .A1(n4331), .A2(n2883), .ZN(n4351) );
  INV_X1 U3122 ( .A(n2727), .ZN(n4349) );
  INV_X1 U3123 ( .A(n4350), .ZN(n2728) );
  INV_X1 U3124 ( .A(n2868), .ZN(n2732) );
  INV_X1 U3125 ( .A(n2854), .ZN(n2736) );
  NAND2_X1 U3126 ( .A1(n3056), .A2(REG1_REG_4__SCAN_IN), .ZN(n3059) );
  NAND2_X1 U3127 ( .A1(n3056), .A2(REG1_REG_0__SCAN_IN), .ZN(n2953) );
  INV_X1 U3128 ( .A(n3971), .ZN(n3970) );
  INV_X1 U3129 ( .A(n2877), .ZN(n2878) );
  INV_X1 U3130 ( .A(n2858), .ZN(n2859) );
  XNOR2_X1 U3131 ( .A(n2858), .B(n3153), .ZN(n4263) );
  NAND2_X2 U3132 ( .A1(n3343), .A2(n3344), .ZN(n3342) );
  AOI21_X1 U3133 ( .B1(n3108), .B2(n3026), .A(n3267), .ZN(n3312) );
  INV_X1 U3134 ( .A(n3026), .ZN(n3324) );
  NOR2_X1 U3135 ( .A1(n3123), .A2(n3138), .ZN(n2740) );
  AND2_X1 U3136 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2741)
         );
  NAND2_X1 U3137 ( .A1(n3144), .A2(n3143), .ZN(n3228) );
  AND2_X1 U3138 ( .A1(n2918), .A2(n2917), .ZN(n2742) );
  OR2_X1 U3139 ( .A1(n5206), .A2(n2797), .ZN(n2743) );
  INV_X1 U3140 ( .A(n3838), .ZN(n3286) );
  OR2_X1 U3141 ( .A1(n3004), .A2(n3024), .ZN(n2744) );
  AND2_X1 U3142 ( .A1(n4122), .A2(n4121), .ZN(n2745) );
  NAND2_X1 U3143 ( .A1(n3285), .A2(n3284), .ZN(n3287) );
  AND3_X1 U3144 ( .A1(n4099), .A2(n4103), .A3(n4098), .ZN(n2746) );
  NAND2_X1 U3145 ( .A1(n3698), .A2(n3697), .ZN(n4481) );
  INV_X1 U3146 ( .A(IR_REG_13__SCAN_IN), .ZN(n4591) );
  NOR2_X1 U3147 ( .A1(n3467), .A2(n3515), .ZN(n3468) );
  INV_X1 U31480 ( .A(IR_REG_21__SCAN_IN), .ZN(n2830) );
  INV_X1 U31490 ( .A(n3194), .ZN(n3028) );
  INV_X1 U3150 ( .A(n3701), .ZN(n3691) );
  INV_X1 U3151 ( .A(n3745), .ZN(n3690) );
  NAND2_X1 U3152 ( .A1(n3120), .A2(n3119), .ZN(n3137) );
  AND2_X1 U3153 ( .A1(n3121), .A2(n3205), .ZN(n3135) );
  NAND2_X1 U3154 ( .A1(n4024), .A2(n3198), .ZN(n3205) );
  OR2_X1 U3155 ( .A1(n3504), .A2(n3503), .ZN(n3505) );
  INV_X1 U3156 ( .A(n3749), .ZN(n3688) );
  NAND2_X1 U3157 ( .A1(n3699), .A2(REG3_REG_25__SCAN_IN), .ZN(n3701) );
  NOR2_X1 U3158 ( .A1(n3733), .A2(n4184), .ZN(n3699) );
  INV_X1 U3159 ( .A(n4203), .ZN(n4071) );
  OR2_X1 U3160 ( .A1(n3779), .A2(n4725), .ZN(n3781) );
  NOR2_X1 U3161 ( .A1(n3358), .A2(n3512), .ZN(n3376) );
  INV_X1 U3162 ( .A(n5066), .ZN(n2925) );
  NOR2_X1 U3163 ( .A1(n4280), .A2(n2867), .ZN(n2868) );
  AND2_X1 U3164 ( .A1(n4383), .A2(n4431), .ZN(n4408) );
  AND2_X1 U3165 ( .A1(n4373), .A2(n4929), .ZN(n4374) );
  AND2_X1 U3166 ( .A1(n4222), .A2(n4944), .ZN(n4901) );
  NAND2_X1 U3167 ( .A1(n3658), .A2(REG3_REG_17__SCAN_IN), .ZN(n3674) );
  INV_X1 U3168 ( .A(n3809), .ZN(n4404) );
  INV_X1 U3169 ( .A(IR_REG_20__SCAN_IN), .ZN(n2957) );
  NAND2_X1 U3170 ( .A1(n3148), .A2(n3147), .ZN(n3257) );
  INV_X1 U3171 ( .A(n3921), .ZN(n3933) );
  NAND2_X1 U3172 ( .A1(n3688), .A2(REG3_REG_19__SCAN_IN), .ZN(n3751) );
  NAND2_X1 U3173 ( .A1(n3426), .A2(REG3_REG_12__SCAN_IN), .ZN(n3455) );
  OR2_X1 U3174 ( .A1(n3455), .A2(n4759), .ZN(n3542) );
  AND2_X1 U3175 ( .A1(n3376), .A2(REG3_REG_11__SCAN_IN), .ZN(n3426) );
  OR2_X1 U3176 ( .A1(n3674), .A2(n4014), .ZN(n3749) );
  OR2_X1 U3177 ( .A1(n4434), .A2(n3790), .ZN(n3778) );
  INV_X1 U3178 ( .A(n5206), .ZN(n3355) );
  XNOR2_X1 U3179 ( .A(n2877), .B(n3547), .ZN(n4314) );
  NAND2_X1 U3180 ( .A1(n4481), .A2(n4377), .ZN(n4378) );
  OR2_X1 U3181 ( .A1(n4373), .A2(n4384), .ZN(n4903) );
  AND2_X1 U3182 ( .A1(n4997), .A2(n3858), .ZN(n3082) );
  NAND2_X1 U3183 ( .A1(n3593), .A2(REG3_REG_16__SCAN_IN), .ZN(n3659) );
  INV_X1 U3184 ( .A(n4957), .ZN(n5282) );
  AND2_X1 U3185 ( .A1(n3075), .A2(n3823), .ZN(n5121) );
  AND2_X1 U3186 ( .A1(n3760), .A2(n3761), .ZN(n3843) );
  AND2_X1 U3187 ( .A1(n3554), .A2(n3461), .ZN(n3820) );
  INV_X1 U3188 ( .A(n3408), .ZN(n4138) );
  OR2_X1 U3189 ( .A1(n2776), .A2(n5064), .ZN(n2777) );
  INV_X1 U3190 ( .A(n4909), .ZN(n4479) );
  AND2_X1 U3191 ( .A1(n3710), .A2(n3709), .ZN(n4893) );
  INV_X1 U3192 ( .A(n3109), .ZN(n3790) );
  AND2_X1 U3193 ( .A1(n3778), .A2(n3777), .ZN(n4383) );
  INV_X1 U3194 ( .A(n2981), .ZN(n2985) );
  INV_X1 U3195 ( .A(n2977), .ZN(n2978) );
  NAND2_X1 U3196 ( .A1(n3118), .A2(n3117), .ZN(n3178) );
  AND2_X1 U3197 ( .A1(n3048), .A2(n3047), .ZN(n5009) );
  INV_X1 U3198 ( .A(n5258), .ZN(n5297) );
  INV_X1 U3199 ( .A(n5009), .ZN(n5049) );
  NOR2_X1 U3200 ( .A1(n5008), .A2(n5007), .ZN(n5050) );
  XNOR2_X1 U3201 ( .A(n2777), .B(IR_REG_5__SCAN_IN), .ZN(n3145) );
  AND2_X1 U3202 ( .A1(n2890), .A2(n2889), .ZN(n5107) );
  INV_X1 U3203 ( .A(n3116), .ZN(n4029) );
  INV_X1 U3204 ( .A(n4383), .ZN(n4448) );
  INV_X1 U3205 ( .A(n4458), .ZN(n4889) );
  NAND2_X1 U3206 ( .A1(n5138), .A2(n3155), .ZN(n5307) );
  NAND2_X2 U3207 ( .A1(n3095), .A2(n4991), .ZN(n5138) );
  INV_X1 U3208 ( .A(n5343), .ZN(n5341) );
  INV_X1 U3209 ( .A(n5347), .ZN(n5344) );
  INV_X1 U32100 ( .A(n5095), .ZN(n5099) );
  AND2_X1 U32110 ( .A1(n3064), .A2(STATE_REG_SCAN_IN), .ZN(n2900) );
  INV_X1 U32120 ( .A(n4235), .ZN(U4043) );
  INV_X2 U32130 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U32140 ( .A(IR_REG_5__SCAN_IN), .ZN(n2769) );
  NOR2_X1 U32150 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2819) );
  INV_X1 U32160 ( .A(n2812), .ZN(n2750) );
  NAND2_X1 U32170 ( .A1(n2750), .A2(IR_REG_31__SCAN_IN), .ZN(n2751) );
  XNOR2_X1 U32180 ( .A(n2751), .B(IR_REG_18__SCAN_IN), .ZN(n5071) );
  NAND2_X1 U32190 ( .A1(n2752), .A2(IR_REG_31__SCAN_IN), .ZN(n2754) );
  NAND2_X1 U32200 ( .A1(n2754), .A2(n4597), .ZN(n2809) );
  NAND2_X1 U32210 ( .A1(n2809), .A2(IR_REG_31__SCAN_IN), .ZN(n2753) );
  XNOR2_X1 U32220 ( .A(n2753), .B(IR_REG_16__SCAN_IN), .ZN(n3654) );
  INV_X1 U32230 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2806) );
  XNOR2_X1 U32240 ( .A(n2754), .B(IR_REG_15__SCAN_IN), .ZN(n5073) );
  INV_X1 U32250 ( .A(n5073), .ZN(n4328) );
  AOI22_X1 U32260 ( .A1(n5073), .A2(REG2_REG_15__SCAN_IN), .B1(n2806), .B2(
        n4328), .ZN(n4323) );
  NAND2_X1 U32270 ( .A1(n2530), .A2(IR_REG_31__SCAN_IN), .ZN(n2755) );
  XNOR2_X1 U32280 ( .A(n2755), .B(IR_REG_14__SCAN_IN), .ZN(n3547) );
  NAND2_X1 U32290 ( .A1(n2756), .A2(IR_REG_31__SCAN_IN), .ZN(n2757) );
  XNOR2_X1 U32300 ( .A(n2757), .B(IR_REG_13__SCAN_IN), .ZN(n3540) );
  NAND2_X1 U32310 ( .A1(n3540), .A2(REG2_REG_13__SCAN_IN), .ZN(n2803) );
  INV_X1 U32320 ( .A(REG2_REG_13__SCAN_IN), .ZN(n2758) );
  INV_X1 U32330 ( .A(n3540), .ZN(n5240) );
  AOI22_X1 U32340 ( .A1(n3540), .A2(REG2_REG_13__SCAN_IN), .B1(n2758), .B2(
        n5240), .ZN(n3942) );
  NAND2_X1 U32350 ( .A1(n2821), .A2(n4775), .ZN(n2759) );
  NAND2_X1 U32360 ( .A1(n2759), .A2(IR_REG_31__SCAN_IN), .ZN(n2762) );
  NAND2_X1 U32370 ( .A1(n2762), .A2(n4781), .ZN(n2760) );
  NAND2_X1 U32380 ( .A1(n2760), .A2(IR_REG_31__SCAN_IN), .ZN(n2761) );
  XNOR2_X1 U32390 ( .A(n2761), .B(IR_REG_12__SCAN_IN), .ZN(n3463) );
  XNOR2_X1 U32400 ( .A(n2762), .B(IR_REG_11__SCAN_IN), .ZN(n3423) );
  NAND2_X1 U32410 ( .A1(n3423), .A2(REG2_REG_11__SCAN_IN), .ZN(n2800) );
  INV_X1 U32420 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2763) );
  INV_X1 U32430 ( .A(n3423), .ZN(n5222) );
  AOI22_X1 U32440 ( .A1(n3423), .A2(REG2_REG_11__SCAN_IN), .B1(n2763), .B2(
        n5222), .ZN(n3482) );
  OR2_X1 U32450 ( .A1(n2821), .A2(n5064), .ZN(n2764) );
  XNOR2_X1 U32460 ( .A(n2764), .B(IR_REG_10__SCAN_IN), .ZN(n3373) );
  NOR2_X1 U32470 ( .A1(n2765), .A2(n5064), .ZN(n2766) );
  MUX2_X1 U32480 ( .A(n5064), .B(n2766), .S(IR_REG_9__SCAN_IN), .Z(n2767) );
  OR2_X1 U32490 ( .A1(n2767), .A2(n2821), .ZN(n5206) );
  INV_X1 U32500 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2797) );
  AOI22_X1 U32510 ( .A1(n3355), .A2(REG2_REG_9__SCAN_IN), .B1(n2797), .B2(
        n5206), .ZN(n4285) );
  NAND2_X1 U32520 ( .A1(n2776), .A2(n2769), .ZN(n2774) );
  NAND2_X1 U32530 ( .A1(n2770), .A2(IR_REG_31__SCAN_IN), .ZN(n2773) );
  NAND2_X1 U32540 ( .A1(n2773), .A2(n4579), .ZN(n2771) );
  NAND2_X1 U32550 ( .A1(n2771), .A2(IR_REG_31__SCAN_IN), .ZN(n2772) );
  XNOR2_X1 U32560 ( .A(n2772), .B(IR_REG_8__SCAN_IN), .ZN(n5074) );
  XNOR2_X1 U32570 ( .A(n2773), .B(IR_REG_7__SCAN_IN), .ZN(n3239) );
  INV_X1 U32580 ( .A(n3239), .ZN(n5191) );
  INV_X1 U32590 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U32600 ( .A1(n3239), .A2(REG2_REG_7__SCAN_IN), .B1(n3253), .B2(
        n5191), .ZN(n2944) );
  NAND2_X1 U32610 ( .A1(n2774), .A2(IR_REG_31__SCAN_IN), .ZN(n2775) );
  XNOR2_X1 U32620 ( .A(n2775), .B(IR_REG_6__SCAN_IN), .ZN(n3153) );
  NAND2_X1 U32630 ( .A1(n3145), .A2(REG2_REG_5__SCAN_IN), .ZN(n2791) );
  INV_X1 U32640 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2778) );
  INV_X1 U32650 ( .A(n3145), .ZN(n5174) );
  AOI22_X1 U32660 ( .A1(n3145), .A2(REG2_REG_5__SCAN_IN), .B1(n2778), .B2(
        n5174), .ZN(n2934) );
  NAND2_X1 U32670 ( .A1(n2779), .A2(IR_REG_31__SCAN_IN), .ZN(n2782) );
  NAND2_X1 U32680 ( .A1(n2782), .A2(n4571), .ZN(n2780) );
  NAND2_X1 U32690 ( .A1(n2780), .A2(IR_REG_31__SCAN_IN), .ZN(n2781) );
  XNOR2_X1 U32700 ( .A(n2781), .B(IR_REG_4__SCAN_IN), .ZN(n5113) );
  INV_X1 U32710 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3184) );
  INV_X1 U32720 ( .A(n2848), .ZN(n2987) );
  INV_X1 U32730 ( .A(n2983), .ZN(n2786) );
  INV_X1 U32740 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2784) );
  MUX2_X1 U32750 ( .A(REG2_REG_1__SCAN_IN), .B(n2784), .S(n2850), .Z(n4242) );
  NAND3_X1 U32760 ( .A1(n4242), .A2(REG2_REG_0__SCAN_IN), .A3(
        IR_REG_0__SCAN_IN), .ZN(n4241) );
  NAND2_X1 U32770 ( .A1(n2850), .A2(REG2_REG_1__SCAN_IN), .ZN(n2982) );
  NAND2_X1 U32780 ( .A1(n4241), .A2(n2982), .ZN(n2785) );
  NAND2_X1 U32790 ( .A1(n4248), .A2(n2787), .ZN(n2788) );
  NAND2_X1 U32800 ( .A1(n5113), .A2(n2789), .ZN(n2790) );
  NAND2_X1 U32810 ( .A1(REG2_REG_4__SCAN_IN), .A2(n5117), .ZN(n5115) );
  NAND2_X1 U32820 ( .A1(n3153), .A2(n2792), .ZN(n2793) );
  NAND2_X1 U32830 ( .A1(REG2_REG_6__SCAN_IN), .A2(n4260), .ZN(n4259) );
  NAND2_X1 U32840 ( .A1(n5074), .A2(n2795), .ZN(n2796) );
  NAND2_X1 U32850 ( .A1(n3373), .A2(n2798), .ZN(n2799) );
  NAND2_X1 U32860 ( .A1(n2799), .A2(n4290), .ZN(n3483) );
  NAND2_X1 U32870 ( .A1(n3482), .A2(n3483), .ZN(n3481) );
  NAND2_X1 U32880 ( .A1(n3463), .A2(n2801), .ZN(n2802) );
  INV_X1 U32890 ( .A(n3463), .ZN(n5231) );
  XNOR2_X1 U32900 ( .A(n2801), .B(n5231), .ZN(n4301) );
  NAND2_X1 U32910 ( .A1(n3547), .A2(n2804), .ZN(n2805) );
  NAND2_X1 U32920 ( .A1(REG2_REG_14__SCAN_IN), .A2(n4311), .ZN(n4310) );
  NOR2_X1 U32930 ( .A1(n3654), .A2(n2807), .ZN(n2808) );
  INV_X1 U32940 ( .A(n3654), .ZN(n5264) );
  OAI21_X1 U32950 ( .B1(n2809), .B2(IR_REG_16__SCAN_IN), .A(IR_REG_31__SCAN_IN), .ZN(n2810) );
  XNOR2_X1 U32960 ( .A(n2810), .B(IR_REG_17__SCAN_IN), .ZN(n5072) );
  OR2_X1 U32970 ( .A1(n5072), .A2(REG2_REG_17__SCAN_IN), .ZN(n4341) );
  XNOR2_X1 U32980 ( .A(n5071), .B(REG2_REG_18__SCAN_IN), .ZN(n4358) );
  INV_X1 U32990 ( .A(REG2_REG_19__SCAN_IN), .ZN(n2814) );
  NAND2_X1 U33000 ( .A1(n2812), .A2(n2811), .ZN(n2813) );
  MUX2_X1 U33010 ( .A(n2814), .B(REG2_REG_19__SCAN_IN), .S(n2961), .Z(n2815)
         );
  NOR2_X1 U33020 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2818) );
  NOR2_X1 U33030 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2817) );
  NAND4_X1 U33040 ( .A1(n2819), .A2(n2818), .A3(n2817), .A4(n2957), .ZN(n2820)
         );
  INV_X1 U33050 ( .A(n2825), .ZN(n2822) );
  INV_X1 U33060 ( .A(IR_REG_23__SCAN_IN), .ZN(n4799) );
  NAND2_X1 U33070 ( .A1(n2833), .A2(n4799), .ZN(n2823) );
  INV_X1 U33080 ( .A(IR_REG_24__SCAN_IN), .ZN(n4800) );
  NAND2_X1 U33090 ( .A1(n2825), .A2(n2828), .ZN(n2826) );
  NAND2_X1 U33100 ( .A1(n2826), .A2(IR_REG_31__SCAN_IN), .ZN(n2827) );
  INV_X1 U33110 ( .A(IR_REG_25__SCAN_IN), .ZN(n4801) );
  NOR2_X1 U33120 ( .A1(n2908), .A2(n3043), .ZN(n2832) );
  XNOR2_X1 U33130 ( .A(n2833), .B(n4799), .ZN(n3064) );
  NAND2_X1 U33140 ( .A1(n2958), .A2(n2900), .ZN(n3090) );
  INV_X1 U33150 ( .A(n3064), .ZN(n2834) );
  NAND2_X1 U33160 ( .A1(n2834), .A2(STATE_REG_SCAN_IN), .ZN(n3916) );
  AND2_X1 U33170 ( .A1(n3090), .A2(n3916), .ZN(n2888) );
  NAND2_X2 U33180 ( .A1(n2846), .A2(n2845), .ZN(n3107) );
  NAND2_X1 U33190 ( .A1(n2566), .A2(IR_REG_31__SCAN_IN), .ZN(n2842) );
  INV_X1 U33200 ( .A(IR_REG_22__SCAN_IN), .ZN(n4604) );
  XNOR2_X1 U33210 ( .A(n2842), .B(n4604), .ZN(n3075) );
  INV_X1 U33220 ( .A(n3075), .ZN(n4997) );
  NAND2_X1 U33230 ( .A1(n2916), .A2(IR_REG_31__SCAN_IN), .ZN(n2843) );
  NAND2_X1 U33240 ( .A1(n3082), .A2(n3064), .ZN(n2844) );
  NAND2_X1 U33250 ( .A1(n3794), .A2(n2844), .ZN(n2889) );
  OR2_X1 U33260 ( .A1(n2495), .A2(n2846), .ZN(n3911) );
  NOR2_X2 U33270 ( .A1(n5104), .A2(n3911), .ZN(n5116) );
  INV_X1 U33280 ( .A(n5116), .ZN(n2895) );
  INV_X1 U33290 ( .A(n5104), .ZN(n2887) );
  NAND2_X1 U33300 ( .A1(n2887), .A2(n2846), .ZN(n5108) );
  INV_X1 U33310 ( .A(REG1_REG_12__SCAN_IN), .ZN(n5236) );
  INV_X1 U33320 ( .A(REG1_REG_4__SCAN_IN), .ZN(n5170) );
  INV_X1 U33330 ( .A(n5113), .ZN(n5164) );
  INV_X1 U33340 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2847) );
  XNOR2_X1 U33350 ( .A(n2848), .B(n2847), .ZN(n2976) );
  INV_X1 U33360 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2849) );
  AND2_X1 U33370 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4238) );
  NAND2_X1 U33380 ( .A1(n2850), .A2(REG1_REG_1__SCAN_IN), .ZN(n2851) );
  NAND2_X1 U33390 ( .A1(n4237), .A2(n2851), .ZN(n2975) );
  NAND2_X1 U33400 ( .A1(n2976), .A2(n2975), .ZN(n2977) );
  NAND2_X1 U33410 ( .A1(n2848), .A2(REG1_REG_2__SCAN_IN), .ZN(n2852) );
  NAND2_X1 U33420 ( .A1(n2977), .A2(n2852), .ZN(n2853) );
  INV_X1 U33430 ( .A(REG1_REG_3__SCAN_IN), .ZN(n5160) );
  XNOR2_X1 U33440 ( .A(n5164), .B(n2855), .ZN(n5110) );
  NOR2_X1 U33450 ( .A1(n5170), .A2(n5110), .ZN(n5109) );
  NOR2_X1 U33460 ( .A1(n2855), .A2(n5164), .ZN(n2856) );
  NAND2_X1 U33470 ( .A1(n3145), .A2(REG1_REG_5__SCAN_IN), .ZN(n2857) );
  OAI21_X1 U33480 ( .B1(n3145), .B2(REG1_REG_5__SCAN_IN), .A(n2857), .ZN(n2931) );
  INV_X1 U33490 ( .A(REG1_REG_6__SCAN_IN), .ZN(n5187) );
  INV_X1 U33500 ( .A(n3153), .ZN(n5183) );
  NOR2_X1 U33510 ( .A1(n2859), .A2(n5183), .ZN(n2860) );
  INV_X1 U33520 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2861) );
  MUX2_X1 U3353 ( .A(n2861), .B(REG1_REG_7__SCAN_IN), .S(n3239), .Z(n2941) );
  INV_X1 U33540 ( .A(n2863), .ZN(n2864) );
  INV_X1 U3355 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2866) );
  MUX2_X1 U3356 ( .A(REG1_REG_9__SCAN_IN), .B(n2866), .S(n5206), .Z(n4281) );
  NOR2_X1 U3357 ( .A1(n2868), .A2(n2601), .ZN(n2869) );
  INV_X1 U3358 ( .A(REG1_REG_10__SCAN_IN), .ZN(n5218) );
  NAND2_X1 U3359 ( .A1(n3423), .A2(REG1_REG_11__SCAN_IN), .ZN(n2870) );
  OAI21_X1 U3360 ( .B1(n3423), .B2(REG1_REG_11__SCAN_IN), .A(n2870), .ZN(n3480) );
  INV_X1 U3361 ( .A(n3479), .ZN(n2871) );
  NOR2_X1 U3362 ( .A1(n2873), .A2(n5231), .ZN(n2874) );
  NAND2_X1 U3363 ( .A1(n3540), .A2(REG1_REG_13__SCAN_IN), .ZN(n2875) );
  OAI21_X1 U3364 ( .B1(n3540), .B2(REG1_REG_13__SCAN_IN), .A(n2875), .ZN(n3939) );
  INV_X1 U3365 ( .A(n3938), .ZN(n2876) );
  INV_X1 U3366 ( .A(REG1_REG_14__SCAN_IN), .ZN(n5252) );
  NOR2_X1 U3367 ( .A1(n2878), .A2(n2587), .ZN(n2879) );
  INV_X1 U3368 ( .A(REG1_REG_15__SCAN_IN), .ZN(n5260) );
  NOR2_X1 U3369 ( .A1(n5073), .A2(n5260), .ZN(n2880) );
  AOI21_X1 U3370 ( .B1(n5073), .B2(n5260), .A(n2880), .ZN(n4320) );
  INV_X1 U3371 ( .A(REG1_REG_16__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U3372 ( .A1(n4332), .A2(n5299), .ZN(n4331) );
  NAND2_X1 U3373 ( .A1(n2882), .A2(n5264), .ZN(n2883) );
  XNOR2_X1 U3374 ( .A(n5072), .B(REG1_REG_17__SCAN_IN), .ZN(n4350) );
  NAND2_X1 U3375 ( .A1(n5072), .A2(REG1_REG_17__SCAN_IN), .ZN(n2884) );
  INV_X1 U3376 ( .A(REG1_REG_18__SCAN_IN), .ZN(n2885) );
  XNOR2_X1 U3377 ( .A(n5071), .B(n2885), .ZN(n4364) );
  NAND2_X1 U3378 ( .A1(n4363), .A2(n4364), .ZN(n4361) );
  NAND2_X1 U3379 ( .A1(n5071), .A2(REG1_REG_18__SCAN_IN), .ZN(n2886) );
  NAND2_X1 U3380 ( .A1(n2887), .A2(n2495), .ZN(n4348) );
  INV_X1 U3381 ( .A(n2888), .ZN(n2890) );
  AND2_X1 U3382 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4162) );
  AOI21_X1 U3383 ( .B1(n5107), .B2(ADDR_REG_19__SCAN_IN), .A(n4162), .ZN(n2891) );
  OAI21_X1 U3384 ( .B1(n4348), .B2(n2961), .A(n2891), .ZN(n2892) );
  INV_X1 U3385 ( .A(n2892), .ZN(n2893) );
  OAI211_X1 U3386 ( .C1(n2510), .C2(n2895), .A(n2894), .B(n2893), .ZN(U3259)
         );
  INV_X1 U3387 ( .A(n2900), .ZN(n2911) );
  OR2_X2 U3388 ( .A1(n2958), .A2(n2911), .ZN(n4235) );
  INV_X1 U3389 ( .A(DATAI_21_), .ZN(n2896) );
  MUX2_X1 U3390 ( .A(n2896), .B(n3823), .S(STATE_REG_SCAN_IN), .Z(n2897) );
  INV_X1 U3391 ( .A(n2897), .ZN(U3331) );
  INV_X1 U3392 ( .A(DATAI_22_), .ZN(n2898) );
  MUX2_X1 U3393 ( .A(n3075), .B(n2898), .S(U3149), .Z(n2899) );
  INV_X1 U3394 ( .A(n2899), .ZN(U3330) );
  INV_X1 U3395 ( .A(DATAI_23_), .ZN(n2901) );
  AOI21_X1 U3396 ( .B1(n2901), .B2(U3149), .A(n2900), .ZN(U3329) );
  INV_X1 U3397 ( .A(DATAI_25_), .ZN(n2902) );
  MUX2_X1 U3398 ( .A(n2902), .B(n3043), .S(STATE_REG_SCAN_IN), .Z(n2903) );
  INV_X1 U3399 ( .A(n2903), .ZN(U3327) );
  INV_X1 U3400 ( .A(DATAI_27_), .ZN(n2904) );
  MUX2_X1 U3401 ( .A(n2904), .B(n2846), .S(STATE_REG_SCAN_IN), .Z(n2905) );
  INV_X1 U3402 ( .A(n2905), .ZN(U3325) );
  INV_X1 U3403 ( .A(DATAI_19_), .ZN(n2906) );
  MUX2_X1 U3404 ( .A(n2906), .B(n2961), .S(STATE_REG_SCAN_IN), .Z(n2907) );
  INV_X1 U3405 ( .A(n2907), .ZN(U3333) );
  INV_X1 U3406 ( .A(n3090), .ZN(n3052) );
  NAND2_X1 U3407 ( .A1(n3043), .A2(n2908), .ZN(n2909) );
  MUX2_X1 U3408 ( .A(n2908), .B(n2909), .S(B_REG_SCAN_IN), .Z(n2910) );
  NAND2_X1 U3409 ( .A1(n2910), .A2(n5069), .ZN(n3049) );
  NAND2_X1 U3410 ( .A1(n3052), .A2(n3049), .ZN(n5095) );
  INV_X1 U3411 ( .A(D_REG_1__SCAN_IN), .ZN(n2912) );
  NOR2_X1 U3412 ( .A1(n5069), .A2(n2911), .ZN(n4030) );
  AOI22_X1 U3413 ( .A1(n5095), .A2(n2912), .B1(n4030), .B2(n3043), .ZN(U3459)
         );
  NAND2_X1 U3414 ( .A1(n2914), .A2(n2918), .ZN(n2915) );
  INV_X1 U3415 ( .A(n2916), .ZN(n2919) );
  NAND2_X1 U3416 ( .A1(n2919), .A2(n2742), .ZN(n2921) );
  NAND2_X1 U3417 ( .A1(n3056), .A2(REG1_REG_30__SCAN_IN), .ZN(n2928) );
  NAND2_X1 U3418 ( .A1(n2494), .A2(REG2_REG_30__SCAN_IN), .ZN(n2927) );
  NAND2_X1 U3419 ( .A1(n3057), .A2(REG0_REG_30__SCAN_IN), .ZN(n2926) );
  AND3_X1 U3420 ( .A1(n2928), .A2(n2927), .A3(n2926), .ZN(n4414) );
  NAND2_X1 U3421 ( .A1(n4235), .A2(DATAO_REG_30__SCAN_IN), .ZN(n2929) );
  OAI21_X1 U3422 ( .B1(n4414), .B2(n4235), .A(n2929), .ZN(U3580) );
  NOR2_X1 U3423 ( .A1(n5107), .A2(U4043), .ZN(U3148) );
  AOI211_X1 U3424 ( .C1(n2932), .C2(n2931), .A(n2930), .B(n5108), .ZN(n2940)
         );
  OAI211_X1 U3425 ( .C1(n2935), .C2(n2934), .A(n5116), .B(n2933), .ZN(n2938)
         );
  INV_X1 U3426 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2936) );
  NOR2_X1 U3427 ( .A1(STATE_REG_SCAN_IN), .A2(n2936), .ZN(n3346) );
  AOI21_X1 U3428 ( .B1(n5107), .B2(ADDR_REG_5__SCAN_IN), .A(n3346), .ZN(n2937)
         );
  OAI211_X1 U3429 ( .C1(n4348), .C2(n5174), .A(n2938), .B(n2937), .ZN(n2939)
         );
  OR2_X1 U3430 ( .A1(n2940), .A2(n2939), .ZN(U3245) );
  AOI211_X1 U3431 ( .C1(n2942), .C2(n2941), .A(n2538), .B(n5108), .ZN(n2950)
         );
  OAI211_X1 U3432 ( .C1(n2945), .C2(n2944), .A(n5116), .B(n2943), .ZN(n2948)
         );
  INV_X1 U3433 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2946) );
  NOR2_X1 U3434 ( .A1(STATE_REG_SCAN_IN), .A2(n2946), .ZN(n4140) );
  AOI21_X1 U3435 ( .B1(n5107), .B2(ADDR_REG_7__SCAN_IN), .A(n4140), .ZN(n2947)
         );
  OAI211_X1 U3436 ( .C1(n4348), .C2(n5191), .A(n2948), .B(n2947), .ZN(n2949)
         );
  OR2_X1 U3437 ( .A1(n2950), .A2(n2949), .ZN(U3247) );
  OR2_X1 U3438 ( .A1(n2846), .A2(REG2_REG_0__SCAN_IN), .ZN(n2951) );
  INV_X1 U3439 ( .A(n2495), .ZN(n5068) );
  NAND2_X1 U3440 ( .A1(n2951), .A2(n5068), .ZN(n5100) );
  NAND2_X1 U3441 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4240) );
  OAI21_X1 U3442 ( .B1(n3911), .B2(n4240), .A(U4043), .ZN(n2974) );
  NAND2_X1 U3443 ( .A1(n3109), .A2(REG3_REG_0__SCAN_IN), .ZN(n2955) );
  NAND2_X1 U3444 ( .A1(n3057), .A2(REG0_REG_0__SCAN_IN), .ZN(n2954) );
  NAND2_X1 U3445 ( .A1(n2494), .A2(REG2_REG_0__SCAN_IN), .ZN(n2952) );
  NAND2_X1 U3446 ( .A1(n4236), .A2(n3492), .ZN(n2960) );
  NAND2_X1 U3447 ( .A1(n3079), .A2(n4050), .ZN(n2959) );
  NAND2_X1 U3448 ( .A1(n2960), .A2(n2959), .ZN(n3004) );
  INV_X1 U3449 ( .A(n2962), .ZN(n3188) );
  NAND2_X1 U3450 ( .A1(n3026), .A2(n4236), .ZN(n2964) );
  NAND2_X1 U3451 ( .A1(n3079), .A2(n3492), .ZN(n2963) );
  NAND2_X1 U3452 ( .A1(n2964), .A2(n2963), .ZN(n2967) );
  INV_X1 U3453 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2965) );
  AOI21_X1 U3454 ( .B1(n2572), .B2(n2965), .A(n2958), .ZN(n2966) );
  NOR3_X1 U3455 ( .A1(n3004), .A2(n2967), .A3(n2966), .ZN(n2971) );
  NAND2_X1 U3456 ( .A1(n2967), .A2(n3004), .ZN(n2970) );
  INV_X1 U3457 ( .A(n2958), .ZN(n2968) );
  NAND3_X1 U34580 ( .A1(n2968), .A2(IR_REG_0__SCAN_IN), .A3(
        REG1_REG_0__SCAN_IN), .ZN(n2969) );
  NAND2_X1 U34590 ( .A1(n2970), .A2(n2969), .ZN(n3003) );
  NOR2_X1 U3460 ( .A1(n2971), .A2(n3003), .ZN(n3235) );
  INV_X1 U3461 ( .A(n2846), .ZN(n2972) );
  NOR3_X1 U3462 ( .A1(n3235), .A2(n2972), .A3(n2495), .ZN(n2973) );
  AOI211_X1 U3463 ( .C1(n2572), .C2(n5100), .A(n2974), .B(n2973), .ZN(n5111)
         );
  INV_X1 U3464 ( .A(n2975), .ZN(n2980) );
  INV_X1 U3465 ( .A(n2976), .ZN(n2979) );
  AOI211_X1 U3466 ( .C1(n2980), .C2(n2979), .A(n2978), .B(n5108), .ZN(n2990)
         );
  AND3_X1 U34670 ( .A1(n2983), .A2(n4241), .A3(n2982), .ZN(n2984) );
  NOR3_X1 U3468 ( .A1(n2895), .A2(n2985), .A3(n2984), .ZN(n2989) );
  AOI22_X1 U34690 ( .A1(n5107), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n2986) );
  OAI21_X1 U3470 ( .B1(n2987), .B2(n4348), .A(n2986), .ZN(n2988) );
  OR4_X1 U34710 ( .A1(n5111), .A2(n2990), .A3(n2989), .A4(n2988), .ZN(U3242)
         );
  INV_X1 U3472 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3068) );
  NAND2_X1 U34730 ( .A1(n3109), .A2(n3068), .ZN(n2994) );
  NAND2_X1 U3474 ( .A1(n3057), .A2(REG0_REG_3__SCAN_IN), .ZN(n2993) );
  NAND2_X1 U34750 ( .A1(n3056), .A2(REG1_REG_3__SCAN_IN), .ZN(n2992) );
  NAND2_X1 U3476 ( .A1(n2494), .A2(REG2_REG_3__SCAN_IN), .ZN(n2991) );
  NAND2_X1 U34770 ( .A1(n4234), .A2(n3492), .ZN(n2996) );
  MUX2_X1 U3478 ( .A(n4248), .B(DATAI_3_), .S(n3107), .Z(n3208) );
  NAND2_X1 U34790 ( .A1(n3208), .A2(n4050), .ZN(n2995) );
  NAND2_X1 U3480 ( .A1(n2996), .A2(n2995), .ZN(n3001) );
  XNOR2_X1 U34810 ( .A(n3001), .B(n3024), .ZN(n3268) );
  AND2_X1 U3482 ( .A1(n3208), .A2(n3492), .ZN(n3002) );
  AOI21_X1 U34830 ( .B1(n4234), .B2(n3026), .A(n3002), .ZN(n3269) );
  XNOR2_X1 U3484 ( .A(n3268), .B(n3269), .ZN(n3273) );
  INV_X1 U34850 ( .A(n3003), .ZN(n3005) );
  NAND2_X1 U3486 ( .A1(n3005), .A2(n2744), .ZN(n4020) );
  NAND2_X1 U34870 ( .A1(n3056), .A2(REG1_REG_1__SCAN_IN), .ZN(n3009) );
  NAND2_X1 U3488 ( .A1(n3109), .A2(REG3_REG_1__SCAN_IN), .ZN(n3008) );
  NAND2_X1 U34890 ( .A1(n2493), .A2(REG0_REG_1__SCAN_IN), .ZN(n3007) );
  NAND2_X1 U3490 ( .A1(n3240), .A2(REG2_REG_1__SCAN_IN), .ZN(n3006) );
  NAND4_X1 U34910 ( .A1(n3009), .A2(n3008), .A3(n3007), .A4(n3006), .ZN(n3078)
         );
  NAND2_X1 U3492 ( .A1(n3078), .A2(n3492), .ZN(n3011) );
  NAND2_X1 U34930 ( .A1(n3116), .A2(n4050), .ZN(n3010) );
  NAND2_X1 U3494 ( .A1(n3011), .A2(n3010), .ZN(n3012) );
  XNOR2_X1 U34950 ( .A(n3012), .B(n3024), .ZN(n3016) );
  AND2_X1 U3496 ( .A1(n3116), .A2(n3492), .ZN(n3013) );
  AOI21_X1 U34970 ( .B1(n3078), .B2(n3026), .A(n3013), .ZN(n3014) );
  XNOR2_X1 U3498 ( .A(n3016), .B(n3014), .ZN(n4022) );
  NAND2_X1 U34990 ( .A1(n4020), .A2(n4022), .ZN(n4021) );
  INV_X1 U3500 ( .A(n3014), .ZN(n3015) );
  NAND2_X1 U35010 ( .A1(n3016), .A2(n3015), .ZN(n3017) );
  NAND2_X1 U3502 ( .A1(n4021), .A2(n3017), .ZN(n3193) );
  INV_X1 U35030 ( .A(n3193), .ZN(n3029) );
  NAND2_X1 U3504 ( .A1(n3057), .A2(REG0_REG_2__SCAN_IN), .ZN(n3021) );
  NAND2_X1 U35050 ( .A1(n3056), .A2(REG1_REG_2__SCAN_IN), .ZN(n3020) );
  NAND2_X1 U35060 ( .A1(n3109), .A2(REG3_REG_2__SCAN_IN), .ZN(n3019) );
  NAND2_X1 U35070 ( .A1(n2494), .A2(REG2_REG_2__SCAN_IN), .ZN(n3018) );
  NAND4_X1 U35080 ( .A1(n3021), .A2(n3020), .A3(n3019), .A4(n3018), .ZN(n3105)
         );
  NAND2_X1 U35090 ( .A1(n3105), .A2(n3492), .ZN(n3023) );
  NAND2_X1 U35100 ( .A1(n3187), .A2(n4050), .ZN(n3022) );
  NAND2_X1 U35110 ( .A1(n3023), .A2(n3022), .ZN(n3025) );
  XNOR2_X1 U35120 ( .A(n3025), .B(n3490), .ZN(n3031) );
  AND2_X1 U35130 ( .A1(n3187), .A2(n3492), .ZN(n3027) );
  AOI21_X1 U35140 ( .B1(n3105), .B2(n3026), .A(n3027), .ZN(n3030) );
  XNOR2_X1 U35150 ( .A(n3031), .B(n3030), .ZN(n3194) );
  NAND2_X1 U35160 ( .A1(n3029), .A2(n3028), .ZN(n3310) );
  NAND2_X1 U35170 ( .A1(n3031), .A2(n3030), .ZN(n3271) );
  NAND2_X1 U35180 ( .A1(n3310), .A2(n3271), .ZN(n3032) );
  XOR2_X1 U35190 ( .A(n3273), .B(n3032), .Z(n3074) );
  NOR4_X1 U35200 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n3033) );
  INV_X1 U35210 ( .A(D_REG_16__SCAN_IN), .ZN(n5086) );
  INV_X1 U35220 ( .A(D_REG_17__SCAN_IN), .ZN(n5087) );
  NAND3_X1 U35230 ( .A1(n3033), .A2(n5086), .A3(n5087), .ZN(n3039) );
  NOR4_X1 U35240 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_23__SCAN_IN), .ZN(n3037) );
  NOR4_X1 U35250 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n3036) );
  NOR4_X1 U35260 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_7__SCAN_IN), .ZN(n3035) );
  NOR4_X1 U35270 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n3034) );
  NAND4_X1 U35280 ( .A1(n3037), .A2(n3036), .A3(n3035), .A4(n3034), .ZN(n3038)
         );
  NOR4_X1 U35290 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(n3039), 
        .A4(n3038), .ZN(n3042) );
  INV_X1 U35300 ( .A(D_REG_6__SCAN_IN), .ZN(n5078) );
  INV_X1 U35310 ( .A(D_REG_5__SCAN_IN), .ZN(n5077) );
  INV_X1 U35320 ( .A(D_REG_12__SCAN_IN), .ZN(n5083) );
  INV_X1 U35330 ( .A(D_REG_8__SCAN_IN), .ZN(n5079) );
  NAND4_X1 U35340 ( .A1(n5078), .A2(n5077), .A3(n5083), .A4(n5079), .ZN(n3040)
         );
  NOR3_X1 U35350 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(n3040), 
        .ZN(n3041) );
  AND2_X1 U35360 ( .A1(n3042), .A2(n3041), .ZN(n3088) );
  INV_X1 U35370 ( .A(n3043), .ZN(n3044) );
  OAI22_X1 U35380 ( .A1(n3049), .A2(D_REG_1__SCAN_IN), .B1(n5069), .B2(n3044), 
        .ZN(n5006) );
  INV_X1 U35390 ( .A(n5006), .ZN(n3093) );
  INV_X1 U35400 ( .A(n3049), .ZN(n3045) );
  INV_X1 U35410 ( .A(D_REG_0__SCAN_IN), .ZN(n4622) );
  NAND2_X1 U35420 ( .A1(n3045), .A2(n4622), .ZN(n3048) );
  INV_X1 U35430 ( .A(n5069), .ZN(n3046) );
  NAND2_X1 U35440 ( .A1(n3046), .A2(n2908), .ZN(n3047) );
  OAI211_X1 U35450 ( .C1(n3088), .C2(n3049), .A(n3093), .B(n5009), .ZN(n3062)
         );
  INV_X1 U35460 ( .A(n3062), .ZN(n3053) );
  NAND2_X1 U35470 ( .A1(n3053), .A2(n3052), .ZN(n3195) );
  INV_X1 U35480 ( .A(n3082), .ZN(n3083) );
  INV_X1 U35490 ( .A(n2997), .ZN(n3907) );
  NAND3_X1 U35500 ( .A1(n5005), .A2(n3083), .A3(n5315), .ZN(n3050) );
  OR2_X2 U35510 ( .A1(n3195), .A2(n3050), .ZN(n5271) );
  NAND2_X1 U35520 ( .A1(n2997), .A2(n2961), .ZN(n3063) );
  INV_X1 U35530 ( .A(n3063), .ZN(n3051) );
  AND3_X1 U35540 ( .A1(n3052), .A2(n3051), .A3(n3082), .ZN(n3913) );
  INV_X1 U35550 ( .A(n3069), .ZN(n3054) );
  NAND2_X1 U35560 ( .A1(n2494), .A2(REG2_REG_4__SCAN_IN), .ZN(n3061) );
  NOR2_X1 U35570 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n3055) );
  NOR2_X1 U35580 ( .A1(n3110), .A2(n3055), .ZN(n3277) );
  NAND2_X1 U35590 ( .A1(n3109), .A2(n3277), .ZN(n3060) );
  NAND2_X1 U35600 ( .A1(n3057), .A2(REG0_REG_4__SCAN_IN), .ZN(n3058) );
  NAND2_X1 U35610 ( .A1(n3062), .A2(n5005), .ZN(n3066) );
  NAND2_X1 U35620 ( .A1(n3063), .A2(n3082), .ZN(n3196) );
  AND3_X1 U35630 ( .A1(n3196), .A2(n2958), .A3(n3064), .ZN(n3065) );
  NAND2_X1 U35640 ( .A1(n3066), .A2(n3065), .ZN(n3067) );
  NAND2_X1 U35650 ( .A1(n3067), .A2(STATE_REG_SCAN_IN), .ZN(n5280) );
  AOI22_X1 U35660 ( .A1(n4219), .A2(n3108), .B1(n4183), .B2(n3068), .ZN(n3073)
         );
  NOR2_X1 U35670 ( .A1(STATE_REG_SCAN_IN), .A2(n3068), .ZN(n4250) );
  OR2_X1 U35680 ( .A1(n3195), .A2(n5315), .ZN(n3070) );
  NAND2_X1 U35690 ( .A1(n3070), .A2(n4991), .ZN(n5266) );
  NOR2_X1 U35700 ( .A1(n4214), .A2(n3215), .ZN(n3071) );
  AOI211_X1 U35710 ( .C1(n5268), .C2(n3105), .A(n4250), .B(n3071), .ZN(n3072)
         );
  OAI211_X1 U35720 ( .C1(n3074), .C2(n5271), .A(n3073), .B(n3072), .ZN(U3215)
         );
  OR2_X1 U35730 ( .A1(n2997), .A2(n3823), .ZN(n3077) );
  OR2_X1 U35740 ( .A1(n2961), .A2(n3075), .ZN(n3076) );
  NAND2_X1 U35750 ( .A1(n3078), .A2(n4029), .ZN(n3856) );
  INV_X1 U35760 ( .A(n3078), .ZN(n3199) );
  NAND2_X1 U35770 ( .A1(n3199), .A2(n3116), .ZN(n3859) );
  INV_X1 U35780 ( .A(n4236), .ZN(n4023) );
  NAND2_X1 U35790 ( .A1(n4023), .A2(n3079), .ZN(n3855) );
  NAND2_X1 U35800 ( .A1(n3080), .A2(n3081), .ZN(n3118) );
  AND2_X1 U35810 ( .A1(n2495), .A2(n3082), .ZN(n5286) );
  AOI22_X1 U3582 ( .A1(n3105), .A2(n5286), .B1(n5325), .B2(n3116), .ZN(n3085)
         );
  NOR2_X2 U3583 ( .A1(n2495), .A2(n3083), .ZN(n4957) );
  NAND2_X1 U3584 ( .A1(n4236), .A2(n4957), .ZN(n3084) );
  OAI211_X1 U3585 ( .C1(n5140), .C2(n4999), .A(n3085), .B(n3084), .ZN(n3086)
         );
  AOI21_X1 U3586 ( .B1(n5124), .B2(n3087), .A(n3086), .ZN(n5141) );
  INV_X1 U3587 ( .A(n3088), .ZN(n3089) );
  OR2_X1 U3588 ( .A1(n3090), .A2(n3089), .ZN(n3091) );
  NAND2_X1 U3589 ( .A1(n5095), .A2(n3091), .ZN(n3092) );
  NAND2_X1 U3590 ( .A1(n3092), .A2(n3196), .ZN(n5008) );
  INV_X1 U3591 ( .A(n5008), .ZN(n3094) );
  NAND3_X1 U3592 ( .A1(n3094), .A2(n3093), .A3(n5049), .ZN(n3095) );
  NOR2_X1 U3593 ( .A1(n5336), .A2(n5130), .ZN(n4390) );
  NAND2_X1 U3594 ( .A1(n3116), .A2(n3079), .ZN(n3096) );
  INV_X1 U3595 ( .A(n5296), .ZN(n5339) );
  NAND2_X1 U3596 ( .A1(n3096), .A2(n5339), .ZN(n3097) );
  NOR2_X1 U3597 ( .A1(n3185), .A2(n3097), .ZN(n5143) );
  INV_X1 U3598 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3098) );
  OAI22_X1 U3599 ( .A1(n5138), .A2(n2784), .B1(n3098), .B2(n4991), .ZN(n3102)
         );
  NAND2_X1 U3600 ( .A1(n3099), .A2(n5130), .ZN(n3154) );
  INV_X1 U3601 ( .A(n3154), .ZN(n3100) );
  AND2_X1 U3602 ( .A1(n5138), .A2(n3100), .ZN(n5134) );
  INV_X1 U3603 ( .A(n5134), .ZN(n3191) );
  NOR2_X1 U3604 ( .A1(n5140), .A2(n3191), .ZN(n3101) );
  AOI211_X1 U3605 ( .C1(n4390), .C2(n5143), .A(n3102), .B(n3101), .ZN(n3103)
         );
  OAI21_X1 U3606 ( .B1(n5141), .B2(n5336), .A(n3103), .ZN(U3289) );
  NAND2_X1 U3607 ( .A1(n3104), .A2(n3859), .ZN(n3179) );
  INV_X1 U3608 ( .A(n3105), .ZN(n4024) );
  NAND2_X1 U3609 ( .A1(n4024), .A2(n3187), .ZN(n3860) );
  NAND2_X1 U3610 ( .A1(n3105), .A2(n3198), .ZN(n3863) );
  INV_X1 U3611 ( .A(n4234), .ZN(n3200) );
  NAND2_X1 U3612 ( .A1(n3200), .A2(n3208), .ZN(n3865) );
  NAND2_X1 U3613 ( .A1(n4234), .A2(n3215), .ZN(n3862) );
  AND2_X1 U3614 ( .A1(n3865), .A2(n3862), .ZN(n3842) );
  NAND2_X1 U3615 ( .A1(n3207), .A2(n3842), .ZN(n3106) );
  XNOR2_X1 U3616 ( .A(n3157), .B(n3138), .ZN(n3127) );
  NAND2_X1 U3617 ( .A1(n3057), .A2(REG0_REG_5__SCAN_IN), .ZN(n3115) );
  OAI21_X1 U3618 ( .B1(n3110), .B2(REG3_REG_5__SCAN_IN), .A(n3161), .ZN(n3111)
         );
  INV_X1 U3619 ( .A(n3111), .ZN(n3345) );
  NAND2_X1 U3620 ( .A1(n3109), .A2(n3345), .ZN(n3114) );
  NAND2_X1 U3621 ( .A1(n3056), .A2(REG1_REG_5__SCAN_IN), .ZN(n3113) );
  NAND2_X1 U3622 ( .A1(n2494), .A2(REG2_REG_5__SCAN_IN), .ZN(n3112) );
  NAND4_X1 U3623 ( .A1(n3115), .A2(n3114), .A3(n3113), .A4(n3112), .ZN(n4233)
         );
  INV_X1 U3624 ( .A(n4233), .ZN(n3167) );
  NAND2_X1 U3625 ( .A1(n3078), .A2(n3116), .ZN(n3117) );
  INV_X1 U3626 ( .A(n3178), .ZN(n3120) );
  INV_X1 U3627 ( .A(n3837), .ZN(n3119) );
  NAND2_X1 U3628 ( .A1(n3200), .A2(n3215), .ZN(n3121) );
  NAND2_X1 U3629 ( .A1(n3137), .A2(n3135), .ZN(n3122) );
  NAND2_X1 U3630 ( .A1(n4234), .A2(n3208), .ZN(n3139) );
  AND2_X1 U3631 ( .A1(n3122), .A2(n3139), .ZN(n3123) );
  AOI21_X1 U3632 ( .B1(n3138), .B2(n3123), .A(n2740), .ZN(n5169) );
  INV_X1 U3633 ( .A(n4999), .ZN(n5125) );
  NAND2_X1 U3634 ( .A1(n5169), .A2(n5125), .ZN(n3125) );
  AOI22_X1 U3635 ( .A1(n4234), .A2(n4957), .B1(n3266), .B2(n5325), .ZN(n3124)
         );
  OAI211_X1 U3636 ( .C1(n3167), .C2(n5127), .A(n3125), .B(n3124), .ZN(n3126)
         );
  AOI21_X1 U3637 ( .B1(n3127), .B2(n5124), .A(n3126), .ZN(n5165) );
  NAND2_X1 U3638 ( .A1(n3216), .A2(n3215), .ZN(n3214) );
  AOI21_X1 U3639 ( .B1(n3214), .B2(n3266), .A(n5296), .ZN(n3128) );
  AND2_X1 U3640 ( .A1(n3128), .A2(n3229), .ZN(n5167) );
  INV_X1 U3641 ( .A(REG2_REG_4__SCAN_IN), .ZN(n3130) );
  INV_X1 U3642 ( .A(n3277), .ZN(n3129) );
  OAI22_X1 U3643 ( .A1(n5138), .A2(n3130), .B1(n3129), .B2(n4991), .ZN(n3131)
         );
  AOI21_X1 U3644 ( .B1(n5167), .B2(n4390), .A(n3131), .ZN(n3133) );
  NAND2_X1 U3645 ( .A1(n5169), .A2(n5134), .ZN(n3132) );
  OAI211_X1 U3646 ( .C1(n5165), .C2(n5333), .A(n3133), .B(n3132), .ZN(U3286)
         );
  AND2_X1 U3647 ( .A1(n3135), .A2(n3134), .ZN(n3136) );
  NAND2_X1 U3648 ( .A1(n3137), .A2(n3136), .ZN(n3144) );
  INV_X1 U3649 ( .A(n3139), .ZN(n3140) );
  NAND2_X1 U3650 ( .A1(n3134), .A2(n3140), .ZN(n3142) );
  NAND2_X1 U3651 ( .A1(n3108), .A2(n3266), .ZN(n3141) );
  AND2_X1 U3652 ( .A1(n3142), .A2(n3141), .ZN(n3143) );
  MUX2_X1 U3653 ( .A(n3145), .B(DATAI_5_), .S(n3794), .Z(n3325) );
  INV_X1 U3654 ( .A(n3325), .ZN(n3349) );
  NAND2_X1 U3655 ( .A1(n3167), .A2(n3349), .ZN(n3146) );
  NAND2_X1 U3656 ( .A1(n3228), .A2(n3146), .ZN(n3148) );
  NAND2_X1 U3657 ( .A1(n4233), .A2(n3325), .ZN(n3147) );
  NAND2_X1 U3658 ( .A1(n2494), .A2(REG2_REG_6__SCAN_IN), .ZN(n3152) );
  XNOR2_X1 U3659 ( .A(n3161), .B(REG3_REG_6__SCAN_IN), .ZN(n3336) );
  NAND2_X1 U3660 ( .A1(n3109), .A2(n3336), .ZN(n3151) );
  NAND2_X1 U3661 ( .A1(n3056), .A2(REG1_REG_6__SCAN_IN), .ZN(n3150) );
  NAND2_X1 U3662 ( .A1(n3057), .A2(REG0_REG_6__SCAN_IN), .ZN(n3149) );
  NAND4_X1 U3663 ( .A1(n3152), .A2(n3151), .A3(n3150), .A4(n3149), .ZN(n4232)
         );
  INV_X1 U3664 ( .A(n4232), .ZN(n3227) );
  MUX2_X1 U3665 ( .A(n3153), .B(DATAI_6_), .S(n3794), .Z(n3334) );
  NAND2_X1 U3666 ( .A1(n3227), .A2(n3334), .ZN(n3872) );
  INV_X1 U3667 ( .A(n3334), .ZN(n3337) );
  NAND2_X1 U3668 ( .A1(n4232), .A2(n3337), .ZN(n3874) );
  XNOR2_X1 U3669 ( .A(n3257), .B(n3840), .ZN(n5186) );
  INV_X1 U3670 ( .A(n5186), .ZN(n3176) );
  NAND2_X1 U3671 ( .A1(n4999), .A2(n3154), .ZN(n3155) );
  INV_X1 U3672 ( .A(n3866), .ZN(n3156) );
  NAND2_X1 U3673 ( .A1(n3167), .A2(n3325), .ZN(n3871) );
  NAND2_X1 U3674 ( .A1(n4233), .A2(n3349), .ZN(n3868) );
  AND2_X1 U3675 ( .A1(n3871), .A2(n3868), .ZN(n3841) );
  NAND2_X1 U3676 ( .A1(n3158), .A2(n3868), .ZN(n3238) );
  XNOR2_X1 U3677 ( .A(n3238), .B(n3840), .ZN(n3170) );
  NAND2_X1 U3678 ( .A1(n2494), .A2(REG2_REG_7__SCAN_IN), .ZN(n3166) );
  INV_X1 U3679 ( .A(n3161), .ZN(n3159) );
  AOI21_X1 U3680 ( .B1(n3159), .B2(REG3_REG_6__SCAN_IN), .A(
        REG3_REG_7__SCAN_IN), .ZN(n3162) );
  NAND2_X1 U3681 ( .A1(REG3_REG_7__SCAN_IN), .A2(REG3_REG_6__SCAN_IN), .ZN(
        n3160) );
  OR2_X1 U3682 ( .A1(n3162), .A2(n3241), .ZN(n3252) );
  INV_X1 U3683 ( .A(n3252), .ZN(n4137) );
  NAND2_X1 U3684 ( .A1(n3109), .A2(n4137), .ZN(n3165) );
  NAND2_X1 U3685 ( .A1(n3056), .A2(REG1_REG_7__SCAN_IN), .ZN(n3164) );
  NAND2_X1 U3686 ( .A1(n3057), .A2(REG0_REG_7__SCAN_IN), .ZN(n3163) );
  NAND4_X1 U3687 ( .A1(n3166), .A2(n3165), .A3(n3164), .A4(n3163), .ZN(n4231)
         );
  OAI22_X1 U3688 ( .A1(n3167), .A2(n5282), .B1(n5315), .B2(n3337), .ZN(n3168)
         );
  AOI21_X1 U3689 ( .B1(n5286), .B2(n4231), .A(n3168), .ZN(n3169) );
  OAI21_X1 U3690 ( .B1(n3170), .B2(n5288), .A(n3169), .ZN(n5184) );
  NAND2_X1 U3691 ( .A1(n5184), .A2(n5138), .ZN(n3175) );
  AOI211_X1 U3692 ( .C1(n3334), .C2(n3230), .A(n5296), .B(n3251), .ZN(n5185)
         );
  INV_X1 U3693 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3172) );
  INV_X1 U3694 ( .A(n3336), .ZN(n3171) );
  OAI22_X1 U3695 ( .A1(n5138), .A2(n3172), .B1(n3171), .B2(n4991), .ZN(n3173)
         );
  AOI21_X1 U3696 ( .B1(n5185), .B2(n4390), .A(n3173), .ZN(n3174) );
  OAI211_X1 U3697 ( .C1(n3176), .C2(n5307), .A(n3175), .B(n3174), .ZN(U3284)
         );
  INV_X1 U3698 ( .A(n3137), .ZN(n3177) );
  AOI21_X1 U3699 ( .B1(n3837), .B2(n3178), .A(n3177), .ZN(n5147) );
  AOI22_X1 U3700 ( .A1(n3078), .A2(n4957), .B1(n3187), .B2(n5325), .ZN(n3180)
         );
  OAI21_X1 U3701 ( .B1(n3200), .B2(n5127), .A(n3180), .ZN(n3182) );
  NOR2_X1 U3702 ( .A1(n5147), .A2(n4999), .ZN(n3181) );
  AOI211_X1 U3703 ( .C1(n5124), .C2(n3183), .A(n3182), .B(n3181), .ZN(n5148)
         );
  MUX2_X1 U3704 ( .A(n3184), .B(n5148), .S(n5138), .Z(n3190) );
  INV_X1 U3705 ( .A(n3185), .ZN(n3186) );
  AOI21_X1 U3706 ( .B1(n3187), .B2(n3186), .A(n3216), .ZN(n5151) );
  NAND2_X1 U3707 ( .A1(n5138), .A2(n2962), .ZN(n5306) );
  INV_X1 U3708 ( .A(n5306), .ZN(n5334) );
  AOI22_X1 U3709 ( .A1(n5151), .A2(n5334), .B1(REG3_REG_2__SCAN_IN), .B2(n5303), .ZN(n3189) );
  OAI211_X1 U3710 ( .C1(n5147), .C2(n3191), .A(n3190), .B(n3189), .ZN(U3288)
         );
  INV_X1 U3711 ( .A(n3310), .ZN(n3192) );
  AOI21_X1 U3712 ( .B1(n3194), .B2(n3193), .A(n3192), .ZN(n3204) );
  INV_X1 U3713 ( .A(n3195), .ZN(n3197) );
  OAI21_X1 U3714 ( .B1(n3197), .B2(n5303), .A(n3196), .ZN(n4026) );
  NOR2_X1 U3715 ( .A1(n4214), .A2(n3198), .ZN(n3202) );
  INV_X1 U3716 ( .A(n4219), .ZN(n4205) );
  OAI22_X1 U3717 ( .A1(n3200), .A2(n4205), .B1(n4216), .B2(n3199), .ZN(n3201)
         );
  AOI211_X1 U3718 ( .C1(REG3_REG_2__SCAN_IN), .C2(n4026), .A(n3202), .B(n3201), 
        .ZN(n3203) );
  OAI21_X1 U3719 ( .B1(n3204), .B2(n5271), .A(n3203), .ZN(U3234) );
  NAND2_X1 U3720 ( .A1(n3137), .A2(n3205), .ZN(n3206) );
  XNOR2_X1 U3721 ( .A(n3206), .B(n3842), .ZN(n5157) );
  XNOR2_X1 U3722 ( .A(n3207), .B(n3842), .ZN(n3212) );
  AOI22_X1 U3723 ( .A1(n3105), .A2(n4957), .B1(n5325), .B2(n3208), .ZN(n3209)
         );
  OAI21_X1 U3724 ( .B1(n3210), .B2(n5127), .A(n3209), .ZN(n3211) );
  AOI21_X1 U3725 ( .B1(n3212), .B2(n5124), .A(n3211), .ZN(n3213) );
  OAI21_X1 U3726 ( .B1(n5157), .B2(n4999), .A(n3213), .ZN(n5159) );
  INV_X1 U3727 ( .A(n5159), .ZN(n3221) );
  INV_X1 U3728 ( .A(n5157), .ZN(n3219) );
  OAI21_X1 U3729 ( .B1(n3216), .B2(n3215), .A(n3214), .ZN(n5155) );
  AOI22_X1 U3730 ( .A1(n5333), .A2(REG2_REG_3__SCAN_IN), .B1(n5303), .B2(n3068), .ZN(n3217) );
  OAI21_X1 U3731 ( .B1(n5155), .B2(n5306), .A(n3217), .ZN(n3218) );
  AOI21_X1 U3732 ( .B1(n3219), .B2(n5134), .A(n3218), .ZN(n3220) );
  OAI21_X1 U3733 ( .B1(n3221), .B2(n5336), .A(n3220), .ZN(U3287) );
  INV_X1 U3734 ( .A(n3841), .ZN(n3222) );
  XNOR2_X1 U3735 ( .A(n3223), .B(n3222), .ZN(n3224) );
  NAND2_X1 U3736 ( .A1(n3224), .A2(n5124), .ZN(n3226) );
  AOI22_X1 U3737 ( .A1(n3108), .A2(n4957), .B1(n3325), .B2(n5325), .ZN(n3225)
         );
  OAI211_X1 U3738 ( .C1(n3227), .C2(n5127), .A(n3226), .B(n3225), .ZN(n5176)
         );
  INV_X1 U3739 ( .A(n5176), .ZN(n3234) );
  XNOR2_X1 U3740 ( .A(n3228), .B(n3841), .ZN(n5178) );
  INV_X1 U3741 ( .A(n5307), .ZN(n4986) );
  OAI21_X1 U3742 ( .B1(n2575), .B2(n3349), .A(n3230), .ZN(n5175) );
  AOI22_X1 U3743 ( .A1(n5333), .A2(REG2_REG_5__SCAN_IN), .B1(n3345), .B2(n5303), .ZN(n3231) );
  OAI21_X1 U3744 ( .B1(n5175), .B2(n5306), .A(n3231), .ZN(n3232) );
  AOI21_X1 U3745 ( .B1(n5178), .B2(n4986), .A(n3232), .ZN(n3233) );
  OAI21_X1 U3746 ( .B1(n3234), .B2(n5336), .A(n3233), .ZN(U3285) );
  INV_X1 U3747 ( .A(n5271), .ZN(n4134) );
  AOI22_X1 U3748 ( .A1(n3235), .A2(n4134), .B1(n5276), .B2(n3078), .ZN(n3237)
         );
  AOI22_X1 U3749 ( .A1(n4026), .A2(REG3_REG_0__SCAN_IN), .B1(n3079), .B2(n5266), .ZN(n3236) );
  NAND2_X1 U3750 ( .A1(n3237), .A2(n3236), .ZN(U3229) );
  MUX2_X1 U3751 ( .A(n3239), .B(DATAI_7_), .S(n3794), .Z(n3408) );
  XNOR2_X1 U3752 ( .A(n4231), .B(n3408), .ZN(n3816) );
  INV_X1 U3753 ( .A(n3816), .ZN(n3258) );
  XNOR2_X1 U3754 ( .A(n3301), .B(n3258), .ZN(n3250) );
  NAND2_X1 U3755 ( .A1(n2494), .A2(REG2_REG_8__SCAN_IN), .ZN(n3246) );
  OR2_X1 U3756 ( .A1(n3241), .A2(REG3_REG_8__SCAN_IN), .ZN(n3242) );
  AND2_X1 U3757 ( .A1(n3295), .A2(n3242), .ZN(n3417) );
  NAND2_X1 U3758 ( .A1(n3109), .A2(n3417), .ZN(n3245) );
  NAND2_X1 U3759 ( .A1(n3056), .A2(REG1_REG_8__SCAN_IN), .ZN(n3244) );
  NAND2_X1 U3760 ( .A1(n3057), .A2(REG0_REG_8__SCAN_IN), .ZN(n3243) );
  NAND4_X1 U3761 ( .A1(n3246), .A2(n3245), .A3(n3244), .A4(n3243), .ZN(n4230)
         );
  NAND2_X1 U3762 ( .A1(n4230), .A2(n5286), .ZN(n3248) );
  NAND2_X1 U3763 ( .A1(n4232), .A2(n4957), .ZN(n3247) );
  OAI211_X1 U3764 ( .C1(n5315), .C2(n4138), .A(n3248), .B(n3247), .ZN(n3249)
         );
  AOI21_X1 U3765 ( .B1(n3250), .B2(n5124), .A(n3249), .ZN(n5195) );
  OAI211_X1 U3766 ( .C1(n3251), .C2(n4138), .A(n5339), .B(n3289), .ZN(n5194)
         );
  INV_X1 U3767 ( .A(n5194), .ZN(n3255) );
  OAI22_X1 U3768 ( .A1(n5138), .A2(n3253), .B1(n3252), .B2(n4991), .ZN(n3254)
         );
  AOI21_X1 U3769 ( .B1(n3255), .B2(n4390), .A(n3254), .ZN(n3262) );
  AND2_X1 U3770 ( .A1(n4232), .A2(n3334), .ZN(n3256) );
  INV_X1 U3771 ( .A(n3260), .ZN(n3259) );
  NAND2_X1 U3772 ( .A1(n3259), .A2(n3258), .ZN(n3285) );
  NAND2_X1 U3773 ( .A1(n3260), .A2(n3816), .ZN(n5192) );
  NAND3_X1 U3774 ( .A1(n3285), .A2(n5192), .A3(n4986), .ZN(n3261) );
  OAI211_X1 U3775 ( .C1(n5195), .C2(n5333), .A(n3262), .B(n3261), .ZN(U3283)
         );
  NAND2_X1 U3776 ( .A1(n3108), .A2(n3492), .ZN(n3264) );
  NAND2_X1 U3777 ( .A1(n3266), .A2(n4050), .ZN(n3263) );
  NAND2_X1 U3778 ( .A1(n3264), .A2(n3263), .ZN(n3265) );
  XNOR2_X1 U3779 ( .A(n3265), .B(n3490), .ZN(n3311) );
  AND2_X1 U3780 ( .A1(n3266), .A2(n3492), .ZN(n3267) );
  XNOR2_X1 U3781 ( .A(n3311), .B(n3312), .ZN(n3316) );
  INV_X1 U3782 ( .A(n3268), .ZN(n3270) );
  NAND2_X1 U3783 ( .A1(n3270), .A2(n3269), .ZN(n3272) );
  AND2_X1 U3784 ( .A1(n3271), .A2(n3272), .ZN(n3307) );
  NAND2_X1 U3785 ( .A1(n3310), .A2(n3307), .ZN(n3275) );
  INV_X1 U3786 ( .A(n3272), .ZN(n3274) );
  OR2_X1 U3787 ( .A1(n3274), .A2(n3273), .ZN(n3317) );
  AND2_X1 U3788 ( .A1(n3275), .A2(n3317), .ZN(n3276) );
  AOI211_X1 U3789 ( .C1(n3316), .C2(n3276), .A(n5271), .B(n2534), .ZN(n3283)
         );
  AOI22_X1 U3790 ( .A1(n5276), .A2(n4233), .B1(n4183), .B2(n3277), .ZN(n3280)
         );
  INV_X1 U3791 ( .A(REG3_REG_4__SCAN_IN), .ZN(n3278) );
  NOR2_X1 U3792 ( .A1(STATE_REG_SCAN_IN), .A2(n3278), .ZN(n5106) );
  AOI21_X1 U3793 ( .B1(n5268), .B2(n4234), .A(n5106), .ZN(n3279) );
  OAI211_X1 U3794 ( .C1(n4214), .C2(n3281), .A(n3280), .B(n3279), .ZN(n3282)
         );
  OR2_X1 U3795 ( .A1(n3283), .A2(n3282), .ZN(U3227) );
  INV_X1 U3796 ( .A(n4230), .ZN(n3364) );
  MUX2_X1 U3797 ( .A(n5074), .B(DATAI_8_), .S(n3794), .Z(n3398) );
  NAND2_X1 U3798 ( .A1(n3364), .A2(n3398), .ZN(n3880) );
  INV_X1 U3799 ( .A(n3398), .ZN(n3418) );
  NAND2_X1 U3800 ( .A1(n4230), .A2(n3418), .ZN(n3876) );
  NAND2_X1 U3801 ( .A1(n4231), .A2(n3408), .ZN(n3284) );
  NOR2_X1 U3802 ( .A1(n3287), .A2(n3838), .ZN(n3288) );
  AOI21_X1 U3803 ( .B1(n3838), .B2(n3287), .A(n3288), .ZN(n5199) );
  INV_X1 U3804 ( .A(n3289), .ZN(n3290) );
  OAI21_X1 U3805 ( .B1(n3290), .B2(n3418), .A(n3368), .ZN(n5198) );
  INV_X1 U3806 ( .A(n5198), .ZN(n3294) );
  INV_X1 U3807 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3292) );
  INV_X1 U3808 ( .A(n3417), .ZN(n3291) );
  OAI22_X1 U3809 ( .A1(n5138), .A2(n3292), .B1(n3291), .B2(n4991), .ZN(n3293)
         );
  AOI21_X1 U3810 ( .B1(n3294), .B2(n5334), .A(n3293), .ZN(n3306) );
  NAND2_X1 U3811 ( .A1(n2494), .A2(REG2_REG_9__SCAN_IN), .ZN(n3300) );
  NAND2_X1 U3812 ( .A1(n3295), .A2(n4561), .ZN(n3296) );
  AND2_X1 U3813 ( .A1(n3358), .A2(n3296), .ZN(n3450) );
  NAND2_X1 U3814 ( .A1(n3109), .A2(n3450), .ZN(n3299) );
  NAND2_X1 U3815 ( .A1(n3056), .A2(REG1_REG_9__SCAN_IN), .ZN(n3298) );
  NAND2_X1 U3816 ( .A1(n3057), .A2(REG0_REG_9__SCAN_IN), .ZN(n3297) );
  XNOR2_X1 U3817 ( .A(n3356), .B(n3286), .ZN(n3302) );
  NAND2_X1 U3818 ( .A1(n3302), .A2(n5124), .ZN(n3304) );
  AOI22_X1 U3819 ( .A1(n4231), .A2(n4957), .B1(n3398), .B2(n5325), .ZN(n3303)
         );
  OAI211_X1 U3820 ( .C1(n3386), .C2(n5127), .A(n3304), .B(n3303), .ZN(n5200)
         );
  NAND2_X1 U3821 ( .A1(n5200), .A2(n5138), .ZN(n3305) );
  OAI211_X1 U3822 ( .C1(n5199), .C2(n5307), .A(n3306), .B(n3305), .ZN(U3282)
         );
  INV_X1 U3823 ( .A(n3307), .ZN(n3308) );
  NOR2_X1 U3824 ( .A1(n3316), .A2(n3308), .ZN(n3309) );
  NAND2_X1 U3825 ( .A1(n3310), .A2(n3309), .ZN(n3320) );
  INV_X1 U3826 ( .A(n3311), .ZN(n3314) );
  INV_X1 U3827 ( .A(n3312), .ZN(n3313) );
  NAND2_X1 U3828 ( .A1(n3314), .A2(n3313), .ZN(n3315) );
  OAI21_X1 U3829 ( .B1(n3317), .B2(n3316), .A(n3315), .ZN(n3318) );
  INV_X1 U3830 ( .A(n3318), .ZN(n3319) );
  NAND2_X1 U3831 ( .A1(n4233), .A2(n3492), .ZN(n3322) );
  NAND2_X1 U3832 ( .A1(n3325), .A2(n4050), .ZN(n3321) );
  NAND2_X1 U3833 ( .A1(n3322), .A2(n3321), .ZN(n3323) );
  XNOR2_X1 U3834 ( .A(n3323), .B(n3024), .ZN(n3327) );
  AND2_X1 U3835 ( .A1(n3325), .A2(n3492), .ZN(n3326) );
  AOI21_X1 U3836 ( .B1(n4233), .B2(n3026), .A(n3326), .ZN(n3328) );
  XNOR2_X1 U3837 ( .A(n3327), .B(n3328), .ZN(n3344) );
  INV_X1 U3838 ( .A(n3327), .ZN(n3329) );
  NAND2_X1 U3839 ( .A1(n3329), .A2(n3328), .ZN(n3330) );
  NAND2_X1 U3840 ( .A1(n4232), .A2(n3492), .ZN(n3332) );
  NAND2_X1 U3841 ( .A1(n3334), .A2(n4050), .ZN(n3331) );
  NAND2_X1 U3842 ( .A1(n3332), .A2(n3331), .ZN(n3333) );
  XNOR2_X1 U3843 ( .A(n3333), .B(n3024), .ZN(n3400) );
  AND2_X1 U3844 ( .A1(n3334), .A2(n3492), .ZN(n3335) );
  AOI21_X1 U3845 ( .B1(n4232), .B2(n3026), .A(n3335), .ZN(n3401) );
  XNOR2_X1 U3846 ( .A(n3400), .B(n3401), .ZN(n3403) );
  XOR2_X1 U3847 ( .A(n3404), .B(n3403), .Z(n3341) );
  AOI22_X1 U3848 ( .A1(n5276), .A2(n4231), .B1(n4183), .B2(n3336), .ZN(n3340)
         );
  AND2_X1 U3849 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n4261) );
  NOR2_X1 U3850 ( .A1(n4214), .A2(n3337), .ZN(n3338) );
  AOI211_X1 U3851 ( .C1(n5268), .C2(n4233), .A(n4261), .B(n3338), .ZN(n3339)
         );
  OAI211_X1 U3852 ( .C1(n3341), .C2(n5271), .A(n3340), .B(n3339), .ZN(U3236)
         );
  OAI21_X1 U3853 ( .B1(n3344), .B2(n3343), .A(n3342), .ZN(n3351) );
  AOI22_X1 U3854 ( .A1(n5276), .A2(n4232), .B1(n4183), .B2(n3345), .ZN(n3348)
         );
  AOI21_X1 U3855 ( .B1(n5268), .B2(n3108), .A(n3346), .ZN(n3347) );
  OAI211_X1 U3856 ( .C1(n4214), .C2(n3349), .A(n3348), .B(n3347), .ZN(n3350)
         );
  AOI21_X1 U3857 ( .B1(n3351), .B2(n4134), .A(n3350), .ZN(n3352) );
  INV_X1 U3858 ( .A(n3352), .ZN(U3224) );
  NAND2_X1 U3859 ( .A1(n3364), .A2(n3418), .ZN(n3353) );
  MUX2_X1 U3860 ( .A(n3355), .B(DATAI_9_), .S(n3794), .Z(n3443) );
  XNOR2_X1 U3861 ( .A(n4229), .B(n3443), .ZN(n3830) );
  XNOR2_X1 U3862 ( .A(n3385), .B(n3830), .ZN(n5207) );
  NAND2_X1 U3863 ( .A1(n3356), .A2(n3838), .ZN(n3357) );
  NAND2_X1 U3864 ( .A1(n3357), .A2(n3876), .ZN(n3374) );
  XNOR2_X1 U3865 ( .A(n3374), .B(n3830), .ZN(n3367) );
  NAND2_X1 U3866 ( .A1(n2494), .A2(REG2_REG_10__SCAN_IN), .ZN(n3363) );
  AND2_X1 U3867 ( .A1(n3358), .A2(n3512), .ZN(n3359) );
  NOR2_X1 U3868 ( .A1(n3376), .A2(n3359), .ZN(n3511) );
  NAND2_X1 U3869 ( .A1(n3109), .A2(n3511), .ZN(n3362) );
  NAND2_X1 U3870 ( .A1(n3056), .A2(REG1_REG_10__SCAN_IN), .ZN(n3361) );
  NAND2_X1 U3871 ( .A1(n3057), .A2(REG0_REG_10__SCAN_IN), .ZN(n3360) );
  NAND4_X1 U3872 ( .A1(n3363), .A2(n3362), .A3(n3361), .A4(n3360), .ZN(n4228)
         );
  OAI22_X1 U3873 ( .A1(n3364), .A2(n5282), .B1(n5315), .B2(n2581), .ZN(n3365)
         );
  AOI21_X1 U3874 ( .B1(n5286), .B2(n4228), .A(n3365), .ZN(n3366) );
  OAI21_X1 U3875 ( .B1(n3367), .B2(n5288), .A(n3366), .ZN(n5209) );
  AOI21_X1 U3876 ( .B1(n3443), .B2(n3368), .A(n3388), .ZN(n5210) );
  INV_X1 U3877 ( .A(n5210), .ZN(n3370) );
  AOI22_X1 U3878 ( .A1(n5333), .A2(REG2_REG_9__SCAN_IN), .B1(n3450), .B2(n5303), .ZN(n3369) );
  OAI21_X1 U3879 ( .B1(n3370), .B2(n5306), .A(n3369), .ZN(n3371) );
  AOI21_X1 U3880 ( .B1(n5209), .B2(n5138), .A(n3371), .ZN(n3372) );
  OAI21_X1 U3881 ( .B1(n5207), .B2(n5307), .A(n3372), .ZN(U3281) );
  INV_X1 U3882 ( .A(n5138), .ZN(n5333) );
  MUX2_X1 U3883 ( .A(n3373), .B(DATAI_10_), .S(n3794), .Z(n3493) );
  NAND2_X1 U3884 ( .A1(n3467), .A2(n3493), .ZN(n3884) );
  NAND2_X1 U3885 ( .A1(n4228), .A2(n3515), .ZN(n3550) );
  NAND2_X1 U3886 ( .A1(n3374), .A2(n3830), .ZN(n3375) );
  NAND2_X1 U3887 ( .A1(n4229), .A2(n2581), .ZN(n3881) );
  NAND2_X1 U3888 ( .A1(n3375), .A2(n3881), .ZN(n3425) );
  XOR2_X1 U3889 ( .A(n3819), .B(n3425), .Z(n3384) );
  NAND2_X1 U3890 ( .A1(n2494), .A2(REG2_REG_11__SCAN_IN), .ZN(n3381) );
  NOR2_X1 U3891 ( .A1(n3376), .A2(REG3_REG_11__SCAN_IN), .ZN(n3377) );
  NOR2_X1 U3892 ( .A1(n3426), .A2(n3377), .ZN(n3531) );
  NAND2_X1 U3893 ( .A1(n3109), .A2(n3531), .ZN(n3380) );
  NAND2_X1 U3894 ( .A1(n3056), .A2(REG1_REG_11__SCAN_IN), .ZN(n3379) );
  NAND2_X1 U3895 ( .A1(n3057), .A2(REG0_REG_11__SCAN_IN), .ZN(n3378) );
  NAND4_X1 U3896 ( .A1(n3381), .A2(n3380), .A3(n3379), .A4(n3378), .ZN(n4227)
         );
  AOI22_X1 U3897 ( .A1(n4227), .A2(n5286), .B1(n5325), .B2(n3493), .ZN(n3382)
         );
  OAI21_X1 U3898 ( .B1(n3386), .B2(n5282), .A(n3382), .ZN(n3383) );
  AOI21_X1 U3899 ( .B1(n3384), .B2(n5124), .A(n3383), .ZN(n5214) );
  XOR2_X1 U3900 ( .A(n3819), .B(n3470), .Z(n5217) );
  NAND2_X1 U3901 ( .A1(n5217), .A2(n4986), .ZN(n3394) );
  INV_X1 U3902 ( .A(n3436), .ZN(n3387) );
  OAI21_X1 U3903 ( .B1(n3388), .B2(n3515), .A(n3387), .ZN(n5215) );
  INV_X1 U3904 ( .A(n5215), .ZN(n3392) );
  INV_X1 U3905 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3390) );
  INV_X1 U3906 ( .A(n3511), .ZN(n3389) );
  OAI22_X1 U3907 ( .A1(n5138), .A2(n3390), .B1(n3389), .B2(n4991), .ZN(n3391)
         );
  AOI21_X1 U3908 ( .B1(n3392), .B2(n5334), .A(n3391), .ZN(n3393) );
  OAI211_X1 U3909 ( .C1(n5333), .C2(n5214), .A(n3394), .B(n3393), .ZN(U3280)
         );
  NAND2_X1 U3910 ( .A1(n4230), .A2(n3492), .ZN(n3396) );
  NAND2_X1 U3911 ( .A1(n3398), .A2(n4050), .ZN(n3395) );
  NAND2_X1 U3912 ( .A1(n3396), .A2(n3395), .ZN(n3397) );
  XNOR2_X1 U3913 ( .A(n3397), .B(n3024), .ZN(n3445) );
  AND2_X1 U3914 ( .A1(n3398), .A2(n3492), .ZN(n3399) );
  AOI21_X1 U3915 ( .B1(n4230), .B2(n3026), .A(n3399), .ZN(n3446) );
  XNOR2_X1 U3916 ( .A(n3445), .B(n3446), .ZN(n3415) );
  INV_X1 U3917 ( .A(n3400), .ZN(n3402) );
  NAND2_X1 U3918 ( .A1(n4231), .A2(n3492), .ZN(n3406) );
  NAND2_X1 U3919 ( .A1(n3408), .A2(n4050), .ZN(n3405) );
  NAND2_X1 U3920 ( .A1(n3406), .A2(n3405), .ZN(n3407) );
  XNOR2_X1 U3921 ( .A(n3407), .B(n3024), .ZN(n3412) );
  AND2_X1 U3922 ( .A1(n3408), .A2(n3492), .ZN(n3409) );
  AOI21_X1 U3923 ( .B1(n4231), .B2(n3026), .A(n3409), .ZN(n3410) );
  XNOR2_X1 U3924 ( .A(n3412), .B(n3410), .ZN(n4136) );
  NAND2_X1 U3925 ( .A1(n3507), .A2(n4136), .ZN(n4135) );
  INV_X1 U3926 ( .A(n3410), .ZN(n3411) );
  NAND2_X1 U3927 ( .A1(n3412), .A2(n3411), .ZN(n3413) );
  AND2_X1 U3928 ( .A1(n4135), .A2(n3413), .ZN(n3414) );
  NAND2_X1 U3929 ( .A1(n4135), .A2(n3500), .ZN(n3448) );
  OAI21_X1 U3930 ( .B1(n3415), .B2(n3414), .A(n3448), .ZN(n3416) );
  INV_X1 U3931 ( .A(n3416), .ZN(n3422) );
  AOI22_X1 U3932 ( .A1(n5276), .A2(n4229), .B1(n4183), .B2(n3417), .ZN(n3421)
         );
  INV_X1 U3933 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4736) );
  NOR2_X1 U3934 ( .A1(STATE_REG_SCAN_IN), .A2(n4736), .ZN(n4271) );
  NOR2_X1 U3935 ( .A1(n4214), .A2(n3418), .ZN(n3419) );
  AOI211_X1 U3936 ( .C1(n5268), .C2(n4231), .A(n4271), .B(n3419), .ZN(n3420)
         );
  OAI211_X1 U3937 ( .C1(n3422), .C2(n5271), .A(n3421), .B(n3420), .ZN(U3218)
         );
  INV_X1 U3938 ( .A(n4227), .ZN(n3424) );
  MUX2_X1 U3939 ( .A(n3423), .B(DATAI_11_), .S(n3794), .Z(n3526) );
  NAND2_X1 U3940 ( .A1(n3424), .A2(n3526), .ZN(n3554) );
  NAND2_X1 U3941 ( .A1(n4227), .A2(n3532), .ZN(n3461) );
  NAND2_X1 U3942 ( .A1(n3425), .A2(n3884), .ZN(n3559) );
  NAND2_X1 U3943 ( .A1(n3559), .A2(n3550), .ZN(n3462) );
  XOR2_X1 U3944 ( .A(n3820), .B(n3462), .Z(n3434) );
  NAND2_X1 U3945 ( .A1(n2494), .A2(REG2_REG_12__SCAN_IN), .ZN(n3431) );
  OR2_X1 U3946 ( .A1(n3426), .A2(REG3_REG_12__SCAN_IN), .ZN(n3427) );
  AND2_X1 U3947 ( .A1(n3455), .A2(n3427), .ZN(n3624) );
  NAND2_X1 U3948 ( .A1(n3109), .A2(n3624), .ZN(n3430) );
  NAND2_X1 U3949 ( .A1(n3056), .A2(REG1_REG_12__SCAN_IN), .ZN(n3429) );
  NAND2_X1 U3950 ( .A1(n3057), .A2(REG0_REG_12__SCAN_IN), .ZN(n3428) );
  NAND4_X1 U3951 ( .A1(n3431), .A2(n3430), .A3(n3429), .A4(n3428), .ZN(n4226)
         );
  INV_X1 U3952 ( .A(n4226), .ZN(n3581) );
  AOI22_X1 U3953 ( .A1(n4228), .A2(n4957), .B1(n3526), .B2(n5325), .ZN(n3432)
         );
  OAI21_X1 U3954 ( .B1(n3581), .B2(n5127), .A(n3432), .ZN(n3433) );
  AOI21_X1 U3955 ( .B1(n3434), .B2(n5124), .A(n3433), .ZN(n5223) );
  OAI22_X1 U3956 ( .A1(n3470), .A2(n3819), .B1(n3467), .B2(n3515), .ZN(n3435)
         );
  XNOR2_X1 U3957 ( .A(n3435), .B(n3820), .ZN(n5226) );
  OAI21_X1 U3958 ( .B1(n3436), .B2(n3532), .A(n3474), .ZN(n5224) );
  AOI22_X1 U3959 ( .A1(n5333), .A2(REG2_REG_11__SCAN_IN), .B1(n3531), .B2(
        n5303), .ZN(n3437) );
  OAI21_X1 U3960 ( .B1(n5224), .B2(n5306), .A(n3437), .ZN(n3438) );
  AOI21_X1 U3961 ( .B1(n5226), .B2(n4986), .A(n3438), .ZN(n3439) );
  OAI21_X1 U3962 ( .B1(n5333), .B2(n5223), .A(n3439), .ZN(U3279) );
  NAND2_X1 U3963 ( .A1(n4229), .A2(n3492), .ZN(n3441) );
  NAND2_X1 U3964 ( .A1(n3443), .A2(n4050), .ZN(n3440) );
  NAND2_X1 U3965 ( .A1(n3441), .A2(n3440), .ZN(n3442) );
  XNOR2_X1 U3966 ( .A(n3442), .B(n3024), .ZN(n3495) );
  AND2_X1 U3967 ( .A1(n3443), .A2(n3492), .ZN(n3444) );
  AOI21_X1 U3968 ( .B1(n4229), .B2(n3026), .A(n3444), .ZN(n3496) );
  XNOR2_X1 U3969 ( .A(n3495), .B(n3496), .ZN(n3503) );
  INV_X1 U3970 ( .A(n3445), .ZN(n3447) );
  NAND2_X1 U3971 ( .A1(n3447), .A2(n3446), .ZN(n3498) );
  NAND2_X1 U3972 ( .A1(n3448), .A2(n3498), .ZN(n3449) );
  XOR2_X1 U3973 ( .A(n3503), .B(n3449), .Z(n3454) );
  AOI22_X1 U3974 ( .A1(n4219), .A2(n4228), .B1(n4183), .B2(n3450), .ZN(n3453)
         );
  NOR2_X1 U3975 ( .A1(STATE_REG_SCAN_IN), .A2(n4561), .ZN(n4279) );
  NOR2_X1 U3976 ( .A1(n4214), .A2(n2581), .ZN(n3451) );
  AOI211_X1 U3977 ( .C1(n5268), .C2(n4230), .A(n4279), .B(n3451), .ZN(n3452)
         );
  OAI211_X1 U3978 ( .C1(n3454), .C2(n5271), .A(n3453), .B(n3452), .ZN(U3228)
         );
  NAND2_X1 U3979 ( .A1(n3057), .A2(REG0_REG_13__SCAN_IN), .ZN(n3460) );
  NAND2_X1 U3980 ( .A1(n3056), .A2(REG1_REG_13__SCAN_IN), .ZN(n3459) );
  NAND2_X1 U3981 ( .A1(n3455), .A2(n4759), .ZN(n3456) );
  AND2_X1 U3982 ( .A1(n3542), .A2(n3456), .ZN(n3648) );
  NAND2_X1 U3983 ( .A1(n3109), .A2(n3648), .ZN(n3458) );
  NAND2_X1 U3984 ( .A1(n2494), .A2(REG2_REG_13__SCAN_IN), .ZN(n3457) );
  NAND4_X1 U3985 ( .A1(n3460), .A2(n3459), .A3(n3458), .A4(n3457), .ZN(n4225)
         );
  INV_X1 U3986 ( .A(n4225), .ZN(n3566) );
  INV_X1 U3987 ( .A(n3461), .ZN(n3552) );
  AOI21_X1 U3988 ( .B1(n3462), .B2(n3820), .A(n3552), .ZN(n3579) );
  MUX2_X1 U3989 ( .A(n3463), .B(DATAI_12_), .S(n3794), .Z(n3611) );
  NAND2_X1 U3990 ( .A1(n3581), .A2(n3611), .ZN(n3553) );
  INV_X1 U3991 ( .A(n3611), .ZN(n3626) );
  NAND2_X1 U3992 ( .A1(n4226), .A2(n3626), .ZN(n3577) );
  NAND2_X1 U3993 ( .A1(n3553), .A2(n3577), .ZN(n3578) );
  INV_X1 U3994 ( .A(n3578), .ZN(n3821) );
  XNOR2_X1 U3995 ( .A(n3579), .B(n3821), .ZN(n3464) );
  NAND2_X1 U3996 ( .A1(n3464), .A2(n5124), .ZN(n3466) );
  AOI22_X1 U3997 ( .A1(n4227), .A2(n4957), .B1(n3611), .B2(n5325), .ZN(n3465)
         );
  OAI211_X1 U3998 ( .C1(n3566), .C2(n5127), .A(n3466), .B(n3465), .ZN(n5233)
         );
  INV_X1 U3999 ( .A(n5233), .ZN(n3478) );
  OAI21_X1 U4000 ( .B1(n3470), .B2(n3819), .A(n3469), .ZN(n3472) );
  NAND2_X1 U4001 ( .A1(n3472), .A2(n3471), .ZN(n3473) );
  NAND2_X1 U4002 ( .A1(n3473), .A2(n3578), .ZN(n3539) );
  OAI21_X1 U4003 ( .B1(n3473), .B2(n3578), .A(n3539), .ZN(n5235) );
  OAI21_X1 U4004 ( .B1(n2577), .B2(n3626), .A(n3586), .ZN(n5232) );
  AOI22_X1 U4005 ( .A1(n5333), .A2(REG2_REG_12__SCAN_IN), .B1(n3624), .B2(
        n5303), .ZN(n3475) );
  OAI21_X1 U4006 ( .B1(n5232), .B2(n5306), .A(n3475), .ZN(n3476) );
  AOI21_X1 U4007 ( .B1(n5235), .B2(n4986), .A(n3476), .ZN(n3477) );
  OAI21_X1 U4008 ( .B1(n5333), .B2(n3478), .A(n3477), .ZN(U3278) );
  AOI211_X1 U4009 ( .C1(n2536), .C2(n3480), .A(n3479), .B(n5108), .ZN(n3487)
         );
  OAI211_X1 U4010 ( .C1(n3483), .C2(n3482), .A(n5116), .B(n3481), .ZN(n3485)
         );
  AND2_X1 U4011 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n3534) );
  AOI21_X1 U4012 ( .B1(n5107), .B2(ADDR_REG_11__SCAN_IN), .A(n3534), .ZN(n3484) );
  OAI211_X1 U4013 ( .C1(n4348), .C2(n5222), .A(n3485), .B(n3484), .ZN(n3486)
         );
  OR2_X1 U4014 ( .A1(n3487), .A2(n3486), .ZN(U3251) );
  NAND2_X1 U4015 ( .A1(n4228), .A2(n3492), .ZN(n3489) );
  NAND2_X1 U4016 ( .A1(n3493), .A2(n4050), .ZN(n3488) );
  NAND2_X1 U4017 ( .A1(n3489), .A2(n3488), .ZN(n3491) );
  XNOR2_X1 U4018 ( .A(n3491), .B(n3490), .ZN(n3518) );
  AND2_X1 U4019 ( .A1(n3493), .A2(n3492), .ZN(n3494) );
  AOI21_X1 U4020 ( .B1(n4228), .B2(n3026), .A(n3494), .ZN(n3519) );
  XNOR2_X1 U4021 ( .A(n3518), .B(n3519), .ZN(n3510) );
  INV_X1 U4022 ( .A(n3495), .ZN(n3497) );
  NAND2_X1 U4023 ( .A1(n3497), .A2(n3496), .ZN(n3502) );
  AND2_X1 U4024 ( .A1(n3498), .A2(n3502), .ZN(n3499) );
  AND2_X1 U4025 ( .A1(n4136), .A2(n3499), .ZN(n3506) );
  INV_X1 U4026 ( .A(n3499), .ZN(n3501) );
  INV_X1 U4027 ( .A(n3502), .ZN(n3504) );
  INV_X1 U4028 ( .A(n3523), .ZN(n3508) );
  AOI211_X1 U4029 ( .C1(n3510), .C2(n3509), .A(n5271), .B(n3508), .ZN(n3517)
         );
  AOI22_X1 U4030 ( .A1(n5276), .A2(n4227), .B1(n4183), .B2(n3511), .ZN(n3514)
         );
  NOR2_X1 U4031 ( .A1(STATE_REG_SCAN_IN), .A2(n3512), .ZN(n4292) );
  AOI21_X1 U4032 ( .B1(n5268), .B2(n4229), .A(n4292), .ZN(n3513) );
  OAI211_X1 U4033 ( .C1(n4214), .C2(n3515), .A(n3514), .B(n3513), .ZN(n3516)
         );
  OR2_X1 U4034 ( .A1(n3517), .A2(n3516), .ZN(U3214) );
  INV_X1 U4035 ( .A(n3518), .ZN(n3521) );
  INV_X1 U4036 ( .A(n3519), .ZN(n3520) );
  NAND2_X1 U4037 ( .A1(n3521), .A2(n3520), .ZN(n3522) );
  NAND2_X1 U4038 ( .A1(n4227), .A2(n3026), .ZN(n3525) );
  NAND2_X1 U4039 ( .A1(n3526), .A2(n3492), .ZN(n3524) );
  NAND2_X1 U4040 ( .A1(n3525), .A2(n3524), .ZN(n3618) );
  NAND2_X1 U4041 ( .A1(n4227), .A2(n3492), .ZN(n3528) );
  NAND2_X1 U4042 ( .A1(n3526), .A2(n4050), .ZN(n3527) );
  NAND2_X1 U40430 ( .A1(n3528), .A2(n3527), .ZN(n3529) );
  XNOR2_X1 U4044 ( .A(n3529), .B(n3024), .ZN(n3619) );
  XOR2_X1 U4045 ( .A(n3618), .B(n3619), .Z(n3530) );
  XNOR2_X1 U4046 ( .A(n3620), .B(n3530), .ZN(n3537) );
  AOI22_X1 U4047 ( .A1(n5276), .A2(n4226), .B1(n4183), .B2(n3531), .ZN(n3536)
         );
  NOR2_X1 U4048 ( .A1(n4214), .A2(n3532), .ZN(n3533) );
  AOI211_X1 U4049 ( .C1(n5268), .C2(n4228), .A(n3534), .B(n3533), .ZN(n3535)
         );
  OAI211_X1 U4050 ( .C1(n3537), .C2(n5271), .A(n3536), .B(n3535), .ZN(U3233)
         );
  NAND2_X1 U4051 ( .A1(n3539), .A2(n3538), .ZN(n3576) );
  MUX2_X1 U4052 ( .A(n3540), .B(DATAI_13_), .S(n3794), .Z(n3634) );
  NAND2_X1 U4053 ( .A1(n4225), .A2(n3634), .ZN(n3541) );
  NAND2_X1 U4054 ( .A1(n2494), .A2(REG2_REG_14__SCAN_IN), .ZN(n3546) );
  AOI21_X1 U4055 ( .B1(n3542), .B2(n4726), .A(n3560), .ZN(n3932) );
  NAND2_X1 U4056 ( .A1(n3109), .A2(n3932), .ZN(n3545) );
  NAND2_X1 U4057 ( .A1(n3056), .A2(REG1_REG_14__SCAN_IN), .ZN(n3544) );
  NAND2_X1 U4058 ( .A1(n3057), .A2(REG0_REG_14__SCAN_IN), .ZN(n3543) );
  NAND4_X1 U4059 ( .A1(n3546), .A2(n3545), .A3(n3544), .A4(n3543), .ZN(n4224)
         );
  INV_X1 U4060 ( .A(n4224), .ZN(n3548) );
  MUX2_X1 U4061 ( .A(n3547), .B(DATAI_14_), .S(n3794), .Z(n3921) );
  NAND2_X1 U4062 ( .A1(n3548), .A2(n3921), .ZN(n3760) );
  NAND2_X1 U4063 ( .A1(n4224), .A2(n3933), .ZN(n3761) );
  XNOR2_X1 U4064 ( .A(n3591), .B(n3843), .ZN(n5251) );
  INV_X1 U4065 ( .A(n5251), .ZN(n3575) );
  NAND2_X1 U4066 ( .A1(n4225), .A2(n3649), .ZN(n3549) );
  NAND2_X1 U4067 ( .A1(n3577), .A2(n3549), .ZN(n3557) );
  INV_X1 U4068 ( .A(n3550), .ZN(n3551) );
  NOR3_X1 U4069 ( .A1(n3557), .A2(n3552), .A3(n3551), .ZN(n3889) );
  INV_X1 U4070 ( .A(n3553), .ZN(n3556) );
  INV_X1 U4071 ( .A(n3554), .ZN(n3555) );
  NOR2_X1 U4072 ( .A1(n3556), .A2(n3555), .ZN(n3558) );
  OAI22_X1 U4073 ( .A1(n3558), .A2(n3557), .B1(n3649), .B2(n4225), .ZN(n3888)
         );
  AOI21_X2 U4074 ( .B1(n3559), .B2(n3889), .A(n3888), .ZN(n3765) );
  AOI21_X1 U4075 ( .B1(n3765), .B2(n2715), .A(n3671), .ZN(n3569) );
  OAI21_X1 U4076 ( .B1(n3560), .B2(REG3_REG_15__SCAN_IN), .A(n3594), .ZN(n3561) );
  INV_X1 U4077 ( .A(n3561), .ZN(n3973) );
  NAND2_X1 U4078 ( .A1(n3109), .A2(n3973), .ZN(n3565) );
  NAND2_X1 U4079 ( .A1(n3057), .A2(REG0_REG_15__SCAN_IN), .ZN(n3564) );
  NAND2_X1 U4080 ( .A1(n3056), .A2(REG1_REG_15__SCAN_IN), .ZN(n3563) );
  NAND2_X1 U4081 ( .A1(n2494), .A2(REG2_REG_15__SCAN_IN), .ZN(n3562) );
  NAND4_X1 U4082 ( .A1(n3565), .A2(n3564), .A3(n3563), .A4(n3562), .ZN(n5267)
         );
  OAI22_X1 U4083 ( .A1(n3566), .A2(n5282), .B1(n3933), .B2(n5315), .ZN(n3567)
         );
  AOI21_X1 U4084 ( .B1(n5286), .B2(n5267), .A(n3567), .ZN(n3568) );
  OAI21_X1 U4085 ( .B1(n3569), .B2(n5288), .A(n3568), .ZN(n5249) );
  INV_X1 U4086 ( .A(n3585), .ZN(n3570) );
  AOI211_X1 U4087 ( .C1(n3921), .C2(n3570), .A(n5296), .B(n3603), .ZN(n5250)
         );
  INV_X1 U4088 ( .A(n5250), .ZN(n3572) );
  INV_X1 U4089 ( .A(n4390), .ZN(n4969) );
  AOI22_X1 U4090 ( .A1(n5333), .A2(REG2_REG_14__SCAN_IN), .B1(n3932), .B2(
        n5303), .ZN(n3571) );
  OAI21_X1 U4091 ( .B1(n3572), .B2(n4969), .A(n3571), .ZN(n3573) );
  AOI21_X1 U4092 ( .B1(n5249), .B2(n5138), .A(n3573), .ZN(n3574) );
  OAI21_X1 U4093 ( .B1(n3575), .B2(n5307), .A(n3574), .ZN(U3276) );
  XNOR2_X1 U4094 ( .A(n4225), .B(n3634), .ZN(n3815) );
  XNOR2_X1 U4095 ( .A(n3576), .B(n3815), .ZN(n5241) );
  OAI21_X1 U4096 ( .B1(n3579), .B2(n3578), .A(n3577), .ZN(n3580) );
  XNOR2_X1 U4097 ( .A(n3580), .B(n3815), .ZN(n3584) );
  OAI22_X1 U4098 ( .A1(n3581), .A2(n5282), .B1(n3649), .B2(n5315), .ZN(n3582)
         );
  AOI21_X1 U4099 ( .B1(n5286), .B2(n4224), .A(n3582), .ZN(n3583) );
  OAI21_X1 U4100 ( .B1(n3584), .B2(n5288), .A(n3583), .ZN(n5243) );
  AOI21_X1 U4101 ( .B1(n3634), .B2(n3586), .A(n3585), .ZN(n5244) );
  INV_X1 U4102 ( .A(n5244), .ZN(n3588) );
  AOI22_X1 U4103 ( .A1(n5333), .A2(REG2_REG_13__SCAN_IN), .B1(n3648), .B2(
        n5303), .ZN(n3587) );
  OAI21_X1 U4104 ( .B1(n3588), .B2(n5306), .A(n3587), .ZN(n3589) );
  AOI21_X1 U4105 ( .B1(n5243), .B2(n5138), .A(n3589), .ZN(n3590) );
  OAI21_X1 U4106 ( .B1(n5241), .B2(n5307), .A(n3590), .ZN(U3277) );
  MUX2_X1 U4107 ( .A(n5073), .B(DATAI_15_), .S(n3794), .Z(n3966) );
  XNOR2_X1 U4108 ( .A(n5267), .B(n3974), .ZN(n3828) );
  XNOR2_X1 U4109 ( .A(n3656), .B(n3828), .ZN(n5259) );
  INV_X1 U4110 ( .A(n3760), .ZN(n3670) );
  NOR2_X1 U4111 ( .A1(n3671), .A2(n3670), .ZN(n3592) );
  XNOR2_X1 U4112 ( .A(n3592), .B(n3828), .ZN(n3602) );
  NAND2_X1 U4113 ( .A1(n3057), .A2(REG0_REG_16__SCAN_IN), .ZN(n3599) );
  NAND2_X1 U4114 ( .A1(n3056), .A2(REG1_REG_16__SCAN_IN), .ZN(n3598) );
  INV_X1 U4115 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4553) );
  NAND2_X1 U4116 ( .A1(n3594), .A2(n4553), .ZN(n3595) );
  AND2_X1 U4117 ( .A1(n3659), .A2(n3595), .ZN(n5304) );
  NAND2_X1 U4118 ( .A1(n3109), .A2(n5304), .ZN(n3597) );
  NAND2_X1 U4119 ( .A1(n2494), .A2(REG2_REG_16__SCAN_IN), .ZN(n3596) );
  NAND4_X1 U4120 ( .A1(n3599), .A2(n3598), .A3(n3597), .A4(n3596), .ZN(n4223)
         );
  AOI22_X1 U4121 ( .A1(n4224), .A2(n4957), .B1(n3966), .B2(n5325), .ZN(n3600)
         );
  OAI21_X1 U4122 ( .B1(n2716), .B2(n5127), .A(n3600), .ZN(n3601) );
  AOI21_X1 U4123 ( .B1(n3602), .B2(n5124), .A(n3601), .ZN(n5255) );
  NOR2_X1 U4124 ( .A1(n5255), .A2(n5333), .ZN(n3606) );
  OAI21_X1 U4125 ( .B1(n3603), .B2(n3974), .A(n5292), .ZN(n5256) );
  AOI22_X1 U4126 ( .A1(n5333), .A2(REG2_REG_15__SCAN_IN), .B1(n5303), .B2(
        n3973), .ZN(n3604) );
  OAI21_X1 U4127 ( .B1(n5256), .B2(n5306), .A(n3604), .ZN(n3605) );
  AOI211_X1 U4128 ( .C1(n5259), .C2(n4986), .A(n3606), .B(n3605), .ZN(n3607)
         );
  INV_X1 U4129 ( .A(n3607), .ZN(U3275) );
  NAND2_X1 U4130 ( .A1(n4226), .A2(n3492), .ZN(n3609) );
  NAND2_X1 U4131 ( .A1(n3611), .A2(n4050), .ZN(n3608) );
  NAND2_X1 U4132 ( .A1(n3609), .A2(n3608), .ZN(n3610) );
  XNOR2_X1 U4133 ( .A(n3610), .B(n3490), .ZN(n3613) );
  AND2_X1 U4134 ( .A1(n3611), .A2(n3492), .ZN(n3612) );
  AOI21_X1 U4135 ( .B1(n4226), .B2(n3026), .A(n3612), .ZN(n3614) );
  NAND2_X1 U4136 ( .A1(n3613), .A2(n3614), .ZN(n3642) );
  INV_X1 U4137 ( .A(n3613), .ZN(n3616) );
  INV_X1 U4138 ( .A(n3614), .ZN(n3615) );
  NAND2_X1 U4139 ( .A1(n3616), .A2(n3615), .ZN(n3617) );
  NAND2_X1 U4140 ( .A1(n3642), .A2(n3617), .ZN(n3623) );
  INV_X1 U4141 ( .A(n3643), .ZN(n3621) );
  AOI21_X1 U4142 ( .B1(n3623), .B2(n3622), .A(n3621), .ZN(n3630) );
  AOI22_X1 U4143 ( .A1(n5276), .A2(n4225), .B1(n4183), .B2(n3624), .ZN(n3629)
         );
  INV_X1 U4144 ( .A(REG3_REG_12__SCAN_IN), .ZN(n3625) );
  NOR2_X1 U4145 ( .A1(STATE_REG_SCAN_IN), .A2(n3625), .ZN(n4302) );
  NOR2_X1 U4146 ( .A1(n4214), .A2(n3626), .ZN(n3627) );
  AOI211_X1 U4147 ( .C1(n5268), .C2(n4227), .A(n4302), .B(n3627), .ZN(n3628)
         );
  OAI211_X1 U4148 ( .C1(n3630), .C2(n5271), .A(n3629), .B(n3628), .ZN(U3221)
         );
  NAND2_X1 U4149 ( .A1(n4225), .A2(n3492), .ZN(n3632) );
  NAND2_X1 U4150 ( .A1(n3634), .A2(n4050), .ZN(n3631) );
  NAND2_X1 U4151 ( .A1(n3632), .A2(n3631), .ZN(n3633) );
  XNOR2_X1 U4152 ( .A(n3633), .B(n3490), .ZN(n3636) );
  AND2_X1 U4153 ( .A1(n3634), .A2(n3492), .ZN(n3635) );
  AOI21_X1 U4154 ( .B1(n4225), .B2(n3026), .A(n3635), .ZN(n3637) );
  NAND2_X1 U4155 ( .A1(n3636), .A2(n3637), .ZN(n3928) );
  INV_X1 U4156 ( .A(n3636), .ZN(n3639) );
  INV_X1 U4157 ( .A(n3637), .ZN(n3638) );
  NAND2_X1 U4158 ( .A1(n3639), .A2(n3638), .ZN(n3640) );
  INV_X1 U4159 ( .A(n3642), .ZN(n3641) );
  NOR2_X1 U4160 ( .A1(n3644), .A2(n3641), .ZN(n3647) );
  NAND2_X1 U4161 ( .A1(n3643), .A2(n3642), .ZN(n3645) );
  NAND2_X1 U4162 ( .A1(n3645), .A2(n3644), .ZN(n3929) );
  INV_X1 U4163 ( .A(n3929), .ZN(n3646) );
  AOI21_X1 U4164 ( .B1(n3647), .B2(n3643), .A(n3646), .ZN(n3653) );
  AOI22_X1 U4165 ( .A1(n4219), .A2(n4224), .B1(n4183), .B2(n3648), .ZN(n3652)
         );
  NOR2_X1 U4166 ( .A1(STATE_REG_SCAN_IN), .A2(n4759), .ZN(n3944) );
  NOR2_X1 U4167 ( .A1(n4214), .A2(n3649), .ZN(n3650) );
  AOI211_X1 U4168 ( .C1(n5268), .C2(n4226), .A(n3944), .B(n3650), .ZN(n3651)
         );
  OAI211_X1 U4169 ( .C1(n3653), .C2(n5271), .A(n3652), .B(n3651), .ZN(U3231)
         );
  MUX2_X1 U4170 ( .A(n3654), .B(DATAI_16_), .S(n3794), .Z(n5265) );
  MUX2_X1 U4171 ( .A(n5072), .B(DATAI_17_), .S(n3794), .Z(n3998) );
  INV_X1 U4172 ( .A(n3998), .ZN(n3667) );
  OAI21_X1 U4173 ( .B1(n2586), .B2(n3667), .A(n3956), .ZN(n5048) );
  NOR2_X1 U4174 ( .A1(n5267), .A2(n3966), .ZN(n3655) );
  INV_X1 U4175 ( .A(n5267), .ZN(n5283) );
  INV_X1 U4176 ( .A(n5265), .ZN(n5294) );
  NAND2_X1 U4177 ( .A1(n4223), .A2(n5294), .ZN(n3766) );
  INV_X1 U4178 ( .A(n3766), .ZN(n3672) );
  NOR2_X1 U4179 ( .A1(n4223), .A2(n5294), .ZN(n3894) );
  INV_X1 U4180 ( .A(n5290), .ZN(n3657) );
  NAND2_X1 U4181 ( .A1(n3057), .A2(REG0_REG_17__SCAN_IN), .ZN(n3665) );
  NAND2_X1 U4182 ( .A1(n3056), .A2(REG1_REG_17__SCAN_IN), .ZN(n3664) );
  INV_X1 U4183 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4749) );
  NAND2_X1 U4184 ( .A1(n3659), .A2(n4749), .ZN(n3660) );
  NAND2_X1 U4185 ( .A1(n3674), .A2(n3660), .ZN(n3995) );
  INV_X1 U4186 ( .A(n3995), .ZN(n3661) );
  NAND2_X1 U4187 ( .A1(n3109), .A2(n3661), .ZN(n3663) );
  NAND2_X1 U4188 ( .A1(n2494), .A2(REG2_REG_17__SCAN_IN), .ZN(n3662) );
  NAND4_X1 U4189 ( .A1(n3665), .A2(n3664), .A3(n3663), .A4(n3662), .ZN(n5285)
         );
  INV_X1 U4190 ( .A(n5285), .ZN(n3666) );
  NAND2_X1 U4191 ( .A1(n3666), .A2(n3998), .ZN(n3951) );
  NAND2_X1 U4192 ( .A1(n5285), .A2(n3667), .ZN(n3767) );
  NAND2_X1 U4193 ( .A1(n3951), .A2(n3767), .ZN(n3669) );
  NAND2_X1 U4194 ( .A1(n3668), .A2(n3669), .ZN(n3950) );
  OAI21_X1 U4195 ( .B1(n3668), .B2(n3669), .A(n3950), .ZN(n5045) );
  NAND2_X1 U4196 ( .A1(n5045), .A2(n4986), .ZN(n3687) );
  INV_X1 U4197 ( .A(n3669), .ZN(n3822) );
  NOR2_X1 U4198 ( .A1(n4395), .A2(n3672), .ZN(n3673) );
  NAND2_X1 U4199 ( .A1(n3673), .A2(n3822), .ZN(n3952) );
  OAI21_X1 U4200 ( .B1(n3822), .B2(n3673), .A(n3952), .ZN(n3682) );
  NAND2_X1 U4201 ( .A1(n2494), .A2(REG2_REG_18__SCAN_IN), .ZN(n3679) );
  INV_X1 U4202 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4014) );
  NAND2_X1 U4203 ( .A1(n3674), .A2(n4014), .ZN(n3675) );
  AND2_X1 U4204 ( .A1(n3749), .A2(n3675), .ZN(n4013) );
  NAND2_X1 U4205 ( .A1(n3109), .A2(n4013), .ZN(n3678) );
  NAND2_X1 U4206 ( .A1(n3056), .A2(REG1_REG_18__SCAN_IN), .ZN(n3677) );
  NAND2_X1 U4207 ( .A1(n3057), .A2(REG0_REG_18__SCAN_IN), .ZN(n3676) );
  NAND4_X1 U4208 ( .A1(n3679), .A2(n3678), .A3(n3677), .A4(n3676), .ZN(n4371)
         );
  INV_X1 U4209 ( .A(n4371), .ZN(n4973) );
  AOI22_X1 U4210 ( .A1(n4223), .A2(n4957), .B1(n5325), .B2(n3998), .ZN(n3680)
         );
  OAI21_X1 U4211 ( .B1(n4973), .B2(n5127), .A(n3680), .ZN(n3681) );
  AOI21_X1 U4212 ( .B1(n3682), .B2(n5124), .A(n3681), .ZN(n5046) );
  OAI21_X1 U4213 ( .B1(n3995), .B2(n4991), .A(n5046), .ZN(n3685) );
  INV_X1 U4214 ( .A(REG2_REG_17__SCAN_IN), .ZN(n3683) );
  NOR2_X1 U4215 ( .A1(n5138), .A2(n3683), .ZN(n3684) );
  AOI21_X1 U4216 ( .B1(n3685), .B2(n5138), .A(n3684), .ZN(n3686) );
  OAI211_X1 U4217 ( .C1(n5048), .C2(n5306), .A(n3687), .B(n3686), .ZN(U3273)
         );
  INV_X1 U4218 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4195) );
  AND2_X1 U4219 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n3689) );
  INV_X1 U4220 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3730) );
  INV_X1 U4221 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4184) );
  INV_X1 U4222 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4215) );
  NAND2_X1 U4223 ( .A1(n3701), .A2(n4215), .ZN(n3692) );
  NAND2_X1 U4224 ( .A1(n3779), .A2(n3692), .ZN(n4468) );
  INV_X1 U4225 ( .A(REG1_REG_26__SCAN_IN), .ZN(n3695) );
  NAND2_X1 U4226 ( .A1(n2494), .A2(REG2_REG_26__SCAN_IN), .ZN(n3694) );
  NAND2_X1 U4227 ( .A1(n3057), .A2(REG0_REG_26__SCAN_IN), .ZN(n3693) );
  OAI211_X1 U4228 ( .C1(n3695), .C2(n2923), .A(n3694), .B(n3693), .ZN(n3696)
         );
  INV_X1 U4229 ( .A(n3696), .ZN(n3697) );
  NAND2_X1 U4230 ( .A1(n3794), .A2(DATAI_26_), .ZN(n4467) );
  NOR2_X1 U4231 ( .A1(n4481), .A2(n4467), .ZN(n3708) );
  INV_X1 U4232 ( .A(n3699), .ZN(n3710) );
  INV_X1 U4233 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4741) );
  NAND2_X1 U4234 ( .A1(n3710), .A2(n4741), .ZN(n3700) );
  NAND2_X1 U4235 ( .A1(n3701), .A2(n3700), .ZN(n4094) );
  INV_X1 U4236 ( .A(REG1_REG_25__SCAN_IN), .ZN(n3704) );
  NAND2_X1 U4237 ( .A1(n2494), .A2(REG2_REG_25__SCAN_IN), .ZN(n3703) );
  NAND2_X1 U4238 ( .A1(n3057), .A2(REG0_REG_25__SCAN_IN), .ZN(n3702) );
  OAI211_X1 U4239 ( .C1(n3704), .C2(n2923), .A(n3703), .B(n3702), .ZN(n3705)
         );
  INV_X1 U4240 ( .A(n3705), .ZN(n3706) );
  NAND2_X1 U4241 ( .A1(n3794), .A2(DATAI_25_), .ZN(n4478) );
  INV_X1 U4242 ( .A(n4478), .ZN(n4485) );
  NOR2_X1 U4243 ( .A1(n3708), .A2(n3809), .ZN(n3854) );
  NAND2_X1 U4244 ( .A1(n4889), .A2(n4478), .ZN(n3810) );
  INV_X1 U4245 ( .A(n3810), .ZN(n4405) );
  NAND2_X1 U4246 ( .A1(n3733), .A2(n4184), .ZN(n3709) );
  NAND2_X1 U4247 ( .A1(n4893), .A2(n3109), .ZN(n3716) );
  INV_X1 U4248 ( .A(REG1_REG_24__SCAN_IN), .ZN(n3713) );
  NAND2_X1 U4249 ( .A1(n2494), .A2(REG2_REG_24__SCAN_IN), .ZN(n3712) );
  NAND2_X1 U4250 ( .A1(n3057), .A2(REG0_REG_24__SCAN_IN), .ZN(n3711) );
  OAI211_X1 U4251 ( .C1(n3713), .C2(n2923), .A(n3712), .B(n3711), .ZN(n3714)
         );
  INV_X1 U4252 ( .A(n3714), .ZN(n3715) );
  NAND2_X1 U4253 ( .A1(n3794), .A2(DATAI_24_), .ZN(n4891) );
  NAND2_X1 U4254 ( .A1(n4909), .A2(n4891), .ZN(n4402) );
  INV_X1 U4255 ( .A(n4402), .ZN(n3833) );
  NOR2_X1 U4256 ( .A1(n4405), .A2(n3833), .ZN(n3900) );
  XNOR2_X1 U4257 ( .A(n3745), .B(REG3_REG_21__SCAN_IN), .ZN(n4946) );
  NAND2_X1 U4258 ( .A1(n4946), .A2(n3109), .ZN(n3722) );
  INV_X1 U4259 ( .A(REG1_REG_21__SCAN_IN), .ZN(n3719) );
  NAND2_X1 U4260 ( .A1(n2494), .A2(REG2_REG_21__SCAN_IN), .ZN(n3718) );
  NAND2_X1 U4261 ( .A1(n3057), .A2(REG0_REG_21__SCAN_IN), .ZN(n3717) );
  OAI211_X1 U4262 ( .C1(n3719), .C2(n2923), .A(n3718), .B(n3717), .ZN(n3720)
         );
  INV_X1 U4263 ( .A(n3720), .ZN(n3721) );
  NAND2_X1 U4264 ( .A1(n3794), .A2(DATAI_21_), .ZN(n4944) );
  INV_X1 U4265 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4173) );
  INV_X1 U4266 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4204) );
  OAI21_X1 U4267 ( .B1(n3745), .B2(n4173), .A(n4204), .ZN(n3723) );
  NAND2_X1 U4268 ( .A1(n3723), .A2(n3731), .ZN(n4922) );
  INV_X1 U4269 ( .A(REG1_REG_22__SCAN_IN), .ZN(n3726) );
  NAND2_X1 U4270 ( .A1(n2494), .A2(REG2_REG_22__SCAN_IN), .ZN(n3725) );
  NAND2_X1 U4271 ( .A1(n3057), .A2(REG0_REG_22__SCAN_IN), .ZN(n3724) );
  OAI211_X1 U4272 ( .C1(n3726), .C2(n2923), .A(n3725), .B(n3724), .ZN(n3727)
         );
  INV_X1 U4273 ( .A(n3727), .ZN(n3728) );
  NAND2_X1 U4274 ( .A1(n3794), .A2(DATAI_22_), .ZN(n4384) );
  AND2_X1 U4275 ( .A1(n4373), .A2(n4384), .ZN(n3811) );
  NAND2_X1 U4276 ( .A1(n3731), .A2(n3730), .ZN(n3732) );
  NAND2_X1 U4277 ( .A1(n3733), .A2(n3732), .ZN(n4913) );
  INV_X1 U4278 ( .A(REG1_REG_23__SCAN_IN), .ZN(n3736) );
  NAND2_X1 U4279 ( .A1(n2494), .A2(REG2_REG_23__SCAN_IN), .ZN(n3735) );
  NAND2_X1 U4280 ( .A1(n3057), .A2(REG0_REG_23__SCAN_IN), .ZN(n3734) );
  OAI211_X1 U4281 ( .C1(n3736), .C2(n2923), .A(n3735), .B(n3734), .ZN(n3737)
         );
  INV_X1 U4282 ( .A(n3737), .ZN(n3738) );
  INV_X1 U4283 ( .A(n4930), .ZN(n4881) );
  NAND2_X1 U4284 ( .A1(n3794), .A2(DATAI_23_), .ZN(n4912) );
  INV_X1 U4285 ( .A(n4912), .ZN(n4375) );
  NOR2_X1 U4286 ( .A1(n4881), .A2(n4375), .ZN(n3834) );
  AOI211_X1 U4287 ( .C1(n4901), .C2(n4903), .A(n3811), .B(n3834), .ZN(n3740)
         );
  INV_X1 U4288 ( .A(n3740), .ZN(n4399) );
  INV_X1 U4289 ( .A(REG1_REG_20__SCAN_IN), .ZN(n3743) );
  NAND2_X1 U4290 ( .A1(n3057), .A2(REG0_REG_20__SCAN_IN), .ZN(n3742) );
  NAND2_X1 U4291 ( .A1(n2494), .A2(REG2_REG_20__SCAN_IN), .ZN(n3741) );
  OAI211_X1 U4292 ( .C1(n2923), .C2(n3743), .A(n3742), .B(n3741), .ZN(n3747)
         );
  NAND2_X1 U4293 ( .A1(n3751), .A2(n4195), .ZN(n3744) );
  NAND2_X1 U4294 ( .A1(n3745), .A2(n3744), .ZN(n4966) );
  NOR2_X1 U4295 ( .A1(n4966), .A2(n3790), .ZN(n3746) );
  NAND2_X1 U4296 ( .A1(n3794), .A2(DATAI_20_), .ZN(n4964) );
  NAND2_X1 U4297 ( .A1(n4982), .A2(n4964), .ZN(n4397) );
  MUX2_X1 U4298 ( .A(n5071), .B(DATAI_18_), .S(n3794), .Z(n4370) );
  NAND2_X1 U4299 ( .A1(n4973), .A2(n4370), .ZN(n4974) );
  NAND2_X1 U4300 ( .A1(n4974), .A2(n3951), .ZN(n3757) );
  INV_X1 U4301 ( .A(n4370), .ZN(n4015) );
  NAND2_X1 U4302 ( .A1(n4371), .A2(n4015), .ZN(n4976) );
  NAND2_X1 U4303 ( .A1(n2494), .A2(REG2_REG_19__SCAN_IN), .ZN(n3755) );
  INV_X1 U4304 ( .A(REG3_REG_19__SCAN_IN), .ZN(n3748) );
  NAND2_X1 U4305 ( .A1(n3749), .A2(n3748), .ZN(n3750) );
  AND2_X1 U4306 ( .A1(n3751), .A2(n3750), .ZN(n4990) );
  NAND2_X1 U4307 ( .A1(n4990), .A2(n3109), .ZN(n3754) );
  NAND2_X1 U4308 ( .A1(n3056), .A2(REG1_REG_19__SCAN_IN), .ZN(n3753) );
  NAND2_X1 U4309 ( .A1(n3057), .A2(REG0_REG_19__SCAN_IN), .ZN(n3752) );
  NAND4_X1 U4310 ( .A1(n3755), .A2(n3754), .A3(n3753), .A4(n3752), .ZN(n4958)
         );
  MUX2_X1 U4311 ( .A(n5130), .B(DATAI_19_), .S(n3794), .Z(n4372) );
  NAND2_X1 U4312 ( .A1(n4958), .A2(n4988), .ZN(n3756) );
  AND2_X1 U4313 ( .A1(n4976), .A2(n3756), .ZN(n3768) );
  NAND2_X1 U4314 ( .A1(n3757), .A2(n3768), .ZN(n3759) );
  INV_X1 U4315 ( .A(n4958), .ZN(n4194) );
  NAND2_X1 U4316 ( .A1(n4194), .A2(n4372), .ZN(n3758) );
  NAND2_X1 U4317 ( .A1(n3759), .A2(n3758), .ZN(n4392) );
  NOR2_X1 U4318 ( .A1(n4982), .A2(n4964), .ZN(n4396) );
  NAND2_X1 U4319 ( .A1(n4903), .A2(n4902), .ZN(n4398) );
  AOI211_X1 U4320 ( .C1(n4397), .C2(n4392), .A(n4396), .B(n4398), .ZN(n3896)
         );
  NAND2_X1 U4321 ( .A1(n5283), .A2(n3966), .ZN(n3763) );
  AND2_X1 U4322 ( .A1(n3760), .A2(n3763), .ZN(n3886) );
  INV_X1 U4323 ( .A(n3761), .ZN(n3762) );
  NAND2_X1 U4324 ( .A1(n3763), .A2(n3762), .ZN(n3764) );
  NAND2_X1 U4325 ( .A1(n3764), .A2(n2535), .ZN(n3892) );
  AOI21_X1 U4326 ( .B1(n3765), .B2(n3886), .A(n3892), .ZN(n3769) );
  AND3_X1 U4327 ( .A1(n3768), .A2(n3767), .A3(n3766), .ZN(n4391) );
  OAI211_X1 U4328 ( .C1(n3769), .C2(n3894), .A(n4391), .B(n4397), .ZN(n3770)
         );
  NOR2_X1 U4329 ( .A1(n4909), .A2(n4891), .ZN(n3832) );
  NOR2_X1 U4330 ( .A1(n4930), .A2(n4912), .ZN(n4882) );
  NOR2_X1 U4331 ( .A1(n3832), .A2(n4882), .ZN(n4401) );
  OAI221_X1 U4332 ( .B1(n4399), .B2(n3896), .C1(n4399), .C2(n3770), .A(n4401), 
        .ZN(n3796) );
  INV_X1 U4333 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4725) );
  INV_X1 U4334 ( .A(n3781), .ZN(n3771) );
  NAND2_X1 U4335 ( .A1(n3771), .A2(REG3_REG_28__SCAN_IN), .ZN(n4388) );
  NAND2_X1 U4336 ( .A1(n3781), .A2(n4734), .ZN(n3772) );
  NAND2_X1 U4337 ( .A1(n4388), .A2(n3772), .ZN(n4434) );
  INV_X1 U4338 ( .A(REG1_REG_28__SCAN_IN), .ZN(n3775) );
  NAND2_X1 U4339 ( .A1(n2494), .A2(REG2_REG_28__SCAN_IN), .ZN(n3774) );
  NAND2_X1 U4340 ( .A1(n3057), .A2(REG0_REG_28__SCAN_IN), .ZN(n3773) );
  OAI211_X1 U4341 ( .C1(n3775), .C2(n2923), .A(n3774), .B(n3773), .ZN(n3776)
         );
  INV_X1 U4342 ( .A(n3776), .ZN(n3777) );
  NAND2_X1 U4343 ( .A1(n3794), .A2(DATAI_28_), .ZN(n4422) );
  INV_X1 U4344 ( .A(n4422), .ZN(n4431) );
  NAND2_X1 U4345 ( .A1(n3779), .A2(n4725), .ZN(n3780) );
  NAND2_X1 U4346 ( .A1(n4451), .A2(n3109), .ZN(n3787) );
  INV_X1 U4347 ( .A(REG1_REG_27__SCAN_IN), .ZN(n3784) );
  NAND2_X1 U4348 ( .A1(n2494), .A2(REG2_REG_27__SCAN_IN), .ZN(n3783) );
  NAND2_X1 U4349 ( .A1(n3057), .A2(REG0_REG_27__SCAN_IN), .ZN(n3782) );
  OAI211_X1 U4350 ( .C1(n3784), .C2(n2923), .A(n3783), .B(n3782), .ZN(n3785)
         );
  INV_X1 U4351 ( .A(n3785), .ZN(n3786) );
  NAND2_X1 U4352 ( .A1(n3794), .A2(DATAI_27_), .ZN(n4450) );
  NOR2_X1 U4353 ( .A1(n4464), .A2(n4450), .ZN(n4407) );
  OR2_X1 U4354 ( .A1(n4408), .A2(n4407), .ZN(n3799) );
  AOI22_X1 U4355 ( .A1(n3056), .A2(REG1_REG_29__SCAN_IN), .B1(n3057), .B2(
        REG0_REG_29__SCAN_IN), .ZN(n3789) );
  NAND2_X1 U4356 ( .A1(n2494), .A2(REG2_REG_29__SCAN_IN), .ZN(n3788) );
  OAI211_X1 U4357 ( .C1(n4388), .C2(n3790), .A(n3789), .B(n3788), .ZN(n4430)
         );
  NAND2_X1 U4358 ( .A1(n3794), .A2(DATAI_29_), .ZN(n4413) );
  NAND2_X1 U4359 ( .A1(n3794), .A2(DATAI_30_), .ZN(n5329) );
  INV_X1 U4360 ( .A(n5329), .ZN(n5317) );
  NAND2_X1 U4361 ( .A1(n4414), .A2(n5317), .ZN(n3795) );
  NAND2_X1 U4362 ( .A1(n3056), .A2(REG1_REG_31__SCAN_IN), .ZN(n3793) );
  NAND2_X1 U4363 ( .A1(n2494), .A2(REG2_REG_31__SCAN_IN), .ZN(n3792) );
  NAND2_X1 U4364 ( .A1(n3057), .A2(REG0_REG_31__SCAN_IN), .ZN(n3791) );
  NAND3_X1 U4365 ( .A1(n3793), .A2(n3792), .A3(n3791), .ZN(n5314) );
  AND2_X1 U4366 ( .A1(n3794), .A2(DATAI_31_), .ZN(n5326) );
  INV_X1 U4367 ( .A(n5326), .ZN(n5331) );
  NAND2_X1 U4368 ( .A1(n5314), .A2(n5331), .ZN(n3902) );
  AND2_X1 U4369 ( .A1(n3795), .A2(n3902), .ZN(n3824) );
  OAI21_X1 U4370 ( .B1(n4430), .B2(n4413), .A(n3824), .ZN(n3798) );
  AOI211_X1 U4371 ( .C1(n3900), .C2(n3796), .A(n3799), .B(n3798), .ZN(n3801)
         );
  NAND2_X1 U4372 ( .A1(n4448), .A2(n4422), .ZN(n3807) );
  INV_X1 U4373 ( .A(n3807), .ZN(n3797) );
  AOI21_X1 U4374 ( .B1(n4430), .B2(n4413), .A(n3797), .ZN(n3800) );
  AOI21_X1 U4375 ( .B1(n3800), .B2(n3799), .A(n3798), .ZN(n3904) );
  NAND2_X1 U4376 ( .A1(n4464), .A2(n4450), .ZN(n3849) );
  NAND2_X1 U4377 ( .A1(n4481), .A2(n4467), .ZN(n4406) );
  NAND3_X1 U4378 ( .A1(n3849), .A2(n4406), .A3(n3800), .ZN(n3897) );
  AOI22_X1 U4379 ( .A1(n3854), .A2(n3801), .B1(n3904), .B2(n3897), .ZN(n3803)
         );
  NOR2_X1 U4380 ( .A1(n5314), .A2(n5329), .ZN(n3802) );
  OAI21_X1 U4381 ( .B1(n3803), .B2(n3802), .A(n3858), .ZN(n3806) );
  INV_X1 U4382 ( .A(n5314), .ZN(n3804) );
  NAND2_X1 U4383 ( .A1(n3804), .A2(n5326), .ZN(n3805) );
  OAI21_X1 U4384 ( .B1(n4414), .B2(n5317), .A(n3805), .ZN(n3903) );
  AOI22_X1 U4385 ( .A1(n3806), .A2(n3907), .B1(n5326), .B2(n3903), .ZN(n3909)
         );
  INV_X1 U4386 ( .A(n4408), .ZN(n3808) );
  NAND2_X1 U4387 ( .A1(n3808), .A2(n3807), .ZN(n4425) );
  NAND2_X1 U4388 ( .A1(n4404), .A2(n3810), .ZN(n4477) );
  INV_X1 U4389 ( .A(n3811), .ZN(n3812) );
  NAND2_X1 U4390 ( .A1(n4903), .A2(n3812), .ZN(n4919) );
  INV_X1 U4391 ( .A(n4397), .ZN(n3813) );
  INV_X1 U4392 ( .A(n3079), .ZN(n5123) );
  NAND2_X1 U4393 ( .A1(n4236), .A2(n5123), .ZN(n3857) );
  NAND2_X1 U4394 ( .A1(n3855), .A2(n3857), .ZN(n5135) );
  NOR4_X1 U4395 ( .A1(n4919), .A2(n4955), .A3(n5290), .A4(n5135), .ZN(n3818)
         );
  INV_X1 U4396 ( .A(n4901), .ZN(n3814) );
  NAND2_X1 U4397 ( .A1(n4902), .A2(n3814), .ZN(n4936) );
  INV_X1 U4398 ( .A(n4936), .ZN(n3817) );
  NAND4_X1 U4399 ( .A1(n3818), .A2(n3817), .A3(n3816), .A4(n3815), .ZN(n3848)
         );
  NAND4_X1 U4400 ( .A1(n3822), .A2(n3821), .A3(n3820), .A4(n3819), .ZN(n3827)
         );
  NAND2_X1 U4401 ( .A1(n4974), .A2(n4976), .ZN(n4368) );
  INV_X1 U4402 ( .A(n3903), .ZN(n3825) );
  NAND4_X1 U4403 ( .A1(n2669), .A2(n3825), .A3(n3824), .A4(n3823), .ZN(n3826)
         );
  NOR2_X1 U4404 ( .A1(n3827), .A2(n3826), .ZN(n3831) );
  XNOR2_X1 U4405 ( .A(n4958), .B(n4988), .ZN(n4984) );
  INV_X1 U4406 ( .A(n3828), .ZN(n3829) );
  NAND4_X1 U4407 ( .A1(n3831), .A2(n2672), .A3(n3830), .A4(n3829), .ZN(n3847)
         );
  OR2_X1 U4408 ( .A1(n3833), .A2(n3832), .ZN(n4885) );
  INV_X1 U4409 ( .A(n4882), .ZN(n3836) );
  INV_X1 U4410 ( .A(n3834), .ZN(n3835) );
  NAND2_X1 U4411 ( .A1(n3836), .A2(n3835), .ZN(n4904) );
  NAND4_X1 U4412 ( .A1(n3839), .A2(n3838), .A3(n3138), .A4(n3837), .ZN(n3845)
         );
  NAND4_X1 U4413 ( .A1(n3843), .A2(n3842), .A3(n3841), .A4(n3840), .ZN(n3844)
         );
  OR4_X1 U4414 ( .A1(n4885), .A2(n4904), .A3(n3845), .A4(n3844), .ZN(n3846) );
  NOR4_X1 U4415 ( .A1(n4477), .A2(n3848), .A3(n3847), .A4(n3846), .ZN(n3852)
         );
  INV_X1 U4416 ( .A(n3849), .ZN(n3850) );
  INV_X1 U4417 ( .A(n4443), .ZN(n3851) );
  NAND2_X1 U4418 ( .A1(n3852), .A2(n3851), .ZN(n3853) );
  XNOR2_X1 U4419 ( .A(n4430), .B(n4413), .ZN(n4409) );
  XNOR2_X1 U4420 ( .A(n4481), .B(n4467), .ZN(n4459) );
  NOR4_X1 U4421 ( .A1(n4425), .A2(n3853), .A3(n4409), .A4(n4459), .ZN(n3908)
         );
  INV_X1 U4422 ( .A(n3854), .ZN(n3901) );
  OAI211_X1 U4423 ( .C1(n2567), .C2(n3858), .A(n3857), .B(n3856), .ZN(n3861)
         );
  NAND3_X1 U4424 ( .A1(n3861), .A2(n3860), .A3(n3859), .ZN(n3864) );
  NAND3_X1 U4425 ( .A1(n3864), .A2(n3863), .A3(n3862), .ZN(n3867) );
  NAND3_X1 U4426 ( .A1(n3867), .A2(n3866), .A3(n3865), .ZN(n3869) );
  NAND4_X1 U4427 ( .A1(n3870), .A2(n3869), .A3(n3874), .A4(n3868), .ZN(n3879)
         );
  INV_X1 U4428 ( .A(n3871), .ZN(n3875) );
  OAI21_X1 U4429 ( .B1(n4138), .B2(n4231), .A(n3872), .ZN(n3873) );
  AOI21_X1 U4430 ( .B1(n3875), .B2(n3874), .A(n3873), .ZN(n3878) );
  INV_X1 U4431 ( .A(n3876), .ZN(n3877) );
  AOI211_X1 U4432 ( .C1(n3879), .C2(n3878), .A(n3877), .B(n2533), .ZN(n3883)
         );
  INV_X1 U4433 ( .A(n3880), .ZN(n3882) );
  OAI21_X1 U4434 ( .B1(n3883), .B2(n3882), .A(n3881), .ZN(n3885) );
  OAI211_X1 U4435 ( .C1(n2581), .C2(n4229), .A(n3885), .B(n3884), .ZN(n3890)
         );
  INV_X1 U4436 ( .A(n3886), .ZN(n3887) );
  AOI211_X1 U4437 ( .C1(n3890), .C2(n3889), .A(n3888), .B(n3887), .ZN(n3891)
         );
  NOR2_X1 U4438 ( .A1(n3892), .A2(n3891), .ZN(n3893) );
  OAI211_X1 U4439 ( .C1(n3894), .C2(n3893), .A(n4391), .B(n4397), .ZN(n3895)
         );
  OAI221_X1 U4440 ( .B1(n4399), .B2(n3896), .C1(n4399), .C2(n3895), .A(n4401), 
        .ZN(n3899) );
  INV_X1 U4441 ( .A(n3897), .ZN(n3898) );
  OAI221_X1 U4442 ( .B1(n3901), .B2(n3900), .C1(n3901), .C2(n3899), .A(n3898), 
        .ZN(n3905) );
  AOI22_X1 U4443 ( .A1(n3905), .A2(n3904), .B1(n3903), .B2(n3902), .ZN(n3906)
         );
  OAI22_X1 U4444 ( .A1(n3909), .A2(n3908), .B1(n3907), .B2(n3906), .ZN(n3910)
         );
  XNOR2_X1 U4445 ( .A(n3910), .B(n2961), .ZN(n3917) );
  INV_X1 U4446 ( .A(n3911), .ZN(n3912) );
  NAND2_X1 U4447 ( .A1(n3913), .A2(n3912), .ZN(n3914) );
  OAI211_X1 U4448 ( .C1(n4997), .C2(n3916), .A(n3914), .B(B_REG_SCAN_IN), .ZN(
        n3915) );
  OAI21_X1 U4449 ( .B1(n3917), .B2(n3916), .A(n3915), .ZN(U3239) );
  NAND2_X1 U4450 ( .A1(n4224), .A2(n3492), .ZN(n3919) );
  NAND2_X1 U4451 ( .A1(n3921), .A2(n4050), .ZN(n3918) );
  NAND2_X1 U4452 ( .A1(n3919), .A2(n3918), .ZN(n3920) );
  XNOR2_X1 U4453 ( .A(n3920), .B(n3490), .ZN(n3923) );
  AND2_X1 U4454 ( .A1(n3921), .A2(n3492), .ZN(n3922) );
  AOI21_X1 U4455 ( .B1(n4224), .B2(n3026), .A(n3922), .ZN(n3924) );
  NAND2_X1 U4456 ( .A1(n3923), .A2(n3924), .ZN(n3965) );
  INV_X1 U4457 ( .A(n3923), .ZN(n3926) );
  INV_X1 U4458 ( .A(n3924), .ZN(n3925) );
  NAND2_X1 U4459 ( .A1(n3926), .A2(n3925), .ZN(n3927) );
  NOR2_X1 U4460 ( .A1(n3930), .A2(n2618), .ZN(n3931) );
  AOI21_X1 U4461 ( .B1(n3931), .B2(n3929), .A(n2521), .ZN(n3937) );
  AOI22_X1 U4462 ( .A1(n4219), .A2(n5267), .B1(n4183), .B2(n3932), .ZN(n3936)
         );
  NOR2_X1 U4463 ( .A1(STATE_REG_SCAN_IN), .A2(n4726), .ZN(n4312) );
  NOR2_X1 U4464 ( .A1(n4214), .A2(n3933), .ZN(n3934) );
  AOI211_X1 U4465 ( .C1(n5268), .C2(n4225), .A(n4312), .B(n3934), .ZN(n3935)
         );
  OAI211_X1 U4466 ( .C1(n3937), .C2(n5271), .A(n3936), .B(n3935), .ZN(U3212)
         );
  AOI211_X1 U4467 ( .C1(n3940), .C2(n3939), .A(n3938), .B(n5108), .ZN(n3948)
         );
  OAI211_X1 U4468 ( .C1(n3943), .C2(n3942), .A(n5116), .B(n3941), .ZN(n3946)
         );
  AOI21_X1 U4469 ( .B1(n5107), .B2(ADDR_REG_13__SCAN_IN), .A(n3944), .ZN(n3945) );
  OAI211_X1 U4470 ( .C1(n4348), .C2(n5240), .A(n3946), .B(n3945), .ZN(n3947)
         );
  OR2_X1 U4471 ( .A1(n3948), .A2(n3947), .ZN(U3253) );
  NAND2_X1 U4472 ( .A1(n3950), .A2(n3949), .ZN(n4369) );
  XNOR2_X1 U4473 ( .A(n4369), .B(n2669), .ZN(n5044) );
  NAND2_X1 U4474 ( .A1(n3952), .A2(n3951), .ZN(n4977) );
  XNOR2_X1 U4475 ( .A(n4977), .B(n2669), .ZN(n3955) );
  AOI22_X1 U4476 ( .A1(n5285), .A2(n4957), .B1(n4370), .B2(n5325), .ZN(n3953)
         );
  OAI21_X1 U4477 ( .B1(n4194), .B2(n5127), .A(n3953), .ZN(n3954) );
  AOI21_X1 U4478 ( .B1(n3955), .B2(n5124), .A(n3954), .ZN(n5043) );
  INV_X1 U4479 ( .A(n5043), .ZN(n3961) );
  INV_X1 U4480 ( .A(n4989), .ZN(n3958) );
  AOI21_X1 U4481 ( .B1(n3956), .B2(n4370), .A(n5296), .ZN(n3957) );
  NAND2_X1 U4482 ( .A1(n3958), .A2(n3957), .ZN(n5042) );
  AOI22_X1 U4483 ( .A1(n5333), .A2(REG2_REG_18__SCAN_IN), .B1(n4013), .B2(
        n5303), .ZN(n3959) );
  OAI21_X1 U4484 ( .B1(n5042), .B2(n4969), .A(n3959), .ZN(n3960) );
  AOI21_X1 U4485 ( .B1(n3961), .B2(n5138), .A(n3960), .ZN(n3962) );
  OAI21_X1 U4486 ( .B1(n5044), .B2(n5307), .A(n3962), .ZN(U3272) );
  NAND2_X1 U4487 ( .A1(n5267), .A2(n3026), .ZN(n3964) );
  NAND2_X1 U4488 ( .A1(n3966), .A2(n3492), .ZN(n3963) );
  NAND2_X1 U4489 ( .A1(n3964), .A2(n3963), .ZN(n3983) );
  NAND2_X1 U4490 ( .A1(n5267), .A2(n3492), .ZN(n3968) );
  NAND2_X1 U4491 ( .A1(n3966), .A2(n4050), .ZN(n3967) );
  NAND2_X1 U4492 ( .A1(n3968), .A2(n3967), .ZN(n3969) );
  NAND2_X1 U4493 ( .A1(n3985), .A2(n3984), .ZN(n3972) );
  XOR2_X1 U4494 ( .A(n3983), .B(n3972), .Z(n3978) );
  AOI22_X1 U4495 ( .A1(n4219), .A2(n4223), .B1(n4183), .B2(n3973), .ZN(n3977)
         );
  AND2_X1 U4496 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4325) );
  NOR2_X1 U4497 ( .A1(n4214), .A2(n3974), .ZN(n3975) );
  AOI211_X1 U4498 ( .C1(n5268), .C2(n4224), .A(n4325), .B(n3975), .ZN(n3976)
         );
  OAI211_X1 U4499 ( .C1(n3978), .C2(n5271), .A(n3977), .B(n3976), .ZN(U3238)
         );
  NAND2_X1 U4500 ( .A1(n5285), .A2(n3492), .ZN(n3980) );
  NAND2_X1 U4501 ( .A1(n3998), .A2(n4050), .ZN(n3979) );
  NAND2_X1 U4502 ( .A1(n3980), .A2(n3979), .ZN(n3981) );
  XNOR2_X1 U4503 ( .A(n3981), .B(n3024), .ZN(n4003) );
  AND2_X1 U4504 ( .A1(n3998), .A2(n3492), .ZN(n3982) );
  AOI21_X1 U4505 ( .B1(n5285), .B2(n3026), .A(n3982), .ZN(n4004) );
  XNOR2_X1 U4506 ( .A(n4003), .B(n4004), .ZN(n4001) );
  NAND2_X1 U4507 ( .A1(n3984), .A2(n3983), .ZN(n3986) );
  NAND2_X1 U4508 ( .A1(n4223), .A2(n3492), .ZN(n3988) );
  NAND2_X1 U4509 ( .A1(n5265), .A2(n4050), .ZN(n3987) );
  NAND2_X1 U4510 ( .A1(n3988), .A2(n3987), .ZN(n3989) );
  XNOR2_X1 U4511 ( .A(n3989), .B(n3490), .ZN(n3993) );
  AND2_X1 U4512 ( .A1(n5265), .A2(n3492), .ZN(n3990) );
  AOI21_X1 U4513 ( .B1(n4223), .B2(n3026), .A(n3990), .ZN(n3992) );
  XNOR2_X1 U4514 ( .A(n3993), .B(n3992), .ZN(n5270) );
  NAND2_X1 U4515 ( .A1(n3993), .A2(n3992), .ZN(n3994) );
  XOR2_X1 U4516 ( .A(n4001), .B(n4002), .Z(n4000) );
  NAND2_X1 U4517 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4346) );
  OAI21_X1 U4518 ( .B1(n4216), .B2(n2716), .A(n4346), .ZN(n3997) );
  OAI22_X1 U4519 ( .A1(n4205), .A2(n4973), .B1(n5280), .B2(n3995), .ZN(n3996)
         );
  AOI211_X1 U4520 ( .C1(n3998), .C2(n5266), .A(n3997), .B(n3996), .ZN(n3999)
         );
  OAI21_X1 U4521 ( .B1(n4000), .B2(n5271), .A(n3999), .ZN(U3225) );
  NAND2_X1 U4522 ( .A1(n4002), .A2(n4001), .ZN(n4007) );
  INV_X1 U4523 ( .A(n4003), .ZN(n4005) );
  NAND2_X1 U4524 ( .A1(n4005), .A2(n4004), .ZN(n4006) );
  NAND2_X1 U4525 ( .A1(n4371), .A2(n3492), .ZN(n4009) );
  NAND2_X1 U4526 ( .A1(n4370), .A2(n4050), .ZN(n4008) );
  NAND2_X1 U4527 ( .A1(n4009), .A2(n4008), .ZN(n4010) );
  XNOR2_X1 U4528 ( .A(n4010), .B(n3490), .ZN(n4033) );
  AND2_X1 U4529 ( .A1(n4370), .A2(n3492), .ZN(n4011) );
  AOI21_X1 U4530 ( .B1(n4371), .B2(n3026), .A(n4011), .ZN(n4034) );
  XNOR2_X1 U4531 ( .A(n4033), .B(n4034), .ZN(n4012) );
  XNOR2_X1 U4532 ( .A(n4039), .B(n4012), .ZN(n4019) );
  AOI22_X1 U4533 ( .A1(n4219), .A2(n4958), .B1(n4183), .B2(n4013), .ZN(n4018)
         );
  NOR2_X1 U4534 ( .A1(STATE_REG_SCAN_IN), .A2(n4014), .ZN(n4360) );
  NOR2_X1 U4535 ( .A1(n4214), .A2(n4015), .ZN(n4016) );
  AOI211_X1 U4536 ( .C1(n5268), .C2(n5285), .A(n4360), .B(n4016), .ZN(n4017)
         );
  OAI211_X1 U4537 ( .C1(n4019), .C2(n5271), .A(n4018), .B(n4017), .ZN(U3235)
         );
  OAI211_X1 U4538 ( .C1(n4022), .C2(n4020), .A(n4021), .B(n4134), .ZN(n4028)
         );
  OAI22_X1 U4539 ( .A1(n4024), .A2(n4205), .B1(n4216), .B2(n4023), .ZN(n4025)
         );
  AOI21_X1 U4540 ( .B1(REG3_REG_1__SCAN_IN), .B2(n4026), .A(n4025), .ZN(n4027)
         );
  OAI211_X1 U4541 ( .C1(n4214), .C2(n4029), .A(n4028), .B(n4027), .ZN(U3219)
         );
  AOI22_X1 U4542 ( .A1(n5095), .A2(n4622), .B1(n4030), .B2(n2908), .ZN(U3458)
         );
  INV_X1 U4543 ( .A(DATAI_20_), .ZN(n4031) );
  MUX2_X1 U4544 ( .A(n4031), .B(n2997), .S(STATE_REG_SCAN_IN), .Z(n4032) );
  INV_X1 U4545 ( .A(n4032), .ZN(U3332) );
  AND2_X1 U4546 ( .A1(n4033), .A2(n4034), .ZN(n4038) );
  INV_X1 U4547 ( .A(n4033), .ZN(n4036) );
  INV_X1 U4548 ( .A(n4034), .ZN(n4035) );
  NAND2_X1 U4549 ( .A1(n4036), .A2(n4035), .ZN(n4037) );
  NAND2_X1 U4550 ( .A1(n4958), .A2(n3492), .ZN(n4041) );
  NAND2_X1 U4551 ( .A1(n4372), .A2(n4050), .ZN(n4040) );
  NAND2_X1 U4552 ( .A1(n4041), .A2(n4040), .ZN(n4042) );
  XNOR2_X1 U4553 ( .A(n4042), .B(n3490), .ZN(n4044) );
  AND2_X1 U4554 ( .A1(n4372), .A2(n3492), .ZN(n4043) );
  AOI21_X1 U4555 ( .B1(n4958), .B2(n3026), .A(n4043), .ZN(n4045) );
  NAND2_X1 U4556 ( .A1(n4044), .A2(n4045), .ZN(n4049) );
  INV_X1 U4557 ( .A(n4044), .ZN(n4047) );
  INV_X1 U4558 ( .A(n4045), .ZN(n4046) );
  NAND2_X1 U4559 ( .A1(n4047), .A2(n4046), .ZN(n4048) );
  NAND2_X1 U4560 ( .A1(n4049), .A2(n4048), .ZN(n4160) );
  NAND2_X1 U4561 ( .A1(n4982), .A2(n3492), .ZN(n4052) );
  OR2_X1 U4562 ( .A1(n4964), .A2(n4123), .ZN(n4051) );
  NAND2_X1 U4563 ( .A1(n4052), .A2(n4051), .ZN(n4053) );
  XNOR2_X1 U4564 ( .A(n4053), .B(n3490), .ZN(n4058) );
  INV_X1 U4565 ( .A(n4058), .ZN(n4056) );
  NOR2_X1 U4566 ( .A1(n4964), .A2(n4112), .ZN(n4054) );
  AOI21_X1 U4567 ( .B1(n4982), .B2(n3026), .A(n4054), .ZN(n4057) );
  INV_X1 U4568 ( .A(n4057), .ZN(n4055) );
  NAND2_X1 U4569 ( .A1(n4056), .A2(n4055), .ZN(n4190) );
  AND2_X1 U4570 ( .A1(n4058), .A2(n4057), .ZN(n4189) );
  NAND2_X1 U4571 ( .A1(n4222), .A2(n3492), .ZN(n4060) );
  OR2_X1 U4572 ( .A1(n4944), .A2(n4123), .ZN(n4059) );
  NAND2_X1 U4573 ( .A1(n4060), .A2(n4059), .ZN(n4061) );
  XNOR2_X1 U4574 ( .A(n4061), .B(n3490), .ZN(n4063) );
  NOR2_X1 U4575 ( .A1(n4944), .A2(n4112), .ZN(n4062) );
  AOI21_X1 U4576 ( .B1(n4222), .B2(n3026), .A(n4062), .ZN(n4064) );
  NAND2_X1 U4577 ( .A1(n4063), .A2(n4064), .ZN(n4167) );
  NAND2_X1 U4578 ( .A1(n4166), .A2(n4167), .ZN(n4171) );
  INV_X1 U4579 ( .A(n4063), .ZN(n4066) );
  INV_X1 U4580 ( .A(n4064), .ZN(n4065) );
  NAND2_X1 U4581 ( .A1(n4066), .A2(n4065), .ZN(n4169) );
  NAND2_X1 U4582 ( .A1(n4171), .A2(n4169), .ZN(n4202) );
  INV_X1 U4583 ( .A(n4202), .ZN(n4072) );
  NAND2_X1 U4584 ( .A1(n4373), .A2(n3492), .ZN(n4068) );
  OR2_X1 U4585 ( .A1(n4384), .A2(n4123), .ZN(n4067) );
  NAND2_X1 U4586 ( .A1(n4068), .A2(n4067), .ZN(n4069) );
  XNOR2_X1 U4587 ( .A(n4069), .B(n3490), .ZN(n4074) );
  NOR2_X1 U4588 ( .A1(n4384), .A2(n4112), .ZN(n4070) );
  AOI21_X1 U4589 ( .B1(n4373), .B2(n3026), .A(n4070), .ZN(n4073) );
  XNOR2_X1 U4590 ( .A(n4074), .B(n4073), .ZN(n4203) );
  NAND2_X1 U4591 ( .A1(n4074), .A2(n4073), .ZN(n4075) );
  NAND2_X1 U4592 ( .A1(n4930), .A2(n3492), .ZN(n4077) );
  OR2_X1 U4593 ( .A1(n4912), .A2(n4123), .ZN(n4076) );
  NAND2_X1 U4594 ( .A1(n4077), .A2(n4076), .ZN(n4078) );
  XNOR2_X1 U4595 ( .A(n4078), .B(n3490), .ZN(n4081) );
  NOR2_X1 U4596 ( .A1(n4912), .A2(n4112), .ZN(n4079) );
  AOI21_X1 U4597 ( .B1(n4930), .B2(n3026), .A(n4079), .ZN(n4082) );
  XNOR2_X1 U4598 ( .A(n4081), .B(n4082), .ZN(n4154) );
  INV_X1 U4599 ( .A(n4081), .ZN(n4084) );
  INV_X1 U4600 ( .A(n4082), .ZN(n4083) );
  NAND2_X1 U4601 ( .A1(n4084), .A2(n4083), .ZN(n4085) );
  NAND2_X2 U4602 ( .A1(n4151), .A2(n4085), .ZN(n4108) );
  INV_X1 U4603 ( .A(n4108), .ZN(n4089) );
  NAND2_X1 U4604 ( .A1(n4909), .A2(n3492), .ZN(n4087) );
  OR2_X1 U4605 ( .A1(n4891), .A2(n4123), .ZN(n4086) );
  NAND2_X1 U4606 ( .A1(n4087), .A2(n4086), .ZN(n4088) );
  XNOR2_X1 U4607 ( .A(n4088), .B(n3490), .ZN(n4099) );
  NOR2_X1 U4608 ( .A1(n4891), .A2(n4112), .ZN(n4090) );
  AOI21_X1 U4609 ( .B1(n4909), .B2(n3026), .A(n4090), .ZN(n4098) );
  INV_X1 U4610 ( .A(n4098), .ZN(n4181) );
  INV_X1 U4611 ( .A(n4099), .ZN(n4100) );
  NOR2_X1 U4612 ( .A1(n4478), .A2(n4112), .ZN(n4091) );
  AOI21_X1 U4613 ( .B1(n4889), .B2(n3026), .A(n4091), .ZN(n4103) );
  OAI22_X1 U4614 ( .A1(n4458), .A2(n4112), .B1(n4123), .B2(n4478), .ZN(n4092)
         );
  XOR2_X1 U4615 ( .A(n3024), .B(n4092), .Z(n4101) );
  XOR2_X1 U4616 ( .A(n4103), .B(n4101), .Z(n4093) );
  INV_X1 U4617 ( .A(n4094), .ZN(n4486) );
  OAI22_X1 U4618 ( .A1(n4479), .A2(n4216), .B1(STATE_REG_SCAN_IN), .B2(n4741), 
        .ZN(n4095) );
  AOI21_X1 U4619 ( .B1(n4486), .B2(n4183), .A(n4095), .ZN(n4097) );
  AOI22_X1 U4620 ( .A1(n4481), .A2(n5276), .B1(n4485), .B2(n5266), .ZN(n4096)
         );
  OAI22_X1 U4621 ( .A1(n4101), .A2(n4103), .B1(n4098), .B2(n4099), .ZN(n4107)
         );
  NOR2_X1 U4622 ( .A1(n4100), .A2(n4181), .ZN(n4102) );
  OAI21_X1 U4623 ( .B1(n4103), .B2(n4102), .A(n4101), .ZN(n4104) );
  NAND2_X1 U4624 ( .A1(n4481), .A2(n3492), .ZN(n4110) );
  OR2_X1 U4625 ( .A1(n4467), .A2(n4123), .ZN(n4109) );
  NAND2_X1 U4626 ( .A1(n4110), .A2(n4109), .ZN(n4111) );
  XNOR2_X1 U4627 ( .A(n4111), .B(n3024), .ZN(n4211) );
  NAND2_X1 U4628 ( .A1(n4481), .A2(n3026), .ZN(n4114) );
  OR2_X1 U4629 ( .A1(n4112), .A2(n4467), .ZN(n4113) );
  NAND2_X1 U4630 ( .A1(n4114), .A2(n4113), .ZN(n4210) );
  NOR2_X1 U4631 ( .A1(n4211), .A2(n4210), .ZN(n4117) );
  INV_X1 U4632 ( .A(n4211), .ZN(n4116) );
  INV_X1 U4633 ( .A(n4210), .ZN(n4115) );
  OAI22_X2 U4634 ( .A1(n4213), .A2(n4117), .B1(n4116), .B2(n4115), .ZN(n4145)
         );
  INV_X1 U4635 ( .A(n4464), .ZN(n4423) );
  OAI22_X1 U4636 ( .A1(n4423), .A2(n3324), .B1(n4112), .B2(n4450), .ZN(n4121)
         );
  NAND2_X1 U4637 ( .A1(n4464), .A2(n3492), .ZN(n4119) );
  OR2_X1 U4638 ( .A1(n4450), .A2(n4123), .ZN(n4118) );
  NAND2_X1 U4639 ( .A1(n4119), .A2(n4118), .ZN(n4120) );
  XNOR2_X1 U4640 ( .A(n4120), .B(n3024), .ZN(n4122) );
  XOR2_X1 U4641 ( .A(n4121), .B(n4122), .Z(n4144) );
  AOI21_X1 U4642 ( .B1(n4145), .B2(n4144), .A(n2745), .ZN(n4128) );
  OAI22_X1 U4643 ( .A1(n4383), .A2(n4112), .B1(n4123), .B2(n4422), .ZN(n4124)
         );
  XNOR2_X1 U4644 ( .A(n4124), .B(n3024), .ZN(n4126) );
  OAI22_X1 U4645 ( .A1(n4383), .A2(n3324), .B1(n4112), .B2(n4422), .ZN(n4125)
         );
  XNOR2_X1 U4646 ( .A(n4126), .B(n4125), .ZN(n4127) );
  XNOR2_X1 U4647 ( .A(n4128), .B(n4127), .ZN(n4133) );
  NAND2_X1 U4648 ( .A1(n4464), .A2(n5268), .ZN(n4130) );
  AOI22_X1 U4649 ( .A1(n5266), .A2(n4431), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n4129) );
  OAI211_X1 U4650 ( .C1(n4434), .C2(n5280), .A(n4130), .B(n4129), .ZN(n4131)
         );
  AOI21_X1 U4651 ( .B1(n4219), .B2(n4430), .A(n4131), .ZN(n4132) );
  OAI21_X1 U4652 ( .B1(n4133), .B2(n5271), .A(n4132), .ZN(U3217) );
  OAI211_X1 U4653 ( .C1(n3507), .C2(n4136), .A(n4135), .B(n4134), .ZN(n4143)
         );
  AOI22_X1 U4654 ( .A1(n4219), .A2(n4230), .B1(n4183), .B2(n4137), .ZN(n4142)
         );
  NOR2_X1 U4655 ( .A1(n4214), .A2(n4138), .ZN(n4139) );
  AOI211_X1 U4656 ( .C1(n5268), .C2(n4232), .A(n4140), .B(n4139), .ZN(n4141)
         );
  NAND3_X1 U4657 ( .A1(n4143), .A2(n4142), .A3(n4141), .ZN(U3210) );
  XNOR2_X1 U4658 ( .A(n4145), .B(n4144), .ZN(n4150) );
  AOI22_X1 U4659 ( .A1(n4451), .A2(n4183), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n4147) );
  NAND2_X1 U4660 ( .A1(n4481), .A2(n5268), .ZN(n4146) );
  OAI211_X1 U4661 ( .C1(n4214), .C2(n4450), .A(n4147), .B(n4146), .ZN(n4148)
         );
  AOI21_X1 U4662 ( .B1(n4448), .B2(n5276), .A(n4148), .ZN(n4149) );
  OAI21_X1 U4663 ( .B1(n4150), .B2(n5271), .A(n4149), .ZN(U3211) );
  INV_X1 U4664 ( .A(n4151), .ZN(n4152) );
  AOI211_X1 U4665 ( .C1(n4154), .C2(n4153), .A(n5271), .B(n4152), .ZN(n4158)
         );
  OAI22_X1 U4666 ( .A1(n4479), .A2(n4205), .B1(n4913), .B2(n5280), .ZN(n4157)
         );
  AOI22_X1 U4667 ( .A1(n5268), .A2(n4373), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n4155) );
  OAI21_X1 U4668 ( .B1(n4214), .B2(n4912), .A(n4155), .ZN(n4156) );
  OR3_X1 U4669 ( .A1(n4158), .A2(n4157), .A3(n4156), .ZN(U3213) );
  AOI21_X1 U4670 ( .B1(n4160), .B2(n4159), .A(n2522), .ZN(n4165) );
  AOI22_X1 U4671 ( .A1(n4219), .A2(n4982), .B1(n4183), .B2(n4990), .ZN(n4164)
         );
  NOR2_X1 U4672 ( .A1(n4214), .A2(n4988), .ZN(n4161) );
  AOI211_X1 U4673 ( .C1(n5268), .C2(n4371), .A(n4162), .B(n4161), .ZN(n4163)
         );
  OAI211_X1 U4674 ( .C1(n4165), .C2(n5271), .A(n4164), .B(n4163), .ZN(U3216)
         );
  AOI21_X1 U4675 ( .B1(n4169), .B2(n4167), .A(n4166), .ZN(n4168) );
  INV_X1 U4676 ( .A(n4168), .ZN(n4172) );
  INV_X1 U4677 ( .A(n4169), .ZN(n4170) );
  AOI22_X1 U4678 ( .A1(n4172), .A2(n4171), .B1(n4170), .B2(n4166), .ZN(n4177)
         );
  AOI22_X1 U4679 ( .A1(n4946), .A2(n4183), .B1(n5268), .B2(n4982), .ZN(n4176)
         );
  INV_X1 U4680 ( .A(n4944), .ZN(n4938) );
  INV_X1 U4681 ( .A(n4373), .ZN(n4940) );
  OAI22_X1 U4682 ( .A1(n4205), .A2(n4940), .B1(STATE_REG_SCAN_IN), .B2(n4173), 
        .ZN(n4174) );
  AOI21_X1 U4683 ( .B1(n4938), .B2(n5266), .A(n4174), .ZN(n4175) );
  OAI211_X1 U4684 ( .C1(n4177), .C2(n5271), .A(n4176), .B(n4175), .ZN(U3220)
         );
  INV_X1 U4685 ( .A(n4178), .ZN(n4182) );
  OR2_X1 U4686 ( .A1(n4179), .A2(n4178), .ZN(n4180) );
  AOI22_X1 U4687 ( .A1(n2507), .A2(n4182), .B1(n4181), .B2(n4180), .ZN(n4188)
         );
  AOI22_X1 U4688 ( .A1(n4889), .A2(n5276), .B1(n4893), .B2(n4183), .ZN(n4187)
         );
  INV_X1 U4689 ( .A(n4891), .ZN(n4385) );
  OAI22_X1 U4690 ( .A1(n4881), .A2(n4216), .B1(STATE_REG_SCAN_IN), .B2(n4184), 
        .ZN(n4185) );
  AOI21_X1 U4691 ( .B1(n4385), .B2(n5266), .A(n4185), .ZN(n4186) );
  OAI211_X1 U4692 ( .C1(n4188), .C2(n5271), .A(n4187), .B(n4186), .ZN(U3226)
         );
  INV_X1 U4693 ( .A(n4189), .ZN(n4191) );
  NAND2_X1 U4694 ( .A1(n4191), .A2(n4190), .ZN(n4192) );
  XNOR2_X1 U4695 ( .A(n4193), .B(n4192), .ZN(n4199) );
  OAI22_X1 U4696 ( .A1(n4216), .A2(n4194), .B1(n4966), .B2(n5280), .ZN(n4197)
         );
  OAI22_X1 U4697 ( .A1(n4205), .A2(n4960), .B1(STATE_REG_SCAN_IN), .B2(n4195), 
        .ZN(n4196) );
  AOI211_X1 U4698 ( .C1(n4956), .C2(n5266), .A(n4197), .B(n4196), .ZN(n4198)
         );
  OAI21_X1 U4699 ( .B1(n4199), .B2(n5271), .A(n4198), .ZN(U3230) );
  INV_X1 U4700 ( .A(n4200), .ZN(n4201) );
  AOI21_X1 U4701 ( .B1(n4203), .B2(n4202), .A(n4201), .ZN(n4209) );
  INV_X1 U4702 ( .A(n4384), .ZN(n4929) );
  OAI22_X1 U4703 ( .A1(n4216), .A2(n4960), .B1(STATE_REG_SCAN_IN), .B2(n4204), 
        .ZN(n4207) );
  OAI22_X1 U4704 ( .A1(n4881), .A2(n4205), .B1(n5280), .B2(n4922), .ZN(n4206)
         );
  AOI211_X1 U4705 ( .C1(n4929), .C2(n5266), .A(n4207), .B(n4206), .ZN(n4208)
         );
  OAI21_X1 U4706 ( .B1(n4209), .B2(n5271), .A(n4208), .ZN(U3232) );
  XNOR2_X1 U4707 ( .A(n4211), .B(n4210), .ZN(n4212) );
  XNOR2_X1 U4708 ( .A(n4213), .B(n4212), .ZN(n4221) );
  OAI22_X1 U4709 ( .A1(n4468), .A2(n5280), .B1(n4214), .B2(n4467), .ZN(n4218)
         );
  OAI22_X1 U4710 ( .A1(n4458), .A2(n4216), .B1(STATE_REG_SCAN_IN), .B2(n4215), 
        .ZN(n4217) );
  AOI211_X1 U4711 ( .C1(n4219), .C2(n4464), .A(n4218), .B(n4217), .ZN(n4220)
         );
  OAI21_X1 U4712 ( .B1(n4221), .B2(n5271), .A(n4220), .ZN(U3237) );
  MUX2_X1 U4713 ( .A(n5314), .B(DATAO_REG_31__SCAN_IN), .S(n4235), .Z(U3581)
         );
  MUX2_X1 U4714 ( .A(DATAO_REG_29__SCAN_IN), .B(n4430), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4715 ( .A(n4448), .B(DATAO_REG_28__SCAN_IN), .S(n4235), .Z(U3578)
         );
  MUX2_X1 U4716 ( .A(n4464), .B(DATAO_REG_27__SCAN_IN), .S(n4235), .Z(U3577)
         );
  MUX2_X1 U4717 ( .A(n4481), .B(DATAO_REG_26__SCAN_IN), .S(n4235), .Z(U3576)
         );
  MUX2_X1 U4718 ( .A(n4889), .B(DATAO_REG_25__SCAN_IN), .S(n4235), .Z(U3575)
         );
  MUX2_X1 U4719 ( .A(n4909), .B(DATAO_REG_24__SCAN_IN), .S(n4235), .Z(U3574)
         );
  MUX2_X1 U4720 ( .A(n4930), .B(DATAO_REG_23__SCAN_IN), .S(n4235), .Z(U3573)
         );
  MUX2_X1 U4721 ( .A(n4373), .B(DATAO_REG_22__SCAN_IN), .S(n4235), .Z(U3572)
         );
  MUX2_X1 U4722 ( .A(DATAO_REG_21__SCAN_IN), .B(n4222), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4723 ( .A(n4982), .B(DATAO_REG_20__SCAN_IN), .S(n4235), .Z(U3570)
         );
  MUX2_X1 U4724 ( .A(n4958), .B(DATAO_REG_19__SCAN_IN), .S(n4235), .Z(U3569)
         );
  MUX2_X1 U4725 ( .A(n4371), .B(DATAO_REG_18__SCAN_IN), .S(n4235), .Z(U3568)
         );
  MUX2_X1 U4726 ( .A(n5285), .B(DATAO_REG_17__SCAN_IN), .S(n4235), .Z(U3567)
         );
  MUX2_X1 U4727 ( .A(n4223), .B(DATAO_REG_16__SCAN_IN), .S(n4235), .Z(U3566)
         );
  MUX2_X1 U4728 ( .A(n5267), .B(DATAO_REG_15__SCAN_IN), .S(n4235), .Z(U3565)
         );
  MUX2_X1 U4729 ( .A(n4224), .B(DATAO_REG_14__SCAN_IN), .S(n4235), .Z(U3564)
         );
  MUX2_X1 U4730 ( .A(n4225), .B(DATAO_REG_13__SCAN_IN), .S(n4235), .Z(U3563)
         );
  MUX2_X1 U4731 ( .A(n4226), .B(DATAO_REG_12__SCAN_IN), .S(n4235), .Z(U3562)
         );
  MUX2_X1 U4732 ( .A(n4227), .B(DATAO_REG_11__SCAN_IN), .S(n4235), .Z(U3561)
         );
  MUX2_X1 U4733 ( .A(n4228), .B(DATAO_REG_10__SCAN_IN), .S(n4235), .Z(U3560)
         );
  MUX2_X1 U4734 ( .A(n4229), .B(DATAO_REG_9__SCAN_IN), .S(n4235), .Z(U3559) );
  MUX2_X1 U4735 ( .A(n4230), .B(DATAO_REG_8__SCAN_IN), .S(n4235), .Z(U3558) );
  MUX2_X1 U4736 ( .A(n4231), .B(DATAO_REG_7__SCAN_IN), .S(n4235), .Z(U3557) );
  MUX2_X1 U4737 ( .A(n4232), .B(DATAO_REG_6__SCAN_IN), .S(n4235), .Z(U3556) );
  MUX2_X1 U4738 ( .A(n4233), .B(DATAO_REG_5__SCAN_IN), .S(n4235), .Z(U3555) );
  MUX2_X1 U4739 ( .A(n3108), .B(DATAO_REG_4__SCAN_IN), .S(n4235), .Z(U3554) );
  MUX2_X1 U4740 ( .A(n4234), .B(DATAO_REG_3__SCAN_IN), .S(n4235), .Z(U3553) );
  MUX2_X1 U4741 ( .A(n3105), .B(DATAO_REG_2__SCAN_IN), .S(n4235), .Z(U3552) );
  MUX2_X1 U4742 ( .A(n3078), .B(DATAO_REG_1__SCAN_IN), .S(n4235), .Z(U3551) );
  MUX2_X1 U4743 ( .A(n4236), .B(DATAO_REG_0__SCAN_IN), .S(n4235), .Z(U3550) );
  INV_X1 U4744 ( .A(n5108), .ZN(n4362) );
  OAI211_X1 U4745 ( .C1(n4239), .C2(n4238), .A(n4362), .B(n4237), .ZN(n4247)
         );
  AOI22_X1 U4746 ( .A1(n5107), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4246) );
  INV_X1 U4747 ( .A(n4348), .ZN(n5114) );
  NAND2_X1 U4748 ( .A1(n5114), .A2(n2850), .ZN(n4245) );
  INV_X1 U4749 ( .A(n4240), .ZN(n4243) );
  OAI211_X1 U4750 ( .C1(n4243), .C2(n4242), .A(n5116), .B(n4241), .ZN(n4244)
         );
  NAND4_X1 U4751 ( .A1(n4247), .A2(n4246), .A3(n4245), .A4(n4244), .ZN(U3241)
         );
  NOR2_X1 U4752 ( .A1(n4348), .A2(n2588), .ZN(n4249) );
  AOI211_X1 U4753 ( .C1(n5107), .C2(ADDR_REG_3__SCAN_IN), .A(n4250), .B(n4249), 
        .ZN(n4258) );
  AOI211_X1 U4754 ( .C1(n5160), .C2(n4252), .A(n4251), .B(n5108), .ZN(n4253)
         );
  INV_X1 U4755 ( .A(n4253), .ZN(n4257) );
  OAI211_X1 U4756 ( .C1(REG2_REG_3__SCAN_IN), .C2(n4255), .A(n5116), .B(n4254), 
        .ZN(n4256) );
  NAND3_X1 U4757 ( .A1(n4258), .A2(n4257), .A3(n4256), .ZN(U3243) );
  OAI211_X1 U4758 ( .C1(n4260), .C2(REG2_REG_6__SCAN_IN), .A(n5116), .B(n4259), 
        .ZN(n4268) );
  AOI21_X1 U4759 ( .B1(n5107), .B2(ADDR_REG_6__SCAN_IN), .A(n4261), .ZN(n4267)
         );
  AOI21_X1 U4760 ( .B1(n4263), .B2(n5187), .A(n4262), .ZN(n4264) );
  NAND2_X1 U4761 ( .A1(n4362), .A2(n4264), .ZN(n4266) );
  OR2_X1 U4762 ( .A1(n4348), .A2(n5183), .ZN(n4265) );
  NAND4_X1 U4763 ( .A1(n4268), .A2(n4267), .A3(n4266), .A4(n4265), .ZN(U3246)
         );
  OAI211_X1 U4764 ( .C1(REG1_REG_8__SCAN_IN), .C2(n4270), .A(n4362), .B(n4269), 
        .ZN(n4277) );
  AOI21_X1 U4765 ( .B1(n5107), .B2(ADDR_REG_8__SCAN_IN), .A(n4271), .ZN(n4276)
         );
  NAND2_X1 U4766 ( .A1(n5114), .A2(n5074), .ZN(n4275) );
  OAI211_X1 U4767 ( .C1(REG2_REG_8__SCAN_IN), .C2(n4273), .A(n5116), .B(n4272), 
        .ZN(n4274) );
  NAND4_X1 U4768 ( .A1(n4277), .A2(n4276), .A3(n4275), .A4(n4274), .ZN(U3248)
         );
  NOR2_X1 U4769 ( .A1(n4348), .A2(n5206), .ZN(n4278) );
  AOI211_X1 U4770 ( .C1(n5107), .C2(ADDR_REG_9__SCAN_IN), .A(n4279), .B(n4278), 
        .ZN(n4289) );
  AOI211_X1 U4771 ( .C1(n4282), .C2(n4281), .A(n4280), .B(n5108), .ZN(n4283)
         );
  INV_X1 U4772 ( .A(n4283), .ZN(n4288) );
  OAI211_X1 U4773 ( .C1(n4286), .C2(n4285), .A(n5116), .B(n4284), .ZN(n4287)
         );
  NAND3_X1 U4774 ( .A1(n4289), .A2(n4288), .A3(n4287), .ZN(U3249) );
  OAI211_X1 U4775 ( .C1(n4291), .C2(REG2_REG_10__SCAN_IN), .A(n5116), .B(n4290), .ZN(n4299) );
  AOI21_X1 U4776 ( .B1(n5107), .B2(ADDR_REG_10__SCAN_IN), .A(n4292), .ZN(n4298) );
  AOI21_X1 U4777 ( .B1(n4294), .B2(n5218), .A(n4293), .ZN(n4295) );
  NAND2_X1 U4778 ( .A1(n4362), .A2(n4295), .ZN(n4297) );
  OR2_X1 U4779 ( .A1(n4348), .A2(n2601), .ZN(n4296) );
  NAND4_X1 U4780 ( .A1(n4299), .A2(n4298), .A3(n4297), .A4(n4296), .ZN(U3250)
         );
  OAI211_X1 U4781 ( .C1(n4301), .C2(REG2_REG_12__SCAN_IN), .A(n5116), .B(n4300), .ZN(n4309) );
  AOI21_X1 U4782 ( .B1(n5107), .B2(ADDR_REG_12__SCAN_IN), .A(n4302), .ZN(n4308) );
  AOI21_X1 U4783 ( .B1(n4304), .B2(n5236), .A(n4303), .ZN(n4305) );
  NAND2_X1 U4784 ( .A1(n4362), .A2(n4305), .ZN(n4307) );
  OR2_X1 U4785 ( .A1(n4348), .A2(n5231), .ZN(n4306) );
  NAND4_X1 U4786 ( .A1(n4309), .A2(n4308), .A3(n4307), .A4(n4306), .ZN(U3252)
         );
  OAI211_X1 U4787 ( .C1(n4311), .C2(REG2_REG_14__SCAN_IN), .A(n5116), .B(n4310), .ZN(n4319) );
  AOI21_X1 U4788 ( .B1(n5107), .B2(ADDR_REG_14__SCAN_IN), .A(n4312), .ZN(n4318) );
  AOI21_X1 U4789 ( .B1(n4314), .B2(n5252), .A(n4313), .ZN(n4315) );
  NAND2_X1 U4790 ( .A1(n4362), .A2(n4315), .ZN(n4317) );
  OR2_X1 U4791 ( .A1(n4348), .A2(n2587), .ZN(n4316) );
  NAND4_X1 U4792 ( .A1(n4319), .A2(n4318), .A3(n4317), .A4(n4316), .ZN(U3254)
         );
  AOI211_X1 U4793 ( .C1(n4321), .C2(n4320), .A(n2509), .B(n5108), .ZN(n4330)
         );
  OAI211_X1 U4794 ( .C1(n4324), .C2(n4323), .A(n5116), .B(n4322), .ZN(n4327)
         );
  AOI21_X1 U4795 ( .B1(n5107), .B2(ADDR_REG_15__SCAN_IN), .A(n4325), .ZN(n4326) );
  OAI211_X1 U4796 ( .C1(n4348), .C2(n4328), .A(n4327), .B(n4326), .ZN(n4329)
         );
  OR2_X1 U4797 ( .A1(n4330), .A2(n4329), .ZN(U3255) );
  OAI21_X1 U4798 ( .B1(n4332), .B2(n5299), .A(n4331), .ZN(n4339) );
  NOR2_X1 U4799 ( .A1(STATE_REG_SCAN_IN), .A2(n4553), .ZN(n5275) );
  AOI21_X1 U4800 ( .B1(n5107), .B2(ADDR_REG_16__SCAN_IN), .A(n5275), .ZN(n4333) );
  OAI21_X1 U4801 ( .B1(n4348), .B2(n5264), .A(n4333), .ZN(n4338) );
  AOI21_X1 U4802 ( .B1(n4335), .B2(REG2_REG_16__SCAN_IN), .A(n4334), .ZN(n4336) );
  NOR2_X1 U4803 ( .A1(n4336), .A2(n2895), .ZN(n4337) );
  AOI211_X1 U4804 ( .C1(n4362), .C2(n4339), .A(n4338), .B(n4337), .ZN(n4340)
         );
  INV_X1 U4805 ( .A(n4340), .ZN(U3256) );
  NAND3_X1 U4806 ( .A1(REG2_REG_17__SCAN_IN), .A2(n4342), .A3(n5072), .ZN(
        n4344) );
  OAI21_X1 U4807 ( .B1(n4342), .B2(n4341), .A(n4357), .ZN(n4343) );
  NAND2_X1 U4808 ( .A1(n4344), .A2(n4343), .ZN(n4354) );
  INV_X1 U4809 ( .A(n5072), .ZN(n4347) );
  NAND2_X1 U4810 ( .A1(n5107), .A2(ADDR_REG_17__SCAN_IN), .ZN(n4345) );
  OAI211_X1 U4811 ( .C1(n4348), .C2(n4347), .A(n4346), .B(n4345), .ZN(n4353)
         );
  AOI211_X1 U4812 ( .C1(n4351), .C2(n4350), .A(n4349), .B(n5108), .ZN(n4352)
         );
  AOI211_X1 U4813 ( .C1(n5116), .C2(n4354), .A(n4353), .B(n4352), .ZN(n4355)
         );
  INV_X1 U4814 ( .A(n4355), .ZN(U3257) );
  AOI21_X1 U4815 ( .B1(n4358), .B2(n4357), .A(n4356), .ZN(n4359) );
  AOI22_X1 U4816 ( .A1(n5114), .A2(n5071), .B1(n5116), .B2(n4359), .ZN(n4367)
         );
  AOI21_X1 U4817 ( .B1(n5107), .B2(ADDR_REG_18__SCAN_IN), .A(n4360), .ZN(n4366) );
  OAI211_X1 U4818 ( .C1(n4364), .C2(n4363), .A(n4362), .B(n4361), .ZN(n4365)
         );
  NAND3_X1 U4819 ( .A1(n4367), .A2(n4366), .A3(n4365), .ZN(U3258) );
  NAND2_X1 U4820 ( .A1(n4952), .A2(n4955), .ZN(n4951) );
  NAND2_X1 U4821 ( .A1(n4951), .A2(n2527), .ZN(n4935) );
  NAND2_X1 U4822 ( .A1(n4909), .A2(n4385), .ZN(n4376) );
  INV_X1 U4823 ( .A(n4481), .ZN(n4441) );
  INV_X1 U4824 ( .A(n4467), .ZN(n4377) );
  INV_X1 U4825 ( .A(n4450), .ZN(n4381) );
  NAND2_X1 U4826 ( .A1(n4464), .A2(n4381), .ZN(n4382) );
  INV_X1 U4827 ( .A(n5000), .ZN(n4420) );
  INV_X1 U4828 ( .A(n4413), .ZN(n4386) );
  NOR2_X2 U4829 ( .A1(n4963), .A2(n4938), .ZN(n4921) );
  AOI211_X1 U4830 ( .C1(n4386), .C2(n4432), .A(n5296), .B(n5330), .ZN(n5001)
         );
  INV_X1 U4831 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4387) );
  OAI22_X1 U4832 ( .A1(n4388), .A2(n4991), .B1(n4387), .B2(n5138), .ZN(n4389)
         );
  AOI21_X1 U4833 ( .B1(n5001), .B2(n4390), .A(n4389), .ZN(n4419) );
  INV_X1 U4834 ( .A(n4391), .ZN(n4394) );
  INV_X1 U4835 ( .A(n4392), .ZN(n4393) );
  OAI21_X1 U4836 ( .B1(n4395), .B2(n4394), .A(n4393), .ZN(n4954) );
  AOI21_X2 U4837 ( .B1(n4954), .B2(n4397), .A(n4396), .ZN(n4937) );
  INV_X1 U4838 ( .A(n4398), .ZN(n4400) );
  AOI21_X1 U4839 ( .B1(n4937), .B2(n4400), .A(n4399), .ZN(n4883) );
  INV_X1 U4840 ( .A(n4401), .ZN(n4403) );
  OAI21_X1 U4841 ( .B1(n4476), .B2(n4405), .A(n4404), .ZN(n4460) );
  NOR2_X1 U4842 ( .A1(n4426), .A2(n4425), .ZN(n4424) );
  NOR2_X1 U4843 ( .A1(n4424), .A2(n4408), .ZN(n4410) );
  XNOR2_X1 U4844 ( .A(n4410), .B(n2693), .ZN(n4417) );
  INV_X1 U4845 ( .A(B_REG_SCAN_IN), .ZN(n4411) );
  OR2_X1 U4846 ( .A1(n2846), .A2(n4411), .ZN(n4412) );
  NAND2_X1 U4847 ( .A1(n5286), .A2(n4412), .ZN(n5312) );
  OAI22_X1 U4848 ( .A1(n4414), .A2(n5312), .B1(n5315), .B2(n4413), .ZN(n4415)
         );
  AOI21_X1 U4849 ( .B1(n4448), .B2(n4957), .A(n4415), .ZN(n4416) );
  OAI21_X1 U4850 ( .B1(n4417), .B2(n5288), .A(n4416), .ZN(n5002) );
  NAND2_X1 U4851 ( .A1(n5002), .A2(n5138), .ZN(n4418) );
  OAI211_X1 U4852 ( .C1(n4420), .C2(n5307), .A(n4419), .B(n4418), .ZN(U3354)
         );
  XNOR2_X1 U4853 ( .A(n4421), .B(n4425), .ZN(n5011) );
  OAI22_X1 U4854 ( .A1(n4423), .A2(n5282), .B1(n5315), .B2(n4422), .ZN(n4429)
         );
  NOR2_X1 U4855 ( .A1(n4427), .A2(n5288), .ZN(n4428) );
  AOI21_X1 U4856 ( .B1(n4449), .B2(n4431), .A(n5296), .ZN(n4433) );
  NAND2_X1 U4857 ( .A1(n4433), .A2(n4432), .ZN(n5010) );
  INV_X1 U4858 ( .A(n4434), .ZN(n4435) );
  AOI22_X1 U4859 ( .A1(n4435), .A2(n5303), .B1(REG2_REG_28__SCAN_IN), .B2(
        n5333), .ZN(n4436) );
  OAI21_X1 U4860 ( .B1(n5010), .B2(n4969), .A(n4436), .ZN(n4437) );
  AOI21_X1 U4861 ( .B1(n4438), .B2(n5138), .A(n4437), .ZN(n4439) );
  OAI21_X1 U4862 ( .B1(n5011), .B2(n5307), .A(n4439), .ZN(U3262) );
  XNOR2_X1 U4863 ( .A(n4440), .B(n4443), .ZN(n5014) );
  OAI22_X1 U4864 ( .A1(n4441), .A2(n5282), .B1(n5315), .B2(n4450), .ZN(n4447)
         );
  AOI21_X1 U4865 ( .B1(n4444), .B2(n4443), .A(n4442), .ZN(n4445) );
  NOR2_X1 U4866 ( .A1(n4445), .A2(n5288), .ZN(n4446) );
  AOI211_X1 U4867 ( .C1(n5286), .C2(n4448), .A(n4447), .B(n4446), .ZN(n5013)
         );
  INV_X1 U4868 ( .A(n2492), .ZN(n4454) );
  OAI211_X1 U4869 ( .C1(n4465), .C2(n4450), .A(n5339), .B(n4449), .ZN(n5012)
         );
  AOI22_X1 U4870 ( .A1(n4451), .A2(n5303), .B1(REG2_REG_27__SCAN_IN), .B2(
        n5333), .ZN(n4452) );
  OAI21_X1 U4871 ( .B1(n5012), .B2(n4969), .A(n4452), .ZN(n4453) );
  AOI21_X1 U4872 ( .B1(n4454), .B2(n5138), .A(n4453), .ZN(n4455) );
  OAI21_X1 U4873 ( .B1(n5014), .B2(n5307), .A(n4455), .ZN(U3263) );
  OAI21_X1 U4874 ( .B1(n4457), .B2(n4459), .A(n4456), .ZN(n5017) );
  OAI22_X1 U4875 ( .A1(n4458), .A2(n5282), .B1(n4467), .B2(n5315), .ZN(n4463)
         );
  XNOR2_X1 U4876 ( .A(n4460), .B(n4459), .ZN(n4461) );
  NOR2_X1 U4877 ( .A1(n4461), .A2(n5288), .ZN(n4462) );
  AOI211_X1 U4878 ( .C1(n5286), .C2(n4464), .A(n4463), .B(n4462), .ZN(n5016)
         );
  INV_X1 U4879 ( .A(n5016), .ZN(n4472) );
  INV_X1 U4880 ( .A(n4465), .ZN(n4466) );
  OAI211_X1 U4881 ( .C1(n4484), .C2(n4467), .A(n4466), .B(n5339), .ZN(n5015)
         );
  INV_X1 U4882 ( .A(n4468), .ZN(n4469) );
  AOI22_X1 U4883 ( .A1(n4469), .A2(n5303), .B1(REG2_REG_26__SCAN_IN), .B2(
        n5333), .ZN(n4470) );
  OAI21_X1 U4884 ( .B1(n5015), .B2(n4969), .A(n4470), .ZN(n4471) );
  AOI21_X1 U4885 ( .B1(n4472), .B2(n5138), .A(n4471), .ZN(n4473) );
  OAI21_X1 U4886 ( .B1(n5017), .B2(n5307), .A(n4473), .ZN(U3264) );
  OAI21_X1 U4887 ( .B1(n4474), .B2(n4477), .A(n4475), .ZN(n5021) );
  XOR2_X1 U4888 ( .A(n4477), .B(n4476), .Z(n4483) );
  OAI22_X1 U4889 ( .A1(n4479), .A2(n5282), .B1(n5315), .B2(n4478), .ZN(n4480)
         );
  AOI21_X1 U4890 ( .B1(n5286), .B2(n4481), .A(n4480), .ZN(n4482) );
  OAI21_X1 U4891 ( .B1(n4483), .B2(n5288), .A(n4482), .ZN(n5018) );
  AOI21_X1 U4892 ( .B1(n4485), .B2(n4890), .A(n4484), .ZN(n5019) );
  INV_X1 U4893 ( .A(n5019), .ZN(n4488) );
  AOI22_X1 U4894 ( .A1(n4486), .A2(n5303), .B1(REG2_REG_25__SCAN_IN), .B2(
        n5336), .ZN(n4487) );
  OAI21_X1 U4895 ( .B1(n4488), .B2(n5306), .A(n4487), .ZN(n4489) );
  AOI21_X1 U4896 ( .B1(n5018), .B2(n5138), .A(n4489), .ZN(n4490) );
  OAI21_X1 U4897 ( .B1(n5021), .B2(n5307), .A(n4490), .ZN(n4879) );
  XOR2_X1 U4898 ( .A(DATAI_29_), .B(keyinput_2), .Z(n4493) );
  XOR2_X1 U4899 ( .A(DATAI_27_), .B(keyinput_4), .Z(n4492) );
  XNOR2_X1 U4900 ( .A(DATAI_30_), .B(keyinput_1), .ZN(n4491) );
  NOR3_X1 U4901 ( .A1(n4493), .A2(n4492), .A3(n4491), .ZN(n4496) );
  XOR2_X1 U4902 ( .A(DATAI_28_), .B(keyinput_3), .Z(n4495) );
  XOR2_X1 U4903 ( .A(DATAI_31_), .B(keyinput_0), .Z(n4494) );
  NAND3_X1 U4904 ( .A1(n4496), .A2(n4495), .A3(n4494), .ZN(n4499) );
  XNOR2_X1 U4905 ( .A(DATAI_26_), .B(keyinput_5), .ZN(n4498) );
  XNOR2_X1 U4906 ( .A(DATAI_25_), .B(keyinput_6), .ZN(n4497) );
  AOI21_X1 U4907 ( .B1(n4499), .B2(n4498), .A(n4497), .ZN(n4502) );
  XOR2_X1 U4908 ( .A(DATAI_23_), .B(keyinput_8), .Z(n4501) );
  XNOR2_X1 U4909 ( .A(DATAI_24_), .B(keyinput_7), .ZN(n4500) );
  NOR3_X1 U4910 ( .A1(n4502), .A2(n4501), .A3(n4500), .ZN(n4513) );
  XNOR2_X1 U4911 ( .A(DATAI_15_), .B(keyinput_16), .ZN(n4506) );
  XNOR2_X1 U4912 ( .A(DATAI_21_), .B(keyinput_10), .ZN(n4505) );
  XNOR2_X1 U4913 ( .A(DATAI_17_), .B(keyinput_14), .ZN(n4504) );
  XNOR2_X1 U4914 ( .A(DATAI_20_), .B(keyinput_11), .ZN(n4503) );
  NAND4_X1 U4915 ( .A1(n4506), .A2(n4505), .A3(n4504), .A4(n4503), .ZN(n4512)
         );
  XOR2_X1 U4916 ( .A(DATAI_16_), .B(keyinput_15), .Z(n4510) );
  XOR2_X1 U4917 ( .A(DATAI_18_), .B(keyinput_13), .Z(n4509) );
  XOR2_X1 U4918 ( .A(DATAI_22_), .B(keyinput_9), .Z(n4508) );
  XOR2_X1 U4919 ( .A(DATAI_19_), .B(keyinput_12), .Z(n4507) );
  NAND4_X1 U4920 ( .A1(n4510), .A2(n4509), .A3(n4508), .A4(n4507), .ZN(n4511)
         );
  NOR3_X1 U4921 ( .A1(n4513), .A2(n4512), .A3(n4511), .ZN(n4516) );
  XNOR2_X1 U4922 ( .A(DATAI_14_), .B(keyinput_17), .ZN(n4515) );
  XNOR2_X1 U4923 ( .A(DATAI_13_), .B(keyinput_18), .ZN(n4514) );
  OAI21_X1 U4924 ( .B1(n4516), .B2(n4515), .A(n4514), .ZN(n4520) );
  XNOR2_X1 U4925 ( .A(DATAI_12_), .B(keyinput_19), .ZN(n4519) );
  INV_X1 U4926 ( .A(DATAI_11_), .ZN(n5221) );
  XNOR2_X1 U4927 ( .A(n5221), .B(keyinput_20), .ZN(n4518) );
  XNOR2_X1 U4928 ( .A(DATAI_10_), .B(keyinput_21), .ZN(n4517) );
  AOI211_X1 U4929 ( .C1(n4520), .C2(n4519), .A(n4518), .B(n4517), .ZN(n4523)
         );
  XOR2_X1 U4930 ( .A(DATAI_8_), .B(keyinput_23), .Z(n4522) );
  XNOR2_X1 U4931 ( .A(DATAI_9_), .B(keyinput_22), .ZN(n4521) );
  NOR3_X1 U4932 ( .A1(n4523), .A2(n4522), .A3(n4521), .ZN(n4527) );
  INV_X1 U4933 ( .A(DATAI_5_), .ZN(n5173) );
  XNOR2_X1 U4934 ( .A(n5173), .B(keyinput_26), .ZN(n4526) );
  INV_X1 U4935 ( .A(DATAI_7_), .ZN(n5190) );
  XNOR2_X1 U4936 ( .A(n5190), .B(keyinput_24), .ZN(n4525) );
  XNOR2_X1 U4937 ( .A(DATAI_6_), .B(keyinput_25), .ZN(n4524) );
  NOR4_X1 U4938 ( .A1(n4527), .A2(n4526), .A3(n4525), .A4(n4524), .ZN(n4530)
         );
  INV_X1 U4939 ( .A(DATAI_4_), .ZN(n5163) );
  XNOR2_X1 U4940 ( .A(n5163), .B(keyinput_27), .ZN(n4529) );
  XNOR2_X1 U4941 ( .A(DATAI_3_), .B(keyinput_28), .ZN(n4528) );
  OAI21_X1 U4942 ( .B1(n4530), .B2(n4529), .A(n4528), .ZN(n4532) );
  XNOR2_X1 U4943 ( .A(DATAI_2_), .B(keyinput_29), .ZN(n4531) );
  NAND2_X1 U4944 ( .A1(n4532), .A2(n4531), .ZN(n4536) );
  XOR2_X1 U4945 ( .A(DATAI_0_), .B(keyinput_31), .Z(n4535) );
  XNOR2_X1 U4946 ( .A(DATAI_1_), .B(keyinput_30), .ZN(n4534) );
  XNOR2_X1 U4947 ( .A(STATE_REG_SCAN_IN), .B(keyinput_32), .ZN(n4533) );
  NAND4_X1 U4948 ( .A1(n4536), .A2(n4535), .A3(n4534), .A4(n4533), .ZN(n4542)
         );
  XOR2_X1 U4949 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_33), .Z(n4541) );
  XNOR2_X1 U4950 ( .A(n4726), .B(keyinput_35), .ZN(n4539) );
  XNOR2_X1 U4951 ( .A(REG3_REG_27__SCAN_IN), .B(keyinput_34), .ZN(n4538) );
  XNOR2_X1 U4952 ( .A(REG3_REG_23__SCAN_IN), .B(keyinput_36), .ZN(n4537) );
  NAND3_X1 U4953 ( .A1(n4539), .A2(n4538), .A3(n4537), .ZN(n4540) );
  AOI21_X1 U4954 ( .B1(n4542), .B2(n4541), .A(n4540), .ZN(n4548) );
  INV_X1 U4955 ( .A(REG3_REG_28__SCAN_IN), .ZN(n4734) );
  AOI22_X1 U4956 ( .A1(n3068), .A2(keyinput_38), .B1(keyinput_40), .B2(n4734), 
        .ZN(n4543) );
  OAI221_X1 U4957 ( .B1(n3068), .B2(keyinput_38), .C1(n4734), .C2(keyinput_40), 
        .A(n4543), .ZN(n4547) );
  AOI22_X1 U4958 ( .A1(REG3_REG_10__SCAN_IN), .A2(keyinput_37), .B1(n4736), 
        .B2(keyinput_41), .ZN(n4544) );
  OAI221_X1 U4959 ( .B1(REG3_REG_10__SCAN_IN), .B2(keyinput_37), .C1(n4736), 
        .C2(keyinput_41), .A(n4544), .ZN(n4546) );
  XNOR2_X1 U4960 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_39), .ZN(n4545) );
  NOR4_X1 U4961 ( .A1(n4548), .A2(n4547), .A3(n4546), .A4(n4545), .ZN(n4556)
         );
  XOR2_X1 U4962 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_42), .Z(n4552) );
  XOR2_X1 U4963 ( .A(REG3_REG_21__SCAN_IN), .B(keyinput_43), .Z(n4551) );
  XNOR2_X1 U4964 ( .A(n4741), .B(keyinput_45), .ZN(n4550) );
  XNOR2_X1 U4965 ( .A(REG3_REG_12__SCAN_IN), .B(keyinput_44), .ZN(n4549) );
  NAND4_X1 U4966 ( .A1(n4552), .A2(n4551), .A3(n4550), .A4(n4549), .ZN(n4555)
         );
  XNOR2_X1 U4967 ( .A(n4553), .B(keyinput_46), .ZN(n4554) );
  OAI21_X1 U4968 ( .B1(n4556), .B2(n4555), .A(n4554), .ZN(n4560) );
  XOR2_X1 U4969 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput_47), .Z(n4559) );
  XNOR2_X1 U4970 ( .A(n4749), .B(keyinput_48), .ZN(n4558) );
  XNOR2_X1 U4971 ( .A(REG3_REG_24__SCAN_IN), .B(keyinput_49), .ZN(n4557) );
  AOI211_X1 U4972 ( .C1(n4560), .C2(n4559), .A(n4558), .B(n4557), .ZN(n4564)
         );
  XOR2_X1 U4973 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_50), .Z(n4563) );
  XNOR2_X1 U4974 ( .A(n4561), .B(keyinput_51), .ZN(n4562) );
  NOR3_X1 U4975 ( .A1(n4564), .A2(n4563), .A3(n4562), .ZN(n4567) );
  XNOR2_X1 U4976 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_52), .ZN(n4566) );
  XNOR2_X1 U4977 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_53), .ZN(n4565) );
  OAI21_X1 U4978 ( .B1(n4567), .B2(n4566), .A(n4565), .ZN(n4570) );
  XOR2_X1 U4979 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_55), .Z(n4569) );
  XNOR2_X1 U4980 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput_54), .ZN(n4568) );
  NAND3_X1 U4981 ( .A1(n4570), .A2(n4569), .A3(n4568), .ZN(n4578) );
  XNOR2_X1 U4982 ( .A(n4571), .B(keyinput_58), .ZN(n4577) );
  XOR2_X1 U4983 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_56), .Z(n4576) );
  XNOR2_X1 U4984 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_57), .ZN(n4574) );
  XNOR2_X1 U4985 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_59), .ZN(n4573) );
  XNOR2_X1 U4986 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_60), .ZN(n4572) );
  NOR3_X1 U4987 ( .A1(n4574), .A2(n4573), .A3(n4572), .ZN(n4575) );
  NAND4_X1 U4988 ( .A1(n4578), .A2(n4577), .A3(n4576), .A4(n4575), .ZN(n4582)
         );
  XNOR2_X1 U4989 ( .A(n4579), .B(keyinput_62), .ZN(n4581) );
  XNOR2_X1 U4990 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_61), .ZN(n4580) );
  NAND3_X1 U4991 ( .A1(n4582), .A2(n4581), .A3(n4580), .ZN(n4586) );
  XNOR2_X1 U4992 ( .A(n4776), .B(keyinput_64), .ZN(n4585) );
  XNOR2_X1 U4993 ( .A(n4775), .B(keyinput_65), .ZN(n4584) );
  XOR2_X1 U4994 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_63), .Z(n4583) );
  NAND4_X1 U4995 ( .A1(n4586), .A2(n4585), .A3(n4584), .A4(n4583), .ZN(n4590)
         );
  XNOR2_X1 U4996 ( .A(IR_REG_11__SCAN_IN), .B(keyinput_66), .ZN(n4589) );
  XNOR2_X1 U4997 ( .A(n4587), .B(keyinput_67), .ZN(n4588) );
  AOI21_X1 U4998 ( .B1(n4590), .B2(n4589), .A(n4588), .ZN(n4594) );
  XNOR2_X1 U4999 ( .A(n4591), .B(keyinput_68), .ZN(n4593) );
  XNOR2_X1 U5000 ( .A(IR_REG_14__SCAN_IN), .B(keyinput_69), .ZN(n4592) );
  OAI21_X1 U5001 ( .B1(n4594), .B2(n4593), .A(n4592), .ZN(n4603) );
  INV_X1 U5002 ( .A(IR_REG_17__SCAN_IN), .ZN(n4596) );
  AOI22_X1 U5003 ( .A1(n4596), .A2(keyinput_72), .B1(keyinput_74), .B2(n4789), 
        .ZN(n4595) );
  OAI221_X1 U5004 ( .B1(n4596), .B2(keyinput_72), .C1(n4789), .C2(keyinput_74), 
        .A(n4595), .ZN(n4601) );
  XNOR2_X1 U5005 ( .A(n4597), .B(keyinput_70), .ZN(n4600) );
  XOR2_X1 U5006 ( .A(IR_REG_16__SCAN_IN), .B(keyinput_71), .Z(n4599) );
  XNOR2_X1 U5007 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_73), .ZN(n4598) );
  NOR4_X1 U5008 ( .A1(n4601), .A2(n4600), .A3(n4599), .A4(n4598), .ZN(n4602)
         );
  NAND2_X1 U5009 ( .A1(n4603), .A2(n4602), .ZN(n4608) );
  XNOR2_X1 U5010 ( .A(n4604), .B(keyinput_77), .ZN(n4607) );
  XNOR2_X1 U5011 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_76), .ZN(n4606) );
  XNOR2_X1 U5012 ( .A(IR_REG_20__SCAN_IN), .B(keyinput_75), .ZN(n4605) );
  NAND4_X1 U5013 ( .A1(n4608), .A2(n4607), .A3(n4606), .A4(n4605), .ZN(n4612)
         );
  XNOR2_X1 U5014 ( .A(IR_REG_23__SCAN_IN), .B(keyinput_78), .ZN(n4611) );
  XNOR2_X1 U5015 ( .A(n4800), .B(keyinput_79), .ZN(n4610) );
  XNOR2_X1 U5016 ( .A(IR_REG_25__SCAN_IN), .B(keyinput_80), .ZN(n4609) );
  AOI211_X1 U5017 ( .C1(n4612), .C2(n4611), .A(n4610), .B(n4609), .ZN(n4617)
         );
  XNOR2_X1 U5018 ( .A(n4806), .B(keyinput_81), .ZN(n4616) );
  XNOR2_X1 U5019 ( .A(n4613), .B(keyinput_82), .ZN(n4615) );
  XNOR2_X1 U5020 ( .A(IR_REG_28__SCAN_IN), .B(keyinput_83), .ZN(n4614) );
  NOR4_X1 U5021 ( .A1(n4617), .A2(n4616), .A3(n4615), .A4(n4614), .ZN(n4621)
         );
  XOR2_X1 U5022 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_86), .Z(n4620) );
  XOR2_X1 U5023 ( .A(IR_REG_30__SCAN_IN), .B(keyinput_85), .Z(n4619) );
  XNOR2_X1 U5024 ( .A(n4811), .B(keyinput_84), .ZN(n4618) );
  NOR4_X1 U5025 ( .A1(n4621), .A2(n4620), .A3(n4619), .A4(n4618), .ZN(n4625)
         );
  XNOR2_X1 U5026 ( .A(n4622), .B(keyinput_87), .ZN(n4624) );
  XOR2_X1 U5027 ( .A(D_REG_1__SCAN_IN), .B(keyinput_88), .Z(n4623) );
  OAI21_X1 U5028 ( .B1(n4625), .B2(n4624), .A(n4623), .ZN(n4629) );
  INV_X1 U5029 ( .A(D_REG_3__SCAN_IN), .ZN(n5076) );
  XNOR2_X1 U5030 ( .A(n5076), .B(keyinput_90), .ZN(n4628) );
  INV_X1 U5031 ( .A(D_REG_2__SCAN_IN), .ZN(n5075) );
  XNOR2_X1 U5032 ( .A(n5075), .B(keyinput_89), .ZN(n4627) );
  XOR2_X1 U5033 ( .A(D_REG_4__SCAN_IN), .B(keyinput_91), .Z(n4626) );
  NAND4_X1 U5034 ( .A1(n4629), .A2(n4628), .A3(n4627), .A4(n4626), .ZN(n4632)
         );
  XNOR2_X1 U5035 ( .A(D_REG_5__SCAN_IN), .B(keyinput_92), .ZN(n4631) );
  XNOR2_X1 U5036 ( .A(D_REG_6__SCAN_IN), .B(keyinput_93), .ZN(n4630) );
  NAND3_X1 U5037 ( .A1(n4632), .A2(n4631), .A3(n4630), .ZN(n4640) );
  INV_X1 U5038 ( .A(D_REG_11__SCAN_IN), .ZN(n5082) );
  XNOR2_X1 U5039 ( .A(n5082), .B(keyinput_98), .ZN(n4639) );
  XOR2_X1 U5040 ( .A(D_REG_7__SCAN_IN), .B(keyinput_94), .Z(n4638) );
  XOR2_X1 U5041 ( .A(D_REG_8__SCAN_IN), .B(keyinput_95), .Z(n4636) );
  XOR2_X1 U5042 ( .A(D_REG_12__SCAN_IN), .B(keyinput_99), .Z(n4635) );
  INV_X1 U5043 ( .A(D_REG_10__SCAN_IN), .ZN(n5081) );
  XNOR2_X1 U5044 ( .A(n5081), .B(keyinput_97), .ZN(n4634) );
  XNOR2_X1 U5045 ( .A(D_REG_9__SCAN_IN), .B(keyinput_96), .ZN(n4633) );
  NOR4_X1 U5046 ( .A1(n4636), .A2(n4635), .A3(n4634), .A4(n4633), .ZN(n4637)
         );
  NAND4_X1 U5047 ( .A1(n4640), .A2(n4639), .A3(n4638), .A4(n4637), .ZN(n4644)
         );
  XNOR2_X1 U5048 ( .A(D_REG_15__SCAN_IN), .B(keyinput_102), .ZN(n4643) );
  XNOR2_X1 U5049 ( .A(D_REG_13__SCAN_IN), .B(keyinput_100), .ZN(n4642) );
  XNOR2_X1 U5050 ( .A(D_REG_14__SCAN_IN), .B(keyinput_101), .ZN(n4641) );
  NAND4_X1 U5051 ( .A1(n4644), .A2(n4643), .A3(n4642), .A4(n4641), .ZN(n4648)
         );
  XNOR2_X1 U5052 ( .A(D_REG_16__SCAN_IN), .B(keyinput_103), .ZN(n4647) );
  XOR2_X1 U5053 ( .A(D_REG_17__SCAN_IN), .B(keyinput_104), .Z(n4646) );
  XNOR2_X1 U5054 ( .A(D_REG_18__SCAN_IN), .B(keyinput_105), .ZN(n4645) );
  AOI211_X1 U5055 ( .C1(n4648), .C2(n4647), .A(n4646), .B(n4645), .ZN(n4654)
         );
  INV_X1 U5056 ( .A(D_REG_19__SCAN_IN), .ZN(n5089) );
  XNOR2_X1 U5057 ( .A(n5089), .B(keyinput_106), .ZN(n4653) );
  INV_X1 U5058 ( .A(D_REG_21__SCAN_IN), .ZN(n5090) );
  XNOR2_X1 U5059 ( .A(n5090), .B(keyinput_108), .ZN(n4651) );
  XNOR2_X1 U5060 ( .A(D_REG_20__SCAN_IN), .B(keyinput_107), .ZN(n4650) );
  XNOR2_X1 U5061 ( .A(D_REG_22__SCAN_IN), .B(keyinput_109), .ZN(n4649) );
  NOR3_X1 U5062 ( .A1(n4651), .A2(n4650), .A3(n4649), .ZN(n4652) );
  OAI21_X1 U5063 ( .B1(n4654), .B2(n4653), .A(n4652), .ZN(n4658) );
  INV_X1 U5064 ( .A(D_REG_23__SCAN_IN), .ZN(n5092) );
  XNOR2_X1 U5065 ( .A(n5092), .B(keyinput_110), .ZN(n4657) );
  XNOR2_X1 U5066 ( .A(D_REG_25__SCAN_IN), .B(keyinput_112), .ZN(n4656) );
  XNOR2_X1 U5067 ( .A(D_REG_24__SCAN_IN), .B(keyinput_111), .ZN(n4655) );
  AOI211_X1 U5068 ( .C1(n4658), .C2(n4657), .A(n4656), .B(n4655), .ZN(n4661)
         );
  INV_X1 U5069 ( .A(D_REG_26__SCAN_IN), .ZN(n5093) );
  XNOR2_X1 U5070 ( .A(n5093), .B(keyinput_113), .ZN(n4660) );
  INV_X1 U5071 ( .A(D_REG_27__SCAN_IN), .ZN(n5094) );
  XNOR2_X1 U5072 ( .A(n5094), .B(keyinput_114), .ZN(n4659) );
  NOR3_X1 U5073 ( .A1(n4661), .A2(n4660), .A3(n4659), .ZN(n4665) );
  INV_X1 U5074 ( .A(D_REG_30__SCAN_IN), .ZN(n5097) );
  XNOR2_X1 U5075 ( .A(n5097), .B(keyinput_117), .ZN(n4664) );
  INV_X1 U5076 ( .A(D_REG_29__SCAN_IN), .ZN(n5096) );
  XNOR2_X1 U5077 ( .A(n5096), .B(keyinput_116), .ZN(n4663) );
  XNOR2_X1 U5078 ( .A(D_REG_28__SCAN_IN), .B(keyinput_115), .ZN(n4662) );
  NOR4_X1 U5079 ( .A1(n4665), .A2(n4664), .A3(n4663), .A4(n4662), .ZN(n4668)
         );
  XOR2_X1 U5080 ( .A(REG0_REG_0__SCAN_IN), .B(keyinput_119), .Z(n4667) );
  XNOR2_X1 U5081 ( .A(D_REG_31__SCAN_IN), .B(keyinput_118), .ZN(n4666) );
  NOR3_X1 U5082 ( .A1(n4668), .A2(n4667), .A3(n4666), .ZN(n4671) );
  XNOR2_X1 U5083 ( .A(REG0_REG_1__SCAN_IN), .B(keyinput_120), .ZN(n4670) );
  XOR2_X1 U5084 ( .A(REG0_REG_2__SCAN_IN), .B(keyinput_121), .Z(n4669) );
  OAI21_X1 U5085 ( .B1(n4671), .B2(n4670), .A(n4669), .ZN(n4674) );
  XOR2_X1 U5086 ( .A(REG0_REG_4__SCAN_IN), .B(keyinput_123), .Z(n4673) );
  XNOR2_X1 U5087 ( .A(REG0_REG_3__SCAN_IN), .B(keyinput_122), .ZN(n4672) );
  NAND3_X1 U5088 ( .A1(n4674), .A2(n4673), .A3(n4672), .ZN(n4677) );
  XNOR2_X1 U5089 ( .A(REG0_REG_5__SCAN_IN), .B(keyinput_124), .ZN(n4676) );
  XNOR2_X1 U5090 ( .A(REG0_REG_6__SCAN_IN), .B(keyinput_125), .ZN(n4675) );
  AOI21_X1 U5091 ( .B1(n4677), .B2(n4676), .A(n4675), .ZN(n4877) );
  XNOR2_X1 U5092 ( .A(REG0_REG_7__SCAN_IN), .B(keyinput_126), .ZN(n4876) );
  XOR2_X1 U5093 ( .A(DATAI_28_), .B(keyinput_131), .Z(n4680) );
  XNOR2_X1 U5094 ( .A(DATAI_30_), .B(keyinput_129), .ZN(n4679) );
  XNOR2_X1 U5095 ( .A(DATAI_29_), .B(keyinput_130), .ZN(n4678) );
  NOR3_X1 U5096 ( .A1(n4680), .A2(n4679), .A3(n4678), .ZN(n4683) );
  XOR2_X1 U5097 ( .A(DATAI_27_), .B(keyinput_132), .Z(n4682) );
  XOR2_X1 U5098 ( .A(DATAI_31_), .B(keyinput_128), .Z(n4681) );
  NAND3_X1 U5099 ( .A1(n4683), .A2(n4682), .A3(n4681), .ZN(n4686) );
  XNOR2_X1 U5100 ( .A(DATAI_26_), .B(keyinput_133), .ZN(n4685) );
  XOR2_X1 U5101 ( .A(DATAI_25_), .B(keyinput_134), .Z(n4684) );
  AOI21_X1 U5102 ( .B1(n4686), .B2(n4685), .A(n4684), .ZN(n4689) );
  XNOR2_X1 U5103 ( .A(DATAI_23_), .B(keyinput_136), .ZN(n4688) );
  XNOR2_X1 U5104 ( .A(DATAI_24_), .B(keyinput_135), .ZN(n4687) );
  NOR3_X1 U5105 ( .A1(n4689), .A2(n4688), .A3(n4687), .ZN(n4701) );
  INV_X1 U5106 ( .A(keyinput_142), .ZN(n4690) );
  XNOR2_X1 U5107 ( .A(n4690), .B(DATAI_17_), .ZN(n4694) );
  XNOR2_X1 U5108 ( .A(DATAI_20_), .B(keyinput_139), .ZN(n4693) );
  XNOR2_X1 U5109 ( .A(DATAI_21_), .B(keyinput_138), .ZN(n4692) );
  XNOR2_X1 U5110 ( .A(DATAI_15_), .B(keyinput_144), .ZN(n4691) );
  NAND4_X1 U5111 ( .A1(n4694), .A2(n4693), .A3(n4692), .A4(n4691), .ZN(n4700)
         );
  XOR2_X1 U5112 ( .A(DATAI_16_), .B(keyinput_143), .Z(n4698) );
  XOR2_X1 U5113 ( .A(DATAI_18_), .B(keyinput_141), .Z(n4697) );
  XOR2_X1 U5114 ( .A(DATAI_22_), .B(keyinput_137), .Z(n4696) );
  XOR2_X1 U5115 ( .A(DATAI_19_), .B(keyinput_140), .Z(n4695) );
  NAND4_X1 U5116 ( .A1(n4698), .A2(n4697), .A3(n4696), .A4(n4695), .ZN(n4699)
         );
  NOR3_X1 U5117 ( .A1(n4701), .A2(n4700), .A3(n4699), .ZN(n4704) );
  XNOR2_X1 U5118 ( .A(DATAI_14_), .B(keyinput_145), .ZN(n4703) );
  INV_X1 U5119 ( .A(DATAI_13_), .ZN(n5239) );
  XNOR2_X1 U5120 ( .A(n5239), .B(keyinput_146), .ZN(n4702) );
  OAI21_X1 U5121 ( .B1(n4704), .B2(n4703), .A(n4702), .ZN(n4708) );
  XNOR2_X1 U5122 ( .A(DATAI_12_), .B(keyinput_147), .ZN(n4707) );
  INV_X1 U5123 ( .A(DATAI_10_), .ZN(n5213) );
  XNOR2_X1 U5124 ( .A(n5213), .B(keyinput_149), .ZN(n4706) );
  XNOR2_X1 U5125 ( .A(n5221), .B(keyinput_148), .ZN(n4705) );
  AOI211_X1 U5126 ( .C1(n4708), .C2(n4707), .A(n4706), .B(n4705), .ZN(n4711)
         );
  XNOR2_X1 U5127 ( .A(DATAI_9_), .B(keyinput_150), .ZN(n4710) );
  XNOR2_X1 U5128 ( .A(DATAI_8_), .B(keyinput_151), .ZN(n4709) );
  NOR3_X1 U5129 ( .A1(n4711), .A2(n4710), .A3(n4709), .ZN(n4715) );
  XNOR2_X1 U5130 ( .A(n5190), .B(keyinput_152), .ZN(n4714) );
  XNOR2_X1 U5131 ( .A(n5173), .B(keyinput_154), .ZN(n4713) );
  XNOR2_X1 U5132 ( .A(DATAI_6_), .B(keyinput_153), .ZN(n4712) );
  NOR4_X1 U5133 ( .A1(n4715), .A2(n4714), .A3(n4713), .A4(n4712), .ZN(n4718)
         );
  XNOR2_X1 U5134 ( .A(n5163), .B(keyinput_155), .ZN(n4717) );
  XNOR2_X1 U5135 ( .A(DATAI_3_), .B(keyinput_156), .ZN(n4716) );
  OAI21_X1 U5136 ( .B1(n4718), .B2(n4717), .A(n4716), .ZN(n4720) );
  XOR2_X1 U5137 ( .A(DATAI_2_), .B(keyinput_157), .Z(n4719) );
  NAND2_X1 U5138 ( .A1(n4720), .A2(n4719), .ZN(n4724) );
  XOR2_X1 U5139 ( .A(DATAI_1_), .B(keyinput_158), .Z(n4723) );
  XOR2_X1 U5140 ( .A(DATAI_0_), .B(keyinput_159), .Z(n4722) );
  XNOR2_X1 U5141 ( .A(U3149), .B(keyinput_160), .ZN(n4721) );
  NAND4_X1 U5142 ( .A1(n4724), .A2(n4723), .A3(n4722), .A4(n4721), .ZN(n4732)
         );
  XOR2_X1 U5143 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_161), .Z(n4731) );
  XNOR2_X1 U5144 ( .A(n4725), .B(keyinput_162), .ZN(n4729) );
  XNOR2_X1 U5145 ( .A(n4726), .B(keyinput_163), .ZN(n4728) );
  XNOR2_X1 U5146 ( .A(REG3_REG_23__SCAN_IN), .B(keyinput_164), .ZN(n4727) );
  NAND3_X1 U5147 ( .A1(n4729), .A2(n4728), .A3(n4727), .ZN(n4730) );
  AOI21_X1 U5148 ( .B1(n4732), .B2(n4731), .A(n4730), .ZN(n4740) );
  AOI22_X1 U5149 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput_167), .B1(n4734), 
        .B2(keyinput_168), .ZN(n4733) );
  OAI221_X1 U5150 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_167), .C1(n4734), 
        .C2(keyinput_168), .A(n4733), .ZN(n4739) );
  AOI22_X1 U5151 ( .A1(n3068), .A2(keyinput_166), .B1(keyinput_169), .B2(n4736), .ZN(n4735) );
  OAI221_X1 U5152 ( .B1(n3068), .B2(keyinput_166), .C1(n4736), .C2(
        keyinput_169), .A(n4735), .ZN(n4738) );
  XNOR2_X1 U5153 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_165), .ZN(n4737) );
  NOR4_X1 U5154 ( .A1(n4740), .A2(n4739), .A3(n4738), .A4(n4737), .ZN(n4748)
         );
  XOR2_X1 U5155 ( .A(REG3_REG_12__SCAN_IN), .B(keyinput_172), .Z(n4745) );
  XNOR2_X1 U5156 ( .A(n4741), .B(keyinput_173), .ZN(n4744) );
  XNOR2_X1 U5157 ( .A(REG3_REG_21__SCAN_IN), .B(keyinput_171), .ZN(n4743) );
  XNOR2_X1 U5158 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_170), .ZN(n4742) );
  NAND4_X1 U5159 ( .A1(n4745), .A2(n4744), .A3(n4743), .A4(n4742), .ZN(n4747)
         );
  XNOR2_X1 U5160 ( .A(REG3_REG_16__SCAN_IN), .B(keyinput_174), .ZN(n4746) );
  OAI21_X1 U5161 ( .B1(n4748), .B2(n4747), .A(n4746), .ZN(n4753) );
  XOR2_X1 U5162 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput_175), .Z(n4752) );
  XNOR2_X1 U5163 ( .A(n4749), .B(keyinput_176), .ZN(n4751) );
  XNOR2_X1 U5164 ( .A(REG3_REG_24__SCAN_IN), .B(keyinput_177), .ZN(n4750) );
  AOI211_X1 U5165 ( .C1(n4753), .C2(n4752), .A(n4751), .B(n4750), .ZN(n4758)
         );
  XNOR2_X1 U5166 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_178), .ZN(n4755) );
  XNOR2_X1 U5167 ( .A(REG3_REG_9__SCAN_IN), .B(keyinput_179), .ZN(n4754) );
  NAND2_X1 U5168 ( .A1(n4755), .A2(n4754), .ZN(n4757) );
  XOR2_X1 U5169 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_180), .Z(n4756) );
  OAI21_X1 U5170 ( .B1(n4758), .B2(n4757), .A(n4756), .ZN(n4763) );
  XNOR2_X1 U5171 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_181), .ZN(n4762) );
  XNOR2_X1 U5172 ( .A(n4759), .B(keyinput_182), .ZN(n4761) );
  XNOR2_X1 U5173 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_183), .ZN(n4760) );
  AOI211_X1 U5174 ( .C1(n4763), .C2(n4762), .A(n4761), .B(n4760), .ZN(n4774)
         );
  XNOR2_X1 U5175 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_188), .ZN(n4765) );
  XNOR2_X1 U5176 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_184), .ZN(n4764) );
  NOR2_X1 U5177 ( .A1(n4765), .A2(n4764), .ZN(n4770) );
  XNOR2_X1 U5178 ( .A(n4766), .B(keyinput_185), .ZN(n4769) );
  XNOR2_X1 U5179 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_186), .ZN(n4768) );
  XNOR2_X1 U5180 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_187), .ZN(n4767) );
  NAND4_X1 U5181 ( .A1(n4770), .A2(n4769), .A3(n4768), .A4(n4767), .ZN(n4773)
         );
  XNOR2_X1 U5182 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_190), .ZN(n4772) );
  XNOR2_X1 U5183 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_189), .ZN(n4771) );
  OAI211_X1 U5184 ( .C1(n4774), .C2(n4773), .A(n4772), .B(n4771), .ZN(n4780)
         );
  XOR2_X1 U5185 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_191), .Z(n4779) );
  XNOR2_X1 U5186 ( .A(n4775), .B(keyinput_193), .ZN(n4778) );
  XNOR2_X1 U5187 ( .A(n4776), .B(keyinput_192), .ZN(n4777) );
  NAND4_X1 U5188 ( .A1(n4780), .A2(n4779), .A3(n4778), .A4(n4777), .ZN(n4784)
         );
  XNOR2_X1 U5189 ( .A(n4781), .B(keyinput_194), .ZN(n4783) );
  XNOR2_X1 U5190 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_195), .ZN(n4782) );
  AOI21_X1 U5191 ( .B1(n4784), .B2(n4783), .A(n4782), .ZN(n4787) );
  XNOR2_X1 U5192 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_196), .ZN(n4786) );
  XNOR2_X1 U5193 ( .A(IR_REG_14__SCAN_IN), .B(keyinput_197), .ZN(n4785) );
  OAI21_X1 U5194 ( .B1(n4787), .B2(n4786), .A(n4785), .ZN(n4794) );
  OAI22_X1 U5195 ( .A1(n2811), .A2(keyinput_201), .B1(IR_REG_17__SCAN_IN), 
        .B2(keyinput_200), .ZN(n4788) );
  AOI221_X1 U5196 ( .B1(n2811), .B2(keyinput_201), .C1(keyinput_200), .C2(
        IR_REG_17__SCAN_IN), .A(n4788), .ZN(n4793) );
  XNOR2_X1 U5197 ( .A(n4789), .B(keyinput_202), .ZN(n4792) );
  OAI22_X1 U5198 ( .A1(IR_REG_16__SCAN_IN), .A2(keyinput_199), .B1(
        IR_REG_15__SCAN_IN), .B2(keyinput_198), .ZN(n4790) );
  AOI221_X1 U5199 ( .B1(IR_REG_16__SCAN_IN), .B2(keyinput_199), .C1(
        keyinput_198), .C2(IR_REG_15__SCAN_IN), .A(n4790), .ZN(n4791) );
  NAND4_X1 U5200 ( .A1(n4794), .A2(n4793), .A3(n4792), .A4(n4791), .ZN(n4798)
         );
  XNOR2_X1 U5201 ( .A(IR_REG_22__SCAN_IN), .B(keyinput_205), .ZN(n4797) );
  XNOR2_X1 U5202 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_204), .ZN(n4796) );
  XNOR2_X1 U5203 ( .A(IR_REG_20__SCAN_IN), .B(keyinput_203), .ZN(n4795) );
  NAND4_X1 U5204 ( .A1(n4798), .A2(n4797), .A3(n4796), .A4(n4795), .ZN(n4805)
         );
  XNOR2_X1 U5205 ( .A(n4799), .B(keyinput_206), .ZN(n4804) );
  XNOR2_X1 U5206 ( .A(n4800), .B(keyinput_207), .ZN(n4803) );
  XNOR2_X1 U5207 ( .A(n4801), .B(keyinput_208), .ZN(n4802) );
  AOI211_X1 U5208 ( .C1(n4805), .C2(n4804), .A(n4803), .B(n4802), .ZN(n4810)
         );
  XNOR2_X1 U5209 ( .A(n4806), .B(keyinput_209), .ZN(n4809) );
  XNOR2_X1 U5210 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_210), .ZN(n4808) );
  XNOR2_X1 U5211 ( .A(IR_REG_28__SCAN_IN), .B(keyinput_211), .ZN(n4807) );
  NOR4_X1 U5212 ( .A1(n4810), .A2(n4809), .A3(n4808), .A4(n4807), .ZN(n4815)
         );
  XNOR2_X1 U5213 ( .A(n4811), .B(keyinput_212), .ZN(n4814) );
  XOR2_X1 U5214 ( .A(IR_REG_30__SCAN_IN), .B(keyinput_213), .Z(n4813) );
  XNOR2_X1 U5215 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_214), .ZN(n4812) );
  NOR4_X1 U5216 ( .A1(n4815), .A2(n4814), .A3(n4813), .A4(n4812), .ZN(n4818)
         );
  XNOR2_X1 U5217 ( .A(D_REG_0__SCAN_IN), .B(keyinput_215), .ZN(n4817) );
  XOR2_X1 U5218 ( .A(D_REG_1__SCAN_IN), .B(keyinput_216), .Z(n4816) );
  OAI21_X1 U5219 ( .B1(n4818), .B2(n4817), .A(n4816), .ZN(n4825) );
  XOR2_X1 U5220 ( .A(D_REG_4__SCAN_IN), .B(keyinput_219), .Z(n4821) );
  XNOR2_X1 U5221 ( .A(n5075), .B(keyinput_217), .ZN(n4820) );
  XNOR2_X1 U5222 ( .A(n5076), .B(keyinput_218), .ZN(n4819) );
  NOR3_X1 U5223 ( .A1(n4821), .A2(n4820), .A3(n4819), .ZN(n4824) );
  XOR2_X1 U5224 ( .A(keyinput_221), .B(D_REG_6__SCAN_IN), .Z(n4823) );
  XOR2_X1 U5225 ( .A(keyinput_220), .B(D_REG_5__SCAN_IN), .Z(n4822) );
  AOI211_X1 U5226 ( .C1(n4825), .C2(n4824), .A(n4823), .B(n4822), .ZN(n4833)
         );
  XNOR2_X1 U5227 ( .A(n5081), .B(keyinput_225), .ZN(n4832) );
  XNOR2_X1 U5228 ( .A(D_REG_7__SCAN_IN), .B(keyinput_222), .ZN(n4831) );
  XNOR2_X1 U5229 ( .A(keyinput_223), .B(D_REG_8__SCAN_IN), .ZN(n4829) );
  XNOR2_X1 U5230 ( .A(keyinput_227), .B(D_REG_12__SCAN_IN), .ZN(n4828) );
  XNOR2_X1 U5231 ( .A(keyinput_224), .B(D_REG_9__SCAN_IN), .ZN(n4827) );
  XNOR2_X1 U5232 ( .A(keyinput_226), .B(D_REG_11__SCAN_IN), .ZN(n4826) );
  NAND4_X1 U5233 ( .A1(n4829), .A2(n4828), .A3(n4827), .A4(n4826), .ZN(n4830)
         );
  NOR4_X1 U5234 ( .A1(n4833), .A2(n4832), .A3(n4831), .A4(n4830), .ZN(n4837)
         );
  INV_X1 U5235 ( .A(D_REG_13__SCAN_IN), .ZN(n5084) );
  XNOR2_X1 U5236 ( .A(n5084), .B(keyinput_228), .ZN(n4836) );
  XNOR2_X1 U5237 ( .A(keyinput_230), .B(D_REG_15__SCAN_IN), .ZN(n4835) );
  XNOR2_X1 U5238 ( .A(D_REG_14__SCAN_IN), .B(keyinput_229), .ZN(n4834) );
  NOR4_X1 U5239 ( .A1(n4837), .A2(n4836), .A3(n4835), .A4(n4834), .ZN(n4841)
         );
  XOR2_X1 U5240 ( .A(keyinput_231), .B(D_REG_16__SCAN_IN), .Z(n4840) );
  XNOR2_X1 U5241 ( .A(keyinput_233), .B(D_REG_18__SCAN_IN), .ZN(n4839) );
  XNOR2_X1 U5242 ( .A(keyinput_232), .B(D_REG_17__SCAN_IN), .ZN(n4838) );
  OAI211_X1 U5243 ( .C1(n4841), .C2(n4840), .A(n4839), .B(n4838), .ZN(n4843)
         );
  XNOR2_X1 U5244 ( .A(n5089), .B(keyinput_234), .ZN(n4842) );
  NAND2_X1 U5245 ( .A1(n4843), .A2(n4842), .ZN(n4847) );
  XNOR2_X1 U5246 ( .A(n5090), .B(keyinput_236), .ZN(n4846) );
  XOR2_X1 U5247 ( .A(D_REG_20__SCAN_IN), .B(keyinput_235), .Z(n4845) );
  XNOR2_X1 U5248 ( .A(keyinput_237), .B(D_REG_22__SCAN_IN), .ZN(n4844) );
  NAND4_X1 U5249 ( .A1(n4847), .A2(n4846), .A3(n4845), .A4(n4844), .ZN(n4851)
         );
  XNOR2_X1 U5250 ( .A(keyinput_238), .B(D_REG_23__SCAN_IN), .ZN(n4850) );
  XNOR2_X1 U5251 ( .A(D_REG_25__SCAN_IN), .B(keyinput_240), .ZN(n4849) );
  XNOR2_X1 U5252 ( .A(D_REG_24__SCAN_IN), .B(keyinput_239), .ZN(n4848) );
  AOI211_X1 U5253 ( .C1(n4851), .C2(n4850), .A(n4849), .B(n4848), .ZN(n4854)
         );
  XNOR2_X1 U5254 ( .A(keyinput_241), .B(D_REG_26__SCAN_IN), .ZN(n4853) );
  XNOR2_X1 U5255 ( .A(keyinput_242), .B(D_REG_27__SCAN_IN), .ZN(n4852) );
  NOR3_X1 U5256 ( .A1(n4854), .A2(n4853), .A3(n4852), .ZN(n4858) );
  XNOR2_X1 U5257 ( .A(keyinput_244), .B(D_REG_29__SCAN_IN), .ZN(n4857) );
  XNOR2_X1 U5258 ( .A(keyinput_245), .B(D_REG_30__SCAN_IN), .ZN(n4856) );
  XNOR2_X1 U5259 ( .A(D_REG_28__SCAN_IN), .B(keyinput_243), .ZN(n4855) );
  NOR4_X1 U5260 ( .A1(n4858), .A2(n4857), .A3(n4856), .A4(n4855), .ZN(n4861)
         );
  INV_X1 U5261 ( .A(D_REG_31__SCAN_IN), .ZN(n5098) );
  XNOR2_X1 U5262 ( .A(n5098), .B(keyinput_246), .ZN(n4860) );
  XNOR2_X1 U5263 ( .A(REG0_REG_0__SCAN_IN), .B(keyinput_247), .ZN(n4859) );
  NOR3_X1 U5264 ( .A1(n4861), .A2(n4860), .A3(n4859), .ZN(n4864) );
  XNOR2_X1 U5265 ( .A(REG0_REG_1__SCAN_IN), .B(keyinput_248), .ZN(n4863) );
  XOR2_X1 U5266 ( .A(REG0_REG_2__SCAN_IN), .B(keyinput_249), .Z(n4862) );
  OAI21_X1 U5267 ( .B1(n4864), .B2(n4863), .A(n4862), .ZN(n4867) );
  XOR2_X1 U5268 ( .A(REG0_REG_4__SCAN_IN), .B(keyinput_251), .Z(n4866) );
  XOR2_X1 U5269 ( .A(REG0_REG_3__SCAN_IN), .B(keyinput_250), .Z(n4865) );
  NAND3_X1 U5270 ( .A1(n4867), .A2(n4866), .A3(n4865), .ZN(n4870) );
  XNOR2_X1 U5271 ( .A(REG0_REG_5__SCAN_IN), .B(keyinput_252), .ZN(n4869) );
  XOR2_X1 U5272 ( .A(REG0_REG_6__SCAN_IN), .B(keyinput_253), .Z(n4868) );
  AOI21_X1 U5273 ( .B1(n4870), .B2(n4869), .A(n4868), .ZN(n4873) );
  XOR2_X1 U5274 ( .A(REG0_REG_7__SCAN_IN), .B(keyinput_254), .Z(n4872) );
  XNOR2_X1 U5275 ( .A(keyinput_127), .B(keyinput_255), .ZN(n4871) );
  OAI21_X1 U5276 ( .B1(n4873), .B2(n4872), .A(n4871), .ZN(n4875) );
  XNOR2_X1 U5277 ( .A(REG0_REG_8__SCAN_IN), .B(keyinput_127), .ZN(n4874) );
  OAI211_X1 U5278 ( .C1(n4877), .C2(n4876), .A(n4875), .B(n4874), .ZN(n4878)
         );
  XNOR2_X1 U5279 ( .A(n4879), .B(n4878), .ZN(U3265) );
  XOR2_X1 U5280 ( .A(n4885), .B(n4880), .Z(n5024) );
  OAI22_X1 U5281 ( .A1(n4881), .A2(n5282), .B1(n5315), .B2(n4891), .ZN(n4888)
         );
  NOR2_X1 U5282 ( .A1(n4883), .A2(n4882), .ZN(n4884) );
  XOR2_X1 U5283 ( .A(n4885), .B(n4884), .Z(n4886) );
  NOR2_X1 U5284 ( .A1(n4886), .A2(n5288), .ZN(n4887) );
  AOI211_X1 U5285 ( .C1(n5286), .C2(n4889), .A(n4888), .B(n4887), .ZN(n5023)
         );
  INV_X1 U5286 ( .A(n5023), .ZN(n4896) );
  INV_X1 U5287 ( .A(n4911), .ZN(n4892) );
  OAI211_X1 U5288 ( .C1(n4892), .C2(n4891), .A(n5339), .B(n4890), .ZN(n5022)
         );
  AOI22_X1 U5289 ( .A1(n4893), .A2(n5303), .B1(n5333), .B2(
        REG2_REG_24__SCAN_IN), .ZN(n4894) );
  OAI21_X1 U5290 ( .B1(n5022), .B2(n4969), .A(n4894), .ZN(n4895) );
  AOI21_X1 U5291 ( .B1(n4896), .B2(n5138), .A(n4895), .ZN(n4897) );
  OAI21_X1 U5292 ( .B1(n5024), .B2(n5307), .A(n4897), .ZN(U3266) );
  OAI21_X1 U5293 ( .B1(n4899), .B2(n4904), .A(n4898), .ZN(n4900) );
  INV_X1 U5294 ( .A(n4900), .ZN(n5027) );
  OAI22_X1 U5295 ( .A1(n4940), .A2(n5282), .B1(n4912), .B2(n5315), .ZN(n4908)
         );
  AOI21_X1 U5296 ( .B1(n4937), .B2(n4902), .A(n4901), .ZN(n4926) );
  INV_X1 U5297 ( .A(n4919), .ZN(n4927) );
  NAND2_X1 U5298 ( .A1(n4926), .A2(n4927), .ZN(n4925) );
  NAND2_X1 U5299 ( .A1(n4925), .A2(n4903), .ZN(n4905) );
  XNOR2_X1 U5300 ( .A(n4905), .B(n4904), .ZN(n4906) );
  NOR2_X1 U5301 ( .A1(n4906), .A2(n5288), .ZN(n4907) );
  AOI211_X1 U5302 ( .C1(n5286), .C2(n4909), .A(n4908), .B(n4907), .ZN(n5026)
         );
  INV_X1 U5303 ( .A(n5026), .ZN(n4917) );
  OAI211_X1 U5304 ( .C1(n4910), .C2(n4912), .A(n5339), .B(n4911), .ZN(n5025)
         );
  INV_X1 U5305 ( .A(n4913), .ZN(n4914) );
  AOI22_X1 U5306 ( .A1(n4914), .A2(n5303), .B1(n5333), .B2(
        REG2_REG_23__SCAN_IN), .ZN(n4915) );
  OAI21_X1 U5307 ( .B1(n5025), .B2(n4969), .A(n4915), .ZN(n4916) );
  AOI21_X1 U5308 ( .B1(n4917), .B2(n5138), .A(n4916), .ZN(n4918) );
  OAI21_X1 U5309 ( .B1(n5027), .B2(n5307), .A(n4918), .ZN(U3267) );
  OAI21_X1 U5310 ( .B1(n4920), .B2(n4919), .A(n2518), .ZN(n5031) );
  INV_X1 U5311 ( .A(n4921), .ZN(n4943) );
  AOI21_X1 U5312 ( .B1(n4929), .B2(n4943), .A(n4910), .ZN(n5029) );
  INV_X1 U5313 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4923) );
  OAI22_X1 U5314 ( .A1(n5138), .A2(n4923), .B1(n4922), .B2(n4991), .ZN(n4924)
         );
  AOI21_X1 U5315 ( .B1(n5029), .B2(n5334), .A(n4924), .ZN(n4934) );
  OAI21_X1 U5316 ( .B1(n4927), .B2(n4926), .A(n4925), .ZN(n4928) );
  NAND2_X1 U5317 ( .A1(n4928), .A2(n5124), .ZN(n4932) );
  AOI22_X1 U5318 ( .A1(n4930), .A2(n5286), .B1(n5325), .B2(n4929), .ZN(n4931)
         );
  OAI211_X1 U5319 ( .C1(n4960), .C2(n5282), .A(n4932), .B(n4931), .ZN(n5028)
         );
  NAND2_X1 U5320 ( .A1(n5028), .A2(n5138), .ZN(n4933) );
  OAI211_X1 U5321 ( .C1(n5031), .C2(n5307), .A(n4934), .B(n4933), .ZN(U3268)
         );
  XOR2_X1 U5322 ( .A(n4936), .B(n4935), .Z(n5034) );
  XNOR2_X1 U5323 ( .A(n4937), .B(n4936), .ZN(n4942) );
  AOI22_X1 U5324 ( .A1(n4982), .A2(n4957), .B1(n4938), .B2(n5325), .ZN(n4939)
         );
  OAI21_X1 U5325 ( .B1(n4940), .B2(n5127), .A(n4939), .ZN(n4941) );
  AOI21_X1 U5326 ( .B1(n4942), .B2(n5124), .A(n4941), .ZN(n5033) );
  INV_X1 U5327 ( .A(n5033), .ZN(n4949) );
  INV_X1 U5328 ( .A(n4963), .ZN(n4945) );
  OAI211_X1 U5329 ( .C1(n4945), .C2(n4944), .A(n4943), .B(n5339), .ZN(n5032)
         );
  AOI22_X1 U5330 ( .A1(n5333), .A2(REG2_REG_21__SCAN_IN), .B1(n4946), .B2(
        n5303), .ZN(n4947) );
  OAI21_X1 U5331 ( .B1(n5032), .B2(n4969), .A(n4947), .ZN(n4948) );
  AOI21_X1 U5332 ( .B1(n4949), .B2(n5138), .A(n4948), .ZN(n4950) );
  OAI21_X1 U5333 ( .B1(n5034), .B2(n5307), .A(n4950), .ZN(U3269) );
  OAI21_X1 U5334 ( .B1(n4952), .B2(n4955), .A(n4951), .ZN(n4953) );
  INV_X1 U5335 ( .A(n4953), .ZN(n5037) );
  XOR2_X1 U5336 ( .A(n4955), .B(n4954), .Z(n4962) );
  AOI22_X1 U5337 ( .A1(n4958), .A2(n4957), .B1(n4956), .B2(n5325), .ZN(n4959)
         );
  OAI21_X1 U5338 ( .B1(n4960), .B2(n5127), .A(n4959), .ZN(n4961) );
  AOI21_X1 U5339 ( .B1(n4962), .B2(n5124), .A(n4961), .ZN(n5036) );
  INV_X1 U5340 ( .A(n5036), .ZN(n4971) );
  INV_X1 U5341 ( .A(n4987), .ZN(n4965) );
  OAI211_X1 U5342 ( .C1(n4965), .C2(n4964), .A(n5339), .B(n4963), .ZN(n5035)
         );
  INV_X1 U5343 ( .A(n4966), .ZN(n4967) );
  AOI22_X1 U5344 ( .A1(n5333), .A2(REG2_REG_20__SCAN_IN), .B1(n4967), .B2(
        n5303), .ZN(n4968) );
  OAI21_X1 U5345 ( .B1(n5035), .B2(n4969), .A(n4968), .ZN(n4970) );
  AOI21_X1 U5346 ( .B1(n4971), .B2(n5138), .A(n4970), .ZN(n4972) );
  OAI21_X1 U5347 ( .B1(n5037), .B2(n5307), .A(n4972), .ZN(U3270) );
  INV_X1 U5348 ( .A(n5138), .ZN(n5336) );
  OAI22_X1 U5349 ( .A1(n4973), .A2(n5282), .B1(n4988), .B2(n5315), .ZN(n4981)
         );
  INV_X1 U5350 ( .A(n4974), .ZN(n4975) );
  AOI21_X1 U5351 ( .B1(n4977), .B2(n4976), .A(n4975), .ZN(n4978) );
  XNOR2_X1 U5352 ( .A(n4978), .B(n2672), .ZN(n4979) );
  NOR2_X1 U5353 ( .A1(n4979), .A2(n5288), .ZN(n4980) );
  AOI211_X1 U5354 ( .C1(n5286), .C2(n4982), .A(n4981), .B(n4980), .ZN(n5039)
         );
  OAI21_X1 U5355 ( .B1(n4985), .B2(n4984), .A(n4983), .ZN(n5038) );
  NAND2_X1 U5356 ( .A1(n5038), .A2(n4986), .ZN(n4996) );
  OAI21_X1 U5357 ( .B1(n4989), .B2(n4988), .A(n4987), .ZN(n5041) );
  INV_X1 U5358 ( .A(n5041), .ZN(n4994) );
  INV_X1 U5359 ( .A(n4990), .ZN(n4992) );
  OAI22_X1 U5360 ( .A1(n5138), .A2(n2814), .B1(n4992), .B2(n4991), .ZN(n4993)
         );
  AOI21_X1 U5361 ( .B1(n4994), .B2(n5334), .A(n4993), .ZN(n4995) );
  OAI211_X1 U5362 ( .C1(n5336), .C2(n5039), .A(n4996), .B(n4995), .ZN(U3271)
         );
  NOR2_X1 U5363 ( .A1(n2961), .A2(n4997), .ZN(n4998) );
  NAND2_X1 U5364 ( .A1(n4998), .A2(n2997), .ZN(n5156) );
  NAND2_X1 U5365 ( .A1(n5000), .A2(n5258), .ZN(n5004) );
  NOR2_X2 U5366 ( .A1(n5002), .A2(n5001), .ZN(n5003) );
  NAND2_X1 U5367 ( .A1(n5004), .A2(n5003), .ZN(n5051) );
  NAND2_X1 U5368 ( .A1(n5006), .A2(n5005), .ZN(n5007) );
  AND2_X2 U5369 ( .A1(n5050), .A2(n5009), .ZN(n5343) );
  MUX2_X1 U5370 ( .A(REG1_REG_29__SCAN_IN), .B(n5051), .S(n5343), .Z(U3547) );
  MUX2_X1 U5371 ( .A(REG1_REG_28__SCAN_IN), .B(n5052), .S(n5343), .Z(U3546) );
  OAI211_X1 U5372 ( .C1(n5014), .C2(n5297), .A(n2492), .B(n5012), .ZN(n5053)
         );
  MUX2_X1 U5373 ( .A(REG1_REG_27__SCAN_IN), .B(n5053), .S(n5343), .Z(U3545) );
  OAI211_X1 U5374 ( .C1(n5017), .C2(n5297), .A(n5016), .B(n5015), .ZN(n5054)
         );
  MUX2_X1 U5375 ( .A(REG1_REG_26__SCAN_IN), .B(n5054), .S(n5343), .Z(U3544) );
  AOI21_X1 U5376 ( .B1(n5339), .B2(n5019), .A(n5018), .ZN(n5020) );
  OAI21_X1 U5377 ( .B1(n5021), .B2(n5297), .A(n5020), .ZN(n5055) );
  MUX2_X1 U5378 ( .A(REG1_REG_25__SCAN_IN), .B(n5055), .S(n5343), .Z(U3543) );
  OAI211_X1 U5379 ( .C1(n5024), .C2(n5297), .A(n5023), .B(n5022), .ZN(n5056)
         );
  MUX2_X1 U5380 ( .A(REG1_REG_24__SCAN_IN), .B(n5056), .S(n5343), .Z(U3542) );
  OAI211_X1 U5381 ( .C1(n5027), .C2(n5297), .A(n5026), .B(n5025), .ZN(n5057)
         );
  MUX2_X1 U5382 ( .A(REG1_REG_23__SCAN_IN), .B(n5057), .S(n5343), .Z(U3541) );
  AOI21_X1 U5383 ( .B1(n5339), .B2(n5029), .A(n5028), .ZN(n5030) );
  OAI21_X1 U5384 ( .B1(n5031), .B2(n5297), .A(n5030), .ZN(n5058) );
  MUX2_X1 U5385 ( .A(REG1_REG_22__SCAN_IN), .B(n5058), .S(n5343), .Z(U3540) );
  OAI211_X1 U5386 ( .C1(n5034), .C2(n5297), .A(n5033), .B(n5032), .ZN(n5059)
         );
  MUX2_X1 U5387 ( .A(REG1_REG_21__SCAN_IN), .B(n5059), .S(n5343), .Z(U3539) );
  OAI211_X1 U5388 ( .C1(n5037), .C2(n5297), .A(n5036), .B(n5035), .ZN(n5060)
         );
  MUX2_X1 U5389 ( .A(REG1_REG_20__SCAN_IN), .B(n5060), .S(n5343), .Z(U3538) );
  NAND2_X1 U5390 ( .A1(n5038), .A2(n5258), .ZN(n5040) );
  OAI211_X1 U5391 ( .C1(n5296), .C2(n5041), .A(n5040), .B(n5039), .ZN(n5061)
         );
  MUX2_X1 U5392 ( .A(REG1_REG_19__SCAN_IN), .B(n5061), .S(n5343), .Z(U3537) );
  OAI211_X1 U5393 ( .C1(n5044), .C2(n5297), .A(n5043), .B(n5042), .ZN(n5062)
         );
  MUX2_X1 U5394 ( .A(REG1_REG_18__SCAN_IN), .B(n5062), .S(n5343), .Z(U3536) );
  NAND2_X1 U5395 ( .A1(n5045), .A2(n5258), .ZN(n5047) );
  OAI211_X1 U5396 ( .C1(n5296), .C2(n5048), .A(n5047), .B(n5046), .ZN(n5063)
         );
  MUX2_X1 U5397 ( .A(REG1_REG_17__SCAN_IN), .B(n5063), .S(n5343), .Z(U3535) );
  MUX2_X1 U5398 ( .A(REG0_REG_29__SCAN_IN), .B(n5051), .S(n5347), .Z(U3515) );
  MUX2_X1 U5399 ( .A(REG0_REG_28__SCAN_IN), .B(n5052), .S(n5347), .Z(U3514) );
  MUX2_X1 U5400 ( .A(REG0_REG_27__SCAN_IN), .B(n5053), .S(n5347), .Z(U3513) );
  MUX2_X1 U5401 ( .A(REG0_REG_26__SCAN_IN), .B(n5054), .S(n5347), .Z(U3512) );
  MUX2_X1 U5402 ( .A(REG0_REG_25__SCAN_IN), .B(n5055), .S(n5347), .Z(U3511) );
  MUX2_X1 U5403 ( .A(REG0_REG_24__SCAN_IN), .B(n5056), .S(n5347), .Z(U3510) );
  MUX2_X1 U5404 ( .A(REG0_REG_23__SCAN_IN), .B(n5057), .S(n5347), .Z(U3509) );
  MUX2_X1 U5405 ( .A(REG0_REG_22__SCAN_IN), .B(n5058), .S(n5347), .Z(U3508) );
  MUX2_X1 U5406 ( .A(REG0_REG_21__SCAN_IN), .B(n5059), .S(n5347), .Z(U3507) );
  MUX2_X1 U5407 ( .A(REG0_REG_20__SCAN_IN), .B(n5060), .S(n5347), .Z(U3506) );
  MUX2_X1 U5408 ( .A(REG0_REG_19__SCAN_IN), .B(n5061), .S(n5347), .Z(U3505) );
  MUX2_X1 U5409 ( .A(REG0_REG_18__SCAN_IN), .B(n5062), .S(n5347), .Z(U3503) );
  MUX2_X1 U5410 ( .A(REG0_REG_17__SCAN_IN), .B(n5063), .S(n5347), .Z(U3501) );
  NOR3_X1 U5411 ( .A1(n2921), .A2(IR_REG_30__SCAN_IN), .A3(n5064), .ZN(n5065)
         );
  MUX2_X1 U5412 ( .A(DATAI_31_), .B(n5065), .S(STATE_REG_SCAN_IN), .Z(U3321)
         );
  MUX2_X1 U5413 ( .A(DATAI_30_), .B(n5066), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U5414 ( .A(n5067), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5415 ( .A(n5068), .B(DATAI_28_), .S(U3149), .Z(U3324) );
  MUX2_X1 U5416 ( .A(DATAI_26_), .B(n5069), .S(STATE_REG_SCAN_IN), .Z(U3326)
         );
  INV_X1 U5417 ( .A(n2908), .ZN(n5070) );
  MUX2_X1 U5418 ( .A(n5070), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5419 ( .A(n5071), .B(DATAI_18_), .S(U3149), .Z(U3334) );
  MUX2_X1 U5420 ( .A(n5072), .B(DATAI_17_), .S(U3149), .Z(U3335) );
  MUX2_X1 U5421 ( .A(n5073), .B(DATAI_15_), .S(U3149), .Z(U3337) );
  MUX2_X1 U5422 ( .A(DATAI_8_), .B(n5074), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5423 ( .A(n2848), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5424 ( .A(n2850), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  NOR2_X1 U5425 ( .A1(n5099), .A2(n5075), .ZN(U3320) );
  NOR2_X1 U5426 ( .A1(n5099), .A2(n5076), .ZN(U3319) );
  AND2_X1 U5427 ( .A1(n5095), .A2(D_REG_4__SCAN_IN), .ZN(U3318) );
  NOR2_X1 U5428 ( .A1(n5099), .A2(n5077), .ZN(U3317) );
  NOR2_X1 U5429 ( .A1(n5099), .A2(n5078), .ZN(U3316) );
  AND2_X1 U5430 ( .A1(n5095), .A2(D_REG_7__SCAN_IN), .ZN(U3315) );
  NOR2_X1 U5431 ( .A1(n5099), .A2(n5079), .ZN(U3314) );
  INV_X1 U5432 ( .A(D_REG_9__SCAN_IN), .ZN(n5080) );
  NOR2_X1 U5433 ( .A1(n5099), .A2(n5080), .ZN(U3313) );
  NOR2_X1 U5434 ( .A1(n5099), .A2(n5081), .ZN(U3312) );
  NOR2_X1 U5435 ( .A1(n5099), .A2(n5082), .ZN(U3311) );
  NOR2_X1 U5436 ( .A1(n5099), .A2(n5083), .ZN(U3310) );
  NOR2_X1 U5437 ( .A1(n5099), .A2(n5084), .ZN(U3309) );
  AND2_X1 U5438 ( .A1(n5095), .A2(D_REG_14__SCAN_IN), .ZN(U3308) );
  INV_X1 U5439 ( .A(D_REG_15__SCAN_IN), .ZN(n5085) );
  NOR2_X1 U5440 ( .A1(n5099), .A2(n5085), .ZN(U3307) );
  NOR2_X1 U5441 ( .A1(n5099), .A2(n5086), .ZN(U3306) );
  NOR2_X1 U5442 ( .A1(n5099), .A2(n5087), .ZN(U3305) );
  INV_X1 U5443 ( .A(D_REG_18__SCAN_IN), .ZN(n5088) );
  NOR2_X1 U5444 ( .A1(n5099), .A2(n5088), .ZN(U3304) );
  NOR2_X1 U5445 ( .A1(n5099), .A2(n5089), .ZN(U3303) );
  AND2_X1 U5446 ( .A1(n5095), .A2(D_REG_20__SCAN_IN), .ZN(U3302) );
  NOR2_X1 U5447 ( .A1(n5099), .A2(n5090), .ZN(U3301) );
  INV_X1 U5448 ( .A(D_REG_22__SCAN_IN), .ZN(n5091) );
  NOR2_X1 U5449 ( .A1(n5099), .A2(n5091), .ZN(U3300) );
  NOR2_X1 U5450 ( .A1(n5099), .A2(n5092), .ZN(U3299) );
  AND2_X1 U5451 ( .A1(n5095), .A2(D_REG_24__SCAN_IN), .ZN(U3298) );
  AND2_X1 U5452 ( .A1(n5095), .A2(D_REG_25__SCAN_IN), .ZN(U3297) );
  NOR2_X1 U5453 ( .A1(n5099), .A2(n5093), .ZN(U3296) );
  NOR2_X1 U5454 ( .A1(n5099), .A2(n5094), .ZN(U3295) );
  AND2_X1 U5455 ( .A1(n5095), .A2(D_REG_28__SCAN_IN), .ZN(U3294) );
  NOR2_X1 U5456 ( .A1(n5099), .A2(n5096), .ZN(U3293) );
  NOR2_X1 U5457 ( .A1(n5099), .A2(n5097), .ZN(U3292) );
  NOR2_X1 U5458 ( .A1(n5099), .A2(n5098), .ZN(U3291) );
  AOI21_X1 U5459 ( .B1(n2965), .B2(n2846), .A(n5100), .ZN(n5101) );
  XNOR2_X1 U5460 ( .A(n5101), .B(IR_REG_0__SCAN_IN), .ZN(n5103) );
  AOI22_X1 U5461 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n5107), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n5102) );
  OAI21_X1 U5462 ( .B1(n5104), .B2(n5103), .A(n5102), .ZN(U3240) );
  INV_X1 U5463 ( .A(DATAI_0_), .ZN(n5105) );
  AOI22_X1 U5464 ( .A1(STATE_REG_SCAN_IN), .A2(n2572), .B1(n5105), .B2(U3149), 
        .ZN(U3352) );
  AOI21_X1 U5465 ( .B1(n5107), .B2(ADDR_REG_4__SCAN_IN), .A(n5106), .ZN(n5120)
         );
  AOI211_X1 U5466 ( .C1(n5110), .C2(n5170), .A(n5109), .B(n5108), .ZN(n5112)
         );
  AOI211_X1 U5467 ( .C1(n5114), .C2(n5113), .A(n5112), .B(n5111), .ZN(n5119)
         );
  OAI211_X1 U5468 ( .C1(REG2_REG_4__SCAN_IN), .C2(n5117), .A(n5116), .B(n5115), 
        .ZN(n5118) );
  NAND3_X1 U5469 ( .A1(n5120), .A2(n5119), .A3(n5118), .ZN(U3244) );
  INV_X1 U5470 ( .A(n5156), .ZN(n5168) );
  INV_X1 U5471 ( .A(n5121), .ZN(n5122) );
  NOR2_X1 U5472 ( .A1(n5123), .A2(n5122), .ZN(n5133) );
  OAI21_X1 U5473 ( .B1(n5125), .B2(n5124), .A(n5135), .ZN(n5126) );
  OAI21_X1 U5474 ( .B1(n3199), .B2(n5127), .A(n5126), .ZN(n5131) );
  AOI211_X1 U5475 ( .C1(n5168), .C2(n5135), .A(n5133), .B(n5131), .ZN(n5129)
         );
  AOI22_X1 U5476 ( .A1(n5343), .A2(n5129), .B1(n2965), .B2(n5341), .ZN(U3518)
         );
  INV_X1 U5477 ( .A(REG0_REG_0__SCAN_IN), .ZN(n5128) );
  AOI22_X1 U5478 ( .A1(n5347), .A2(n5129), .B1(n5128), .B2(n5344), .ZN(U3467)
         );
  NAND2_X1 U5479 ( .A1(n2997), .A2(n5130), .ZN(n5132) );
  AOI21_X1 U5480 ( .B1(n5133), .B2(n5132), .A(n5131), .ZN(n5139) );
  INV_X1 U5481 ( .A(REG2_REG_0__SCAN_IN), .ZN(n5137) );
  AOI22_X1 U5482 ( .A1(n5135), .A2(n5134), .B1(REG3_REG_0__SCAN_IN), .B2(n5303), .ZN(n5136) );
  OAI221_X1 U5483 ( .B1(n5336), .B2(n5139), .C1(n5138), .C2(n5137), .A(n5136), 
        .ZN(U3290) );
  INV_X1 U5484 ( .A(n5140), .ZN(n5144) );
  INV_X1 U5485 ( .A(n5141), .ZN(n5142) );
  AOI211_X1 U5486 ( .C1(n5144), .C2(n5168), .A(n5143), .B(n5142), .ZN(n5146)
         );
  AOI22_X1 U5487 ( .A1(n5343), .A2(n5146), .B1(n2849), .B2(n5341), .ZN(U3519)
         );
  INV_X1 U5488 ( .A(REG0_REG_1__SCAN_IN), .ZN(n5145) );
  AOI22_X1 U5489 ( .A1(n5347), .A2(n5146), .B1(n5145), .B2(n5344), .ZN(U3469)
         );
  NOR2_X1 U5490 ( .A1(n5147), .A2(n5156), .ZN(n5150) );
  INV_X1 U5491 ( .A(n5148), .ZN(n5149) );
  AOI211_X1 U5492 ( .C1(n5339), .C2(n5151), .A(n5150), .B(n5149), .ZN(n5153)
         );
  AOI22_X1 U5493 ( .A1(n5343), .A2(n5153), .B1(n2847), .B2(n5341), .ZN(U3520)
         );
  INV_X1 U5494 ( .A(REG0_REG_2__SCAN_IN), .ZN(n5152) );
  AOI22_X1 U5495 ( .A1(n5347), .A2(n5153), .B1(n5152), .B2(n5344), .ZN(U3471)
         );
  INV_X1 U5496 ( .A(DATAI_3_), .ZN(n5154) );
  AOI22_X1 U5497 ( .A1(STATE_REG_SCAN_IN), .A2(n2588), .B1(n5154), .B2(U3149), 
        .ZN(U3349) );
  OAI22_X1 U5498 ( .A1(n5157), .A2(n5156), .B1(n5296), .B2(n5155), .ZN(n5158)
         );
  NOR2_X1 U5499 ( .A1(n5159), .A2(n5158), .ZN(n5162) );
  AOI22_X1 U5500 ( .A1(n5343), .A2(n5162), .B1(n5160), .B2(n5341), .ZN(U3521)
         );
  INV_X1 U5501 ( .A(REG0_REG_3__SCAN_IN), .ZN(n5161) );
  AOI22_X1 U5502 ( .A1(n5347), .A2(n5162), .B1(n5161), .B2(n5344), .ZN(U3473)
         );
  AOI22_X1 U5503 ( .A1(STATE_REG_SCAN_IN), .A2(n5164), .B1(n5163), .B2(U3149), 
        .ZN(U3348) );
  INV_X1 U5504 ( .A(n5165), .ZN(n5166) );
  AOI211_X1 U5505 ( .C1(n5169), .C2(n5168), .A(n5167), .B(n5166), .ZN(n5172)
         );
  AOI22_X1 U5506 ( .A1(n5343), .A2(n5172), .B1(n5170), .B2(n5341), .ZN(U3522)
         );
  INV_X1 U5507 ( .A(REG0_REG_4__SCAN_IN), .ZN(n5171) );
  AOI22_X1 U5508 ( .A1(n5347), .A2(n5172), .B1(n5171), .B2(n5344), .ZN(U3475)
         );
  AOI22_X1 U5509 ( .A1(STATE_REG_SCAN_IN), .A2(n5174), .B1(n5173), .B2(U3149), 
        .ZN(U3347) );
  NOR2_X1 U5510 ( .A1(n5175), .A2(n5296), .ZN(n5177) );
  AOI211_X1 U5511 ( .C1(n5178), .C2(n5258), .A(n5177), .B(n5176), .ZN(n5181)
         );
  INV_X1 U5512 ( .A(REG1_REG_5__SCAN_IN), .ZN(n5179) );
  AOI22_X1 U5513 ( .A1(n5343), .A2(n5181), .B1(n5179), .B2(n5341), .ZN(U3523)
         );
  INV_X1 U5514 ( .A(REG0_REG_5__SCAN_IN), .ZN(n5180) );
  AOI22_X1 U5515 ( .A1(n5347), .A2(n5181), .B1(n5180), .B2(n5344), .ZN(U3477)
         );
  INV_X1 U5516 ( .A(DATAI_6_), .ZN(n5182) );
  AOI22_X1 U5517 ( .A1(STATE_REG_SCAN_IN), .A2(n5183), .B1(n5182), .B2(U3149), 
        .ZN(U3346) );
  AOI211_X1 U5518 ( .C1(n5186), .C2(n5258), .A(n5185), .B(n5184), .ZN(n5189)
         );
  AOI22_X1 U5519 ( .A1(n5343), .A2(n5189), .B1(n5187), .B2(n5341), .ZN(U3524)
         );
  INV_X1 U5520 ( .A(REG0_REG_6__SCAN_IN), .ZN(n5188) );
  AOI22_X1 U5521 ( .A1(n5347), .A2(n5189), .B1(n5188), .B2(n5344), .ZN(U3479)
         );
  AOI22_X1 U5522 ( .A1(STATE_REG_SCAN_IN), .A2(n5191), .B1(n5190), .B2(U3149), 
        .ZN(U3345) );
  NAND3_X1 U5523 ( .A1(n3285), .A2(n5192), .A3(n5258), .ZN(n5193) );
  AND3_X1 U5524 ( .A1(n5195), .A2(n5194), .A3(n5193), .ZN(n5197) );
  AOI22_X1 U5525 ( .A1(n5343), .A2(n5197), .B1(n2861), .B2(n5341), .ZN(U3525)
         );
  INV_X1 U5526 ( .A(REG0_REG_7__SCAN_IN), .ZN(n5196) );
  AOI22_X1 U5527 ( .A1(n5347), .A2(n5197), .B1(n5196), .B2(n5344), .ZN(U3481)
         );
  OAI22_X1 U5528 ( .A1(n5199), .A2(n5297), .B1(n5296), .B2(n5198), .ZN(n5201)
         );
  NOR2_X1 U5529 ( .A1(n5201), .A2(n5200), .ZN(n5204) );
  INV_X1 U5530 ( .A(REG1_REG_8__SCAN_IN), .ZN(n5202) );
  AOI22_X1 U5531 ( .A1(n5343), .A2(n5204), .B1(n5202), .B2(n5341), .ZN(U3526)
         );
  INV_X1 U5532 ( .A(REG0_REG_8__SCAN_IN), .ZN(n5203) );
  AOI22_X1 U5533 ( .A1(n5347), .A2(n5204), .B1(n5203), .B2(n5344), .ZN(U3483)
         );
  INV_X1 U5534 ( .A(DATAI_9_), .ZN(n5205) );
  AOI22_X1 U5535 ( .A1(STATE_REG_SCAN_IN), .A2(n5206), .B1(n5205), .B2(U3149), 
        .ZN(U3343) );
  NOR2_X1 U5536 ( .A1(n5207), .A2(n5297), .ZN(n5208) );
  AOI211_X1 U5537 ( .C1(n5339), .C2(n5210), .A(n5209), .B(n5208), .ZN(n5212)
         );
  AOI22_X1 U5538 ( .A1(n5343), .A2(n5212), .B1(n2866), .B2(n5341), .ZN(U3527)
         );
  INV_X1 U5539 ( .A(REG0_REG_9__SCAN_IN), .ZN(n5211) );
  AOI22_X1 U5540 ( .A1(n5347), .A2(n5212), .B1(n5211), .B2(n5344), .ZN(U3485)
         );
  AOI22_X1 U5541 ( .A1(STATE_REG_SCAN_IN), .A2(n2601), .B1(n5213), .B2(U3149), 
        .ZN(U3342) );
  OAI21_X1 U5542 ( .B1(n5296), .B2(n5215), .A(n5214), .ZN(n5216) );
  AOI21_X1 U5543 ( .B1(n5217), .B2(n5258), .A(n5216), .ZN(n5220) );
  AOI22_X1 U5544 ( .A1(n5343), .A2(n5220), .B1(n5218), .B2(n5341), .ZN(U3528)
         );
  INV_X1 U5545 ( .A(REG0_REG_10__SCAN_IN), .ZN(n5219) );
  AOI22_X1 U5546 ( .A1(n5347), .A2(n5220), .B1(n5219), .B2(n5344), .ZN(U3487)
         );
  AOI22_X1 U5547 ( .A1(STATE_REG_SCAN_IN), .A2(n5222), .B1(n5221), .B2(U3149), 
        .ZN(U3341) );
  OAI21_X1 U5548 ( .B1(n5296), .B2(n5224), .A(n5223), .ZN(n5225) );
  AOI21_X1 U5549 ( .B1(n5226), .B2(n5258), .A(n5225), .ZN(n5229) );
  INV_X1 U5550 ( .A(REG1_REG_11__SCAN_IN), .ZN(n5227) );
  AOI22_X1 U5551 ( .A1(n5343), .A2(n5229), .B1(n5227), .B2(n5341), .ZN(U3529)
         );
  INV_X1 U5552 ( .A(REG0_REG_11__SCAN_IN), .ZN(n5228) );
  AOI22_X1 U5553 ( .A1(n5347), .A2(n5229), .B1(n5228), .B2(n5344), .ZN(U3489)
         );
  INV_X1 U5554 ( .A(DATAI_12_), .ZN(n5230) );
  AOI22_X1 U5555 ( .A1(STATE_REG_SCAN_IN), .A2(n5231), .B1(n5230), .B2(U3149), 
        .ZN(U3340) );
  NOR2_X1 U5556 ( .A1(n5232), .A2(n5296), .ZN(n5234) );
  AOI211_X1 U5557 ( .C1(n5235), .C2(n5258), .A(n5234), .B(n5233), .ZN(n5238)
         );
  AOI22_X1 U5558 ( .A1(n5343), .A2(n5238), .B1(n5236), .B2(n5341), .ZN(U3530)
         );
  INV_X1 U5559 ( .A(REG0_REG_12__SCAN_IN), .ZN(n5237) );
  AOI22_X1 U5560 ( .A1(n5347), .A2(n5238), .B1(n5237), .B2(n5344), .ZN(U3491)
         );
  AOI22_X1 U5561 ( .A1(STATE_REG_SCAN_IN), .A2(n5240), .B1(n5239), .B2(U3149), 
        .ZN(U3339) );
  NOR2_X1 U5562 ( .A1(n5241), .A2(n5297), .ZN(n5242) );
  AOI211_X1 U5563 ( .C1(n5339), .C2(n5244), .A(n5243), .B(n5242), .ZN(n5247)
         );
  INV_X1 U5564 ( .A(REG1_REG_13__SCAN_IN), .ZN(n5245) );
  AOI22_X1 U5565 ( .A1(n5343), .A2(n5247), .B1(n5245), .B2(n5341), .ZN(U3531)
         );
  INV_X1 U5566 ( .A(REG0_REG_13__SCAN_IN), .ZN(n5246) );
  AOI22_X1 U5567 ( .A1(n5347), .A2(n5247), .B1(n5246), .B2(n5344), .ZN(U3493)
         );
  INV_X1 U5568 ( .A(DATAI_14_), .ZN(n5248) );
  AOI22_X1 U5569 ( .A1(STATE_REG_SCAN_IN), .A2(n2587), .B1(n5248), .B2(U3149), 
        .ZN(U3338) );
  AOI211_X1 U5570 ( .C1(n5251), .C2(n5258), .A(n5250), .B(n5249), .ZN(n5254)
         );
  AOI22_X1 U5571 ( .A1(n5343), .A2(n5254), .B1(n5252), .B2(n5341), .ZN(U3532)
         );
  INV_X1 U5572 ( .A(REG0_REG_14__SCAN_IN), .ZN(n5253) );
  AOI22_X1 U5573 ( .A1(n5347), .A2(n5254), .B1(n5253), .B2(n5344), .ZN(U3495)
         );
  OAI21_X1 U5574 ( .B1(n5296), .B2(n5256), .A(n5255), .ZN(n5257) );
  AOI21_X1 U5575 ( .B1(n5259), .B2(n5258), .A(n5257), .ZN(n5262) );
  AOI22_X1 U5576 ( .A1(n5343), .A2(n5262), .B1(n5260), .B2(n5341), .ZN(U3533)
         );
  INV_X1 U5577 ( .A(REG0_REG_15__SCAN_IN), .ZN(n5261) );
  AOI22_X1 U5578 ( .A1(n5347), .A2(n5262), .B1(n5261), .B2(n5344), .ZN(U3497)
         );
  INV_X1 U5579 ( .A(DATAI_16_), .ZN(n5263) );
  AOI22_X1 U5580 ( .A1(STATE_REG_SCAN_IN), .A2(n5264), .B1(n5263), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5581 ( .A(n5304), .ZN(n5279) );
  AOI22_X1 U5582 ( .A1(n5268), .A2(n5267), .B1(n5266), .B2(n5265), .ZN(n5278)
         );
  NAND2_X1 U5583 ( .A1(n5269), .A2(n5270), .ZN(n5272) );
  AOI21_X1 U5584 ( .B1(n5273), .B2(n5272), .A(n5271), .ZN(n5274) );
  AOI211_X1 U5585 ( .C1(n5276), .C2(n5285), .A(n5275), .B(n5274), .ZN(n5277)
         );
  OAI211_X1 U5586 ( .C1(n5280), .C2(n5279), .A(n5278), .B(n5277), .ZN(U3223)
         );
  XNOR2_X1 U5587 ( .A(n5281), .B(n5290), .ZN(n5289) );
  OAI22_X1 U5588 ( .A1(n5283), .A2(n5282), .B1(n5294), .B2(n5315), .ZN(n5284)
         );
  AOI21_X1 U5589 ( .B1(n5286), .B2(n5285), .A(n5284), .ZN(n5287) );
  OAI21_X1 U5590 ( .B1(n5289), .B2(n5288), .A(n5287), .ZN(n5302) );
  XNOR2_X1 U5591 ( .A(n5291), .B(n5290), .ZN(n5308) );
  INV_X1 U5592 ( .A(n5292), .ZN(n5295) );
  OAI21_X1 U5593 ( .B1(n5295), .B2(n5294), .A(n5293), .ZN(n5305) );
  OAI22_X1 U5594 ( .A1(n5308), .A2(n5297), .B1(n5296), .B2(n5305), .ZN(n5298)
         );
  NOR2_X1 U5595 ( .A1(n5302), .A2(n5298), .ZN(n5301) );
  AOI22_X1 U5596 ( .A1(n5343), .A2(n5301), .B1(n5299), .B2(n5341), .ZN(U3534)
         );
  INV_X1 U5597 ( .A(REG0_REG_16__SCAN_IN), .ZN(n5300) );
  AOI22_X1 U5598 ( .A1(n5347), .A2(n5301), .B1(n5300), .B2(n5344), .ZN(U3499)
         );
  AOI21_X1 U5599 ( .B1(n5304), .B2(n5303), .A(n5302), .ZN(n5311) );
  OAI22_X1 U5600 ( .A1(n5308), .A2(n5307), .B1(n5306), .B2(n5305), .ZN(n5309)
         );
  AOI21_X1 U5601 ( .B1(n5336), .B2(REG2_REG_16__SCAN_IN), .A(n5309), .ZN(n5310) );
  OAI21_X1 U5602 ( .B1(n5311), .B2(n5336), .A(n5310), .ZN(U3274) );
  INV_X1 U5603 ( .A(n5312), .ZN(n5313) );
  NAND2_X1 U5604 ( .A1(n5314), .A2(n5313), .ZN(n5328) );
  OR2_X1 U5605 ( .A1(n5329), .A2(n5315), .ZN(n5316) );
  AND2_X1 U5606 ( .A1(n5328), .A2(n5316), .ZN(n5319) );
  XNOR2_X1 U5607 ( .A(n5330), .B(n5317), .ZN(n5321) );
  AOI22_X1 U5608 ( .A1(n5321), .A2(n5334), .B1(REG2_REG_30__SCAN_IN), .B2(
        n5333), .ZN(n5318) );
  OAI21_X1 U5609 ( .B1(n5336), .B2(n5319), .A(n5318), .ZN(U3261) );
  INV_X1 U5610 ( .A(n5319), .ZN(n5320) );
  AOI21_X1 U5611 ( .B1(n5321), .B2(n5339), .A(n5320), .ZN(n5324) );
  INV_X1 U5612 ( .A(REG1_REG_30__SCAN_IN), .ZN(n5322) );
  AOI22_X1 U5613 ( .A1(n5343), .A2(n5324), .B1(n5322), .B2(n5341), .ZN(U3548)
         );
  INV_X1 U5614 ( .A(REG0_REG_30__SCAN_IN), .ZN(n5323) );
  AOI22_X1 U5615 ( .A1(n5347), .A2(n5324), .B1(n5323), .B2(n5344), .ZN(U3516)
         );
  NAND2_X1 U5616 ( .A1(n5326), .A2(n5325), .ZN(n5327) );
  AND2_X1 U5617 ( .A1(n5328), .A2(n5327), .ZN(n5337) );
  NAND2_X1 U5618 ( .A1(n5330), .A2(n5329), .ZN(n5332) );
  XNOR2_X1 U5619 ( .A(n5332), .B(n5331), .ZN(n5340) );
  AOI22_X1 U5620 ( .A1(n5340), .A2(n5334), .B1(n5333), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n5335) );
  OAI21_X1 U5621 ( .B1(n5336), .B2(n5337), .A(n5335), .ZN(U3260) );
  INV_X1 U5622 ( .A(n5337), .ZN(n5338) );
  AOI21_X1 U5623 ( .B1(n5340), .B2(n5339), .A(n5338), .ZN(n5346) );
  INV_X1 U5624 ( .A(REG1_REG_31__SCAN_IN), .ZN(n5342) );
  AOI22_X1 U5625 ( .A1(n5343), .A2(n5346), .B1(n5342), .B2(n5341), .ZN(U3549)
         );
  INV_X1 U5626 ( .A(REG0_REG_31__SCAN_IN), .ZN(n5345) );
  AOI22_X1 U5627 ( .A1(n5347), .A2(n5346), .B1(n5345), .B2(n5344), .ZN(U3517)
         );
  CLKBUF_X1 U2541 ( .A(n2845), .Z(n2495) );
endmodule

