

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput127, keyinput126,
         keyinput125, keyinput124, keyinput123, keyinput122, keyinput121,
         keyinput120, keyinput119, keyinput118, keyinput117, keyinput116,
         keyinput115, keyinput114, keyinput113, keyinput112, keyinput111,
         keyinput110, keyinput109, keyinput108, keyinput107, keyinput106,
         keyinput105, keyinput104, keyinput103, keyinput102, keyinput101,
         keyinput100, keyinput99, keyinput98, keyinput97, keyinput96,
         keyinput95, keyinput94, keyinput93, keyinput92, keyinput91,
         keyinput90, keyinput89, keyinput88, keyinput87, keyinput86,
         keyinput85, keyinput84, keyinput83, keyinput82, keyinput81,
         keyinput80, keyinput79, keyinput78, keyinput77, keyinput76,
         keyinput75, keyinput74, keyinput73, keyinput72, keyinput71,
         keyinput70, keyinput69, keyinput68, keyinput67, keyinput66,
         keyinput65, keyinput64, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901;

  AOI21_X1 U3539 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n6870), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3654) );
  AND2_X1 U3540 ( .A1(n4498), .A2(n4499), .ZN(n4496) );
  NAND2_X1 U3541 ( .A1(n3383), .A2(n3382), .ZN(n3418) );
  OAI21_X1 U3542 ( .B1(n3494), .B2(n3135), .A(n3133), .ZN(n3383) );
  CLKBUF_X2 U3543 ( .A(n3346), .Z(n4008) );
  CLKBUF_X2 U3544 ( .A(n3384), .Z(n4007) );
  BUF_X2 U3545 ( .A(n3368), .Z(n3985) );
  CLKBUF_X2 U3546 ( .A(n3349), .Z(n4013) );
  BUF_X2 U3547 ( .A(n3302), .Z(n3999) );
  CLKBUF_X2 U3548 ( .A(n3367), .Z(n3984) );
  CLKBUF_X2 U3549 ( .A(n3360), .Z(n3348) );
  CLKBUF_X2 U3550 ( .A(n3288), .Z(n4002) );
  BUF_X1 U3551 ( .A(n3317), .Z(n5139) );
  AND2_X1 U3552 ( .A1(n4034), .A2(n3376), .ZN(n4068) );
  NAND4_X1 U3553 ( .A1(n6872), .A2(n3153), .A3(n6871), .A4(n6870), .ZN(n6880)
         );
  NAND2_X1 U3554 ( .A1(n4226), .A2(n4225), .ZN(n6098) );
  XNOR2_X1 U3555 ( .A(n3418), .B(n3416), .ZN(n3482) );
  OAI221_X1 U3556 ( .B1(n6757), .B2(keyinput0), .C1(n6756), .C2(keyinput28), 
        .A(n6755), .ZN(n6764) );
  INV_X1 U3558 ( .A(n5044), .ZN(n5998) );
  INV_X1 U3559 ( .A(n3296), .ZN(n4189) );
  INV_X1 U3560 ( .A(n4207), .ZN(n4623) );
  AND2_X2 U3561 ( .A1(n3099), .A2(n4510), .ZN(n4373) );
  AND2_X1 U3562 ( .A1(n6078), .A2(n4423), .ZN(n6097) );
  INV_X1 U3563 ( .A(n6006), .ZN(n5993) );
  AND3_X1 U3564 ( .A1(n3505), .A2(n4443), .A3(n4444), .ZN(n3091) );
  OR2_X2 U3565 ( .A1(n5310), .A2(n5120), .ZN(n5121) );
  AND4_X4 U3566 ( .A1(n3227), .A2(n3226), .A3(n3225), .A4(n3224), .ZN(n3403)
         );
  AND4_X2 U3567 ( .A1(n3223), .A2(n3222), .A3(n3221), .A4(n3220), .ZN(n3224)
         );
  NAND3_X4 U3568 ( .A1(n3275), .A2(n3274), .A3(n3273), .ZN(n3339) );
  XNOR2_X2 U3569 ( .A(n3549), .B(n3550), .ZN(n4235) );
  NOR2_X2 U3570 ( .A1(n3549), .A2(n3553), .ZN(n3578) );
  NOR2_X2 U3571 ( .A1(n5700), .A2(n5701), .ZN(n5699) );
  AND2_X4 U3572 ( .A1(n3407), .A2(n3099), .ZN(n4202) );
  BUF_X4 U3573 ( .A(n3340), .Z(n3099) );
  AND2_X4 U3575 ( .A1(n4048), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3201)
         );
  NAND2_X2 U3576 ( .A1(n3467), .A2(n3468), .ZN(n3549) );
  INV_X4 U3577 ( .A(n5716), .ZN(n5557) );
  AOI22_X2 U3578 ( .A1(n6099), .A2(n4228), .B1(n4227), .B2(n6181), .ZN(n4842)
         );
  INV_X2 U3579 ( .A(n5842), .ZN(n5964) );
  NAND2_X1 U3580 ( .A1(n6588), .A2(n4352), .ZN(n5044) );
  OR2_X1 U3581 ( .A1(n3374), .A2(n3373), .ZN(n4264) );
  NOR2_X1 U3582 ( .A1(n4084), .A2(n4623), .ZN(n3095) );
  OR2_X1 U3583 ( .A1(n4084), .A2(n4623), .ZN(n4213) );
  AND2_X1 U3584 ( .A1(n3264), .A2(n3263), .ZN(n3275) );
  INV_X1 U3585 ( .A(n3316), .ZN(n3493) );
  NAND2_X1 U3586 ( .A1(n3284), .A2(n3106), .ZN(n3340) );
  INV_X2 U3587 ( .A(n3390), .ZN(n4011) );
  CLKBUF_X2 U3588 ( .A(n3304), .Z(n4001) );
  BUF_X2 U3589 ( .A(n3347), .Z(n4009) );
  INV_X2 U3590 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3195) );
  XNOR2_X1 U3591 ( .A(n5153), .B(n5152), .ZN(n5196) );
  OR2_X1 U3592 ( .A1(n5310), .A2(n5309), .ZN(n5794) );
  AND2_X1 U3593 ( .A1(n3160), .A2(n3159), .ZN(n5444) );
  OAI21_X1 U3594 ( .B1(n4280), .B2(n3188), .A(n3154), .ZN(n5422) );
  NAND2_X1 U3595 ( .A1(n3908), .A2(n3907), .ZN(n5319) );
  NAND2_X1 U3596 ( .A1(n3148), .A2(n3145), .ZN(n5546) );
  NOR2_X1 U3597 ( .A1(n4610), .A2(n4609), .ZN(n3576) );
  NOR2_X1 U3598 ( .A1(n5268), .A2(n5281), .ZN(n5907) );
  AOI21_X1 U3599 ( .B1(n3547), .B2(n3708), .A(n3546), .ZN(n4655) );
  OR2_X1 U3600 ( .A1(n5983), .A2(n4358), .ZN(n5281) );
  AND2_X2 U3601 ( .A1(n4251), .A2(n4200), .ZN(n5716) );
  INV_X1 U3602 ( .A(n3468), .ZN(n4589) );
  OR2_X1 U3603 ( .A1(n5263), .A2(n4146), .ZN(n5362) );
  NOR2_X2 U3604 ( .A1(n6583), .A2(n5998), .ZN(n5024) );
  BUF_X2 U3605 ( .A(n4210), .Z(n4576) );
  INV_X1 U3606 ( .A(n5728), .ZN(n6226) );
  INV_X2 U3607 ( .A(n6023), .ZN(n3092) );
  AND2_X1 U3608 ( .A1(n4392), .A2(n4390), .ZN(n6588) );
  OR2_X1 U3609 ( .A1(n3886), .A2(n5072), .ZN(n3887) );
  NAND2_X1 U3610 ( .A1(n3446), .A2(n3445), .ZN(n4561) );
  NAND2_X1 U3611 ( .A1(n3111), .A2(n3489), .ZN(n3492) );
  AND2_X1 U3612 ( .A1(n3132), .A2(n3488), .ZN(n3111) );
  NOR2_X1 U3613 ( .A1(n3851), .A2(n6772), .ZN(n3853) );
  CLKBUF_X1 U3614 ( .A(n3494), .Z(n3102) );
  OR2_X1 U3615 ( .A1(n3803), .A2(n5829), .ZN(n3851) );
  AOI21_X1 U3616 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6586), .A(n4071), 
        .ZN(n4077) );
  AND2_X1 U3617 ( .A1(n3134), .A2(n3489), .ZN(n3133) );
  AND2_X1 U3618 ( .A1(n3297), .A2(n4524), .ZN(n3336) );
  NAND2_X1 U3619 ( .A1(n3453), .A2(n3452), .ZN(n4073) );
  INV_X2 U3620 ( .A(n4081), .ZN(n3296) );
  NOR2_X1 U3621 ( .A1(n4213), .A2(n5139), .ZN(n4292) );
  NAND2_X1 U3622 ( .A1(n4207), .A2(n3339), .ZN(n4081) );
  INV_X1 U3624 ( .A(n3340), .ZN(n3324) );
  NOR2_X1 U3625 ( .A1(n4084), .A2(n4207), .ZN(n4097) );
  NOR2_X1 U3626 ( .A1(n6757), .A2(n3601), .ZN(n3633) );
  NAND2_X2 U3627 ( .A1(n3311), .A2(n3310), .ZN(n4084) );
  NOR2_X1 U3628 ( .A1(n3569), .A2(n3571), .ZN(n3595) );
  AND4_X1 U3629 ( .A1(n3199), .A2(n3198), .A3(n3197), .A4(n3196), .ZN(n3207)
         );
  AND4_X1 U3630 ( .A1(n3219), .A2(n3218), .A3(n3217), .A4(n3216), .ZN(n3225)
         );
  AND4_X1 U3631 ( .A1(n3215), .A2(n3214), .A3(n3213), .A4(n3212), .ZN(n3226)
         );
  AND4_X1 U3632 ( .A1(n3262), .A2(n3261), .A3(n3260), .A4(n3259), .ZN(n3263)
         );
  AND4_X1 U3633 ( .A1(n3309), .A2(n3308), .A3(n3307), .A4(n3306), .ZN(n3310)
         );
  AND4_X1 U3634 ( .A1(n3268), .A2(n3267), .A3(n3266), .A4(n3265), .ZN(n3274)
         );
  AND4_X1 U3635 ( .A1(n3272), .A2(n3271), .A3(n3270), .A4(n3269), .ZN(n3273)
         );
  AND4_X1 U3636 ( .A1(n3279), .A2(n3278), .A3(n3277), .A4(n3276), .ZN(n3284)
         );
  AND4_X1 U3637 ( .A1(n3292), .A2(n3291), .A3(n3290), .A4(n3289), .ZN(n3185)
         );
  AND3_X1 U3638 ( .A1(n3287), .A2(n3286), .A3(n3285), .ZN(n3294) );
  AND4_X1 U3639 ( .A1(n3205), .A2(n3204), .A3(n3203), .A4(n3202), .ZN(n3206)
         );
  AND4_X1 U3640 ( .A1(n3231), .A2(n3230), .A3(n3229), .A4(n3228), .ZN(n3237)
         );
  AND4_X1 U3641 ( .A1(n3235), .A2(n3234), .A3(n3233), .A4(n3232), .ZN(n3236)
         );
  AND4_X1 U3642 ( .A1(n3211), .A2(n3210), .A3(n3209), .A4(n3208), .ZN(n3227)
         );
  AOI22_X1 U3643 ( .A1(n3827), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3347), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3198) );
  AND2_X2 U3644 ( .A1(n5176), .A2(n4560), .ZN(n3349) );
  AND2_X2 U3645 ( .A1(n5172), .A2(n4545), .ZN(n3302) );
  AND2_X2 U3646 ( .A1(n5176), .A2(n3200), .ZN(n3367) );
  AND2_X2 U3647 ( .A1(n3200), .A2(n4534), .ZN(n3827) );
  AND2_X2 U3648 ( .A1(n4571), .A2(n3200), .ZN(n3347) );
  AND2_X2 U3649 ( .A1(n5172), .A2(n3200), .ZN(n3360) );
  AND2_X2 U3650 ( .A1(n4545), .A2(n5176), .ZN(n3454) );
  AND2_X2 U3651 ( .A1(n5172), .A2(n4560), .ZN(n3350) );
  AND2_X2 U3652 ( .A1(n3195), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5172)
         );
  AND2_X2 U3653 ( .A1(n5107), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5176)
         );
  AND2_X2 U3654 ( .A1(n3470), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3200)
         );
  AND2_X2 U3655 ( .A1(n4560), .A2(n4534), .ZN(n3305) );
  AND2_X2 U3656 ( .A1(n4571), .A2(n4545), .ZN(n3288) );
  AND2_X2 U3657 ( .A1(n4571), .A2(n4560), .ZN(n3366) );
  AND2_X2 U3658 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4560) );
  CLKBUF_X1 U3659 ( .A(n4855), .Z(n3093) );
  NAND2_X1 U3660 ( .A1(n4857), .A2(n4856), .ZN(n4855) );
  NAND2_X2 U3662 ( .A1(n3317), .A2(n3295), .ZN(n3341) );
  NAND2_X2 U3663 ( .A1(n3237), .A2(n3236), .ZN(n3316) );
  AOI21_X2 U3664 ( .B1(n3482), .B2(n3481), .A(n3419), .ZN(n3479) );
  CLKBUF_X1 U3665 ( .A(n3298), .Z(n3959) );
  AOI21_X2 U3666 ( .B1(n5023), .B2(n5024), .A(n5964), .ZN(n6002) );
  NAND2_X2 U3667 ( .A1(n3698), .A2(n3697), .ZN(n5287) );
  NAND2_X1 U3668 ( .A1(n3093), .A2(n4263), .ZN(n3094) );
  CLKBUF_X1 U3669 ( .A(n6333), .Z(n3101) );
  NAND2_X1 U3670 ( .A1(n4623), .A2(n3099), .ZN(n4184) );
  NAND2_X1 U3671 ( .A1(n5713), .A2(n3149), .ZN(n3148) );
  NOR2_X1 U3672 ( .A1(n3406), .A2(n3104), .ZN(n3096) );
  OR2_X1 U3673 ( .A1(n5499), .A2(n3097), .ZN(n4274) );
  OR2_X1 U3674 ( .A1(n3112), .A2(n5644), .ZN(n3097) );
  OAI22_X2 U3675 ( .A1(n5544), .A2(n3136), .B1(n3138), .B2(n5528), .ZN(n3098)
         );
  NOR2_X2 U3676 ( .A1(n3406), .A2(n3104), .ZN(n4298) );
  OAI22_X1 U3677 ( .A1(n5544), .A2(n3136), .B1(n3138), .B2(n5528), .ZN(n5499)
         );
  NOR2_X1 U3678 ( .A1(n4525), .A2(n3404), .ZN(n4326) );
  NAND2_X1 U3679 ( .A1(n3317), .A2(n3493), .ZN(n3322) );
  XNOR2_X1 U3680 ( .A(n4229), .B(n4205), .ZN(n4843) );
  NAND2_X1 U3681 ( .A1(n3143), .A2(n4204), .ZN(n4229) );
  NAND2_X1 U3682 ( .A1(n4589), .A2(n3469), .ZN(n3144) );
  AND2_X1 U3683 ( .A1(n5172), .A2(n4560), .ZN(n3100) );
  AOI21_X1 U3684 ( .B1(n3406), .B2(n5023), .A(n3342), .ZN(n4089) );
  AOI21_X1 U3685 ( .B1(n3423), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3411), 
        .ZN(n3412) );
  INV_X2 U3686 ( .A(n3341), .ZN(n4307) );
  XNOR2_X1 U3687 ( .A(n4561), .B(n4618), .ZN(n6333) );
  NAND2_X2 U3688 ( .A1(n3326), .A2(n3325), .ZN(n3423) );
  XNOR2_X1 U3689 ( .A(n3402), .B(n3345), .ZN(n3494) );
  AOI211_X1 U3690 ( .C1(n4202), .C2(n6584), .A(n6583), .B(n6582), .ZN(n6587)
         );
  NAND2_X2 U3691 ( .A1(n5492), .A2(n5060), .ZN(n5459) );
  NAND2_X2 U3692 ( .A1(n3414), .A2(n3420), .ZN(n3422) );
  NAND2_X2 U3693 ( .A1(n3413), .A2(n3412), .ZN(n3420) );
  AND2_X1 U3694 ( .A1(n4373), .A2(n4081), .ZN(n4181) );
  NOR2_X2 U3695 ( .A1(n5319), .A2(n5228), .ZN(n5227) );
  NAND2_X2 U3696 ( .A1(n4298), .A2(n3407), .ZN(n4309) );
  NAND2_X2 U3697 ( .A1(n5546), .A2(n5545), .ZN(n5544) );
  NAND2_X1 U3698 ( .A1(n3549), .A2(n3144), .ZN(n4720) );
  AOI21_X4 U3699 ( .B1(n5081), .B2(n5082), .A(n5084), .ZN(n5713) );
  NAND2_X2 U3700 ( .A1(n4968), .A2(n4269), .ZN(n5081) );
  OAI22_X2 U3701 ( .A1(n4235), .A2(n4260), .B1(n4234), .B2(n4258), .ZN(n4236)
         );
  AND2_X2 U3702 ( .A1(n4560), .A2(n4534), .ZN(n3103) );
  INV_X1 U3703 ( .A(n3385), .ZN(n4012) );
  NAND2_X1 U3704 ( .A1(n3578), .A2(n3577), .ZN(n4251) );
  NAND2_X1 U3705 ( .A1(n4491), .A2(n4490), .ZN(n4520) );
  INV_X1 U3706 ( .A(n3146), .ZN(n3145) );
  OAI22_X1 U3707 ( .A1(n5552), .A2(n3147), .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n5716), .ZN(n3146) );
  AND2_X1 U3708 ( .A1(n4306), .A2(n6481), .ZN(n4329) );
  NAND2_X1 U3709 ( .A1(n3565), .A2(n3564), .ZN(n3577) );
  NAND2_X1 U3710 ( .A1(n3377), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3453) );
  INV_X1 U3711 ( .A(n4028), .ZN(n3996) );
  NOR2_X1 U3712 ( .A1(n4299), .A2(n6586), .ZN(n4028) );
  NOR2_X1 U3713 ( .A1(n5361), .A2(n3115), .ZN(n3122) );
  NAND2_X1 U3714 ( .A1(n5699), .A2(n4139), .ZN(n5263) );
  OR2_X1 U3715 ( .A1(n4529), .A2(n4092), .ZN(n4312) );
  INV_X1 U3716 ( .A(n3453), .ZN(n4199) );
  INV_X1 U3717 ( .A(n4026), .ZN(n3952) );
  AND2_X1 U3718 ( .A1(n3178), .A2(n5308), .ZN(n3176) );
  NOR2_X1 U3719 ( .A1(n5128), .A2(n3296), .ZN(n4193) );
  NAND2_X1 U3720 ( .A1(n5716), .A2(n3117), .ZN(n3151) );
  NOR2_X1 U3721 ( .A1(n5716), .A2(n3116), .ZN(n3152) );
  OR2_X1 U3722 ( .A1(n4077), .A2(n4288), .ZN(n4078) );
  NAND2_X1 U3723 ( .A1(n4076), .A2(n4075), .ZN(n4079) );
  OR2_X1 U3724 ( .A1(n5220), .A2(n5947), .ZN(n3127) );
  OAI21_X1 U3725 ( .B1(n4049), .B2(n3541), .A(n3540), .ZN(n3552) );
  OAI21_X1 U3726 ( .B1(n3107), .B2(n3140), .A(n5526), .ZN(n3139) );
  NAND2_X1 U3727 ( .A1(n4373), .A2(n6027), .ZN(n3124) );
  OR2_X1 U3728 ( .A1(n3396), .A2(n3395), .ZN(n4212) );
  NAND2_X1 U3729 ( .A1(n3252), .A2(n3251), .ZN(n4083) );
  INV_X1 U3730 ( .A(n3452), .ZN(n3441) );
  NAND2_X1 U3731 ( .A1(n3324), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3452) );
  AND2_X1 U3732 ( .A1(n3099), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4034) );
  NOR2_X1 U3733 ( .A1(n4344), .A2(n3179), .ZN(n3178) );
  INV_X1 U3734 ( .A(n5120), .ZN(n3179) );
  NOR2_X1 U3735 ( .A1(n3869), .A2(n5339), .ZN(n3164) );
  OR2_X1 U3736 ( .A1(n5328), .A2(n5237), .ZN(n3869) );
  NOR2_X1 U3737 ( .A1(n3174), .A2(n3173), .ZN(n3172) );
  INV_X1 U3738 ( .A(n5360), .ZN(n3173) );
  NAND2_X1 U3739 ( .A1(n3175), .A2(n5261), .ZN(n3174) );
  INV_X1 U3740 ( .A(n5276), .ZN(n3175) );
  NAND2_X1 U3741 ( .A1(n3169), .A2(n5411), .ZN(n3168) );
  INV_X1 U3742 ( .A(n5370), .ZN(n3169) );
  NOR2_X1 U3743 ( .A1(n5454), .A2(n3157), .ZN(n3156) );
  INV_X1 U3744 ( .A(n4279), .ZN(n3157) );
  INV_X1 U3745 ( .A(n4454), .ZN(n3130) );
  OR2_X1 U3746 ( .A1(n3438), .A2(n3437), .ZN(n4206) );
  NAND2_X1 U3747 ( .A1(n3451), .A2(n3450), .ZN(n4618) );
  INV_X1 U3748 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6334) );
  INV_X1 U3749 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6456) );
  AND2_X1 U3750 ( .A1(n4558), .A2(n4557), .ZN(n6462) );
  AND2_X1 U3751 ( .A1(n3950), .A2(n3949), .ZN(n5308) );
  AND2_X1 U3752 ( .A1(n4493), .A2(n4492), .ZN(n5140) );
  NAND2_X1 U3753 ( .A1(n4348), .A2(n4456), .ZN(n4392) );
  INV_X1 U3754 ( .A(n3880), .ZN(n5150) );
  INV_X1 U3755 ( .A(n5317), .ZN(n3907) );
  OR2_X1 U3756 ( .A1(n5854), .A2(n4025), .ZN(n3768) );
  NAND2_X1 U3757 ( .A1(n3736), .A2(n3735), .ZN(n3769) );
  INV_X1 U3758 ( .A(n5285), .ZN(n3697) );
  NAND2_X1 U3759 ( .A1(n4236), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4237)
         );
  XNOR2_X1 U3760 ( .A(n4242), .B(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4850)
         );
  NOR2_X1 U3761 ( .A1(n5188), .A2(n4421), .ZN(n6464) );
  AND2_X1 U3762 ( .A1(n5610), .A2(n4323), .ZN(n5584) );
  NAND2_X1 U3763 ( .A1(n4159), .A2(n3122), .ZN(n3121) );
  INV_X1 U3764 ( .A(n3122), .ZN(n3119) );
  AND2_X1 U3765 ( .A1(n6134), .A2(n4316), .ZN(n5703) );
  AND3_X1 U3766 ( .A1(n4199), .A2(n4250), .A3(n4264), .ZN(n4200) );
  NAND2_X1 U3767 ( .A1(n4329), .A2(n5183), .ZN(n5641) );
  NAND2_X1 U3768 ( .A1(n4329), .A2(n6452), .ZN(n5690) );
  INV_X1 U3769 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6451) );
  INV_X1 U3770 ( .A(n4697), .ZN(n4757) );
  AND2_X1 U3771 ( .A1(n4523), .A2(n4580), .ZN(n6264) );
  AND2_X1 U3772 ( .A1(n4576), .A2(n5728), .ZN(n5731) );
  INV_X1 U3773 ( .A(n4713), .ZN(n4770) );
  INV_X2 U3774 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6583) );
  AND2_X1 U3775 ( .A1(n6006), .A2(n5222), .ZN(n3128) );
  INV_X1 U3776 ( .A(n5980), .ZN(n5947) );
  XNOR2_X1 U3777 ( .A(n4195), .B(n5201), .ZN(n5220) );
  NOR2_X1 U3778 ( .A1(n4193), .A2(n4192), .ZN(n4195) );
  NAND2_X2 U3779 ( .A1(n4099), .A2(n4098), .ZN(n6026) );
  OR2_X1 U3780 ( .A1(n4494), .A2(n5203), .ZN(n4098) );
  INV_X1 U3781 ( .A(n5148), .ZN(n4032) );
  NAND2_X1 U3782 ( .A1(n4329), .A2(n4311), .ZN(n6184) );
  CLKBUF_X1 U3783 ( .A(n4522), .Z(n4523) );
  INV_X1 U3784 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6460) );
  NAND2_X1 U3785 ( .A1(n3488), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3134) );
  NAND2_X1 U3786 ( .A1(n3552), .A2(n3551), .ZN(n3553) );
  OR2_X1 U3787 ( .A1(n3563), .A2(n3562), .ZN(n4256) );
  OR2_X1 U3788 ( .A1(n3515), .A2(n3514), .ZN(n4246) );
  AND3_X1 U3789 ( .A1(n3400), .A2(n3399), .A3(n3398), .ZN(n3416) );
  AOI21_X1 U3790 ( .B1(n4580), .B2(n6586), .A(n3415), .ZN(n3481) );
  AND2_X1 U3791 ( .A1(n4199), .A2(n4212), .ZN(n3415) );
  AND3_X1 U3792 ( .A1(n4301), .A2(n3095), .A3(n4300), .ZN(n4308) );
  NOR2_X1 U3793 ( .A1(n3258), .A2(n3257), .ZN(n3264) );
  AOI21_X1 U3794 ( .B1(n3302), .B2(INSTQUEUE_REG_1__2__SCAN_IN), .A(n3161), 
        .ZN(n3303) );
  AOI21_X1 U3795 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6460), .A(n4066), 
        .ZN(n4072) );
  INV_X1 U3796 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6834) );
  AOI22_X1 U3797 ( .A1(n3367), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3278) );
  NAND2_X1 U3798 ( .A1(n3692), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3699)
         );
  NOR2_X1 U3799 ( .A1(n3497), .A2(n6834), .ZN(n3519) );
  NAND2_X1 U3800 ( .A1(n5716), .A2(n3184), .ZN(n4279) );
  NAND2_X1 U3801 ( .A1(n3141), .A2(n3142), .ZN(n3136) );
  INV_X1 U3802 ( .A(n3139), .ZN(n3138) );
  NAND2_X1 U3803 ( .A1(n3152), .A2(n3151), .ZN(n3147) );
  NOR2_X1 U3804 ( .A1(n5552), .A2(n3150), .ZN(n3149) );
  INV_X1 U3805 ( .A(n3151), .ZN(n3150) );
  NOR2_X1 U3806 ( .A1(n4453), .A2(n4113), .ZN(n3129) );
  NAND2_X1 U3807 ( .A1(n4101), .A2(n3123), .ZN(n4103) );
  INV_X1 U3808 ( .A(n4083), .ZN(n4291) );
  NAND2_X1 U3809 ( .A1(n3406), .A2(n3441), .ZN(n3325) );
  INV_X1 U3810 ( .A(n4068), .ZN(n4049) );
  XNOR2_X1 U3811 ( .A(n3443), .B(n3442), .ZN(n3477) );
  NAND2_X1 U3812 ( .A1(n3440), .A2(n3439), .ZN(n3443) );
  OR2_X1 U3813 ( .A1(n3322), .A2(n3718), .ZN(n4299) );
  AND4_X1 U3814 ( .A1(n4087), .A2(n4302), .A3(n4086), .A4(n4085), .ZN(n4088)
         );
  AND2_X1 U3815 ( .A1(n3447), .A2(n4768), .ZN(n4690) );
  OAI21_X1 U3816 ( .B1(n6495), .B2(n5725), .A(n6564), .ZN(n4622) );
  NAND2_X1 U3817 ( .A1(n6586), .A2(n4622), .ZN(n4697) );
  NAND2_X1 U3818 ( .A1(n4068), .A2(n4250), .ZN(n4075) );
  AND2_X1 U3819 ( .A1(n4360), .A2(n5921), .ZN(n5838) );
  NAND2_X1 U3820 ( .A1(n3324), .A2(n3339), .ZN(n5026) );
  AND2_X1 U3821 ( .A1(n4371), .A2(n5024), .ZN(n4353) );
  AND2_X1 U3822 ( .A1(n4130), .A2(n4129), .ZN(n5373) );
  XNOR2_X1 U3823 ( .A(n4103), .B(n4395), .ZN(n4436) );
  AND2_X1 U3824 ( .A1(n3178), .A2(n3114), .ZN(n3177) );
  AND2_X1 U3825 ( .A1(n3971), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3972)
         );
  NAND2_X1 U3826 ( .A1(n5310), .A2(n5120), .ZN(n5122) );
  AND2_X1 U3827 ( .A1(n3927), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3928)
         );
  AND2_X1 U3828 ( .A1(n3164), .A2(n5077), .ZN(n3163) );
  NAND2_X1 U3829 ( .A1(n3853), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3886)
         );
  NAND2_X1 U3830 ( .A1(n3820), .A2(n3819), .ZN(n5337) );
  OR2_X1 U3831 ( .A1(n3786), .A2(n6702), .ZN(n3803) );
  NAND2_X1 U3832 ( .A1(n3113), .A2(n3172), .ZN(n3171) );
  NOR2_X1 U3833 ( .A1(n3769), .A2(n6615), .ZN(n3770) );
  NOR2_X1 U3834 ( .A1(n3717), .A2(n3716), .ZN(n3736) );
  AND2_X1 U3835 ( .A1(n3752), .A2(n3751), .ZN(n5360) );
  NAND2_X1 U3836 ( .A1(n3170), .A2(n3172), .ZN(n5359) );
  INV_X1 U3837 ( .A(n5287), .ZN(n3170) );
  OR2_X1 U3838 ( .A1(n3699), .A2(n5538), .ZN(n3717) );
  AND3_X1 U3839 ( .A1(n3696), .A2(n3695), .A3(n3694), .ZN(n5285) );
  NOR2_X1 U3840 ( .A1(n3168), .A2(n3167), .ZN(n3166) );
  INV_X1 U3841 ( .A(n5053), .ZN(n3167) );
  OR2_X1 U3842 ( .A1(n3649), .A2(n5938), .ZN(n3650) );
  NOR2_X1 U3843 ( .A1(n6870), .A2(n3650), .ZN(n3692) );
  NAND2_X1 U3844 ( .A1(n3633), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3649)
         );
  INV_X1 U3845 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5938) );
  NOR2_X1 U3846 ( .A1(n5371), .A2(n5370), .ZN(n5412) );
  NAND2_X1 U3847 ( .A1(n3600), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3601)
         );
  INV_X1 U3848 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6757) );
  AND2_X1 U3849 ( .A1(n3595), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3600)
         );
  AOI21_X1 U3850 ( .B1(n3584), .B2(n3708), .A(n3583), .ZN(n4614) );
  NAND2_X1 U3851 ( .A1(n3568), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3569)
         );
  NAND2_X1 U3852 ( .A1(n3091), .A2(n3162), .ZN(n4610) );
  AND2_X1 U3853 ( .A1(n3548), .A2(n4507), .ZN(n3162) );
  AOI21_X1 U3854 ( .B1(n4249), .B2(n3708), .A(n3575), .ZN(n4609) );
  AND2_X1 U3855 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3519), .ZN(n3568)
         );
  INV_X1 U3856 ( .A(n3155), .ZN(n3154) );
  OAI21_X1 U3857 ( .B1(n3156), .B2(n3188), .A(n3158), .ZN(n3155) );
  INV_X1 U3858 ( .A(n5145), .ZN(n3158) );
  NOR2_X1 U3859 ( .A1(n5422), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5426)
         );
  OR2_X1 U3860 ( .A1(n5323), .A2(n5229), .ZN(n5313) );
  INV_X1 U3861 ( .A(n3160), .ZN(n5453) );
  NOR2_X1 U3862 ( .A1(n5342), .A2(n4165), .ZN(n5332) );
  AND2_X1 U3863 ( .A1(n4149), .A2(n4148), .ZN(n5361) );
  NOR2_X1 U3864 ( .A1(n5362), .A2(n5361), .ZN(n5364) );
  NAND2_X1 U3865 ( .A1(n5544), .A2(n3107), .ZN(n3137) );
  NAND2_X1 U3866 ( .A1(n3126), .A2(n3125), .ZN(n5700) );
  INV_X1 U3867 ( .A(n5373), .ZN(n3125) );
  OR2_X1 U3868 ( .A1(n6179), .A2(n4332), .ZN(n5642) );
  OR2_X1 U3869 ( .A1(n5641), .A2(n4333), .ZN(n5871) );
  AND2_X1 U3870 ( .A1(n4735), .A2(n4734), .ZN(n5035) );
  AND2_X1 U3871 ( .A1(n4120), .A2(n4119), .ZN(n4633) );
  NOR2_X1 U3872 ( .A1(n5958), .A2(n4633), .ZN(n4735) );
  OR2_X1 U3873 ( .A1(n5956), .A2(n5955), .ZN(n5958) );
  NAND2_X1 U3874 ( .A1(n4243), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4244)
         );
  NAND2_X1 U3875 ( .A1(n3130), .A2(n3131), .ZN(n4452) );
  NAND2_X1 U3876 ( .A1(n4222), .A2(n4221), .ZN(n4399) );
  NOR2_X1 U3877 ( .A1(n3338), .A2(n3337), .ZN(n3343) );
  NAND2_X1 U3878 ( .A1(n3494), .A2(n6586), .ZN(n3132) );
  INV_X1 U3879 ( .A(n4299), .ZN(n5167) );
  NOR2_X1 U3880 ( .A1(n4521), .A2(n4520), .ZN(n6449) );
  NAND2_X1 U3881 ( .A1(n5102), .A2(n4622), .ZN(n4758) );
  AND2_X1 U3882 ( .A1(n6858), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4095) );
  INV_X1 U3883 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5829) );
  INV_X1 U3884 ( .A(n5995), .ZN(n5969) );
  AND2_X1 U3885 ( .A1(n5966), .A2(REIP_REG_5__SCAN_IN), .ZN(n5960) );
  AND2_X1 U3886 ( .A1(n4373), .A2(n4372), .ZN(n5980) );
  AND2_X1 U3887 ( .A1(n5044), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5990) );
  AND2_X1 U3888 ( .A1(n5155), .A2(n4379), .ZN(n6006) );
  AND2_X1 U3889 ( .A1(n5419), .A2(n4500), .ZN(n6832) );
  INV_X2 U3890 ( .A(n5419), .ZN(n6830) );
  AND2_X1 U3891 ( .A1(n5419), .A2(n4501), .ZN(n6831) );
  INV_X2 U3892 ( .A(n6832), .ZN(n5418) );
  INV_X1 U3893 ( .A(n6831), .ZN(n5421) );
  AND2_X1 U3894 ( .A1(n4459), .A2(n4509), .ZN(n6055) );
  INV_X1 U3895 ( .A(n6055), .ZN(n6060) );
  INV_X1 U3896 ( .A(n4458), .ZN(n6069) );
  OR3_X1 U3897 ( .A1(n4392), .A2(n3407), .A3(READY_N), .ZN(n4493) );
  INV_X1 U3898 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6772) );
  INV_X1 U3899 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6702) );
  NAND2_X1 U3900 ( .A1(n5544), .A2(n3182), .ZN(n5536) );
  INV_X1 U3901 ( .A(n6097), .ZN(n5548) );
  INV_X1 U3902 ( .A(n6108), .ZN(n6074) );
  INV_X1 U3903 ( .A(n4193), .ZN(n5199) );
  AND2_X1 U3904 ( .A1(n5621), .A2(n4322), .ZN(n5610) );
  XNOR2_X1 U3905 ( .A(n5066), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5080)
         );
  NAND2_X1 U3906 ( .A1(n5065), .A2(n5064), .ZN(n5066) );
  AND2_X1 U3907 ( .A1(n5637), .A2(n5461), .ZN(n5623) );
  NOR2_X1 U3908 ( .A1(n5674), .A2(n4336), .ZN(n5637) );
  OR2_X1 U3909 ( .A1(n5670), .A2(n4320), .ZN(n5636) );
  NOR2_X1 U3910 ( .A1(n5362), .A2(n3119), .ZN(n5347) );
  INV_X1 U3911 ( .A(n5493), .ZN(n5060) );
  OAI21_X1 U3912 ( .B1(n5713), .B2(n3152), .A(n3151), .ZN(n5553) );
  INV_X1 U3913 ( .A(n6190), .ZN(n6156) );
  INV_X1 U3914 ( .A(n6184), .ZN(n6167) );
  INV_X1 U3915 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6858) );
  AND2_X1 U3916 ( .A1(n3096), .A2(n4510), .ZN(n6452) );
  NOR2_X1 U3917 ( .A1(n5102), .A2(n5883), .ZN(n5164) );
  INV_X1 U3918 ( .A(n6477), .ZN(n6564) );
  NOR2_X1 U3919 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n5881) );
  INV_X1 U3920 ( .A(n4979), .ZN(n5014) );
  OAI21_X1 U3921 ( .B1(n6200), .B2(n6215), .A(n6336), .ZN(n6218) );
  INV_X1 U3922 ( .A(n6221), .ZN(n6197) );
  OAI21_X1 U3923 ( .B1(n6230), .B2(n4620), .A(n4619), .ZN(n4919) );
  INV_X1 U3924 ( .A(n6231), .ZN(n6250) );
  OR4_X1 U3925 ( .A1(n6269), .A2(n6268), .A3(n6340), .A4(n6267), .ZN(n6294) );
  INV_X1 U3926 ( .A(n6262), .ZN(n6293) );
  INV_X1 U3927 ( .A(n6302), .ZN(n6324) );
  OR3_X1 U3928 ( .A1(n4645), .A2(n6269), .A3(n4644), .ZN(n4964) );
  INV_X1 U3929 ( .A(n6400), .ZN(n6344) );
  AND2_X1 U3930 ( .A1(n6101), .A2(DATAI_24_), .ZN(n6397) );
  INV_X1 U3931 ( .A(n6406), .ZN(n6347) );
  NOR2_X1 U3932 ( .A1(n4758), .A2(n3407), .ZN(n6401) );
  INV_X1 U3933 ( .A(n6412), .ZN(n6351) );
  AND2_X1 U3934 ( .A1(n6101), .A2(DATAI_26_), .ZN(n6409) );
  INV_X1 U3935 ( .A(n6418), .ZN(n6355) );
  NOR2_X1 U3936 ( .A1(n4758), .A2(n4623), .ZN(n6413) );
  INV_X1 U3937 ( .A(n6424), .ZN(n6359) );
  AND2_X1 U3938 ( .A1(n6101), .A2(DATAI_28_), .ZN(n6420) );
  INV_X1 U3939 ( .A(n6430), .ZN(n6363) );
  AND2_X1 U3940 ( .A1(n6101), .A2(DATAI_29_), .ZN(n6426) );
  INV_X1 U3941 ( .A(n6436), .ZN(n6367) );
  AND2_X1 U3942 ( .A1(n6101), .A2(DATAI_30_), .ZN(n6432) );
  NOR2_X1 U3943 ( .A1(n4758), .A2(n3250), .ZN(n6438) );
  AND2_X1 U3944 ( .A1(n4713), .A2(n4637), .ZN(n4963) );
  AND2_X1 U3945 ( .A1(n4713), .A2(n4657), .ZN(n4942) );
  AND2_X1 U3946 ( .A1(n6101), .A2(DATAI_31_), .ZN(n6442) );
  AND2_X1 U3947 ( .A1(n4095), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6481) );
  AND2_X1 U3948 ( .A1(n6476), .A2(n6475), .ZN(n6484) );
  NOR2_X1 U3949 ( .A1(n6688), .A2(n5188), .ZN(n6477) );
  INV_X1 U3950 ( .A(n6481), .ZN(n6485) );
  INV_X1 U3951 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6504) );
  INV_X1 U3952 ( .A(n6547), .ZN(n6593) );
  OAI211_X1 U3953 ( .C1(n5223), .C2(REIP_REG_30__SCAN_IN), .A(n3110), .B(n3127), .ZN(n5224) );
  OAI22_X1 U3954 ( .A1(n5220), .A2(n5376), .B1(n5219), .B2(n6026), .ZN(n4196)
         );
  AND2_X1 U3955 ( .A1(n4342), .A2(n4341), .ZN(n4343) );
  OR2_X1 U3956 ( .A1(n3341), .A2(n3099), .ZN(n3104) );
  AND2_X1 U3957 ( .A1(n3402), .A2(n3401), .ZN(n3421) );
  NAND2_X1 U3958 ( .A1(n5557), .A2(n6624), .ZN(n3105) );
  INV_X1 U3959 ( .A(n4025), .ZN(n3969) );
  INV_X1 U3960 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5107) );
  AND2_X1 U3961 ( .A1(n3820), .A2(n3164), .ZN(n5075) );
  AND4_X1 U3962 ( .A1(n3283), .A2(n3282), .A3(n3281), .A4(n3280), .ZN(n3106)
         );
  AND2_X1 U3963 ( .A1(n3105), .A2(n3182), .ZN(n3107) );
  OR2_X1 U3964 ( .A1(n5163), .A2(n5842), .ZN(n3108) );
  INV_X1 U3965 ( .A(n3488), .ZN(n3135) );
  AND2_X1 U3966 ( .A1(n5716), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3109)
         );
  INV_X1 U3967 ( .A(n5528), .ZN(n3142) );
  INV_X1 U3968 ( .A(n4453), .ZN(n3131) );
  NOR2_X1 U3969 ( .A1(n5221), .A2(n3128), .ZN(n3110) );
  INV_X1 U3970 ( .A(n3141), .ZN(n3140) );
  NAND2_X1 U3971 ( .A1(n3105), .A2(n3109), .ZN(n3141) );
  NAND2_X1 U3972 ( .A1(n3091), .A2(n4507), .ZN(n4506) );
  NOR2_X1 U3973 ( .A1(n5287), .A2(n5276), .ZN(n5258) );
  NOR2_X1 U3974 ( .A1(n5371), .A2(n3168), .ZN(n5051) );
  NAND2_X1 U3975 ( .A1(n3165), .A2(n3166), .ZN(n5052) );
  NAND2_X1 U3976 ( .A1(n3137), .A2(n3141), .ZN(n5525) );
  INV_X1 U3977 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6586) );
  INV_X1 U3978 ( .A(n5339), .ZN(n3819) );
  INV_X1 U3979 ( .A(n3120), .ZN(n5342) );
  NOR2_X1 U3980 ( .A1(n5362), .A2(n3121), .ZN(n3120) );
  AND2_X1 U3981 ( .A1(n5557), .A2(n5500), .ZN(n3112) );
  NOR2_X1 U3982 ( .A1(n5334), .A2(n5068), .ZN(n5067) );
  NOR2_X1 U3983 ( .A1(n5351), .A2(n5246), .ZN(n3113) );
  AND2_X1 U3984 ( .A1(n5148), .A2(n5308), .ZN(n3114) );
  INV_X1 U3985 ( .A(n4250), .ZN(n4260) );
  AND2_X1 U3986 ( .A1(n5139), .A2(n4510), .ZN(n4250) );
  NOR2_X1 U3987 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4031) );
  INV_X1 U3988 ( .A(n4031), .ZN(n4025) );
  INV_X1 U3989 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3470) );
  INV_X1 U3990 ( .A(n3126), .ZN(n5374) );
  NOR2_X1 U3991 ( .A1(n5037), .A2(n4866), .ZN(n3126) );
  NAND2_X1 U3992 ( .A1(n3466), .A2(n3465), .ZN(n3468) );
  NAND2_X1 U3993 ( .A1(n4420), .A2(n6380), .ZN(n5564) );
  NAND2_X1 U3994 ( .A1(n4560), .A2(n4534), .ZN(n3385) );
  NAND2_X1 U3995 ( .A1(n4153), .A2(n4152), .ZN(n3115) );
  AND2_X1 U3996 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3116) );
  NAND2_X1 U3997 ( .A1(n4270), .A2(n3153), .ZN(n3117) );
  AND2_X1 U3998 ( .A1(n3130), .A2(n3129), .ZN(n3118) );
  INV_X2 U3999 ( .A(n4373), .ZN(n5203) );
  NAND3_X1 U4000 ( .A1(n3124), .A2(n4184), .A3(n4100), .ZN(n3123) );
  NAND3_X1 U4001 ( .A1(n3130), .A2(n3129), .A3(n4654), .ZN(n5956) );
  NAND2_X1 U4002 ( .A1(n6010), .A2(n4104), .ZN(n4454) );
  NOR2_X2 U4003 ( .A1(n5313), .A2(n4188), .ZN(n5128) );
  NOR2_X2 U4004 ( .A1(n3098), .A2(n3112), .ZN(n5501) );
  NAND3_X1 U4005 ( .A1(n3549), .A2(n3144), .A3(n4250), .ZN(n3143) );
  NAND2_X1 U4006 ( .A1(n5713), .A2(n4270), .ZN(n5715) );
  INV_X1 U4007 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3153) );
  NAND2_X1 U4008 ( .A1(n4280), .A2(n3156), .ZN(n3160) );
  NAND2_X1 U4009 ( .A1(n4280), .A2(n4279), .ZN(n5116) );
  INV_X1 U4010 ( .A(n3188), .ZN(n3159) );
  NAND3_X1 U4011 ( .A1(n4097), .A2(n5023), .A3(n3403), .ZN(n4525) );
  INV_X1 U4012 ( .A(n3366), .ZN(n3979) );
  AND2_X1 U4013 ( .A1(n3366), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3161) );
  INV_X1 U4014 ( .A(n4720), .ZN(n3476) );
  INV_X1 U4015 ( .A(n5076), .ZN(n3908) );
  NAND2_X1 U4016 ( .A1(n3820), .A2(n3163), .ZN(n5076) );
  INV_X1 U4017 ( .A(n5371), .ZN(n3165) );
  INV_X1 U4018 ( .A(n5052), .ZN(n3698) );
  NOR2_X2 U4019 ( .A1(n5287), .A2(n3171), .ZN(n5353) );
  NOR2_X1 U4020 ( .A1(n5287), .A2(n3174), .ZN(n5259) );
  AND2_X1 U4021 ( .A1(n5227), .A2(n3176), .ZN(n5149) );
  AND2_X2 U4022 ( .A1(n5227), .A2(n5308), .ZN(n5310) );
  NAND2_X1 U4023 ( .A1(n5227), .A2(n3177), .ZN(n5153) );
  XNOR2_X1 U4024 ( .A(n4236), .B(n6163), .ZN(n6089) );
  OAI21_X1 U4025 ( .B1(n5425), .B2(n5424), .A(n5423), .ZN(n5427) );
  NAND2_X1 U4026 ( .A1(n5217), .A2(n6023), .ZN(n4198) );
  AOI211_X2 U4027 ( .C1(n6074), .C2(n5132), .A(n5124), .B(n5123), .ZN(n5125)
         );
  NOR2_X2 U4028 ( .A1(n5478), .A2(n5479), .ZN(n5477) );
  NAND2_X1 U4029 ( .A1(n4275), .A2(n4274), .ZN(n5492) );
  NAND2_X1 U4030 ( .A1(n5444), .A2(n5442), .ZN(n5435) );
  CLKBUF_X1 U4031 ( .A(n3098), .Z(n5517) );
  INV_X1 U4032 ( .A(n5432), .ZN(n5163) );
  NOR2_X1 U4033 ( .A1(n4720), .A2(n4713), .ZN(n6379) );
  CLKBUF_X1 U4034 ( .A(n4575), .Z(n4713) );
  AND2_X1 U4035 ( .A1(n3186), .A2(n3303), .ZN(n3311) );
  INV_X1 U4036 ( .A(n4084), .ZN(n4746) );
  NOR2_X4 U4037 ( .A1(n3099), .A2(n3339), .ZN(n5023) );
  AND2_X1 U4038 ( .A1(n5319), .A2(n5318), .ZN(n5804) );
  XNOR2_X1 U4039 ( .A(n5149), .B(n4032), .ZN(n5217) );
  AND3_X1 U4040 ( .A1(n4292), .A2(n4291), .A3(n3099), .ZN(n4348) );
  OR2_X1 U4041 ( .A1(n3411), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3180)
         );
  OR2_X1 U4042 ( .A1(n5716), .A2(n4276), .ZN(n3181) );
  OR2_X1 U4043 ( .A1(n5716), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3182)
         );
  OR2_X1 U4044 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3183)
         );
  NOR2_X1 U4045 ( .A1(n3472), .A2(n6583), .ZN(n3543) );
  INV_X1 U4046 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4271) );
  OR4_X1 U4047 ( .A1(n5645), .A2(n5629), .A3(INSTADDRPOINTER_REG_24__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3184) );
  AND3_X1 U4048 ( .A1(n3301), .A2(n3300), .A3(n3299), .ZN(n3186) );
  AND4_X1 U4049 ( .A1(n3358), .A2(n3357), .A3(n3356), .A4(n3355), .ZN(n3187)
         );
  AND2_X1 U4050 ( .A1(n5557), .A2(n6731), .ZN(n3188) );
  AND2_X1 U4051 ( .A1(n5557), .A2(n3192), .ZN(n3189) );
  AND2_X1 U4052 ( .A1(n5557), .A2(n6760), .ZN(n3190) );
  INV_X1 U4053 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3716) );
  INV_X1 U4054 ( .A(n6590), .ZN(n6051) );
  OR2_X1 U4055 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3191)
         );
  INV_X1 U4056 ( .A(n6061), .ZN(n4464) );
  INV_X1 U4057 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3571) );
  AND2_X1 U4058 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3192) );
  AND3_X1 U4059 ( .A1(n3353), .A2(n3352), .A3(n3351), .ZN(n3193) );
  OR2_X1 U4060 ( .A1(n5197), .A2(n5428), .ZN(n3194) );
  INV_X1 U4061 ( .A(n5376), .ZN(n6022) );
  NAND2_X1 U4062 ( .A1(n6026), .A2(n3250), .ZN(n5376) );
  AND2_X1 U4063 ( .A1(n6026), .A2(n3472), .ZN(n6023) );
  INV_X1 U4064 ( .A(n3404), .ZN(n3319) );
  NOR2_X1 U4065 ( .A1(n5023), .A2(n4036), .ZN(n4060) );
  AND2_X1 U4066 ( .A1(n3251), .A2(n3472), .ZN(n3248) );
  INV_X1 U4067 ( .A(n3472), .ZN(n3250) );
  INV_X1 U4068 ( .A(n3376), .ZN(n3295) );
  INV_X1 U4069 ( .A(n3550), .ZN(n3551) );
  NOR2_X1 U4070 ( .A1(n3250), .A2(n3376), .ZN(n3252) );
  OR2_X1 U4071 ( .A1(n3464), .A2(n3463), .ZN(n4232) );
  AND2_X1 U4072 ( .A1(n3517), .A2(n3516), .ZN(n3550) );
  OR2_X1 U4073 ( .A1(n3539), .A2(n3538), .ZN(n4245) );
  AND2_X1 U4074 ( .A1(n4056), .A2(n4055), .ZN(n4066) );
  NAND2_X1 U4075 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6451), .ZN(n4043) );
  INV_X1 U4076 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6615) );
  INV_X1 U4077 ( .A(n3543), .ZN(n4026) );
  INV_X1 U4078 ( .A(n4080), .ZN(n4301) );
  INV_X1 U4079 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4205) );
  AND2_X1 U4080 ( .A1(n5885), .A2(n4072), .ZN(n4067) );
  NOR2_X1 U4081 ( .A1(n5848), .A2(n5850), .ZN(n5839) );
  AND2_X1 U4082 ( .A1(n3099), .A2(n4353), .ZN(n4354) );
  OR2_X1 U4083 ( .A1(n5790), .A2(n4025), .ZN(n3950) );
  NAND2_X1 U4084 ( .A1(n3972), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4345)
         );
  NAND2_X1 U4085 ( .A1(n3770), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3786)
         );
  INV_X1 U4086 ( .A(n4946), .ZN(n3617) );
  INV_X1 U4087 ( .A(n4181), .ZN(n4180) );
  OR2_X1 U4088 ( .A1(n4268), .A2(n6739), .ZN(n4269) );
  XNOR2_X1 U4089 ( .A(n3482), .B(n3481), .ZN(n4210) );
  NOR2_X1 U4090 ( .A1(n4312), .A2(n4093), .ZN(n5183) );
  OR2_X1 U4091 ( .A1(n4523), .A2(n4580), .ZN(n4696) );
  INV_X1 U4092 ( .A(n3489), .ZN(n3490) );
  NAND2_X1 U4093 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4067), .ZN(n4287) );
  NOR2_X1 U4094 ( .A1(n3887), .A2(n3902), .ZN(n3927) );
  INV_X1 U4095 ( .A(n5067), .ZN(n5321) );
  AND2_X1 U4096 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3735) );
  INV_X1 U4097 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6870) );
  OR2_X1 U4098 ( .A1(n4345), .A2(n6869), .ZN(n4347) );
  INV_X1 U4099 ( .A(n5990), .ZN(n6000) );
  NAND2_X1 U4100 ( .A1(n4355), .A2(n4354), .ZN(n5983) );
  OR2_X1 U4101 ( .A1(n5810), .A2(n4025), .ZN(n3885) );
  NOR2_X1 U4102 ( .A1(n5188), .A2(n6485), .ZN(n4456) );
  NAND2_X1 U4103 ( .A1(n3928), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3970)
         );
  OR2_X1 U4104 ( .A1(n5916), .A2(n4025), .ZN(n3752) );
  INV_X1 U4105 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5538) );
  AND2_X1 U4106 ( .A1(n3616), .A2(n3615), .ZN(n4946) );
  NAND2_X1 U4107 ( .A1(n4254), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4255)
         );
  OR2_X1 U4108 ( .A1(n4449), .A2(n4496), .ZN(n4443) );
  NOR2_X2 U4109 ( .A1(n5435), .A2(n4339), .ZN(n5425) );
  NAND2_X1 U4110 ( .A1(n5716), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5061) );
  NAND2_X1 U4111 ( .A1(n5875), .A2(n4335), .ZN(n5674) );
  NOR2_X1 U4112 ( .A1(n5557), .A2(n4318), .ZN(n5528) );
  INV_X1 U4113 ( .A(n6174), .ZN(n6127) );
  NAND2_X1 U4114 ( .A1(n4079), .A2(n4078), .ZN(n5188) );
  OR2_X1 U4115 ( .A1(n4981), .A2(n6226), .ZN(n6196) );
  INV_X1 U4116 ( .A(n4576), .ZN(n4769) );
  INV_X1 U4117 ( .A(n6379), .ZN(n6330) );
  NAND2_X1 U4118 ( .A1(n3135), .A2(n3490), .ZN(n3491) );
  AOI21_X1 U4119 ( .B1(n6451), .B2(STATE2_REG_3__SCAN_IN), .A(n4697), .ZN(
        n6306) );
  NAND2_X1 U4120 ( .A1(n5067), .A2(n4177), .ZN(n5323) );
  NOR2_X1 U4121 ( .A1(n6541), .A2(n5825), .ZN(n5805) );
  XNOR2_X1 U4122 ( .A(n4347), .B(n4346), .ZN(n5155) );
  INV_X1 U4123 ( .A(n5944), .ZN(n5984) );
  AND2_X1 U4124 ( .A1(n4377), .A2(n5024), .ZN(n5995) );
  INV_X1 U4125 ( .A(n6059), .ZN(n6054) );
  INV_X1 U4126 ( .A(n4464), .ZN(n6070) );
  INV_X1 U4127 ( .A(n4493), .ZN(n6063) );
  NAND2_X1 U4128 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3497) );
  INV_X1 U4129 ( .A(n6078), .ZN(n6104) );
  NOR2_X1 U4130 ( .A1(n5477), .A2(n3190), .ZN(n5470) );
  NAND2_X1 U4131 ( .A1(n5642), .A2(n5871), .ZN(n5875) );
  NAND2_X1 U4132 ( .A1(n4313), .A2(n5690), .ZN(n6137) );
  INV_X1 U4133 ( .A(n5641), .ZN(n6178) );
  AND2_X1 U4134 ( .A1(n4329), .A2(n4328), .ZN(n6174) );
  INV_X1 U4135 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4048) );
  OAI21_X1 U4136 ( .B1(n4978), .B2(n4661), .A(n4660), .ZN(n4938) );
  INV_X1 U4137 ( .A(n4980), .ZN(n5012) );
  INV_X1 U4138 ( .A(n6196), .ZN(n6217) );
  OAI21_X1 U4139 ( .B1(n4725), .B2(n4724), .A(n4723), .ZN(n4884) );
  INV_X1 U4140 ( .A(n4881), .ZN(n4923) );
  INV_X1 U4141 ( .A(n6380), .ZN(n6393) );
  AND2_X1 U4142 ( .A1(n4713), .A2(n4589), .ZN(n6257) );
  AND2_X1 U4143 ( .A1(n6257), .A2(n5731), .ZN(n6322) );
  NOR2_X1 U4144 ( .A1(n6330), .A2(n5732), .ZN(n6440) );
  NOR2_X1 U4145 ( .A1(n4758), .A2(n4746), .ZN(n6407) );
  NOR2_X1 U4146 ( .A1(n4758), .A2(n3403), .ZN(n6425) );
  INV_X1 U4147 ( .A(n6446), .ZN(n6373) );
  NOR2_X1 U4148 ( .A1(n6583), .A2(n6858), .ZN(n5725) );
  INV_X1 U4149 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6507) );
  NAND2_X1 U4150 ( .A1(n6507), .A2(STATE_REG_1__SCAN_IN), .ZN(n6580) );
  NOR2_X1 U4151 ( .A1(n5838), .A2(n4362), .ZN(n5826) );
  OR2_X1 U4152 ( .A1(n5155), .A2(n4378), .ZN(n5842) );
  INV_X1 U4153 ( .A(n4196), .ZN(n4197) );
  INV_X1 U4154 ( .A(n5217), .ZN(n5380) );
  INV_X1 U4155 ( .A(n5804), .ZN(n5388) );
  NAND2_X1 U4156 ( .A1(n5140), .A2(n4495), .ZN(n5419) );
  OR2_X1 U4157 ( .A1(n6055), .A2(n6051), .ZN(n6059) );
  OR2_X1 U4158 ( .A1(n4392), .A2(n4510), .ZN(n4458) );
  OR2_X1 U4159 ( .A1(n6097), .A2(n4825), .ZN(n6108) );
  NAND2_X1 U4160 ( .A1(n6464), .A2(n6481), .ZN(n6078) );
  OR2_X1 U4161 ( .A1(n5612), .A2(n5603), .ZN(n5598) );
  OR2_X1 U4162 ( .A1(n4422), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6190) );
  NOR2_X1 U4163 ( .A1(n4574), .A2(n4757), .ZN(n6191) );
  INV_X1 U4164 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5885) );
  OR2_X1 U4165 ( .A1(n4981), .A2(n5728), .ZN(n4980) );
  AOI21_X1 U4166 ( .B1(n6393), .B2(n6228), .A(n6225), .ZN(n6255) );
  NAND2_X1 U4167 ( .A1(n6257), .A2(n6256), .ZN(n6302) );
  NAND2_X1 U4168 ( .A1(n4676), .A2(n6226), .ZN(n4906) );
  AOI21_X1 U4169 ( .B1(n6338), .B2(n6342), .A(n6337), .ZN(n6377) );
  AND2_X1 U4170 ( .A1(n6387), .A2(n6386), .ZN(n6447) );
  INV_X1 U4171 ( .A(n6440), .ZN(n5788) );
  NAND2_X1 U4172 ( .A1(n4636), .A2(n5728), .ZN(n4967) );
  AOI21_X1 U4173 ( .B1(n4776), .B2(n4774), .A(n4773), .ZN(n4802) );
  INV_X1 U4174 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6688) );
  INV_X1 U4175 ( .A(n6560), .ZN(n6496) );
  INV_X1 U4176 ( .A(n6580), .ZN(n6547) );
  INV_X1 U4177 ( .A(n6553), .ZN(n6552) );
  NAND2_X1 U4178 ( .A1(n4198), .A2(n4197), .ZN(U2829) );
  NOR2_X4 U4179 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4571) );
  NOR2_X4 U4180 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4545) );
  AOI22_X1 U4181 ( .A1(n3360), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3199) );
  AND2_X4 U4182 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4534) );
  AND2_X4 U4183 ( .A1(n3201), .A2(n5172), .ZN(n3304) );
  AND2_X4 U4184 ( .A1(n3201), .A2(n4571), .ZN(n3346) );
  AOI22_X1 U4185 ( .A1(n3304), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3197) );
  AOI22_X1 U4186 ( .A1(n3349), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3196) );
  AOI22_X1 U4187 ( .A1(n3350), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3205) );
  AND2_X4 U4188 ( .A1(n3201), .A2(n5176), .ZN(n3384) );
  AOI22_X1 U4189 ( .A1(n3367), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3384), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3204) );
  AOI22_X1 U4190 ( .A1(n3302), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3366), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3203) );
  AND2_X4 U4191 ( .A1(n3201), .A2(n4534), .ZN(n3368) );
  AND2_X4 U4192 ( .A1(n4545), .A2(n4534), .ZN(n3298) );
  AOI22_X1 U4193 ( .A1(n3368), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3202) );
  NAND2_X2 U4194 ( .A1(n3207), .A2(n3206), .ZN(n3376) );
  NAND2_X1 U4195 ( .A1(n3827), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3211) );
  NAND2_X1 U4196 ( .A1(n3347), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3210) );
  NAND2_X1 U4197 ( .A1(n3304), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3209) );
  NAND2_X1 U4198 ( .A1(n3346), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3208) );
  NAND2_X1 U4199 ( .A1(n3367), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3215) );
  NAND2_X1 U4200 ( .A1(n3384), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3214)
         );
  NAND2_X1 U4201 ( .A1(n3368), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3213)
         );
  NAND2_X1 U4202 ( .A1(n3298), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3212) );
  NAND2_X1 U4203 ( .A1(n3454), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3219) );
  NAND2_X1 U4204 ( .A1(n3302), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3218) );
  NAND2_X1 U4205 ( .A1(n3350), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3217)
         );
  NAND2_X1 U4206 ( .A1(n3366), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3216)
         );
  NAND2_X1 U4207 ( .A1(n3360), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3223) );
  NAND2_X1 U4208 ( .A1(n3349), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3222)
         );
  NAND2_X1 U4209 ( .A1(n3288), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3221) );
  NAND2_X1 U4210 ( .A1(n3103), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3220)
         );
  INV_X2 U4211 ( .A(n3403), .ZN(n3317) );
  AOI22_X1 U4212 ( .A1(n3347), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3231) );
  AOI22_X1 U4213 ( .A1(n3454), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3230) );
  AOI22_X1 U4214 ( .A1(n3367), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3368), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3229) );
  AOI22_X1 U4215 ( .A1(n3360), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3228) );
  AOI22_X1 U4216 ( .A1(n3304), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3235) );
  AOI22_X1 U4217 ( .A1(n3349), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3234) );
  AOI22_X1 U4218 ( .A1(n3384), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3233) );
  AOI22_X1 U4219 ( .A1(n3350), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3366), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3232) );
  NAND2_X1 U4220 ( .A1(n3316), .A2(n3403), .ZN(n3251) );
  AOI22_X1 U4221 ( .A1(n3304), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3241) );
  AOI22_X1 U4222 ( .A1(n3349), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3347), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3240) );
  AOI22_X1 U4223 ( .A1(n3367), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3360), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3239) );
  AOI22_X1 U4224 ( .A1(n3384), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3366), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3238) );
  NAND4_X1 U4225 ( .A1(n3241), .A2(n3240), .A3(n3239), .A4(n3238), .ZN(n3247)
         );
  AOI22_X1 U4226 ( .A1(n3350), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3245) );
  AOI22_X1 U4227 ( .A1(n3454), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3244) );
  AOI22_X1 U4228 ( .A1(n3368), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3243) );
  AOI22_X1 U4229 ( .A1(n3346), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3242) );
  NAND4_X1 U4230 ( .A1(n3245), .A2(n3244), .A3(n3243), .A4(n3242), .ZN(n3246)
         );
  OR2_X2 U4231 ( .A1(n3247), .A2(n3246), .ZN(n3472) );
  OAI21_X1 U4232 ( .B1(n3376), .B2(n3322), .A(n3248), .ZN(n4080) );
  AND2_X1 U4233 ( .A1(n3322), .A2(n3376), .ZN(n3249) );
  NOR2_X1 U4234 ( .A1(n4080), .A2(n3249), .ZN(n3329) );
  NAND2_X1 U4235 ( .A1(n3298), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3254) );
  NAND2_X1 U4236 ( .A1(n3454), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3253) );
  NAND2_X1 U4237 ( .A1(n3254), .A2(n3253), .ZN(n3258) );
  NAND2_X1 U4238 ( .A1(n3100), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3256)
         );
  NAND2_X1 U4239 ( .A1(n3288), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3255) );
  NAND2_X1 U4240 ( .A1(n3256), .A2(n3255), .ZN(n3257) );
  NAND2_X1 U4241 ( .A1(n3368), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3262)
         );
  NAND2_X1 U4242 ( .A1(n3346), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3261) );
  NAND2_X1 U4243 ( .A1(n3827), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3260) );
  NAND2_X1 U4244 ( .A1(n3305), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3259)
         );
  NAND2_X1 U4245 ( .A1(n3349), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3268)
         );
  NAND2_X1 U4246 ( .A1(n3360), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3267) );
  NAND2_X1 U4247 ( .A1(n3304), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3266) );
  NAND2_X1 U4248 ( .A1(n3347), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3265) );
  NAND2_X1 U4249 ( .A1(n3367), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3272) );
  NAND2_X1 U4250 ( .A1(n3384), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3271)
         );
  NAND2_X1 U4251 ( .A1(n3302), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3270) );
  NAND2_X1 U4252 ( .A1(n3366), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3269)
         );
  AOI22_X1 U4253 ( .A1(n3304), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3347), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3279) );
  AOI22_X1 U4254 ( .A1(n3100), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3366), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3277) );
  AOI22_X1 U4255 ( .A1(n3349), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3276) );
  AOI22_X1 U4256 ( .A1(n3360), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3283) );
  AOI22_X1 U4257 ( .A1(n3368), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3282) );
  AOI22_X1 U4258 ( .A1(n3346), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3281) );
  AOI22_X1 U4259 ( .A1(n3384), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3280) );
  NAND2_X1 U4260 ( .A1(n4083), .A2(n4202), .ZN(n3297) );
  AOI22_X1 U4261 ( .A1(n3347), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3287) );
  AOI22_X1 U4262 ( .A1(n3349), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4263 ( .A1(n3304), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4264 ( .A1(n3454), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3293) );
  AOI22_X1 U4265 ( .A1(n3384), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U4266 ( .A1(n3367), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3368), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3291) );
  AOI22_X1 U4267 ( .A1(n3302), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3366), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3290) );
  AOI22_X1 U4268 ( .A1(n3360), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3289) );
  NAND3_X2 U4269 ( .A1(n3294), .A2(n3293), .A3(n3185), .ZN(n4207) );
  XNOR2_X1 U4270 ( .A(n6504), .B(STATE_REG_2__SCAN_IN), .ZN(n4283) );
  OR2_X1 U4271 ( .A1(n3339), .A2(n4283), .ZN(n3405) );
  INV_X1 U4272 ( .A(n3405), .ZN(n3312) );
  AOI22_X1 U4273 ( .A1(n3368), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4274 ( .A1(n3350), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3454), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4275 ( .A1(n3367), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3384), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4276 ( .A1(n3304), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4277 ( .A1(n3347), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4278 ( .A1(n3360), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U4279 ( .A1(n3349), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3306) );
  OAI211_X1 U4280 ( .C1(n3312), .C2(n5139), .A(n3095), .B(n5026), .ZN(n3313)
         );
  INV_X1 U4281 ( .A(n3313), .ZN(n3314) );
  NAND3_X1 U4282 ( .A1(n3329), .A2(n3336), .A3(n3314), .ZN(n3315) );
  NAND2_X1 U4283 ( .A1(n3315), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3326) );
  NAND2_X1 U4284 ( .A1(n3472), .A2(n3376), .ZN(n3718) );
  NAND2_X2 U4285 ( .A1(n3472), .A2(n3316), .ZN(n3404) );
  OAI22_X1 U4286 ( .A1(n3331), .A2(n3718), .B1(n3404), .B2(n3317), .ZN(n3318)
         );
  NAND2_X1 U4287 ( .A1(n3318), .A2(n4746), .ZN(n3321) );
  NAND3_X1 U4288 ( .A1(n4307), .A2(n4084), .A3(n3319), .ZN(n3320) );
  NAND2_X1 U4289 ( .A1(n3321), .A2(n3320), .ZN(n3323) );
  NAND2_X1 U4290 ( .A1(n3322), .A2(n4207), .ZN(n3332) );
  NAND2_X2 U4291 ( .A1(n3323), .A2(n3332), .ZN(n3406) );
  NAND2_X1 U4292 ( .A1(n3423), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3328) );
  NAND2_X1 U4293 ( .A1(n5881), .A2(n6586), .ZN(n4422) );
  MUX2_X1 U4294 ( .A(n4422), .B(n4095), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3327) );
  NAND2_X1 U4295 ( .A1(n3328), .A2(n3327), .ZN(n3402) );
  INV_X1 U4296 ( .A(n3329), .ZN(n3330) );
  OAI21_X1 U4297 ( .B1(n3330), .B2(n4623), .A(n4510), .ZN(n3344) );
  INV_X1 U4298 ( .A(n4097), .ZN(n3335) );
  NAND2_X1 U4299 ( .A1(n3332), .A2(n4202), .ZN(n3334) );
  NAND2_X1 U4300 ( .A1(n5881), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6486) );
  AOI21_X1 U4301 ( .B1(n3099), .B2(n4084), .A(n6486), .ZN(n3333) );
  OAI211_X1 U4302 ( .C1(n3335), .C2(n3331), .A(n3334), .B(n3333), .ZN(n3338)
         );
  INV_X1 U4303 ( .A(n3336), .ZN(n3337) );
  INV_X1 U4304 ( .A(n5026), .ZN(n4386) );
  AND2_X1 U4305 ( .A1(n4386), .A2(n3341), .ZN(n3342) );
  NAND3_X1 U4306 ( .A1(n3344), .A2(n3343), .A3(n4089), .ZN(n3401) );
  INV_X1 U4307 ( .A(n3401), .ZN(n3345) );
  AOI22_X1 U4308 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4008), .B1(n4009), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4309 ( .A1(n3348), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4310 ( .A1(n4013), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3352) );
  INV_X1 U4311 ( .A(n3350), .ZN(n3390) );
  AOI22_X1 U4312 ( .A1(n3984), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4011), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3351) );
  INV_X1 U4313 ( .A(n3454), .ZN(n3361) );
  AOI22_X1 U4314 ( .A1(n4007), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3358) );
  INV_X1 U4315 ( .A(n3827), .ZN(n3354) );
  INV_X2 U4316 ( .A(n3354), .ZN(n3938) );
  AOI22_X1 U4317 ( .A1(n3304), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3357) );
  AOI22_X1 U4318 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n3999), .B1(n3366), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3356) );
  AOI22_X1 U4319 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n3985), .B1(n4002), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3355) );
  NAND3_X1 U4320 ( .A1(n3359), .A2(n3193), .A3(n3187), .ZN(n4219) );
  INV_X1 U4321 ( .A(n4219), .ZN(n3375) );
  AOI22_X1 U4322 ( .A1(n4011), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3999), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3365) );
  AOI22_X1 U4323 ( .A1(n3348), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4324 ( .A1(n3304), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4009), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3363) );
  AOI22_X1 U4325 ( .A1(n4000), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3362) );
  NAND4_X1 U4326 ( .A1(n3365), .A2(n3364), .A3(n3363), .A4(n3362), .ZN(n3374)
         );
  AOI22_X1 U4327 ( .A1(n4008), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3372) );
  AOI22_X1 U4328 ( .A1(n4007), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3366), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3371) );
  AOI22_X1 U4329 ( .A1(n3984), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4330 ( .A1(n3985), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3369) );
  NAND4_X1 U4331 ( .A1(n3372), .A2(n3371), .A3(n3370), .A4(n3369), .ZN(n3373)
         );
  XNOR2_X1 U4332 ( .A(n3375), .B(n4264), .ZN(n3378) );
  INV_X1 U4333 ( .A(n3376), .ZN(n3377) );
  NAND2_X1 U4334 ( .A1(n3378), .A2(n4199), .ZN(n3488) );
  INV_X1 U4335 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3381) );
  AOI21_X1 U4336 ( .B1(n3377), .B2(n4264), .A(n6586), .ZN(n3380) );
  NAND2_X1 U4337 ( .A1(n3324), .A2(n4219), .ZN(n3379) );
  OAI211_X1 U4338 ( .C1(n4049), .C2(n3381), .A(n3380), .B(n3379), .ZN(n3489)
         );
  NAND2_X1 U4339 ( .A1(n4199), .A2(n4264), .ZN(n3382) );
  NAND2_X1 U4340 ( .A1(n4068), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4341 ( .A1(n3984), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4007), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3389) );
  AOI22_X1 U4342 ( .A1(n4008), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4343 ( .A1(n3348), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3387) );
  AOI22_X1 U4344 ( .A1(n4013), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3386) );
  NAND4_X1 U4345 ( .A1(n3389), .A2(n3388), .A3(n3387), .A4(n3386), .ZN(n3396)
         );
  AOI22_X1 U4346 ( .A1(n4011), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4347 ( .A1(n4001), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4009), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3393) );
  INV_X2 U4348 ( .A(n3979), .ZN(n4010) );
  AOI22_X1 U4349 ( .A1(n3999), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3392) );
  AOI22_X1 U4350 ( .A1(n3985), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3391) );
  NAND4_X1 U4351 ( .A1(n3394), .A2(n3393), .A3(n3392), .A4(n3391), .ZN(n3395)
         );
  NAND2_X1 U4352 ( .A1(n3441), .A2(n4212), .ZN(n3399) );
  INV_X1 U4353 ( .A(n4264), .ZN(n3397) );
  NAND2_X1 U4354 ( .A1(n4199), .A2(n3397), .ZN(n3398) );
  AOI21_X1 U4355 ( .B1(n4348), .B2(n3405), .A(n4326), .ZN(n3408) );
  NAND2_X1 U4356 ( .A1(n3408), .A2(n4309), .ZN(n3409) );
  NAND2_X1 U4357 ( .A1(n3409), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3413) );
  INV_X1 U4358 ( .A(n3413), .ZN(n3410) );
  XNOR2_X1 U4359 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4689) );
  OAI22_X1 U4360 ( .A1(n4422), .A2(n4689), .B1(n4095), .B2(n6456), .ZN(n3411)
         );
  NAND2_X1 U4361 ( .A1(n3410), .A2(n3180), .ZN(n3414) );
  XNOR2_X2 U4362 ( .A(n3421), .B(n3422), .ZN(n4580) );
  INV_X1 U4363 ( .A(n3416), .ZN(n3417) );
  NOR2_X1 U4364 ( .A1(n3418), .A2(n3417), .ZN(n3419) );
  OAI21_X2 U4365 ( .B1(n3422), .B2(n3421), .A(n3420), .ZN(n3444) );
  NAND2_X1 U4366 ( .A1(n3423), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3428) );
  INV_X1 U4367 ( .A(n4422), .ZN(n3449) );
  AND2_X1 U4368 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3424) );
  NAND2_X1 U4369 ( .A1(n3424), .A2(n6334), .ZN(n6382) );
  INV_X1 U4370 ( .A(n3424), .ZN(n3425) );
  NAND2_X1 U4371 ( .A1(n3425), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3426) );
  NAND2_X1 U4372 ( .A1(n6382), .A2(n3426), .ZN(n4621) );
  INV_X1 U4373 ( .A(n4095), .ZN(n3448) );
  AOI22_X1 U4374 ( .A1(n3449), .A2(n4621), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3448), .ZN(n3427) );
  NAND2_X1 U4375 ( .A1(n3428), .A2(n3427), .ZN(n3445) );
  XNOR2_X1 U4376 ( .A(n3444), .B(n3445), .ZN(n4522) );
  NAND2_X1 U4377 ( .A1(n4522), .A2(n6586), .ZN(n3440) );
  AOI22_X1 U4378 ( .A1(n3984), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4007), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3432) );
  AOI22_X1 U4379 ( .A1(n4011), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4380 ( .A1(n3999), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4381 ( .A1(n3985), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3429) );
  NAND4_X1 U4382 ( .A1(n3432), .A2(n3431), .A3(n3430), .A4(n3429), .ZN(n3438)
         );
  INV_X1 U4383 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n6728) );
  AOI22_X1 U4384 ( .A1(n4009), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3436) );
  AOI22_X1 U4385 ( .A1(n4001), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3435) );
  AOI22_X1 U4386 ( .A1(n3348), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3434) );
  AOI22_X1 U4387 ( .A1(n4013), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3433) );
  NAND4_X1 U4388 ( .A1(n3436), .A2(n3435), .A3(n3434), .A4(n3433), .ZN(n3437)
         );
  NAND2_X1 U4389 ( .A1(n4199), .A2(n4206), .ZN(n3439) );
  AOI22_X1 U4390 ( .A1(n4068), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3441), 
        .B2(n4206), .ZN(n3442) );
  NAND2_X1 U4391 ( .A1(n3479), .A2(n3477), .ZN(n3469) );
  INV_X1 U4392 ( .A(n3469), .ZN(n3467) );
  INV_X1 U4393 ( .A(n3444), .ZN(n3446) );
  NAND2_X1 U4394 ( .A1(n3423), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3451) );
  NOR3_X1 U4395 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6334), .A3(n6456), 
        .ZN(n6307) );
  NAND2_X1 U4396 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6307), .ZN(n6299) );
  NAND2_X1 U4397 ( .A1(n6460), .A2(n6299), .ZN(n3447) );
  NOR3_X1 U4398 ( .A1(n6460), .A2(n6334), .A3(n6456), .ZN(n4772) );
  NAND2_X1 U4399 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4772), .ZN(n4768) );
  AOI22_X1 U4400 ( .A1(n3449), .A2(n4690), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3448), .ZN(n3450) );
  NAND2_X1 U4401 ( .A1(n6333), .A2(n6586), .ZN(n3466) );
  INV_X1 U4402 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n6627) );
  AOI22_X1 U4403 ( .A1(n3984), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4007), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3458) );
  INV_X2 U4404 ( .A(n3361), .ZN(n4000) );
  AOI22_X1 U4405 ( .A1(n4011), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3457) );
  AOI22_X1 U4406 ( .A1(n3999), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3456) );
  AOI22_X1 U4407 ( .A1(n3985), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3455) );
  NAND4_X1 U4408 ( .A1(n3458), .A2(n3457), .A3(n3456), .A4(n3455), .ZN(n3464)
         );
  AOI22_X1 U4409 ( .A1(n4009), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3462) );
  AOI22_X1 U4410 ( .A1(n4001), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3461) );
  AOI22_X1 U4411 ( .A1(n3348), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3460) );
  AOI22_X1 U4412 ( .A1(n4013), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3459) );
  NAND4_X1 U4413 ( .A1(n3462), .A2(n3461), .A3(n3460), .A4(n3459), .ZN(n3463)
         );
  AOI22_X1 U4414 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n4068), .B1(n4073), 
        .B2(n4232), .ZN(n3465) );
  NOR2_X2 U4415 ( .A1(n3331), .A2(n6583), .ZN(n3708) );
  NAND2_X1 U4416 ( .A1(n3319), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3526) );
  INV_X1 U4417 ( .A(n3497), .ZN(n3471) );
  INV_X1 U4418 ( .A(n3519), .ZN(n3520) );
  OAI21_X1 U4419 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3471), .A(n3520), 
        .ZN(n5041) );
  NAND2_X1 U4420 ( .A1(n6583), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4421 ( .A1(n4031), .A2(n5041), .B1(n5150), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3474) );
  NAND2_X1 U4422 ( .A1(n3952), .A2(EAX_REG_3__SCAN_IN), .ZN(n3473) );
  OAI211_X1 U4423 ( .C1(n3526), .C2(n3470), .A(n3474), .B(n3473), .ZN(n3475)
         );
  AOI21_X1 U4424 ( .B1(n3476), .B2(n3708), .A(n3475), .ZN(n4445) );
  INV_X1 U4425 ( .A(n4445), .ZN(n3505) );
  INV_X1 U4426 ( .A(n3477), .ZN(n3478) );
  XNOR2_X1 U4427 ( .A(n3479), .B(n3478), .ZN(n4575) );
  NAND2_X1 U4428 ( .A1(n4575), .A2(n3708), .ZN(n3480) );
  NAND2_X1 U4429 ( .A1(n3480), .A2(n3880), .ZN(n4449) );
  NAND2_X1 U4430 ( .A1(n4576), .A2(n3708), .ZN(n3487) );
  NAND2_X1 U4431 ( .A1(n6583), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3484)
         );
  NAND2_X1 U4432 ( .A1(n3543), .A2(EAX_REG_1__SCAN_IN), .ZN(n3483) );
  OAI211_X1 U4433 ( .C1(n3526), .C2(n3195), .A(n3484), .B(n3483), .ZN(n3485)
         );
  INV_X1 U4434 ( .A(n3485), .ZN(n3486) );
  NAND2_X1 U4435 ( .A1(n3487), .A2(n3486), .ZN(n4498) );
  NAND2_X2 U4436 ( .A1(n3492), .A2(n3491), .ZN(n5728) );
  AOI21_X1 U4437 ( .B1(n6226), .B2(n3493), .A(n6583), .ZN(n4398) );
  NAND2_X1 U4438 ( .A1(n3102), .A2(n3708), .ZN(n3496) );
  AOI22_X1 U4439 ( .A1(n3543), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6583), .ZN(n3495) );
  OAI211_X1 U4440 ( .C1(n3526), .C2(n5107), .A(n3496), .B(n3495), .ZN(n4397)
         );
  MUX2_X1 U4441 ( .A(n3969), .B(n4398), .S(n4397), .Z(n4499) );
  NAND2_X1 U4442 ( .A1(n4449), .A2(n4496), .ZN(n3504) );
  INV_X1 U4443 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3499) );
  OAI21_X1 U4444 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3497), .ZN(n6107) );
  NAND2_X1 U4445 ( .A1(n3969), .A2(n6107), .ZN(n3498) );
  OAI21_X1 U4446 ( .B1(n3880), .B2(n3499), .A(n3498), .ZN(n3500) );
  AOI21_X1 U4447 ( .B1(n3952), .B2(EAX_REG_2__SCAN_IN), .A(n3500), .ZN(n3503)
         );
  INV_X1 U4448 ( .A(n3526), .ZN(n3501) );
  NAND2_X1 U4449 ( .A1(n3501), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3502) );
  AND2_X1 U4450 ( .A1(n3503), .A2(n3502), .ZN(n4447) );
  NAND2_X1 U4451 ( .A1(n3504), .A2(n4447), .ZN(n4444) );
  NAND2_X1 U4452 ( .A1(n4068), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U4453 ( .A1(n3984), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4007), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3509) );
  AOI22_X1 U4454 ( .A1(n4011), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3508) );
  AOI22_X1 U4455 ( .A1(n3999), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3507) );
  AOI22_X1 U4456 ( .A1(n3985), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3506) );
  NAND4_X1 U4457 ( .A1(n3509), .A2(n3508), .A3(n3507), .A4(n3506), .ZN(n3515)
         );
  AOI22_X1 U4458 ( .A1(n4009), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4459 ( .A1(n4001), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4460 ( .A1(n3348), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3511) );
  AOI22_X1 U4461 ( .A1(n4013), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3510) );
  NAND4_X1 U4462 ( .A1(n3513), .A2(n3512), .A3(n3511), .A4(n3510), .ZN(n3514)
         );
  NAND2_X1 U4463 ( .A1(n4073), .A2(n4246), .ZN(n3516) );
  INV_X1 U4464 ( .A(n4235), .ZN(n3518) );
  NAND2_X1 U4465 ( .A1(n3518), .A2(n3708), .ZN(n3529) );
  INV_X1 U4466 ( .A(n3568), .ZN(n3523) );
  INV_X1 U4467 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3521) );
  NAND2_X1 U4468 ( .A1(n3521), .A2(n3520), .ZN(n3522) );
  NAND2_X1 U4469 ( .A1(n3523), .A2(n3522), .ZN(n6096) );
  INV_X1 U4470 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6584) );
  OAI21_X1 U4471 ( .B1(n6584), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6583), 
        .ZN(n3525) );
  NAND2_X1 U4472 ( .A1(n3952), .A2(EAX_REG_4__SCAN_IN), .ZN(n3524) );
  OAI211_X1 U4473 ( .C1(n3526), .C2(n5885), .A(n3525), .B(n3524), .ZN(n3527)
         );
  OAI21_X1 U4474 ( .B1(n4025), .B2(n6096), .A(n3527), .ZN(n3528) );
  NAND2_X1 U4475 ( .A1(n3529), .A2(n3528), .ZN(n4507) );
  NOR2_X1 U4476 ( .A1(n3549), .A2(n3550), .ZN(n3542) );
  INV_X1 U4477 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4478 ( .A1(n3984), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4007), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3533) );
  AOI22_X1 U4479 ( .A1(n4011), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3532) );
  AOI22_X1 U4480 ( .A1(n3999), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3531) );
  AOI22_X1 U4481 ( .A1(n3985), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3530) );
  NAND4_X1 U4482 ( .A1(n3533), .A2(n3532), .A3(n3531), .A4(n3530), .ZN(n3539)
         );
  INV_X1 U4483 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n6843) );
  AOI22_X1 U4484 ( .A1(n4009), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4485 ( .A1(n4001), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3536) );
  AOI22_X1 U4486 ( .A1(n3348), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3535) );
  AOI22_X1 U4487 ( .A1(n4013), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3534) );
  NAND4_X1 U4488 ( .A1(n3537), .A2(n3536), .A3(n3535), .A4(n3534), .ZN(n3538)
         );
  NAND2_X1 U4489 ( .A1(n4073), .A2(n4245), .ZN(n3540) );
  XNOR2_X1 U4490 ( .A(n3542), .B(n3552), .ZN(n4241) );
  INV_X1 U4491 ( .A(n4241), .ZN(n3547) );
  INV_X1 U4492 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3545) );
  XNOR2_X1 U4493 ( .A(n3568), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5971) );
  AOI22_X1 U4494 ( .A1(n5971), .A2(n3969), .B1(n5150), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3544) );
  OAI21_X1 U4495 ( .B1(n4026), .B2(n3545), .A(n3544), .ZN(n3546) );
  INV_X1 U4496 ( .A(n4655), .ZN(n3548) );
  INV_X1 U4497 ( .A(n3578), .ZN(n3567) );
  NAND2_X1 U4498 ( .A1(n4068), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4499 ( .A1(n3984), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4007), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U4500 ( .A1(n4011), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3556) );
  AOI22_X1 U4501 ( .A1(n3999), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3555) );
  AOI22_X1 U4502 ( .A1(n3985), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3554) );
  NAND4_X1 U4503 ( .A1(n3557), .A2(n3556), .A3(n3555), .A4(n3554), .ZN(n3563)
         );
  AOI22_X1 U4504 ( .A1(n4009), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4505 ( .A1(n4001), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4506 ( .A1(n3348), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U4507 ( .A1(n4013), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3558) );
  NAND4_X1 U4508 ( .A1(n3561), .A2(n3560), .A3(n3559), .A4(n3558), .ZN(n3562)
         );
  NAND2_X1 U4509 ( .A1(n4073), .A2(n4256), .ZN(n3564) );
  INV_X1 U4510 ( .A(n3577), .ZN(n3566) );
  NAND2_X1 U4511 ( .A1(n3567), .A2(n3566), .ZN(n4249) );
  INV_X1 U4512 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3574) );
  AND2_X1 U4513 ( .A1(n3569), .A2(n3571), .ZN(n3570) );
  OR2_X1 U4514 ( .A1(n3570), .A2(n3595), .ZN(n6087) );
  NOR2_X1 U4515 ( .A1(n3880), .A2(n3571), .ZN(n3572) );
  AOI21_X1 U4516 ( .B1(n6087), .B2(n3969), .A(n3572), .ZN(n3573) );
  OAI21_X1 U4517 ( .B1(n4026), .B2(n3574), .A(n3573), .ZN(n3575) );
  INV_X1 U4518 ( .A(n3576), .ZN(n4608) );
  AOI22_X1 U4519 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n4068), .B1(n4073), 
        .B2(n4264), .ZN(n3579) );
  XNOR2_X1 U4520 ( .A(n4251), .B(n3579), .ZN(n4261) );
  INV_X1 U4521 ( .A(n4261), .ZN(n3584) );
  INV_X1 U4522 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3582) );
  XNOR2_X1 U4523 ( .A(n3595), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4859) );
  INV_X1 U4524 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4819) );
  NOR2_X1 U4525 ( .A1(n3880), .A2(n4819), .ZN(n3580) );
  AOI21_X1 U4526 ( .B1(n4859), .B2(n3969), .A(n3580), .ZN(n3581) );
  OAI21_X1 U4527 ( .B1(n4026), .B2(n3582), .A(n3581), .ZN(n3583) );
  NOR2_X2 U4528 ( .A1(n4608), .A2(n4614), .ZN(n4674) );
  AOI22_X1 U4529 ( .A1(n4011), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3588) );
  AOI22_X1 U4530 ( .A1(n3999), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4531 ( .A1(n3348), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4532 ( .A1(n3938), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3585) );
  NAND4_X1 U4533 ( .A1(n3588), .A2(n3587), .A3(n3586), .A4(n3585), .ZN(n3594)
         );
  AOI22_X1 U4534 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n4007), .B1(n3984), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3592) );
  AOI22_X1 U4535 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n4009), .B1(n4013), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4536 ( .A1(n4001), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3590) );
  AOI22_X1 U4537 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n3985), .B1(n3959), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3589) );
  NAND4_X1 U4538 ( .A1(n3592), .A2(n3591), .A3(n3590), .A4(n3589), .ZN(n3593)
         );
  OAI21_X1 U4539 ( .B1(n3594), .B2(n3593), .A(n3708), .ZN(n3599) );
  NAND2_X1 U4540 ( .A1(n3952), .A2(EAX_REG_8__SCAN_IN), .ZN(n3598) );
  XNOR2_X1 U4541 ( .A(n3600), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4973) );
  NAND2_X1 U4542 ( .A1(n4973), .A2(n3969), .ZN(n3597) );
  NAND2_X1 U4543 ( .A1(n5150), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3596)
         );
  NAND4_X1 U4544 ( .A1(n3599), .A2(n3598), .A3(n3597), .A4(n3596), .ZN(n4673)
         );
  NAND2_X1 U4545 ( .A1(n4674), .A2(n4673), .ZN(n4672) );
  INV_X1 U4546 ( .A(n4672), .ZN(n3618) );
  AOI21_X1 U4547 ( .B1(n6757), .B2(n3601), .A(n3633), .ZN(n5951) );
  OR2_X1 U4548 ( .A1(n5951), .A2(n4025), .ZN(n3616) );
  AOI22_X1 U4549 ( .A1(n4011), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3605) );
  AOI22_X1 U4550 ( .A1(n4001), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4009), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3604) );
  AOI22_X1 U4551 ( .A1(n3999), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3603) );
  AOI22_X1 U4552 ( .A1(n4007), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3602) );
  NAND4_X1 U4553 ( .A1(n3605), .A2(n3604), .A3(n3603), .A4(n3602), .ZN(n3611)
         );
  AOI22_X1 U4554 ( .A1(n3348), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4555 ( .A1(n4008), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3608) );
  AOI22_X1 U4556 ( .A1(n3984), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3607) );
  AOI22_X1 U4557 ( .A1(n3985), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3606) );
  NAND4_X1 U4558 ( .A1(n3609), .A2(n3608), .A3(n3607), .A4(n3606), .ZN(n3610)
         );
  OAI21_X1 U4559 ( .B1(n3611), .B2(n3610), .A(n3708), .ZN(n3614) );
  NAND2_X1 U4560 ( .A1(n3952), .A2(EAX_REG_9__SCAN_IN), .ZN(n3613) );
  NAND2_X1 U4561 ( .A1(n5150), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3612)
         );
  AND3_X1 U4562 ( .A1(n3614), .A2(n3613), .A3(n3612), .ZN(n3615) );
  NAND2_X1 U4563 ( .A1(n3618), .A2(n3617), .ZN(n4863) );
  XNOR2_X1 U4564 ( .A(n3633), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5559)
         );
  AOI22_X1 U4565 ( .A1(n4001), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4566 ( .A1(n3999), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4567 ( .A1(n4011), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4568 ( .A1(n4009), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3619) );
  NAND4_X1 U4569 ( .A1(n3622), .A2(n3621), .A3(n3620), .A4(n3619), .ZN(n3628)
         );
  AOI22_X1 U4570 ( .A1(n4007), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4571 ( .A1(n3984), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3985), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4572 ( .A1(n4013), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4573 ( .A1(n3348), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3623) );
  NAND4_X1 U4574 ( .A1(n3626), .A2(n3625), .A3(n3624), .A4(n3623), .ZN(n3627)
         );
  OAI21_X1 U4575 ( .B1(n3628), .B2(n3627), .A(n3708), .ZN(n3631) );
  NAND2_X1 U4576 ( .A1(n3952), .A2(EAX_REG_10__SCAN_IN), .ZN(n3630) );
  NAND2_X1 U4577 ( .A1(n5150), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3629)
         );
  NAND3_X1 U4578 ( .A1(n3631), .A2(n3630), .A3(n3629), .ZN(n3632) );
  AOI21_X1 U4579 ( .B1(n5559), .B2(n3969), .A(n3632), .ZN(n4864) );
  OR2_X2 U4580 ( .A1(n4863), .A2(n4864), .ZN(n5371) );
  XOR2_X1 U4581 ( .A(n5938), .B(n3649), .Z(n6073) );
  INV_X1 U4582 ( .A(n6073), .ZN(n3648) );
  AOI22_X1 U4583 ( .A1(n4009), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4584 ( .A1(n4000), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3636) );
  AOI22_X1 U4585 ( .A1(n3984), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3635) );
  AOI22_X1 U4586 ( .A1(n3985), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3634) );
  NAND4_X1 U4587 ( .A1(n3637), .A2(n3636), .A3(n3635), .A4(n3634), .ZN(n3643)
         );
  AOI22_X1 U4588 ( .A1(n4011), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3999), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4589 ( .A1(n3348), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4590 ( .A1(n4001), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4591 ( .A1(n4007), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3638) );
  NAND4_X1 U4592 ( .A1(n3641), .A2(n3640), .A3(n3639), .A4(n3638), .ZN(n3642)
         );
  OAI21_X1 U4593 ( .B1(n3643), .B2(n3642), .A(n3708), .ZN(n3646) );
  NAND2_X1 U4594 ( .A1(n3952), .A2(EAX_REG_11__SCAN_IN), .ZN(n3645) );
  NAND2_X1 U4595 ( .A1(n5150), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3644)
         );
  NAND3_X1 U4596 ( .A1(n3646), .A2(n3645), .A3(n3644), .ZN(n3647) );
  AOI21_X1 U4597 ( .B1(n3648), .B2(n3969), .A(n3647), .ZN(n5370) );
  NAND2_X1 U4598 ( .A1(n3650), .A2(n6870), .ZN(n3652) );
  INV_X1 U4599 ( .A(n3692), .ZN(n3651) );
  NAND2_X1 U4600 ( .A1(n3652), .A2(n3651), .ZN(n5931) );
  AND2_X1 U4601 ( .A1(n3952), .A2(EAX_REG_12__SCAN_IN), .ZN(n3653) );
  OAI22_X1 U4602 ( .A1(n5931), .A2(n4025), .B1(n3654), .B2(n3653), .ZN(n3666)
         );
  AOI22_X1 U4603 ( .A1(n4001), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4604 ( .A1(n3999), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4605 ( .A1(n3348), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4606 ( .A1(n4013), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3655) );
  NAND4_X1 U4607 ( .A1(n3658), .A2(n3657), .A3(n3656), .A4(n3655), .ZN(n3664)
         );
  AOI22_X1 U4608 ( .A1(n4011), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4609 ( .A1(n3984), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4007), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3661) );
  AOI22_X1 U4610 ( .A1(n4009), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4611 ( .A1(n3985), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3659) );
  NAND4_X1 U4612 ( .A1(n3662), .A2(n3661), .A3(n3660), .A4(n3659), .ZN(n3663)
         );
  OAI21_X1 U4613 ( .B1(n3664), .B2(n3663), .A(n3708), .ZN(n3665) );
  NAND2_X1 U4614 ( .A1(n3666), .A2(n3665), .ZN(n5411) );
  INV_X1 U4615 ( .A(n3708), .ZN(n3681) );
  AOI22_X1 U4616 ( .A1(n4007), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4617 ( .A1(n4013), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3985), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4618 ( .A1(n4001), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4619 ( .A1(n4009), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3667) );
  NAND4_X1 U4620 ( .A1(n3670), .A2(n3669), .A3(n3668), .A4(n3667), .ZN(n3676)
         );
  AOI22_X1 U4621 ( .A1(n3984), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4011), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3674) );
  AOI22_X1 U4622 ( .A1(n3348), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3673) );
  AOI22_X1 U4623 ( .A1(n3999), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4624 ( .A1(n4002), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3671) );
  NAND4_X1 U4625 ( .A1(n3674), .A2(n3673), .A3(n3672), .A4(n3671), .ZN(n3675)
         );
  NOR2_X1 U4626 ( .A1(n3676), .A2(n3675), .ZN(n3680) );
  XOR2_X1 U4627 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n3692), .Z(n5918) );
  INV_X1 U4628 ( .A(n5918), .ZN(n3677) );
  AOI22_X1 U4629 ( .A1(n5150), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .B1(n4031), 
        .B2(n3677), .ZN(n3679) );
  NAND2_X1 U4630 ( .A1(n3952), .A2(EAX_REG_13__SCAN_IN), .ZN(n3678) );
  OAI211_X1 U4631 ( .C1(n3681), .C2(n3680), .A(n3679), .B(n3678), .ZN(n5053)
         );
  AOI22_X1 U4632 ( .A1(n3984), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3999), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4633 ( .A1(n4009), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4634 ( .A1(n3985), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4635 ( .A1(n4002), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3682) );
  NAND4_X1 U4636 ( .A1(n3685), .A2(n3684), .A3(n3683), .A4(n3682), .ZN(n3691)
         );
  AOI22_X1 U4637 ( .A1(n4007), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4638 ( .A1(n3348), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3688) );
  AOI22_X1 U4639 ( .A1(n4001), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4640 ( .A1(n4011), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3686) );
  NAND4_X1 U4641 ( .A1(n3689), .A2(n3688), .A3(n3687), .A4(n3686), .ZN(n3690)
         );
  OAI21_X1 U4642 ( .B1(n3691), .B2(n3690), .A(n3708), .ZN(n3696) );
  INV_X1 U4643 ( .A(n3699), .ZN(n3693) );
  XNOR2_X1 U4644 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3693), .ZN(n5290)
         );
  AOI22_X1 U4645 ( .A1(n4031), .A2(n5290), .B1(n5150), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3695) );
  NAND2_X1 U4646 ( .A1(n3952), .A2(EAX_REG_14__SCAN_IN), .ZN(n3694) );
  XOR2_X1 U4647 ( .A(n3716), .B(n3717), .Z(n5530) );
  INV_X1 U4648 ( .A(n5530), .ZN(n3715) );
  AOI22_X1 U4649 ( .A1(n3348), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4650 ( .A1(n4009), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4651 ( .A1(n4000), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4652 ( .A1(n4007), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3700) );
  NAND4_X1 U4653 ( .A1(n3703), .A2(n3702), .A3(n3701), .A4(n3700), .ZN(n3710)
         );
  AOI22_X1 U4654 ( .A1(n4011), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3999), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3707) );
  AOI22_X1 U4655 ( .A1(n3984), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3985), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3706) );
  AOI22_X1 U4656 ( .A1(n4001), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4657 ( .A1(n4002), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3704) );
  NAND4_X1 U4658 ( .A1(n3707), .A2(n3706), .A3(n3705), .A4(n3704), .ZN(n3709)
         );
  OAI21_X1 U4659 ( .B1(n3710), .B2(n3709), .A(n3708), .ZN(n3713) );
  NAND2_X1 U4660 ( .A1(n3952), .A2(EAX_REG_15__SCAN_IN), .ZN(n3712) );
  NAND2_X1 U4661 ( .A1(n5150), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3711)
         );
  NAND3_X1 U4662 ( .A1(n3713), .A2(n3712), .A3(n3711), .ZN(n3714) );
  AOI21_X1 U4663 ( .B1(n3715), .B2(n3969), .A(n3714), .ZN(n5276) );
  XNOR2_X1 U4664 ( .A(n3736), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5262)
         );
  NAND2_X1 U4665 ( .A1(n5262), .A2(n4031), .ZN(n3733) );
  AOI22_X1 U4666 ( .A1(n4011), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4667 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4007), .B1(n3984), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4668 ( .A1(n3348), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4669 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n4001), .B1(n4009), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3719) );
  NAND4_X1 U4670 ( .A1(n3722), .A2(n3721), .A3(n3720), .A4(n3719), .ZN(n3728)
         );
  AOI22_X1 U4671 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n3827), .B1(n4008), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4672 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n3999), .B1(n4010), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4673 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n3985), .B1(n3959), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4674 ( .A1(n4002), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3723) );
  NAND4_X1 U4675 ( .A1(n3726), .A2(n3725), .A3(n3724), .A4(n3723), .ZN(n3727)
         );
  OR2_X1 U4676 ( .A1(n3728), .A2(n3727), .ZN(n3731) );
  INV_X1 U4677 ( .A(EAX_REG_16__SCAN_IN), .ZN(n3729) );
  INV_X1 U4678 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5519) );
  OAI22_X1 U4679 ( .A1(n4026), .A2(n3729), .B1(n3880), .B2(n5519), .ZN(n3730)
         );
  AOI21_X1 U4680 ( .B1(n4028), .B2(n3731), .A(n3730), .ZN(n3732) );
  NAND2_X1 U4681 ( .A1(n3733), .A2(n3732), .ZN(n5261) );
  NAND2_X1 U4682 ( .A1(n3736), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3734)
         );
  INV_X1 U4683 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U4684 ( .A1(n3734), .A2(n5908), .ZN(n3737) );
  NAND2_X1 U4685 ( .A1(n3737), .A2(n3769), .ZN(n5916) );
  AOI22_X1 U4686 ( .A1(n4000), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3999), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3741) );
  AOI22_X1 U4687 ( .A1(n3348), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3985), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4688 ( .A1(n4013), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4689 ( .A1(n4007), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3738) );
  NAND4_X1 U4690 ( .A1(n3741), .A2(n3740), .A3(n3739), .A4(n3738), .ZN(n3747)
         );
  AOI22_X1 U4691 ( .A1(n4001), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3745) );
  AOI22_X1 U4692 ( .A1(n4011), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4693 ( .A1(n3984), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4694 ( .A1(n4009), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3742) );
  NAND4_X1 U4695 ( .A1(n3745), .A2(n3744), .A3(n3743), .A4(n3742), .ZN(n3746)
         );
  NOR2_X1 U4696 ( .A1(n3747), .A2(n3746), .ZN(n3750) );
  OAI21_X1 U4697 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6584), .A(n6583), 
        .ZN(n3749) );
  NAND2_X1 U4698 ( .A1(n3952), .A2(EAX_REG_17__SCAN_IN), .ZN(n3748) );
  OAI211_X1 U4699 ( .C1(n3996), .C2(n3750), .A(n3749), .B(n3748), .ZN(n3751)
         );
  OR2_X1 U4700 ( .A1(n3770), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3753)
         );
  NAND2_X1 U4701 ( .A1(n3786), .A2(n3753), .ZN(n5854) );
  AOI22_X1 U4702 ( .A1(n4011), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3999), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3757) );
  AOI22_X1 U4703 ( .A1(n3984), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4704 ( .A1(n3985), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4705 ( .A1(n4008), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3754) );
  NAND4_X1 U4706 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3763)
         );
  AOI22_X1 U4707 ( .A1(n3348), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4708 ( .A1(n4001), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4709 ( .A1(n4007), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4710 ( .A1(n4009), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3758) );
  NAND4_X1 U4711 ( .A1(n3761), .A2(n3760), .A3(n3759), .A4(n3758), .ZN(n3762)
         );
  NOR2_X1 U4712 ( .A1(n3763), .A2(n3762), .ZN(n3766) );
  OAI21_X1 U4713 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6584), .A(n6583), 
        .ZN(n3765) );
  NAND2_X1 U4714 ( .A1(n3952), .A2(EAX_REG_19__SCAN_IN), .ZN(n3764) );
  OAI211_X1 U4715 ( .C1(n3996), .C2(n3766), .A(n3765), .B(n3764), .ZN(n3767)
         );
  NAND2_X1 U4716 ( .A1(n3768), .A2(n3767), .ZN(n5351) );
  AND2_X1 U4717 ( .A1(n3769), .A2(n6615), .ZN(n3771) );
  OR2_X1 U4718 ( .A1(n3771), .A2(n3770), .ZN(n5504) );
  AOI22_X1 U4719 ( .A1(n4011), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4720 ( .A1(n4008), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4721 ( .A1(n3999), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4722 ( .A1(n4009), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3772) );
  NAND4_X1 U4723 ( .A1(n3775), .A2(n3774), .A3(n3773), .A4(n3772), .ZN(n3781)
         );
  AOI22_X1 U4724 ( .A1(n3984), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4007), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4725 ( .A1(n4001), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4726 ( .A1(n3985), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4727 ( .A1(n3348), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3776) );
  NAND4_X1 U4728 ( .A1(n3779), .A2(n3778), .A3(n3777), .A4(n3776), .ZN(n3780)
         );
  NOR2_X1 U4729 ( .A1(n3781), .A2(n3780), .ZN(n3784) );
  OAI21_X1 U4730 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6615), .A(n4025), .ZN(
        n3782) );
  AOI21_X1 U4731 ( .B1(n3952), .B2(EAX_REG_18__SCAN_IN), .A(n3782), .ZN(n3783)
         );
  OAI21_X1 U4732 ( .B1(n3996), .B2(n3784), .A(n3783), .ZN(n3785) );
  OAI21_X1 U4733 ( .B1(n5504), .B2(n4025), .A(n3785), .ZN(n5246) );
  NAND2_X1 U4734 ( .A1(n3786), .A2(n6702), .ZN(n3787) );
  AND2_X1 U4735 ( .A1(n3803), .A2(n3787), .ZN(n5845) );
  AOI22_X1 U4736 ( .A1(n4007), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4011), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4737 ( .A1(n4009), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4738 ( .A1(n3999), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3789) );
  AOI22_X1 U4739 ( .A1(n4013), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3788) );
  NAND4_X1 U4740 ( .A1(n3791), .A2(n3790), .A3(n3789), .A4(n3788), .ZN(n3797)
         );
  AOI22_X1 U4741 ( .A1(n3984), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4742 ( .A1(n4001), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4743 ( .A1(n3985), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4744 ( .A1(n3348), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3792) );
  NAND4_X1 U4745 ( .A1(n3795), .A2(n3794), .A3(n3793), .A4(n3792), .ZN(n3796)
         );
  OR2_X1 U4746 ( .A1(n3797), .A2(n3796), .ZN(n3801) );
  INV_X1 U4747 ( .A(EAX_REG_20__SCAN_IN), .ZN(n3799) );
  NAND2_X1 U4748 ( .A1(n6583), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3798)
         );
  OAI211_X1 U4749 ( .C1(n4026), .C2(n3799), .A(n4025), .B(n3798), .ZN(n3800)
         );
  AOI21_X1 U4750 ( .B1(n4028), .B2(n3801), .A(n3800), .ZN(n3802) );
  AOI21_X1 U4751 ( .B1(n5845), .B2(n4031), .A(n3802), .ZN(n5345) );
  NAND2_X1 U4752 ( .A1(n5353), .A2(n5345), .ZN(n5344) );
  INV_X1 U4753 ( .A(n5344), .ZN(n3820) );
  NAND2_X1 U4754 ( .A1(n3803), .A2(n5829), .ZN(n3804) );
  NAND2_X1 U4755 ( .A1(n3851), .A2(n3804), .ZN(n5837) );
  AOI22_X1 U4756 ( .A1(n4007), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4011), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4757 ( .A1(n4001), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4758 ( .A1(n3984), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4759 ( .A1(n3348), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3805) );
  NAND4_X1 U4760 ( .A1(n3808), .A2(n3807), .A3(n3806), .A4(n3805), .ZN(n3814)
         );
  AOI22_X1 U4761 ( .A1(n4000), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3985), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4762 ( .A1(n4009), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4763 ( .A1(n3999), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4764 ( .A1(n4013), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3809) );
  NAND4_X1 U4765 ( .A1(n3812), .A2(n3811), .A3(n3810), .A4(n3809), .ZN(n3813)
         );
  NOR2_X1 U4766 ( .A1(n3814), .A2(n3813), .ZN(n3817) );
  OAI21_X1 U4767 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5829), .A(n4025), .ZN(
        n3815) );
  AOI21_X1 U4768 ( .B1(n3952), .B2(EAX_REG_21__SCAN_IN), .A(n3815), .ZN(n3816)
         );
  OAI21_X1 U4769 ( .B1(n3996), .B2(n3817), .A(n3816), .ZN(n3818) );
  OAI21_X1 U4770 ( .B1(n5837), .B2(n4025), .A(n3818), .ZN(n5339) );
  OR2_X1 U4771 ( .A1(n3853), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3821)
         );
  NAND2_X1 U4772 ( .A1(n3886), .A2(n3821), .ZN(n5818) );
  AOI22_X1 U4773 ( .A1(n3984), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4007), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4774 ( .A1(n4011), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3825) );
  INV_X1 U4775 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4776 ( .A1(n3999), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4777 ( .A1(n3985), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3823) );
  NAND4_X1 U4778 ( .A1(n3826), .A2(n3825), .A3(n3824), .A4(n3823), .ZN(n3833)
         );
  AOI22_X1 U4779 ( .A1(n4009), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4780 ( .A1(n4001), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3830) );
  AOI22_X1 U4781 ( .A1(n3348), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4782 ( .A1(n4013), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3828) );
  NAND4_X1 U4783 ( .A1(n3831), .A2(n3830), .A3(n3829), .A4(n3828), .ZN(n3832)
         );
  OR2_X1 U4784 ( .A1(n3833), .A2(n3832), .ZN(n3845) );
  AOI22_X1 U4785 ( .A1(n3984), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4007), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4786 ( .A1(n4011), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4787 ( .A1(n3999), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4788 ( .A1(n3985), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3834) );
  NAND4_X1 U4789 ( .A1(n3837), .A2(n3836), .A3(n3835), .A4(n3834), .ZN(n3843)
         );
  AOI22_X1 U4790 ( .A1(n4009), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4791 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4001), .B1(n4008), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4792 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n3348), .B1(n4002), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4793 ( .A1(n4013), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3838) );
  NAND4_X1 U4794 ( .A1(n3841), .A2(n3840), .A3(n3839), .A4(n3838), .ZN(n3842)
         );
  OR2_X1 U4795 ( .A1(n3843), .A2(n3842), .ZN(n3844) );
  NAND2_X1 U4796 ( .A1(n3844), .A2(n3845), .ZN(n3900) );
  OAI21_X1 U4797 ( .B1(n3845), .B2(n3844), .A(n3900), .ZN(n3846) );
  NOR2_X1 U4798 ( .A1(n3996), .A2(n3846), .ZN(n3850) );
  INV_X1 U4799 ( .A(EAX_REG_23__SCAN_IN), .ZN(n3848) );
  NAND2_X1 U4800 ( .A1(n6583), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3847)
         );
  OAI211_X1 U4801 ( .C1(n4026), .C2(n3848), .A(n4025), .B(n3847), .ZN(n3849)
         );
  OAI22_X1 U4802 ( .A1(n5818), .A2(n4025), .B1(n3850), .B2(n3849), .ZN(n5328)
         );
  AND2_X1 U4803 ( .A1(n3851), .A2(n6772), .ZN(n3852) );
  NOR2_X1 U4804 ( .A1(n3853), .A2(n3852), .ZN(n5473) );
  NAND2_X1 U4805 ( .A1(n5473), .A2(n4031), .ZN(n3868) );
  AOI22_X1 U4806 ( .A1(n3984), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4007), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3857) );
  INV_X1 U4807 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4808 ( .A1(n4011), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4809 ( .A1(n3999), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4810 ( .A1(n3985), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3854) );
  NAND4_X1 U4811 ( .A1(n3857), .A2(n3856), .A3(n3855), .A4(n3854), .ZN(n3863)
         );
  AOI22_X1 U4812 ( .A1(n4009), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4813 ( .A1(n4001), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4814 ( .A1(n3348), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4815 ( .A1(n4013), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3858) );
  NAND4_X1 U4816 ( .A1(n3861), .A2(n3860), .A3(n3859), .A4(n3858), .ZN(n3862)
         );
  NOR2_X1 U4817 ( .A1(n3863), .A2(n3862), .ZN(n3866) );
  AOI21_X1 U4818 ( .B1(n6772), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3864) );
  AOI21_X1 U4819 ( .B1(n3952), .B2(EAX_REG_22__SCAN_IN), .A(n3864), .ZN(n3865)
         );
  OAI21_X1 U4820 ( .B1(n3996), .B2(n3866), .A(n3865), .ZN(n3867) );
  NAND2_X1 U4821 ( .A1(n3868), .A2(n3867), .ZN(n5237) );
  XNOR2_X1 U4822 ( .A(n3886), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5810)
         );
  AOI22_X1 U4823 ( .A1(n3984), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4011), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4824 ( .A1(n3348), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3985), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4825 ( .A1(n4001), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4826 ( .A1(n3938), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3870) );
  NAND4_X1 U4827 ( .A1(n3873), .A2(n3872), .A3(n3871), .A4(n3870), .ZN(n3879)
         );
  AOI22_X1 U4828 ( .A1(n4007), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4829 ( .A1(n4013), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4009), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4830 ( .A1(n3999), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4831 ( .A1(n4002), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3874) );
  NAND4_X1 U4832 ( .A1(n3877), .A2(n3876), .A3(n3875), .A4(n3874), .ZN(n3878)
         );
  OR2_X1 U4833 ( .A1(n3879), .A2(n3878), .ZN(n3899) );
  XNOR2_X1 U4834 ( .A(n3900), .B(n3899), .ZN(n3883) );
  INV_X1 U4835 ( .A(EAX_REG_24__SCAN_IN), .ZN(n3881) );
  INV_X1 U4836 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5072) );
  OAI22_X1 U4837 ( .A1(n4026), .A2(n3881), .B1(n3880), .B2(n5072), .ZN(n3882)
         );
  AOI21_X1 U4838 ( .B1(n4028), .B2(n3883), .A(n3882), .ZN(n3884) );
  NAND2_X1 U4839 ( .A1(n3885), .A2(n3884), .ZN(n5077) );
  INV_X1 U4840 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3902) );
  AND2_X1 U4841 ( .A1(n3887), .A2(n3902), .ZN(n3888) );
  OR2_X1 U4842 ( .A1(n3888), .A2(n3927), .ZN(n5802) );
  AOI22_X1 U4843 ( .A1(n3984), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4007), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4844 ( .A1(n4011), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4845 ( .A1(n3999), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4846 ( .A1(n3985), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3889) );
  NAND4_X1 U4847 ( .A1(n3892), .A2(n3891), .A3(n3890), .A4(n3889), .ZN(n3898)
         );
  AOI22_X1 U4848 ( .A1(n4009), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4849 ( .A1(n4001), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4850 ( .A1(n3348), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4851 ( .A1(n4013), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3893) );
  NAND4_X1 U4852 ( .A1(n3896), .A2(n3895), .A3(n3894), .A4(n3893), .ZN(n3897)
         );
  OR2_X1 U4853 ( .A1(n3898), .A2(n3897), .ZN(n3919) );
  INV_X1 U4854 ( .A(n3899), .ZN(n3901) );
  NOR2_X1 U4855 ( .A1(n3901), .A2(n3900), .ZN(n3920) );
  XNOR2_X1 U4856 ( .A(n3919), .B(n3920), .ZN(n3905) );
  OAI21_X1 U4857 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n3902), .A(n4025), .ZN(
        n3903) );
  AOI21_X1 U4858 ( .B1(n3952), .B2(EAX_REG_25__SCAN_IN), .A(n3903), .ZN(n3904)
         );
  OAI21_X1 U4859 ( .B1(n3996), .B2(n3905), .A(n3904), .ZN(n3906) );
  OAI21_X1 U4860 ( .B1(n5802), .B2(n4025), .A(n3906), .ZN(n5317) );
  INV_X1 U4861 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5448) );
  XNOR2_X1 U4862 ( .A(n3927), .B(n5448), .ZN(n5446) );
  NAND2_X1 U4863 ( .A1(n5446), .A2(n4031), .ZN(n3926) );
  AOI22_X1 U4864 ( .A1(n3348), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4013), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4865 ( .A1(n4001), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4866 ( .A1(n3984), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4867 ( .A1(n4009), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4012), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3909) );
  NAND4_X1 U4868 ( .A1(n3912), .A2(n3911), .A3(n3910), .A4(n3909), .ZN(n3918)
         );
  AOI22_X1 U4869 ( .A1(n4011), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3999), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4870 ( .A1(n4007), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4871 ( .A1(n3985), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4872 ( .A1(n3938), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3913) );
  NAND4_X1 U4873 ( .A1(n3916), .A2(n3915), .A3(n3914), .A4(n3913), .ZN(n3917)
         );
  NOR2_X1 U4874 ( .A1(n3918), .A2(n3917), .ZN(n3933) );
  NAND2_X1 U4875 ( .A1(n3920), .A2(n3919), .ZN(n3932) );
  XOR2_X1 U4876 ( .A(n3933), .B(n3932), .Z(n3921) );
  NAND2_X1 U4877 ( .A1(n3921), .A2(n4028), .ZN(n3924) );
  OAI21_X1 U4878 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5448), .A(n4025), .ZN(
        n3922) );
  AOI21_X1 U4879 ( .B1(n3952), .B2(EAX_REG_26__SCAN_IN), .A(n3922), .ZN(n3923)
         );
  NAND2_X1 U4880 ( .A1(n3924), .A2(n3923), .ZN(n3925) );
  NAND2_X1 U4881 ( .A1(n3926), .A2(n3925), .ZN(n5228) );
  INV_X1 U4882 ( .A(n3928), .ZN(n3930) );
  INV_X1 U4883 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3929) );
  NAND2_X1 U4884 ( .A1(n3930), .A2(n3929), .ZN(n3931) );
  NAND2_X1 U4885 ( .A1(n3970), .A2(n3931), .ZN(n5790) );
  NOR2_X1 U4886 ( .A1(n3933), .A2(n3932), .ZN(n3954) );
  AOI22_X1 U4887 ( .A1(n3984), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4007), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4888 ( .A1(n4011), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4000), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3936) );
  AOI22_X1 U4889 ( .A1(n3999), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4890 ( .A1(n3985), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3934) );
  NAND4_X1 U4891 ( .A1(n3937), .A2(n3936), .A3(n3935), .A4(n3934), .ZN(n3944)
         );
  AOI22_X1 U4892 ( .A1(n4009), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4893 ( .A1(n4001), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4894 ( .A1(n3348), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3940) );
  AOI22_X1 U4895 ( .A1(n4013), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3939) );
  NAND4_X1 U4896 ( .A1(n3942), .A2(n3941), .A3(n3940), .A4(n3939), .ZN(n3943)
         );
  OR2_X1 U4897 ( .A1(n3944), .A2(n3943), .ZN(n3953) );
  XNOR2_X1 U4898 ( .A(n3954), .B(n3953), .ZN(n3948) );
  NAND2_X1 U4899 ( .A1(n6583), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n3945)
         );
  NAND2_X1 U4900 ( .A1(n4025), .A2(n3945), .ZN(n3946) );
  AOI21_X1 U4901 ( .B1(n3952), .B2(EAX_REG_27__SCAN_IN), .A(n3946), .ZN(n3947)
         );
  OAI21_X1 U4902 ( .B1(n3948), .B2(n3996), .A(n3947), .ZN(n3949) );
  XNOR2_X1 U4903 ( .A(n3970), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5132)
         );
  INV_X1 U4904 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5119) );
  NOR2_X1 U4905 ( .A1(n5119), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3951) );
  AOI211_X1 U4906 ( .C1(n3952), .C2(EAX_REG_28__SCAN_IN), .A(n3969), .B(n3951), 
        .ZN(n3968) );
  NAND2_X1 U4907 ( .A1(n3954), .A2(n3953), .ZN(n3976) );
  AOI22_X1 U4908 ( .A1(n3984), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3985), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4909 ( .A1(n4001), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4910 ( .A1(n4007), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4911 ( .A1(n4009), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3955) );
  NAND4_X1 U4912 ( .A1(n3958), .A2(n3957), .A3(n3956), .A4(n3955), .ZN(n3965)
         );
  AOI22_X1 U4913 ( .A1(n4011), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3999), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4914 ( .A1(n4013), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4915 ( .A1(n4000), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3959), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4916 ( .A1(n3348), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3960) );
  NAND4_X1 U4917 ( .A1(n3963), .A2(n3962), .A3(n3961), .A4(n3960), .ZN(n3964)
         );
  NOR2_X1 U4918 ( .A1(n3965), .A2(n3964), .ZN(n3977) );
  XOR2_X1 U4919 ( .A(n3976), .B(n3977), .Z(n3966) );
  NAND2_X1 U4920 ( .A1(n3966), .A2(n4028), .ZN(n3967) );
  AOI22_X1 U4921 ( .A1(n5132), .A2(n3969), .B1(n3968), .B2(n3967), .ZN(n5120)
         );
  INV_X1 U4922 ( .A(n3970), .ZN(n3971) );
  INV_X1 U4923 ( .A(n3972), .ZN(n3974) );
  INV_X1 U4924 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3973) );
  NAND2_X1 U4925 ( .A1(n3974), .A2(n3973), .ZN(n3975) );
  NAND2_X1 U4926 ( .A1(n4345), .A2(n3975), .ZN(n5430) );
  NOR2_X1 U4927 ( .A1(n3977), .A2(n3976), .ZN(n4021) );
  NOR2_X1 U4928 ( .A1(n3979), .A2(n3978), .ZN(n3983) );
  INV_X1 U4929 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3981) );
  INV_X1 U4930 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3980) );
  OAI22_X1 U4931 ( .A1(n3390), .A2(n3981), .B1(n3361), .B2(n3980), .ZN(n3982)
         );
  AOI211_X1 U4932 ( .C1(INSTQUEUE_REG_5__6__SCAN_IN), .C2(n3999), .A(n3983), 
        .B(n3982), .ZN(n3993) );
  AOI22_X1 U4933 ( .A1(n3984), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4007), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U4934 ( .A1(n3985), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4935 ( .A1(n4009), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U4936 ( .A1(n4001), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U4937 ( .A1(n3348), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U4938 ( .A1(n4013), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3986) );
  AND4_X1 U4939 ( .A1(n3989), .A2(n3988), .A3(n3987), .A4(n3986), .ZN(n3990)
         );
  NAND4_X1 U4940 ( .A1(n3993), .A2(n3992), .A3(n3991), .A4(n3990), .ZN(n4020)
         );
  XNOR2_X1 U4941 ( .A(n4021), .B(n4020), .ZN(n3997) );
  AOI21_X1 U4942 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6583), .A(n4031), 
        .ZN(n3995) );
  NAND2_X1 U4943 ( .A1(n3952), .A2(EAX_REG_29__SCAN_IN), .ZN(n3994) );
  OAI211_X1 U4944 ( .C1(n3997), .C2(n3996), .A(n3995), .B(n3994), .ZN(n3998)
         );
  OAI21_X1 U4945 ( .B1(n5430), .B2(n4025), .A(n3998), .ZN(n4344) );
  XNOR2_X1 U4946 ( .A(n4345), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5222)
         );
  AOI22_X1 U4947 ( .A1(n4000), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3999), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4948 ( .A1(n4001), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3938), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U4949 ( .A1(n3985), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4950 ( .A1(n3348), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4002), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4003) );
  NAND4_X1 U4951 ( .A1(n4006), .A2(n4005), .A3(n4004), .A4(n4003), .ZN(n4019)
         );
  AOI22_X1 U4952 ( .A1(n3984), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4007), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4953 ( .A1(n4009), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4008), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U4954 ( .A1(n4011), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4010), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U4955 ( .A1(n4013), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4014) );
  NAND4_X1 U4956 ( .A1(n4017), .A2(n4016), .A3(n4015), .A4(n4014), .ZN(n4018)
         );
  NOR2_X1 U4957 ( .A1(n4019), .A2(n4018), .ZN(n4023) );
  NAND2_X1 U4958 ( .A1(n4021), .A2(n4020), .ZN(n4022) );
  XOR2_X1 U4959 ( .A(n4023), .B(n4022), .Z(n4029) );
  INV_X1 U4960 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4462) );
  NAND2_X1 U4961 ( .A1(n6583), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4024)
         );
  OAI211_X1 U4962 ( .C1(n4026), .C2(n4462), .A(n4025), .B(n4024), .ZN(n4027)
         );
  AOI21_X1 U4963 ( .B1(n4029), .B2(n4028), .A(n4027), .ZN(n4030) );
  AOI21_X1 U4964 ( .B1(n5222), .B2(n4031), .A(n4030), .ZN(n5148) );
  OAI21_X1 U4965 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6451), .A(n4043), 
        .ZN(n4035) );
  INV_X1 U4966 ( .A(n4035), .ZN(n4033) );
  NAND2_X1 U4967 ( .A1(n4073), .A2(n4033), .ZN(n4038) );
  XNOR2_X1 U4968 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4045) );
  XNOR2_X1 U4969 ( .A(n4045), .B(n4043), .ZN(n4286) );
  NAND2_X1 U4970 ( .A1(n4286), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4039) );
  AOI21_X1 U4971 ( .B1(n4073), .B2(n4510), .A(n3403), .ZN(n4040) );
  OAI21_X1 U4972 ( .B1(n4307), .B2(n4035), .A(n4034), .ZN(n4037) );
  AND2_X1 U4973 ( .A1(n3407), .A2(n5139), .ZN(n4036) );
  AOI222_X1 U4974 ( .A1(n4038), .A2(n4075), .B1(n4039), .B2(n4040), .C1(n4037), 
        .C2(n4060), .ZN(n4042) );
  AOI22_X1 U4975 ( .A1(n4040), .A2(n4286), .B1(n4075), .B2(n4039), .ZN(n4041)
         );
  NOR2_X1 U4976 ( .A1(n4042), .A2(n4041), .ZN(n4061) );
  INV_X1 U4977 ( .A(n4061), .ZN(n4065) );
  INV_X1 U4978 ( .A(n4043), .ZN(n4044) );
  NAND2_X1 U4979 ( .A1(n4045), .A2(n4044), .ZN(n4047) );
  NAND2_X1 U4980 ( .A1(n6456), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4046) );
  NAND2_X1 U4981 ( .A1(n4047), .A2(n4046), .ZN(n4051) );
  XNOR2_X1 U4982 ( .A(n4048), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4050)
         );
  XNOR2_X1 U4983 ( .A(n4051), .B(n4050), .ZN(n4285) );
  OAI21_X1 U4984 ( .B1(n4049), .B2(n4285), .A(n4060), .ZN(n4064) );
  INV_X1 U4985 ( .A(n4050), .ZN(n4052) );
  NAND2_X1 U4986 ( .A1(n4052), .A2(n4051), .ZN(n4054) );
  NAND2_X1 U4987 ( .A1(n6334), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4053) );
  NAND2_X1 U4988 ( .A1(n4054), .A2(n4053), .ZN(n4056) );
  XNOR2_X1 U4989 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4055) );
  NOR2_X1 U4990 ( .A1(n4056), .A2(n4055), .ZN(n4057) );
  NOR2_X1 U4991 ( .A1(n4066), .A2(n4057), .ZN(n4284) );
  NOR2_X1 U4992 ( .A1(n4260), .A2(n4284), .ZN(n4063) );
  INV_X1 U4993 ( .A(n4073), .ZN(n4059) );
  INV_X1 U4994 ( .A(n4285), .ZN(n4058) );
  AOI211_X1 U4995 ( .C1(n4061), .C2(n4060), .A(n4059), .B(n4058), .ZN(n4062)
         );
  AOI211_X1 U4996 ( .C1(n4065), .C2(n4064), .A(n4063), .B(n4062), .ZN(n4070)
         );
  AOI21_X1 U4997 ( .B1(n4287), .B2(n4284), .A(n4068), .ZN(n4069) );
  OAI22_X1 U4998 ( .A1(n4070), .A2(n4069), .B1(n4075), .B2(n4287), .ZN(n4071)
         );
  AOI222_X1 U4999 ( .A1(n4072), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B1(
        n4072), .B2(n5885), .C1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n5885), 
        .ZN(n4288) );
  NAND2_X1 U5000 ( .A1(n4288), .A2(n4073), .ZN(n4074) );
  NAND2_X1 U5001 ( .A1(n4077), .A2(n4074), .ZN(n4076) );
  NAND2_X1 U5002 ( .A1(n4080), .A2(n3296), .ZN(n4087) );
  INV_X1 U5003 ( .A(n3322), .ZN(n4082) );
  NAND2_X1 U5004 ( .A1(n4250), .A2(n3493), .ZN(n4093) );
  OAI211_X1 U5005 ( .C1(n4083), .C2(n4082), .A(n3099), .B(n4093), .ZN(n4302)
         );
  NOR2_X1 U5006 ( .A1(n5026), .A2(n4084), .ZN(n4514) );
  NAND2_X2 U5007 ( .A1(n4184), .A2(n4189), .ZN(n5204) );
  OAI21_X1 U5008 ( .B1(n4514), .B2(n5204), .A(n4213), .ZN(n4086) );
  OAI21_X1 U5009 ( .B1(n3404), .B2(n3099), .A(n4084), .ZN(n4085) );
  NAND2_X1 U5010 ( .A1(n4089), .A2(n4088), .ZN(n4529) );
  NAND2_X1 U5011 ( .A1(n5167), .A2(n4097), .ZN(n4550) );
  INV_X1 U5012 ( .A(n4524), .ZN(n4090) );
  NAND2_X1 U5013 ( .A1(n4090), .A2(n3324), .ZN(n4091) );
  OAI211_X1 U5014 ( .C1(n4525), .C2(n3331), .A(n4550), .B(n4091), .ZN(n4092)
         );
  AND2_X1 U5015 ( .A1(n5183), .A2(n6481), .ZN(n4094) );
  NAND2_X1 U5016 ( .A1(n5188), .A2(n4094), .ZN(n4099) );
  AND4_X1 U5017 ( .A1(n3250), .A2(n3403), .A3(n4095), .A4(n3331), .ZN(n4096)
         );
  NAND3_X1 U5018 ( .A1(n4199), .A2(n4097), .A3(n4096), .ZN(n4494) );
  INV_X1 U5019 ( .A(EBX_REG_1__SCAN_IN), .ZN(n6027) );
  NAND2_X1 U5020 ( .A1(n4181), .A2(n6027), .ZN(n4101) );
  NAND2_X1 U5021 ( .A1(n4081), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4100)
         );
  INV_X1 U5022 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4102) );
  OAI22_X1 U5023 ( .A1(n4184), .A2(n4102), .B1(n4081), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n4395) );
  NAND2_X1 U5024 ( .A1(n4436), .A2(n4373), .ZN(n6010) );
  INV_X1 U5025 ( .A(n4103), .ZN(n4104) );
  MUX2_X1 U5026 ( .A(n4180), .B(n4189), .S(EBX_REG_2__SCAN_IN), .Z(n4106) );
  OR2_X1 U5027 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4105)
         );
  NAND2_X1 U5028 ( .A1(n4106), .A2(n4105), .ZN(n4453) );
  MUX2_X1 U5029 ( .A(n4181), .B(n3296), .S(EBX_REG_4__SCAN_IN), .Z(n4108) );
  NOR2_X1 U5030 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4107)
         );
  NOR2_X1 U5031 ( .A1(n4108), .A2(n4107), .ZN(n4584) );
  NAND2_X1 U5032 ( .A1(n3296), .A2(n4373), .ZN(n4185) );
  MUX2_X1 U5033 ( .A(n4185), .B(n4184), .S(EBX_REG_3__SCAN_IN), .Z(n4112) );
  INV_X1 U5034 ( .A(n4184), .ZN(n4109) );
  NAND2_X1 U5035 ( .A1(n4109), .A2(n5203), .ZN(n4167) );
  NAND2_X1 U5036 ( .A1(n5203), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4110)
         );
  AND2_X1 U5037 ( .A1(n4167), .A2(n4110), .ZN(n4111) );
  NAND2_X1 U5038 ( .A1(n4112), .A2(n4111), .ZN(n4585) );
  NAND2_X1 U5039 ( .A1(n4584), .A2(n4585), .ZN(n4113) );
  INV_X1 U5040 ( .A(EBX_REG_5__SCAN_IN), .ZN(n6811) );
  MUX2_X1 U5041 ( .A(n4184), .B(n4185), .S(n6811), .Z(n4116) );
  NAND2_X1 U5042 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n5203), .ZN(n4114)
         );
  AND2_X1 U5043 ( .A1(n4167), .A2(n4114), .ZN(n4115) );
  NAND2_X1 U5044 ( .A1(n4116), .A2(n4115), .ZN(n4654) );
  MUX2_X1 U5045 ( .A(n4180), .B(n4189), .S(EBX_REG_6__SCAN_IN), .Z(n4117) );
  NAND2_X1 U5046 ( .A1(n3183), .A2(n4117), .ZN(n5955) );
  MUX2_X1 U5047 ( .A(n4185), .B(n4184), .S(EBX_REG_7__SCAN_IN), .Z(n4120) );
  NAND2_X1 U5048 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n5203), .ZN(n4118)
         );
  AND2_X1 U5049 ( .A1(n4167), .A2(n4118), .ZN(n4119) );
  MUX2_X1 U5050 ( .A(n4180), .B(n4189), .S(EBX_REG_8__SCAN_IN), .Z(n4121) );
  INV_X1 U5051 ( .A(n4121), .ZN(n4123) );
  NOR2_X1 U5052 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4122)
         );
  NOR2_X1 U5053 ( .A1(n4123), .A2(n4122), .ZN(n4734) );
  MUX2_X1 U5054 ( .A(n4185), .B(n4184), .S(EBX_REG_9__SCAN_IN), .Z(n4126) );
  NAND2_X1 U5055 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n5203), .ZN(n4124)
         );
  AND2_X1 U5056 ( .A1(n4167), .A2(n4124), .ZN(n4125) );
  NAND2_X1 U5057 ( .A1(n4126), .A2(n4125), .ZN(n5034) );
  NAND2_X1 U5058 ( .A1(n5035), .A2(n5034), .ZN(n5037) );
  MUX2_X1 U5059 ( .A(n4180), .B(n4189), .S(EBX_REG_10__SCAN_IN), .Z(n4127) );
  NAND2_X1 U5060 ( .A1(n3191), .A2(n4127), .ZN(n4866) );
  MUX2_X1 U5061 ( .A(n4185), .B(n4184), .S(EBX_REG_11__SCAN_IN), .Z(n4130) );
  NAND2_X1 U5062 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n5203), .ZN(n4128) );
  AND2_X1 U5063 ( .A1(n4167), .A2(n4128), .ZN(n4129) );
  NAND2_X1 U5064 ( .A1(n4189), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4131) );
  OAI211_X1 U5065 ( .C1(n5203), .C2(EBX_REG_12__SCAN_IN), .A(n4184), .B(n4131), 
        .ZN(n4132) );
  OAI21_X1 U5066 ( .B1(n4180), .B2(EBX_REG_12__SCAN_IN), .A(n4132), .ZN(n5701)
         );
  MUX2_X1 U5067 ( .A(n4181), .B(n3296), .S(EBX_REG_14__SCAN_IN), .Z(n4134) );
  NOR2_X1 U5068 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4133)
         );
  NOR2_X1 U5069 ( .A1(n4134), .A2(n4133), .ZN(n5291) );
  INV_X1 U5070 ( .A(n4185), .ZN(n4172) );
  INV_X1 U5071 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U5072 ( .A1(n4172), .A2(n6014), .ZN(n4138) );
  INV_X1 U5073 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4317) );
  NAND2_X1 U5074 ( .A1(n4184), .A2(n4317), .ZN(n4136) );
  NAND2_X1 U5075 ( .A1(n4373), .A2(n6014), .ZN(n4135) );
  NAND3_X1 U5076 ( .A1(n4136), .A2(n4189), .A3(n4135), .ZN(n4137) );
  NAND2_X1 U5077 ( .A1(n4138), .A2(n4137), .ZN(n5691) );
  AND2_X1 U5078 ( .A1(n5291), .A2(n5691), .ZN(n4139) );
  MUX2_X1 U5079 ( .A(n4181), .B(n3296), .S(EBX_REG_16__SCAN_IN), .Z(n4141) );
  NOR2_X1 U5080 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4140)
         );
  NOR2_X1 U5081 ( .A1(n4141), .A2(n4140), .ZN(n5264) );
  INV_X1 U5082 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U5083 ( .A1(n4172), .A2(n5367), .ZN(n4145) );
  INV_X1 U5084 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4318) );
  NAND2_X1 U5085 ( .A1(n4184), .A2(n4318), .ZN(n4143) );
  NAND2_X1 U5086 ( .A1(n4373), .A2(n5367), .ZN(n4142) );
  NAND3_X1 U5087 ( .A1(n4143), .A2(n4189), .A3(n4142), .ZN(n4144) );
  NAND2_X1 U5088 ( .A1(n4145), .A2(n4144), .ZN(n5278) );
  NAND2_X1 U5089 ( .A1(n5264), .A2(n5278), .ZN(n4146) );
  MUX2_X1 U5090 ( .A(n4185), .B(n4184), .S(EBX_REG_17__SCAN_IN), .Z(n4149) );
  NAND2_X1 U5091 ( .A1(n5203), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4147) );
  AND2_X1 U5092 ( .A1(n4167), .A2(n4147), .ZN(n4148) );
  INV_X1 U5093 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U5094 ( .A1(n4181), .A2(n5859), .ZN(n4153) );
  NAND2_X1 U5095 ( .A1(n4373), .A2(n5859), .ZN(n4151) );
  NAND2_X1 U5096 ( .A1(n4189), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4150) );
  NAND3_X1 U5097 ( .A1(n4151), .A2(n4184), .A3(n4150), .ZN(n4152) );
  NAND2_X1 U5098 ( .A1(n5204), .A2(EBX_REG_18__SCAN_IN), .ZN(n4155) );
  NAND2_X1 U5099 ( .A1(n5203), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4154) );
  NAND2_X1 U5100 ( .A1(n4155), .A2(n4154), .ZN(n5346) );
  AND2_X1 U5101 ( .A1(n5346), .A2(n4189), .ZN(n5250) );
  NOR2_X1 U5102 ( .A1(n5346), .A2(n4189), .ZN(n5251) );
  OR2_X1 U5103 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4158)
         );
  INV_X1 U5104 ( .A(EBX_REG_20__SCAN_IN), .ZN(n4156) );
  NAND2_X1 U5105 ( .A1(n4373), .A2(n4156), .ZN(n4157) );
  NAND2_X1 U5106 ( .A1(n4158), .A2(n4157), .ZN(n5349) );
  MUX2_X1 U5107 ( .A(n5250), .B(n5251), .S(n5349), .Z(n4159) );
  MUX2_X1 U5108 ( .A(n4181), .B(n3296), .S(EBX_REG_22__SCAN_IN), .Z(n4161) );
  NOR2_X1 U5109 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4160)
         );
  NOR2_X1 U5110 ( .A1(n4161), .A2(n4160), .ZN(n5241) );
  MUX2_X1 U5111 ( .A(n4185), .B(n4184), .S(EBX_REG_21__SCAN_IN), .Z(n4164) );
  NAND2_X1 U5112 ( .A1(n5203), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4162) );
  AND2_X1 U5113 ( .A1(n4167), .A2(n4162), .ZN(n4163) );
  NAND2_X1 U5114 ( .A1(n4164), .A2(n4163), .ZN(n5340) );
  NAND2_X1 U5115 ( .A1(n5241), .A2(n5340), .ZN(n4165) );
  MUX2_X1 U5116 ( .A(n4185), .B(n4184), .S(EBX_REG_23__SCAN_IN), .Z(n4169) );
  NAND2_X1 U5117 ( .A1(n5203), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4166) );
  AND2_X1 U5118 ( .A1(n4167), .A2(n4166), .ZN(n4168) );
  NAND2_X1 U5119 ( .A1(n4169), .A2(n4168), .ZN(n5331) );
  NAND2_X1 U5120 ( .A1(n5332), .A2(n5331), .ZN(n5334) );
  NAND2_X1 U5121 ( .A1(n4189), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4170) );
  OAI211_X1 U5122 ( .C1(n5203), .C2(EBX_REG_24__SCAN_IN), .A(n4184), .B(n4170), 
        .ZN(n4171) );
  OAI21_X1 U5123 ( .B1(n4180), .B2(EBX_REG_24__SCAN_IN), .A(n4171), .ZN(n5068)
         );
  INV_X1 U5124 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U5125 ( .A1(n4172), .A2(n5324), .ZN(n4176) );
  INV_X1 U5126 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6731) );
  NAND2_X1 U5127 ( .A1(n4184), .A2(n6731), .ZN(n4174) );
  NAND2_X1 U5128 ( .A1(n4373), .A2(n5324), .ZN(n4173) );
  NAND3_X1 U5129 ( .A1(n4174), .A2(n4189), .A3(n4173), .ZN(n4175) );
  AND2_X1 U5130 ( .A1(n4176), .A2(n4175), .ZN(n5320) );
  INV_X1 U5131 ( .A(n5320), .ZN(n4177) );
  NAND2_X1 U5132 ( .A1(n4189), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4178) );
  OAI211_X1 U5133 ( .C1(n5203), .C2(EBX_REG_26__SCAN_IN), .A(n4184), .B(n4178), 
        .ZN(n4179) );
  OAI21_X1 U5134 ( .B1(n4180), .B2(EBX_REG_26__SCAN_IN), .A(n4179), .ZN(n5229)
         );
  MUX2_X1 U5135 ( .A(n4181), .B(n3296), .S(EBX_REG_28__SCAN_IN), .Z(n4183) );
  NOR2_X1 U5136 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4182)
         );
  NOR2_X1 U5137 ( .A1(n4183), .A2(n4182), .ZN(n5126) );
  MUX2_X1 U5138 ( .A(n4185), .B(n4184), .S(EBX_REG_27__SCAN_IN), .Z(n4187) );
  NAND2_X1 U5139 ( .A1(n5203), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4186) );
  NAND2_X1 U5140 ( .A1(n4187), .A2(n4186), .ZN(n5311) );
  NAND2_X1 U5141 ( .A1(n5126), .A2(n5311), .ZN(n4188) );
  OR2_X1 U5142 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4191)
         );
  INV_X1 U5143 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5162) );
  NAND2_X1 U5144 ( .A1(n4373), .A2(n5162), .ZN(n4190) );
  NAND2_X1 U5145 ( .A1(n4191), .A2(n4190), .ZN(n4367) );
  AND2_X1 U5146 ( .A1(n5128), .A2(n4367), .ZN(n4192) );
  INV_X1 U5147 ( .A(n5204), .ZN(n4194) );
  INV_X1 U5148 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5219) );
  INV_X1 U5149 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4340) );
  OAI22_X1 U5150 ( .A1(n4194), .A2(n5219), .B1(n4373), .B2(n4340), .ZN(n5201)
         );
  INV_X1 U5151 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U5152 ( .A1(n4219), .A2(n4212), .ZN(n4211) );
  INV_X1 U5153 ( .A(n4206), .ZN(n4201) );
  NAND2_X1 U5154 ( .A1(n4211), .A2(n4201), .ZN(n4233) );
  XNOR2_X1 U5155 ( .A(n4233), .B(n4232), .ZN(n4203) );
  INV_X1 U5156 ( .A(n4202), .ZN(n4258) );
  OR2_X1 U5157 ( .A1(n4203), .A2(n4258), .ZN(n4204) );
  XNOR2_X1 U5158 ( .A(n4211), .B(n4206), .ZN(n4208) );
  NAND2_X1 U5159 ( .A1(n3324), .A2(n4207), .ZN(n4218) );
  OAI21_X1 U5160 ( .B1(n4208), .B2(n4258), .A(n4218), .ZN(n4209) );
  AOI21_X1 U5161 ( .B1(n4575), .B2(n4250), .A(n4209), .ZN(n6099) );
  NAND2_X1 U5162 ( .A1(n4210), .A2(n4250), .ZN(n4217) );
  OAI21_X1 U5163 ( .B1(n4212), .B2(n4219), .A(n4211), .ZN(n4214) );
  OAI211_X1 U5164 ( .C1(n4214), .C2(n4258), .A(n3095), .B(n5139), .ZN(n4215)
         );
  INV_X1 U5165 ( .A(n4215), .ZN(n4216) );
  NAND2_X1 U5166 ( .A1(n4217), .A2(n4216), .ZN(n4432) );
  NAND2_X1 U5167 ( .A1(n5728), .A2(n4250), .ZN(n4222) );
  OAI21_X1 U5168 ( .B1(n4258), .B2(n4219), .A(n4218), .ZN(n4220) );
  INV_X1 U5169 ( .A(n4220), .ZN(n4221) );
  NAND2_X1 U5170 ( .A1(n4399), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4223)
         );
  INV_X1 U5171 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U5172 ( .A1(n4223), .A2(n6180), .ZN(n4224) );
  AND2_X1 U5173 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U5174 ( .A1(n4399), .A2(n6177), .ZN(n4225) );
  AND2_X1 U5175 ( .A1(n4224), .A2(n4225), .ZN(n4431) );
  NAND2_X1 U5176 ( .A1(n4432), .A2(n4431), .ZN(n4226) );
  NAND2_X1 U5177 ( .A1(n6098), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4228)
         );
  INV_X1 U5178 ( .A(n6098), .ZN(n4227) );
  INV_X1 U5179 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U5180 ( .A1(n4843), .A2(n4842), .ZN(n4841) );
  INV_X1 U5181 ( .A(n4229), .ZN(n4230) );
  OR2_X1 U5182 ( .A1(n4230), .A2(n4205), .ZN(n4231) );
  NAND2_X1 U5183 ( .A1(n4841), .A2(n4231), .ZN(n6090) );
  NAND2_X1 U5184 ( .A1(n4233), .A2(n4232), .ZN(n4248) );
  XOR2_X1 U5185 ( .A(n4246), .B(n4248), .Z(n4234) );
  NAND2_X1 U5186 ( .A1(n6090), .A2(n6089), .ZN(n6088) );
  INV_X1 U5187 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U5188 ( .A1(n6088), .A2(n4237), .ZN(n4851) );
  INV_X1 U5189 ( .A(n4248), .ZN(n4238) );
  NAND2_X1 U5190 ( .A1(n4238), .A2(n4246), .ZN(n4239) );
  XOR2_X1 U5191 ( .A(n4245), .B(n4239), .Z(n4240) );
  OAI22_X1 U5192 ( .A1(n4241), .A2(n4260), .B1(n4240), .B2(n4258), .ZN(n4243)
         );
  INV_X1 U5193 ( .A(n4243), .ZN(n4242) );
  NAND2_X1 U5194 ( .A1(n4851), .A2(n4850), .ZN(n4849) );
  INV_X1 U5195 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U5196 ( .A1(n4849), .A2(n4244), .ZN(n6082) );
  NAND2_X1 U5197 ( .A1(n4246), .A2(n4245), .ZN(n4247) );
  NOR2_X1 U5198 ( .A1(n4248), .A2(n4247), .ZN(n4257) );
  XNOR2_X1 U5199 ( .A(n4257), .B(n4256), .ZN(n4253) );
  NAND3_X1 U5200 ( .A1(n4251), .A2(n4250), .A3(n4249), .ZN(n4252) );
  OAI21_X1 U5201 ( .B1(n4253), .B2(n4258), .A(n4252), .ZN(n4254) );
  XOR2_X1 U5202 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .B(n4254), .Z(n6081) );
  NAND2_X1 U5203 ( .A1(n6082), .A2(n6081), .ZN(n6080) );
  INV_X1 U5204 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U5205 ( .A1(n6080), .A2(n4255), .ZN(n4857) );
  NAND2_X1 U5206 ( .A1(n4257), .A2(n4256), .ZN(n4266) );
  XOR2_X1 U5207 ( .A(n4264), .B(n4266), .Z(n4259) );
  OAI22_X1 U5208 ( .A1(n4261), .A2(n4260), .B1(n4259), .B2(n4258), .ZN(n4262)
         );
  XOR2_X1 U5209 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .B(n4262), .Z(n4856) );
  INV_X1 U5210 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U5211 ( .A1(n4262), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4263)
         );
  NAND2_X1 U5212 ( .A1(n4855), .A2(n4263), .ZN(n4970) );
  NAND2_X1 U5213 ( .A1(n4202), .A2(n4264), .ZN(n4265) );
  OAI21_X1 U5214 ( .B1(n4266), .B2(n4265), .A(n5557), .ZN(n4267) );
  XOR2_X1 U5215 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .B(n4267), .Z(n4969) );
  NAND2_X1 U5216 ( .A1(n4970), .A2(n4969), .ZN(n4968) );
  INV_X1 U5217 ( .A(n4267), .ZN(n4268) );
  INV_X1 U5218 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6739) );
  INV_X1 U5219 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5094) );
  NAND2_X1 U5220 ( .A1(n5557), .A2(n5094), .ZN(n5082) );
  NOR2_X1 U5221 ( .A1(n5557), .A2(n5094), .ZN(n5084) );
  INV_X1 U5222 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4270) );
  INV_X1 U5223 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5706) );
  XNOR2_X1 U5224 ( .A(n5557), .B(n5706), .ZN(n5552) );
  XNOR2_X1 U5225 ( .A(n5557), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5545)
         );
  INV_X1 U5226 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6624) );
  NAND2_X1 U5227 ( .A1(n5557), .A2(n4318), .ZN(n5526) );
  NAND3_X1 U5228 ( .A1(n5665), .A2(n5500), .A3(n4271), .ZN(n4272) );
  OAI21_X1 U5229 ( .B1(n5501), .B2(n4272), .A(n5716), .ZN(n4275) );
  NAND2_X1 U5230 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5644) );
  INV_X1 U5231 ( .A(n5644), .ZN(n4273) );
  NAND2_X1 U5232 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U5233 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U5234 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4337) );
  NOR3_X1 U5235 ( .A1(n5630), .A2(n5646), .A3(n4337), .ZN(n4276) );
  NAND2_X1 U5236 ( .A1(n5492), .A2(n3181), .ZN(n4280) );
  INV_X1 U5237 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6871) );
  INV_X1 U5238 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4277) );
  NAND2_X1 U5239 ( .A1(n6871), .A2(n4277), .ZN(n5645) );
  INV_X1 U5240 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6760) );
  INV_X1 U5241 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4278) );
  NAND2_X1 U5242 ( .A1(n6760), .A2(n4278), .ZN(n5629) );
  XOR2_X1 U5243 ( .A(n5557), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .Z(n5454) );
  AND2_X1 U5244 ( .A1(n5557), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5442)
         );
  NAND2_X1 U5245 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4339) );
  NOR2_X1 U5246 ( .A1(n5557), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5443)
         );
  NOR2_X1 U5247 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4281) );
  NAND2_X1 U5248 ( .A1(n5443), .A2(n4281), .ZN(n5145) );
  AOI21_X1 U5249 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5425), .A(n5426), 
        .ZN(n4282) );
  XNOR2_X1 U5250 ( .A(n4282), .B(n4340), .ZN(n5059) );
  NAND2_X1 U5251 ( .A1(n4283), .A2(n6507), .ZN(n6503) );
  NAND2_X1 U5252 ( .A1(n4510), .A2(n6503), .ZN(n4290) );
  INV_X1 U5253 ( .A(READY_N), .ZN(n6506) );
  AND3_X1 U5254 ( .A1(n4286), .A2(n4285), .A3(n4284), .ZN(n4289) );
  OAI21_X1 U5255 ( .B1(n4289), .B2(n4288), .A(n4287), .ZN(n5189) );
  AND2_X1 U5256 ( .A1(n6506), .A2(n5189), .ZN(n4489) );
  NAND2_X1 U5257 ( .A1(n4290), .A2(n4489), .ZN(n4297) );
  INV_X1 U5258 ( .A(n5188), .ZN(n4295) );
  AND2_X1 U5259 ( .A1(n4292), .A2(n4291), .ZN(n4527) );
  INV_X1 U5260 ( .A(n6503), .ZN(n4509) );
  OR2_X1 U5261 ( .A1(n4510), .A2(n4509), .ZN(n4355) );
  NAND3_X1 U5262 ( .A1(n4527), .A2(n4355), .A3(n6506), .ZN(n4293) );
  NAND3_X1 U5263 ( .A1(n4293), .A2(n3099), .A3(n3404), .ZN(n4294) );
  NAND2_X1 U5264 ( .A1(n4295), .A2(n4294), .ZN(n4296) );
  MUX2_X1 U5265 ( .A(n4297), .B(n4296), .S(n4746), .Z(n4305) );
  INV_X1 U5266 ( .A(n3096), .ZN(n5180) );
  NAND2_X1 U5267 ( .A1(n4299), .A2(n3324), .ZN(n4300) );
  NAND2_X1 U5268 ( .A1(n4308), .A2(n4302), .ZN(n4303) );
  NAND2_X1 U5269 ( .A1(n5180), .A2(n4303), .ZN(n4516) );
  NAND3_X1 U5270 ( .A1(n5188), .A2(n5167), .A3(n4510), .ZN(n4304) );
  NAND3_X1 U5271 ( .A1(n4305), .A2(n4516), .A3(n4304), .ZN(n4306) );
  NAND2_X1 U5272 ( .A1(n4308), .A2(n5023), .ZN(n4532) );
  NAND2_X1 U5273 ( .A1(n4308), .A2(n4307), .ZN(n4421) );
  AND2_X1 U5274 ( .A1(n4532), .A2(n4421), .ZN(n5179) );
  AOI22_X1 U5275 ( .A1(n4373), .A2(n4527), .B1(n4326), .B2(n3376), .ZN(n4310)
         );
  NAND3_X1 U5276 ( .A1(n5179), .A2(n4310), .A3(n4309), .ZN(n4311) );
  AND2_X1 U5277 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5566) );
  INV_X1 U5278 ( .A(n5566), .ZN(n4325) );
  NAND2_X1 U5279 ( .A1(n4329), .A2(n4312), .ZN(n5872) );
  NAND2_X1 U5280 ( .A1(n5641), .A2(n5872), .ZN(n5688) );
  INV_X1 U5281 ( .A(n5688), .ZN(n4313) );
  INV_X1 U5282 ( .A(n4339), .ZN(n4324) );
  INV_X1 U5283 ( .A(n6137), .ZN(n5679) );
  INV_X1 U5284 ( .A(n4329), .ZN(n4314) );
  NAND2_X1 U5285 ( .A1(n4314), .A2(n6190), .ZN(n4435) );
  OAI21_X1 U5286 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n5872), .A(n4435), 
        .ZN(n5090) );
  INV_X1 U5287 ( .A(n5090), .ZN(n6134) );
  AOI21_X1 U5288 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6175) );
  NAND2_X1 U5289 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6159) );
  NOR2_X1 U5290 ( .A1(n6175), .A2(n6159), .ZN(n6148) );
  NAND2_X1 U5291 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6148), .ZN(n6138)
         );
  NOR2_X1 U5292 ( .A1(n6144), .A2(n6138), .ZN(n5088) );
  NOR2_X1 U5293 ( .A1(n6132), .A2(n6739), .ZN(n6120) );
  INV_X1 U5294 ( .A(n6120), .ZN(n5093) );
  NAND2_X1 U5295 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6113) );
  NOR2_X1 U5296 ( .A1(n5093), .A2(n6113), .ZN(n4315) );
  NAND2_X1 U5297 ( .A1(n5088), .A2(n4315), .ZN(n4333) );
  NAND2_X1 U5298 ( .A1(n5690), .A2(n5872), .ZN(n5086) );
  NAND4_X1 U5299 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6146) );
  NOR3_X1 U5300 ( .A1(n6145), .A2(n6144), .A3(n6146), .ZN(n5087) );
  NAND2_X1 U5301 ( .A1(n4315), .A2(n5087), .ZN(n4332) );
  AOI22_X1 U5302 ( .A1(n4333), .A2(n6178), .B1(n5086), .B2(n4332), .ZN(n4316)
         );
  NAND2_X1 U5303 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5704) );
  NOR2_X1 U5304 ( .A1(n4317), .A2(n5704), .ZN(n5876) );
  NAND2_X1 U5305 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5876), .ZN(n5680) );
  NOR2_X1 U5306 ( .A1(n4318), .A2(n5680), .ZN(n5864) );
  NAND2_X1 U5307 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n5864), .ZN(n4334) );
  NAND2_X1 U5308 ( .A1(n6137), .A2(n4334), .ZN(n4319) );
  NAND2_X1 U5309 ( .A1(n5703), .A2(n4319), .ZN(n5670) );
  INV_X1 U5310 ( .A(n5646), .ZN(n5460) );
  NAND2_X1 U5311 ( .A1(n5460), .A2(n4273), .ZN(n4336) );
  AND2_X1 U5312 ( .A1(n6137), .A2(n4336), .ZN(n4320) );
  AND2_X1 U5313 ( .A1(n6137), .A2(n5630), .ZN(n4321) );
  NOR2_X1 U5314 ( .A1(n5636), .A2(n4321), .ZN(n5621) );
  INV_X1 U5315 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5109) );
  NAND2_X1 U5316 ( .A1(n5109), .A2(n5690), .ZN(n4433) );
  NAND2_X1 U5317 ( .A1(n4433), .A2(n5086), .ZN(n6179) );
  NAND2_X1 U5318 ( .A1(n5641), .A2(n6179), .ZN(n5092) );
  NAND2_X1 U5319 ( .A1(n5092), .A2(n4337), .ZN(n4322) );
  NAND2_X1 U5320 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U5321 ( .A1(n6137), .A2(n5603), .ZN(n4323) );
  OAI21_X1 U5322 ( .B1(n4324), .B2(n5679), .A(n5584), .ZN(n5578) );
  AOI21_X1 U5323 ( .B1(n4325), .B2(n6137), .A(n5578), .ZN(n5569) );
  INV_X1 U5324 ( .A(n5569), .ZN(n4331) );
  NAND2_X1 U5325 ( .A1(n4527), .A2(n4202), .ZN(n6474) );
  NAND2_X1 U5326 ( .A1(n4326), .A2(n3377), .ZN(n4327) );
  NAND2_X1 U5327 ( .A1(n6474), .A2(n4327), .ZN(n4328) );
  NAND2_X1 U5328 ( .A1(n6156), .A2(REIP_REG_30__SCAN_IN), .ZN(n5055) );
  OAI21_X1 U5329 ( .B1(n5220), .B2(n6127), .A(n5055), .ZN(n4330) );
  AOI21_X1 U5330 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n4331), .A(n4330), 
        .ZN(n4342) );
  INV_X1 U5331 ( .A(n4334), .ZN(n4335) );
  INV_X1 U5332 ( .A(n5630), .ZN(n5461) );
  INV_X1 U5333 ( .A(n4337), .ZN(n4338) );
  NAND2_X1 U5334 ( .A1(n5623), .A2(n4338), .ZN(n5612) );
  NOR2_X1 U5335 ( .A1(n5598), .A2(n4339), .ZN(n5580) );
  NAND3_X1 U5336 ( .A1(n5580), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n4340), .ZN(n4341) );
  OAI21_X1 U5337 ( .B1(n5059), .B2(n6184), .A(n4343), .ZN(U2988) );
  AOI21_X1 U5338 ( .B1(n4344), .B2(n5122), .A(n5149), .ZN(n5432) );
  INV_X1 U5339 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6869) );
  INV_X1 U5340 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4346) );
  AND2_X1 U5341 ( .A1(n3096), .A2(n6481), .ZN(n4349) );
  NAND2_X1 U5342 ( .A1(n5189), .A2(n4349), .ZN(n4390) );
  NAND2_X1 U5343 ( .A1(n6586), .A2(n6583), .ZN(n6492) );
  NOR3_X1 U5344 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6858), .A3(n6492), .ZN(
        n6487) );
  NOR2_X1 U5345 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6495) );
  INV_X1 U5346 ( .A(n6495), .ZN(n6585) );
  NOR3_X1 U5347 ( .A1(n6586), .A2(n6688), .A3(n6585), .ZN(n6479) );
  INV_X1 U5348 ( .A(n6479), .ZN(n4350) );
  NAND2_X1 U5349 ( .A1(n6190), .A2(n4350), .ZN(n4351) );
  NOR2_X1 U5350 ( .A1(n6487), .A2(n4351), .ZN(n4352) );
  NAND2_X1 U5351 ( .A1(n5044), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4378) );
  INV_X1 U5352 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6541) );
  INV_X1 U5353 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U5354 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5848) );
  NAND2_X1 U5355 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n5268) );
  NOR2_X1 U5356 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4371) );
  INV_X1 U5357 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6657) );
  NAND4_X1 U5358 ( .A1(REIP_REG_4__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .A4(REIP_REG_1__SCAN_IN), .ZN(n4816) );
  NOR2_X1 U5359 ( .A1(n6657), .A2(n4816), .ZN(n4814) );
  NAND4_X1 U5360 ( .A1(n4814), .A2(REIP_REG_8__SCAN_IN), .A3(
        REIP_REG_7__SCAN_IN), .A4(REIP_REG_6__SCAN_IN), .ZN(n5919) );
  NAND3_X1 U5361 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .ZN(n5920) );
  NOR2_X1 U5362 ( .A1(n5919), .A2(n5920), .ZN(n4356) );
  NAND4_X1 U5363 ( .A1(REIP_REG_12__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_14__SCAN_IN), .A4(n4356), .ZN(n4358) );
  NAND2_X1 U5364 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5907), .ZN(n5850) );
  NAND2_X1 U5365 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5839), .ZN(n5827) );
  NOR2_X1 U5366 ( .A1(n6539), .A2(n5827), .ZN(n5240) );
  NAND2_X1 U5367 ( .A1(REIP_REG_22__SCAN_IN), .A2(n5240), .ZN(n5825) );
  AND3_X1 U5368 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4363) );
  NAND2_X1 U5369 ( .A1(n5805), .A2(n4363), .ZN(n5798) );
  INV_X1 U5370 ( .A(REIP_REG_29__SCAN_IN), .ZN(n5428) );
  AND2_X1 U5371 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5210) );
  NAND2_X1 U5372 ( .A1(n5428), .A2(n5210), .ZN(n4357) );
  OR2_X1 U5373 ( .A1(n5798), .A2(n4357), .ZN(n5198) );
  NOR2_X1 U5374 ( .A1(n5998), .A2(n4358), .ZN(n5269) );
  NAND4_X1 U5375 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5269), .A3(
        REIP_REG_16__SCAN_IN), .A4(REIP_REG_15__SCAN_IN), .ZN(n5248) );
  NOR2_X1 U5376 ( .A1(n5248), .A2(n5848), .ZN(n4359) );
  NAND2_X1 U5377 ( .A1(n4359), .A2(REIP_REG_20__SCAN_IN), .ZN(n4360) );
  NAND2_X1 U5378 ( .A1(n5044), .A2(n5983), .ZN(n5921) );
  AND3_X1 U5379 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4361) );
  NOR2_X1 U5380 ( .A1(n5983), .A2(n4361), .ZN(n4362) );
  INV_X1 U5381 ( .A(n5983), .ZN(n5300) );
  INV_X1 U5382 ( .A(n4363), .ZN(n4364) );
  NAND2_X1 U5383 ( .A1(n5300), .A2(n4364), .ZN(n4365) );
  NAND2_X1 U5384 ( .A1(n5826), .A2(n4365), .ZN(n5792) );
  NOR2_X1 U5385 ( .A1(n5983), .A2(n5210), .ZN(n4366) );
  NOR2_X1 U5386 ( .A1(n5792), .A2(n4366), .ZN(n5197) );
  NAND2_X1 U5387 ( .A1(n4367), .A2(n4189), .ZN(n5200) );
  NAND2_X1 U5388 ( .A1(n3296), .A2(EBX_REG_29__SCAN_IN), .ZN(n4368) );
  AND2_X1 U5389 ( .A1(n5200), .A2(n4368), .ZN(n4369) );
  NAND2_X1 U5390 ( .A1(n5128), .A2(n4369), .ZN(n5202) );
  OR2_X1 U5391 ( .A1(n5128), .A2(n4369), .ZN(n4370) );
  NAND2_X1 U5392 ( .A1(n5202), .A2(n4370), .ZN(n5575) );
  AND2_X1 U5393 ( .A1(EBX_REG_31__SCAN_IN), .A2(n5024), .ZN(n5208) );
  INV_X1 U5394 ( .A(n4371), .ZN(n4374) );
  NAND2_X1 U5395 ( .A1(n5208), .A2(n4374), .ZN(n6009) );
  INV_X1 U5396 ( .A(n6009), .ZN(n4372) );
  OR2_X1 U5397 ( .A1(n6503), .A2(n4374), .ZN(n6473) );
  AND2_X1 U5398 ( .A1(n4202), .A2(n6473), .ZN(n5207) );
  INV_X1 U5399 ( .A(n5207), .ZN(n4376) );
  INV_X1 U5400 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5307) );
  NAND3_X1 U5401 ( .A1(n3099), .A2(n5307), .A3(n4374), .ZN(n4375) );
  NAND2_X1 U5402 ( .A1(n4376), .A2(n4375), .ZN(n4377) );
  AOI22_X1 U5403 ( .A1(n5990), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n5995), .ZN(n4382) );
  INV_X1 U5404 ( .A(n4378), .ZN(n4379) );
  INV_X1 U5405 ( .A(n5430), .ZN(n4380) );
  NAND2_X1 U5406 ( .A1(n6006), .A2(n4380), .ZN(n4381) );
  OAI211_X1 U5407 ( .C1(n5575), .C2(n5947), .A(n4382), .B(n4381), .ZN(n4383)
         );
  INV_X1 U5408 ( .A(n4383), .ZN(n4384) );
  NAND4_X1 U5409 ( .A1(n3108), .A2(n5198), .A3(n3194), .A4(n4384), .ZN(U2798)
         );
  NOR2_X2 U5410 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6380) );
  OAI21_X1 U5411 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n6393), .A(n4392), .ZN(
        n4387) );
  AOI21_X1 U5412 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n4390), .A(n4387), .ZN(
        n4385) );
  INV_X1 U5413 ( .A(n4385), .ZN(U2788) );
  OR2_X1 U5414 ( .A1(n4202), .A2(n4386), .ZN(n5194) );
  INV_X1 U5415 ( .A(n5194), .ZN(n4388) );
  OAI22_X1 U5416 ( .A1(n6588), .A2(n4388), .B1(n4387), .B2(
        READREQUEST_REG_SCAN_IN), .ZN(n4389) );
  OAI21_X1 U5417 ( .B1(n5194), .B2(n4390), .A(n4389), .ZN(U3474) );
  INV_X1 U5418 ( .A(DATAI_15_), .ZN(n4394) );
  INV_X1 U5419 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4393) );
  INV_X1 U5420 ( .A(n4392), .ZN(n4391) );
  OAI21_X2 U5421 ( .B1(n4202), .B2(n6506), .A(n4391), .ZN(n6061) );
  INV_X1 U5422 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6040) );
  OAI222_X1 U5423 ( .A1(n4394), .A2(n4493), .B1(n4393), .B2(n4464), .C1(n4458), 
        .C2(n6040), .ZN(U2954) );
  NOR2_X1 U5424 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4396)
         );
  OR2_X1 U5425 ( .A1(n4396), .A2(n4395), .ZN(n5028) );
  XNOR2_X1 U5426 ( .A(n4398), .B(n4397), .ZN(n5033) );
  OAI222_X1 U5427 ( .A1(n5028), .A2(n5376), .B1(n6026), .B2(n4102), .C1(n3092), 
        .C2(n5033), .ZN(U2859) );
  XNOR2_X1 U5428 ( .A(n4399), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4427)
         );
  INV_X1 U5429 ( .A(n5028), .ZN(n4402) );
  INV_X1 U5430 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6576) );
  NOR2_X1 U5431 ( .A1(n6190), .A2(n6576), .ZN(n4401) );
  AOI21_X1 U5432 ( .B1(n5690), .B2(n4435), .A(n5109), .ZN(n4400) );
  AOI211_X1 U5433 ( .C1(n4402), .C2(n6174), .A(n4401), .B(n4400), .ZN(n4403)
         );
  NAND2_X1 U5434 ( .A1(n5109), .A2(n5688), .ZN(n4434) );
  OAI211_X1 U5435 ( .C1(n4427), .C2(n6184), .A(n4403), .B(n4434), .ZN(U3018)
         );
  AOI22_X1 U5436 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n6061), .B1(n6069), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n4405) );
  INV_X1 U5437 ( .A(DATAI_5_), .ZN(n4404) );
  OR2_X1 U5438 ( .A1(n4493), .A2(n4404), .ZN(n4465) );
  NAND2_X1 U5439 ( .A1(n4405), .A2(n4465), .ZN(U2944) );
  AOI22_X1 U5440 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6061), .B1(n6069), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n4406) );
  INV_X1 U5441 ( .A(DATAI_6_), .ZN(n4612) );
  OR2_X1 U5442 ( .A1(n4493), .A2(n4612), .ZN(n4467) );
  NAND2_X1 U5443 ( .A1(n4406), .A2(n4467), .ZN(U2945) );
  AOI22_X1 U5444 ( .A1(UWORD_REG_0__SCAN_IN), .A2(n6070), .B1(n6069), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n4407) );
  INV_X1 U5445 ( .A(DATAI_0_), .ZN(n4503) );
  OR2_X1 U5446 ( .A1(n4493), .A2(n4503), .ZN(n4476) );
  NAND2_X1 U5447 ( .A1(n4407), .A2(n4476), .ZN(U2924) );
  AOI22_X1 U5448 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6061), .B1(n6069), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n4408) );
  INV_X1 U5449 ( .A(DATAI_7_), .ZN(n4616) );
  OR2_X1 U5450 ( .A1(n4493), .A2(n4616), .ZN(n4469) );
  NAND2_X1 U5451 ( .A1(n4408), .A2(n4469), .ZN(U2946) );
  AOI22_X1 U5452 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n6061), .B1(n6069), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n4409) );
  NAND2_X1 U5453 ( .A1(n6063), .A2(DATAI_4_), .ZN(n4481) );
  NAND2_X1 U5454 ( .A1(n4409), .A2(n4481), .ZN(U2943) );
  INV_X1 U5455 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6742) );
  NAND2_X1 U5456 ( .A1(n6063), .A2(DATAI_13_), .ZN(n6071) );
  NAND2_X1 U5457 ( .A1(n6070), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4410) );
  OAI211_X1 U5458 ( .C1(n6742), .C2(n4458), .A(n6071), .B(n4410), .ZN(U2937)
         );
  INV_X1 U5459 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6744) );
  NAND2_X1 U5460 ( .A1(n6070), .A2(LWORD_REG_9__SCAN_IN), .ZN(n4411) );
  NAND2_X1 U5461 ( .A1(n6063), .A2(DATAI_9_), .ZN(n4415) );
  OAI211_X1 U5462 ( .C1(n6744), .C2(n4458), .A(n4411), .B(n4415), .ZN(U2948)
         );
  INV_X1 U5463 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U5464 ( .A1(n6070), .A2(LWORD_REG_12__SCAN_IN), .ZN(n4412) );
  NAND2_X1 U5465 ( .A1(n6063), .A2(DATAI_12_), .ZN(n4413) );
  OAI211_X1 U5466 ( .C1(n6045), .C2(n4458), .A(n4412), .B(n4413), .ZN(U2951)
         );
  INV_X1 U5467 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4460) );
  NAND2_X1 U5468 ( .A1(n6070), .A2(UWORD_REG_12__SCAN_IN), .ZN(n4414) );
  OAI211_X1 U5469 ( .C1(n4460), .C2(n4458), .A(n4414), .B(n4413), .ZN(U2936)
         );
  INV_X1 U5470 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4605) );
  NAND2_X1 U5471 ( .A1(n6070), .A2(UWORD_REG_9__SCAN_IN), .ZN(n4416) );
  OAI211_X1 U5472 ( .C1(n4605), .C2(n4458), .A(n4416), .B(n4415), .ZN(U2933)
         );
  INV_X1 U5473 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6717) );
  NAND2_X1 U5474 ( .A1(n6070), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4417) );
  NAND2_X1 U5475 ( .A1(n6063), .A2(DATAI_8_), .ZN(n4418) );
  OAI211_X1 U5476 ( .C1(n6717), .C2(n4458), .A(n4417), .B(n4418), .ZN(U2947)
         );
  NAND2_X1 U5477 ( .A1(n6070), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4419) );
  OAI211_X1 U5478 ( .C1(n3881), .C2(n4458), .A(n4419), .B(n4418), .ZN(U2932)
         );
  NAND3_X1 U5479 ( .A1(n6586), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6493) );
  INV_X1 U5480 ( .A(n6493), .ZN(n4420) );
  AND2_X1 U5481 ( .A1(n6393), .A2(n4422), .ZN(n6589) );
  OR2_X1 U5482 ( .A1(n6589), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4423) );
  NAND2_X1 U5483 ( .A1(n6586), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4425) );
  NAND2_X1 U5484 ( .A1(n6584), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4424) );
  AND2_X1 U5485 ( .A1(n4425), .A2(n4424), .ZN(n4825) );
  INV_X1 U5486 ( .A(n4825), .ZN(n4426) );
  OAI21_X1 U5487 ( .B1(n6097), .B2(n4426), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4430) );
  INV_X1 U5488 ( .A(n4427), .ZN(n4428) );
  AOI22_X1 U5489 ( .A1(n6104), .A2(n4428), .B1(n6156), .B2(REIP_REG_0__SCAN_IN), .ZN(n4429) );
  OAI211_X1 U5490 ( .C1(n5033), .C2(n5564), .A(n4430), .B(n4429), .ZN(U2986)
         );
  XNOR2_X1 U5491 ( .A(n4432), .B(n4431), .ZN(n4829) );
  AND3_X1 U5492 ( .A1(n6137), .A2(n4433), .A3(n6180), .ZN(n4441) );
  AOI21_X1 U5493 ( .B1(n4435), .B2(n4434), .A(n6180), .ZN(n4440) );
  INV_X1 U5494 ( .A(n4436), .ZN(n4438) );
  INV_X1 U5495 ( .A(n6010), .ZN(n4437) );
  AOI21_X1 U5496 ( .B1(n4438), .B2(n5203), .A(n4437), .ZN(n6020) );
  INV_X1 U5497 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6570) );
  OAI22_X1 U5498 ( .A1(n6127), .A2(n6020), .B1(n6570), .B2(n6190), .ZN(n4439)
         );
  NOR3_X1 U5499 ( .A1(n4441), .A2(n4440), .A3(n4439), .ZN(n4442) );
  OAI21_X1 U5500 ( .B1(n4829), .B2(n6184), .A(n4442), .ZN(U3017) );
  NAND2_X1 U5501 ( .A1(n4444), .A2(n4443), .ZN(n4451) );
  XNOR2_X1 U5502 ( .A(n4445), .B(n4451), .ZN(n5050) );
  XNOR2_X1 U5503 ( .A(n4452), .B(n4585), .ZN(n6165) );
  INV_X1 U5504 ( .A(n6026), .ZN(n5368) );
  AOI22_X1 U5505 ( .A1(n6022), .A2(n6165), .B1(n5368), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4446) );
  OAI21_X1 U5506 ( .B1(n5050), .B2(n3092), .A(n4446), .ZN(U2856) );
  INV_X1 U5507 ( .A(n4447), .ZN(n4448) );
  OR3_X1 U5508 ( .A1(n4496), .A2(n4449), .A3(n4448), .ZN(n4450) );
  AND2_X1 U5509 ( .A1(n4451), .A2(n4450), .ZN(n6102) );
  INV_X1 U5510 ( .A(n6102), .ZN(n4505) );
  INV_X1 U5511 ( .A(n4452), .ZN(n4586) );
  AOI21_X1 U5512 ( .B1(n4454), .B2(n4453), .A(n4586), .ZN(n6173) );
  AOI22_X1 U5513 ( .A1(n6022), .A2(n6173), .B1(n5368), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4455) );
  OAI21_X1 U5514 ( .B1(n4505), .B2(n3092), .A(n4455), .ZN(U2857) );
  NAND2_X1 U5515 ( .A1(n4456), .A2(n6452), .ZN(n4457) );
  NAND2_X1 U5516 ( .A1(n4458), .A2(n4457), .ZN(n4459) );
  NAND2_X1 U5517 ( .A1(n6586), .A2(n5725), .ZN(n6590) );
  INV_X1 U5518 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n6662) );
  NAND2_X1 U5519 ( .A1(n6055), .A2(n3099), .ZN(n6033) );
  INV_X1 U5520 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n6613) );
  OAI222_X1 U5521 ( .A1(n6059), .A2(n6662), .B1(n6033), .B2(n4460), .C1(n6590), 
        .C2(n6613), .ZN(U2895) );
  INV_X1 U5522 ( .A(UWORD_REG_14__SCAN_IN), .ZN(n4463) );
  INV_X1 U5523 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4461) );
  OAI222_X1 U5524 ( .A1(n4463), .A2(n6590), .B1(n6033), .B2(n4462), .C1(n4461), 
        .C2(n6059), .ZN(U2893) );
  AOI22_X1 U5525 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n6061), .B1(n6069), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n4466) );
  NAND2_X1 U5526 ( .A1(n4466), .A2(n4465), .ZN(U2929) );
  AOI22_X1 U5527 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n6061), .B1(n6069), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n4468) );
  NAND2_X1 U5528 ( .A1(n4468), .A2(n4467), .ZN(U2930) );
  AOI22_X1 U5529 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n6061), .B1(n6069), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n4470) );
  NAND2_X1 U5530 ( .A1(n4470), .A2(n4469), .ZN(U2931) );
  AOI22_X1 U5531 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n6061), .B1(n6069), .B2(
        EAX_REG_3__SCAN_IN), .ZN(n4472) );
  INV_X1 U5532 ( .A(DATAI_3_), .ZN(n4471) );
  OR2_X1 U5533 ( .A1(n4493), .A2(n4471), .ZN(n4483) );
  NAND2_X1 U5534 ( .A1(n4472), .A2(n4483), .ZN(U2942) );
  AOI22_X1 U5535 ( .A1(LWORD_REG_14__SCAN_IN), .A2(n6061), .B1(n6069), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n4473) );
  NAND2_X1 U5536 ( .A1(n6063), .A2(DATAI_14_), .ZN(n4474) );
  NAND2_X1 U5537 ( .A1(n4473), .A2(n4474), .ZN(U2953) );
  AOI22_X1 U5538 ( .A1(UWORD_REG_14__SCAN_IN), .A2(n6061), .B1(n6069), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n4475) );
  NAND2_X1 U5539 ( .A1(n4475), .A2(n4474), .ZN(U2938) );
  AOI22_X1 U5540 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n6061), .B1(n6069), .B2(
        EAX_REG_0__SCAN_IN), .ZN(n4477) );
  NAND2_X1 U5541 ( .A1(n4477), .A2(n4476), .ZN(U2939) );
  AOI22_X1 U5542 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n6061), .B1(n6069), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n4479) );
  INV_X1 U5543 ( .A(DATAI_1_), .ZN(n4478) );
  OR2_X1 U5544 ( .A1(n4493), .A2(n4478), .ZN(n4485) );
  NAND2_X1 U5545 ( .A1(n4479), .A2(n4485), .ZN(U2940) );
  AOI22_X1 U5546 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n6061), .B1(n6069), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n4480) );
  NAND2_X1 U5547 ( .A1(n6063), .A2(DATAI_2_), .ZN(n4487) );
  NAND2_X1 U5548 ( .A1(n4480), .A2(n4487), .ZN(U2941) );
  AOI22_X1 U5549 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n6061), .B1(n6069), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n4482) );
  NAND2_X1 U5550 ( .A1(n4482), .A2(n4481), .ZN(U2928) );
  AOI22_X1 U5551 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n6061), .B1(n6069), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n4484) );
  NAND2_X1 U5552 ( .A1(n4484), .A2(n4483), .ZN(U2927) );
  AOI22_X1 U5553 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n6061), .B1(n6069), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n4486) );
  NAND2_X1 U5554 ( .A1(n4486), .A2(n4485), .ZN(U2925) );
  AOI22_X1 U5555 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n6061), .B1(n6069), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n4488) );
  NAND2_X1 U5556 ( .A1(n4488), .A2(n4487), .ZN(U2926) );
  OR2_X1 U5557 ( .A1(n5188), .A2(n4532), .ZN(n4491) );
  INV_X1 U5558 ( .A(n4309), .ZN(n5882) );
  NAND2_X1 U5559 ( .A1(n5882), .A2(n4489), .ZN(n4490) );
  NAND2_X1 U5560 ( .A1(n4520), .A2(n6481), .ZN(n4492) );
  INV_X1 U5561 ( .A(n5023), .ZN(n5187) );
  OR2_X1 U5562 ( .A1(n4494), .A2(n5187), .ZN(n4495) );
  NAND2_X1 U5563 ( .A1(n3322), .A2(n3472), .ZN(n4500) );
  INV_X1 U5564 ( .A(n4496), .ZN(n4497) );
  OAI21_X1 U5565 ( .B1(n4499), .B2(n4498), .A(n4497), .ZN(n6001) );
  INV_X1 U5566 ( .A(n4500), .ZN(n4501) );
  AOI22_X1 U5567 ( .A1(n6831), .A2(DATAI_1_), .B1(n6830), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n4502) );
  OAI21_X1 U5568 ( .B1(n5418), .B2(n6001), .A(n4502), .ZN(U2890) );
  INV_X1 U5569 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6696) );
  OAI222_X1 U5570 ( .A1(n5418), .A2(n5033), .B1(n5421), .B2(n4503), .C1(n5419), 
        .C2(n6696), .ZN(U2891) );
  AOI22_X1 U5571 ( .A1(n6831), .A2(DATAI_3_), .B1(n6830), .B2(
        EAX_REG_3__SCAN_IN), .ZN(n4504) );
  OAI21_X1 U5572 ( .B1(n5050), .B2(n5418), .A(n4504), .ZN(U2888) );
  INV_X1 U5573 ( .A(DATAI_2_), .ZN(n6674) );
  INV_X1 U5574 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6057) );
  OAI222_X1 U5575 ( .A1(n4505), .A2(n5418), .B1(n5421), .B2(n6674), .C1(n5419), 
        .C2(n6057), .ZN(U2889) );
  OAI21_X1 U5576 ( .B1(n3091), .B2(n4507), .A(n4506), .ZN(n6092) );
  INV_X1 U5577 ( .A(DATAI_4_), .ZN(n6756) );
  INV_X1 U5578 ( .A(EAX_REG_4__SCAN_IN), .ZN(n4508) );
  OAI222_X1 U5579 ( .A1(n6092), .A2(n5418), .B1(n5421), .B2(n6756), .C1(n4508), 
        .C2(n5419), .ZN(U2887) );
  OAI21_X1 U5580 ( .B1(n6452), .B2(n4527), .A(n4509), .ZN(n4512) );
  NAND2_X1 U5581 ( .A1(n4348), .A2(n4510), .ZN(n4511) );
  NAND2_X1 U5582 ( .A1(n4512), .A2(n4511), .ZN(n4513) );
  NAND2_X1 U5583 ( .A1(n4513), .A2(n6506), .ZN(n4519) );
  NAND2_X1 U5584 ( .A1(n5188), .A2(n5183), .ZN(n4518) );
  INV_X1 U5585 ( .A(n4514), .ZN(n4515) );
  AND2_X1 U5586 ( .A1(n4516), .A2(n4515), .ZN(n4517) );
  OAI211_X1 U5587 ( .C1(n5188), .C2(n4519), .A(n4518), .B(n4517), .ZN(n4521)
         );
  NAND2_X1 U5588 ( .A1(n4525), .A2(n4524), .ZN(n4526) );
  NOR2_X1 U5589 ( .A1(n4527), .A2(n4526), .ZN(n4528) );
  AND2_X1 U5590 ( .A1(n4309), .A2(n4528), .ZN(n4531) );
  INV_X1 U5591 ( .A(n4529), .ZN(n4530) );
  NAND2_X1 U5592 ( .A1(n4531), .A2(n4530), .ZN(n5171) );
  NAND2_X1 U5593 ( .A1(n4523), .A2(n5171), .ZN(n4540) );
  INV_X1 U5594 ( .A(n4532), .ZN(n4533) );
  OR2_X1 U5595 ( .A1(n5183), .A2(n4533), .ZN(n4548) );
  XNOR2_X1 U5596 ( .A(n4534), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4538)
         );
  XNOR2_X1 U5597 ( .A(n3195), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4535)
         );
  NAND2_X1 U5598 ( .A1(n6452), .A2(n4535), .ZN(n4536) );
  OAI21_X1 U5599 ( .B1(n4538), .B2(n4550), .A(n4536), .ZN(n4537) );
  AOI21_X1 U5600 ( .B1(n4548), .B2(n4538), .A(n4537), .ZN(n4539) );
  NAND2_X1 U5601 ( .A1(n4540), .A2(n4539), .ZN(n5113) );
  OR2_X1 U5602 ( .A1(n6449), .A2(n5113), .ZN(n4542) );
  NAND2_X1 U5603 ( .A1(n6449), .A2(n4048), .ZN(n4541) );
  NAND2_X1 U5604 ( .A1(n4542), .A2(n4541), .ZN(n6459) );
  INV_X1 U5605 ( .A(n6459), .ZN(n4559) );
  NAND2_X1 U5606 ( .A1(n6449), .A2(n3470), .ZN(n4558) );
  INV_X1 U5607 ( .A(n6449), .ZN(n4556) );
  NAND2_X1 U5608 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4544) );
  INV_X1 U5609 ( .A(n4544), .ZN(n4543) );
  MUX2_X1 U5610 ( .A(n4544), .B(n4543), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4554) );
  INV_X1 U5611 ( .A(n6452), .ZN(n4553) );
  MUX2_X1 U5612 ( .A(n4545), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4534), 
        .Z(n4546) );
  NOR2_X1 U5613 ( .A1(n4546), .A2(n4560), .ZN(n4547) );
  NAND2_X1 U5614 ( .A1(n4548), .A2(n4547), .ZN(n4552) );
  INV_X1 U5615 ( .A(n4545), .ZN(n4549) );
  OAI211_X1 U5616 ( .C1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n4534), .A(n3385), .B(n4549), .ZN(n6565) );
  OR2_X1 U5617 ( .A1(n4550), .A2(n6565), .ZN(n4551) );
  OAI211_X1 U5618 ( .C1(n4554), .C2(n4553), .A(n4552), .B(n4551), .ZN(n4555)
         );
  AOI21_X1 U5619 ( .B1(n3101), .B2(n5171), .A(n4555), .ZN(n6567) );
  NAND2_X1 U5620 ( .A1(n4556), .A2(n6567), .ZN(n4557) );
  NAND3_X1 U5621 ( .A1(n4559), .A2(n6462), .A3(n6858), .ZN(n4570) );
  INV_X1 U5622 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6753) );
  NAND2_X1 U5623 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6753), .ZN(n4566) );
  INV_X1 U5624 ( .A(n4560), .ZN(n4565) );
  INV_X1 U5625 ( .A(n4618), .ZN(n6263) );
  NOR2_X1 U5626 ( .A1(n4561), .A2(n6263), .ZN(n4562) );
  XNOR2_X1 U5627 ( .A(n4562), .B(n5885), .ZN(n5981) );
  NOR2_X1 U5628 ( .A1(n4309), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4563) );
  NAND2_X1 U5629 ( .A1(n5981), .A2(n4563), .ZN(n4564) );
  OAI21_X1 U5630 ( .B1(n4566), .B2(n4565), .A(n4564), .ZN(n4567) );
  INV_X1 U5631 ( .A(n4567), .ZN(n4569) );
  MUX2_X1 U5632 ( .A(n6449), .B(n6753), .S(STATE2_REG_1__SCAN_IN), .Z(n4568)
         );
  NAND2_X1 U5633 ( .A1(n4568), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4572) );
  NAND3_X1 U5634 ( .A1(n4570), .A2(n4569), .A3(n4572), .ZN(n6470) );
  NAND2_X1 U5635 ( .A1(n4571), .A2(n4572), .ZN(n4573) );
  NAND2_X1 U5636 ( .A1(n6470), .A2(n4573), .ZN(n5726) );
  NAND2_X1 U5637 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5725), .ZN(n6561) );
  AOI21_X1 U5638 ( .B1(n5726), .B2(n6753), .A(n6561), .ZN(n4574) );
  NAND2_X1 U5639 ( .A1(n4576), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4712) );
  XNOR2_X1 U5640 ( .A(n4713), .B(n4712), .ZN(n4577) );
  NAND2_X1 U5641 ( .A1(n6688), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5727) );
  AOI22_X1 U5642 ( .A1(n4577), .A2(n6380), .B1(n5727), .B2(n4523), .ZN(n4579)
         );
  NAND2_X1 U5643 ( .A1(n6191), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4578) );
  OAI21_X1 U5644 ( .B1(n6191), .B2(n4579), .A(n4578), .ZN(U3463) );
  AOI21_X1 U5645 ( .B1(n4769), .B2(n6584), .A(n6393), .ZN(n4581) );
  AOI22_X1 U5646 ( .A1(n4581), .A2(n4712), .B1(n4580), .B2(n5727), .ZN(n4583)
         );
  NAND2_X1 U5647 ( .A1(n6191), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4582) );
  OAI21_X1 U5648 ( .B1(n6191), .B2(n4583), .A(n4582), .ZN(U3464) );
  AOI21_X1 U5649 ( .B1(n4586), .B2(n4585), .A(n4584), .ZN(n4587) );
  OR2_X1 U5650 ( .A1(n4587), .A2(n3118), .ZN(n5978) );
  INV_X1 U5651 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4588) );
  OAI222_X1 U5652 ( .A1(n5978), .A2(n5376), .B1(n4588), .B2(n6026), .C1(n3092), 
        .C2(n6092), .ZN(U2855) );
  INV_X1 U5653 ( .A(n6191), .ZN(n4596) );
  NOR2_X1 U5654 ( .A1(n4576), .A2(n4589), .ZN(n4590) );
  NAND2_X1 U5655 ( .A1(n4713), .A2(n4590), .ZN(n4743) );
  INV_X1 U5656 ( .A(n4743), .ZN(n4636) );
  NAND2_X1 U5657 ( .A1(n4636), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4740) );
  INV_X1 U5658 ( .A(n4740), .ZN(n4591) );
  NOR2_X1 U5659 ( .A1(n4591), .A2(n6379), .ZN(n4715) );
  INV_X1 U5660 ( .A(n4712), .ZN(n6378) );
  NAND2_X1 U5661 ( .A1(n6257), .A2(n6378), .ZN(n6298) );
  AOI21_X1 U5662 ( .B1(n4715), .B2(n6298), .A(n6393), .ZN(n4594) );
  NAND2_X1 U5663 ( .A1(n6380), .A2(n6584), .ZN(n6265) );
  INV_X1 U5664 ( .A(n3101), .ZN(n5040) );
  INV_X1 U5665 ( .A(n5727), .ZN(n4592) );
  OAI22_X1 U5666 ( .A1(n4720), .A2(n6265), .B1(n5040), .B2(n4592), .ZN(n4593)
         );
  OAI21_X1 U5667 ( .B1(n4594), .B2(n4593), .A(n4596), .ZN(n4595) );
  OAI21_X1 U5668 ( .B1(n4596), .B2(n6460), .A(n4595), .ZN(U3462) );
  INV_X1 U5669 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6618) );
  AOI22_X1 U5670 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n6051), .B1(n6054), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4597) );
  OAI21_X1 U5671 ( .B1(n6618), .B2(n6033), .A(n4597), .ZN(U2904) );
  AOI22_X1 U5672 ( .A1(n6051), .A2(UWORD_REG_0__SCAN_IN), .B1(n6054), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4598) );
  OAI21_X1 U5673 ( .B1(n3729), .B2(n6033), .A(n4598), .ZN(U2907) );
  INV_X1 U5674 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6800) );
  AOI22_X1 U5675 ( .A1(n6051), .A2(UWORD_REG_6__SCAN_IN), .B1(n6054), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4599) );
  OAI21_X1 U5676 ( .B1(n6800), .B2(n6033), .A(n4599), .ZN(U2901) );
  AOI22_X1 U5677 ( .A1(n6051), .A2(UWORD_REG_8__SCAN_IN), .B1(n6054), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4600) );
  OAI21_X1 U5678 ( .B1(n3881), .B2(n6033), .A(n4600), .ZN(U2899) );
  AOI22_X1 U5679 ( .A1(n6051), .A2(UWORD_REG_7__SCAN_IN), .B1(n6054), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4601) );
  OAI21_X1 U5680 ( .B1(n3848), .B2(n6033), .A(n4601), .ZN(U2900) );
  INV_X1 U5681 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4603) );
  AOI22_X1 U5682 ( .A1(n6051), .A2(UWORD_REG_5__SCAN_IN), .B1(n6054), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4602) );
  OAI21_X1 U5683 ( .B1(n4603), .B2(n6033), .A(n4602), .ZN(U2902) );
  AOI22_X1 U5684 ( .A1(n6051), .A2(UWORD_REG_9__SCAN_IN), .B1(n6054), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4604) );
  OAI21_X1 U5685 ( .B1(n4605), .B2(n6033), .A(n4604), .ZN(U2898) );
  INV_X1 U5686 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6603) );
  AOI22_X1 U5687 ( .A1(n6051), .A2(UWORD_REG_1__SCAN_IN), .B1(n6054), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4606) );
  OAI21_X1 U5688 ( .B1(n6603), .B2(n6033), .A(n4606), .ZN(U2906) );
  AOI22_X1 U5689 ( .A1(n6051), .A2(UWORD_REG_13__SCAN_IN), .B1(n6054), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4607) );
  OAI21_X1 U5690 ( .B1(n6742), .B2(n6033), .A(n4607), .ZN(U2894) );
  NAND2_X1 U5691 ( .A1(n4610), .A2(n4609), .ZN(n4611) );
  AND2_X1 U5692 ( .A1(n4608), .A2(n4611), .ZN(n6084) );
  INV_X1 U5693 ( .A(n6084), .ZN(n4613) );
  OAI222_X1 U5694 ( .A1(n4613), .A2(n5418), .B1(n5421), .B2(n4612), .C1(n5419), 
        .C2(n3574), .ZN(U2885) );
  INV_X1 U5695 ( .A(n4614), .ZN(n4615) );
  XNOR2_X1 U5696 ( .A(n4608), .B(n4615), .ZN(n4861) );
  INV_X1 U5697 ( .A(n4861), .ZN(n4824) );
  OAI222_X1 U5698 ( .A1(n5418), .A2(n4824), .B1(n5421), .B2(n4616), .C1(n5419), 
        .C2(n3582), .ZN(U2884) );
  NAND2_X1 U5699 ( .A1(n6257), .A2(n4769), .ZN(n6227) );
  OR2_X1 U5700 ( .A1(n6227), .A2(n5728), .ZN(n6231) );
  AND2_X1 U5701 ( .A1(n6101), .A2(DATAI_19_), .ZN(n6415) );
  INV_X1 U5702 ( .A(n6415), .ZN(n6281) );
  OR2_X1 U5703 ( .A1(n6227), .A2(n6584), .ZN(n4617) );
  NAND2_X1 U5704 ( .A1(n4617), .A2(n6380), .ZN(n6230) );
  NAND3_X1 U5705 ( .A1(n4770), .A2(n5731), .A3(n4720), .ZN(n4881) );
  INV_X1 U5706 ( .A(n6265), .ZN(n6331) );
  INV_X1 U5707 ( .A(n4580), .ZN(n4716) );
  NAND2_X1 U5708 ( .A1(n4523), .A2(n4716), .ZN(n5733) );
  OR2_X1 U5709 ( .A1(n5733), .A2(n4618), .ZN(n6222) );
  OAI21_X1 U5710 ( .B1(n4881), .B2(n6331), .A(n6222), .ZN(n4620) );
  NAND3_X1 U5711 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6460), .A3(n6456), .ZN(n6228) );
  OR2_X1 U5712 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6228), .ZN(n4920)
         );
  NOR2_X1 U5713 ( .A1(n4621), .A2(n6583), .ZN(n6340) );
  INV_X1 U5714 ( .A(n4689), .ZN(n6339) );
  NOR2_X1 U5715 ( .A1(n6339), .A2(n4690), .ZN(n4662) );
  OAI21_X1 U5716 ( .B1(n4662), .B2(n6583), .A(n4757), .ZN(n4659) );
  AOI211_X1 U5717 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4920), .A(n6340), .B(
        n4659), .ZN(n4619) );
  NAND2_X1 U5718 ( .A1(n4919), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4626) );
  INV_X2 U5719 ( .A(n5564), .ZN(n6101) );
  AND2_X1 U5720 ( .A1(n6101), .A2(DATAI_27_), .ZN(n6414) );
  NAND2_X1 U5721 ( .A1(DATAI_3_), .A2(n4757), .ZN(n6418) );
  NOR2_X1 U5722 ( .A1(n3101), .A2(n6393), .ZN(n6192) );
  INV_X1 U5723 ( .A(n5733), .ZN(n5741) );
  AND2_X1 U5724 ( .A1(n4621), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6258) );
  AOI22_X1 U5725 ( .A1(n6192), .A2(n5741), .B1(n6258), .B2(n4662), .ZN(n4921)
         );
  NAND2_X1 U5726 ( .A1(n6586), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6562) );
  INV_X1 U5727 ( .A(n6562), .ZN(n5102) );
  INV_X1 U5728 ( .A(n6413), .ZN(n5759) );
  OAI22_X1 U5729 ( .A1(n6418), .A2(n4921), .B1(n5759), .B2(n4920), .ZN(n4624)
         );
  AOI21_X1 U5730 ( .B1(n6414), .B2(n4923), .A(n4624), .ZN(n4625) );
  OAI211_X1 U5731 ( .C1(n6231), .C2(n6281), .A(n4626), .B(n4625), .ZN(U3055)
         );
  NAND2_X1 U5732 ( .A1(n6101), .A2(DATAI_23_), .ZN(n6297) );
  NAND2_X1 U5733 ( .A1(n4919), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4629) );
  NAND2_X1 U5734 ( .A1(DATAI_7_), .A2(n4757), .ZN(n6446) );
  INV_X1 U5735 ( .A(n6438), .ZN(n5781) );
  OAI22_X1 U5736 ( .A1(n6446), .A2(n4921), .B1(n5781), .B2(n4920), .ZN(n4627)
         );
  AOI21_X1 U5737 ( .B1(n6442), .B2(n4923), .A(n4627), .ZN(n4628) );
  OAI211_X1 U5738 ( .C1(n6231), .C2(n6297), .A(n4629), .B(n4628), .ZN(U3059)
         );
  AND2_X1 U5739 ( .A1(n6101), .A2(DATAI_17_), .ZN(n6403) );
  INV_X1 U5740 ( .A(n6403), .ZN(n6275) );
  NAND2_X1 U5741 ( .A1(n4919), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4632) );
  NAND2_X1 U5742 ( .A1(n6101), .A2(DATAI_25_), .ZN(n5753) );
  INV_X1 U5743 ( .A(n5753), .ZN(n6402) );
  NAND2_X1 U5744 ( .A1(DATAI_1_), .A2(n4757), .ZN(n6406) );
  INV_X1 U5745 ( .A(n6401), .ZN(n5749) );
  OAI22_X1 U5746 ( .A1(n6406), .A2(n4921), .B1(n5749), .B2(n4920), .ZN(n4630)
         );
  AOI21_X1 U5747 ( .B1(n6402), .B2(n4923), .A(n4630), .ZN(n4631) );
  OAI211_X1 U5748 ( .C1(n6231), .C2(n6275), .A(n4632), .B(n4631), .ZN(U3053)
         );
  AND2_X1 U5749 ( .A1(n5958), .A2(n4633), .ZN(n4634) );
  OR2_X1 U5750 ( .A1(n4634), .A2(n4735), .ZN(n6128) );
  INV_X1 U5751 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4635) );
  OAI222_X1 U5752 ( .A1(n6128), .A2(n5376), .B1(n6026), .B2(n4635), .C1(n3092), 
        .C2(n4824), .ZN(U2852) );
  INV_X1 U5753 ( .A(n6442), .ZN(n5787) );
  INV_X1 U5754 ( .A(n6297), .ZN(n6439) );
  NAND2_X1 U5755 ( .A1(n4576), .A2(n6226), .ZN(n6329) );
  NOR2_X1 U5756 ( .A1(n6329), .A2(n4589), .ZN(n4637) );
  NOR2_X1 U5757 ( .A1(n5040), .A2(n6393), .ZN(n5742) );
  INV_X1 U5758 ( .A(n6258), .ZN(n4699) );
  NOR3_X1 U5759 ( .A1(n4699), .A2(n6460), .A3(n4689), .ZN(n4638) );
  AOI21_X1 U5760 ( .B1(n5742), .B2(n6264), .A(n4638), .ZN(n4961) );
  INV_X1 U5761 ( .A(n4772), .ZN(n4775) );
  NOR2_X1 U5762 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4775), .ZN(n4643)
         );
  INV_X1 U5763 ( .A(n4643), .ZN(n4960) );
  OAI22_X1 U5764 ( .A1(n6446), .A2(n4961), .B1(n5781), .B2(n4960), .ZN(n4639)
         );
  AOI21_X1 U5765 ( .B1(n6439), .B2(n4963), .A(n4639), .ZN(n4647) );
  INV_X1 U5766 ( .A(n4963), .ZN(n4640) );
  NAND3_X1 U5767 ( .A1(n4967), .A2(n4640), .A3(n6380), .ZN(n4641) );
  AOI22_X1 U5768 ( .A1(n4641), .A2(n6265), .B1(n6264), .B2(n3101), .ZN(n4645)
         );
  NAND2_X1 U5769 ( .A1(n4689), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4642) );
  NAND2_X1 U5770 ( .A1(n4757), .A2(n4642), .ZN(n6269) );
  INV_X1 U5771 ( .A(n6340), .ZN(n5737) );
  NAND2_X1 U5772 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6460), .ZN(n6335) );
  OAI211_X1 U5773 ( .C1(n4643), .C2(n6688), .A(n5737), .B(n6335), .ZN(n4644)
         );
  NAND2_X1 U5774 ( .A1(n4964), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4646)
         );
  OAI211_X1 U5775 ( .C1(n4967), .C2(n5787), .A(n4647), .B(n4646), .ZN(U3139)
         );
  OAI22_X1 U5776 ( .A1(n6406), .A2(n4961), .B1(n5749), .B2(n4960), .ZN(n4648)
         );
  AOI21_X1 U5777 ( .B1(n6403), .B2(n4963), .A(n4648), .ZN(n4650) );
  NAND2_X1 U5778 ( .A1(n4964), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4649)
         );
  OAI211_X1 U5779 ( .C1(n4967), .C2(n5753), .A(n4650), .B(n4649), .ZN(U3133)
         );
  INV_X1 U5780 ( .A(n6414), .ZN(n5763) );
  OAI22_X1 U5781 ( .A1(n6418), .A2(n4961), .B1(n5759), .B2(n4960), .ZN(n4651)
         );
  AOI21_X1 U5782 ( .B1(n6415), .B2(n4963), .A(n4651), .ZN(n4653) );
  NAND2_X1 U5783 ( .A1(n4964), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4652)
         );
  OAI211_X1 U5784 ( .C1(n4967), .C2(n5763), .A(n4653), .B(n4652), .ZN(U3135)
         );
  OAI21_X1 U5785 ( .B1(n3118), .B2(n4654), .A(n5956), .ZN(n5967) );
  XOR2_X1 U5786 ( .A(n4506), .B(n4655), .Z(n6833) );
  INV_X1 U5787 ( .A(n6833), .ZN(n4656) );
  OAI222_X1 U5788 ( .A1(n5376), .A2(n5967), .B1(n6026), .B2(n6811), .C1(n3092), 
        .C2(n4656), .ZN(U2854) );
  NAND3_X1 U5789 ( .A1(n4770), .A2(n4769), .A3(n4720), .ZN(n4981) );
  NOR2_X1 U5790 ( .A1(n4696), .A2(n3101), .ZN(n4978) );
  AND2_X1 U5791 ( .A1(n5731), .A2(n3468), .ZN(n4657) );
  NOR2_X1 U5792 ( .A1(n4942), .A2(n6393), .ZN(n4658) );
  AOI21_X1 U5793 ( .B1(n4980), .B2(n4658), .A(n6331), .ZN(n4661) );
  NAND3_X1 U5794 ( .A1(n6460), .A2(n6334), .A3(n6456), .ZN(n4983) );
  OR2_X1 U5795 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4983), .ZN(n4939)
         );
  AOI211_X1 U5796 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4939), .A(n6258), .B(
        n4659), .ZN(n4660) );
  NAND2_X1 U5797 ( .A1(n4938), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4665) );
  AOI22_X1 U5798 ( .A1(n4978), .A2(n6380), .B1(n6340), .B2(n4662), .ZN(n4940)
         );
  OAI22_X1 U5799 ( .A1(n6406), .A2(n4940), .B1(n5749), .B2(n4939), .ZN(n4663)
         );
  AOI21_X1 U5800 ( .B1(n6402), .B2(n4942), .A(n4663), .ZN(n4664) );
  OAI211_X1 U5801 ( .C1(n4980), .C2(n6275), .A(n4665), .B(n4664), .ZN(U3021)
         );
  NAND2_X1 U5802 ( .A1(n4938), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4668) );
  OAI22_X1 U5803 ( .A1(n6446), .A2(n4940), .B1(n5781), .B2(n4939), .ZN(n4666)
         );
  AOI21_X1 U5804 ( .B1(n6442), .B2(n4942), .A(n4666), .ZN(n4667) );
  OAI211_X1 U5805 ( .C1(n4980), .C2(n6297), .A(n4668), .B(n4667), .ZN(U3027)
         );
  NAND2_X1 U5806 ( .A1(n4938), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4671) );
  OAI22_X1 U5807 ( .A1(n6418), .A2(n4940), .B1(n5759), .B2(n4939), .ZN(n4669)
         );
  AOI21_X1 U5808 ( .B1(n6414), .B2(n4942), .A(n4669), .ZN(n4670) );
  OAI211_X1 U5809 ( .C1(n4980), .C2(n6281), .A(n4671), .B(n4670), .ZN(U3023)
         );
  OAI21_X1 U5810 ( .B1(n4674), .B2(n4673), .A(n4672), .ZN(n4977) );
  AOI22_X1 U5811 ( .A1(n6831), .A2(DATAI_8_), .B1(n6830), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4675) );
  OAI21_X1 U5812 ( .B1(n4977), .B2(n5418), .A(n4675), .ZN(U2883) );
  NAND2_X1 U5813 ( .A1(n6379), .A2(n4769), .ZN(n4682) );
  INV_X1 U5814 ( .A(n4682), .ZN(n4676) );
  AND2_X1 U5815 ( .A1(n3101), .A2(n3102), .ZN(n6384) );
  INV_X1 U5816 ( .A(n4696), .ZN(n4691) );
  NAND3_X1 U5817 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6334), .A3(n6456), .ZN(n4692) );
  NOR2_X1 U5818 ( .A1(n6451), .A2(n4692), .ZN(n4811) );
  AOI21_X1 U5819 ( .B1(n6384), .B2(n4691), .A(n4811), .ZN(n4681) );
  NAND3_X1 U5820 ( .A1(n6379), .A2(n4769), .A3(STATEBS16_REG_SCAN_IN), .ZN(
        n4677) );
  AND2_X1 U5821 ( .A1(n4677), .A2(n6380), .ZN(n4679) );
  AOI22_X1 U5822 ( .A1(n4681), .A2(n4679), .B1(n6393), .B2(n4692), .ZN(n4678)
         );
  NAND2_X1 U5823 ( .A1(n6306), .A2(n4678), .ZN(n4810) );
  INV_X1 U5824 ( .A(n4679), .ZN(n4680) );
  OAI22_X1 U5825 ( .A1(n4681), .A2(n4680), .B1(n6583), .B2(n4692), .ZN(n4809)
         );
  AOI22_X1 U5826 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4810), .B1(n6347), 
        .B2(n4809), .ZN(n4684) );
  NOR2_X2 U5827 ( .A1(n4682), .A2(n6226), .ZN(n6372) );
  AOI22_X1 U5828 ( .A1(n6372), .A2(n6403), .B1(n4811), .B2(n6401), .ZN(n4683)
         );
  OAI211_X1 U5829 ( .C1(n4906), .C2(n5753), .A(n4684), .B(n4683), .ZN(U3093)
         );
  AOI22_X1 U5830 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4810), .B1(n6373), 
        .B2(n4809), .ZN(n4686) );
  AOI22_X1 U5831 ( .A1(n6372), .A2(n6439), .B1(n4811), .B2(n6438), .ZN(n4685)
         );
  OAI211_X1 U5832 ( .C1(n4906), .C2(n5787), .A(n4686), .B(n4685), .ZN(U3099)
         );
  AOI22_X1 U5833 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4810), .B1(n6355), 
        .B2(n4809), .ZN(n4688) );
  AOI22_X1 U5834 ( .A1(n6372), .A2(n6415), .B1(n4811), .B2(n6413), .ZN(n4687)
         );
  OAI211_X1 U5835 ( .C1(n4906), .C2(n5763), .A(n4688), .B(n4687), .ZN(U3095)
         );
  NAND2_X1 U5836 ( .A1(n4690), .A2(n4689), .ZN(n4698) );
  INV_X1 U5837 ( .A(n4698), .ZN(n5740) );
  AOI22_X1 U5838 ( .A1(n5742), .A2(n4691), .B1(n6340), .B2(n5740), .ZN(n4901)
         );
  NOR2_X1 U5839 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4692), .ZN(n4700)
         );
  INV_X1 U5840 ( .A(n4700), .ZN(n4900) );
  OAI22_X1 U5841 ( .A1(n6418), .A2(n4901), .B1(n5759), .B2(n4900), .ZN(n4693)
         );
  AOI21_X1 U5842 ( .B1(n6414), .B2(n6322), .A(n4693), .ZN(n4705) );
  INV_X1 U5843 ( .A(n4906), .ZN(n4694) );
  OAI21_X1 U5844 ( .B1(n4694), .B2(n6322), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4695) );
  OAI211_X1 U5845 ( .C1(n5040), .C2(n4696), .A(n4695), .B(n6380), .ZN(n4703)
         );
  AOI21_X1 U5846 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4698), .A(n4697), .ZN(
        n5738) );
  OAI21_X1 U5847 ( .B1(n6688), .B2(n4700), .A(n4699), .ZN(n4701) );
  INV_X1 U5848 ( .A(n4701), .ZN(n4702) );
  NAND3_X1 U5849 ( .A1(n4703), .A2(n5738), .A3(n4702), .ZN(n4903) );
  NAND2_X1 U5850 ( .A1(n4903), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4704) );
  OAI211_X1 U5851 ( .C1(n6281), .C2(n4906), .A(n4705), .B(n4704), .ZN(U3087)
         );
  OAI22_X1 U5852 ( .A1(n6446), .A2(n4901), .B1(n5781), .B2(n4900), .ZN(n4706)
         );
  AOI21_X1 U5853 ( .B1(n6442), .B2(n6322), .A(n4706), .ZN(n4708) );
  NAND2_X1 U5854 ( .A1(n4903), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4707) );
  OAI211_X1 U5855 ( .C1(n6297), .C2(n4906), .A(n4708), .B(n4707), .ZN(U3091)
         );
  OAI22_X1 U5856 ( .A1(n6406), .A2(n4901), .B1(n5749), .B2(n4900), .ZN(n4709)
         );
  AOI21_X1 U5857 ( .B1(n6402), .B2(n6322), .A(n4709), .ZN(n4711) );
  NAND2_X1 U5858 ( .A1(n4903), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4710) );
  OAI211_X1 U5859 ( .C1(n6275), .C2(n4906), .A(n4711), .B(n4710), .ZN(U3085)
         );
  NOR2_X1 U5860 ( .A1(n4713), .A2(n4712), .ZN(n4714) );
  AOI21_X1 U5861 ( .B1(n4715), .B2(n4714), .A(n6393), .ZN(n4722) );
  OR2_X1 U5862 ( .A1(n4523), .A2(n4716), .ZN(n6194) );
  INV_X1 U5863 ( .A(n6194), .ZN(n6383) );
  NAND2_X1 U5864 ( .A1(n6383), .A2(n5040), .ZN(n6198) );
  INV_X1 U5865 ( .A(n3102), .ZN(n5027) );
  OR2_X1 U5866 ( .A1(n6198), .A2(n5027), .ZN(n4718) );
  INV_X1 U5867 ( .A(n6382), .ZN(n4717) );
  NAND2_X1 U5868 ( .A1(n4717), .A2(n6460), .ZN(n4882) );
  NAND2_X1 U5869 ( .A1(n4718), .A2(n4882), .ZN(n4724) );
  NAND3_X1 U5870 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6460), .A3(n6334), .ZN(n6195) );
  INV_X1 U5871 ( .A(n6195), .ZN(n4719) );
  AOI22_X1 U5872 ( .A1(n4722), .A2(n4724), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4719), .ZN(n4887) );
  INV_X1 U5873 ( .A(n6329), .ZN(n6256) );
  NAND3_X1 U5874 ( .A1(n4770), .A2(n6256), .A3(n4720), .ZN(n6221) );
  OAI22_X1 U5875 ( .A1(n5781), .A2(n4882), .B1(n6297), .B2(n4881), .ZN(n4721)
         );
  AOI21_X1 U5876 ( .B1(n6442), .B2(n6197), .A(n4721), .ZN(n4727) );
  INV_X1 U5877 ( .A(n4722), .ZN(n4725) );
  INV_X1 U5878 ( .A(n6306), .ZN(n6391) );
  AOI21_X1 U5879 ( .B1(n6393), .B2(n6195), .A(n6391), .ZN(n4723) );
  NAND2_X1 U5880 ( .A1(n4884), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4726) );
  OAI211_X1 U5881 ( .C1(n4887), .C2(n6446), .A(n4727), .B(n4726), .ZN(U3051)
         );
  OAI22_X1 U5882 ( .A1(n5759), .A2(n4882), .B1(n6281), .B2(n4881), .ZN(n4728)
         );
  AOI21_X1 U5883 ( .B1(n6414), .B2(n6197), .A(n4728), .ZN(n4730) );
  NAND2_X1 U5884 ( .A1(n4884), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4729) );
  OAI211_X1 U5885 ( .C1(n4887), .C2(n6418), .A(n4730), .B(n4729), .ZN(U3047)
         );
  OAI22_X1 U5886 ( .A1(n5749), .A2(n4882), .B1(n6275), .B2(n4881), .ZN(n4731)
         );
  AOI21_X1 U5887 ( .B1(n6402), .B2(n6197), .A(n4731), .ZN(n4733) );
  NAND2_X1 U5888 ( .A1(n4884), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4732) );
  OAI211_X1 U5889 ( .C1(n4887), .C2(n6406), .A(n4733), .B(n4732), .ZN(U3045)
         );
  INV_X1 U5890 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4737) );
  NOR2_X1 U5891 ( .A1(n4735), .A2(n4734), .ZN(n4736) );
  OR2_X1 U5892 ( .A1(n5035), .A2(n4736), .ZN(n4830) );
  OAI222_X1 U5893 ( .A1(n4977), .A2(n3092), .B1(n6026), .B2(n4737), .C1(n5376), 
        .C2(n4830), .ZN(U2851) );
  AND2_X1 U5894 ( .A1(n6101), .A2(DATAI_22_), .ZN(n6433) );
  INV_X1 U5895 ( .A(n6433), .ZN(n6290) );
  NOR3_X1 U5896 ( .A1(n6334), .A2(n6460), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4739) );
  INV_X1 U5897 ( .A(n4739), .ZN(n5735) );
  NOR2_X1 U5898 ( .A1(n6451), .A2(n5735), .ZN(n4763) );
  AOI21_X1 U5899 ( .B1(n6384), .B2(n5741), .A(n4763), .ZN(n4742) );
  NAND3_X1 U5900 ( .A1(n6380), .A2(n4742), .A3(n4740), .ZN(n4738) );
  OAI211_X1 U5901 ( .C1(n6380), .C2(n4739), .A(n6306), .B(n4738), .ZN(n4762)
         );
  NAND2_X1 U5902 ( .A1(DATAI_6_), .A2(n4757), .ZN(n6436) );
  NAND2_X1 U5903 ( .A1(n6380), .A2(n4740), .ZN(n4741) );
  OAI22_X1 U5904 ( .A1(n4742), .A2(n4741), .B1(n6583), .B2(n5735), .ZN(n4761)
         );
  AOI22_X1 U5905 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4762), .B1(n6367), 
        .B2(n4761), .ZN(n4745) );
  NOR2_X1 U5906 ( .A1(n4758), .A2(n3493), .ZN(n6431) );
  NOR2_X2 U5907 ( .A1(n4743), .A2(n5728), .ZN(n5784) );
  AOI22_X1 U5908 ( .A1(n6431), .A2(n4763), .B1(n6432), .B2(n5784), .ZN(n4744)
         );
  OAI211_X1 U5909 ( .C1(n6290), .C2(n4967), .A(n4745), .B(n4744), .ZN(U3130)
         );
  NAND2_X1 U5910 ( .A1(n6101), .A2(DATAI_18_), .ZN(n6278) );
  NAND2_X1 U5911 ( .A1(DATAI_2_), .A2(n4757), .ZN(n6412) );
  AOI22_X1 U5912 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4762), .B1(n6351), 
        .B2(n4761), .ZN(n4748) );
  AOI22_X1 U5913 ( .A1(n6407), .A2(n4763), .B1(n6409), .B2(n5784), .ZN(n4747)
         );
  OAI211_X1 U5914 ( .C1(n6278), .C2(n4967), .A(n4748), .B(n4747), .ZN(U3126)
         );
  AOI22_X1 U5915 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4762), .B1(n6355), 
        .B2(n4761), .ZN(n4750) );
  AOI22_X1 U5916 ( .A1(n6413), .A2(n4763), .B1(n6414), .B2(n5784), .ZN(n4749)
         );
  OAI211_X1 U5917 ( .C1(n6281), .C2(n4967), .A(n4750), .B(n4749), .ZN(U3127)
         );
  AND2_X1 U5918 ( .A1(n6101), .A2(DATAI_21_), .ZN(n6427) );
  INV_X1 U5919 ( .A(n6427), .ZN(n6287) );
  NAND2_X1 U5920 ( .A1(DATAI_5_), .A2(n4757), .ZN(n6430) );
  AOI22_X1 U5921 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4762), .B1(n6363), 
        .B2(n4761), .ZN(n4752) );
  AOI22_X1 U5922 ( .A1(n6425), .A2(n4763), .B1(n6426), .B2(n5784), .ZN(n4751)
         );
  OAI211_X1 U5923 ( .C1(n6287), .C2(n4967), .A(n4752), .B(n4751), .ZN(U3129)
         );
  AND2_X1 U5924 ( .A1(n6101), .A2(DATAI_20_), .ZN(n6421) );
  INV_X1 U5925 ( .A(n6421), .ZN(n6284) );
  NAND2_X1 U5926 ( .A1(DATAI_4_), .A2(n4757), .ZN(n6424) );
  AOI22_X1 U5927 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4762), .B1(n6359), 
        .B2(n4761), .ZN(n4754) );
  NOR2_X1 U5928 ( .A1(n4758), .A2(n3377), .ZN(n6419) );
  AOI22_X1 U5929 ( .A1(n6419), .A2(n4763), .B1(n6420), .B2(n5784), .ZN(n4753)
         );
  OAI211_X1 U5930 ( .C1(n6284), .C2(n4967), .A(n4754), .B(n4753), .ZN(U3128)
         );
  AOI22_X1 U5931 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4762), .B1(n6373), 
        .B2(n4761), .ZN(n4756) );
  AOI22_X1 U5932 ( .A1(n6438), .A2(n4763), .B1(n6442), .B2(n5784), .ZN(n4755)
         );
  OAI211_X1 U5933 ( .C1(n6297), .C2(n4967), .A(n4756), .B(n4755), .ZN(U3131)
         );
  AND2_X1 U5934 ( .A1(n6101), .A2(DATAI_16_), .ZN(n6389) );
  INV_X1 U5935 ( .A(n6389), .ZN(n6272) );
  NAND2_X1 U5936 ( .A1(DATAI_0_), .A2(n4757), .ZN(n6400) );
  AOI22_X1 U5937 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4762), .B1(n6344), 
        .B2(n4761), .ZN(n4760) );
  NOR2_X1 U5938 ( .A1(n4758), .A2(n3324), .ZN(n6388) );
  AOI22_X1 U5939 ( .A1(n6388), .A2(n4763), .B1(n6397), .B2(n5784), .ZN(n4759)
         );
  OAI211_X1 U5940 ( .C1(n6272), .C2(n4967), .A(n4760), .B(n4759), .ZN(U3124)
         );
  AOI22_X1 U5941 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4762), .B1(n6347), 
        .B2(n4761), .ZN(n4765) );
  AOI22_X1 U5942 ( .A1(n6401), .A2(n4763), .B1(n6402), .B2(n5784), .ZN(n4764)
         );
  OAI211_X1 U5943 ( .C1(n6275), .C2(n4967), .A(n4765), .B(n4764), .ZN(U3125)
         );
  INV_X1 U5944 ( .A(n6397), .ZN(n5748) );
  AOI22_X1 U5945 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4810), .B1(n6344), 
        .B2(n4809), .ZN(n4767) );
  AOI22_X1 U5946 ( .A1(n6372), .A2(n6389), .B1(n6388), .B2(n4811), .ZN(n4766)
         );
  OAI211_X1 U5947 ( .C1(n5748), .C2(n4906), .A(n4767), .B(n4766), .ZN(U3092)
         );
  INV_X1 U5948 ( .A(n4768), .ZN(n4797) );
  AOI21_X1 U5949 ( .B1(n6384), .B2(n6264), .A(n4797), .ZN(n4776) );
  NOR3_X1 U5950 ( .A1(n4770), .A2(n4589), .A3(n4769), .ZN(n4771) );
  OAI21_X1 U5951 ( .B1(n4771), .B2(n5564), .A(n6265), .ZN(n4774) );
  OAI21_X1 U5952 ( .B1(n4772), .B2(n6380), .A(n6306), .ZN(n4773) );
  INV_X1 U5953 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4779) );
  OAI22_X1 U5954 ( .A1(n4776), .A2(n6393), .B1(n4775), .B2(n6583), .ZN(n4798)
         );
  AOI22_X1 U5955 ( .A1(n6359), .A2(n4798), .B1(n4797), .B2(n6419), .ZN(n4778)
         );
  AOI22_X1 U5956 ( .A1(n6421), .A2(n4942), .B1(n4963), .B2(n6420), .ZN(n4777)
         );
  OAI211_X1 U5957 ( .C1(n4802), .C2(n4779), .A(n4778), .B(n4777), .ZN(U3144)
         );
  INV_X1 U5958 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4782) );
  AOI22_X1 U5959 ( .A1(n6344), .A2(n4798), .B1(n4797), .B2(n6388), .ZN(n4781)
         );
  AOI22_X1 U5960 ( .A1(n6389), .A2(n4942), .B1(n4963), .B2(n6397), .ZN(n4780)
         );
  OAI211_X1 U5961 ( .C1(n4802), .C2(n4782), .A(n4781), .B(n4780), .ZN(U3140)
         );
  INV_X1 U5962 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4785) );
  AOI22_X1 U5963 ( .A1(n6363), .A2(n4798), .B1(n4797), .B2(n6425), .ZN(n4784)
         );
  AOI22_X1 U5964 ( .A1(n6427), .A2(n4942), .B1(n4963), .B2(n6426), .ZN(n4783)
         );
  OAI211_X1 U5965 ( .C1(n4802), .C2(n4785), .A(n4784), .B(n4783), .ZN(U3145)
         );
  INV_X1 U5966 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4788) );
  AOI22_X1 U5967 ( .A1(n6351), .A2(n4798), .B1(n4797), .B2(n6407), .ZN(n4787)
         );
  INV_X1 U5968 ( .A(n6278), .ZN(n6408) );
  AOI22_X1 U5969 ( .A1(n6408), .A2(n4942), .B1(n4963), .B2(n6409), .ZN(n4786)
         );
  OAI211_X1 U5970 ( .C1(n4802), .C2(n4788), .A(n4787), .B(n4786), .ZN(U3142)
         );
  INV_X1 U5971 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4791) );
  AOI22_X1 U5972 ( .A1(n6367), .A2(n4798), .B1(n4797), .B2(n6431), .ZN(n4790)
         );
  AOI22_X1 U5973 ( .A1(n6433), .A2(n4942), .B1(n4963), .B2(n6432), .ZN(n4789)
         );
  OAI211_X1 U5974 ( .C1(n4802), .C2(n4791), .A(n4790), .B(n4789), .ZN(U3146)
         );
  INV_X1 U5975 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4794) );
  AOI22_X1 U5976 ( .A1(n6355), .A2(n4798), .B1(n4797), .B2(n6413), .ZN(n4793)
         );
  AOI22_X1 U5977 ( .A1(n6415), .A2(n4942), .B1(n4963), .B2(n6414), .ZN(n4792)
         );
  OAI211_X1 U5978 ( .C1(n4802), .C2(n4794), .A(n4793), .B(n4792), .ZN(U3143)
         );
  AOI22_X1 U5979 ( .A1(n6373), .A2(n4798), .B1(n4797), .B2(n6438), .ZN(n4796)
         );
  AOI22_X1 U5980 ( .A1(n6439), .A2(n4942), .B1(n4963), .B2(n6442), .ZN(n4795)
         );
  OAI211_X1 U5981 ( .C1(n4802), .C2(n3822), .A(n4796), .B(n4795), .ZN(U3147)
         );
  INV_X1 U5982 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4801) );
  AOI22_X1 U5983 ( .A1(n6347), .A2(n4798), .B1(n4797), .B2(n6401), .ZN(n4800)
         );
  AOI22_X1 U5984 ( .A1(n6403), .A2(n4942), .B1(n4963), .B2(n6402), .ZN(n4799)
         );
  OAI211_X1 U5985 ( .C1(n4802), .C2(n4801), .A(n4800), .B(n4799), .ZN(U3141)
         );
  INV_X1 U5986 ( .A(n6432), .ZN(n5778) );
  AOI22_X1 U5987 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4810), .B1(n6367), 
        .B2(n4809), .ZN(n4804) );
  AOI22_X1 U5988 ( .A1(n6372), .A2(n6433), .B1(n4811), .B2(n6431), .ZN(n4803)
         );
  OAI211_X1 U5989 ( .C1(n4906), .C2(n5778), .A(n4804), .B(n4803), .ZN(U3098)
         );
  INV_X1 U5990 ( .A(n6426), .ZN(n5773) );
  AOI22_X1 U5991 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4810), .B1(n6363), 
        .B2(n4809), .ZN(n4806) );
  AOI22_X1 U5992 ( .A1(n6372), .A2(n6427), .B1(n4811), .B2(n6425), .ZN(n4805)
         );
  OAI211_X1 U5993 ( .C1(n4906), .C2(n5773), .A(n4806), .B(n4805), .ZN(U3097)
         );
  INV_X1 U5994 ( .A(n6420), .ZN(n5768) );
  AOI22_X1 U5995 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4810), .B1(n6359), 
        .B2(n4809), .ZN(n4808) );
  AOI22_X1 U5996 ( .A1(n6372), .A2(n6421), .B1(n4811), .B2(n6419), .ZN(n4807)
         );
  OAI211_X1 U5997 ( .C1(n4906), .C2(n5768), .A(n4808), .B(n4807), .ZN(U3096)
         );
  INV_X1 U5998 ( .A(n6409), .ZN(n5758) );
  AOI22_X1 U5999 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4810), .B1(n6351), 
        .B2(n4809), .ZN(n4813) );
  AOI22_X1 U6000 ( .A1(n6372), .A2(n6408), .B1(n4811), .B2(n6407), .ZN(n4812)
         );
  OAI211_X1 U6001 ( .C1(n4906), .C2(n5758), .A(n4813), .B(n4812), .ZN(U3094)
         );
  INV_X1 U6002 ( .A(n4859), .ZN(n4822) );
  INV_X1 U6003 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6126) );
  NAND2_X1 U6004 ( .A1(n5044), .A2(n4814), .ZN(n4815) );
  NAND2_X1 U6005 ( .A1(n5921), .A2(n4815), .ZN(n5976) );
  OAI22_X1 U6006 ( .A1(n5947), .A2(n6128), .B1(n6126), .B2(n5976), .ZN(n4821)
         );
  NOR2_X1 U6007 ( .A1(n5983), .A2(n4816), .ZN(n5966) );
  INV_X1 U6008 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6518) );
  NOR2_X1 U6009 ( .A1(n6126), .A2(n6518), .ZN(n4834) );
  AOI21_X1 U6010 ( .B1(n6126), .B2(n6518), .A(n4834), .ZN(n4817) );
  AOI22_X1 U6011 ( .A1(EBX_REG_7__SCAN_IN), .A2(n5995), .B1(n5960), .B2(n4817), 
        .ZN(n4818) );
  NAND3_X1 U6012 ( .A1(n6858), .A2(n5044), .A3(n6380), .ZN(n5944) );
  OAI211_X1 U6013 ( .C1(n6000), .C2(n4819), .A(n4818), .B(n5944), .ZN(n4820)
         );
  AOI211_X1 U6014 ( .C1(n6006), .C2(n4822), .A(n4821), .B(n4820), .ZN(n4823)
         );
  OAI21_X1 U6015 ( .B1(n4824), .B2(n5842), .A(n4823), .ZN(U2820) );
  INV_X1 U6016 ( .A(n6001), .ZN(n6024) );
  AOI22_X1 U6017 ( .A1(n6097), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6156), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4826) );
  OAI21_X1 U6018 ( .B1(n6108), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4826), 
        .ZN(n4827) );
  AOI21_X1 U6019 ( .B1(n6101), .B2(n6024), .A(n4827), .ZN(n4828) );
  OAI21_X1 U6020 ( .B1(n4829), .B2(n6078), .A(n4828), .ZN(U2985) );
  INV_X1 U6021 ( .A(n4973), .ZN(n4839) );
  INV_X1 U6022 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4832) );
  INV_X1 U6023 ( .A(n4830), .ZN(n6119) );
  AOI22_X1 U6024 ( .A1(EBX_REG_8__SCAN_IN), .A2(n5995), .B1(n5980), .B2(n6119), 
        .ZN(n4831) );
  OAI211_X1 U6025 ( .C1(n6000), .C2(n4832), .A(n4831), .B(n5944), .ZN(n4838)
         );
  INV_X1 U6026 ( .A(n5921), .ZN(n5270) );
  NOR2_X1 U6027 ( .A1(n5998), .A2(n5919), .ZN(n4833) );
  NOR2_X1 U6028 ( .A1(n5270), .A2(n4833), .ZN(n5950) );
  INV_X1 U6029 ( .A(n5950), .ZN(n4836) );
  AOI21_X1 U6030 ( .B1(n5960), .B2(n4834), .A(REIP_REG_8__SCAN_IN), .ZN(n4835)
         );
  NOR2_X1 U6031 ( .A1(n4836), .A2(n4835), .ZN(n4837) );
  AOI211_X1 U6032 ( .C1(n6006), .C2(n4839), .A(n4838), .B(n4837), .ZN(n4840)
         );
  OAI21_X1 U6033 ( .B1(n5842), .B2(n4977), .A(n4840), .ZN(U2819) );
  OAI21_X1 U6034 ( .B1(n4843), .B2(n4842), .A(n4841), .ZN(n4844) );
  INV_X1 U6035 ( .A(n4844), .ZN(n6168) );
  INV_X1 U6036 ( .A(REIP_REG_3__SCAN_IN), .ZN(n4845) );
  NOR2_X1 U6037 ( .A1(n6190), .A2(n4845), .ZN(n6164) );
  AOI21_X1 U6038 ( .B1(n6097), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n6164), 
        .ZN(n4846) );
  OAI21_X1 U6039 ( .B1(n6108), .B2(n5041), .A(n4846), .ZN(n4847) );
  AOI21_X1 U6040 ( .B1(n6168), .B2(n6104), .A(n4847), .ZN(n4848) );
  OAI21_X1 U6041 ( .B1(n5050), .B2(n5564), .A(n4848), .ZN(U2983) );
  OAI21_X1 U6042 ( .B1(n4851), .B2(n4850), .A(n4849), .ZN(n6149) );
  AOI22_X1 U6043 ( .A1(n6097), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .B1(n6156), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n4852) );
  OAI21_X1 U6044 ( .B1(n6108), .B2(n5971), .A(n4852), .ZN(n4853) );
  AOI21_X1 U6045 ( .B1(n6833), .B2(n6101), .A(n4853), .ZN(n4854) );
  OAI21_X1 U6046 ( .B1(n6149), .B2(n6078), .A(n4854), .ZN(U2981) );
  OAI21_X1 U6047 ( .B1(n4857), .B2(n4856), .A(n3093), .ZN(n6125) );
  AOI22_X1 U6048 ( .A1(n6097), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .B1(n6156), 
        .B2(REIP_REG_7__SCAN_IN), .ZN(n4858) );
  OAI21_X1 U6049 ( .B1(n6108), .B2(n4859), .A(n4858), .ZN(n4860) );
  AOI21_X1 U6050 ( .B1(n4861), .B2(n6101), .A(n4860), .ZN(n4862) );
  OAI21_X1 U6051 ( .B1(n6125), .B2(n6078), .A(n4862), .ZN(U2979) );
  INV_X1 U6052 ( .A(n4863), .ZN(n4945) );
  INV_X1 U6053 ( .A(n4864), .ZN(n4865) );
  OAI21_X1 U6054 ( .B1(n4945), .B2(n4865), .A(n5371), .ZN(n5563) );
  AOI21_X1 U6055 ( .B1(n4866), .B2(n5037), .A(n3126), .ZN(n6110) );
  AOI22_X1 U6056 ( .A1(n6022), .A2(n6110), .B1(EBX_REG_10__SCAN_IN), .B2(n5368), .ZN(n4867) );
  OAI21_X1 U6057 ( .B1(n5563), .B2(n3092), .A(n4867), .ZN(U2849) );
  AOI22_X1 U6058 ( .A1(n6831), .A2(DATAI_10_), .B1(n6830), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n4868) );
  OAI21_X1 U6059 ( .B1(n5563), .B2(n5418), .A(n4868), .ZN(U2881) );
  INV_X1 U6060 ( .A(n6388), .ZN(n5744) );
  OAI22_X1 U6061 ( .A1(n5744), .A2(n4882), .B1(n6272), .B2(n4881), .ZN(n4869)
         );
  AOI21_X1 U6062 ( .B1(n6397), .B2(n6197), .A(n4869), .ZN(n4871) );
  NAND2_X1 U6063 ( .A1(n4884), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4870) );
  OAI211_X1 U6064 ( .C1(n4887), .C2(n6400), .A(n4871), .B(n4870), .ZN(U3044)
         );
  INV_X1 U6065 ( .A(n6407), .ZN(n5754) );
  OAI22_X1 U6066 ( .A1(n5754), .A2(n4882), .B1(n6278), .B2(n4881), .ZN(n4872)
         );
  AOI21_X1 U6067 ( .B1(n6409), .B2(n6197), .A(n4872), .ZN(n4874) );
  NAND2_X1 U6068 ( .A1(n4884), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4873) );
  OAI211_X1 U6069 ( .C1(n4887), .C2(n6412), .A(n4874), .B(n4873), .ZN(U3046)
         );
  INV_X1 U6070 ( .A(n6425), .ZN(n5769) );
  OAI22_X1 U6071 ( .A1(n5769), .A2(n4882), .B1(n6287), .B2(n4881), .ZN(n4875)
         );
  AOI21_X1 U6072 ( .B1(n6426), .B2(n6197), .A(n4875), .ZN(n4877) );
  NAND2_X1 U6073 ( .A1(n4884), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4876) );
  OAI211_X1 U6074 ( .C1(n4887), .C2(n6430), .A(n4877), .B(n4876), .ZN(U3049)
         );
  INV_X1 U6075 ( .A(n6431), .ZN(n5774) );
  OAI22_X1 U6076 ( .A1(n5774), .A2(n4882), .B1(n6290), .B2(n4881), .ZN(n4878)
         );
  AOI21_X1 U6077 ( .B1(n6432), .B2(n6197), .A(n4878), .ZN(n4880) );
  NAND2_X1 U6078 ( .A1(n4884), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4879) );
  OAI211_X1 U6079 ( .C1(n4887), .C2(n6436), .A(n4880), .B(n4879), .ZN(U3050)
         );
  INV_X1 U6080 ( .A(n6419), .ZN(n5764) );
  OAI22_X1 U6081 ( .A1(n5764), .A2(n4882), .B1(n6284), .B2(n4881), .ZN(n4883)
         );
  AOI21_X1 U6082 ( .B1(n6420), .B2(n6197), .A(n4883), .ZN(n4886) );
  NAND2_X1 U6083 ( .A1(n4884), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4885) );
  OAI211_X1 U6084 ( .C1(n4887), .C2(n6424), .A(n4886), .B(n4885), .ZN(U3048)
         );
  OAI22_X1 U6085 ( .A1(n6400), .A2(n4901), .B1(n5744), .B2(n4900), .ZN(n4888)
         );
  AOI21_X1 U6086 ( .B1(n6397), .B2(n6322), .A(n4888), .ZN(n4890) );
  NAND2_X1 U6087 ( .A1(n4903), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4889) );
  OAI211_X1 U6088 ( .C1(n6272), .C2(n4906), .A(n4890), .B(n4889), .ZN(U3084)
         );
  OAI22_X1 U6089 ( .A1(n6412), .A2(n4901), .B1(n5754), .B2(n4900), .ZN(n4891)
         );
  AOI21_X1 U6090 ( .B1(n6409), .B2(n6322), .A(n4891), .ZN(n4893) );
  NAND2_X1 U6091 ( .A1(n4903), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4892) );
  OAI211_X1 U6092 ( .C1(n6278), .C2(n4906), .A(n4893), .B(n4892), .ZN(U3086)
         );
  OAI22_X1 U6093 ( .A1(n6430), .A2(n4901), .B1(n5769), .B2(n4900), .ZN(n4894)
         );
  AOI21_X1 U6094 ( .B1(n6426), .B2(n6322), .A(n4894), .ZN(n4896) );
  NAND2_X1 U6095 ( .A1(n4903), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4895) );
  OAI211_X1 U6096 ( .C1(n6287), .C2(n4906), .A(n4896), .B(n4895), .ZN(U3089)
         );
  OAI22_X1 U6097 ( .A1(n6436), .A2(n4901), .B1(n5774), .B2(n4900), .ZN(n4897)
         );
  AOI21_X1 U6098 ( .B1(n6432), .B2(n6322), .A(n4897), .ZN(n4899) );
  NAND2_X1 U6099 ( .A1(n4903), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4898) );
  OAI211_X1 U6100 ( .C1(n6290), .C2(n4906), .A(n4899), .B(n4898), .ZN(U3090)
         );
  OAI22_X1 U6101 ( .A1(n6424), .A2(n4901), .B1(n5764), .B2(n4900), .ZN(n4902)
         );
  AOI21_X1 U6102 ( .B1(n6420), .B2(n6322), .A(n4902), .ZN(n4905) );
  NAND2_X1 U6103 ( .A1(n4903), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4904) );
  OAI211_X1 U6104 ( .C1(n6284), .C2(n4906), .A(n4905), .B(n4904), .ZN(U3088)
         );
  NAND2_X1 U6105 ( .A1(n4919), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4909) );
  OAI22_X1 U6106 ( .A1(n6400), .A2(n4921), .B1(n5744), .B2(n4920), .ZN(n4907)
         );
  AOI21_X1 U6107 ( .B1(n6397), .B2(n4923), .A(n4907), .ZN(n4908) );
  OAI211_X1 U6108 ( .C1(n6231), .C2(n6272), .A(n4909), .B(n4908), .ZN(U3052)
         );
  NAND2_X1 U6109 ( .A1(n4919), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4912) );
  OAI22_X1 U6110 ( .A1(n6412), .A2(n4921), .B1(n5754), .B2(n4920), .ZN(n4910)
         );
  AOI21_X1 U6111 ( .B1(n6409), .B2(n4923), .A(n4910), .ZN(n4911) );
  OAI211_X1 U6112 ( .C1(n6231), .C2(n6278), .A(n4912), .B(n4911), .ZN(U3054)
         );
  NAND2_X1 U6113 ( .A1(n4919), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4915) );
  OAI22_X1 U6114 ( .A1(n6430), .A2(n4921), .B1(n5769), .B2(n4920), .ZN(n4913)
         );
  AOI21_X1 U6115 ( .B1(n6426), .B2(n4923), .A(n4913), .ZN(n4914) );
  OAI211_X1 U6116 ( .C1(n6231), .C2(n6287), .A(n4915), .B(n4914), .ZN(U3057)
         );
  NAND2_X1 U6117 ( .A1(n4919), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4918) );
  OAI22_X1 U6118 ( .A1(n6436), .A2(n4921), .B1(n5774), .B2(n4920), .ZN(n4916)
         );
  AOI21_X1 U6119 ( .B1(n6432), .B2(n4923), .A(n4916), .ZN(n4917) );
  OAI211_X1 U6120 ( .C1(n6231), .C2(n6290), .A(n4918), .B(n4917), .ZN(U3058)
         );
  NAND2_X1 U6121 ( .A1(n4919), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4925) );
  OAI22_X1 U6122 ( .A1(n6424), .A2(n4921), .B1(n5764), .B2(n4920), .ZN(n4922)
         );
  AOI21_X1 U6123 ( .B1(n6420), .B2(n4923), .A(n4922), .ZN(n4924) );
  OAI211_X1 U6124 ( .C1(n6231), .C2(n6284), .A(n4925), .B(n4924), .ZN(U3056)
         );
  NAND2_X1 U6125 ( .A1(n4938), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4928) );
  OAI22_X1 U6126 ( .A1(n6400), .A2(n4940), .B1(n5744), .B2(n4939), .ZN(n4926)
         );
  AOI21_X1 U6127 ( .B1(n6397), .B2(n4942), .A(n4926), .ZN(n4927) );
  OAI211_X1 U6128 ( .C1(n4980), .C2(n6272), .A(n4928), .B(n4927), .ZN(U3020)
         );
  NAND2_X1 U6129 ( .A1(n4938), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4931) );
  OAI22_X1 U6130 ( .A1(n6424), .A2(n4940), .B1(n5764), .B2(n4939), .ZN(n4929)
         );
  AOI21_X1 U6131 ( .B1(n6420), .B2(n4942), .A(n4929), .ZN(n4930) );
  OAI211_X1 U6132 ( .C1(n4980), .C2(n6284), .A(n4931), .B(n4930), .ZN(U3024)
         );
  NAND2_X1 U6133 ( .A1(n4938), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4934) );
  OAI22_X1 U6134 ( .A1(n6412), .A2(n4940), .B1(n5754), .B2(n4939), .ZN(n4932)
         );
  AOI21_X1 U6135 ( .B1(n6409), .B2(n4942), .A(n4932), .ZN(n4933) );
  OAI211_X1 U6136 ( .C1(n4980), .C2(n6278), .A(n4934), .B(n4933), .ZN(U3022)
         );
  NAND2_X1 U6137 ( .A1(n4938), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4937) );
  OAI22_X1 U6138 ( .A1(n6436), .A2(n4940), .B1(n5774), .B2(n4939), .ZN(n4935)
         );
  AOI21_X1 U6139 ( .B1(n6432), .B2(n4942), .A(n4935), .ZN(n4936) );
  OAI211_X1 U6140 ( .C1(n4980), .C2(n6290), .A(n4937), .B(n4936), .ZN(U3026)
         );
  NAND2_X1 U6141 ( .A1(n4938), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4944) );
  OAI22_X1 U6142 ( .A1(n6430), .A2(n4940), .B1(n5769), .B2(n4939), .ZN(n4941)
         );
  AOI21_X1 U6143 ( .B1(n6426), .B2(n4942), .A(n4941), .ZN(n4943) );
  OAI211_X1 U6144 ( .C1(n4980), .C2(n6287), .A(n4944), .B(n4943), .ZN(U3025)
         );
  AOI21_X1 U6145 ( .B1(n4946), .B2(n4672), .A(n4945), .ZN(n5952) );
  INV_X1 U6146 ( .A(n5952), .ZN(n5038) );
  AOI22_X1 U6147 ( .A1(n6831), .A2(DATAI_9_), .B1(n6830), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4947) );
  OAI21_X1 U6148 ( .B1(n5038), .B2(n5418), .A(n4947), .ZN(U2882) );
  OAI22_X1 U6149 ( .A1(n6400), .A2(n4961), .B1(n5744), .B2(n4960), .ZN(n4948)
         );
  AOI21_X1 U6150 ( .B1(n6389), .B2(n4963), .A(n4948), .ZN(n4950) );
  NAND2_X1 U6151 ( .A1(n4964), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4949)
         );
  OAI211_X1 U6152 ( .C1(n4967), .C2(n5748), .A(n4950), .B(n4949), .ZN(U3132)
         );
  OAI22_X1 U6153 ( .A1(n6412), .A2(n4961), .B1(n5754), .B2(n4960), .ZN(n4951)
         );
  AOI21_X1 U6154 ( .B1(n6408), .B2(n4963), .A(n4951), .ZN(n4953) );
  NAND2_X1 U6155 ( .A1(n4964), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4952)
         );
  OAI211_X1 U6156 ( .C1(n4967), .C2(n5758), .A(n4953), .B(n4952), .ZN(U3134)
         );
  OAI22_X1 U6157 ( .A1(n6430), .A2(n4961), .B1(n5769), .B2(n4960), .ZN(n4954)
         );
  AOI21_X1 U6158 ( .B1(n6427), .B2(n4963), .A(n4954), .ZN(n4956) );
  NAND2_X1 U6159 ( .A1(n4964), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4955)
         );
  OAI211_X1 U6160 ( .C1(n4967), .C2(n5773), .A(n4956), .B(n4955), .ZN(U3137)
         );
  OAI22_X1 U6161 ( .A1(n6436), .A2(n4961), .B1(n5774), .B2(n4960), .ZN(n4957)
         );
  AOI21_X1 U6162 ( .B1(n6433), .B2(n4963), .A(n4957), .ZN(n4959) );
  NAND2_X1 U6163 ( .A1(n4964), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4958)
         );
  OAI211_X1 U6164 ( .C1(n4967), .C2(n5778), .A(n4959), .B(n4958), .ZN(U3138)
         );
  OAI22_X1 U6165 ( .A1(n6424), .A2(n4961), .B1(n5764), .B2(n4960), .ZN(n4962)
         );
  AOI21_X1 U6166 ( .B1(n6421), .B2(n4963), .A(n4962), .ZN(n4966) );
  NAND2_X1 U6167 ( .A1(n4964), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4965)
         );
  OAI211_X1 U6168 ( .C1(n4967), .C2(n5768), .A(n4966), .B(n4965), .ZN(U3136)
         );
  OAI21_X1 U6169 ( .B1(n3094), .B2(n4969), .A(n4968), .ZN(n4971) );
  INV_X1 U6170 ( .A(n4971), .ZN(n6122) );
  NAND2_X1 U6171 ( .A1(n6122), .A2(n6104), .ZN(n4976) );
  INV_X1 U6172 ( .A(REIP_REG_8__SCAN_IN), .ZN(n4972) );
  NOR2_X1 U6173 ( .A1(n6190), .A2(n4972), .ZN(n6118) );
  NOR2_X1 U6174 ( .A1(n6108), .A2(n4973), .ZN(n4974) );
  AOI211_X1 U6175 ( .C1(n6097), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6118), 
        .B(n4974), .ZN(n4975) );
  OAI211_X1 U6176 ( .C1(n5564), .C2(n4977), .A(n4976), .B(n4975), .ZN(U2978)
         );
  AOI21_X1 U6177 ( .B1(n4981), .B2(n6380), .A(n6331), .ZN(n4982) );
  NOR2_X1 U6178 ( .A1(n6451), .A2(n4983), .ZN(n5009) );
  AOI21_X1 U6179 ( .B1(n4978), .B2(n3102), .A(n5009), .ZN(n4985) );
  OAI22_X1 U6180 ( .A1(n4982), .A2(n4985), .B1(n4983), .B2(n6583), .ZN(n4979)
         );
  INV_X1 U6181 ( .A(n4982), .ZN(n4984) );
  AOI22_X1 U6182 ( .A1(n4985), .A2(n4984), .B1(n4983), .B2(n6393), .ZN(n4986)
         );
  NAND2_X1 U6183 ( .A1(n6306), .A2(n4986), .ZN(n5008) );
  AOI22_X1 U6184 ( .A1(n6413), .A2(n5009), .B1(INSTQUEUE_REG_1__3__SCAN_IN), 
        .B2(n5008), .ZN(n4987) );
  OAI21_X1 U6185 ( .B1(n6281), .B2(n6196), .A(n4987), .ZN(n4988) );
  AOI21_X1 U6186 ( .B1(n6414), .B2(n5012), .A(n4988), .ZN(n4989) );
  OAI21_X1 U6187 ( .B1(n5014), .B2(n6418), .A(n4989), .ZN(U3031) );
  AOI22_X1 U6188 ( .A1(n6438), .A2(n5009), .B1(INSTQUEUE_REG_1__7__SCAN_IN), 
        .B2(n5008), .ZN(n4990) );
  OAI21_X1 U6189 ( .B1(n6297), .B2(n6196), .A(n4990), .ZN(n4991) );
  AOI21_X1 U6190 ( .B1(n6442), .B2(n5012), .A(n4991), .ZN(n4992) );
  OAI21_X1 U6191 ( .B1(n5014), .B2(n6446), .A(n4992), .ZN(U3035) );
  AOI22_X1 U6192 ( .A1(n6431), .A2(n5009), .B1(INSTQUEUE_REG_1__6__SCAN_IN), 
        .B2(n5008), .ZN(n4993) );
  OAI21_X1 U6193 ( .B1(n6290), .B2(n6196), .A(n4993), .ZN(n4994) );
  AOI21_X1 U6194 ( .B1(n6432), .B2(n5012), .A(n4994), .ZN(n4995) );
  OAI21_X1 U6195 ( .B1(n5014), .B2(n6436), .A(n4995), .ZN(U3034) );
  AOI22_X1 U6196 ( .A1(n6401), .A2(n5009), .B1(INSTQUEUE_REG_1__1__SCAN_IN), 
        .B2(n5008), .ZN(n4996) );
  OAI21_X1 U6197 ( .B1(n6275), .B2(n6196), .A(n4996), .ZN(n4997) );
  AOI21_X1 U6198 ( .B1(n6402), .B2(n5012), .A(n4997), .ZN(n4998) );
  OAI21_X1 U6199 ( .B1(n5014), .B2(n6406), .A(n4998), .ZN(U3029) );
  AOI22_X1 U6200 ( .A1(n6419), .A2(n5009), .B1(INSTQUEUE_REG_1__4__SCAN_IN), 
        .B2(n5008), .ZN(n4999) );
  OAI21_X1 U6201 ( .B1(n6284), .B2(n6196), .A(n4999), .ZN(n5000) );
  AOI21_X1 U6202 ( .B1(n6420), .B2(n5012), .A(n5000), .ZN(n5001) );
  OAI21_X1 U6203 ( .B1(n5014), .B2(n6424), .A(n5001), .ZN(U3032) );
  AOI22_X1 U6204 ( .A1(n6425), .A2(n5009), .B1(INSTQUEUE_REG_1__5__SCAN_IN), 
        .B2(n5008), .ZN(n5002) );
  OAI21_X1 U6205 ( .B1(n6287), .B2(n6196), .A(n5002), .ZN(n5003) );
  AOI21_X1 U6206 ( .B1(n6426), .B2(n5012), .A(n5003), .ZN(n5004) );
  OAI21_X1 U6207 ( .B1(n5014), .B2(n6430), .A(n5004), .ZN(U3033) );
  AOI22_X1 U6208 ( .A1(n6407), .A2(n5009), .B1(INSTQUEUE_REG_1__2__SCAN_IN), 
        .B2(n5008), .ZN(n5005) );
  OAI21_X1 U6209 ( .B1(n6278), .B2(n6196), .A(n5005), .ZN(n5006) );
  AOI21_X1 U6210 ( .B1(n6409), .B2(n5012), .A(n5006), .ZN(n5007) );
  OAI21_X1 U6211 ( .B1(n5014), .B2(n6412), .A(n5007), .ZN(U3030) );
  AOI22_X1 U6212 ( .A1(n6388), .A2(n5009), .B1(INSTQUEUE_REG_1__0__SCAN_IN), 
        .B2(n5008), .ZN(n5010) );
  OAI21_X1 U6213 ( .B1(n6272), .B2(n6196), .A(n5010), .ZN(n5011) );
  AOI21_X1 U6214 ( .B1(n6397), .B2(n5012), .A(n5011), .ZN(n5013) );
  OAI21_X1 U6215 ( .B1(n5014), .B2(n6400), .A(n5013), .ZN(U3028) );
  NAND4_X1 U6216 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .A4(n5960), .ZN(n5288) );
  NOR2_X1 U6217 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5288), .ZN(n5949) );
  OAI21_X1 U6218 ( .B1(n5950), .B2(n5949), .A(REIP_REG_10__SCAN_IN), .ZN(n5019) );
  INV_X1 U6219 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5016) );
  AOI22_X1 U6220 ( .A1(EBX_REG_10__SCAN_IN), .A2(n5995), .B1(n5980), .B2(n6110), .ZN(n5015) );
  OAI211_X1 U6221 ( .C1(n6000), .C2(n5016), .A(n5015), .B(n5944), .ZN(n5017)
         );
  INV_X1 U6222 ( .A(n5017), .ZN(n5018) );
  OAI211_X1 U6223 ( .C1(n5993), .C2(n5559), .A(n5019), .B(n5018), .ZN(n5021)
         );
  INV_X1 U6224 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6522) );
  NOR3_X1 U6225 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6522), .A3(n5288), .ZN(n5020) );
  NOR2_X1 U6226 ( .A1(n5021), .A2(n5020), .ZN(n5022) );
  OAI21_X1 U6227 ( .B1(n5842), .B2(n5563), .A(n5022), .ZN(U2817) );
  INV_X1 U6228 ( .A(n5024), .ZN(n5025) );
  OR2_X1 U6229 ( .A1(n5026), .A2(n5025), .ZN(n5996) );
  NOR2_X1 U6230 ( .A1(n5027), .A2(n5996), .ZN(n5030) );
  OAI22_X1 U6231 ( .A1(n5969), .A2(n4102), .B1(n5028), .B2(n5947), .ZN(n5029)
         );
  AOI211_X1 U6232 ( .C1(n5921), .C2(REIP_REG_0__SCAN_IN), .A(n5030), .B(n5029), 
        .ZN(n5032) );
  OAI21_X1 U6233 ( .B1(n6006), .B2(n5990), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5031) );
  OAI211_X1 U6234 ( .C1(n6002), .C2(n5033), .A(n5032), .B(n5031), .ZN(U2827)
         );
  OR2_X1 U6235 ( .A1(n5035), .A2(n5034), .ZN(n5036) );
  NAND2_X1 U6236 ( .A1(n5037), .A2(n5036), .ZN(n5946) );
  INV_X1 U6237 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6872) );
  OAI222_X1 U6238 ( .A1(n5946), .A2(n5376), .B1(n6026), .B2(n6872), .C1(n3092), 
        .C2(n5038), .ZN(U2850) );
  AOI22_X1 U6239 ( .A1(n6165), .A2(n5980), .B1(n5995), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n5039) );
  OAI21_X1 U6240 ( .B1(n5040), .B2(n5996), .A(n5039), .ZN(n5043) );
  NOR2_X1 U6241 ( .A1(n5993), .A2(n5041), .ZN(n5042) );
  AOI211_X1 U6242 ( .C1(n5990), .C2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n5043), 
        .B(n5042), .ZN(n5049) );
  NAND2_X1 U6243 ( .A1(n5044), .A2(REIP_REG_2__SCAN_IN), .ZN(n5045) );
  NOR2_X1 U6244 ( .A1(n5983), .A2(REIP_REG_1__SCAN_IN), .ZN(n5994) );
  NOR2_X1 U6245 ( .A1(n5045), .A2(n5994), .ZN(n5301) );
  NOR2_X1 U6246 ( .A1(n4845), .A2(n6570), .ZN(n5047) );
  INV_X1 U6247 ( .A(n5045), .ZN(n5046) );
  AOI21_X1 U6248 ( .B1(n5047), .B2(n5046), .A(n5270), .ZN(n5979) );
  OAI21_X1 U6249 ( .B1(REIP_REG_3__SCAN_IN), .B2(n5301), .A(n5979), .ZN(n5048)
         );
  OAI211_X1 U6250 ( .C1(n6002), .C2(n5050), .A(n5049), .B(n5048), .ZN(U2824)
         );
  OAI21_X1 U6251 ( .B1(n5051), .B2(n5053), .A(n5052), .ZN(n5917) );
  AOI22_X1 U6252 ( .A1(n6831), .A2(DATAI_13_), .B1(n6830), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5054) );
  OAI21_X1 U6253 ( .B1(n5917), .B2(n5418), .A(n5054), .ZN(U2878) );
  NAND2_X1 U6254 ( .A1(n5222), .A2(n6074), .ZN(n5056) );
  OAI211_X1 U6255 ( .C1(n6869), .C2(n5548), .A(n5056), .B(n5055), .ZN(n5057)
         );
  AOI21_X1 U6256 ( .B1(n5217), .B2(n6101), .A(n5057), .ZN(n5058) );
  OAI21_X1 U6257 ( .B1(n5059), .B2(n6078), .A(n5058), .ZN(U2956) );
  XNOR2_X1 U6258 ( .A(n5557), .B(n6871), .ZN(n5493) );
  AND2_X2 U6259 ( .A1(n5459), .A2(n5061), .ZN(n5487) );
  NOR2_X1 U6260 ( .A1(n5716), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5483)
         );
  NAND2_X1 U6261 ( .A1(n5716), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5484) );
  OAI21_X2 U6262 ( .B1(n5487), .B2(n5483), .A(n5484), .ZN(n5478) );
  XNOR2_X1 U6263 ( .A(n5557), .B(n6760), .ZN(n5479) );
  NOR2_X1 U6264 ( .A1(n5557), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5469)
         );
  NAND2_X1 U6265 ( .A1(n5477), .A2(n5469), .ZN(n5463) );
  INV_X1 U6266 ( .A(n5463), .ZN(n5063) );
  INV_X1 U6267 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5062) );
  NAND2_X1 U6268 ( .A1(n5063), .A2(n5062), .ZN(n5065) );
  NAND2_X1 U6269 ( .A1(n5470), .A2(n3189), .ZN(n5064) );
  AOI21_X1 U6270 ( .B1(n5068), .B2(n5334), .A(n5067), .ZN(n5812) );
  AND2_X1 U6271 ( .A1(n6156), .A2(REIP_REG_24__SCAN_IN), .ZN(n5074) );
  AOI21_X1 U6272 ( .B1(n5623), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5069) );
  NOR2_X1 U6273 ( .A1(n5610), .A2(n5069), .ZN(n5070) );
  AOI211_X1 U6274 ( .C1(n6174), .C2(n5812), .A(n5074), .B(n5070), .ZN(n5071)
         );
  OAI21_X1 U6275 ( .B1(n5080), .B2(n6184), .A(n5071), .ZN(U2994) );
  NOR2_X1 U6276 ( .A1(n5548), .A2(n5072), .ZN(n5073) );
  AOI211_X1 U6277 ( .C1(n6074), .C2(n5810), .A(n5074), .B(n5073), .ZN(n5079)
         );
  OAI21_X1 U6278 ( .B1(n5075), .B2(n5077), .A(n5076), .ZN(n5391) );
  INV_X1 U6279 ( .A(n5391), .ZN(n5813) );
  NAND2_X1 U6280 ( .A1(n5813), .A2(n6101), .ZN(n5078) );
  OAI211_X1 U6281 ( .C1(n5080), .C2(n6078), .A(n5079), .B(n5078), .ZN(U2962)
         );
  INV_X1 U6282 ( .A(n5082), .ZN(n5083) );
  NOR2_X1 U6283 ( .A1(n5084), .A2(n5083), .ZN(n5085) );
  XNOR2_X1 U6284 ( .A(n5081), .B(n5085), .ZN(n5101) );
  INV_X1 U6285 ( .A(n5086), .ZN(n6136) );
  OAI22_X1 U6286 ( .A1(n5088), .A2(n5641), .B1(n6136), .B2(n5087), .ZN(n5089)
         );
  NOR2_X1 U6287 ( .A1(n5090), .A2(n5089), .ZN(n6131) );
  OAI21_X1 U6288 ( .B1(n5679), .B2(n6120), .A(n6131), .ZN(n6111) );
  OAI22_X1 U6289 ( .A1(n6127), .A2(n5946), .B1(n6522), .B2(n6190), .ZN(n5091)
         );
  AOI21_X1 U6290 ( .B1(n6111), .B2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n5091), 
        .ZN(n5096) );
  NOR2_X1 U6291 ( .A1(n6181), .A2(n6180), .ZN(n6135) );
  OAI21_X1 U6292 ( .B1(n6178), .B2(n6135), .A(n5092), .ZN(n6166) );
  NOR2_X1 U6293 ( .A1(n6138), .A2(n6166), .ZN(n6140) );
  NAND2_X1 U6294 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6140), .ZN(n6133)
         );
  NOR2_X1 U6295 ( .A1(n5093), .A2(n6133), .ZN(n6114) );
  NAND2_X1 U6296 ( .A1(n6114), .A2(n5094), .ZN(n5095) );
  OAI211_X1 U6297 ( .C1(n5101), .C2(n6184), .A(n5096), .B(n5095), .ZN(U3009)
         );
  INV_X1 U6298 ( .A(n5951), .ZN(n5098) );
  AOI22_X1 U6299 ( .A1(n6097), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .B1(n6156), 
        .B2(REIP_REG_9__SCAN_IN), .ZN(n5097) );
  OAI21_X1 U6300 ( .B1(n6108), .B2(n5098), .A(n5097), .ZN(n5099) );
  AOI21_X1 U6301 ( .B1(n5952), .B2(n6101), .A(n5099), .ZN(n5100) );
  OAI21_X1 U6302 ( .B1(n5101), .B2(n6078), .A(n5100), .ZN(U2977) );
  OAI22_X1 U6303 ( .A1(n6449), .A2(n6485), .B1(n6561), .B2(n6753), .ZN(n5883)
         );
  AOI21_X1 U6304 ( .B1(n6452), .B2(n5881), .A(n5164), .ZN(n5108) );
  NAND2_X1 U6305 ( .A1(n3102), .A2(n5171), .ZN(n5104) );
  NAND2_X1 U6306 ( .A1(n5167), .A2(n5107), .ZN(n5103) );
  NAND2_X1 U6307 ( .A1(n5104), .A2(n5103), .ZN(n6450) );
  OAI22_X1 U6308 ( .A1(n6858), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6564), .ZN(n5105) );
  AOI21_X1 U6309 ( .B1(n6450), .B2(n5881), .A(n5105), .ZN(n5106) );
  OAI22_X1 U6310 ( .A1(n5108), .A2(n5107), .B1(n5164), .B2(n5106), .ZN(U3461)
         );
  INV_X1 U6311 ( .A(n4534), .ZN(n5165) );
  AOI21_X1 U6312 ( .B1(n6477), .B2(n5165), .A(n5164), .ZN(n5115) );
  INV_X1 U6313 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5568) );
  AOI22_X1 U6314 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5568), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6180), .ZN(n5173) );
  NOR2_X1 U6315 ( .A1(n6858), .A2(n5109), .ZN(n5174) );
  INV_X1 U6316 ( .A(n5174), .ZN(n5111) );
  NAND3_X1 U6317 ( .A1(n4534), .A2(n6477), .A3(n4048), .ZN(n5110) );
  OAI21_X1 U6318 ( .B1(n5173), .B2(n5111), .A(n5110), .ZN(n5112) );
  AOI21_X1 U6319 ( .B1(n5113), .B2(n5881), .A(n5112), .ZN(n5114) );
  OAI22_X1 U6320 ( .A1(n5115), .A2(n4048), .B1(n5164), .B2(n5114), .ZN(U3459)
         );
  NAND3_X1 U6321 ( .A1(n5444), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5557), .ZN(n5117) );
  INV_X1 U6322 ( .A(n5116), .ZN(n5452) );
  NAND3_X1 U6323 ( .A1(n5452), .A2(n5443), .A3(n6731), .ZN(n5434) );
  INV_X1 U6324 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5605) );
  AOI22_X1 U6325 ( .A1(n5117), .A2(n5434), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5605), .ZN(n5118) );
  XNOR2_X1 U6326 ( .A(n5118), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5591)
         );
  NAND2_X1 U6327 ( .A1(n6156), .A2(REIP_REG_28__SCAN_IN), .ZN(n5586) );
  OAI21_X1 U6328 ( .B1(n5548), .B2(n5119), .A(n5586), .ZN(n5124) );
  NAND2_X2 U6329 ( .A1(n5122), .A2(n5121), .ZN(n5143) );
  NOR2_X1 U6330 ( .A1(n5143), .A2(n5564), .ZN(n5123) );
  OAI21_X1 U6331 ( .B1(n5591), .B2(n6078), .A(n5125), .ZN(U2958) );
  INV_X1 U6332 ( .A(n5798), .ZN(n5211) );
  INV_X1 U6333 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6548) );
  NOR2_X1 U6334 ( .A1(n6548), .A2(REIP_REG_28__SCAN_IN), .ZN(n5137) );
  INV_X1 U6335 ( .A(n5313), .ZN(n5127) );
  AOI21_X1 U6336 ( .B1(n5127), .B2(n5311), .A(n5126), .ZN(n5129) );
  OR2_X1 U6337 ( .A1(n5129), .A2(n5128), .ZN(n5587) );
  INV_X1 U6338 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5144) );
  NAND2_X1 U6339 ( .A1(n5990), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5130)
         );
  OAI21_X1 U6340 ( .B1(n5144), .B2(n5969), .A(n5130), .ZN(n5131) );
  AOI21_X1 U6341 ( .B1(n6006), .B2(n5132), .A(n5131), .ZN(n5135) );
  INV_X1 U6342 ( .A(REIP_REG_28__SCAN_IN), .ZN(n5133) );
  OR2_X1 U6343 ( .A1(n5197), .A2(n5133), .ZN(n5134) );
  OAI211_X1 U6344 ( .C1(n5587), .C2(n5947), .A(n5135), .B(n5134), .ZN(n5136)
         );
  AOI21_X1 U6345 ( .B1(n5211), .B2(n5137), .A(n5136), .ZN(n5138) );
  OAI21_X1 U6346 ( .B1(n5143), .B2(n5842), .A(n5138), .ZN(U2799) );
  NOR2_X2 U6347 ( .A1(n5140), .A2(n5139), .ZN(n6030) );
  AOI22_X1 U6348 ( .A1(n6030), .A2(DATAI_12_), .B1(n6830), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5142) );
  NOR2_X2 U6349 ( .A1(n6830), .A2(n3404), .ZN(n6028) );
  NAND2_X1 U6350 ( .A1(n6028), .A2(DATAI_28_), .ZN(n5141) );
  OAI211_X1 U6351 ( .C1(n5143), .C2(n5418), .A(n5142), .B(n5141), .ZN(U2863)
         );
  OAI222_X1 U6352 ( .A1(n5144), .A2(n6026), .B1(n5376), .B2(n5587), .C1(n5143), 
        .C2(n3092), .ZN(U2831) );
  NOR3_X1 U6353 ( .A1(n5145), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5146) );
  AOI22_X1 U6354 ( .A1(n5425), .A2(n5566), .B1(n5453), .B2(n5146), .ZN(n5147)
         );
  XNOR2_X1 U6355 ( .A(n5147), .B(n5568), .ZN(n5574) );
  AOI22_X1 U6356 ( .A1(n3952), .A2(EAX_REG_31__SCAN_IN), .B1(n5150), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5151) );
  INV_X1 U6357 ( .A(n5151), .ZN(n5152) );
  INV_X1 U6358 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6876) );
  NOR2_X1 U6359 ( .A1(n6190), .A2(n6876), .ZN(n5571) );
  AOI21_X1 U6360 ( .B1(n6097), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5571), 
        .ZN(n5154) );
  OAI21_X1 U6361 ( .B1(n5155), .B2(n6108), .A(n5154), .ZN(n5156) );
  AOI21_X1 U6362 ( .B1(n5196), .B2(n6101), .A(n5156), .ZN(n5157) );
  OAI21_X1 U6363 ( .B1(n5574), .B2(n6078), .A(n5157), .ZN(U2955) );
  NAND3_X1 U6364 ( .A1(n5196), .A2(n3250), .A3(n5419), .ZN(n5159) );
  AOI22_X1 U6365 ( .A1(n6028), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6830), .ZN(n5158) );
  NAND2_X1 U6366 ( .A1(n5159), .A2(n5158), .ZN(U2860) );
  AOI22_X1 U6367 ( .A1(n6030), .A2(DATAI_13_), .B1(n6830), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5161) );
  NAND2_X1 U6368 ( .A1(n6028), .A2(DATAI_29_), .ZN(n5160) );
  OAI211_X1 U6369 ( .C1(n5163), .C2(n5418), .A(n5161), .B(n5160), .ZN(U2862)
         );
  OAI222_X1 U6370 ( .A1(n3092), .A2(n5163), .B1(n6026), .B2(n5162), .C1(n5575), 
        .C2(n5376), .ZN(U2830) );
  INV_X1 U6371 ( .A(n5164), .ZN(n6568) );
  NAND2_X1 U6372 ( .A1(n6452), .A2(n3195), .ZN(n5169) );
  INV_X1 U6373 ( .A(n4571), .ZN(n5166) );
  NAND3_X1 U6374 ( .A1(n5167), .A2(n5166), .A3(n5165), .ZN(n5168) );
  NAND2_X1 U6375 ( .A1(n5169), .A2(n5168), .ZN(n5170) );
  AOI21_X1 U6376 ( .B1(n4580), .B2(n5171), .A(n5170), .ZN(n6448) );
  INV_X1 U6377 ( .A(n5881), .ZN(n6566) );
  AOI22_X1 U6378 ( .A1(n5174), .A2(n5173), .B1(n5172), .B2(n6477), .ZN(n5175)
         );
  OAI21_X1 U6379 ( .B1(n6448), .B2(n6566), .A(n5175), .ZN(n5177) );
  AOI22_X1 U6380 ( .A1(n6568), .A2(n5177), .B1(n5176), .B2(n6477), .ZN(n5178)
         );
  OAI21_X1 U6381 ( .B1(n3195), .B2(n6568), .A(n5178), .ZN(U3460) );
  INV_X1 U6382 ( .A(n4348), .ZN(n5190) );
  NAND2_X1 U6383 ( .A1(n5179), .A2(n5190), .ZN(n5182) );
  NOR2_X1 U6384 ( .A1(n5189), .A2(n5180), .ZN(n5181) );
  AOI21_X1 U6385 ( .B1(n5188), .B2(n5182), .A(n5181), .ZN(n5186) );
  INV_X1 U6386 ( .A(n5183), .ZN(n5184) );
  OR2_X1 U6387 ( .A1(n5188), .A2(n5184), .ZN(n5185) );
  AND2_X1 U6388 ( .A1(n5186), .A2(n5185), .ZN(n6466) );
  INV_X1 U6389 ( .A(n6466), .ZN(n5195) );
  NAND2_X1 U6390 ( .A1(n5188), .A2(n5187), .ZN(n5193) );
  NAND2_X1 U6391 ( .A1(n5189), .A2(n3096), .ZN(n5191) );
  NAND2_X1 U6392 ( .A1(n5191), .A2(n5190), .ZN(n5192) );
  NAND2_X1 U6393 ( .A1(n5193), .A2(n5192), .ZN(n5887) );
  AOI21_X1 U6394 ( .B1(n5194), .B2(n6503), .A(READY_N), .ZN(n6581) );
  OR2_X1 U6395 ( .A1(n5887), .A2(n6581), .ZN(n6468) );
  AND2_X1 U6396 ( .A1(n6468), .A2(n6481), .ZN(n5892) );
  MUX2_X1 U6397 ( .A(MORE_REG_SCAN_IN), .B(n5195), .S(n5892), .Z(U3471) );
  INV_X1 U6398 ( .A(n5196), .ZN(n5216) );
  AND2_X1 U6399 ( .A1(n5198), .A2(n5197), .ZN(n5218) );
  OAI21_X1 U6400 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5983), .A(n5218), .ZN(n5214) );
  OAI211_X1 U6401 ( .C1(n5202), .C2(n5201), .A(n5200), .B(n5199), .ZN(n5206)
         );
  OAI22_X1 U6402 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n5203), .ZN(n5205) );
  XNOR2_X1 U6403 ( .A(n5206), .B(n5205), .ZN(n5565) );
  AOI22_X1 U6404 ( .A1(n5990), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .B1(n5208), 
        .B2(n5207), .ZN(n5209) );
  OAI21_X1 U6405 ( .B1(n5565), .B2(n5947), .A(n5209), .ZN(n5213) );
  NAND3_X1 U6406 ( .A1(n5211), .A2(REIP_REG_29__SCAN_IN), .A3(n5210), .ZN(
        n5223) );
  INV_X1 U6407 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6556) );
  NOR3_X1 U6408 ( .A1(n5223), .A2(REIP_REG_31__SCAN_IN), .A3(n6556), .ZN(n5212) );
  AOI211_X1 U6409 ( .C1(REIP_REG_31__SCAN_IN), .C2(n5214), .A(n5213), .B(n5212), .ZN(n5215) );
  OAI21_X1 U6410 ( .B1(n5216), .B2(n5842), .A(n5215), .ZN(U2796) );
  INV_X1 U6411 ( .A(n5218), .ZN(n5225) );
  OAI22_X1 U6412 ( .A1(n6000), .A2(n6869), .B1(n5219), .B2(n5969), .ZN(n5221)
         );
  AOI21_X1 U6413 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5225), .A(n5224), .ZN(n5226) );
  OAI21_X1 U6414 ( .B1(n5380), .B2(n5842), .A(n5226), .ZN(U2797) );
  AOI21_X1 U6415 ( .B1(n5228), .B2(n5319), .A(n5227), .ZN(n5450) );
  INV_X1 U6416 ( .A(n5450), .ZN(n5385) );
  INV_X1 U6417 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6877) );
  OAI22_X1 U6418 ( .A1(n6877), .A2(n5969), .B1(n5448), .B2(n6000), .ZN(n5232)
         );
  NAND2_X1 U6419 ( .A1(n5323), .A2(n5229), .ZN(n5230) );
  NAND2_X1 U6420 ( .A1(n5313), .A2(n5230), .ZN(n5599) );
  NOR2_X1 U6421 ( .A1(n5599), .A2(n5947), .ZN(n5231) );
  AOI211_X1 U6422 ( .C1(n6006), .C2(n5446), .A(n5232), .B(n5231), .ZN(n5235)
         );
  INV_X1 U6423 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6544) );
  NAND2_X1 U6424 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5805), .ZN(n5799) );
  INV_X1 U6425 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6546) );
  OAI21_X1 U6426 ( .B1(n6544), .B2(n5799), .A(n6546), .ZN(n5233) );
  NAND2_X1 U6427 ( .A1(n5233), .A2(n5792), .ZN(n5234) );
  OAI211_X1 U6428 ( .C1(n5385), .C2(n5842), .A(n5235), .B(n5234), .ZN(U2801)
         );
  OR2_X1 U6429 ( .A1(n5337), .A2(n5237), .ZN(n5329) );
  INV_X1 U6430 ( .A(n5329), .ZN(n5236) );
  AOI21_X1 U6431 ( .B1(n5237), .B2(n5337), .A(n5236), .ZN(n5474) );
  INV_X1 U6432 ( .A(n5474), .ZN(n5396) );
  INV_X1 U6433 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6875) );
  INV_X1 U6434 ( .A(n5838), .ZN(n5828) );
  OAI21_X1 U6435 ( .B1(REIP_REG_21__SCAN_IN), .B2(n5827), .A(n5828), .ZN(n5239) );
  NAND2_X1 U6436 ( .A1(STATE2_REG_3__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6837) );
  INV_X1 U6437 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5336) );
  OAI22_X1 U6438 ( .A1(n5998), .A2(n6837), .B1(n5336), .B2(n5969), .ZN(n5238)
         );
  AOI221_X1 U6439 ( .B1(n5240), .B2(n6875), .C1(n5239), .C2(
        REIP_REG_22__SCAN_IN), .A(n5238), .ZN(n5245) );
  AOI21_X1 U6440 ( .B1(n3120), .B2(n5340), .A(n5241), .ZN(n5242) );
  OR2_X1 U6441 ( .A1(n5242), .A2(n5332), .ZN(n5626) );
  NOR2_X1 U6442 ( .A1(n5626), .A2(n5947), .ZN(n5243) );
  AOI21_X1 U6443 ( .B1(n6006), .B2(n5473), .A(n5243), .ZN(n5244) );
  OAI211_X1 U6444 ( .C1(n5396), .C2(n5842), .A(n5245), .B(n5244), .ZN(U2805)
         );
  OR2_X1 U6445 ( .A1(n5359), .A2(n5246), .ZN(n5352) );
  NAND2_X1 U6446 ( .A1(n5359), .A2(n5246), .ZN(n5247) );
  NAND2_X1 U6447 ( .A1(n5352), .A2(n5247), .ZN(n5508) );
  INV_X1 U6448 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6535) );
  NAND2_X1 U6449 ( .A1(n5921), .A2(n5248), .ZN(n5909) );
  AOI21_X1 U6450 ( .B1(n5990), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5984), 
        .ZN(n5249) );
  OAI221_X1 U6451 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5850), .C1(n6535), .C2(
        n5909), .A(n5249), .ZN(n5256) );
  OR2_X1 U6452 ( .A1(n5251), .A2(n5250), .ZN(n5252) );
  NAND2_X1 U6453 ( .A1(n5364), .A2(n5252), .ZN(n5355) );
  OR2_X1 U6454 ( .A1(n5364), .A2(n5252), .ZN(n5253) );
  AND2_X1 U6455 ( .A1(n5355), .A2(n5253), .ZN(n5661) );
  AOI22_X1 U6456 ( .A1(n5661), .A2(n5980), .B1(EBX_REG_18__SCAN_IN), .B2(n5995), .ZN(n5254) );
  OAI21_X1 U6457 ( .B1(n5993), .B2(n5504), .A(n5254), .ZN(n5255) );
  NOR2_X1 U6458 ( .A1(n5256), .A2(n5255), .ZN(n5257) );
  OAI21_X1 U6459 ( .B1(n5508), .B2(n5842), .A(n5257), .ZN(U2809) );
  INV_X1 U6460 ( .A(n5259), .ZN(n5260) );
  OAI21_X1 U6461 ( .B1(n5258), .B2(n5261), .A(n5260), .ZN(n5524) );
  INV_X1 U6462 ( .A(n5262), .ZN(n5521) );
  INV_X1 U6463 ( .A(n5263), .ZN(n5293) );
  AOI21_X1 U6464 ( .B1(n5293), .B2(n5278), .A(n5264), .ZN(n5266) );
  INV_X1 U6465 ( .A(n5362), .ZN(n5265) );
  NOR2_X1 U6466 ( .A1(n5266), .A2(n5265), .ZN(n5860) );
  AOI21_X1 U6467 ( .B1(n5860), .B2(n5980), .A(n5984), .ZN(n5267) );
  OAI21_X1 U6468 ( .B1(n6000), .B2(n5519), .A(n5267), .ZN(n5274) );
  OAI21_X1 U6469 ( .B1(REIP_REG_16__SCAN_IN), .B2(REIP_REG_15__SCAN_IN), .A(
        n5268), .ZN(n5272) );
  NOR2_X1 U6470 ( .A1(n5270), .A2(n5269), .ZN(n5289) );
  AOI22_X1 U6471 ( .A1(EBX_REG_16__SCAN_IN), .A2(n5995), .B1(
        REIP_REG_16__SCAN_IN), .B2(n5289), .ZN(n5271) );
  OAI21_X1 U6472 ( .B1(n5281), .B2(n5272), .A(n5271), .ZN(n5273) );
  AOI211_X1 U6473 ( .C1(n6006), .C2(n5521), .A(n5274), .B(n5273), .ZN(n5275)
         );
  OAI21_X1 U6474 ( .B1(n5524), .B2(n5842), .A(n5275), .ZN(U2811) );
  AND2_X1 U6475 ( .A1(n5287), .A2(n5276), .ZN(n5277) );
  NOR2_X1 U6476 ( .A1(n5258), .A2(n5277), .ZN(n5533) );
  INV_X1 U6477 ( .A(n5533), .ZN(n5409) );
  XNOR2_X1 U6478 ( .A(n5293), .B(n5278), .ZN(n5683) );
  NAND2_X1 U6479 ( .A1(n5990), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5279)
         );
  OAI211_X1 U6480 ( .C1(n5683), .C2(n5947), .A(n5279), .B(n5944), .ZN(n5283)
         );
  AOI22_X1 U6481 ( .A1(EBX_REG_15__SCAN_IN), .A2(n5995), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5289), .ZN(n5280) );
  OAI21_X1 U6482 ( .B1(REIP_REG_15__SCAN_IN), .B2(n5281), .A(n5280), .ZN(n5282) );
  AOI211_X1 U6483 ( .C1(n5530), .C2(n6006), .A(n5283), .B(n5282), .ZN(n5284)
         );
  OAI21_X1 U6484 ( .B1(n5409), .B2(n5842), .A(n5284), .ZN(U2812) );
  NAND2_X1 U6485 ( .A1(n5052), .A2(n5285), .ZN(n5286) );
  NAND2_X1 U6486 ( .A1(n5287), .A2(n5286), .ZN(n5543) );
  INV_X1 U6487 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6527) );
  INV_X1 U6488 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6521) );
  NOR3_X1 U6489 ( .A1(n6521), .A2(n6522), .A3(n5288), .ZN(n5936) );
  NAND2_X1 U6490 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5936), .ZN(n5935) );
  NOR2_X1 U6491 ( .A1(n6527), .A2(n5935), .ZN(n5926) );
  OAI221_X1 U6492 ( .B1(REIP_REG_14__SCAN_IN), .B2(REIP_REG_13__SCAN_IN), .C1(
        REIP_REG_14__SCAN_IN), .C2(n5926), .A(n5289), .ZN(n5297) );
  INV_X1 U6493 ( .A(n5290), .ZN(n5540) );
  AOI21_X1 U6494 ( .B1(n5699), .B2(n5691), .A(n5291), .ZN(n5292) );
  NOR2_X1 U6495 ( .A1(n5293), .A2(n5292), .ZN(n5869) );
  AOI22_X1 U6496 ( .A1(EBX_REG_14__SCAN_IN), .A2(n5995), .B1(n5980), .B2(n5869), .ZN(n5294) );
  OAI21_X1 U6497 ( .B1(n5538), .B2(n6000), .A(n5294), .ZN(n5295) );
  AOI211_X1 U6498 ( .C1(n6006), .C2(n5540), .A(n5984), .B(n5295), .ZN(n5296)
         );
  OAI211_X1 U6499 ( .C1(n5543), .C2(n5842), .A(n5297), .B(n5296), .ZN(U2813)
         );
  INV_X1 U6500 ( .A(n6002), .ZN(n5973) );
  NAND2_X1 U6501 ( .A1(n5973), .A2(n6102), .ZN(n5306) );
  INV_X1 U6502 ( .A(n4523), .ZN(n5299) );
  AOI22_X1 U6503 ( .A1(n6173), .A2(n5980), .B1(n5995), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n5298) );
  OAI21_X1 U6504 ( .B1(n5299), .B2(n5996), .A(n5298), .ZN(n5304) );
  INV_X1 U6505 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6698) );
  NAND2_X1 U6506 ( .A1(n5300), .A2(REIP_REG_1__SCAN_IN), .ZN(n5302) );
  AOI21_X1 U6507 ( .B1(n6698), .B2(n5302), .A(n5301), .ZN(n5303) );
  AOI211_X1 U6508 ( .C1(n5990), .C2(PHYADDRPOINTER_REG_2__SCAN_IN), .A(n5304), 
        .B(n5303), .ZN(n5305) );
  OAI211_X1 U6509 ( .C1(n6107), .C2(n5993), .A(n5306), .B(n5305), .ZN(U2825)
         );
  OAI22_X1 U6510 ( .A1(n5565), .A2(n5376), .B1(n5307), .B2(n6026), .ZN(U2828)
         );
  NOR2_X1 U6511 ( .A1(n5227), .A2(n5308), .ZN(n5309) );
  INV_X1 U6512 ( .A(n5311), .ZN(n5312) );
  XNOR2_X1 U6513 ( .A(n5313), .B(n5312), .ZN(n5793) );
  INV_X1 U6514 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5314) );
  OAI222_X1 U6515 ( .A1(n3092), .A2(n5794), .B1(n5376), .B2(n5793), .C1(n5314), 
        .C2(n6026), .ZN(U2832) );
  OAI22_X1 U6516 ( .A1(n5599), .A2(n5376), .B1(n6877), .B2(n6026), .ZN(n5315)
         );
  INV_X1 U6517 ( .A(n5315), .ZN(n5316) );
  OAI21_X1 U6518 ( .B1(n5385), .B2(n3092), .A(n5316), .ZN(U2833) );
  NAND2_X1 U6519 ( .A1(n5076), .A2(n5317), .ZN(n5318) );
  NAND2_X1 U6520 ( .A1(n5321), .A2(n5320), .ZN(n5322) );
  NAND2_X1 U6521 ( .A1(n5323), .A2(n5322), .ZN(n5809) );
  OAI22_X1 U6522 ( .A1(n5809), .A2(n5376), .B1(n5324), .B2(n6026), .ZN(n5325)
         );
  INV_X1 U6523 ( .A(n5325), .ZN(n5326) );
  OAI21_X1 U6524 ( .B1(n5388), .B2(n3092), .A(n5326), .ZN(U2834) );
  AOI22_X1 U6525 ( .A1(n5812), .A2(n6022), .B1(EBX_REG_24__SCAN_IN), .B2(n5368), .ZN(n5327) );
  OAI21_X1 U6526 ( .B1(n5391), .B2(n3092), .A(n5327), .ZN(U2835) );
  AND2_X1 U6527 ( .A1(n5329), .A2(n5328), .ZN(n5330) );
  NOR2_X1 U6528 ( .A1(n5075), .A2(n5330), .ZN(n5467) );
  INV_X1 U6529 ( .A(n5467), .ZN(n5821) );
  INV_X1 U6530 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5335) );
  OR2_X1 U6531 ( .A1(n5332), .A2(n5331), .ZN(n5333) );
  AND2_X1 U6532 ( .A1(n5334), .A2(n5333), .ZN(n5619) );
  INV_X1 U6533 ( .A(n5619), .ZN(n5820) );
  OAI222_X1 U6534 ( .A1(n3092), .A2(n5821), .B1(n6026), .B2(n5335), .C1(n5820), 
        .C2(n5376), .ZN(U2836) );
  OAI222_X1 U6535 ( .A1(n3092), .A2(n5396), .B1(n6026), .B2(n5336), .C1(n5626), 
        .C2(n5376), .ZN(U2837) );
  INV_X1 U6536 ( .A(n5337), .ZN(n5338) );
  AOI21_X1 U6537 ( .B1(n5339), .B2(n5344), .A(n5338), .ZN(n5834) );
  INV_X1 U6538 ( .A(n5834), .ZN(n5399) );
  INV_X1 U6539 ( .A(n5340), .ZN(n5341) );
  XNOR2_X1 U6540 ( .A(n5342), .B(n5341), .ZN(n5832) );
  INV_X1 U6541 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5343) );
  OAI222_X1 U6542 ( .A1(n3092), .A2(n5399), .B1(n5376), .B2(n5832), .C1(n5343), 
        .C2(n6026), .ZN(U2838) );
  OAI21_X1 U6543 ( .B1(n5353), .B2(n5345), .A(n5344), .ZN(n5843) );
  INV_X1 U6544 ( .A(n5346), .ZN(n5348) );
  MUX2_X1 U6545 ( .A(n4189), .B(n5348), .S(n5347), .Z(n5350) );
  XNOR2_X1 U6546 ( .A(n5350), .B(n5349), .ZN(n5847) );
  OAI222_X1 U6547 ( .A1(n5843), .A2(n3092), .B1(n5376), .B2(n5847), .C1(n6026), 
        .C2(n4156), .ZN(U2839) );
  AND2_X1 U6548 ( .A1(n5352), .A2(n5351), .ZN(n5354) );
  OR2_X1 U6549 ( .A1(n5354), .A2(n5353), .ZN(n5852) );
  XNOR2_X1 U6550 ( .A(n5355), .B(n3115), .ZN(n5853) );
  OAI22_X1 U6551 ( .A1(n5853), .A2(n5376), .B1(n5859), .B2(n6026), .ZN(n5356)
         );
  INV_X1 U6552 ( .A(n5356), .ZN(n5357) );
  OAI21_X1 U6553 ( .B1(n5852), .B2(n3092), .A(n5357), .ZN(U2840) );
  AOI22_X1 U6554 ( .A1(n5661), .A2(n6022), .B1(EBX_REG_18__SCAN_IN), .B2(n5368), .ZN(n5358) );
  OAI21_X1 U6555 ( .B1(n5508), .B2(n3092), .A(n5358), .ZN(U2841) );
  OAI21_X1 U6556 ( .B1(n5259), .B2(n5360), .A(n5359), .ZN(n5912) );
  AND2_X1 U6557 ( .A1(n5362), .A2(n5361), .ZN(n5363) );
  NOR2_X1 U6558 ( .A1(n5364), .A2(n5363), .ZN(n5913) );
  AOI22_X1 U6559 ( .A1(n5913), .A2(n6022), .B1(EBX_REG_17__SCAN_IN), .B2(n5368), .ZN(n5365) );
  OAI21_X1 U6560 ( .B1(n5912), .B2(n3092), .A(n5365), .ZN(U2842) );
  AOI22_X1 U6561 ( .A1(n5860), .A2(n6022), .B1(EBX_REG_16__SCAN_IN), .B2(n5368), .ZN(n5366) );
  OAI21_X1 U6562 ( .B1(n5524), .B2(n3092), .A(n5366), .ZN(U2843) );
  OAI222_X1 U6563 ( .A1(n5409), .A2(n3092), .B1(n5376), .B2(n5683), .C1(n5367), 
        .C2(n6026), .ZN(U2844) );
  AOI22_X1 U6564 ( .A1(n5869), .A2(n6022), .B1(EBX_REG_14__SCAN_IN), .B2(n5368), .ZN(n5369) );
  OAI21_X1 U6565 ( .B1(n5543), .B2(n3092), .A(n5369), .ZN(U2845) );
  AND2_X1 U6566 ( .A1(n5371), .A2(n5370), .ZN(n5372) );
  NOR2_X1 U6567 ( .A1(n5412), .A2(n5372), .ZN(n6075) );
  INV_X1 U6568 ( .A(n6075), .ZN(n5417) );
  INV_X1 U6569 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U6570 ( .A1(n5374), .A2(n5373), .ZN(n5375) );
  NAND2_X1 U6571 ( .A1(n5700), .A2(n5375), .ZN(n5937) );
  OAI222_X1 U6572 ( .A1(n5417), .A2(n3092), .B1(n6026), .B2(n5377), .C1(n5937), 
        .C2(n5376), .ZN(U2848) );
  AOI22_X1 U6573 ( .A1(n6030), .A2(DATAI_14_), .B1(n6830), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U6574 ( .A1(n6028), .A2(DATAI_30_), .ZN(n5378) );
  OAI211_X1 U6575 ( .C1(n5380), .C2(n5418), .A(n5379), .B(n5378), .ZN(U2861)
         );
  AOI22_X1 U6576 ( .A1(n6030), .A2(DATAI_11_), .B1(n6830), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U6577 ( .A1(n6028), .A2(DATAI_27_), .ZN(n5381) );
  OAI211_X1 U6578 ( .C1(n5794), .C2(n5418), .A(n5382), .B(n5381), .ZN(U2864)
         );
  AOI22_X1 U6579 ( .A1(n6030), .A2(DATAI_10_), .B1(n6830), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U6580 ( .A1(n6028), .A2(DATAI_26_), .ZN(n5383) );
  OAI211_X1 U6581 ( .C1(n5385), .C2(n5418), .A(n5384), .B(n5383), .ZN(U2865)
         );
  AOI22_X1 U6582 ( .A1(n6030), .A2(DATAI_9_), .B1(n6830), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U6583 ( .A1(n6028), .A2(DATAI_25_), .ZN(n5386) );
  OAI211_X1 U6584 ( .C1(n5388), .C2(n5418), .A(n5387), .B(n5386), .ZN(U2866)
         );
  AOI22_X1 U6585 ( .A1(n6030), .A2(DATAI_8_), .B1(n6830), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6586 ( .A1(n6028), .A2(DATAI_24_), .ZN(n5389) );
  OAI211_X1 U6587 ( .C1(n5391), .C2(n5418), .A(n5390), .B(n5389), .ZN(U2867)
         );
  AOI22_X1 U6588 ( .A1(n6030), .A2(DATAI_7_), .B1(n6830), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5393) );
  NAND2_X1 U6589 ( .A1(n6028), .A2(DATAI_23_), .ZN(n5392) );
  OAI211_X1 U6590 ( .C1(n5821), .C2(n5418), .A(n5393), .B(n5392), .ZN(U2868)
         );
  AOI22_X1 U6591 ( .A1(n6030), .A2(DATAI_6_), .B1(n6830), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U6592 ( .A1(n6028), .A2(DATAI_22_), .ZN(n5394) );
  OAI211_X1 U6593 ( .C1(n5396), .C2(n5418), .A(n5395), .B(n5394), .ZN(U2869)
         );
  AOI22_X1 U6594 ( .A1(n6030), .A2(DATAI_5_), .B1(n6830), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U6595 ( .A1(n6028), .A2(DATAI_21_), .ZN(n5397) );
  OAI211_X1 U6596 ( .C1(n5399), .C2(n5418), .A(n5398), .B(n5397), .ZN(U2870)
         );
  AOI22_X1 U6597 ( .A1(n6030), .A2(DATAI_4_), .B1(n6830), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6598 ( .A1(n6028), .A2(DATAI_20_), .ZN(n5400) );
  OAI211_X1 U6599 ( .C1(n5843), .C2(n5418), .A(n5401), .B(n5400), .ZN(U2871)
         );
  AOI22_X1 U6600 ( .A1(n6030), .A2(DATAI_3_), .B1(n6830), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U6601 ( .A1(n6028), .A2(DATAI_19_), .ZN(n5402) );
  OAI211_X1 U6602 ( .C1(n5852), .C2(n5418), .A(n5403), .B(n5402), .ZN(U2872)
         );
  AOI22_X1 U6603 ( .A1(n6030), .A2(DATAI_2_), .B1(n6830), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6604 ( .A1(n6028), .A2(DATAI_18_), .ZN(n5404) );
  OAI211_X1 U6605 ( .C1(n5508), .C2(n5418), .A(n5405), .B(n5404), .ZN(U2873)
         );
  AOI22_X1 U6606 ( .A1(n6030), .A2(DATAI_0_), .B1(n6830), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5407) );
  NAND2_X1 U6607 ( .A1(n6028), .A2(DATAI_16_), .ZN(n5406) );
  OAI211_X1 U6608 ( .C1(n5524), .C2(n5418), .A(n5407), .B(n5406), .ZN(U2875)
         );
  AOI22_X1 U6609 ( .A1(n6831), .A2(DATAI_15_), .B1(n6830), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5408) );
  OAI21_X1 U6610 ( .B1(n5409), .B2(n5418), .A(n5408), .ZN(U2876) );
  AOI22_X1 U6611 ( .A1(n6831), .A2(DATAI_14_), .B1(n6830), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5410) );
  OAI21_X1 U6612 ( .B1(n5543), .B2(n5418), .A(n5410), .ZN(U2877) );
  INV_X1 U6613 ( .A(n5411), .ZN(n5414) );
  INV_X1 U6614 ( .A(n5412), .ZN(n5413) );
  AOI21_X1 U6615 ( .B1(n5414), .B2(n5413), .A(n5051), .ZN(n6016) );
  INV_X1 U6616 ( .A(n6016), .ZN(n5416) );
  AOI22_X1 U6617 ( .A1(n6831), .A2(DATAI_12_), .B1(n6830), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5415) );
  OAI21_X1 U6618 ( .B1(n5416), .B2(n5418), .A(n5415), .ZN(U2879) );
  INV_X1 U6619 ( .A(DATAI_11_), .ZN(n5420) );
  INV_X1 U6620 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6784) );
  OAI222_X1 U6621 ( .A1(n5421), .A2(n5420), .B1(n5419), .B2(n6784), .C1(n5418), 
        .C2(n5417), .ZN(U2880) );
  NAND2_X1 U6622 ( .A1(n5422), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5424) );
  INV_X1 U6623 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U6624 ( .A1(n5425), .A2(n5579), .ZN(n5423) );
  NOR2_X1 U6625 ( .A1(n5427), .A2(n5426), .ZN(n5583) );
  NOR2_X1 U6626 ( .A1(n6190), .A2(n5428), .ZN(n5577) );
  AOI21_X1 U6627 ( .B1(n6097), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5577), 
        .ZN(n5429) );
  OAI21_X1 U6628 ( .B1(n5430), .B2(n6108), .A(n5429), .ZN(n5431) );
  AOI21_X1 U6629 ( .B1(n5432), .B2(n6101), .A(n5431), .ZN(n5433) );
  OAI21_X1 U6630 ( .B1(n5583), .B2(n6078), .A(n5433), .ZN(U2957) );
  NAND2_X1 U6631 ( .A1(n5435), .A2(n5434), .ZN(n5436) );
  XOR2_X1 U6632 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .B(n5436), .Z(n5592) );
  INV_X1 U6633 ( .A(n5592), .ZN(n5441) );
  INV_X1 U6634 ( .A(n5794), .ZN(n5439) );
  NOR2_X1 U6635 ( .A1(n6190), .A2(n6548), .ZN(n5594) );
  AOI21_X1 U6636 ( .B1(n6097), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5594), 
        .ZN(n5437) );
  OAI21_X1 U6637 ( .B1(n5790), .B2(n6108), .A(n5437), .ZN(n5438) );
  AOI21_X1 U6638 ( .B1(n5439), .B2(n6101), .A(n5438), .ZN(n5440) );
  OAI21_X1 U6639 ( .B1(n5441), .B2(n6078), .A(n5440), .ZN(U2959) );
  NOR2_X1 U6640 ( .A1(n5443), .A2(n5442), .ZN(n5445) );
  XOR2_X1 U6641 ( .A(n5445), .B(n5444), .Z(n5609) );
  NAND2_X1 U6642 ( .A1(n6074), .A2(n5446), .ZN(n5447) );
  NAND2_X1 U6643 ( .A1(n6156), .A2(REIP_REG_26__SCAN_IN), .ZN(n5600) );
  OAI211_X1 U6644 ( .C1(n5548), .C2(n5448), .A(n5447), .B(n5600), .ZN(n5449)
         );
  AOI21_X1 U6645 ( .B1(n5450), .B2(n6101), .A(n5449), .ZN(n5451) );
  OAI21_X1 U6646 ( .B1(n5609), .B2(n6078), .A(n5451), .ZN(U2960) );
  AOI21_X1 U6647 ( .B1(n5454), .B2(n5116), .A(n5453), .ZN(n5617) );
  NAND2_X1 U6648 ( .A1(n6156), .A2(REIP_REG_25__SCAN_IN), .ZN(n5611) );
  INV_X1 U6649 ( .A(n5611), .ZN(n5455) );
  AOI21_X1 U6650 ( .B1(n6097), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5455), 
        .ZN(n5456) );
  OAI21_X1 U6651 ( .B1(n6108), .B2(n5802), .A(n5456), .ZN(n5457) );
  AOI21_X1 U6652 ( .B1(n5804), .B2(n6101), .A(n5457), .ZN(n5458) );
  OAI21_X1 U6653 ( .B1(n5617), .B2(n6078), .A(n5458), .ZN(U2961) );
  INV_X1 U6654 ( .A(n5459), .ZN(n5491) );
  NAND3_X1 U6655 ( .A1(n5491), .A2(n5461), .A3(n5460), .ZN(n5462) );
  NAND2_X1 U6656 ( .A1(n5463), .A2(n5462), .ZN(n5464) );
  XNOR2_X1 U6657 ( .A(n5464), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5625)
         );
  NOR2_X1 U6658 ( .A1(n6190), .A2(n6541), .ZN(n5618) );
  AOI21_X1 U6659 ( .B1(n6097), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n5618), 
        .ZN(n5465) );
  OAI21_X1 U6660 ( .B1(n6108), .B2(n5818), .A(n5465), .ZN(n5466) );
  AOI21_X1 U6661 ( .B1(n5467), .B2(n6101), .A(n5466), .ZN(n5468) );
  OAI21_X1 U6662 ( .B1(n5625), .B2(n6078), .A(n5468), .ZN(U2963) );
  AOI21_X1 U6663 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5557), .A(n5469), 
        .ZN(n5471) );
  XOR2_X1 U6664 ( .A(n5471), .B(n5470), .Z(n5633) );
  NOR2_X1 U6665 ( .A1(n6190), .A2(n6875), .ZN(n5628) );
  NOR2_X1 U6666 ( .A1(n5548), .A2(n6772), .ZN(n5472) );
  AOI211_X1 U6667 ( .C1(n6074), .C2(n5473), .A(n5628), .B(n5472), .ZN(n5476)
         );
  NAND2_X1 U6668 ( .A1(n5474), .A2(n6101), .ZN(n5475) );
  OAI211_X1 U6669 ( .C1(n5633), .C2(n6078), .A(n5476), .B(n5475), .ZN(U2964)
         );
  AOI21_X1 U6670 ( .B1(n5479), .B2(n5478), .A(n5477), .ZN(n5640) );
  NOR2_X1 U6671 ( .A1(n6190), .A2(n6539), .ZN(n5635) );
  AOI21_X1 U6672 ( .B1(n6097), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5635), 
        .ZN(n5480) );
  OAI21_X1 U6673 ( .B1(n6108), .B2(n5837), .A(n5480), .ZN(n5481) );
  AOI21_X1 U6674 ( .B1(n5834), .B2(n6101), .A(n5481), .ZN(n5482) );
  OAI21_X1 U6675 ( .B1(n5640), .B2(n6078), .A(n5482), .ZN(U2965) );
  INV_X1 U6676 ( .A(n5483), .ZN(n5485) );
  NAND2_X1 U6677 ( .A1(n5485), .A2(n5484), .ZN(n5486) );
  XNOR2_X1 U6678 ( .A(n5487), .B(n5486), .ZN(n5651) );
  NAND2_X1 U6679 ( .A1(n6156), .A2(REIP_REG_20__SCAN_IN), .ZN(n5647) );
  OAI21_X1 U6680 ( .B1(n5548), .B2(n6702), .A(n5647), .ZN(n5489) );
  NOR2_X1 U6681 ( .A1(n5843), .A2(n5564), .ZN(n5488) );
  AOI211_X1 U6682 ( .C1(n6074), .C2(n5845), .A(n5489), .B(n5488), .ZN(n5490)
         );
  OAI21_X1 U6683 ( .B1(n5651), .B2(n6078), .A(n5490), .ZN(U2966) );
  INV_X1 U6684 ( .A(n5492), .ZN(n5494) );
  NAND2_X1 U6685 ( .A1(n5494), .A2(n5493), .ZN(n5653) );
  NAND3_X1 U6686 ( .A1(n5459), .A2(n6104), .A3(n5653), .ZN(n5498) );
  INV_X1 U6687 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5495) );
  NOR2_X1 U6688 ( .A1(n6190), .A2(n5495), .ZN(n5654) );
  NOR2_X1 U6689 ( .A1(n6108), .A2(n5854), .ZN(n5496) );
  AOI211_X1 U6690 ( .C1(n6097), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5654), 
        .B(n5496), .ZN(n5497) );
  OAI211_X1 U6691 ( .C1(n5564), .C2(n5852), .A(n5498), .B(n5497), .ZN(U2967)
         );
  NAND3_X1 U6692 ( .A1(n5517), .A2(n5716), .A3(n5500), .ZN(n5509) );
  NAND3_X1 U6693 ( .A1(n5501), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5557), .ZN(n5502) );
  OAI21_X1 U6694 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5509), .A(n5502), 
        .ZN(n5503) );
  XOR2_X1 U6695 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .B(n5503), .Z(n5668) );
  NAND2_X1 U6696 ( .A1(n5668), .A2(n6104), .ZN(n5507) );
  NOR2_X1 U6697 ( .A1(n6190), .A2(n6535), .ZN(n5660) );
  NOR2_X1 U6698 ( .A1(n6108), .A2(n5504), .ZN(n5505) );
  AOI211_X1 U6699 ( .C1(n6097), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5660), 
        .B(n5505), .ZN(n5506) );
  OAI211_X1 U6700 ( .C1(n5564), .C2(n5508), .A(n5507), .B(n5506), .ZN(U2968)
         );
  NAND2_X1 U6701 ( .A1(n5557), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5510) );
  OAI21_X1 U6702 ( .B1(n5517), .B2(n5510), .A(n5509), .ZN(n5511) );
  XNOR2_X1 U6703 ( .A(n5511), .B(n4271), .ZN(n5676) );
  NAND2_X1 U6704 ( .A1(n5676), .A2(n6104), .ZN(n5515) );
  INV_X1 U6705 ( .A(REIP_REG_17__SCAN_IN), .ZN(n5512) );
  NOR2_X1 U6706 ( .A1(n6190), .A2(n5512), .ZN(n5671) );
  NOR2_X1 U6707 ( .A1(n6108), .A2(n5916), .ZN(n5513) );
  AOI211_X1 U6708 ( .C1(n6097), .C2(PHYADDRPOINTER_REG_17__SCAN_IN), .A(n5671), 
        .B(n5513), .ZN(n5514) );
  OAI211_X1 U6709 ( .C1(n5564), .C2(n5912), .A(n5515), .B(n5514), .ZN(U2969)
         );
  XNOR2_X1 U6710 ( .A(n5557), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5516)
         );
  XNOR2_X1 U6711 ( .A(n5517), .B(n5516), .ZN(n5861) );
  NAND2_X1 U6712 ( .A1(n5861), .A2(n6104), .ZN(n5523) );
  INV_X1 U6713 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5518) );
  OAI22_X1 U6714 ( .A1(n5548), .A2(n5519), .B1(n6190), .B2(n5518), .ZN(n5520)
         );
  AOI21_X1 U6715 ( .B1(n5521), .B2(n6074), .A(n5520), .ZN(n5522) );
  OAI211_X1 U6716 ( .C1(n5564), .C2(n5524), .A(n5523), .B(n5522), .ZN(U2970)
         );
  INV_X1 U6717 ( .A(n5526), .ZN(n5527) );
  NOR2_X1 U6718 ( .A1(n5528), .A2(n5527), .ZN(n5529) );
  XNOR2_X1 U6719 ( .A(n5525), .B(n5529), .ZN(n5686) );
  NAND2_X1 U6720 ( .A1(n6074), .A2(n5530), .ZN(n5531) );
  NAND2_X1 U6721 ( .A1(n6156), .A2(REIP_REG_15__SCAN_IN), .ZN(n5682) );
  OAI211_X1 U6722 ( .C1(n5548), .C2(n3716), .A(n5531), .B(n5682), .ZN(n5532)
         );
  AOI21_X1 U6723 ( .B1(n5533), .B2(n6101), .A(n5532), .ZN(n5534) );
  OAI21_X1 U6724 ( .B1(n5686), .B2(n6078), .A(n5534), .ZN(U2971) );
  XNOR2_X1 U6725 ( .A(n5557), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5535)
         );
  XNOR2_X1 U6726 ( .A(n5536), .B(n5535), .ZN(n5870) );
  NAND2_X1 U6727 ( .A1(n5870), .A2(n6104), .ZN(n5542) );
  INV_X1 U6728 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5537) );
  OAI22_X1 U6729 ( .A1(n5548), .A2(n5538), .B1(n6190), .B2(n5537), .ZN(n5539)
         );
  AOI21_X1 U6730 ( .B1(n6074), .B2(n5540), .A(n5539), .ZN(n5541) );
  OAI211_X1 U6731 ( .C1(n5564), .C2(n5543), .A(n5542), .B(n5541), .ZN(U2972)
         );
  OAI21_X1 U6732 ( .B1(n5546), .B2(n5545), .A(n5544), .ZN(n5687) );
  NAND2_X1 U6733 ( .A1(n5687), .A2(n6104), .ZN(n5551) );
  INV_X1 U6734 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U6735 ( .A1(n6156), .A2(REIP_REG_13__SCAN_IN), .ZN(n5693) );
  OAI21_X1 U6736 ( .B1(n5548), .B2(n5547), .A(n5693), .ZN(n5549) );
  AOI21_X1 U6737 ( .B1(n6074), .B2(n5918), .A(n5549), .ZN(n5550) );
  OAI211_X1 U6738 ( .C1(n5564), .C2(n5917), .A(n5551), .B(n5550), .ZN(U2973)
         );
  XOR2_X1 U6739 ( .A(n5553), .B(n5552), .Z(n5712) );
  NOR2_X1 U6740 ( .A1(n6190), .A2(n6527), .ZN(n5702) );
  AOI21_X1 U6741 ( .B1(n6097), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n5702), 
        .ZN(n5554) );
  OAI21_X1 U6742 ( .B1(n6108), .B2(n5931), .A(n5554), .ZN(n5555) );
  AOI21_X1 U6743 ( .B1(n6016), .B2(n6101), .A(n5555), .ZN(n5556) );
  OAI21_X1 U6744 ( .B1(n5712), .B2(n6078), .A(n5556), .ZN(U2974) );
  XNOR2_X1 U6745 ( .A(n5557), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5558)
         );
  XNOR2_X1 U6746 ( .A(n5713), .B(n5558), .ZN(n6112) );
  NAND2_X1 U6747 ( .A1(n6112), .A2(n6104), .ZN(n5562) );
  NOR2_X1 U6748 ( .A1(n6190), .A2(n6521), .ZN(n6109) );
  NOR2_X1 U6749 ( .A1(n6108), .A2(n5559), .ZN(n5560) );
  AOI211_X1 U6750 ( .C1(n6097), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6109), 
        .B(n5560), .ZN(n5561) );
  OAI211_X1 U6751 ( .C1(n5564), .C2(n5563), .A(n5562), .B(n5561), .ZN(U2976)
         );
  INV_X1 U6752 ( .A(n5565), .ZN(n5572) );
  NAND3_X1 U6753 ( .A1(n5580), .A2(n5566), .A3(n5568), .ZN(n5567) );
  OAI21_X1 U6754 ( .B1(n5569), .B2(n5568), .A(n5567), .ZN(n5570) );
  AOI211_X1 U6755 ( .C1(n5572), .C2(n6174), .A(n5571), .B(n5570), .ZN(n5573)
         );
  OAI21_X1 U6756 ( .B1(n5574), .B2(n6184), .A(n5573), .ZN(U2987) );
  NOR2_X1 U6757 ( .A1(n5575), .A2(n6127), .ZN(n5576) );
  AOI211_X1 U6758 ( .C1(INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n5578), .A(n5577), .B(n5576), .ZN(n5582) );
  NAND2_X1 U6759 ( .A1(n5580), .A2(n5579), .ZN(n5581) );
  OAI211_X1 U6760 ( .C1(n5583), .C2(n6184), .A(n5582), .B(n5581), .ZN(U2989)
         );
  INV_X1 U6761 ( .A(n5584), .ZN(n5595) );
  XNOR2_X1 U6762 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .B(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5585) );
  NOR2_X1 U6763 ( .A1(n5598), .A2(n5585), .ZN(n5589) );
  OAI21_X1 U6764 ( .B1(n5587), .B2(n6127), .A(n5586), .ZN(n5588) );
  AOI211_X1 U6765 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n5595), .A(n5589), .B(n5588), .ZN(n5590) );
  OAI21_X1 U6766 ( .B1(n5591), .B2(n6184), .A(n5590), .ZN(U2990) );
  NAND2_X1 U6767 ( .A1(n5592), .A2(n6167), .ZN(n5597) );
  NOR2_X1 U6768 ( .A1(n5793), .A2(n6127), .ZN(n5593) );
  AOI211_X1 U6769 ( .C1(n5595), .C2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5594), .B(n5593), .ZN(n5596) );
  OAI211_X1 U6770 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5598), .A(n5597), .B(n5596), .ZN(U2991) );
  INV_X1 U6771 ( .A(n5599), .ZN(n5602) );
  INV_X1 U6772 ( .A(n5600), .ZN(n5601) );
  AOI21_X1 U6773 ( .B1(n5602), .B2(n6174), .A(n5601), .ZN(n5608) );
  INV_X1 U6774 ( .A(n5603), .ZN(n5604) );
  OAI22_X1 U6775 ( .A1(n5610), .A2(n5605), .B1(n5604), .B2(n5612), .ZN(n5606)
         );
  OAI21_X1 U6776 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5606), .ZN(n5607) );
  OAI211_X1 U6777 ( .C1(n5609), .C2(n6184), .A(n5608), .B(n5607), .ZN(U2992)
         );
  INV_X1 U6778 ( .A(n5610), .ZN(n5615) );
  OAI21_X1 U6779 ( .B1(n5809), .B2(n6127), .A(n5611), .ZN(n5614) );
  NOR2_X1 U6780 ( .A1(n5612), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5613)
         );
  AOI211_X1 U6781 ( .C1(n5615), .C2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5614), .B(n5613), .ZN(n5616) );
  OAI21_X1 U6782 ( .B1(n5617), .B2(n6184), .A(n5616), .ZN(U2993) );
  AOI21_X1 U6783 ( .B1(n5619), .B2(n6174), .A(n5618), .ZN(n5620) );
  OAI21_X1 U6784 ( .B1(n5621), .B2(n5062), .A(n5620), .ZN(n5622) );
  AOI21_X1 U6785 ( .B1(n5623), .B2(n5062), .A(n5622), .ZN(n5624) );
  OAI21_X1 U6786 ( .B1(n5625), .B2(n6184), .A(n5624), .ZN(U2995) );
  NOR2_X1 U6787 ( .A1(n5626), .A2(n6127), .ZN(n5627) );
  AOI211_X1 U6788 ( .C1(n5636), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5628), .B(n5627), .ZN(n5632) );
  NAND3_X1 U6789 ( .A1(n5637), .A2(n5630), .A3(n5629), .ZN(n5631) );
  OAI211_X1 U6790 ( .C1(n5633), .C2(n6184), .A(n5632), .B(n5631), .ZN(U2996)
         );
  NOR2_X1 U6791 ( .A1(n5832), .A2(n6127), .ZN(n5634) );
  AOI211_X1 U6792 ( .C1(n5636), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5635), .B(n5634), .ZN(n5639) );
  NAND2_X1 U6793 ( .A1(n5637), .A2(n6760), .ZN(n5638) );
  OAI211_X1 U6794 ( .C1(n5640), .C2(n6184), .A(n5639), .B(n5638), .ZN(U2997)
         );
  NAND2_X1 U6795 ( .A1(n5642), .A2(n5641), .ZN(n5705) );
  AND2_X1 U6796 ( .A1(n5705), .A2(n4271), .ZN(n5643) );
  NOR2_X1 U6797 ( .A1(n5670), .A2(n5643), .ZN(n5666) );
  OAI21_X1 U6798 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5679), .A(n5666), 
        .ZN(n5652) );
  NOR2_X1 U6799 ( .A1(n5674), .A2(n5644), .ZN(n5656) );
  NAND3_X1 U6800 ( .A1(n5656), .A2(n5646), .A3(n5645), .ZN(n5648) );
  OAI211_X1 U6801 ( .C1(n5847), .C2(n6127), .A(n5648), .B(n5647), .ZN(n5649)
         );
  AOI21_X1 U6802 ( .B1(n5652), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5649), 
        .ZN(n5650) );
  OAI21_X1 U6803 ( .B1(n5651), .B2(n6184), .A(n5650), .ZN(U2998) );
  INV_X1 U6804 ( .A(n5652), .ZN(n5659) );
  NAND3_X1 U6805 ( .A1(n5459), .A2(n6167), .A3(n5653), .ZN(n5658) );
  NOR2_X1 U6806 ( .A1(n5853), .A2(n6127), .ZN(n5655) );
  AOI211_X1 U6807 ( .C1(n5656), .C2(n6871), .A(n5655), .B(n5654), .ZN(n5657)
         );
  OAI211_X1 U6808 ( .C1(n5659), .C2(n6871), .A(n5658), .B(n5657), .ZN(U2999)
         );
  INV_X1 U6809 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5665) );
  AOI21_X1 U6810 ( .B1(n5661), .B2(n6174), .A(n5660), .ZN(n5664) );
  INV_X1 U6811 ( .A(n5674), .ZN(n5662) );
  NAND3_X1 U6812 ( .A1(n5662), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5665), .ZN(n5663) );
  OAI211_X1 U6813 ( .C1(n5666), .C2(n5665), .A(n5664), .B(n5663), .ZN(n5667)
         );
  AOI21_X1 U6814 ( .B1(n5668), .B2(n6167), .A(n5667), .ZN(n5669) );
  INV_X1 U6815 ( .A(n5669), .ZN(U3000) );
  NAND2_X1 U6816 ( .A1(n5670), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5673) );
  AOI21_X1 U6817 ( .B1(n5913), .B2(n6174), .A(n5671), .ZN(n5672) );
  OAI211_X1 U6818 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5674), .A(n5673), .B(n5672), .ZN(n5675) );
  AOI21_X1 U6819 ( .B1(n5676), .B2(n6167), .A(n5675), .ZN(n5677) );
  INV_X1 U6820 ( .A(n5677), .ZN(U3001) );
  INV_X1 U6821 ( .A(n5680), .ZN(n5678) );
  OAI21_X1 U6822 ( .B1(n5679), .B2(n5678), .A(n5703), .ZN(n5862) );
  INV_X1 U6823 ( .A(n5875), .ZN(n5707) );
  NOR3_X1 U6824 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n5707), .A3(n5680), 
        .ZN(n5863) );
  INV_X1 U6825 ( .A(n5863), .ZN(n5681) );
  OAI211_X1 U6826 ( .C1(n6127), .C2(n5683), .A(n5682), .B(n5681), .ZN(n5684)
         );
  AOI21_X1 U6827 ( .B1(n5862), .B2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5684), 
        .ZN(n5685) );
  OAI21_X1 U6828 ( .B1(n5686), .B2(n6184), .A(n5685), .ZN(U3003) );
  INV_X1 U6829 ( .A(n5687), .ZN(n5698) );
  NAND2_X1 U6830 ( .A1(n5704), .A2(n5688), .ZN(n5689) );
  OAI211_X1 U6831 ( .C1(n5876), .C2(n5690), .A(n5703), .B(n5689), .ZN(n5873)
         );
  XOR2_X1 U6832 ( .A(n5691), .B(n5699), .Z(n6011) );
  INV_X1 U6833 ( .A(n6011), .ZN(n5695) );
  NOR2_X1 U6834 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5704), .ZN(n5692)
         );
  NAND2_X1 U6835 ( .A1(n5875), .A2(n5692), .ZN(n5694) );
  OAI211_X1 U6836 ( .C1(n5695), .C2(n6127), .A(n5694), .B(n5693), .ZN(n5696)
         );
  AOI21_X1 U6837 ( .B1(n5873), .B2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(n5696), 
        .ZN(n5697) );
  OAI21_X1 U6838 ( .B1(n5698), .B2(n6184), .A(n5697), .ZN(U3005) );
  AOI21_X1 U6839 ( .B1(n5701), .B2(n5700), .A(n5699), .ZN(n6015) );
  AOI21_X1 U6840 ( .B1(n6174), .B2(n6015), .A(n5702), .ZN(n5711) );
  INV_X1 U6841 ( .A(n5703), .ZN(n5722) );
  AND2_X1 U6842 ( .A1(n5705), .A2(n5704), .ZN(n5709) );
  OAI21_X1 U6843 ( .B1(n5707), .B2(n3153), .A(n5706), .ZN(n5708) );
  OAI21_X1 U6844 ( .B1(n5722), .B2(n5709), .A(n5708), .ZN(n5710) );
  OAI211_X1 U6845 ( .C1(n5712), .C2(n6184), .A(n5711), .B(n5710), .ZN(U3006)
         );
  INV_X1 U6846 ( .A(n5713), .ZN(n5714) );
  AOI22_X1 U6847 ( .A1(n5716), .A2(n5715), .B1(n5714), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5718) );
  XNOR2_X1 U6848 ( .A(n5716), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5717)
         );
  XNOR2_X1 U6849 ( .A(n5718), .B(n5717), .ZN(n6079) );
  INV_X1 U6850 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6525) );
  INV_X1 U6851 ( .A(n5937), .ZN(n5719) );
  NAND2_X1 U6852 ( .A1(n6174), .A2(n5719), .ZN(n5720) );
  OAI21_X1 U6853 ( .B1(n6525), .B2(n6190), .A(n5720), .ZN(n5721) );
  AOI21_X1 U6854 ( .B1(n5722), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n5721), 
        .ZN(n5724) );
  NAND2_X1 U6855 ( .A1(n5875), .A2(n3153), .ZN(n5723) );
  OAI211_X1 U6856 ( .C1(n6079), .C2(n6184), .A(n5724), .B(n5723), .ZN(U3007)
         );
  NAND2_X1 U6857 ( .A1(n5726), .A2(n5725), .ZN(n6483) );
  AOI22_X1 U6858 ( .A1(n5728), .A2(n6380), .B1(n3102), .B2(n5727), .ZN(n5729)
         );
  NAND2_X1 U6859 ( .A1(n6483), .A2(n5729), .ZN(n5730) );
  MUX2_X1 U6860 ( .A(n5730), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .S(n6191), 
        .Z(U3465) );
  INV_X1 U6861 ( .A(n5731), .ZN(n5732) );
  NOR3_X1 U6862 ( .A1(n6440), .A2(n5784), .A3(n6393), .ZN(n5734) );
  OAI22_X1 U6863 ( .A1(n5734), .A2(n6331), .B1(n6263), .B2(n5733), .ZN(n5739)
         );
  NOR2_X1 U6864 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5735), .ZN(n5743)
         );
  OR2_X1 U6865 ( .A1(n5743), .A2(n6688), .ZN(n5736) );
  NAND4_X1 U6866 ( .A1(n5739), .A2(n5738), .A3(n5737), .A4(n5736), .ZN(n5779)
         );
  NAND2_X1 U6867 ( .A1(n5779), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5747)
         );
  AOI22_X1 U6868 ( .A1(n5742), .A2(n5741), .B1(n5740), .B2(n6258), .ZN(n5782)
         );
  INV_X1 U6869 ( .A(n5743), .ZN(n5780) );
  OAI22_X1 U6870 ( .A1(n6400), .A2(n5782), .B1(n5744), .B2(n5780), .ZN(n5745)
         );
  AOI21_X1 U6871 ( .B1(n6389), .B2(n5784), .A(n5745), .ZN(n5746) );
  OAI211_X1 U6872 ( .C1(n5788), .C2(n5748), .A(n5747), .B(n5746), .ZN(U3116)
         );
  NAND2_X1 U6873 ( .A1(n5779), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5752)
         );
  OAI22_X1 U6874 ( .A1(n6406), .A2(n5782), .B1(n5749), .B2(n5780), .ZN(n5750)
         );
  AOI21_X1 U6875 ( .B1(n6403), .B2(n5784), .A(n5750), .ZN(n5751) );
  OAI211_X1 U6876 ( .C1(n5788), .C2(n5753), .A(n5752), .B(n5751), .ZN(U3117)
         );
  NAND2_X1 U6877 ( .A1(n5779), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5757)
         );
  OAI22_X1 U6878 ( .A1(n6412), .A2(n5782), .B1(n5754), .B2(n5780), .ZN(n5755)
         );
  AOI21_X1 U6879 ( .B1(n6408), .B2(n5784), .A(n5755), .ZN(n5756) );
  OAI211_X1 U6880 ( .C1(n5788), .C2(n5758), .A(n5757), .B(n5756), .ZN(U3118)
         );
  NAND2_X1 U6881 ( .A1(n5779), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5762)
         );
  OAI22_X1 U6882 ( .A1(n6418), .A2(n5782), .B1(n5759), .B2(n5780), .ZN(n5760)
         );
  AOI21_X1 U6883 ( .B1(n6415), .B2(n5784), .A(n5760), .ZN(n5761) );
  OAI211_X1 U6884 ( .C1(n5788), .C2(n5763), .A(n5762), .B(n5761), .ZN(U3119)
         );
  NAND2_X1 U6885 ( .A1(n5779), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5767)
         );
  OAI22_X1 U6886 ( .A1(n6424), .A2(n5782), .B1(n5764), .B2(n5780), .ZN(n5765)
         );
  AOI21_X1 U6887 ( .B1(n6421), .B2(n5784), .A(n5765), .ZN(n5766) );
  OAI211_X1 U6888 ( .C1(n5788), .C2(n5768), .A(n5767), .B(n5766), .ZN(U3120)
         );
  NAND2_X1 U6889 ( .A1(n5779), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5772)
         );
  OAI22_X1 U6890 ( .A1(n6430), .A2(n5782), .B1(n5769), .B2(n5780), .ZN(n5770)
         );
  AOI21_X1 U6891 ( .B1(n6427), .B2(n5784), .A(n5770), .ZN(n5771) );
  OAI211_X1 U6892 ( .C1(n5788), .C2(n5773), .A(n5772), .B(n5771), .ZN(U3121)
         );
  NAND2_X1 U6893 ( .A1(n5779), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5777)
         );
  OAI22_X1 U6894 ( .A1(n6436), .A2(n5782), .B1(n5774), .B2(n5780), .ZN(n5775)
         );
  AOI21_X1 U6895 ( .B1(n6433), .B2(n5784), .A(n5775), .ZN(n5776) );
  OAI211_X1 U6896 ( .C1(n5788), .C2(n5778), .A(n5777), .B(n5776), .ZN(U3122)
         );
  NAND2_X1 U6897 ( .A1(n5779), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5786)
         );
  OAI22_X1 U6898 ( .A1(n6446), .A2(n5782), .B1(n5781), .B2(n5780), .ZN(n5783)
         );
  AOI21_X1 U6899 ( .B1(n6439), .B2(n5784), .A(n5783), .ZN(n5785) );
  OAI211_X1 U6900 ( .C1(n5788), .C2(n5787), .A(n5786), .B(n5785), .ZN(U3123)
         );
  INV_X1 U6901 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n6641) );
  NOR2_X1 U6902 ( .A1(n6641), .A2(n6059), .ZN(U2892) );
  AOI22_X1 U6903 ( .A1(EBX_REG_27__SCAN_IN), .A2(n5995), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n5990), .ZN(n5789) );
  OAI21_X1 U6904 ( .B1(n5790), .B2(n5993), .A(n5789), .ZN(n5791) );
  AOI21_X1 U6905 ( .B1(REIP_REG_27__SCAN_IN), .B2(n5792), .A(n5791), .ZN(n5797) );
  OAI22_X1 U6906 ( .A1(n5794), .A2(n5842), .B1(n5793), .B2(n5947), .ZN(n5795)
         );
  INV_X1 U6907 ( .A(n5795), .ZN(n5796) );
  OAI211_X1 U6908 ( .C1(REIP_REG_27__SCAN_IN), .C2(n5798), .A(n5797), .B(n5796), .ZN(U2800) );
  OAI22_X1 U6909 ( .A1(n5969), .A2(n5324), .B1(REIP_REG_25__SCAN_IN), .B2(
        n5799), .ZN(n5800) );
  AOI21_X1 U6910 ( .B1(n5990), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5800), 
        .ZN(n5801) );
  OAI21_X1 U6911 ( .B1(n5993), .B2(n5802), .A(n5801), .ZN(n5803) );
  AOI21_X1 U6912 ( .B1(n5804), .B2(n5964), .A(n5803), .ZN(n5808) );
  INV_X1 U6913 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U6914 ( .A1(n6542), .A2(n5805), .ZN(n5814) );
  AOI21_X1 U6915 ( .B1(n5814), .B2(n5826), .A(n6544), .ZN(n5806) );
  INV_X1 U6916 ( .A(n5806), .ZN(n5807) );
  OAI211_X1 U6917 ( .C1(n5947), .C2(n5809), .A(n5808), .B(n5807), .ZN(U2802)
         );
  AOI22_X1 U6918 ( .A1(EBX_REG_24__SCAN_IN), .A2(n5995), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n5990), .ZN(n5817) );
  INV_X1 U6919 ( .A(n5826), .ZN(n5811) );
  AOI22_X1 U6920 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5811), .B1(n5810), .B2(
        n6006), .ZN(n5816) );
  AOI22_X1 U6921 ( .A1(n5813), .A2(n5964), .B1(n5812), .B2(n5980), .ZN(n5815)
         );
  NAND4_X1 U6922 ( .A1(n5817), .A2(n5816), .A3(n5815), .A4(n5814), .ZN(U2803)
         );
  INV_X1 U6923 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5819) );
  OAI22_X1 U6924 ( .A1(n5819), .A2(n6000), .B1(n5818), .B2(n5993), .ZN(n5823)
         );
  OAI22_X1 U6925 ( .A1(n5821), .A2(n5842), .B1(n5820), .B2(n5947), .ZN(n5822)
         );
  AOI211_X1 U6926 ( .C1(EBX_REG_23__SCAN_IN), .C2(n5995), .A(n5823), .B(n5822), 
        .ZN(n5824) );
  OAI221_X1 U6927 ( .B1(n5826), .B2(n6541), .C1(n5826), .C2(n5825), .A(n5824), 
        .ZN(U2804) );
  NOR2_X1 U6928 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5827), .ZN(n5831) );
  OAI22_X1 U6929 ( .A1(n5829), .A2(n6000), .B1(n6539), .B2(n5828), .ZN(n5830)
         );
  AOI211_X1 U6930 ( .C1(n5995), .C2(EBX_REG_21__SCAN_IN), .A(n5831), .B(n5830), 
        .ZN(n5836) );
  INV_X1 U6931 ( .A(n5832), .ZN(n5833) );
  AOI22_X1 U6932 ( .A1(n5834), .A2(n5964), .B1(n5980), .B2(n5833), .ZN(n5835)
         );
  OAI211_X1 U6933 ( .C1(n5837), .C2(n5993), .A(n5836), .B(n5835), .ZN(U2806)
         );
  OAI21_X1 U6934 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5839), .A(n5838), .ZN(n5841) );
  AOI22_X1 U6935 ( .A1(n5990), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n5995), .ZN(n5840) );
  OAI211_X1 U6936 ( .C1(n5843), .C2(n5842), .A(n5841), .B(n5840), .ZN(n5844)
         );
  AOI21_X1 U6937 ( .B1(n5845), .B2(n6006), .A(n5844), .ZN(n5846) );
  OAI21_X1 U6938 ( .B1(n5847), .B2(n5947), .A(n5846), .ZN(U2807) );
  OAI21_X1 U6939 ( .B1(REIP_REG_19__SCAN_IN), .B2(REIP_REG_18__SCAN_IN), .A(
        n5848), .ZN(n5849) );
  OAI22_X1 U6940 ( .A1(n5495), .A2(n5909), .B1(n5850), .B2(n5849), .ZN(n5851)
         );
  AOI211_X1 U6941 ( .C1(n5990), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5984), 
        .B(n5851), .ZN(n5858) );
  INV_X1 U6942 ( .A(n5852), .ZN(n5856) );
  OAI22_X1 U6943 ( .A1(n5993), .A2(n5854), .B1(n5947), .B2(n5853), .ZN(n5855)
         );
  AOI21_X1 U6944 ( .B1(n5856), .B2(n5964), .A(n5855), .ZN(n5857) );
  OAI211_X1 U6945 ( .C1(n5859), .C2(n5969), .A(n5858), .B(n5857), .ZN(U2808)
         );
  AOI22_X1 U6946 ( .A1(n5861), .A2(n6167), .B1(n6174), .B2(n5860), .ZN(n5868)
         );
  NAND2_X1 U6947 ( .A1(n6156), .A2(REIP_REG_16__SCAN_IN), .ZN(n5867) );
  OAI21_X1 U6948 ( .B1(n5863), .B2(n5862), .A(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n5866) );
  NAND3_X1 U6949 ( .A1(n5864), .A2(n5500), .A3(n5875), .ZN(n5865) );
  NAND4_X1 U6950 ( .A1(n5868), .A2(n5867), .A3(n5866), .A4(n5865), .ZN(U3002)
         );
  AOI22_X1 U6951 ( .A1(n5870), .A2(n6167), .B1(n6174), .B2(n5869), .ZN(n5880)
         );
  NAND2_X1 U6952 ( .A1(n6156), .A2(REIP_REG_14__SCAN_IN), .ZN(n5879) );
  AOI21_X1 U6953 ( .B1(n5872), .B2(n5871), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5874) );
  OAI21_X1 U6954 ( .B1(n5874), .B2(n5873), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5878) );
  NAND3_X1 U6955 ( .A1(n5876), .A2(n6624), .A3(n5875), .ZN(n5877) );
  NAND4_X1 U6956 ( .A1(n5880), .A2(n5879), .A3(n5878), .A4(n5877), .ZN(U3004)
         );
  NAND4_X1 U6957 ( .A1(n5883), .A2(n5882), .A3(n5881), .A4(n5981), .ZN(n5884)
         );
  OAI21_X1 U6958 ( .B1(n6568), .B2(n5885), .A(n5884), .ZN(U3455) );
  INV_X1 U6959 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6513) );
  AOI21_X1 U6960 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6513), .A(n6507), .ZN(n5890) );
  INV_X1 U6961 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5886) );
  AOI21_X1 U6962 ( .B1(n5890), .B2(n5886), .A(n6547), .ZN(U2789) );
  NOR2_X1 U6963 ( .A1(n5887), .A2(n6485), .ZN(n5888) );
  INV_X1 U6964 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6867) );
  OAI22_X1 U6965 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6486), .B1(n5888), .B2(
        n6867), .ZN(U2790) );
  NOR2_X1 U6966 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n5891) );
  OAI21_X1 U6967 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5891), .A(n6593), .ZN(n5889)
         );
  OAI21_X1 U6968 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6580), .A(n5889), .ZN(
        U2791) );
  NOR2_X1 U6969 ( .A1(n6547), .A2(n5890), .ZN(n6560) );
  OAI21_X1 U6970 ( .B1(n5891), .B2(BS16_N), .A(n6560), .ZN(n6558) );
  OAI21_X1 U6971 ( .B1(n6560), .B2(n6584), .A(n6558), .ZN(U2792) );
  OAI21_X1 U6972 ( .B1(n5892), .B2(n6753), .A(n6078), .ZN(U2793) );
  NOR4_X1 U6973 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n5896) );
  NOR4_X1 U6974 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n5895) );
  NOR4_X1 U6975 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n5894) );
  NOR4_X1 U6976 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_22__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n5893) );
  NAND4_X1 U6977 ( .A1(n5896), .A2(n5895), .A3(n5894), .A4(n5893), .ZN(n5902)
         );
  NOR4_X1 U6978 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(
        DATAWIDTH_REG_2__SCAN_IN), .ZN(n5900) );
  AOI211_X1 U6979 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_10__SCAN_IN), .B(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5899) );
  NOR4_X1 U6980 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(
        n5898) );
  NOR4_X1 U6981 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_5__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n5897) );
  NAND4_X1 U6982 ( .A1(n5900), .A2(n5899), .A3(n5898), .A4(n5897), .ZN(n5901)
         );
  NOR2_X1 U6983 ( .A1(n5902), .A2(n5901), .ZN(n6574) );
  INV_X1 U6984 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6600) );
  NOR3_X1 U6985 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5904) );
  OAI21_X1 U6986 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5904), .A(n6574), .ZN(n5903)
         );
  OAI21_X1 U6987 ( .B1(n6574), .B2(n6600), .A(n5903), .ZN(U2794) );
  INV_X1 U6988 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6559) );
  AOI21_X1 U6989 ( .B1(n6570), .B2(n6559), .A(n5904), .ZN(n5906) );
  INV_X1 U6990 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5905) );
  INV_X1 U6991 ( .A(n6574), .ZN(n6577) );
  AOI22_X1 U6992 ( .A1(n6574), .A2(n5906), .B1(n5905), .B2(n6577), .ZN(U2795)
         );
  NOR2_X1 U6993 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5907), .ZN(n5910) );
  OAI22_X1 U6994 ( .A1(n5910), .A2(n5909), .B1(n5908), .B2(n6000), .ZN(n5911)
         );
  AOI211_X1 U6995 ( .C1(n5995), .C2(EBX_REG_17__SCAN_IN), .A(n5984), .B(n5911), 
        .ZN(n5915) );
  INV_X1 U6996 ( .A(n5912), .ZN(n6029) );
  AOI22_X1 U6997 ( .A1(n6029), .A2(n5964), .B1(n5980), .B2(n5913), .ZN(n5914)
         );
  OAI211_X1 U6998 ( .C1(n5916), .C2(n5993), .A(n5915), .B(n5914), .ZN(U2810)
         );
  INV_X1 U6999 ( .A(n5917), .ZN(n6012) );
  AOI22_X1 U7000 ( .A1(n6012), .A2(n5964), .B1(n6006), .B2(n5918), .ZN(n5928)
         );
  INV_X1 U7001 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6686) );
  OR3_X1 U7002 ( .A1(n5998), .A2(n5920), .A3(n5919), .ZN(n5922) );
  NAND2_X1 U7003 ( .A1(n5922), .A2(n5921), .ZN(n5942) );
  OAI21_X1 U7004 ( .B1(REIP_REG_12__SCAN_IN), .B2(n5935), .A(n5942), .ZN(n5925) );
  AOI22_X1 U7005 ( .A1(EBX_REG_13__SCAN_IN), .A2(n5995), .B1(n5980), .B2(n6011), .ZN(n5923) );
  OAI211_X1 U7006 ( .C1(n6000), .C2(n5547), .A(n5923), .B(n5944), .ZN(n5924)
         );
  AOI221_X1 U7007 ( .B1(n5926), .B2(n6686), .C1(n5925), .C2(
        REIP_REG_13__SCAN_IN), .A(n5924), .ZN(n5927) );
  NAND2_X1 U7008 ( .A1(n5928), .A2(n5927), .ZN(U2814) );
  OAI21_X1 U7009 ( .B1(n6000), .B2(n6870), .A(n5944), .ZN(n5930) );
  INV_X1 U7010 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6018) );
  OAI22_X1 U7011 ( .A1(n6018), .A2(n5969), .B1(n6527), .B2(n5942), .ZN(n5929)
         );
  AOI211_X1 U7012 ( .C1(n5980), .C2(n6015), .A(n5930), .B(n5929), .ZN(n5934)
         );
  INV_X1 U7013 ( .A(n5931), .ZN(n5932) );
  AOI22_X1 U7014 ( .A1(n6016), .A2(n5964), .B1(n5932), .B2(n6006), .ZN(n5933)
         );
  OAI211_X1 U7015 ( .C1(REIP_REG_12__SCAN_IN), .C2(n5935), .A(n5934), .B(n5933), .ZN(U2815) );
  NOR2_X1 U7016 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5936), .ZN(n5943) );
  OAI22_X1 U7017 ( .A1(n5938), .A2(n6000), .B1(n5947), .B2(n5937), .ZN(n5939)
         );
  AOI211_X1 U7018 ( .C1(n5995), .C2(EBX_REG_11__SCAN_IN), .A(n5984), .B(n5939), 
        .ZN(n5941) );
  AOI22_X1 U7019 ( .A1(n6075), .A2(n5964), .B1(n6006), .B2(n6073), .ZN(n5940)
         );
  OAI211_X1 U7020 ( .C1(n5943), .C2(n5942), .A(n5941), .B(n5940), .ZN(U2816)
         );
  AOI22_X1 U7021 ( .A1(EBX_REG_9__SCAN_IN), .A2(n5995), .B1(
        PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n5990), .ZN(n5945) );
  OAI211_X1 U7022 ( .C1(n5947), .C2(n5946), .A(n5945), .B(n5944), .ZN(n5948)
         );
  AOI211_X1 U7023 ( .C1(n5950), .C2(REIP_REG_9__SCAN_IN), .A(n5949), .B(n5948), 
        .ZN(n5954) );
  AOI22_X1 U7024 ( .A1(n5952), .A2(n5964), .B1(n6006), .B2(n5951), .ZN(n5953)
         );
  NAND2_X1 U7025 ( .A1(n5954), .A2(n5953), .ZN(U2818) );
  NAND2_X1 U7026 ( .A1(n5956), .A2(n5955), .ZN(n5957) );
  AND2_X1 U7027 ( .A1(n5958), .A2(n5957), .ZN(n6139) );
  INV_X1 U7028 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6745) );
  OAI22_X1 U7029 ( .A1(n6745), .A2(n5969), .B1(n3571), .B2(n6000), .ZN(n5959)
         );
  AOI211_X1 U7030 ( .C1(n5980), .C2(n6139), .A(n5984), .B(n5959), .ZN(n5962)
         );
  NAND2_X1 U7031 ( .A1(n5960), .A2(n6518), .ZN(n5961) );
  OAI211_X1 U7032 ( .C1(n6518), .C2(n5976), .A(n5962), .B(n5961), .ZN(n5963)
         );
  AOI21_X1 U7033 ( .B1(n5964), .B2(n6084), .A(n5963), .ZN(n5965) );
  OAI21_X1 U7034 ( .B1(n6087), .B2(n5993), .A(n5965), .ZN(U2821) );
  NOR2_X1 U7035 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5966), .ZN(n5977) );
  INV_X1 U7036 ( .A(n5967), .ZN(n6150) );
  INV_X1 U7037 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5968) );
  OAI22_X1 U7038 ( .A1(n6811), .A2(n5969), .B1(n5968), .B2(n6000), .ZN(n5970)
         );
  AOI211_X1 U7039 ( .C1(n5980), .C2(n6150), .A(n5984), .B(n5970), .ZN(n5975)
         );
  INV_X1 U7040 ( .A(n5971), .ZN(n5972) );
  AOI22_X1 U7041 ( .A1(n5973), .A2(n6833), .B1(n5972), .B2(n6006), .ZN(n5974)
         );
  OAI211_X1 U7042 ( .C1(n5977), .C2(n5976), .A(n5975), .B(n5974), .ZN(U2822)
         );
  INV_X1 U7043 ( .A(n5978), .ZN(n6157) );
  AOI22_X1 U7044 ( .A1(n5980), .A2(n6157), .B1(REIP_REG_4__SCAN_IN), .B2(n5979), .ZN(n5992) );
  INV_X1 U7045 ( .A(n5981), .ZN(n5987) );
  NAND3_X1 U7046 ( .A1(REIP_REG_2__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_1__SCAN_IN), .ZN(n5982) );
  NOR3_X1 U7047 ( .A1(n5983), .A2(REIP_REG_4__SCAN_IN), .A3(n5982), .ZN(n5985)
         );
  AOI211_X1 U7048 ( .C1(n5995), .C2(EBX_REG_4__SCAN_IN), .A(n5985), .B(n5984), 
        .ZN(n5986) );
  OAI21_X1 U7049 ( .B1(n5987), .B2(n5996), .A(n5986), .ZN(n5989) );
  NOR2_X1 U7050 ( .A1(n6002), .A2(n6092), .ZN(n5988) );
  AOI211_X1 U7051 ( .C1(n5990), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5989), 
        .B(n5988), .ZN(n5991) );
  OAI211_X1 U7052 ( .C1(n6096), .C2(n5993), .A(n5992), .B(n5991), .ZN(U2823)
         );
  AOI21_X1 U7053 ( .B1(n5995), .B2(EBX_REG_1__SCAN_IN), .A(n5994), .ZN(n6008)
         );
  INV_X1 U7054 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6005) );
  INV_X1 U7055 ( .A(n5996), .ZN(n5997) );
  AOI22_X1 U7056 ( .A1(n5998), .A2(REIP_REG_1__SCAN_IN), .B1(n4580), .B2(n5997), .ZN(n5999) );
  OAI21_X1 U7057 ( .B1(n6000), .B2(n6005), .A(n5999), .ZN(n6004) );
  NOR2_X1 U7058 ( .A1(n6002), .A2(n6001), .ZN(n6003) );
  AOI211_X1 U7059 ( .C1(n6006), .C2(n6005), .A(n6004), .B(n6003), .ZN(n6007)
         );
  OAI211_X1 U7060 ( .C1(n6010), .C2(n6009), .A(n6008), .B(n6007), .ZN(U2826)
         );
  AOI22_X1 U7061 ( .A1(n6012), .A2(n6023), .B1(n6022), .B2(n6011), .ZN(n6013)
         );
  OAI21_X1 U7062 ( .B1(n6014), .B2(n6026), .A(n6013), .ZN(U2846) );
  AOI22_X1 U7063 ( .A1(n6016), .A2(n6023), .B1(n6022), .B2(n6015), .ZN(n6017)
         );
  OAI21_X1 U7064 ( .B1(n6018), .B2(n6026), .A(n6017), .ZN(U2847) );
  AOI22_X1 U7065 ( .A1(n6084), .A2(n6023), .B1(n6022), .B2(n6139), .ZN(n6019)
         );
  OAI21_X1 U7066 ( .B1(n6745), .B2(n6026), .A(n6019), .ZN(U2853) );
  INV_X1 U7067 ( .A(n6020), .ZN(n6021) );
  AOI22_X1 U7068 ( .A1(n6024), .A2(n6023), .B1(n6022), .B2(n6021), .ZN(n6025)
         );
  OAI21_X1 U7069 ( .B1(n6027), .B2(n6026), .A(n6025), .ZN(U2858) );
  AOI22_X1 U7070 ( .A1(n6029), .A2(n6832), .B1(n6028), .B2(DATAI_17_), .ZN(
        n6032) );
  AOI22_X1 U7071 ( .A1(n6030), .A2(DATAI_1_), .B1(n6830), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7072 ( .A1(n6032), .A2(n6031), .ZN(U2874) );
  INV_X1 U7073 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n6713) );
  INV_X1 U7074 ( .A(n6033), .ZN(n6037) );
  AOI22_X1 U7075 ( .A1(n6037), .A2(EAX_REG_27__SCAN_IN), .B1(n6051), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n6034) );
  OAI21_X1 U7076 ( .B1(n6713), .B2(n6059), .A(n6034), .ZN(U2896) );
  INV_X1 U7077 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n6778) );
  AOI22_X1 U7078 ( .A1(n6037), .A2(EAX_REG_26__SCAN_IN), .B1(n6051), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6035) );
  OAI21_X1 U7079 ( .B1(n6778), .B2(n6059), .A(n6035), .ZN(U2897) );
  INV_X1 U7080 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n6671) );
  AOI22_X1 U7081 ( .A1(n6054), .A2(DATAO_REG_20__SCAN_IN), .B1(n6037), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6036) );
  OAI21_X1 U7082 ( .B1(n6671), .B2(n6590), .A(n6036), .ZN(U2903) );
  INV_X1 U7083 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n6789) );
  AOI22_X1 U7084 ( .A1(n6037), .A2(EAX_REG_18__SCAN_IN), .B1(n6051), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n6038) );
  OAI21_X1 U7085 ( .B1(n6789), .B2(n6059), .A(n6038), .ZN(U2905) );
  AOI22_X1 U7086 ( .A1(n6051), .A2(LWORD_REG_15__SCAN_IN), .B1(n6054), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6039) );
  OAI21_X1 U7087 ( .B1(n6040), .B2(n6060), .A(n6039), .ZN(U2908) );
  INV_X1 U7088 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6042) );
  AOI22_X1 U7089 ( .A1(n6051), .A2(LWORD_REG_14__SCAN_IN), .B1(n6054), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6041) );
  OAI21_X1 U7090 ( .B1(n6042), .B2(n6060), .A(n6041), .ZN(U2909) );
  INV_X1 U7091 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n6601) );
  AOI22_X1 U7092 ( .A1(EAX_REG_13__SCAN_IN), .A2(n6055), .B1(n6051), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n6043) );
  OAI21_X1 U7093 ( .B1(n6601), .B2(n6059), .A(n6043), .ZN(U2910) );
  AOI22_X1 U7094 ( .A1(n6051), .A2(LWORD_REG_12__SCAN_IN), .B1(n6054), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6044) );
  OAI21_X1 U7095 ( .B1(n6045), .B2(n6060), .A(n6044), .ZN(U2911) );
  AOI222_X1 U7096 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6051), .B1(n6055), .B2(
        EAX_REG_11__SCAN_IN), .C1(n6054), .C2(DATAO_REG_11__SCAN_IN), .ZN(
        n6046) );
  INV_X1 U7097 ( .A(n6046), .ZN(U2912) );
  INV_X1 U7098 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6048) );
  AOI22_X1 U7099 ( .A1(n6051), .A2(LWORD_REG_10__SCAN_IN), .B1(n6054), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6047) );
  OAI21_X1 U7100 ( .B1(n6048), .B2(n6060), .A(n6047), .ZN(U2913) );
  AOI22_X1 U7101 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n6051), .B1(n6054), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6049) );
  OAI21_X1 U7102 ( .B1(n6744), .B2(n6060), .A(n6049), .ZN(U2914) );
  AOI222_X1 U7103 ( .A1(LWORD_REG_8__SCAN_IN), .A2(n6051), .B1(n6055), .B2(
        EAX_REG_8__SCAN_IN), .C1(n6054), .C2(DATAO_REG_8__SCAN_IN), .ZN(n6050)
         );
  INV_X1 U7104 ( .A(n6050), .ZN(U2915) );
  INV_X1 U7105 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n6617) );
  INV_X1 U7106 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n6663) );
  OAI222_X1 U7107 ( .A1(n6059), .A2(n6617), .B1(n6060), .B2(n3582), .C1(n6663), 
        .C2(n6590), .ZN(U2916) );
  INV_X1 U7108 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n6669) );
  INV_X1 U7109 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n6754) );
  OAI222_X1 U7110 ( .A1(n6590), .A2(n6669), .B1(n6060), .B2(n3574), .C1(n6754), 
        .C2(n6059), .ZN(U2917) );
  AOI22_X1 U7111 ( .A1(n6051), .A2(LWORD_REG_5__SCAN_IN), .B1(n6054), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6052) );
  OAI21_X1 U7112 ( .B1(n3545), .B2(n6060), .A(n6052), .ZN(U2918) );
  INV_X1 U7113 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n6655) );
  AOI22_X1 U7114 ( .A1(EAX_REG_4__SCAN_IN), .A2(n6055), .B1(n6054), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6053) );
  OAI21_X1 U7115 ( .B1(n6655), .B2(n6590), .A(n6053), .ZN(U2919) );
  INV_X1 U7116 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n6725) );
  AOI22_X1 U7117 ( .A1(EAX_REG_3__SCAN_IN), .A2(n6055), .B1(n6054), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6056) );
  OAI21_X1 U7118 ( .B1(n6725), .B2(n6590), .A(n6056), .ZN(U2920) );
  INV_X1 U7119 ( .A(LWORD_REG_2__SCAN_IN), .ZN(n6677) );
  INV_X1 U7120 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n6609) );
  OAI222_X1 U7121 ( .A1(n6590), .A2(n6677), .B1(n6060), .B2(n6057), .C1(n6609), 
        .C2(n6059), .ZN(U2921) );
  INV_X1 U7122 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n6700) );
  INV_X1 U7123 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6058) );
  INV_X1 U7124 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n6660) );
  OAI222_X1 U7125 ( .A1(n6059), .A2(n6700), .B1(n6060), .B2(n6058), .C1(n6660), 
        .C2(n6590), .ZN(U2922) );
  INV_X1 U7126 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n6598) );
  INV_X1 U7127 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n6684) );
  OAI222_X1 U7128 ( .A1(n6590), .A2(n6598), .B1(n6060), .B2(n6696), .C1(n6684), 
        .C2(n6059), .ZN(U2923) );
  AOI22_X1 U7129 ( .A1(UWORD_REG_10__SCAN_IN), .A2(n6061), .B1(n6069), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7130 ( .A1(n6063), .A2(DATAI_10_), .ZN(n6065) );
  NAND2_X1 U7131 ( .A1(n6062), .A2(n6065), .ZN(U2934) );
  AOI22_X1 U7132 ( .A1(UWORD_REG_11__SCAN_IN), .A2(n6070), .B1(n6069), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7133 ( .A1(n6063), .A2(DATAI_11_), .ZN(n6067) );
  NAND2_X1 U7134 ( .A1(n6064), .A2(n6067), .ZN(U2935) );
  AOI22_X1 U7135 ( .A1(LWORD_REG_10__SCAN_IN), .A2(n6070), .B1(n6069), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U7136 ( .A1(n6066), .A2(n6065), .ZN(U2949) );
  AOI22_X1 U7137 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6070), .B1(n6069), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7138 ( .A1(n6068), .A2(n6067), .ZN(U2950) );
  AOI22_X1 U7139 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n6070), .B1(n6069), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7140 ( .A1(n6072), .A2(n6071), .ZN(U2952) );
  AOI22_X1 U7141 ( .A1(n6156), .A2(REIP_REG_11__SCAN_IN), .B1(n6097), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6077) );
  AOI22_X1 U7142 ( .A1(n6075), .A2(n6101), .B1(n6074), .B2(n6073), .ZN(n6076)
         );
  OAI211_X1 U7143 ( .C1(n6079), .C2(n6078), .A(n6077), .B(n6076), .ZN(U2975)
         );
  AOI22_X1 U7144 ( .A1(n6156), .A2(REIP_REG_6__SCAN_IN), .B1(n6097), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6086) );
  OAI21_X1 U7145 ( .B1(n6082), .B2(n6081), .A(n6080), .ZN(n6083) );
  INV_X1 U7146 ( .A(n6083), .ZN(n6141) );
  AOI22_X1 U7147 ( .A1(n6141), .A2(n6104), .B1(n6101), .B2(n6084), .ZN(n6085)
         );
  OAI211_X1 U7148 ( .C1(n6108), .C2(n6087), .A(n6086), .B(n6085), .ZN(U2980)
         );
  AOI22_X1 U7149 ( .A1(n6156), .A2(REIP_REG_4__SCAN_IN), .B1(n6097), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6095) );
  OAI21_X1 U7150 ( .B1(n6090), .B2(n6089), .A(n6088), .ZN(n6091) );
  INV_X1 U7151 ( .A(n6091), .ZN(n6158) );
  INV_X1 U7152 ( .A(n6092), .ZN(n6093) );
  AOI22_X1 U7153 ( .A1(n6158), .A2(n6104), .B1(n6101), .B2(n6093), .ZN(n6094)
         );
  OAI211_X1 U7154 ( .C1(n6108), .C2(n6096), .A(n6095), .B(n6094), .ZN(U2982)
         );
  AOI22_X1 U7155 ( .A1(n6156), .A2(REIP_REG_2__SCAN_IN), .B1(n6097), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6106) );
  XNOR2_X1 U7156 ( .A(n6098), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6100)
         );
  XNOR2_X1 U7157 ( .A(n6100), .B(n6099), .ZN(n6185) );
  INV_X1 U7158 ( .A(n6185), .ZN(n6103) );
  AOI22_X1 U7159 ( .A1(n6104), .A2(n6103), .B1(n6102), .B2(n6101), .ZN(n6105)
         );
  OAI211_X1 U7160 ( .C1(n6108), .C2(n6107), .A(n6106), .B(n6105), .ZN(U2984)
         );
  AOI21_X1 U7161 ( .B1(n6174), .B2(n6110), .A(n6109), .ZN(n6117) );
  AOI22_X1 U7162 ( .A1(n6112), .A2(n6167), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6111), .ZN(n6116) );
  OAI211_X1 U7163 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6114), .B(n6113), .ZN(n6115) );
  NAND3_X1 U7164 ( .A1(n6117), .A2(n6116), .A3(n6115), .ZN(U3008) );
  AOI21_X1 U7165 ( .B1(n6174), .B2(n6119), .A(n6118), .ZN(n6124) );
  AOI211_X1 U7166 ( .C1(n6132), .C2(n6739), .A(n6120), .B(n6133), .ZN(n6121)
         );
  AOI21_X1 U7167 ( .B1(n6122), .B2(n6167), .A(n6121), .ZN(n6123) );
  OAI211_X1 U7168 ( .C1(n6131), .C2(n6739), .A(n6124), .B(n6123), .ZN(U3010)
         );
  OAI222_X1 U7169 ( .A1(n6128), .A2(n6127), .B1(n6190), .B2(n6126), .C1(n6184), 
        .C2(n6125), .ZN(n6129) );
  INV_X1 U7170 ( .A(n6129), .ZN(n6130) );
  OAI221_X1 U7171 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n6133), .C1(n6132), .C2(n6131), .A(n6130), .ZN(U3011) );
  OAI21_X1 U7172 ( .B1(n6136), .B2(n6135), .A(n6134), .ZN(n6176) );
  AOI21_X1 U7173 ( .B1(n6138), .B2(n6137), .A(n6176), .ZN(n6155) );
  AOI22_X1 U7174 ( .A1(n6174), .A2(n6139), .B1(n6156), .B2(REIP_REG_6__SCAN_IN), .ZN(n6143) );
  AOI22_X1 U7175 ( .A1(n6141), .A2(n6167), .B1(n6140), .B2(n6144), .ZN(n6142)
         );
  OAI211_X1 U7176 ( .C1(n6155), .C2(n6144), .A(n6143), .B(n6142), .ZN(U3012)
         );
  OAI21_X1 U7177 ( .B1(n6179), .B2(n6146), .A(n6145), .ZN(n6147) );
  AOI21_X1 U7178 ( .B1(n6178), .B2(n6148), .A(n6147), .ZN(n6154) );
  INV_X1 U7179 ( .A(n6149), .ZN(n6151) );
  AOI22_X1 U7180 ( .A1(n6151), .A2(n6167), .B1(n6174), .B2(n6150), .ZN(n6153)
         );
  NAND2_X1 U7181 ( .A1(n6156), .A2(REIP_REG_5__SCAN_IN), .ZN(n6152) );
  OAI211_X1 U7182 ( .C1(n6155), .C2(n6154), .A(n6153), .B(n6152), .ZN(U3013)
         );
  AOI21_X1 U7183 ( .B1(n6178), .B2(n6175), .A(n6176), .ZN(n6172) );
  AOI22_X1 U7184 ( .A1(n6174), .A2(n6157), .B1(n6156), .B2(REIP_REG_4__SCAN_IN), .ZN(n6162) );
  AOI211_X1 U7185 ( .C1(n4205), .C2(n6163), .A(n6175), .B(n6166), .ZN(n6160)
         );
  AOI22_X1 U7186 ( .A1(n6160), .A2(n6159), .B1(n6167), .B2(n6158), .ZN(n6161)
         );
  OAI211_X1 U7187 ( .C1(n6172), .C2(n6163), .A(n6162), .B(n6161), .ZN(U3014)
         );
  AOI21_X1 U7188 ( .B1(n6174), .B2(n6165), .A(n6164), .ZN(n6171) );
  NOR2_X1 U7189 ( .A1(n6175), .A2(n6166), .ZN(n6169) );
  AOI22_X1 U7190 ( .A1(n6169), .A2(n4205), .B1(n6168), .B2(n6167), .ZN(n6170)
         );
  OAI211_X1 U7191 ( .C1(n6172), .C2(n4205), .A(n6171), .B(n6170), .ZN(U3015)
         );
  AOI22_X1 U7192 ( .A1(n6178), .A2(n6175), .B1(n6174), .B2(n6173), .ZN(n6189)
         );
  AOI21_X1 U7194 ( .B1(n6178), .B2(n6177), .A(n6176), .ZN(n6182) );
  OAI33_X1 U7195 ( .A1(1'b0), .A2(n6182), .A3(n6181), .B1(
        INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6180), .B3(n6179), .ZN(n6187) );
  NOR2_X1 U7196 ( .A1(n6185), .A2(n6184), .ZN(n6186) );
  NOR2_X1 U7197 ( .A1(n6187), .A2(n6186), .ZN(n6188) );
  OAI211_X1 U7198 ( .C1(n6190), .C2(n6698), .A(n6189), .B(n6188), .ZN(U3016)
         );
  AND2_X1 U7199 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6191), .ZN(U3019)
         );
  INV_X1 U7200 ( .A(n6192), .ZN(n6261) );
  NAND3_X1 U7201 ( .A1(n6340), .A2(n6339), .A3(n6460), .ZN(n6193) );
  OAI21_X1 U7202 ( .B1(n6261), .B2(n6194), .A(n6193), .ZN(n6216) );
  NOR2_X1 U7203 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6195), .ZN(n6215)
         );
  AOI22_X1 U7204 ( .A1(n6344), .A2(n6216), .B1(n6388), .B2(n6215), .ZN(n6202)
         );
  OAI21_X1 U7205 ( .B1(n6217), .B2(n6197), .A(n6265), .ZN(n6199) );
  AOI21_X1 U7206 ( .B1(n6199), .B2(n6198), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n6200) );
  NOR2_X1 U7207 ( .A1(n6258), .A2(n6269), .ZN(n6336) );
  AOI22_X1 U7208 ( .A1(n6218), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n6397), 
        .B2(n6217), .ZN(n6201) );
  OAI211_X1 U7209 ( .C1(n6272), .C2(n6221), .A(n6202), .B(n6201), .ZN(U3036)
         );
  AOI22_X1 U7210 ( .A1(n6347), .A2(n6216), .B1(n6401), .B2(n6215), .ZN(n6204)
         );
  AOI22_X1 U7211 ( .A1(n6218), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n6402), 
        .B2(n6217), .ZN(n6203) );
  OAI211_X1 U7212 ( .C1(n6221), .C2(n6275), .A(n6204), .B(n6203), .ZN(U3037)
         );
  AOI22_X1 U7213 ( .A1(n6351), .A2(n6216), .B1(n6407), .B2(n6215), .ZN(n6206)
         );
  AOI22_X1 U7214 ( .A1(n6218), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n6409), 
        .B2(n6217), .ZN(n6205) );
  OAI211_X1 U7215 ( .C1(n6221), .C2(n6278), .A(n6206), .B(n6205), .ZN(U3038)
         );
  AOI22_X1 U7216 ( .A1(n6355), .A2(n6216), .B1(n6413), .B2(n6215), .ZN(n6208)
         );
  AOI22_X1 U7217 ( .A1(n6218), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n6414), 
        .B2(n6217), .ZN(n6207) );
  OAI211_X1 U7218 ( .C1(n6221), .C2(n6281), .A(n6208), .B(n6207), .ZN(U3039)
         );
  AOI22_X1 U7219 ( .A1(n6359), .A2(n6216), .B1(n6419), .B2(n6215), .ZN(n6210)
         );
  AOI22_X1 U7220 ( .A1(n6218), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n6420), 
        .B2(n6217), .ZN(n6209) );
  OAI211_X1 U7221 ( .C1(n6221), .C2(n6284), .A(n6210), .B(n6209), .ZN(U3040)
         );
  AOI22_X1 U7222 ( .A1(n6363), .A2(n6216), .B1(n6425), .B2(n6215), .ZN(n6212)
         );
  AOI22_X1 U7223 ( .A1(n6218), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n6426), 
        .B2(n6217), .ZN(n6211) );
  OAI211_X1 U7224 ( .C1(n6221), .C2(n6287), .A(n6212), .B(n6211), .ZN(U3041)
         );
  AOI22_X1 U7225 ( .A1(n6367), .A2(n6216), .B1(n6431), .B2(n6215), .ZN(n6214)
         );
  AOI22_X1 U7226 ( .A1(n6218), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n6432), 
        .B2(n6217), .ZN(n6213) );
  OAI211_X1 U7227 ( .C1(n6221), .C2(n6290), .A(n6214), .B(n6213), .ZN(U3042)
         );
  AOI22_X1 U7228 ( .A1(n6373), .A2(n6216), .B1(n6438), .B2(n6215), .ZN(n6220)
         );
  AOI22_X1 U7229 ( .A1(n6218), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n6442), 
        .B2(n6217), .ZN(n6219) );
  OAI211_X1 U7230 ( .C1(n6221), .C2(n6297), .A(n6220), .B(n6219), .ZN(U3043)
         );
  INV_X1 U7231 ( .A(n6222), .ZN(n6223) );
  NOR2_X1 U7232 ( .A1(n6451), .A2(n6228), .ZN(n6249) );
  AOI21_X1 U7233 ( .B1(n6223), .B2(n3102), .A(n6249), .ZN(n6229) );
  INV_X1 U7234 ( .A(n6229), .ZN(n6224) );
  OAI21_X1 U7235 ( .B1(n6230), .B2(n6224), .A(n6306), .ZN(n6225) );
  INV_X1 U7236 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n6690) );
  OR2_X1 U7237 ( .A1(n6227), .A2(n6226), .ZN(n6262) );
  AOI22_X1 U7238 ( .A1(n6389), .A2(n6293), .B1(n6388), .B2(n6249), .ZN(n6233)
         );
  OAI22_X1 U7239 ( .A1(n6230), .A2(n6229), .B1(n6228), .B2(n6583), .ZN(n6251)
         );
  AOI22_X1 U7240 ( .A1(n6251), .A2(n6344), .B1(n6397), .B2(n6250), .ZN(n6232)
         );
  OAI211_X1 U7241 ( .C1(n6255), .C2(n6690), .A(n6233), .B(n6232), .ZN(U3060)
         );
  INV_X1 U7242 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6236) );
  AOI22_X1 U7243 ( .A1(n6403), .A2(n6293), .B1(n6401), .B2(n6249), .ZN(n6235)
         );
  AOI22_X1 U7244 ( .A1(n6251), .A2(n6347), .B1(n6402), .B2(n6250), .ZN(n6234)
         );
  OAI211_X1 U7245 ( .C1(n6255), .C2(n6236), .A(n6235), .B(n6234), .ZN(U3061)
         );
  INV_X1 U7246 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6239) );
  AOI22_X1 U7247 ( .A1(n6408), .A2(n6293), .B1(n6407), .B2(n6249), .ZN(n6238)
         );
  AOI22_X1 U7248 ( .A1(n6251), .A2(n6351), .B1(n6409), .B2(n6250), .ZN(n6237)
         );
  OAI211_X1 U7249 ( .C1(n6255), .C2(n6239), .A(n6238), .B(n6237), .ZN(U3062)
         );
  INV_X1 U7250 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n6242) );
  AOI22_X1 U7251 ( .A1(n6415), .A2(n6293), .B1(n6413), .B2(n6249), .ZN(n6241)
         );
  AOI22_X1 U7252 ( .A1(n6251), .A2(n6355), .B1(n6414), .B2(n6250), .ZN(n6240)
         );
  OAI211_X1 U7253 ( .C1(n6255), .C2(n6242), .A(n6241), .B(n6240), .ZN(U3063)
         );
  INV_X1 U7254 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n6638) );
  AOI22_X1 U7255 ( .A1(n6421), .A2(n6293), .B1(n6419), .B2(n6249), .ZN(n6244)
         );
  AOI22_X1 U7256 ( .A1(n6251), .A2(n6359), .B1(n6420), .B2(n6250), .ZN(n6243)
         );
  OAI211_X1 U7257 ( .C1(n6255), .C2(n6638), .A(n6244), .B(n6243), .ZN(U3064)
         );
  AOI22_X1 U7258 ( .A1(n6427), .A2(n6293), .B1(n6425), .B2(n6249), .ZN(n6246)
         );
  AOI22_X1 U7259 ( .A1(n6251), .A2(n6363), .B1(n6426), .B2(n6250), .ZN(n6245)
         );
  OAI211_X1 U7260 ( .C1(n6255), .C2(n6843), .A(n6246), .B(n6245), .ZN(U3065)
         );
  INV_X1 U7261 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6659) );
  AOI22_X1 U7262 ( .A1(n6433), .A2(n6293), .B1(n6431), .B2(n6249), .ZN(n6248)
         );
  AOI22_X1 U7263 ( .A1(n6251), .A2(n6367), .B1(n6432), .B2(n6250), .ZN(n6247)
         );
  OAI211_X1 U7264 ( .C1(n6255), .C2(n6659), .A(n6248), .B(n6247), .ZN(U3066)
         );
  INV_X1 U7265 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n6254) );
  AOI22_X1 U7266 ( .A1(n6439), .A2(n6293), .B1(n6438), .B2(n6249), .ZN(n6253)
         );
  AOI22_X1 U7267 ( .A1(n6251), .A2(n6373), .B1(n6442), .B2(n6250), .ZN(n6252)
         );
  OAI211_X1 U7268 ( .C1(n6255), .C2(n6254), .A(n6253), .B(n6252), .ZN(U3067)
         );
  INV_X1 U7269 ( .A(n6264), .ZN(n6260) );
  NAND3_X1 U7270 ( .A1(n6258), .A2(n6339), .A3(n6460), .ZN(n6259) );
  OAI21_X1 U7271 ( .B1(n6261), .B2(n6260), .A(n6259), .ZN(n6292) );
  AND2_X1 U7272 ( .A1(n6451), .A2(n6307), .ZN(n6291) );
  AOI22_X1 U7273 ( .A1(n6344), .A2(n6292), .B1(n6388), .B2(n6291), .ZN(n6271)
         );
  NAND3_X1 U7274 ( .A1(n6262), .A2(n6380), .A3(n6302), .ZN(n6266) );
  AND2_X1 U7275 ( .A1(n6264), .A2(n6263), .ZN(n6300) );
  AOI21_X1 U7276 ( .B1(n6266), .B2(n6265), .A(n6300), .ZN(n6268) );
  OAI21_X1 U7277 ( .B1(n6688), .B2(n6291), .A(n6460), .ZN(n6267) );
  AOI22_X1 U7278 ( .A1(n6294), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6397), 
        .B2(n6293), .ZN(n6270) );
  OAI211_X1 U7279 ( .C1(n6272), .C2(n6302), .A(n6271), .B(n6270), .ZN(U3068)
         );
  AOI22_X1 U7280 ( .A1(n6347), .A2(n6292), .B1(n6401), .B2(n6291), .ZN(n6274)
         );
  AOI22_X1 U7281 ( .A1(n6294), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6402), 
        .B2(n6293), .ZN(n6273) );
  OAI211_X1 U7282 ( .C1(n6275), .C2(n6302), .A(n6274), .B(n6273), .ZN(U3069)
         );
  AOI22_X1 U7283 ( .A1(n6351), .A2(n6292), .B1(n6407), .B2(n6291), .ZN(n6277)
         );
  AOI22_X1 U7284 ( .A1(n6294), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6409), 
        .B2(n6293), .ZN(n6276) );
  OAI211_X1 U7285 ( .C1(n6278), .C2(n6302), .A(n6277), .B(n6276), .ZN(U3070)
         );
  AOI22_X1 U7286 ( .A1(n6355), .A2(n6292), .B1(n6413), .B2(n6291), .ZN(n6280)
         );
  AOI22_X1 U7287 ( .A1(n6294), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6414), 
        .B2(n6293), .ZN(n6279) );
  OAI211_X1 U7288 ( .C1(n6281), .C2(n6302), .A(n6280), .B(n6279), .ZN(U3071)
         );
  AOI22_X1 U7289 ( .A1(n6359), .A2(n6292), .B1(n6419), .B2(n6291), .ZN(n6283)
         );
  AOI22_X1 U7290 ( .A1(n6294), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6420), 
        .B2(n6293), .ZN(n6282) );
  OAI211_X1 U7291 ( .C1(n6284), .C2(n6302), .A(n6283), .B(n6282), .ZN(U3072)
         );
  AOI22_X1 U7292 ( .A1(n6363), .A2(n6292), .B1(n6425), .B2(n6291), .ZN(n6286)
         );
  AOI22_X1 U7293 ( .A1(n6294), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6426), 
        .B2(n6293), .ZN(n6285) );
  OAI211_X1 U7294 ( .C1(n6287), .C2(n6302), .A(n6286), .B(n6285), .ZN(U3073)
         );
  AOI22_X1 U7295 ( .A1(n6367), .A2(n6292), .B1(n6431), .B2(n6291), .ZN(n6289)
         );
  AOI22_X1 U7296 ( .A1(n6294), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6432), 
        .B2(n6293), .ZN(n6288) );
  OAI211_X1 U7297 ( .C1(n6290), .C2(n6302), .A(n6289), .B(n6288), .ZN(U3074)
         );
  AOI22_X1 U7298 ( .A1(n6373), .A2(n6292), .B1(n6438), .B2(n6291), .ZN(n6296)
         );
  AOI22_X1 U7299 ( .A1(n6294), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6442), 
        .B2(n6293), .ZN(n6295) );
  OAI211_X1 U7300 ( .C1(n6297), .C2(n6302), .A(n6296), .B(n6295), .ZN(U3075)
         );
  AND2_X1 U7301 ( .A1(n6298), .A2(n6380), .ZN(n6304) );
  INV_X1 U7302 ( .A(n6299), .ZN(n6323) );
  AOI21_X1 U7303 ( .B1(n6300), .B2(n3102), .A(n6323), .ZN(n6303) );
  INV_X1 U7304 ( .A(n6303), .ZN(n6301) );
  AOI22_X1 U7305 ( .A1(n6304), .A2(n6301), .B1(n6307), .B2(
        STATE2_REG_2__SCAN_IN), .ZN(n6328) );
  AOI22_X1 U7306 ( .A1(n6388), .A2(n6323), .B1(n6324), .B2(n6397), .ZN(n6309)
         );
  NAND2_X1 U7307 ( .A1(n6304), .A2(n6303), .ZN(n6305) );
  OAI211_X1 U7308 ( .C1(n6307), .C2(n6380), .A(n6306), .B(n6305), .ZN(n6325)
         );
  AOI22_X1 U7309 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6325), .B1(n6389), 
        .B2(n6322), .ZN(n6308) );
  OAI211_X1 U7310 ( .C1(n6328), .C2(n6400), .A(n6309), .B(n6308), .ZN(U3076)
         );
  AOI22_X1 U7311 ( .A1(n6401), .A2(n6323), .B1(n6324), .B2(n6402), .ZN(n6311)
         );
  AOI22_X1 U7312 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6325), .B1(n6403), 
        .B2(n6322), .ZN(n6310) );
  OAI211_X1 U7313 ( .C1(n6328), .C2(n6406), .A(n6311), .B(n6310), .ZN(U3077)
         );
  AOI22_X1 U7314 ( .A1(n6407), .A2(n6323), .B1(n6408), .B2(n6322), .ZN(n6313)
         );
  AOI22_X1 U7315 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6325), .B1(n6409), 
        .B2(n6324), .ZN(n6312) );
  OAI211_X1 U7316 ( .C1(n6328), .C2(n6412), .A(n6313), .B(n6312), .ZN(U3078)
         );
  AOI22_X1 U7317 ( .A1(n6413), .A2(n6323), .B1(n6415), .B2(n6322), .ZN(n6315)
         );
  AOI22_X1 U7318 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6325), .B1(n6414), 
        .B2(n6324), .ZN(n6314) );
  OAI211_X1 U7319 ( .C1(n6328), .C2(n6418), .A(n6315), .B(n6314), .ZN(U3079)
         );
  AOI22_X1 U7320 ( .A1(n6419), .A2(n6323), .B1(n6421), .B2(n6322), .ZN(n6317)
         );
  AOI22_X1 U7321 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6325), .B1(n6420), 
        .B2(n6324), .ZN(n6316) );
  OAI211_X1 U7322 ( .C1(n6328), .C2(n6424), .A(n6317), .B(n6316), .ZN(U3080)
         );
  AOI22_X1 U7323 ( .A1(n6425), .A2(n6323), .B1(n6427), .B2(n6322), .ZN(n6319)
         );
  AOI22_X1 U7324 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6325), .B1(n6426), 
        .B2(n6324), .ZN(n6318) );
  OAI211_X1 U7325 ( .C1(n6328), .C2(n6430), .A(n6319), .B(n6318), .ZN(U3081)
         );
  AOI22_X1 U7326 ( .A1(n6431), .A2(n6323), .B1(n6433), .B2(n6322), .ZN(n6321)
         );
  AOI22_X1 U7327 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6325), .B1(n6432), 
        .B2(n6324), .ZN(n6320) );
  OAI211_X1 U7328 ( .C1(n6328), .C2(n6436), .A(n6321), .B(n6320), .ZN(U3082)
         );
  AOI22_X1 U7329 ( .A1(n6438), .A2(n6323), .B1(n6439), .B2(n6322), .ZN(n6327)
         );
  AOI22_X1 U7330 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6325), .B1(n6442), 
        .B2(n6324), .ZN(n6326) );
  OAI211_X1 U7331 ( .C1(n6328), .C2(n6446), .A(n6327), .B(n6326), .ZN(U3083)
         );
  NOR2_X2 U7332 ( .A1(n6330), .A2(n6329), .ZN(n6441) );
  NOR3_X1 U7333 ( .A1(n6441), .A2(n6372), .A3(n6393), .ZN(n6332) );
  NOR2_X1 U7334 ( .A1(n6332), .A2(n6331), .ZN(n6343) );
  INV_X1 U7335 ( .A(n6343), .ZN(n6338) );
  NAND2_X1 U7336 ( .A1(n6383), .A2(n3101), .ZN(n6342) );
  NAND3_X1 U7337 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6334), .ZN(n6392) );
  NOR2_X1 U7338 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6392), .ZN(n6371)
         );
  OAI211_X1 U7339 ( .C1(n6371), .C2(n6688), .A(n6336), .B(n6335), .ZN(n6337)
         );
  INV_X1 U7340 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n6629) );
  AOI22_X1 U7341 ( .A1(n6441), .A2(n6389), .B1(n6388), .B2(n6371), .ZN(n6346)
         );
  NAND3_X1 U7342 ( .A1(n6340), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6339), .ZN(n6341) );
  OAI21_X1 U7343 ( .B1(n6343), .B2(n6342), .A(n6341), .ZN(n6374) );
  AOI22_X1 U7344 ( .A1(n6374), .A2(n6344), .B1(n6397), .B2(n6372), .ZN(n6345)
         );
  OAI211_X1 U7345 ( .C1(n6377), .C2(n6629), .A(n6346), .B(n6345), .ZN(U3100)
         );
  INV_X1 U7346 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n6350) );
  AOI22_X1 U7347 ( .A1(n6441), .A2(n6403), .B1(n6401), .B2(n6371), .ZN(n6349)
         );
  AOI22_X1 U7348 ( .A1(n6374), .A2(n6347), .B1(n6372), .B2(n6402), .ZN(n6348)
         );
  OAI211_X1 U7349 ( .C1(n6377), .C2(n6350), .A(n6349), .B(n6348), .ZN(U3101)
         );
  INV_X1 U7350 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n6354) );
  AOI22_X1 U7351 ( .A1(n6441), .A2(n6408), .B1(n6407), .B2(n6371), .ZN(n6353)
         );
  AOI22_X1 U7352 ( .A1(n6374), .A2(n6351), .B1(n6372), .B2(n6409), .ZN(n6352)
         );
  OAI211_X1 U7353 ( .C1(n6377), .C2(n6354), .A(n6353), .B(n6352), .ZN(U3102)
         );
  INV_X1 U7354 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6358) );
  AOI22_X1 U7355 ( .A1(n6441), .A2(n6415), .B1(n6413), .B2(n6371), .ZN(n6357)
         );
  AOI22_X1 U7356 ( .A1(n6374), .A2(n6355), .B1(n6372), .B2(n6414), .ZN(n6356)
         );
  OAI211_X1 U7357 ( .C1(n6377), .C2(n6358), .A(n6357), .B(n6356), .ZN(U3103)
         );
  INV_X1 U7358 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n6362) );
  AOI22_X1 U7359 ( .A1(n6441), .A2(n6421), .B1(n6419), .B2(n6371), .ZN(n6361)
         );
  AOI22_X1 U7360 ( .A1(n6374), .A2(n6359), .B1(n6372), .B2(n6420), .ZN(n6360)
         );
  OAI211_X1 U7361 ( .C1(n6377), .C2(n6362), .A(n6361), .B(n6360), .ZN(U3104)
         );
  INV_X1 U7362 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n6366) );
  AOI22_X1 U7363 ( .A1(n6441), .A2(n6427), .B1(n6425), .B2(n6371), .ZN(n6365)
         );
  AOI22_X1 U7364 ( .A1(n6374), .A2(n6363), .B1(n6372), .B2(n6426), .ZN(n6364)
         );
  OAI211_X1 U7365 ( .C1(n6377), .C2(n6366), .A(n6365), .B(n6364), .ZN(U3105)
         );
  INV_X1 U7366 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6370) );
  AOI22_X1 U7367 ( .A1(n6441), .A2(n6433), .B1(n6431), .B2(n6371), .ZN(n6369)
         );
  AOI22_X1 U7368 ( .A1(n6374), .A2(n6367), .B1(n6372), .B2(n6432), .ZN(n6368)
         );
  OAI211_X1 U7369 ( .C1(n6377), .C2(n6370), .A(n6369), .B(n6368), .ZN(U3106)
         );
  INV_X1 U7370 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n6838) );
  AOI22_X1 U7371 ( .A1(n6441), .A2(n6439), .B1(n6438), .B2(n6371), .ZN(n6376)
         );
  AOI22_X1 U7372 ( .A1(n6374), .A2(n6373), .B1(n6372), .B2(n6442), .ZN(n6375)
         );
  OAI211_X1 U7373 ( .C1(n6377), .C2(n6838), .A(n6376), .B(n6375), .ZN(U3107)
         );
  NAND2_X1 U7374 ( .A1(n6379), .A2(n6378), .ZN(n6381) );
  NAND2_X1 U7375 ( .A1(n6381), .A2(n6380), .ZN(n6396) );
  NOR2_X1 U7376 ( .A1(n6382), .A2(n6460), .ZN(n6437) );
  AOI21_X1 U7377 ( .B1(n6384), .B2(n6383), .A(n6437), .ZN(n6390) );
  OR2_X1 U7378 ( .A1(n6396), .A2(n6390), .ZN(n6387) );
  INV_X1 U7379 ( .A(n6392), .ZN(n6385) );
  NAND2_X1 U7380 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6385), .ZN(n6386) );
  AOI22_X1 U7381 ( .A1(n6440), .A2(n6389), .B1(n6388), .B2(n6437), .ZN(n6399)
         );
  INV_X1 U7382 ( .A(n6390), .ZN(n6395) );
  AOI21_X1 U7383 ( .B1(n6393), .B2(n6392), .A(n6391), .ZN(n6394) );
  OAI21_X1 U7384 ( .B1(n6396), .B2(n6395), .A(n6394), .ZN(n6443) );
  AOI22_X1 U7385 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6443), .B1(n6397), 
        .B2(n6441), .ZN(n6398) );
  OAI211_X1 U7386 ( .C1(n6447), .C2(n6400), .A(n6399), .B(n6398), .ZN(U3108)
         );
  AOI22_X1 U7387 ( .A1(n6441), .A2(n6402), .B1(n6401), .B2(n6437), .ZN(n6405)
         );
  AOI22_X1 U7388 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6443), .B1(n6403), 
        .B2(n6440), .ZN(n6404) );
  OAI211_X1 U7389 ( .C1(n6447), .C2(n6406), .A(n6405), .B(n6404), .ZN(U3109)
         );
  AOI22_X1 U7390 ( .A1(n6440), .A2(n6408), .B1(n6407), .B2(n6437), .ZN(n6411)
         );
  AOI22_X1 U7391 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6443), .B1(n6409), 
        .B2(n6441), .ZN(n6410) );
  OAI211_X1 U7392 ( .C1(n6447), .C2(n6412), .A(n6411), .B(n6410), .ZN(U3110)
         );
  AOI22_X1 U7393 ( .A1(n6441), .A2(n6414), .B1(n6413), .B2(n6437), .ZN(n6417)
         );
  AOI22_X1 U7394 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6443), .B1(n6415), 
        .B2(n6440), .ZN(n6416) );
  OAI211_X1 U7395 ( .C1(n6447), .C2(n6418), .A(n6417), .B(n6416), .ZN(U3111)
         );
  AOI22_X1 U7396 ( .A1(n6441), .A2(n6420), .B1(n6419), .B2(n6437), .ZN(n6423)
         );
  AOI22_X1 U7397 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6443), .B1(n6421), 
        .B2(n6440), .ZN(n6422) );
  OAI211_X1 U7398 ( .C1(n6447), .C2(n6424), .A(n6423), .B(n6422), .ZN(U3112)
         );
  AOI22_X1 U7399 ( .A1(n6441), .A2(n6426), .B1(n6425), .B2(n6437), .ZN(n6429)
         );
  AOI22_X1 U7400 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6443), .B1(n6427), 
        .B2(n6440), .ZN(n6428) );
  OAI211_X1 U7401 ( .C1(n6447), .C2(n6430), .A(n6429), .B(n6428), .ZN(U3113)
         );
  AOI22_X1 U7402 ( .A1(n6441), .A2(n6432), .B1(n6431), .B2(n6437), .ZN(n6435)
         );
  AOI22_X1 U7403 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6443), .B1(n6433), 
        .B2(n6440), .ZN(n6434) );
  OAI211_X1 U7404 ( .C1(n6447), .C2(n6436), .A(n6435), .B(n6434), .ZN(U3114)
         );
  AOI22_X1 U7405 ( .A1(n6440), .A2(n6439), .B1(n6438), .B2(n6437), .ZN(n6445)
         );
  AOI22_X1 U7406 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6443), .B1(n6442), 
        .B2(n6441), .ZN(n6444) );
  OAI211_X1 U7407 ( .C1(n6447), .C2(n6446), .A(n6445), .B(n6444), .ZN(U3115)
         );
  OR2_X1 U7408 ( .A1(n6449), .A2(n6448), .ZN(n6454) );
  INV_X1 U7409 ( .A(n6454), .ZN(n6457) );
  AOI211_X1 U7410 ( .C1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n6452), .A(n6451), .B(n6450), .ZN(n6453) );
  OAI21_X1 U7411 ( .B1(n6454), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6453), 
        .ZN(n6455) );
  OAI21_X1 U7412 ( .B1(n6457), .B2(n6456), .A(n6455), .ZN(n6458) );
  AOI222_X1 U7413 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6459), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6458), .C1(n6459), .C2(n6458), 
        .ZN(n6461) );
  AOI222_X1 U7414 ( .A1(n6462), .A2(n6461), .B1(n6462), .B2(n6460), .C1(n6461), 
        .C2(n6460), .ZN(n6463) );
  OR2_X1 U7415 ( .A1(n6463), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6472)
         );
  NOR2_X1 U7416 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6467) );
  INV_X1 U7417 ( .A(n6464), .ZN(n6465) );
  OAI211_X1 U7418 ( .C1(n6468), .C2(n6467), .A(n6466), .B(n6465), .ZN(n6469)
         );
  NOR2_X1 U7419 ( .A1(n6470), .A2(n6469), .ZN(n6471) );
  NAND2_X1 U7420 ( .A1(n6472), .A2(n6471), .ZN(n6480) );
  OAI22_X1 U7421 ( .A1(n6480), .A2(n6485), .B1(n6506), .B2(n6590), .ZN(n6476)
         );
  OR2_X1 U7422 ( .A1(n6474), .A2(n6473), .ZN(n6475) );
  AOI21_X1 U7423 ( .B1(READY_N), .B2(n6583), .A(n6484), .ZN(n6491) );
  AOI211_X1 U7424 ( .C1(n6495), .C2(n6477), .A(STATE2_REG_0__SCAN_IN), .B(
        n6484), .ZN(n6478) );
  AOI211_X1 U7425 ( .C1(n6481), .C2(n6480), .A(n6479), .B(n6478), .ZN(n6482)
         );
  OAI221_X1 U7426 ( .B1(n6586), .B2(n6491), .C1(n6586), .C2(n6483), .A(n6482), 
        .ZN(U3148) );
  NAND2_X1 U7427 ( .A1(n6492), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6490) );
  INV_X1 U7428 ( .A(n6484), .ZN(n6563) );
  OAI21_X1 U7429 ( .B1(READY_N), .B2(n6486), .A(n6485), .ZN(n6488) );
  AOI21_X1 U7430 ( .B1(n6563), .B2(n6488), .A(n6487), .ZN(n6489) );
  OAI21_X1 U7431 ( .B1(n6491), .B2(n6490), .A(n6489), .ZN(U3149) );
  OAI211_X1 U7432 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6506), .A(n6561), .B(
        n6492), .ZN(n6494) );
  OAI21_X1 U7433 ( .B1(n6495), .B2(n6494), .A(n6493), .ZN(U3150) );
  INV_X1 U7434 ( .A(DATAWIDTH_REG_31__SCAN_IN), .ZN(n6726) );
  NOR2_X1 U7435 ( .A1(n6560), .A2(n6726), .ZN(U3151) );
  AND2_X1 U7436 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6496), .ZN(U3152) );
  AND2_X1 U7437 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6496), .ZN(U3153) );
  AND2_X1 U7438 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6496), .ZN(U3154) );
  INV_X1 U7439 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n6672) );
  NOR2_X1 U7440 ( .A1(n6560), .A2(n6672), .ZN(U3155) );
  AND2_X1 U7441 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6496), .ZN(U3156) );
  AND2_X1 U7442 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6496), .ZN(U3157) );
  INV_X1 U7443 ( .A(DATAWIDTH_REG_24__SCAN_IN), .ZN(n6597) );
  NOR2_X1 U7444 ( .A1(n6560), .A2(n6597), .ZN(U3158) );
  AND2_X1 U7445 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6496), .ZN(U3159) );
  AND2_X1 U7446 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6496), .ZN(U3160) );
  AND2_X1 U7447 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6496), .ZN(U3161) );
  AND2_X1 U7448 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6496), .ZN(U3162) );
  AND2_X1 U7449 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6496), .ZN(U3163) );
  AND2_X1 U7450 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6496), .ZN(U3164) );
  AND2_X1 U7451 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6496), .ZN(U3165) );
  AND2_X1 U7452 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6496), .ZN(U3166) );
  AND2_X1 U7453 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6496), .ZN(U3167) );
  AND2_X1 U7454 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6496), .ZN(U3168) );
  AND2_X1 U7455 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6496), .ZN(U3169) );
  AND2_X1 U7456 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6496), .ZN(U3170) );
  INV_X1 U7457 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6761) );
  NOR2_X1 U7458 ( .A1(n6560), .A2(n6761), .ZN(U3171) );
  INV_X1 U7459 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6645) );
  NOR2_X1 U7460 ( .A1(n6560), .A2(n6645), .ZN(U3172) );
  AND2_X1 U7461 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6496), .ZN(U3173) );
  AND2_X1 U7462 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6496), .ZN(U3174) );
  AND2_X1 U7463 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6496), .ZN(U3175) );
  AND2_X1 U7464 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6496), .ZN(U3176) );
  AND2_X1 U7465 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6496), .ZN(U3177) );
  AND2_X1 U7466 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6496), .ZN(U3178) );
  AND2_X1 U7467 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6496), .ZN(U3179) );
  AND2_X1 U7468 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6496), .ZN(U3180) );
  NOR2_X1 U7469 ( .A1(n6504), .A2(n6513), .ZN(n6498) );
  AOI22_X1 U7470 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6512) );
  AND2_X1 U7471 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6501) );
  INV_X1 U7472 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6499) );
  INV_X1 U7473 ( .A(NA_N), .ZN(n6625) );
  AOI221_X1 U7474 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6625), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6509) );
  AOI221_X1 U7475 ( .B1(n6501), .B2(n6593), .C1(n6499), .C2(n6593), .A(n6509), 
        .ZN(n6497) );
  OAI21_X1 U7476 ( .B1(n6498), .B2(n6512), .A(n6497), .ZN(U3181) );
  NOR2_X1 U7477 ( .A1(n6507), .A2(n6499), .ZN(n6505) );
  NAND2_X1 U7478 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6500) );
  OAI21_X1 U7479 ( .B1(n6505), .B2(n6501), .A(n6500), .ZN(n6502) );
  OAI211_X1 U7480 ( .C1(n6504), .C2(n6506), .A(n6503), .B(n6502), .ZN(U3182)
         );
  AOI22_X1 U7481 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .B1(
        n6505), .B2(n6625), .ZN(n6511) );
  AOI221_X1 U7482 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6506), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6508) );
  AOI221_X1 U7483 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6508), .C2(HOLD), .A(n6507), .ZN(n6510) );
  OAI22_X1 U7484 ( .A1(n6512), .A2(n6511), .B1(n6510), .B2(n6509), .ZN(U3183)
         );
  NOR2_X1 U7485 ( .A1(n6513), .A2(n6593), .ZN(n6550) );
  INV_X1 U7486 ( .A(n6550), .ZN(n6555) );
  INV_X1 U7487 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6637) );
  NOR2_X2 U7488 ( .A1(n6593), .A2(STATE_REG_2__SCAN_IN), .ZN(n6553) );
  OAI222_X1 U7489 ( .A1(n6555), .A2(n6570), .B1(n6637), .B2(n6547), .C1(n6698), 
        .C2(n6552), .ZN(U3184) );
  AOI22_X1 U7490 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6553), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6580), .ZN(n6514) );
  OAI21_X1 U7491 ( .B1(n6698), .B2(n6555), .A(n6514), .ZN(U3185) );
  AOI22_X1 U7492 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6553), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6593), .ZN(n6515) );
  OAI21_X1 U7493 ( .B1(n4845), .B2(n6555), .A(n6515), .ZN(U3186) );
  AOI22_X1 U7494 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6593), .ZN(n6516) );
  OAI21_X1 U7495 ( .B1(n6657), .B2(n6552), .A(n6516), .ZN(U3187) );
  INV_X1 U7496 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n6809) );
  OAI222_X1 U7497 ( .A1(n6552), .A2(n6518), .B1(n6809), .B2(n6547), .C1(n6657), 
        .C2(n6555), .ZN(U3188) );
  AOI22_X1 U7498 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6553), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6593), .ZN(n6517) );
  OAI21_X1 U7499 ( .B1(n6518), .B2(n6555), .A(n6517), .ZN(U3189) );
  AOI22_X1 U7500 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6593), .ZN(n6519) );
  OAI21_X1 U7501 ( .B1(n4972), .B2(n6552), .A(n6519), .ZN(U3190) );
  AOI22_X1 U7502 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6553), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6580), .ZN(n6520) );
  OAI21_X1 U7503 ( .B1(n4972), .B2(n6555), .A(n6520), .ZN(U3191) );
  INV_X1 U7504 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6610) );
  OAI222_X1 U7505 ( .A1(n6555), .A2(n6522), .B1(n6610), .B2(n6547), .C1(n6521), 
        .C2(n6552), .ZN(U3192) );
  AOI22_X1 U7506 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6580), .ZN(n6523) );
  OAI21_X1 U7507 ( .B1(n6525), .B2(n6552), .A(n6523), .ZN(U3193) );
  AOI22_X1 U7508 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6553), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6580), .ZN(n6524) );
  OAI21_X1 U7509 ( .B1(n6525), .B2(n6555), .A(n6524), .ZN(U3194) );
  AOI22_X1 U7510 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6553), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6580), .ZN(n6526) );
  OAI21_X1 U7511 ( .B1(n6527), .B2(n6555), .A(n6526), .ZN(U3195) );
  AOI22_X1 U7512 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6553), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6580), .ZN(n6528) );
  OAI21_X1 U7513 ( .B1(n6686), .B2(n6555), .A(n6528), .ZN(U3196) );
  INV_X1 U7514 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6531) );
  AOI22_X1 U7515 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6580), .ZN(n6529) );
  OAI21_X1 U7516 ( .B1(n6531), .B2(n6552), .A(n6529), .ZN(U3197) );
  AOI22_X1 U7517 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6553), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6580), .ZN(n6530) );
  OAI21_X1 U7518 ( .B1(n6531), .B2(n6555), .A(n6530), .ZN(U3198) );
  AOI22_X1 U7519 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6553), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6580), .ZN(n6532) );
  OAI21_X1 U7520 ( .B1(n5518), .B2(n6555), .A(n6532), .ZN(U3199) );
  AOI22_X1 U7521 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6580), .ZN(n6533) );
  OAI21_X1 U7522 ( .B1(n6535), .B2(n6552), .A(n6533), .ZN(U3200) );
  AOI22_X1 U7523 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6553), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6580), .ZN(n6534) );
  OAI21_X1 U7524 ( .B1(n6535), .B2(n6555), .A(n6534), .ZN(U3201) );
  AOI22_X1 U7525 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6553), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6580), .ZN(n6536) );
  OAI21_X1 U7526 ( .B1(n5495), .B2(n6555), .A(n6536), .ZN(U3202) );
  AOI22_X1 U7527 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6580), .ZN(n6537) );
  OAI21_X1 U7528 ( .B1(n6539), .B2(n6552), .A(n6537), .ZN(U3203) );
  AOI22_X1 U7529 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6553), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6580), .ZN(n6538) );
  OAI21_X1 U7530 ( .B1(n6539), .B2(n6555), .A(n6538), .ZN(U3204) );
  AOI22_X1 U7531 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6580), .ZN(n6540) );
  OAI21_X1 U7532 ( .B1(n6541), .B2(n6552), .A(n6540), .ZN(U3205) );
  INV_X1 U7533 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n6802) );
  OAI222_X1 U7534 ( .A1(n6555), .A2(n6541), .B1(n6802), .B2(n6547), .C1(n6542), 
        .C2(n6552), .ZN(U3206) );
  INV_X1 U7535 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6791) );
  OAI222_X1 U7536 ( .A1(n6552), .A2(n6544), .B1(n6791), .B2(n6547), .C1(n6542), 
        .C2(n6555), .ZN(U3207) );
  AOI22_X1 U7537 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6553), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6593), .ZN(n6543) );
  OAI21_X1 U7538 ( .B1(n6544), .B2(n6555), .A(n6543), .ZN(U3208) );
  AOI22_X1 U7539 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6553), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6580), .ZN(n6545) );
  OAI21_X1 U7540 ( .B1(n6546), .B2(n6555), .A(n6545), .ZN(U3209) );
  INV_X1 U7541 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6815) );
  OAI222_X1 U7542 ( .A1(n6555), .A2(n6548), .B1(n6815), .B2(n6547), .C1(n5133), 
        .C2(n6552), .ZN(U3210) );
  AOI22_X1 U7543 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6553), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6580), .ZN(n6549) );
  OAI21_X1 U7544 ( .B1(n5133), .B2(n6555), .A(n6549), .ZN(U3211) );
  AOI22_X1 U7545 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6550), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6580), .ZN(n6551) );
  OAI21_X1 U7546 ( .B1(n6556), .B2(n6552), .A(n6551), .ZN(U3212) );
  AOI22_X1 U7547 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6553), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6580), .ZN(n6554) );
  OAI21_X1 U7548 ( .B1(n6556), .B2(n6555), .A(n6554), .ZN(U3213) );
  MUX2_X1 U7549 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6593), .Z(U3445) );
  MUX2_X1 U7550 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6593), .Z(U3446) );
  MUX2_X1 U7551 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6593), .Z(U3447) );
  MUX2_X1 U7552 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6593), .Z(U3448) );
  OAI21_X1 U7553 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6560), .A(n6558), .ZN(
        n6557) );
  INV_X1 U7554 ( .A(n6557), .ZN(U3451) );
  OAI21_X1 U7555 ( .B1(n6560), .B2(n6559), .A(n6558), .ZN(U3452) );
  OAI211_X1 U7556 ( .C1(n6688), .C2(n6563), .A(n6562), .B(n6561), .ZN(U3453)
         );
  OAI22_X1 U7557 ( .A1(n6567), .A2(n6566), .B1(n6565), .B2(n6564), .ZN(n6569)
         );
  MUX2_X1 U7558 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6569), .S(n6568), 
        .Z(U3456) );
  AOI21_X1 U7559 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6571) );
  AOI22_X1 U7560 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6571), .B2(n6570), .ZN(n6573) );
  INV_X1 U7561 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6572) );
  AOI22_X1 U7562 ( .A1(n6574), .A2(n6573), .B1(n6572), .B2(n6577), .ZN(U3468)
         );
  INV_X1 U7563 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6578) );
  NOR2_X1 U7564 ( .A1(n6577), .A2(REIP_REG_1__SCAN_IN), .ZN(n6575) );
  AOI22_X1 U7565 ( .A1(n6578), .A2(n6577), .B1(n6576), .B2(n6575), .ZN(U3469)
         );
  NAND2_X1 U7566 ( .A1(n6580), .A2(W_R_N_REG_SCAN_IN), .ZN(n6579) );
  OAI21_X1 U7567 ( .B1(n6580), .B2(READREQUEST_REG_SCAN_IN), .A(n6579), .ZN(
        U3470) );
  INV_X1 U7568 ( .A(n6581), .ZN(n6582) );
  OAI21_X1 U7569 ( .B1(n6587), .B2(n6586), .A(n6585), .ZN(n6592) );
  OAI211_X1 U7570 ( .C1(READY_N), .C2(n6590), .A(n6589), .B(n6588), .ZN(n6591)
         );
  MUX2_X1 U7571 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(n6592), .S(n6591), .Z(
        U3472) );
  MUX2_X1 U7572 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6593), .Z(U3473) );
  INV_X1 U7573 ( .A(DATAI_14_), .ZN(n6595) );
  AOI22_X1 U7574 ( .A1(n6595), .A2(keyinput6), .B1(n3571), .B2(keyinput24), 
        .ZN(n6594) );
  OAI221_X1 U7575 ( .B1(n6595), .B2(keyinput6), .C1(n3571), .C2(keyinput24), 
        .A(n6594), .ZN(n6607) );
  AOI22_X1 U7576 ( .A1(n6598), .A2(keyinput29), .B1(n6597), .B2(keyinput104), 
        .ZN(n6596) );
  OAI221_X1 U7577 ( .B1(n6598), .B2(keyinput29), .C1(n6597), .C2(keyinput104), 
        .A(n6596), .ZN(n6606) );
  AOI22_X1 U7578 ( .A1(n6601), .A2(keyinput98), .B1(n6600), .B2(keyinput31), 
        .ZN(n6599) );
  OAI221_X1 U7579 ( .B1(n6601), .B2(keyinput98), .C1(n6600), .C2(keyinput31), 
        .A(n6599), .ZN(n6605) );
  AOI22_X1 U7580 ( .A1(n6843), .A2(keyinput5), .B1(keyinput114), .B2(n6603), 
        .ZN(n6602) );
  OAI221_X1 U7581 ( .B1(n6843), .B2(keyinput5), .C1(n6603), .C2(keyinput114), 
        .A(n6602), .ZN(n6604) );
  NOR4_X1 U7582 ( .A1(n6607), .A2(n6606), .A3(n6605), .A4(n6604), .ZN(n6653)
         );
  AOI22_X1 U7583 ( .A1(n6610), .A2(keyinput119), .B1(n6609), .B2(keyinput61), 
        .ZN(n6608) );
  OAI221_X1 U7584 ( .B1(n6610), .B2(keyinput119), .C1(n6609), .C2(keyinput61), 
        .A(n6608), .ZN(n6622) );
  INV_X1 U7585 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n6612) );
  AOI22_X1 U7586 ( .A1(n6613), .A2(keyinput78), .B1(keyinput45), .B2(n6612), 
        .ZN(n6611) );
  OAI221_X1 U7587 ( .B1(n6613), .B2(keyinput78), .C1(n6612), .C2(keyinput45), 
        .A(n6611), .ZN(n6621) );
  INV_X1 U7588 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6873) );
  AOI22_X1 U7589 ( .A1(n6615), .A2(keyinput20), .B1(n6873), .B2(keyinput25), 
        .ZN(n6614) );
  OAI221_X1 U7590 ( .B1(n6615), .B2(keyinput20), .C1(n6873), .C2(keyinput25), 
        .A(n6614), .ZN(n6620) );
  AOI22_X1 U7591 ( .A1(n6618), .A2(keyinput105), .B1(keyinput103), .B2(n6617), 
        .ZN(n6616) );
  OAI221_X1 U7592 ( .B1(n6618), .B2(keyinput105), .C1(n6617), .C2(keyinput103), 
        .A(n6616), .ZN(n6619) );
  NOR4_X1 U7593 ( .A1(n6622), .A2(n6621), .A3(n6620), .A4(n6619), .ZN(n6652)
         );
  AOI22_X1 U7594 ( .A1(n6625), .A2(keyinput67), .B1(n6624), .B2(keyinput110), 
        .ZN(n6623) );
  OAI221_X1 U7595 ( .B1(n6625), .B2(keyinput67), .C1(n6624), .C2(keyinput110), 
        .A(n6623), .ZN(n6635) );
  AOI22_X1 U7596 ( .A1(n6838), .A2(keyinput40), .B1(keyinput101), .B2(n6627), 
        .ZN(n6626) );
  OAI221_X1 U7597 ( .B1(n6838), .B2(keyinput40), .C1(n6627), .C2(keyinput101), 
        .A(n6626), .ZN(n6634) );
  INV_X1 U7598 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n6835) );
  AOI22_X1 U7599 ( .A1(n6835), .A2(keyinput112), .B1(n6629), .B2(keyinput38), 
        .ZN(n6628) );
  OAI221_X1 U7600 ( .B1(n6835), .B2(keyinput112), .C1(n6629), .C2(keyinput38), 
        .A(n6628), .ZN(n6633) );
  INV_X1 U7601 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6631) );
  INV_X1 U7602 ( .A(DATAI_28_), .ZN(n6874) );
  AOI22_X1 U7603 ( .A1(n6631), .A2(keyinput117), .B1(keyinput11), .B2(n6874), 
        .ZN(n6630) );
  OAI221_X1 U7604 ( .B1(n6631), .B2(keyinput117), .C1(n6874), .C2(keyinput11), 
        .A(n6630), .ZN(n6632) );
  NOR4_X1 U7605 ( .A1(n6635), .A2(n6634), .A3(n6633), .A4(n6632), .ZN(n6651)
         );
  AOI22_X1 U7606 ( .A1(n6638), .A2(keyinput88), .B1(keyinput68), .B2(n6637), 
        .ZN(n6636) );
  OAI221_X1 U7607 ( .B1(n6638), .B2(keyinput88), .C1(n6637), .C2(keyinput68), 
        .A(n6636), .ZN(n6649) );
  INV_X1 U7608 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n6640) );
  AOI22_X1 U7609 ( .A1(n6641), .A2(keyinput34), .B1(n6640), .B2(keyinput73), 
        .ZN(n6639) );
  OAI221_X1 U7610 ( .B1(n6641), .B2(keyinput34), .C1(n6640), .C2(keyinput73), 
        .A(n6639), .ZN(n6648) );
  INV_X1 U7611 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n6643) );
  AOI22_X1 U7612 ( .A1(n6643), .A2(keyinput66), .B1(keyinput16), .B2(n3582), 
        .ZN(n6642) );
  OAI221_X1 U7613 ( .B1(n6643), .B2(keyinput66), .C1(n3582), .C2(keyinput16), 
        .A(n6642), .ZN(n6647) );
  AOI22_X1 U7614 ( .A1(n6645), .A2(keyinput17), .B1(n4205), .B2(keyinput116), 
        .ZN(n6644) );
  OAI221_X1 U7615 ( .B1(n6645), .B2(keyinput17), .C1(n4205), .C2(keyinput116), 
        .A(n6644), .ZN(n6646) );
  NOR4_X1 U7616 ( .A1(n6649), .A2(n6648), .A3(n6647), .A4(n6646), .ZN(n6650)
         );
  NAND4_X1 U7617 ( .A1(n6653), .A2(n6652), .A3(n6651), .A4(n6650), .ZN(n6829)
         );
  AOI22_X1 U7618 ( .A1(n3574), .A2(keyinput63), .B1(keyinput46), .B2(n6655), 
        .ZN(n6654) );
  OAI221_X1 U7619 ( .B1(n3574), .B2(keyinput63), .C1(n6655), .C2(keyinput46), 
        .A(n6654), .ZN(n6667) );
  AOI22_X1 U7620 ( .A1(n6876), .A2(keyinput1), .B1(keyinput115), .B2(n6657), 
        .ZN(n6656) );
  OAI221_X1 U7621 ( .B1(n6876), .B2(keyinput1), .C1(n6657), .C2(keyinput115), 
        .A(n6656), .ZN(n6666) );
  AOI22_X1 U7622 ( .A1(n6660), .A2(keyinput47), .B1(n6659), .B2(keyinput111), 
        .ZN(n6658) );
  OAI221_X1 U7623 ( .B1(n6660), .B2(keyinput47), .C1(n6659), .C2(keyinput111), 
        .A(n6658), .ZN(n6665) );
  AOI22_X1 U7624 ( .A1(n6663), .A2(keyinput19), .B1(n6662), .B2(keyinput94), 
        .ZN(n6661) );
  OAI221_X1 U7625 ( .B1(n6663), .B2(keyinput19), .C1(n6662), .C2(keyinput94), 
        .A(n6661), .ZN(n6664) );
  NOR4_X1 U7626 ( .A1(n6667), .A2(n6666), .A3(n6665), .A4(n6664), .ZN(n6711)
         );
  AOI22_X1 U7627 ( .A1(n6834), .A2(keyinput49), .B1(keyinput41), .B2(n6669), 
        .ZN(n6668) );
  OAI221_X1 U7628 ( .B1(n6834), .B2(keyinput49), .C1(n6669), .C2(keyinput41), 
        .A(n6668), .ZN(n6681) );
  AOI22_X1 U7629 ( .A1(n6672), .A2(keyinput10), .B1(keyinput50), .B2(n6671), 
        .ZN(n6670) );
  OAI221_X1 U7630 ( .B1(n6672), .B2(keyinput10), .C1(n6671), .C2(keyinput50), 
        .A(n6670), .ZN(n6680) );
  AOI22_X1 U7631 ( .A1(n4463), .A2(keyinput102), .B1(n6674), .B2(keyinput118), 
        .ZN(n6673) );
  OAI221_X1 U7632 ( .B1(n4463), .B2(keyinput102), .C1(n6674), .C2(keyinput118), 
        .A(n6673), .ZN(n6679) );
  INV_X1 U7633 ( .A(DATAI_17_), .ZN(n6676) );
  AOI22_X1 U7634 ( .A1(n6677), .A2(keyinput57), .B1(n6676), .B2(keyinput27), 
        .ZN(n6675) );
  OAI221_X1 U7635 ( .B1(n6677), .B2(keyinput57), .C1(n6676), .C2(keyinput27), 
        .A(n6675), .ZN(n6678) );
  NOR4_X1 U7636 ( .A1(n6681), .A2(n6680), .A3(n6679), .A4(n6678), .ZN(n6710)
         );
  INV_X1 U7637 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n6683) );
  AOI22_X1 U7638 ( .A1(n6684), .A2(keyinput95), .B1(n6683), .B2(keyinput23), 
        .ZN(n6682) );
  OAI221_X1 U7639 ( .B1(n6684), .B2(keyinput95), .C1(n6683), .C2(keyinput23), 
        .A(n6682), .ZN(n6694) );
  AOI22_X1 U7640 ( .A1(n6686), .A2(keyinput79), .B1(n6869), .B2(keyinput91), 
        .ZN(n6685) );
  OAI221_X1 U7641 ( .B1(n6686), .B2(keyinput79), .C1(n6869), .C2(keyinput91), 
        .A(n6685), .ZN(n6693) );
  AOI22_X1 U7642 ( .A1(n6870), .A2(keyinput7), .B1(n6688), .B2(keyinput48), 
        .ZN(n6687) );
  OAI221_X1 U7643 ( .B1(n6870), .B2(keyinput7), .C1(n6688), .C2(keyinput48), 
        .A(n6687), .ZN(n6692) );
  INV_X1 U7644 ( .A(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n6857) );
  AOI22_X1 U7645 ( .A1(n6857), .A2(keyinput65), .B1(n6690), .B2(keyinput89), 
        .ZN(n6689) );
  OAI221_X1 U7646 ( .B1(n6857), .B2(keyinput65), .C1(n6690), .C2(keyinput89), 
        .A(n6689), .ZN(n6691) );
  NOR4_X1 U7647 ( .A1(n6694), .A2(n6693), .A3(n6692), .A4(n6691), .ZN(n6709)
         );
  AOI22_X1 U7648 ( .A1(n6696), .A2(keyinput99), .B1(keyinput125), .B2(n4461), 
        .ZN(n6695) );
  OAI221_X1 U7649 ( .B1(n6696), .B2(keyinput99), .C1(n4461), .C2(keyinput125), 
        .A(n6695), .ZN(n6707) );
  AOI22_X1 U7650 ( .A1(n4791), .A2(keyinput84), .B1(keyinput72), .B2(n6698), 
        .ZN(n6697) );
  OAI221_X1 U7651 ( .B1(n4791), .B2(keyinput84), .C1(n6698), .C2(keyinput72), 
        .A(n6697), .ZN(n6706) );
  AOI22_X1 U7652 ( .A1(n6700), .A2(keyinput64), .B1(n6858), .B2(keyinput4), 
        .ZN(n6699) );
  OAI221_X1 U7653 ( .B1(n6700), .B2(keyinput64), .C1(n6858), .C2(keyinput4), 
        .A(n6699), .ZN(n6705) );
  INV_X1 U7654 ( .A(DATAI_27_), .ZN(n6703) );
  AOI22_X1 U7655 ( .A1(n6703), .A2(keyinput18), .B1(n6702), .B2(keyinput96), 
        .ZN(n6701) );
  OAI221_X1 U7656 ( .B1(n6703), .B2(keyinput18), .C1(n6702), .C2(keyinput96), 
        .A(n6701), .ZN(n6704) );
  NOR4_X1 U7657 ( .A1(n6707), .A2(n6706), .A3(n6705), .A4(n6704), .ZN(n6708)
         );
  NAND4_X1 U7658 ( .A1(n6711), .A2(n6710), .A3(n6709), .A4(n6708), .ZN(n6828)
         );
  AOI22_X1 U7659 ( .A1(n6713), .A2(keyinput120), .B1(n4972), .B2(keyinput42), 
        .ZN(n6712) );
  OAI221_X1 U7660 ( .B1(n6713), .B2(keyinput120), .C1(n4972), .C2(keyinput42), 
        .A(n6712), .ZN(n6723) );
  INV_X1 U7661 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n6715) );
  AOI22_X1 U7662 ( .A1(n6715), .A2(keyinput14), .B1(n5500), .B2(keyinput87), 
        .ZN(n6714) );
  OAI221_X1 U7663 ( .B1(n6715), .B2(keyinput14), .C1(n5500), .C2(keyinput87), 
        .A(n6714), .ZN(n6722) );
  INV_X1 U7664 ( .A(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n6839) );
  AOI22_X1 U7665 ( .A1(n6839), .A2(keyinput75), .B1(keyinput12), .B2(n6717), 
        .ZN(n6716) );
  OAI221_X1 U7666 ( .B1(n6839), .B2(keyinput75), .C1(n6717), .C2(keyinput12), 
        .A(n6716), .ZN(n6721) );
  INV_X1 U7667 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n6719) );
  AOI22_X1 U7668 ( .A1(n6872), .A2(keyinput71), .B1(keyinput15), .B2(n6719), 
        .ZN(n6718) );
  OAI221_X1 U7669 ( .B1(n6872), .B2(keyinput71), .C1(n6719), .C2(keyinput15), 
        .A(n6718), .ZN(n6720) );
  NOR4_X1 U7670 ( .A1(n6723), .A2(n6722), .A3(n6721), .A4(n6720), .ZN(n6769)
         );
  AOI22_X1 U7671 ( .A1(n6726), .A2(keyinput85), .B1(keyinput58), .B2(n6725), 
        .ZN(n6724) );
  OAI221_X1 U7672 ( .B1(n6726), .B2(keyinput85), .C1(n6725), .C2(keyinput58), 
        .A(n6724), .ZN(n6737) );
  AOI22_X1 U7673 ( .A1(n4845), .A2(keyinput3), .B1(n6728), .B2(keyinput26), 
        .ZN(n6727) );
  OAI221_X1 U7674 ( .B1(n4845), .B2(keyinput3), .C1(n6728), .C2(keyinput26), 
        .A(n6727), .ZN(n6736) );
  INV_X1 U7675 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n6730) );
  AOI22_X1 U7676 ( .A1(n6731), .A2(keyinput77), .B1(n6730), .B2(keyinput126), 
        .ZN(n6729) );
  OAI221_X1 U7677 ( .B1(n6731), .B2(keyinput77), .C1(n6730), .C2(keyinput126), 
        .A(n6729), .ZN(n6735) );
  XNOR2_X1 U7678 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .B(keyinput13), .ZN(
        n6733) );
  XNOR2_X1 U7679 ( .A(INSTQUEUE_REG_9__4__SCAN_IN), .B(keyinput127), .ZN(n6732) );
  NAND2_X1 U7680 ( .A1(n6733), .A2(n6732), .ZN(n6734) );
  NOR4_X1 U7681 ( .A1(n6737), .A2(n6736), .A3(n6735), .A4(n6734), .ZN(n6768)
         );
  AOI22_X1 U7682 ( .A1(n6739), .A2(keyinput32), .B1(keyinput35), .B2(n3153), 
        .ZN(n6738) );
  OAI221_X1 U7683 ( .B1(n6739), .B2(keyinput32), .C1(n3153), .C2(keyinput35), 
        .A(n6738), .ZN(n6751) );
  INV_X1 U7684 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n6741) );
  AOI22_X1 U7685 ( .A1(n6742), .A2(keyinput123), .B1(n6741), .B2(keyinput21), 
        .ZN(n6740) );
  OAI221_X1 U7686 ( .B1(n6742), .B2(keyinput123), .C1(n6741), .C2(keyinput21), 
        .A(n6740), .ZN(n6750) );
  AOI22_X1 U7687 ( .A1(n6744), .A2(keyinput44), .B1(n5062), .B2(keyinput93), 
        .ZN(n6743) );
  OAI221_X1 U7688 ( .B1(n6744), .B2(keyinput44), .C1(n5062), .C2(keyinput93), 
        .A(n6743), .ZN(n6749) );
  XOR2_X1 U7689 ( .A(n6745), .B(keyinput86), .Z(n6747) );
  XNOR2_X1 U7690 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .B(keyinput43), .ZN(n6746)
         );
  NAND2_X1 U7691 ( .A1(n6747), .A2(n6746), .ZN(n6748) );
  NOR4_X1 U7692 ( .A1(n6751), .A2(n6750), .A3(n6749), .A4(n6748), .ZN(n6767)
         );
  AOI22_X1 U7693 ( .A1(n6754), .A2(keyinput109), .B1(keyinput54), .B2(n6753), 
        .ZN(n6752) );
  OAI221_X1 U7694 ( .B1(n6754), .B2(keyinput109), .C1(n6753), .C2(keyinput54), 
        .A(n6752), .ZN(n6765) );
  AOI22_X1 U7695 ( .A1(n6757), .A2(keyinput0), .B1(keyinput28), .B2(n6756), 
        .ZN(n6755) );
  INV_X1 U7696 ( .A(DATAI_21_), .ZN(n6868) );
  AOI22_X1 U7697 ( .A1(n6868), .A2(keyinput9), .B1(n4270), .B2(keyinput121), 
        .ZN(n6758) );
  OAI221_X1 U7698 ( .B1(n6868), .B2(keyinput9), .C1(n4270), .C2(keyinput121), 
        .A(n6758), .ZN(n6763) );
  AOI22_X1 U7699 ( .A1(n6761), .A2(keyinput30), .B1(n6760), .B2(keyinput82), 
        .ZN(n6759) );
  OAI221_X1 U7700 ( .B1(n6761), .B2(keyinput30), .C1(n6760), .C2(keyinput82), 
        .A(n6759), .ZN(n6762) );
  NOR4_X1 U7701 ( .A1(n6765), .A2(n6764), .A3(n6763), .A4(n6762), .ZN(n6766)
         );
  NAND4_X1 U7702 ( .A1(n6769), .A2(n6768), .A3(n6767), .A4(n6766), .ZN(n6827)
         );
  INV_X1 U7703 ( .A(LWORD_REG_9__SCAN_IN), .ZN(n6771) );
  AOI22_X1 U7704 ( .A1(n6772), .A2(keyinput108), .B1(keyinput70), .B2(n6771), 
        .ZN(n6770) );
  OAI221_X1 U7705 ( .B1(n6772), .B2(keyinput108), .C1(n6771), .C2(keyinput70), 
        .A(n6770), .ZN(n6782) );
  INV_X1 U7706 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6774) );
  AOI22_X1 U7707 ( .A1(n6774), .A2(keyinput124), .B1(n3381), .B2(keyinput106), 
        .ZN(n6773) );
  OAI221_X1 U7708 ( .B1(n6774), .B2(keyinput124), .C1(n3381), .C2(keyinput106), 
        .A(n6773), .ZN(n6781) );
  AOI22_X1 U7709 ( .A1(n3729), .A2(keyinput53), .B1(n6877), .B2(keyinput60), 
        .ZN(n6775) );
  OAI221_X1 U7710 ( .B1(n3729), .B2(keyinput53), .C1(n6877), .C2(keyinput60), 
        .A(n6775), .ZN(n6780) );
  INV_X1 U7711 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n6777) );
  AOI22_X1 U7712 ( .A1(n6778), .A2(keyinput62), .B1(n6777), .B2(keyinput39), 
        .ZN(n6776) );
  OAI221_X1 U7713 ( .B1(n6778), .B2(keyinput62), .C1(n6777), .C2(keyinput39), 
        .A(n6776), .ZN(n6779) );
  NOR4_X1 U7714 ( .A1(n6782), .A2(n6781), .A3(n6780), .A4(n6779), .ZN(n6825)
         );
  INV_X1 U7715 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6785) );
  AOI22_X1 U7716 ( .A1(n6785), .A2(keyinput92), .B1(keyinput56), .B2(n6784), 
        .ZN(n6783) );
  OAI221_X1 U7717 ( .B1(n6785), .B2(keyinput92), .C1(n6784), .C2(keyinput56), 
        .A(n6783), .ZN(n6795) );
  INV_X1 U7718 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n6787) );
  AOI22_X1 U7719 ( .A1(n6867), .A2(keyinput90), .B1(n6787), .B2(keyinput83), 
        .ZN(n6786) );
  OAI221_X1 U7720 ( .B1(n6867), .B2(keyinput90), .C1(n6787), .C2(keyinput83), 
        .A(n6786), .ZN(n6794) );
  AOI22_X1 U7721 ( .A1(n6789), .A2(keyinput74), .B1(n6875), .B2(keyinput69), 
        .ZN(n6788) );
  OAI221_X1 U7722 ( .B1(n6789), .B2(keyinput74), .C1(n6875), .C2(keyinput69), 
        .A(n6788), .ZN(n6793) );
  INV_X1 U7723 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n6841) );
  AOI22_X1 U7724 ( .A1(n6791), .A2(keyinput33), .B1(n6841), .B2(keyinput51), 
        .ZN(n6790) );
  OAI221_X1 U7725 ( .B1(n6791), .B2(keyinput33), .C1(n6841), .C2(keyinput51), 
        .A(n6790), .ZN(n6792) );
  NOR4_X1 U7726 ( .A1(n6795), .A2(n6794), .A3(n6793), .A4(n6792), .ZN(n6824)
         );
  AOI22_X1 U7727 ( .A1(n4782), .A2(keyinput80), .B1(keyinput59), .B2(n3848), 
        .ZN(n6796) );
  OAI221_X1 U7728 ( .B1(n4782), .B2(keyinput80), .C1(n3848), .C2(keyinput59), 
        .A(n6796), .ZN(n6806) );
  INV_X1 U7729 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n6840) );
  AOI22_X1 U7730 ( .A1(n6871), .A2(keyinput107), .B1(n6840), .B2(keyinput122), 
        .ZN(n6797) );
  OAI221_X1 U7731 ( .B1(n6871), .B2(keyinput107), .C1(n6840), .C2(keyinput122), 
        .A(n6797), .ZN(n6805) );
  INV_X1 U7732 ( .A(EAX_REG_31__SCAN_IN), .ZN(n6799) );
  AOI22_X1 U7733 ( .A1(n6800), .A2(keyinput97), .B1(keyinput81), .B2(n6799), 
        .ZN(n6798) );
  OAI221_X1 U7734 ( .B1(n6800), .B2(keyinput97), .C1(n6799), .C2(keyinput81), 
        .A(n6798), .ZN(n6804) );
  INV_X1 U7735 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n6842) );
  AOI22_X1 U7736 ( .A1(n6842), .A2(keyinput76), .B1(keyinput2), .B2(n6802), 
        .ZN(n6801) );
  OAI221_X1 U7737 ( .B1(n6842), .B2(keyinput76), .C1(n6802), .C2(keyinput2), 
        .A(n6801), .ZN(n6803) );
  NOR4_X1 U7738 ( .A1(n6806), .A2(n6805), .A3(n6804), .A4(n6803), .ZN(n6823)
         );
  INV_X1 U7739 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n6808) );
  AOI22_X1 U7740 ( .A1(n6809), .A2(keyinput37), .B1(n6808), .B2(keyinput36), 
        .ZN(n6807) );
  OAI221_X1 U7741 ( .B1(n6809), .B2(keyinput37), .C1(n6808), .C2(keyinput36), 
        .A(n6807), .ZN(n6821) );
  INV_X1 U7742 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n6812) );
  AOI22_X1 U7743 ( .A1(n6812), .A2(keyinput22), .B1(keyinput113), .B2(n6811), 
        .ZN(n6810) );
  OAI221_X1 U7744 ( .B1(n6812), .B2(keyinput22), .C1(n6811), .C2(keyinput113), 
        .A(n6810), .ZN(n6820) );
  INV_X1 U7745 ( .A(DATAI_24_), .ZN(n6814) );
  AOI22_X1 U7746 ( .A1(n6815), .A2(keyinput100), .B1(n6814), .B2(keyinput52), 
        .ZN(n6813) );
  OAI221_X1 U7747 ( .B1(n6815), .B2(keyinput100), .C1(n6814), .C2(keyinput52), 
        .A(n6813), .ZN(n6819) );
  XNOR2_X1 U7748 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .B(keyinput55), .ZN(n6817) );
  XNOR2_X1 U7749 ( .A(keyinput8), .B(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n6816)
         );
  NAND2_X1 U7750 ( .A1(n6817), .A2(n6816), .ZN(n6818) );
  NOR4_X1 U7751 ( .A1(n6821), .A2(n6820), .A3(n6819), .A4(n6818), .ZN(n6822)
         );
  NAND4_X1 U7752 ( .A1(n6825), .A2(n6824), .A3(n6823), .A4(n6822), .ZN(n6826)
         );
  NOR4_X1 U7753 ( .A1(n6829), .A2(n6828), .A3(n6827), .A4(n6826), .ZN(n6901)
         );
  AOI222_X1 U7754 ( .A1(n6833), .A2(n6832), .B1(DATAI_5_), .B2(n6831), .C1(
        EAX_REG_5__SCAN_IN), .C2(n6830), .ZN(n6899) );
  NAND4_X1 U7755 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(
        INSTQUEUE_REG_0__7__SCAN_IN), .A3(n6835), .A4(n6834), .ZN(n6836) );
  NOR4_X1 U7756 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(
        INSTQUEUE_REG_14__7__SCAN_IN), .A3(n6837), .A4(n6836), .ZN(n6852) );
  NOR4_X1 U7757 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(
        INSTQUEUE_REG_14__4__SCAN_IN), .A3(INSTQUEUE_REG_5__4__SCAN_IN), .A4(
        INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6851) );
  NOR4_X1 U7758 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(
        INSTQUEUE_REG_4__6__SCAN_IN), .A3(n6838), .A4(n4791), .ZN(n6850) );
  NAND4_X1 U7759 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(
        INSTQUEUE_REG_11__3__SCAN_IN), .A3(n6840), .A4(n6839), .ZN(n6848) );
  NAND4_X1 U7760 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(
        INSTQUEUE_REG_5__0__SCAN_IN), .A3(n6841), .A4(n3381), .ZN(n6847) );
  NAND4_X1 U7761 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(
        INSTQUEUE_REG_14__1__SCAN_IN), .A3(INSTQUEUE_REG_2__1__SCAN_IN), .A4(
        n6842), .ZN(n6846) );
  INV_X1 U7762 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n6844) );
  NAND4_X1 U7763 ( .A1(n6844), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .A3(
        INSTQUEUE_REG_15__0__SCAN_IN), .A4(n6843), .ZN(n6845) );
  NOR4_X1 U7764 ( .A1(n6848), .A2(n6847), .A3(n6846), .A4(n6845), .ZN(n6849)
         );
  NAND4_X1 U7765 ( .A1(n6852), .A2(n6851), .A3(n6850), .A4(n6849), .ZN(n6897)
         );
  NOR4_X1 U7766 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(LWORD_REG_7__SCAN_IN), .A3(LWORD_REG_4__SCAN_IN), .A4(LWORD_REG_2__SCAN_IN), .ZN(n6856) );
  NOR4_X1 U7767 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(EAX_REG_6__SCAN_IN), 
        .A3(EAX_REG_7__SCAN_IN), .A4(ADDRESS_REG_26__SCAN_IN), .ZN(n6855) );
  NOR4_X1 U7768 ( .A1(EAX_REG_17__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        DATAI_2_), .A4(DATAO_REG_11__SCAN_IN), .ZN(n6854) );
  NOR4_X1 U7769 ( .A1(EAX_REG_9__SCAN_IN), .A2(LWORD_REG_1__SCAN_IN), .A3(
        UWORD_REG_14__SCAN_IN), .A4(DATAO_REG_8__SCAN_IN), .ZN(n6853) );
  NAND4_X1 U7770 ( .A1(n6856), .A2(n6855), .A3(n6854), .A4(n6853), .ZN(n6896)
         );
  NOR4_X1 U7771 ( .A1(EAX_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), 
        .A3(DATAWIDTH_REG_27__SCAN_IN), .A4(ADDRESS_REG_22__SCAN_IN), .ZN(
        n6862) );
  NOR4_X1 U7772 ( .A1(DATAO_REG_28__SCAN_IN), .A2(DATAO_REG_0__SCAN_IN), .A3(
        DATAO_REG_2__SCAN_IN), .A4(FLUSH_REG_SCAN_IN), .ZN(n6861) );
  NOR4_X1 U7773 ( .A1(DATAO_REG_6__SCAN_IN), .A2(UWORD_REG_4__SCAN_IN), .A3(
        DATAO_REG_26__SCAN_IN), .A4(DATAO_REG_27__SCAN_IN), .ZN(n6860) );
  AND4_X1 U7774 ( .A1(n6858), .A2(n6728), .A3(INSTQUEUE_REG_12__2__SCAN_IN), 
        .A4(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n6859) );
  NAND4_X1 U7775 ( .A1(n6862), .A2(n6861), .A3(n6860), .A4(n6859), .ZN(n6895)
         );
  NAND4_X1 U7776 ( .A1(ADDRESS_REG_4__SCAN_IN), .A2(ADDRESS_REG_0__SCAN_IN), 
        .A3(DATAWIDTH_REG_31__SCAN_IN), .A4(DATAO_REG_18__SCAN_IN), .ZN(n6866)
         );
  NAND4_X1 U7777 ( .A1(DATAO_REG_30__SCAN_IN), .A2(DATAO_REG_7__SCAN_IN), .A3(
        ADDRESS_REG_23__SCAN_IN), .A4(DATAO_REG_31__SCAN_IN), .ZN(n6865) );
  NAND4_X1 U7778 ( .A1(EBX_REG_5__SCAN_IN), .A2(EBX_REG_10__SCAN_IN), .A3(
        LWORD_REG_6__SCAN_IN), .A4(LWORD_REG_9__SCAN_IN), .ZN(n6864) );
  NAND4_X1 U7779 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(NA_N), .A4(BYTEENABLE_REG_1__SCAN_IN), 
        .ZN(n6863) );
  NOR4_X1 U7780 ( .A1(n6866), .A2(n6865), .A3(n6864), .A4(n6863), .ZN(n6893)
         );
  NAND4_X1 U7781 ( .A1(n4270), .A2(n6869), .A3(n6868), .A4(n6867), .ZN(n6881)
         );
  NAND4_X1 U7782 ( .A1(DATAO_REG_1__SCAN_IN), .A2(ADDRESS_REG_8__SCAN_IN), 
        .A3(n6873), .A4(n4205), .ZN(n6879) );
  NAND4_X1 U7783 ( .A1(n6877), .A2(n6876), .A3(n6875), .A4(n6874), .ZN(n6878)
         );
  NOR4_X1 U7784 ( .A1(n6881), .A2(n6880), .A3(n6879), .A4(n6878), .ZN(n6892)
         );
  NAND4_X1 U7785 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .A3(EAX_REG_19__SCAN_IN), .A4(
        EAX_REG_22__SCAN_IN), .ZN(n6885) );
  NAND4_X1 U7786 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .A3(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6884) );
  NAND4_X1 U7787 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        EAX_REG_31__SCAN_IN), .A3(DATAI_14_), .A4(DATAI_27_), .ZN(n6883) );
  NAND4_X1 U7788 ( .A1(EAX_REG_23__SCAN_IN), .A2(EAX_REG_29__SCAN_IN), .A3(
        DATAI_24_), .A4(DATAI_4_), .ZN(n6882) );
  NOR4_X1 U7789 ( .A1(n6885), .A2(n6884), .A3(n6883), .A4(n6882), .ZN(n6891)
         );
  NAND4_X1 U7790 ( .A1(EAX_REG_8__SCAN_IN), .A2(EAX_REG_11__SCAN_IN), .A3(
        EAX_REG_16__SCAN_IN), .A4(UWORD_REG_3__SCAN_IN), .ZN(n6889) );
  NAND4_X1 U7791 ( .A1(LWORD_REG_0__SCAN_IN), .A2(LWORD_REG_3__SCAN_IN), .A3(
        DATAO_REG_13__SCAN_IN), .A4(UWORD_REG_12__SCAN_IN), .ZN(n6888) );
  NAND4_X1 U7792 ( .A1(EBX_REG_6__SCAN_IN), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), 
        .A3(REIP_REG_8__SCAN_IN), .A4(REIP_REG_13__SCAN_IN), .ZN(n6887) );
  NAND4_X1 U7793 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        REIP_REG_5__SCAN_IN), .A3(REIP_REG_2__SCAN_IN), .A4(DATAI_17_), .ZN(
        n6886) );
  NOR4_X1 U7794 ( .A1(n6889), .A2(n6888), .A3(n6887), .A4(n6886), .ZN(n6890)
         );
  NAND4_X1 U7795 ( .A1(n6893), .A2(n6892), .A3(n6891), .A4(n6890), .ZN(n6894)
         );
  NOR4_X1 U7796 ( .A1(n6897), .A2(n6896), .A3(n6895), .A4(n6894), .ZN(n6898)
         );
  XOR2_X1 U7797 ( .A(n6899), .B(n6898), .Z(n6900) );
  XNOR2_X1 U7798 ( .A(n6901), .B(n6900), .ZN(U2886) );
  INV_X1 U3574 ( .A(n3339), .ZN(n3407) );
  OR2_X1 U3661 ( .A1(n4081), .A2(n3341), .ZN(n4524) );
  CLKBUF_X1 U3557 ( .A(n3316), .Z(n3331) );
  CLKBUF_X2 U3623 ( .A(n3339), .Z(n4510) );
endmodule

