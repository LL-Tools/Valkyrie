

module b14_C_AntiSAT_k_128_6 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4709, n4710;

  CLKBUF_X2 U2297 ( .A(n3328), .Z(n2056) );
  INV_X2 U2298 ( .A(n3343), .ZN(n3334) );
  INV_X1 U2299 ( .A(n3340), .ZN(n3328) );
  NAND3_X1 U2300 ( .A1(n2157), .A2(n2335), .A3(n2336), .ZN(n2942) );
  NAND2_X1 U2301 ( .A1(n2319), .A2(n2318), .ZN(n3810) );
  NAND2_X1 U2303 ( .A1(n2295), .A2(n4344), .ZN(n2609) );
  INV_X1 U2304 ( .A(n3340), .ZN(n2057) );
  INV_X1 U2305 ( .A(n3299), .ZN(n3342) );
  NOR2_X1 U2306 ( .A1(n4404), .A2(n4405), .ZN(n4403) );
  AND2_X1 U2307 ( .A1(n2708), .A2(n2707), .ZN(n4496) );
  OAI21_X2 U2308 ( .B1(n2673), .B2(IR_REG_22__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2686) );
  NAND2_X2 U2309 ( .A1(n2295), .A2(n2288), .ZN(n2351) );
  CLKBUF_X1 U2310 ( .A(n3328), .Z(n2055) );
  NAND2_X2 U2311 ( .A1(n2990), .A2(n2989), .ZN(n3177) );
  NAND2_X2 U2312 ( .A1(n3997), .A2(n3998), .ZN(n3996) );
  AOI21_X2 U2313 ( .B1(n4012), .B2(n2535), .A(n2259), .ZN(n3997) );
  NAND2_X2 U2314 ( .A1(n2524), .A2(n3748), .ZN(n4012) );
  XNOR2_X1 U2315 ( .A(n2967), .B(n2968), .ZN(n2949) );
  AOI21_X1 U2316 ( .B1(n2941), .B2(n2940), .A(n2939), .ZN(n2950) );
  XNOR2_X2 U2317 ( .A(n2154), .B(IR_REG_2__SCAN_IN), .ZN(n4352) );
  NAND4_X2 U2318 ( .A1(n2325), .A2(n2324), .A3(n2323), .A4(n2322), .ZN(n3524)
         );
  AOI21_X2 U2319 ( .B1(n4123), .B2(n2471), .A(n2470), .ZN(n4107) );
  NAND2_X2 U2320 ( .A1(n2158), .A2(n2159), .ZN(n4123) );
  CLKBUF_X2 U2321 ( .A(n3300), .Z(n2061) );
  INV_X1 U2322 ( .A(n3524), .ZN(n2975) );
  NAND4_X1 U2323 ( .A1(n2356), .A2(n2355), .A3(n2354), .A4(n2353), .ZN(n3491)
         );
  INV_X1 U2324 ( .A(n2997), .ZN(n2910) );
  CLKBUF_X2 U2325 ( .A(n2338), .Z(n2060) );
  NAND2_X1 U2326 ( .A1(n2201), .A2(n2088), .ZN(n3399) );
  OR2_X1 U2327 ( .A1(n3445), .A2(n3438), .ZN(n2204) );
  OR2_X1 U2328 ( .A1(n2657), .A2(n4108), .ZN(n2128) );
  NAND2_X1 U2329 ( .A1(n4106), .A2(n2485), .ZN(n4089) );
  OR2_X1 U2330 ( .A1(n3139), .A2(n3138), .ZN(n3835) );
  OAI21_X1 U2331 ( .B1(n3087), .B2(n3670), .A(n3654), .ZN(n3099) );
  NAND2_X1 U2332 ( .A1(n2134), .A2(n3651), .ZN(n3087) );
  AOI21_X1 U2333 ( .B1(n2252), .B2(n2247), .A(n2067), .ZN(n2245) );
  CLKBUF_X1 U2334 ( .A(n3579), .Z(n3627) );
  XNOR2_X1 U2335 ( .A(n2870), .B(n2812), .ZN(n2810) );
  OAI21_X1 U2336 ( .B1(n2856), .B2(n2854), .A(n4187), .ZN(n3579) );
  OAI21_X1 U2337 ( .B1(n2806), .B2(n2805), .A(n2809), .ZN(n2870) );
  AND2_X1 U2338 ( .A1(n3644), .A2(n3647), .ZN(n3735) );
  AND2_X1 U2339 ( .A1(n3643), .A2(n3640), .ZN(n3733) );
  NOR2_X1 U2340 ( .A1(n2317), .A2(n2316), .ZN(n2319) );
  NAND2_X1 U2341 ( .A1(n2684), .A2(IR_REG_31__SCAN_IN), .ZN(n2675) );
  INV_X1 U2342 ( .A(n2895), .ZN(n2936) );
  INV_X4 U2343 ( .A(n2425), .ZN(n3692) );
  AND2_X1 U2344 ( .A1(n2620), .A2(n2673), .ZN(n3786) );
  INV_X1 U2345 ( .A(n2288), .ZN(n4344) );
  MUX2_X1 U2346 ( .A(n2750), .B(n2749), .S(IR_REG_28__SCAN_IN), .Z(n2346) );
  OAI211_X1 U2347 ( .C1(n2680), .C2(n2282), .A(n2679), .B(n2678), .ZN(n2703)
         );
  NAND2_X1 U2348 ( .A1(n2071), .A2(n2304), .ZN(n2750) );
  XNOR2_X1 U2349 ( .A(n2285), .B(n2257), .ZN(n2288) );
  NAND2_X1 U2350 ( .A1(n2284), .A2(IR_REG_31__SCAN_IN), .ZN(n2285) );
  AND4_X1 U2351 ( .A1(n2273), .A2(n2272), .A3(n2271), .A4(n2270), .ZN(n2274)
         );
  AND4_X1 U2352 ( .A1(n2276), .A2(n2482), .A3(n2275), .A4(n2467), .ZN(n2064)
         );
  NOR2_X1 U2353 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2320)
         );
  INV_X1 U2354 ( .A(IR_REG_16__SCAN_IN), .ZN(n2482) );
  INV_X1 U2355 ( .A(IR_REG_15__SCAN_IN), .ZN(n2467) );
  OAI21_X2 U2356 ( .B1(n4089), .B2(n2164), .A(n2162), .ZN(n4049) );
  NAND2_X1 U2357 ( .A1(n2295), .A2(n4344), .ZN(n2059) );
  OAI21_X2 U2358 ( .B1(n3589), .B2(n2236), .A(n2234), .ZN(n3441) );
  AOI21_X2 U2359 ( .B1(n3501), .B2(n3497), .A(n3499), .ZN(n3589) );
  OAI22_X2 U2360 ( .A1(n3062), .A2(n2179), .B1(n2178), .B2(n2181), .ZN(n3092)
         );
  XNOR2_X2 U2361 ( .A(n2675), .B(n2674), .ZN(n2683) );
  NAND2_X1 U2362 ( .A1(n4343), .A2(n4344), .ZN(n2342) );
  NAND2_X2 U2363 ( .A1(n2821), .A2(n2895), .ZN(n3188) );
  OR2_X4 U2364 ( .A1(n2683), .A2(n2682), .ZN(n2821) );
  INV_X1 U2365 ( .A(IR_REG_2__SCAN_IN), .ZN(n2268) );
  OR2_X1 U2366 ( .A1(n2506), .A2(n4649), .ZN(n2527) );
  NAND2_X1 U2367 ( .A1(n2221), .A2(n3237), .ZN(n2216) );
  AOI21_X1 U2368 ( .B1(n2219), .B2(n2221), .A(n2218), .ZN(n2217) );
  INV_X1 U2369 ( .A(n2225), .ZN(n2219) );
  INV_X1 U2370 ( .A(n3452), .ZN(n2218) );
  XNOR2_X1 U2371 ( .A(n2287), .B(n2286), .ZN(n2295) );
  OR2_X1 U2372 ( .A1(n3491), .A2(n3181), .ZN(n3644) );
  AND2_X1 U2373 ( .A1(n3786), .A2(n2707), .ZN(n2895) );
  INV_X1 U2374 ( .A(n2346), .ZN(n2425) );
  INV_X1 U2375 ( .A(n2058), .ZN(n2589) );
  INV_X1 U2376 ( .A(n3704), .ZN(n2590) );
  NOR2_X1 U2377 ( .A1(n2793), .A2(n2189), .ZN(n2775) );
  AND2_X1 U2378 ( .A1(n4350), .A2(REG2_REG_5__SCAN_IN), .ZN(n2189) );
  NOR2_X1 U2379 ( .A1(n2875), .A2(n2874), .ZN(n3130) );
  INV_X1 U2380 ( .A(n2143), .ZN(n3135) );
  OR2_X1 U2381 ( .A1(n3851), .A2(n3850), .ZN(n3867) );
  AND2_X1 U2382 ( .A1(n3927), .A2(n4130), .ZN(n2140) );
  OR2_X1 U2383 ( .A1(n2581), .A2(n3612), .ZN(n2603) );
  OR2_X1 U2384 ( .A1(n2527), .A2(n2525), .ZN(n2537) );
  AND2_X1 U2385 ( .A1(n2185), .A2(n2082), .ZN(n2184) );
  INV_X1 U2386 ( .A(IR_REG_5__SCAN_IN), .ZN(n2301) );
  INV_X1 U2387 ( .A(n2213), .ZN(n2212) );
  OAI21_X1 U2388 ( .B1(n2217), .B2(n2215), .A(n2214), .ZN(n2213) );
  INV_X1 U2389 ( .A(n3552), .ZN(n2214) );
  NAND2_X1 U2390 ( .A1(n2227), .A2(n2226), .ZN(n2225) );
  INV_X1 U2391 ( .A(n3574), .ZN(n2227) );
  INV_X1 U2392 ( .A(n3573), .ZN(n2226) );
  XNOR2_X1 U2393 ( .A(n2993), .B(n3343), .ZN(n3173) );
  NAND2_X1 U2394 ( .A1(n2992), .A2(n2991), .ZN(n2993) );
  INV_X1 U2395 ( .A(n2224), .ZN(n2222) );
  INV_X1 U2396 ( .A(n3188), .ZN(n3299) );
  OR2_X1 U2397 ( .A1(n3800), .A2(n3564), .ZN(n3979) );
  INV_X1 U2398 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2427) );
  OAI21_X1 U2399 ( .B1(n3061), .B2(n2399), .A(n2076), .ZN(n2182) );
  INV_X1 U2400 ( .A(n2399), .ZN(n2180) );
  NAND2_X1 U2401 ( .A1(n3806), .A2(n3431), .ZN(n2183) );
  NAND2_X1 U2402 ( .A1(n2942), .A2(n2952), .ZN(n3636) );
  NOR2_X1 U2403 ( .A1(n4032), .A2(n3420), .ZN(n2110) );
  AND2_X1 U2404 ( .A1(n4144), .A2(n2085), .ZN(n2160) );
  INV_X1 U2405 ( .A(n3073), .ZN(n2103) );
  INV_X1 U2406 ( .A(n3490), .ZN(n3187) );
  AND2_X1 U2407 ( .A1(n2281), .A2(n2282), .ZN(n2185) );
  NAND2_X1 U2408 ( .A1(n2668), .A2(n2185), .ZN(n2679) );
  INV_X1 U2409 ( .A(IR_REG_14__SCAN_IN), .ZN(n2276) );
  INV_X1 U2410 ( .A(IR_REG_23__SCAN_IN), .ZN(n2685) );
  AND2_X1 U2411 ( .A1(n2511), .A2(n2510), .ZN(n2615) );
  INV_X1 U2412 ( .A(IR_REG_18__SCAN_IN), .ZN(n2510) );
  NOR2_X1 U2413 ( .A1(n3198), .A2(n3196), .ZN(n2248) );
  NAND2_X1 U2414 ( .A1(n2251), .A2(n2250), .ZN(n2249) );
  INV_X1 U2415 ( .A(n3600), .ZN(n2251) );
  NOR2_X1 U2416 ( .A1(n3417), .A2(n2238), .ZN(n2237) );
  INV_X1 U2417 ( .A(n2241), .ZN(n2238) );
  NAND2_X1 U2418 ( .A1(n2945), .A2(n2944), .ZN(n2946) );
  NAND2_X1 U2419 ( .A1(n3574), .A2(n3573), .ZN(n2224) );
  NAND2_X1 U2420 ( .A1(n3572), .A2(n2225), .ZN(n2223) );
  NAND2_X1 U2421 ( .A1(n3183), .A2(n3185), .ZN(n3186) );
  AOI21_X1 U2422 ( .B1(n2207), .B2(n2209), .A(n3264), .ZN(n2205) );
  AND2_X1 U2423 ( .A1(n3262), .A2(n2210), .ZN(n2209) );
  OR2_X1 U2424 ( .A1(n2560), .A2(n3512), .ZN(n2571) );
  XNOR2_X1 U2425 ( .A(n4353), .B(n2115), .ZN(n3814) );
  INV_X1 U2426 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2115) );
  NAND2_X1 U2427 ( .A1(n2754), .A2(n2753), .ZN(n2756) );
  NAND2_X1 U2428 ( .A1(n2121), .A2(n2188), .ZN(n2187) );
  NAND2_X1 U2429 ( .A1(n2776), .A2(n2777), .ZN(n2188) );
  NAND2_X1 U2430 ( .A1(n2778), .A2(REG2_REG_6__SCAN_IN), .ZN(n2121) );
  NAND2_X1 U2431 ( .A1(n2796), .A2(n2763), .ZN(n2771) );
  NAND2_X1 U2432 ( .A1(n2113), .A2(n2089), .ZN(n3122) );
  INV_X1 U2433 ( .A(n3119), .ZN(n2113) );
  OR2_X1 U2434 ( .A1(n3130), .A2(n2095), .ZN(n2148) );
  NOR2_X1 U2435 ( .A1(n4410), .A2(n2147), .ZN(n2146) );
  NAND2_X1 U2436 ( .A1(n2120), .A2(n2118), .ZN(n3844) );
  NAND2_X1 U2437 ( .A1(n2119), .A2(n4189), .ZN(n2118) );
  AND2_X1 U2438 ( .A1(n3126), .A2(n2117), .ZN(n2116) );
  NAND2_X1 U2439 ( .A1(n3867), .A2(n3866), .ZN(n2190) );
  NAND2_X1 U2440 ( .A1(n4448), .A2(n4447), .ZN(n2197) );
  INV_X1 U2441 ( .A(n3985), .ZN(n3945) );
  NAND2_X1 U2442 ( .A1(n2536), .A2(REG3_REG_22__SCAN_IN), .ZN(n2549) );
  OR2_X1 U2443 ( .A1(n4110), .A2(n4098), .ZN(n2494) );
  AND2_X1 U2444 ( .A1(n2166), .A2(n2260), .ZN(n2165) );
  INV_X1 U2445 ( .A(n4072), .ZN(n2166) );
  OR2_X1 U2446 ( .A1(n2451), .A2(n2450), .ZN(n2460) );
  OR2_X1 U2447 ( .A1(n3580), .A2(n3457), .ZN(n2438) );
  AND2_X1 U2448 ( .A1(n3149), .A2(n3220), .ZN(n2177) );
  AND2_X1 U2449 ( .A1(n3144), .A2(n2086), .ZN(n2175) );
  OR2_X1 U2450 ( .A1(n3068), .A2(n3093), .ZN(n2263) );
  INV_X1 U2451 ( .A(n3535), .ZN(n3093) );
  INV_X1 U2452 ( .A(n2123), .ZN(n2122) );
  OAI21_X1 U2453 ( .B1(n2124), .B2(n3733), .A(n3647), .ZN(n2123) );
  NAND2_X1 U2454 ( .A1(n2821), .A2(n4464), .ZN(n2858) );
  NAND2_X1 U2455 ( .A1(n2626), .A2(n3876), .ZN(n4182) );
  OR2_X1 U2456 ( .A1(n2847), .A2(n4354), .ZN(n4127) );
  AND2_X1 U2457 ( .A1(n3062), .A2(n3061), .ZN(n4498) );
  NAND2_X1 U2458 ( .A1(n2681), .A2(n4345), .ZN(n2839) );
  INV_X1 U2459 ( .A(IR_REG_28__SCAN_IN), .ZN(n2283) );
  NOR2_X1 U2460 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2269)
         );
  AND2_X1 U2461 ( .A1(n2330), .A2(n2357), .ZN(n2755) );
  AOI21_X1 U2462 ( .B1(n2231), .B2(n2230), .A(n2087), .ZN(n2229) );
  INV_X1 U2463 ( .A(n3464), .ZN(n2230) );
  AND2_X1 U2464 ( .A1(n2634), .A2(n2633), .ZN(n3710) );
  AND2_X1 U2465 ( .A1(n2603), .A2(n2582), .ZN(n3934) );
  AND2_X1 U2466 ( .A1(n2951), .A2(n4354), .ZN(n3628) );
  NAND2_X1 U2467 ( .A1(n2596), .A2(n2595), .ZN(n3927) );
  XNOR2_X1 U2468 ( .A(n3122), .B(n4383), .ZN(n4380) );
  NAND2_X1 U2469 ( .A1(n4380), .A2(REG2_REG_10__SCAN_IN), .ZN(n4379) );
  XNOR2_X1 U2470 ( .A(n2148), .B(n4472), .ZN(n4375) );
  NOR2_X1 U2471 ( .A1(n4375), .A2(n4376), .ZN(n4374) );
  XNOR2_X1 U2472 ( .A(n3844), .B(n2192), .ZN(n4407) );
  NOR2_X1 U2473 ( .A1(n4407), .A2(n4159), .ZN(n4406) );
  XNOR2_X1 U2474 ( .A(n2190), .B(n4468), .ZN(n4419) );
  NAND2_X1 U2475 ( .A1(n4419), .A2(n4116), .ZN(n4418) );
  NAND2_X1 U2476 ( .A1(n4430), .A2(n4431), .ZN(n4429) );
  INV_X1 U2477 ( .A(n3621), .ZN(n2210) );
  AND2_X1 U2478 ( .A1(n3477), .A2(n2208), .ZN(n2207) );
  NAND2_X1 U2479 ( .A1(n3263), .A2(n3621), .ZN(n2208) );
  INV_X1 U2480 ( .A(n2497), .ZN(n2495) );
  OR2_X1 U2481 ( .A1(n2486), .A2(n4556), .ZN(n2497) );
  INV_X1 U2482 ( .A(n3834), .ZN(n2147) );
  INV_X1 U2483 ( .A(n3842), .ZN(n2117) );
  AND2_X1 U2484 ( .A1(n3858), .A2(n3857), .ZN(n3859) );
  INV_X1 U2485 ( .A(n2579), .ZN(n2171) );
  NOR2_X1 U2486 ( .A1(n3757), .A2(n2127), .ZN(n2126) );
  INV_X1 U2487 ( .A(n2129), .ZN(n2127) );
  AOI21_X1 U2488 ( .B1(n3728), .B2(n2131), .A(n2130), .ZN(n2129) );
  INV_X1 U2489 ( .A(n3659), .ZN(n2131) );
  NAND2_X1 U2490 ( .A1(n2472), .A2(REG3_REG_16__SCAN_IN), .ZN(n2486) );
  INV_X1 U2491 ( .A(n2474), .ZN(n2472) );
  OR2_X1 U2492 ( .A1(n2460), .A2(n3625), .ZN(n2474) );
  OR2_X1 U2493 ( .A1(n2403), .A2(n2291), .ZN(n2404) );
  INV_X1 U2494 ( .A(n3643), .ZN(n2125) );
  NAND2_X1 U2495 ( .A1(n2103), .A2(n2102), .ZN(n3104) );
  NOR2_X1 U2496 ( .A1(n2105), .A2(n3409), .ZN(n2102) );
  NOR2_X1 U2497 ( .A1(n3692), .A2(n2597), .ZN(n3915) );
  INV_X1 U2498 ( .A(n3609), .ZN(n2232) );
  INV_X1 U2499 ( .A(n2211), .ZN(n3238) );
  OAI21_X1 U2500 ( .B1(n3572), .B2(n2216), .A(n2212), .ZN(n2211) );
  NAND2_X1 U2501 ( .A1(n2202), .A2(n3438), .ZN(n2200) );
  AOI22_X1 U2502 ( .A1(n3531), .A2(n3532), .B1(n3216), .B2(n3215), .ZN(n3408)
         );
  NAND2_X1 U2503 ( .A1(n2987), .A2(n2988), .ZN(n2989) );
  NAND2_X1 U2504 ( .A1(n3589), .A2(n2240), .ZN(n2239) );
  NAND2_X1 U2505 ( .A1(n3587), .A2(n3586), .ZN(n2241) );
  INV_X1 U2506 ( .A(n3202), .ZN(n2254) );
  INV_X1 U2507 ( .A(n3203), .ZN(n2253) );
  NAND2_X1 U2508 ( .A1(n2547), .A2(REG3_REG_23__SCAN_IN), .ZN(n2560) );
  NAND2_X1 U2509 ( .A1(n2822), .A2(REG1_REG_0__SCAN_IN), .ZN(n2826) );
  AOI21_X1 U2510 ( .B1(n2237), .B2(n2242), .A(n2235), .ZN(n2234) );
  INV_X1 U2511 ( .A(n2237), .ZN(n2236) );
  INV_X1 U2512 ( .A(n3280), .ZN(n2235) );
  NOR2_X1 U2513 ( .A1(n3563), .A2(n2203), .ZN(n2202) );
  INV_X1 U2514 ( .A(n3439), .ZN(n2203) );
  NAND2_X1 U2515 ( .A1(n2628), .A2(REG2_REG_1__SCAN_IN), .ZN(n2335) );
  AND2_X1 U2516 ( .A1(n2613), .A2(n2612), .ZN(n3381) );
  NAND2_X1 U2517 ( .A1(n2315), .A2(n2314), .ZN(n2316) );
  AND2_X1 U2518 ( .A1(n3814), .A2(n2081), .ZN(n3811) );
  NAND2_X1 U2519 ( .A1(n2142), .A2(n2757), .ZN(n2759) );
  AOI21_X1 U2520 ( .B1(n2872), .B2(n4348), .A(n2871), .ZN(n2875) );
  NAND2_X1 U2521 ( .A1(n4389), .A2(n3124), .ZN(n3125) );
  OR2_X1 U2522 ( .A1(n4384), .A2(n2144), .ZN(n2143) );
  AND2_X1 U2523 ( .A1(n4470), .A2(REG1_REG_11__SCAN_IN), .ZN(n2144) );
  NOR2_X1 U2524 ( .A1(n4403), .A2(n3836), .ZN(n3838) );
  OR2_X1 U2525 ( .A1(n3838), .A2(n3839), .ZN(n3858) );
  INV_X1 U2526 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3625) );
  XNOR2_X1 U2527 ( .A(n3859), .B(n2484), .ZN(n4417) );
  NAND2_X1 U2528 ( .A1(n4429), .A2(n2098), .ZN(n4442) );
  OAI21_X1 U2529 ( .B1(n3870), .B2(REG1_REG_17__SCAN_IN), .A(n4426), .ZN(n4446) );
  NOR2_X1 U2530 ( .A1(n3692), .A2(n3691), .ZN(n3898) );
  OAI21_X1 U2531 ( .B1(n3939), .B2(n2169), .A(n2168), .ZN(n3894) );
  OR2_X1 U2532 ( .A1(n2075), .A2(n2170), .ZN(n2168) );
  OR2_X1 U2533 ( .A1(n2075), .A2(n2580), .ZN(n2169) );
  NOR2_X1 U2534 ( .A1(n2598), .A2(n2171), .ZN(n2170) );
  NAND2_X1 U2535 ( .A1(n2172), .A2(n2579), .ZN(n3921) );
  OR2_X1 U2536 ( .A1(n3939), .A2(n2580), .ZN(n2172) );
  NOR2_X1 U2537 ( .A1(n3692), .A2(n2545), .ZN(n4007) );
  AOI21_X1 U2538 ( .B1(n2165), .B2(n2163), .A(n2094), .ZN(n2162) );
  INV_X1 U2539 ( .A(n2165), .ZN(n2164) );
  INV_X1 U2540 ( .A(n2494), .ZN(n2163) );
  INV_X1 U2541 ( .A(n3802), .ZN(n4093) );
  NAND2_X1 U2542 ( .A1(n2128), .A2(n2129), .ZN(n4090) );
  NAND2_X1 U2543 ( .A1(n2657), .A2(n3659), .ZN(n4109) );
  INV_X1 U2544 ( .A(n3480), .ZN(n4118) );
  AOI21_X1 U2545 ( .B1(n2160), .B2(n2070), .A(n2091), .ZN(n2159) );
  INV_X1 U2546 ( .A(n2441), .ZN(n2440) );
  OR2_X1 U2547 ( .A1(n2428), .A2(n2427), .ZN(n2441) );
  AOI21_X1 U2548 ( .B1(n2175), .B2(n2177), .A(n2092), .ZN(n2174) );
  NAND2_X1 U2549 ( .A1(n3067), .A2(n3653), .ZN(n2134) );
  INV_X1 U2550 ( .A(n2183), .ZN(n2178) );
  NAND2_X1 U2551 ( .A1(n2180), .A2(n2183), .ZN(n2179) );
  INV_X1 U2552 ( .A(n2182), .ZN(n2181) );
  INV_X1 U2553 ( .A(n4176), .ZN(n4130) );
  INV_X1 U2554 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2387) );
  NAND2_X1 U2555 ( .A1(n2903), .A2(n3643), .ZN(n3002) );
  AND2_X1 U2556 ( .A1(n2910), .A2(n2112), .ZN(n3038) );
  AND2_X1 U2557 ( .A1(n2925), .A2(n3181), .ZN(n2112) );
  NAND2_X1 U2558 ( .A1(n2910), .A2(n2925), .ZN(n3001) );
  NAND2_X1 U2559 ( .A1(n2904), .A2(n3733), .ZN(n2903) );
  INV_X1 U2560 ( .A(n4127), .ZN(n4173) );
  NAND2_X1 U2561 ( .A1(n2133), .A2(n2132), .ZN(n2919) );
  AND2_X1 U2562 ( .A1(n2889), .A2(n3637), .ZN(n3736) );
  NOR2_X1 U2563 ( .A1(n3931), .A2(n2106), .ZN(n4204) );
  OR2_X1 U2564 ( .A1(n2107), .A2(n3892), .ZN(n2106) );
  OR2_X1 U2565 ( .A1(n3915), .A2(n3898), .ZN(n2107) );
  NOR2_X1 U2566 ( .A1(n3931), .A2(n3915), .ZN(n3914) );
  INV_X1 U2567 ( .A(n3926), .ZN(n3932) );
  OR2_X1 U2568 ( .A1(n3952), .A2(n3926), .ZN(n3931) );
  NOR2_X1 U2569 ( .A1(n3692), .A2(n2578), .ZN(n3950) );
  OR2_X1 U2570 ( .A1(n3967), .A2(n3950), .ZN(n3952) );
  NOR2_X1 U2571 ( .A1(n2062), .A2(n3988), .ZN(n3989) );
  NAND2_X1 U2572 ( .A1(n2110), .A2(n4019), .ZN(n2109) );
  INV_X1 U2573 ( .A(n3446), .ZN(n4019) );
  NOR2_X1 U2574 ( .A1(n4080), .A2(n2108), .ZN(n4038) );
  INV_X1 U2575 ( .A(n2110), .ZN(n2108) );
  OR2_X1 U2576 ( .A1(n4100), .A2(n4079), .ZN(n4080) );
  INV_X1 U2577 ( .A(n3420), .ZN(n4064) );
  NOR2_X1 U2578 ( .A1(n4080), .A2(n3420), .ZN(n4062) );
  OR2_X1 U2579 ( .A1(n4256), .A2(n4098), .ZN(n4100) );
  NAND2_X1 U2580 ( .A1(n4134), .A2(n4118), .ZN(n4256) );
  NAND2_X1 U2581 ( .A1(n4184), .A2(n2084), .ZN(n4157) );
  NAND2_X1 U2582 ( .A1(n2161), .A2(n2160), .ZN(n4143) );
  AND2_X1 U2583 ( .A1(n2161), .A2(n2085), .ZN(n4145) );
  OR2_X1 U2584 ( .A1(n4165), .A2(n2070), .ZN(n2161) );
  NAND2_X1 U2585 ( .A1(n4184), .A2(n4183), .ZN(n4186) );
  AND2_X1 U2586 ( .A1(n3166), .A2(n3232), .ZN(n4184) );
  INV_X1 U2587 ( .A(n3457), .ZN(n3232) );
  NOR2_X1 U2588 ( .A1(n3104), .A2(n3578), .ZN(n3166) );
  NAND2_X1 U2589 ( .A1(n2103), .A2(n2104), .ZN(n3105) );
  OR2_X1 U2590 ( .A1(n3058), .A2(n3371), .ZN(n3073) );
  NOR2_X1 U2591 ( .A1(n3073), .A2(n3431), .ZN(n3094) );
  NOR2_X1 U2592 ( .A1(n2997), .A2(n3523), .ZN(n2111) );
  OR2_X1 U2593 ( .A1(n3039), .A2(n3603), .ZN(n3058) );
  AND2_X1 U2594 ( .A1(n2885), .A2(n2974), .ZN(n2925) );
  NAND2_X1 U2595 ( .A1(n2704), .A2(n2732), .ZN(n2881) );
  OR2_X1 U2596 ( .A1(n2839), .A2(D_REG_0__SCAN_IN), .ZN(n2704) );
  AND3_X1 U2597 ( .A1(n2702), .A2(n2701), .A3(n2700), .ZN(n2710) );
  AND2_X1 U2598 ( .A1(n2679), .A2(n2305), .ZN(n2749) );
  AND2_X1 U2599 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2305)
         );
  NAND2_X1 U2600 ( .A1(n2282), .A2(n2480), .ZN(n2678) );
  XNOR2_X1 U2601 ( .A(n2625), .B(n2624), .ZN(n2635) );
  INV_X1 U2602 ( .A(IR_REG_22__SCAN_IN), .ZN(n2624) );
  NAND2_X1 U2603 ( .A1(n2673), .A2(IR_REG_31__SCAN_IN), .ZN(n2625) );
  NOR2_X1 U2604 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2614)
         );
  XNOR2_X1 U2605 ( .A(n2623), .B(n2622), .ZN(n2707) );
  INV_X1 U2606 ( .A(IR_REG_20__SCAN_IN), .ZN(n2622) );
  NAND2_X1 U2607 ( .A1(n2621), .A2(IR_REG_31__SCAN_IN), .ZN(n2623) );
  OR2_X1 U2608 ( .A1(n2615), .A2(n2480), .ZN(n2513) );
  INV_X1 U2609 ( .A(IR_REG_19__SCAN_IN), .ZN(n2512) );
  NAND2_X1 U2610 ( .A1(n2513), .A2(n2512), .ZN(n2621) );
  OR2_X1 U2611 ( .A1(n2423), .A2(IR_REG_10__SCAN_IN), .ZN(n2424) );
  INV_X1 U2612 ( .A(IR_REG_7__SCAN_IN), .ZN(n2394) );
  NAND2_X1 U2613 ( .A1(n2249), .A2(n2246), .ZN(n3368) );
  INV_X1 U2614 ( .A(n2248), .ZN(n2246) );
  NOR2_X1 U2615 ( .A1(n3692), .A2(n2556), .ZN(n3988) );
  OR2_X1 U2616 ( .A1(n3338), .A2(n3337), .ZN(n3339) );
  NAND2_X1 U2617 ( .A1(n2223), .A2(n2224), .ZN(n3455) );
  NAND2_X1 U2618 ( .A1(n3708), .A2(DATAI_24_), .ZN(n3968) );
  NAND2_X1 U2619 ( .A1(n2204), .A2(n3439), .ZN(n3562) );
  INV_X1 U2620 ( .A(n2965), .ZN(n2974) );
  INV_X1 U2621 ( .A(n3628), .ZN(n3567) );
  INV_X1 U2622 ( .A(n3619), .ZN(n3623) );
  NAND2_X1 U2623 ( .A1(n2233), .A2(n3465), .ZN(n3611) );
  NAND2_X1 U2624 ( .A1(n3466), .A2(n3464), .ZN(n2233) );
  INV_X1 U2625 ( .A(n3566), .ZN(n3629) );
  OR2_X1 U2626 ( .A1(n3188), .A2(n2843), .ZN(n3793) );
  NAND2_X1 U2627 ( .A1(n2587), .A2(n2586), .ZN(n3947) );
  NAND2_X1 U2628 ( .A1(n2566), .A2(n2565), .ZN(n3985) );
  NAND2_X1 U2629 ( .A1(n2544), .A2(n2543), .ZN(n3800) );
  NAND2_X1 U2630 ( .A1(n2533), .A2(n2532), .ZN(n4001) );
  NAND2_X1 U2631 ( .A1(n2522), .A2(n2521), .ZN(n4059) );
  OR2_X1 U2632 ( .A1(n2609), .A2(n2352), .ZN(n2353) );
  OR2_X1 U2633 ( .A1(n2058), .A2(REG3_REG_3__SCAN_IN), .ZN(n2324) );
  NOR2_X1 U2634 ( .A1(n3811), .A2(n2114), .ZN(n3828) );
  AND2_X1 U2635 ( .A1(n4353), .A2(REG2_REG_1__SCAN_IN), .ZN(n2114) );
  XNOR2_X1 U2636 ( .A(n2744), .B(n2791), .ZN(n2191) );
  XNOR2_X1 U2637 ( .A(n2759), .B(n2758), .ZN(n2831) );
  XNOR2_X1 U2638 ( .A(n2775), .B(n2777), .ZN(n2778) );
  NAND2_X1 U2639 ( .A1(n2187), .A2(n2186), .ZN(n2804) );
  INV_X1 U2640 ( .A(n2779), .ZN(n2186) );
  INV_X1 U2641 ( .A(n2187), .ZN(n2780) );
  NAND2_X1 U2642 ( .A1(n2773), .A2(n2772), .ZN(n2806) );
  NOR2_X1 U2643 ( .A1(n2868), .A2(n2867), .ZN(n3119) );
  NAND2_X1 U2644 ( .A1(n4379), .A2(n3123), .ZN(n4390) );
  NAND2_X1 U2645 ( .A1(n4390), .A2(n4391), .ZN(n4389) );
  NOR2_X1 U2646 ( .A1(n3133), .A2(n4374), .ZN(n4386) );
  INV_X1 U2647 ( .A(n2148), .ZN(n3132) );
  NOR2_X1 U2648 ( .A1(n4386), .A2(n4385), .ZN(n4384) );
  XNOR2_X1 U2649 ( .A(n3125), .B(n4469), .ZN(n4400) );
  NAND2_X1 U2650 ( .A1(n4400), .A2(REG2_REG_12__SCAN_IN), .ZN(n4399) );
  XNOR2_X1 U2651 ( .A(n2143), .B(n3134), .ZN(n4396) );
  NOR2_X1 U2652 ( .A1(n4396), .A2(n4536), .ZN(n4395) );
  NAND2_X1 U2653 ( .A1(n4399), .A2(n3126), .ZN(n3843) );
  NOR2_X1 U2654 ( .A1(n4406), .A2(n3845), .ZN(n3851) );
  NAND2_X1 U2655 ( .A1(n4418), .A2(n3869), .ZN(n4430) );
  INV_X1 U2656 ( .A(n2190), .ZN(n3868) );
  NOR2_X1 U2657 ( .A1(n4442), .A2(n4441), .ZN(n4439) );
  NAND2_X1 U2658 ( .A1(n2199), .A2(n4433), .ZN(n2198) );
  NAND2_X1 U2659 ( .A1(n4442), .A2(n4441), .ZN(n2199) );
  NOR2_X1 U2660 ( .A1(n2196), .A2(n2195), .ZN(n2194) );
  NOR2_X1 U2661 ( .A1(n4451), .A2(n4450), .ZN(n2195) );
  NAND2_X1 U2662 ( .A1(n2197), .A2(n4449), .ZN(n2196) );
  NAND2_X1 U2663 ( .A1(n2153), .A2(n2152), .ZN(n4443) );
  INV_X1 U2664 ( .A(n4445), .ZN(n2152) );
  INV_X1 U2665 ( .A(n4446), .ZN(n2153) );
  AOI21_X1 U2666 ( .B1(n4446), .B2(n4445), .A(n4444), .ZN(n2151) );
  AOI21_X1 U2667 ( .B1(n2063), .B2(n3898), .A(n4204), .ZN(n4212) );
  XNOR2_X1 U2668 ( .A(n3894), .B(n3893), .ZN(n3366) );
  AOI21_X1 U2669 ( .B1(n2065), .B2(n4179), .A(n2139), .ZN(n3359) );
  OR2_X1 U2670 ( .A1(n2667), .A2(n2140), .ZN(n2139) );
  NAND2_X1 U2671 ( .A1(n2167), .A2(n2260), .ZN(n4071) );
  NAND2_X1 U2672 ( .A1(n4089), .A2(n2494), .ZN(n2167) );
  NAND2_X1 U2673 ( .A1(n2176), .A2(n2175), .ZN(n3143) );
  AND2_X1 U2674 ( .A1(n2176), .A2(n2086), .ZN(n3145) );
  OR2_X1 U2675 ( .A1(n3103), .A2(n2177), .ZN(n2176) );
  NOR2_X1 U2676 ( .A1(n4498), .A2(n2399), .ZN(n3072) );
  AND2_X1 U2677 ( .A1(n4357), .A2(n3023), .ZN(n3897) );
  OR2_X1 U2678 ( .A1(n2858), .A2(n2853), .ZN(n4187) );
  INV_X1 U2679 ( .A(n4187), .ZN(n4456) );
  NAND2_X1 U2680 ( .A1(n3359), .A2(n2137), .ZN(n2711) );
  NAND2_X1 U2681 ( .A1(n2138), .A2(n4508), .ZN(n2137) );
  INV_X1 U2682 ( .A(n3366), .ZN(n2138) );
  INV_X1 U2683 ( .A(n4519), .ZN(n4517) );
  NAND2_X1 U2684 ( .A1(n2711), .A2(n4511), .ZN(n2136) );
  NOR2_X1 U2685 ( .A1(n2256), .A2(IR_REG_26__SCAN_IN), .ZN(n2255) );
  NAND2_X1 U2686 ( .A1(n2082), .A2(n2257), .ZN(n2256) );
  XNOR2_X1 U2687 ( .A(n2627), .B(IR_REG_28__SCAN_IN), .ZN(n4354) );
  NAND2_X1 U2688 ( .A1(n2672), .A2(n2677), .ZN(n2718) );
  INV_X1 U2689 ( .A(n2635), .ZN(n3794) );
  NAND2_X1 U2690 ( .A1(n2621), .A2(n2514), .ZN(n3876) );
  OR2_X1 U2691 ( .A1(n2513), .A2(n2512), .ZN(n2514) );
  XNOR2_X1 U2692 ( .A(n2435), .B(IR_REG_11__SCAN_IN), .ZN(n4470) );
  NOR2_X1 U2693 ( .A1(n2370), .A2(n2369), .ZN(n4350) );
  INV_X1 U2694 ( .A(n2755), .ZN(n2791) );
  NAND2_X1 U2695 ( .A1(n2155), .A2(IR_REG_31__SCAN_IN), .ZN(n2154) );
  INV_X2 U2696 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U2697 ( .A1(n2150), .A2(n2149), .ZN(U3258) );
  INV_X1 U2698 ( .A(n2193), .ZN(n2149) );
  NAND2_X1 U2699 ( .A1(n4443), .A2(n2151), .ZN(n2150) );
  OAI21_X1 U2700 ( .B1(n4439), .B2(n2198), .A(n2194), .ZN(n2193) );
  OR2_X1 U2701 ( .A1(n2073), .A2(n4007), .ZN(n2062) );
  OR2_X2 U2702 ( .A1(n3311), .A2(n4496), .ZN(n3340) );
  OR2_X1 U2703 ( .A1(n3261), .A2(n3262), .ZN(n3474) );
  OR3_X1 U2704 ( .A1(n3931), .A2(n3915), .A3(n3892), .ZN(n2063) );
  NAND2_X1 U2705 ( .A1(n2239), .A2(n2241), .ZN(n3416) );
  XNOR2_X1 U2706 ( .A(n3893), .B(n3885), .ZN(n2065) );
  AND2_X1 U2707 ( .A1(n2970), .A2(n2969), .ZN(n2066) );
  AND2_X1 U2708 ( .A1(n2254), .A2(n2253), .ZN(n2067) );
  AND2_X1 U2709 ( .A1(n2791), .A2(n2745), .ZN(n2068) );
  AND2_X1 U2710 ( .A1(n4344), .A2(REG3_REG_1__SCAN_IN), .ZN(n2069) );
  AND2_X1 U2711 ( .A1(n4151), .A2(n4183), .ZN(n2070) );
  INV_X1 U2712 ( .A(n3237), .ZN(n2215) );
  INV_X1 U2713 ( .A(n2887), .ZN(n2133) );
  INV_X1 U2714 ( .A(n3626), .ZN(n2100) );
  INV_X1 U2715 ( .A(n4410), .ZN(n2192) );
  OR2_X1 U2716 ( .A1(n2679), .A2(IR_REG_27__SCAN_IN), .ZN(n2071) );
  AND2_X1 U2717 ( .A1(n2326), .A2(n2269), .ZN(n2300) );
  AND2_X1 U2718 ( .A1(n2204), .A2(n2202), .ZN(n2072) );
  OR2_X1 U2719 ( .A1(n4080), .A2(n2109), .ZN(n2073) );
  NAND2_X1 U2720 ( .A1(n4343), .A2(n2288), .ZN(n2338) );
  INV_X1 U2721 ( .A(n2988), .ZN(n2966) );
  NAND3_X1 U2722 ( .A1(n2345), .A2(n2344), .A3(n2343), .ZN(n2825) );
  AND4_X1 U2723 ( .A1(n2280), .A2(n2279), .A3(n2278), .A4(n2277), .ZN(n2074)
         );
  AND2_X1 U2724 ( .A1(n2320), .A2(n2268), .ZN(n2326) );
  NOR2_X1 U2725 ( .A1(n2601), .A2(n2600), .ZN(n2075) );
  OR2_X1 U2726 ( .A1(n3806), .A2(n3431), .ZN(n2076) );
  AND2_X1 U2727 ( .A1(n2668), .A2(n2281), .ZN(n2671) );
  NOR2_X1 U2728 ( .A1(n3367), .A2(n2248), .ZN(n2247) );
  AND2_X1 U2729 ( .A1(n2239), .A2(n2237), .ZN(n2077) );
  AND2_X1 U2730 ( .A1(n2942), .A2(n2943), .ZN(n2078) );
  XNOR2_X1 U2731 ( .A(n2946), .B(n3334), .ZN(n2967) );
  AND4_X1 U2732 ( .A1(n2300), .A2(n2074), .A3(n2274), .A4(n2064), .ZN(n2668)
         );
  AND2_X1 U2733 ( .A1(n2136), .A2(n2135), .ZN(n2079) );
  INV_X1 U2734 ( .A(n2252), .ZN(n2250) );
  AND2_X1 U2735 ( .A1(n3198), .A2(n3196), .ZN(n2252) );
  INV_X1 U2736 ( .A(IR_REG_31__SCAN_IN), .ZN(n2480) );
  AND2_X1 U2737 ( .A1(n3835), .A2(n3834), .ZN(n2080) );
  AND2_X1 U2738 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2081)
         );
  AND2_X1 U2739 ( .A1(n2283), .A2(n2258), .ZN(n2082) );
  OR2_X1 U2740 ( .A1(n2791), .A2(n2745), .ZN(n2083) );
  INV_X1 U2741 ( .A(IR_REG_27__SCAN_IN), .ZN(n2258) );
  OR2_X1 U2742 ( .A1(n2639), .A2(n2125), .ZN(n2124) );
  INV_X1 U2743 ( .A(IR_REG_26__SCAN_IN), .ZN(n2282) );
  INV_X1 U2744 ( .A(IR_REG_29__SCAN_IN), .ZN(n2257) );
  NAND2_X1 U2745 ( .A1(n3261), .A2(n3262), .ZN(n3475) );
  INV_X1 U2746 ( .A(n3188), .ZN(n3331) );
  INV_X1 U2747 ( .A(n2889), .ZN(n2132) );
  AND2_X1 U2748 ( .A1(n4183), .A2(n2459), .ZN(n2084) );
  NAND2_X1 U2749 ( .A1(n2300), .A2(n2274), .ZN(n2447) );
  INV_X1 U2750 ( .A(n3679), .ZN(n2130) );
  NAND2_X1 U2751 ( .A1(n3803), .A2(n4172), .ZN(n2085) );
  NAND2_X1 U2752 ( .A1(n3804), .A2(n3409), .ZN(n2086) );
  AND2_X1 U2753 ( .A1(n3330), .A2(n3329), .ZN(n2087) );
  AND2_X1 U2754 ( .A1(n3307), .A2(n2200), .ZN(n2088) );
  INV_X1 U2755 ( .A(n2242), .ZN(n2240) );
  NOR2_X1 U2756 ( .A1(n3587), .A2(n3586), .ZN(n2242) );
  OR2_X1 U2757 ( .A1(n3120), .A2(n3121), .ZN(n2089) );
  AND2_X1 U2758 ( .A1(n2084), .A2(n2100), .ZN(n2090) );
  NOR2_X1 U2759 ( .A1(n4174), .A2(n4155), .ZN(n2091) );
  NOR2_X1 U2760 ( .A1(n3458), .A2(n3578), .ZN(n2092) );
  AND2_X1 U2761 ( .A1(n2167), .A2(n2165), .ZN(n2093) );
  INV_X1 U2762 ( .A(n2105), .ZN(n2104) );
  NAND2_X1 U2763 ( .A1(n3093), .A2(n3207), .ZN(n2105) );
  AND2_X1 U2764 ( .A1(n4093), .A2(n3272), .ZN(n2094) );
  NOR2_X1 U2765 ( .A1(n2503), .A2(IR_REG_17__SCAN_IN), .ZN(n2511) );
  INV_X1 U2766 ( .A(n2221), .ZN(n2220) );
  NOR2_X1 U2767 ( .A1(n2222), .A2(n3451), .ZN(n2221) );
  AND2_X1 U2768 ( .A1(n3131), .A2(REG1_REG_9__SCAN_IN), .ZN(n2095) );
  AND2_X1 U2769 ( .A1(n2232), .A2(n3465), .ZN(n2231) );
  NAND2_X1 U2770 ( .A1(n2244), .A2(n2245), .ZN(n3426) );
  INV_X1 U2771 ( .A(n4032), .ZN(n4040) );
  NOR2_X1 U2772 ( .A1(n3692), .A2(n2523), .ZN(n4032) );
  INV_X1 U2773 ( .A(n2101), .ZN(n4134) );
  NAND2_X1 U2774 ( .A1(n4184), .A2(n2090), .ZN(n2101) );
  AND2_X1 U2775 ( .A1(n2635), .A2(n2688), .ZN(n2708) );
  INV_X1 U2776 ( .A(n2942), .ZN(n2817) );
  INV_X1 U2777 ( .A(n4440), .ZN(n4433) );
  AND2_X2 U2778 ( .A1(n2710), .A2(n2881), .ZN(n4511) );
  NAND2_X1 U2779 ( .A1(n2821), .A2(n2936), .ZN(n3311) );
  AND2_X1 U2780 ( .A1(n2666), .A2(n2665), .ZN(n4132) );
  NAND2_X1 U2781 ( .A1(n3636), .A2(n3638), .ZN(n2887) );
  OR2_X1 U2782 ( .A1(n3210), .A2(n3209), .ZN(n2096) );
  AND2_X1 U2783 ( .A1(n4182), .A2(n4482), .ZN(n4499) );
  OR2_X1 U2784 ( .A1(n2192), .A2(n3834), .ZN(n2097) );
  INV_X1 U2785 ( .A(IR_REG_30__SCAN_IN), .ZN(n2286) );
  INV_X1 U2786 ( .A(n3841), .ZN(n2119) );
  OR2_X1 U2787 ( .A1(n3870), .A2(REG2_REG_17__SCAN_IN), .ZN(n2098) );
  AND2_X1 U2788 ( .A1(n2671), .A2(n2255), .ZN(n3355) );
  OAI211_X1 U2789 ( .C1(n2609), .C2(n4247), .A(n2509), .B(n2508), .ZN(n2099)
         );
  NAND3_X1 U2790 ( .A1(n3187), .A2(n2925), .A3(n2111), .ZN(n3039) );
  XNOR2_X2 U2791 ( .A(n2334), .B(IR_REG_1__SCAN_IN), .ZN(n4353) );
  NAND2_X1 U2792 ( .A1(n4399), .A2(n2116), .ZN(n2120) );
  OAI21_X1 U2793 ( .B1(n2904), .B2(n2124), .A(n2122), .ZN(n3032) );
  NAND2_X1 U2794 ( .A1(n2128), .A2(n2126), .ZN(n4029) );
  OR2_X2 U2795 ( .A1(n2942), .A2(n2952), .ZN(n3638) );
  NAND2_X1 U2796 ( .A1(n4510), .A2(REG0_REG_28__SCAN_IN), .ZN(n2135) );
  XNOR2_X2 U2797 ( .A(n2287), .B(IR_REG_30__SCAN_IN), .ZN(n4343) );
  NAND2_X1 U2798 ( .A1(n2069), .A2(n4343), .ZN(n2141) );
  OAI21_X1 U2799 ( .B1(n2333), .B2(n4343), .A(n2141), .ZN(n2156) );
  NAND2_X1 U2800 ( .A1(n2831), .A2(REG1_REG_4__SCAN_IN), .ZN(n2761) );
  NAND2_X1 U2801 ( .A1(n2786), .A2(REG1_REG_3__SCAN_IN), .ZN(n2142) );
  NAND2_X1 U2802 ( .A1(n3835), .A2(n2146), .ZN(n2145) );
  OAI211_X1 U2803 ( .C1(n3835), .C2(n2192), .A(n2097), .B(n2145), .ZN(n4404)
         );
  INV_X1 U2804 ( .A(n2320), .ZN(n2155) );
  NOR2_X1 U2805 ( .A1(n2810), .A2(n2309), .ZN(n2871) );
  INV_X1 U2806 ( .A(n2156), .ZN(n2157) );
  AOI21_X2 U2807 ( .B1(n2887), .B2(n2888), .A(n2078), .ZN(n2917) );
  NAND2_X1 U2808 ( .A1(n4165), .A2(n2160), .ZN(n2158) );
  NAND2_X1 U2809 ( .A1(n3103), .A2(n2175), .ZN(n2173) );
  NAND2_X1 U2810 ( .A1(n2173), .A2(n2174), .ZN(n3165) );
  NAND2_X1 U2811 ( .A1(n2668), .A2(n2184), .ZN(n2284) );
  AOI21_X1 U2812 ( .B1(n2744), .B2(n2083), .A(n2068), .ZN(n2746) );
  XNOR2_X1 U2813 ( .A(n2191), .B(REG2_REG_3__SCAN_IN), .ZN(n2787) );
  NAND2_X1 U2814 ( .A1(n3445), .A2(n2202), .ZN(n2201) );
  NAND2_X1 U2815 ( .A1(n3261), .A2(n2207), .ZN(n2206) );
  NAND2_X2 U2816 ( .A1(n2206), .A2(n2205), .ZN(n3501) );
  OAI21_X1 U2817 ( .B1(n3572), .B2(n2220), .A(n2217), .ZN(n3554) );
  NAND2_X1 U2818 ( .A1(n3317), .A2(n3509), .ZN(n3466) );
  NAND2_X1 U2819 ( .A1(n2228), .A2(n2229), .ZN(n3378) );
  NAND3_X1 U2820 ( .A1(n3317), .A2(n2231), .A3(n3509), .ZN(n2228) );
  NAND3_X1 U2821 ( .A1(n2300), .A2(n2274), .A3(n2064), .ZN(n2503) );
  NAND2_X1 U2822 ( .A1(n2243), .A2(n3427), .ZN(n3531) );
  NAND3_X1 U2823 ( .A1(n2244), .A2(n2096), .A3(n2245), .ZN(n2243) );
  NAND2_X1 U2824 ( .A1(n2247), .A2(n3600), .ZN(n2244) );
  OR2_X1 U2825 ( .A1(n3921), .A2(n3902), .ZN(n3904) );
  NAND2_X1 U2826 ( .A1(n2619), .A2(n2618), .ZN(n2673) );
  INV_X1 U2827 ( .A(n2617), .ZN(n2619) );
  NAND2_X1 U2828 ( .A1(n3399), .A2(n2266), .ZN(n3508) );
  NAND2_X1 U2829 ( .A1(n3704), .A2(REG0_REG_1__SCAN_IN), .ZN(n2336) );
  INV_X1 U2830 ( .A(n3003), .ZN(n3004) );
  NOR2_X1 U2831 ( .A1(n2949), .A2(n2950), .ZN(n2971) );
  AND2_X1 U2832 ( .A1(n4034), .A2(n4019), .ZN(n2259) );
  OR2_X1 U2833 ( .A1(n4076), .A2(n4092), .ZN(n2260) );
  OR2_X1 U2834 ( .A1(n4177), .A2(n3232), .ZN(n2261) );
  AND2_X1 U2835 ( .A1(n3175), .A2(n3174), .ZN(n2262) );
  OR2_X1 U2836 ( .A1(n2821), .A2(n2712), .ZN(n3801) );
  INV_X2 U2837 ( .A(n3801), .ZN(U4043) );
  OR2_X1 U2838 ( .A1(n3362), .A2(n4341), .ZN(n2264) );
  OR2_X1 U2839 ( .A1(n3362), .A2(n4281), .ZN(n2265) );
  AND2_X1 U2840 ( .A1(n3979), .A2(n2663), .ZN(n3978) );
  AND2_X1 U2841 ( .A1(n3313), .A2(n3314), .ZN(n2266) );
  INV_X1 U2842 ( .A(n2636), .ZN(n3734) );
  OR2_X1 U2843 ( .A1(n3945), .A2(n3968), .ZN(n2267) );
  INV_X1 U2844 ( .A(IR_REG_13__SCAN_IN), .ZN(n2275) );
  INV_X1 U2845 ( .A(n3223), .ZN(n3224) );
  NAND2_X1 U2846 ( .A1(n3300), .A2(n2943), .ZN(n2944) );
  NAND2_X1 U2847 ( .A1(n3222), .A2(n3224), .ZN(n3225) );
  INV_X1 U2848 ( .A(IR_REG_25__SCAN_IN), .ZN(n2281) );
  INV_X1 U2849 ( .A(n3192), .ZN(n3193) );
  INV_X1 U2850 ( .A(IR_REG_24__SCAN_IN), .ZN(n2674) );
  NOR2_X1 U2851 ( .A1(n2060), .A2(n4460), .ZN(n2341) );
  INV_X1 U2852 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2450) );
  INV_X1 U2853 ( .A(IR_REG_21__SCAN_IN), .ZN(n2618) );
  INV_X1 U2854 ( .A(n3184), .ZN(n3185) );
  INV_X1 U2855 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4649) );
  INV_X1 U2856 ( .A(n2537), .ZN(n2536) );
  NAND2_X1 U2857 ( .A1(n2570), .A2(REG3_REG_25__SCAN_IN), .ZN(n2581) );
  OR2_X1 U2858 ( .A1(n2718), .A2(n2703), .ZN(n2682) );
  NAND2_X1 U2859 ( .A1(n2495), .A2(REG3_REG_18__SCAN_IN), .ZN(n2506) );
  AND2_X1 U2860 ( .A1(n3947), .A2(n3932), .ZN(n3716) );
  NAND2_X1 U2861 ( .A1(n2555), .A2(n2554), .ZN(n4000) );
  NAND2_X1 U2862 ( .A1(n2440), .A2(REG3_REG_13__SCAN_IN), .ZN(n2451) );
  OR2_X1 U2863 ( .A1(n2388), .A2(n2387), .ZN(n2403) );
  NAND2_X1 U2864 ( .A1(n2349), .A2(n2348), .ZN(n3003) );
  OR2_X1 U2865 ( .A1(n3805), .A2(n3535), .ZN(n2413) );
  AND2_X1 U2866 ( .A1(n3807), .A2(n3371), .ZN(n2399) );
  INV_X1 U2867 ( .A(n3786), .ZN(n2688) );
  INV_X1 U2868 ( .A(n3876), .ZN(n2894) );
  INV_X1 U2869 ( .A(n3947), .ZN(n3909) );
  INV_X1 U2870 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3512) );
  INV_X1 U2871 ( .A(n4001), .ZN(n4034) );
  OR2_X1 U2872 ( .A1(n2881), .A2(n2879), .ZN(n2856) );
  INV_X1 U2873 ( .A(n4000), .ZN(n4706) );
  NOR2_X1 U2874 ( .A1(n2059), .A2(n2929), .ZN(n2317) );
  INV_X1 U2875 ( .A(n4354), .ZN(n2852) );
  OR2_X1 U2876 ( .A1(n2410), .A2(IR_REG_9__SCAN_IN), .ZN(n2423) );
  INV_X1 U2877 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4556) );
  INV_X1 U2878 ( .A(n3698), .ZN(n3883) );
  NOR2_X1 U2879 ( .A1(n4149), .A2(n3626), .ZN(n2470) );
  MUX2_X1 U2880 ( .A(DATAI_1_), .B(n4353), .S(n2346), .Z(n2943) );
  INV_X1 U2881 ( .A(n4207), .ZN(n4198) );
  NOR2_X1 U2882 ( .A1(n3692), .A2(n2588), .ZN(n3926) );
  INV_X1 U2883 ( .A(n4172), .ZN(n4183) );
  AND2_X1 U2884 ( .A1(n3086), .A2(n3654), .ZN(n3724) );
  OR2_X1 U2885 ( .A1(n2852), .A2(n2847), .ZN(n4176) );
  INV_X1 U2886 ( .A(n4489), .ZN(n4482) );
  NAND2_X1 U2887 ( .A1(n2951), .A2(n2852), .ZN(n3566) );
  NOR2_X1 U2888 ( .A1(n3692), .A2(n2534), .ZN(n3446) );
  AND2_X1 U2889 ( .A1(n2571), .A2(n2561), .ZN(n3969) );
  AOI21_X1 U2890 ( .B1(n3177), .B2(n3176), .A(n2262), .ZN(n3520) );
  NAND2_X2 U2891 ( .A1(n2986), .A2(n2985), .ZN(n3631) );
  OR2_X1 U2892 ( .A1(n3468), .A2(n2058), .ZN(n2577) );
  AND2_X1 U2893 ( .A1(n2412), .A2(n2423), .ZN(n3131) );
  INV_X1 U2894 ( .A(n4444), .ZN(n4435) );
  AND2_X1 U2895 ( .A1(n2708), .A2(n4346), .ZN(n4207) );
  INV_X1 U2896 ( .A(n3978), .ZN(n3998) );
  AND2_X1 U2897 ( .A1(n4053), .A2(n4054), .ZN(n4072) );
  INV_X1 U2898 ( .A(n4132), .ZN(n4179) );
  AND2_X1 U2899 ( .A1(n3646), .A2(n3662), .ZN(n3723) );
  AND2_X1 U2900 ( .A1(n4082), .A2(n4496), .ZN(n4362) );
  INV_X1 U2901 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4536) );
  INV_X1 U2902 ( .A(n4499), .ZN(n4508) );
  AND2_X1 U2903 ( .A1(n4452), .A2(n2635), .ZN(n4489) );
  INV_X1 U2904 ( .A(n2858), .ZN(n2882) );
  NAND2_X1 U2905 ( .A1(n2684), .A2(n2687), .ZN(n2982) );
  AND2_X1 U2906 ( .A1(n2449), .A2(n2466), .ZN(n3841) );
  AND2_X1 U2907 ( .A1(n2748), .A2(n2735), .ZN(n4425) );
  NAND2_X1 U2908 ( .A1(n2860), .A2(n2859), .ZN(n3619) );
  INV_X1 U2909 ( .A(n3381), .ZN(n3911) );
  NAND2_X1 U2910 ( .A1(n2577), .A2(n2576), .ZN(n3964) );
  OR2_X1 U2911 ( .A1(n4369), .A2(n3792), .ZN(n4440) );
  OR2_X1 U2912 ( .A1(n4369), .A2(n4354), .ZN(n4438) );
  OR2_X1 U2913 ( .A1(n4369), .A2(n4367), .ZN(n4444) );
  INV_X1 U2914 ( .A(n3897), .ZN(n4141) );
  INV_X1 U2915 ( .A(n4362), .ZN(n4138) );
  NAND2_X1 U2916 ( .A1(n4519), .A2(n4496), .ZN(n4281) );
  AND2_X2 U2917 ( .A1(n2710), .A2(n2705), .ZN(n4519) );
  NAND2_X1 U2918 ( .A1(n4511), .A2(n4496), .ZN(n4341) );
  INV_X1 U2919 ( .A(n4511), .ZN(n4510) );
  INV_X1 U2920 ( .A(n4462), .ZN(n4463) );
  NAND2_X1 U2921 ( .A1(n2839), .A2(n2882), .ZN(n4462) );
  AND2_X1 U2922 ( .A1(n2982), .A2(STATE_REG_SCAN_IN), .ZN(n4464) );
  AND2_X1 U2923 ( .A1(n2481), .A2(n2469), .ZN(n4347) );
  AND2_X1 U2924 ( .A1(n2397), .A2(n2396), .ZN(n4349) );
  NOR2_X1 U2925 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2273)
         );
  NOR2_X1 U2926 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2272)
         );
  NOR2_X1 U2927 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2271)
         );
  NOR2_X1 U2928 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2270)
         );
  NOR2_X1 U2929 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2280)
         );
  NOR2_X1 U2930 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2279)
         );
  NOR2_X1 U2931 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2278)
         );
  NOR2_X1 U2932 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2277)
         );
  OR2_X2 U2933 ( .A1(n3355), .A2(n2480), .ZN(n2287) );
  INV_X4 U2934 ( .A(n2351), .ZN(n3704) );
  NAND2_X1 U2935 ( .A1(n3704), .A2(REG0_REG_10__SCAN_IN), .ZN(n2299) );
  INV_X1 U2936 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3106) );
  OR2_X1 U2937 ( .A1(n2060), .A2(n3106), .ZN(n2298) );
  NAND2_X1 U2938 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2362) );
  INV_X1 U2939 ( .A(n2362), .ZN(n2289) );
  NAND2_X1 U2940 ( .A1(n2289), .A2(REG3_REG_5__SCAN_IN), .ZN(n2375) );
  INV_X1 U2941 ( .A(n2375), .ZN(n2290) );
  NAND2_X1 U2942 ( .A1(n2290), .A2(REG3_REG_6__SCAN_IN), .ZN(n2388) );
  NAND2_X1 U2943 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2291) );
  INV_X1 U2944 ( .A(n2404), .ZN(n2292) );
  NAND2_X1 U2945 ( .A1(n2292), .A2(REG3_REG_10__SCAN_IN), .ZN(n2417) );
  INV_X1 U2946 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2293) );
  NAND2_X1 U2947 ( .A1(n2404), .A2(n2293), .ZN(n2294) );
  NAND2_X1 U2948 ( .A1(n2417), .A2(n2294), .ZN(n3410) );
  OR2_X1 U2949 ( .A1(n2058), .A2(n3410), .ZN(n2297) );
  OR2_X1 U2950 ( .A1(n2059), .A2(n4376), .ZN(n2296) );
  NAND4_X1 U2951 ( .A1(n2299), .A2(n2298), .A3(n2297), .A4(n2296), .ZN(n3804)
         );
  INV_X1 U2952 ( .A(n3804), .ZN(n3149) );
  NAND2_X1 U2953 ( .A1(n2300), .A2(n2301), .ZN(n2382) );
  NOR2_X1 U2954 ( .A1(n2382), .A2(IR_REG_6__SCAN_IN), .ZN(n2306) );
  NOR2_X1 U2955 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2302)
         );
  NAND2_X1 U2956 ( .A1(n2306), .A2(n2302), .ZN(n2410) );
  NAND2_X1 U2957 ( .A1(n2423), .A2(IR_REG_31__SCAN_IN), .ZN(n2303) );
  XNOR2_X1 U2958 ( .A(n2303), .B(IR_REG_10__SCAN_IN), .ZN(n4472) );
  NAND2_X1 U2959 ( .A1(n2258), .A2(n2480), .ZN(n2304) );
  MUX2_X1 U2960 ( .A(DATAI_10_), .B(n4472), .S(n3692), .Z(n3409) );
  INV_X1 U2961 ( .A(n3409), .ZN(n3220) );
  OR2_X1 U2962 ( .A1(n2306), .A2(n2480), .ZN(n2395) );
  NAND2_X1 U2963 ( .A1(n2395), .A2(n2394), .ZN(n2397) );
  NAND2_X1 U2964 ( .A1(n2397), .A2(IR_REG_31__SCAN_IN), .ZN(n2307) );
  XNOR2_X1 U2965 ( .A(n2307), .B(IR_REG_8__SCAN_IN), .ZN(n4348) );
  MUX2_X1 U2966 ( .A(DATAI_8_), .B(n4348), .S(n3692), .Z(n3431) );
  INV_X4 U2967 ( .A(n2338), .ZN(n2628) );
  NAND2_X1 U2968 ( .A1(n2628), .A2(REG2_REG_8__SCAN_IN), .ZN(n2313) );
  INV_X1 U2969 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2308) );
  OR2_X1 U2970 ( .A1(n2590), .A2(n2308), .ZN(n2312) );
  INV_X1 U2971 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2402) );
  XNOR2_X1 U2972 ( .A(n2403), .B(n2402), .ZN(n3432) );
  OR2_X1 U2973 ( .A1(n2058), .A2(n3432), .ZN(n2311) );
  INV_X1 U2974 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2309) );
  OR2_X1 U2975 ( .A1(n2059), .A2(n2309), .ZN(n2310) );
  NAND4_X1 U2976 ( .A1(n2313), .A2(n2312), .A3(n2311), .A4(n2310), .ZN(n3806)
         );
  INV_X1 U2977 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2929) );
  INV_X1 U2978 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2959) );
  OR2_X1 U2979 ( .A1(n2338), .A2(n2959), .ZN(n2315) );
  INV_X1 U2980 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2976) );
  OR2_X1 U2981 ( .A1(n2342), .A2(n2976), .ZN(n2314) );
  NAND2_X1 U2982 ( .A1(n3704), .A2(REG0_REG_2__SCAN_IN), .ZN(n2318) );
  INV_X1 U2983 ( .A(n3810), .ZN(n2905) );
  MUX2_X1 U2984 ( .A(DATAI_2_), .B(n4352), .S(n2346), .Z(n2965) );
  NAND2_X1 U2985 ( .A1(n2905), .A2(n2974), .ZN(n2901) );
  NAND2_X1 U2986 ( .A1(n3704), .A2(REG0_REG_3__SCAN_IN), .ZN(n2325) );
  INV_X1 U2987 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2321) );
  OR2_X1 U2988 ( .A1(n2609), .A2(n2321), .ZN(n2323) );
  INV_X1 U2989 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2745) );
  OR2_X1 U2990 ( .A1(n2060), .A2(n2745), .ZN(n2322) );
  NOR2_X1 U2991 ( .A1(n2326), .A2(n2480), .ZN(n2327) );
  NAND2_X1 U2992 ( .A1(n2327), .A2(IR_REG_3__SCAN_IN), .ZN(n2330) );
  INV_X1 U2993 ( .A(n2327), .ZN(n2329) );
  INV_X1 U2994 ( .A(IR_REG_3__SCAN_IN), .ZN(n2328) );
  NAND2_X1 U2995 ( .A1(n2329), .A2(n2328), .ZN(n2357) );
  MUX2_X1 U2996 ( .A(DATAI_3_), .B(n2755), .S(n3692), .Z(n2997) );
  NAND2_X1 U2997 ( .A1(n2975), .A2(n2910), .ZN(n2331) );
  AND2_X1 U2998 ( .A1(n2901), .A2(n2331), .ZN(n2347) );
  INV_X1 U2999 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2954) );
  INV_X1 U3000 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2332) );
  OR2_X1 U3001 ( .A1(n2332), .A2(n2288), .ZN(n2333) );
  NAND2_X1 U3002 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2334)
         );
  INV_X1 U3003 ( .A(n2943), .ZN(n2952) );
  INV_X1 U3004 ( .A(n2609), .ZN(n2337) );
  NAND2_X1 U3005 ( .A1(n2337), .A2(REG1_REG_0__SCAN_IN), .ZN(n2345) );
  INV_X1 U3006 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4460) );
  INV_X1 U3007 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2339) );
  NOR2_X1 U3008 ( .A1(n2351), .A2(n2339), .ZN(n2340) );
  NOR2_X1 U3009 ( .A1(n2341), .A2(n2340), .ZN(n2344) );
  INV_X1 U3010 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2864) );
  OR2_X1 U3011 ( .A1(n2058), .A2(n2864), .ZN(n2343) );
  MUX2_X1 U3012 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(n2346), .Z(n2855) );
  AND2_X1 U3013 ( .A1(n2825), .A2(n2855), .ZN(n2888) );
  NAND2_X1 U3014 ( .A1(n2905), .A2(n2965), .ZN(n2638) );
  NAND2_X1 U3015 ( .A1(n3810), .A2(n2974), .ZN(n3641) );
  NAND2_X1 U3016 ( .A1(n2638), .A2(n3641), .ZN(n2636) );
  NAND2_X1 U3017 ( .A1(n2917), .A2(n2636), .ZN(n2900) );
  NAND2_X1 U3018 ( .A1(n2347), .A2(n2900), .ZN(n2349) );
  NAND2_X1 U3019 ( .A1(n3524), .A2(n2997), .ZN(n2348) );
  NAND2_X1 U3020 ( .A1(n2628), .A2(REG2_REG_4__SCAN_IN), .ZN(n2356) );
  INV_X1 U3021 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2350) );
  OR2_X1 U3022 ( .A1(n2351), .A2(n2350), .ZN(n2355) );
  OAI21_X1 U3023 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2362), .ZN(n3525) );
  OR2_X1 U3024 ( .A1(n2058), .A2(n3525), .ZN(n2354) );
  INV_X1 U3025 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2352) );
  NAND2_X1 U3026 ( .A1(n2357), .A2(IR_REG_31__SCAN_IN), .ZN(n2358) );
  XNOR2_X1 U3027 ( .A(n2358), .B(IR_REG_4__SCAN_IN), .ZN(n4351) );
  MUX2_X1 U3028 ( .A(DATAI_4_), .B(n4351), .S(n3692), .Z(n3523) );
  INV_X1 U3029 ( .A(n3523), .ZN(n3181) );
  NAND2_X1 U3030 ( .A1(n3491), .A2(n3181), .ZN(n3647) );
  INV_X1 U3031 ( .A(n3735), .ZN(n2359) );
  NAND2_X1 U3032 ( .A1(n3003), .A2(n2359), .ZN(n3006) );
  NAND2_X1 U3033 ( .A1(n3491), .A2(n3523), .ZN(n2360) );
  NAND2_X1 U3034 ( .A1(n3006), .A2(n2360), .ZN(n3031) );
  NAND2_X1 U3035 ( .A1(n3704), .A2(REG0_REG_5__SCAN_IN), .ZN(n2367) );
  INV_X1 U3036 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3037) );
  OR2_X1 U3037 ( .A1(n2060), .A2(n3037), .ZN(n2366) );
  INV_X1 U3038 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2361) );
  NAND2_X1 U3039 ( .A1(n2362), .A2(n2361), .ZN(n2363) );
  NAND2_X1 U3040 ( .A1(n2375), .A2(n2363), .ZN(n3042) );
  OR2_X1 U3041 ( .A1(n2058), .A2(n3042), .ZN(n2365) );
  INV_X1 U3042 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2762) );
  OR2_X1 U3043 ( .A1(n2609), .A2(n2762), .ZN(n2364) );
  NAND4_X1 U3044 ( .A1(n2367), .A2(n2366), .A3(n2365), .A4(n2364), .ZN(n3809)
         );
  INV_X1 U3045 ( .A(n3809), .ZN(n3020) );
  NOR2_X1 U3046 ( .A1(n2300), .A2(n2480), .ZN(n2368) );
  MUX2_X1 U3047 ( .A(n2480), .B(n2368), .S(IR_REG_5__SCAN_IN), .Z(n2370) );
  INV_X1 U3048 ( .A(n2382), .ZN(n2369) );
  MUX2_X1 U3049 ( .A(DATAI_5_), .B(n4350), .S(n3692), .Z(n3490) );
  NAND2_X1 U3050 ( .A1(n3020), .A2(n3187), .ZN(n2372) );
  AND2_X1 U3051 ( .A1(n3809), .A2(n3490), .ZN(n2371) );
  AOI21_X2 U3052 ( .B1(n3031), .B2(n2372), .A(n2371), .ZN(n3021) );
  NAND2_X1 U3053 ( .A1(n2628), .A2(REG2_REG_6__SCAN_IN), .ZN(n2381) );
  INV_X1 U3054 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2373) );
  OR2_X1 U3055 ( .A1(n2590), .A2(n2373), .ZN(n2380) );
  INV_X1 U3056 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2374) );
  NAND2_X1 U3057 ( .A1(n2375), .A2(n2374), .ZN(n2376) );
  NAND2_X1 U3058 ( .A1(n2388), .A2(n2376), .ZN(n3025) );
  OR2_X1 U3059 ( .A1(n2058), .A2(n3025), .ZN(n2379) );
  INV_X1 U3060 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2377) );
  OR2_X1 U3061 ( .A1(n2609), .A2(n2377), .ZN(n2378) );
  NAND4_X1 U3062 ( .A1(n2381), .A2(n2380), .A3(n2379), .A4(n2378), .ZN(n3808)
         );
  NAND2_X1 U3063 ( .A1(n2382), .A2(IR_REG_31__SCAN_IN), .ZN(n2383) );
  XNOR2_X1 U3064 ( .A(n2383), .B(IR_REG_6__SCAN_IN), .ZN(n2777) );
  MUX2_X1 U3065 ( .A(DATAI_6_), .B(n2777), .S(n3692), .Z(n3603) );
  NAND2_X1 U3066 ( .A1(n3808), .A2(n3603), .ZN(n2385) );
  NOR2_X1 U3067 ( .A1(n3808), .A2(n3603), .ZN(n2384) );
  AOI21_X2 U3068 ( .B1(n3021), .B2(n2385), .A(n2384), .ZN(n3062) );
  NAND2_X1 U3069 ( .A1(n2628), .A2(REG2_REG_7__SCAN_IN), .ZN(n2393) );
  INV_X1 U3070 ( .A(REG0_REG_7__SCAN_IN), .ZN(n2386) );
  OR2_X1 U3071 ( .A1(n2590), .A2(n2386), .ZN(n2392) );
  NAND2_X1 U3072 ( .A1(n2388), .A2(n2387), .ZN(n2389) );
  NAND2_X1 U3073 ( .A1(n2403), .A2(n2389), .ZN(n3372) );
  OR2_X1 U3074 ( .A1(n2058), .A2(n3372), .ZN(n2391) );
  INV_X1 U3075 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2807) );
  OR2_X1 U3076 ( .A1(n2609), .A2(n2807), .ZN(n2390) );
  NAND4_X1 U3077 ( .A1(n2393), .A2(n2392), .A3(n2391), .A4(n2390), .ZN(n3807)
         );
  INV_X1 U3078 ( .A(n3807), .ZN(n2398) );
  OR2_X1 U3079 ( .A1(n2395), .A2(n2394), .ZN(n2396) );
  MUX2_X1 U3080 ( .A(DATAI_7_), .B(n4349), .S(n3692), .Z(n3371) );
  NAND2_X1 U3081 ( .A1(n2398), .A2(n3371), .ZN(n2643) );
  INV_X1 U3082 ( .A(n3371), .ZN(n3200) );
  NAND2_X1 U3083 ( .A1(n3807), .A2(n3200), .ZN(n3652) );
  NAND2_X1 U3084 ( .A1(n2643), .A2(n3652), .ZN(n3061) );
  INV_X1 U3085 ( .A(n3806), .ZN(n3089) );
  INV_X1 U3086 ( .A(n3431), .ZN(n3207) );
  NAND2_X1 U3087 ( .A1(n2628), .A2(REG2_REG_9__SCAN_IN), .ZN(n2409) );
  INV_X1 U3088 ( .A(REG0_REG_9__SCAN_IN), .ZN(n2400) );
  OR2_X1 U3089 ( .A1(n2590), .A2(n2400), .ZN(n2408) );
  INV_X1 U3090 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2401) );
  OAI21_X1 U3091 ( .B1(n2403), .B2(n2402), .A(n2401), .ZN(n2405) );
  NAND2_X1 U3092 ( .A1(n2405), .A2(n2404), .ZN(n3095) );
  OR2_X1 U3093 ( .A1(n2058), .A2(n3095), .ZN(n2407) );
  INV_X1 U3094 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2873) );
  OR2_X1 U3095 ( .A1(n2609), .A2(n2873), .ZN(n2406) );
  NAND4_X1 U3096 ( .A1(n2409), .A2(n2408), .A3(n2407), .A4(n2406), .ZN(n3805)
         );
  INV_X1 U3097 ( .A(n3805), .ZN(n3068) );
  NAND2_X1 U3098 ( .A1(n2410), .A2(IR_REG_31__SCAN_IN), .ZN(n2411) );
  MUX2_X1 U3099 ( .A(IR_REG_31__SCAN_IN), .B(n2411), .S(IR_REG_9__SCAN_IN), 
        .Z(n2412) );
  MUX2_X1 U3100 ( .A(DATAI_9_), .B(n3131), .S(n3692), .Z(n3535) );
  NAND2_X1 U3101 ( .A1(n3092), .A2(n2263), .ZN(n2414) );
  NAND2_X1 U3102 ( .A1(n2414), .A2(n2413), .ZN(n3103) );
  NAND2_X1 U3103 ( .A1(n3704), .A2(REG0_REG_11__SCAN_IN), .ZN(n2422) );
  INV_X1 U3104 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2415) );
  OR2_X1 U3105 ( .A1(n2060), .A2(n2415), .ZN(n2421) );
  INV_X1 U3106 ( .A(n2417), .ZN(n2416) );
  NAND2_X1 U3107 ( .A1(n2416), .A2(REG3_REG_11__SCAN_IN), .ZN(n2428) );
  INV_X1 U3108 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3577) );
  NAND2_X1 U3109 ( .A1(n2417), .A2(n3577), .ZN(n2418) );
  NAND2_X1 U3110 ( .A1(n2428), .A2(n2418), .ZN(n3154) );
  OR2_X1 U3111 ( .A1(n2058), .A2(n3154), .ZN(n2420) );
  INV_X1 U3112 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4279) );
  OR2_X1 U3113 ( .A1(n2059), .A2(n4279), .ZN(n2419) );
  NAND4_X1 U3114 ( .A1(n2422), .A2(n2421), .A3(n2420), .A4(n2419), .ZN(n3458)
         );
  INV_X1 U3115 ( .A(n3458), .ZN(n3227) );
  NAND2_X1 U3116 ( .A1(n2424), .A2(IR_REG_31__SCAN_IN), .ZN(n2435) );
  MUX2_X1 U3117 ( .A(DATAI_11_), .B(n4470), .S(n3692), .Z(n3578) );
  NAND2_X1 U3118 ( .A1(n3227), .A2(n3578), .ZN(n3158) );
  INV_X1 U3119 ( .A(n3578), .ZN(n3226) );
  NAND2_X1 U3120 ( .A1(n3458), .A2(n3226), .ZN(n3160) );
  NAND2_X1 U3121 ( .A1(n3158), .A2(n3160), .ZN(n3144) );
  INV_X1 U3122 ( .A(REG2_REG_12__SCAN_IN), .ZN(n2426) );
  OR2_X1 U3123 ( .A1(n2060), .A2(n2426), .ZN(n2433) );
  INV_X1 U3124 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4335) );
  OR2_X1 U3125 ( .A1(n2590), .A2(n4335), .ZN(n2432) );
  NAND2_X1 U3126 ( .A1(n2428), .A2(n2427), .ZN(n2429) );
  NAND2_X1 U3127 ( .A1(n2441), .A2(n2429), .ZN(n3168) );
  OR2_X1 U3128 ( .A1(n2058), .A2(n3168), .ZN(n2431) );
  OR2_X1 U3129 ( .A1(n2609), .A2(n4536), .ZN(n2430) );
  NAND4_X1 U3130 ( .A1(n2433), .A2(n2432), .A3(n2431), .A4(n2430), .ZN(n3580)
         );
  INV_X1 U3131 ( .A(n3580), .ZN(n4177) );
  INV_X1 U3132 ( .A(IR_REG_11__SCAN_IN), .ZN(n2434) );
  NAND2_X1 U3133 ( .A1(n2435), .A2(n2434), .ZN(n2436) );
  NAND2_X1 U3134 ( .A1(n2436), .A2(IR_REG_31__SCAN_IN), .ZN(n2437) );
  XNOR2_X1 U3135 ( .A(n2437), .B(IR_REG_12__SCAN_IN), .ZN(n3134) );
  MUX2_X1 U3136 ( .A(DATAI_12_), .B(n3134), .S(n3692), .Z(n3457) );
  NAND2_X1 U3137 ( .A1(n3165), .A2(n2261), .ZN(n2439) );
  NAND2_X1 U3138 ( .A1(n2439), .A2(n2438), .ZN(n4165) );
  NAND2_X1 U3139 ( .A1(n3704), .A2(REG0_REG_13__SCAN_IN), .ZN(n2446) );
  INV_X1 U3140 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4189) );
  OR2_X1 U3141 ( .A1(n2060), .A2(n4189), .ZN(n2445) );
  INV_X1 U3142 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3129) );
  NAND2_X1 U3143 ( .A1(n2441), .A2(n3129), .ZN(n2442) );
  NAND2_X1 U3144 ( .A1(n2451), .A2(n2442), .ZN(n4188) );
  OR2_X1 U3145 ( .A1(n2058), .A2(n4188), .ZN(n2444) );
  INV_X1 U3146 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4271) );
  OR2_X1 U3147 ( .A1(n2059), .A2(n4271), .ZN(n2443) );
  NAND4_X1 U31480 ( .A1(n2446), .A2(n2445), .A3(n2444), .A4(n2443), .ZN(n3803)
         );
  INV_X1 U31490 ( .A(n3803), .ZN(n4151) );
  NAND2_X1 U3150 ( .A1(n2447), .A2(IR_REG_31__SCAN_IN), .ZN(n2448) );
  MUX2_X1 U3151 ( .A(IR_REG_31__SCAN_IN), .B(n2448), .S(IR_REG_13__SCAN_IN), 
        .Z(n2449) );
  OR2_X1 U3152 ( .A1(n2447), .A2(IR_REG_13__SCAN_IN), .ZN(n2466) );
  MUX2_X1 U3153 ( .A(DATAI_13_), .B(n3841), .S(n3692), .Z(n4172) );
  NAND2_X1 U3154 ( .A1(n3704), .A2(REG0_REG_14__SCAN_IN), .ZN(n2456) );
  INV_X1 U3155 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4159) );
  OR2_X1 U3156 ( .A1(n2060), .A2(n4159), .ZN(n2455) );
  NAND2_X1 U3157 ( .A1(n2451), .A2(n2450), .ZN(n2452) );
  NAND2_X1 U3158 ( .A1(n2460), .A2(n2452), .ZN(n4158) );
  OR2_X1 U3159 ( .A1(n2058), .A2(n4158), .ZN(n2454) );
  INV_X1 U3160 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4405) );
  OR2_X1 U3161 ( .A1(n2609), .A2(n4405), .ZN(n2453) );
  NAND4_X1 U3162 ( .A1(n2456), .A2(n2455), .A3(n2454), .A4(n2453), .ZN(n4174)
         );
  INV_X1 U3163 ( .A(n4174), .ZN(n2458) );
  NAND2_X1 U3164 ( .A1(n2466), .A2(IR_REG_31__SCAN_IN), .ZN(n2457) );
  XNOR2_X1 U3165 ( .A(n2457), .B(IR_REG_14__SCAN_IN), .ZN(n4410) );
  MUX2_X1 U3166 ( .A(DATAI_14_), .B(n4410), .S(n3692), .Z(n4155) );
  NAND2_X1 U3167 ( .A1(n2458), .A2(n4155), .ZN(n4124) );
  INV_X1 U3168 ( .A(n4155), .ZN(n2459) );
  NAND2_X1 U3169 ( .A1(n4174), .A2(n2459), .ZN(n3658) );
  NAND2_X1 U3170 ( .A1(n4124), .A2(n3658), .ZN(n4144) );
  NAND2_X1 U3171 ( .A1(n2628), .A2(REG2_REG_15__SCAN_IN), .ZN(n2465) );
  INV_X1 U3172 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4323) );
  OR2_X1 U3173 ( .A1(n2590), .A2(n4323), .ZN(n2464) );
  NAND2_X1 U3174 ( .A1(n2460), .A2(n3625), .ZN(n2461) );
  NAND2_X1 U3175 ( .A1(n2474), .A2(n2461), .ZN(n3630) );
  OR2_X1 U3176 ( .A1(n2058), .A2(n3630), .ZN(n2463) );
  INV_X1 U3177 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4263) );
  OR2_X1 U3178 ( .A1(n2059), .A2(n4263), .ZN(n2462) );
  NAND4_X1 U3179 ( .A1(n2465), .A2(n2464), .A3(n2463), .A4(n2462), .ZN(n4149)
         );
  OAI21_X1 U3180 ( .B1(n2466), .B2(IR_REG_14__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2468) );
  NAND2_X1 U3181 ( .A1(n2468), .A2(n2467), .ZN(n2481) );
  OR2_X1 U3182 ( .A1(n2468), .A2(n2467), .ZN(n2469) );
  MUX2_X1 U3183 ( .A(DATAI_15_), .B(n4347), .S(n3692), .Z(n3626) );
  NAND2_X1 U3184 ( .A1(n4149), .A2(n3626), .ZN(n2471) );
  INV_X1 U3185 ( .A(n4149), .ZN(n2654) );
  NAND2_X1 U3186 ( .A1(n3704), .A2(REG0_REG_16__SCAN_IN), .ZN(n2479) );
  INV_X1 U3187 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4116) );
  OR2_X1 U3188 ( .A1(n2060), .A2(n4116), .ZN(n2478) );
  INV_X1 U3189 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2473) );
  NAND2_X1 U3190 ( .A1(n2474), .A2(n2473), .ZN(n2475) );
  NAND2_X1 U3191 ( .A1(n2486), .A2(n2475), .ZN(n4115) );
  OR2_X1 U3192 ( .A1(n2058), .A2(n4115), .ZN(n2477) );
  INV_X1 U3193 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4416) );
  OR2_X1 U3194 ( .A1(n2609), .A2(n4416), .ZN(n2476) );
  NAND4_X1 U3195 ( .A1(n2479), .A2(n2478), .A3(n2477), .A4(n2476), .ZN(n4095)
         );
  INV_X1 U3196 ( .A(n4095), .ZN(n4128) );
  NAND2_X1 U3197 ( .A1(n2481), .A2(IR_REG_31__SCAN_IN), .ZN(n2483) );
  XNOR2_X1 U3198 ( .A(n2483), .B(n2482), .ZN(n4468) );
  INV_X1 U3199 ( .A(n4468), .ZN(n2484) );
  MUX2_X1 U3200 ( .A(DATAI_16_), .B(n2484), .S(n3692), .Z(n3480) );
  NAND2_X1 U3201 ( .A1(n4128), .A2(n3480), .ZN(n3759) );
  NAND2_X1 U3202 ( .A1(n4095), .A2(n4118), .ZN(n3679) );
  NAND2_X1 U3203 ( .A1(n3759), .A2(n3679), .ZN(n4108) );
  NAND2_X1 U3204 ( .A1(n4107), .A2(n4108), .ZN(n4106) );
  NAND2_X1 U3205 ( .A1(n4095), .A2(n3480), .ZN(n2485) );
  NAND2_X1 U3206 ( .A1(n2486), .A2(n4556), .ZN(n2487) );
  NAND2_X1 U3207 ( .A1(n2497), .A2(n2487), .ZN(n3503) );
  OR2_X1 U3208 ( .A1(n3503), .A2(n2058), .ZN(n2492) );
  INV_X1 U3209 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2488) );
  OR2_X1 U32100 ( .A1(n2060), .A2(n2488), .ZN(n2491) );
  INV_X1 U32110 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4318) );
  OR2_X1 U32120 ( .A1(n2590), .A2(n4318), .ZN(n2490) );
  INV_X1 U32130 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4254) );
  OR2_X1 U32140 ( .A1(n2609), .A2(n4254), .ZN(n2489) );
  NAND4_X1 U32150 ( .A1(n2492), .A2(n2491), .A3(n2490), .A4(n2489), .ZN(n4110)
         );
  NAND2_X1 U32160 ( .A1(n2503), .A2(IR_REG_31__SCAN_IN), .ZN(n2493) );
  XNOR2_X1 U32170 ( .A(n2493), .B(IR_REG_17__SCAN_IN), .ZN(n3870) );
  MUX2_X1 U32180 ( .A(DATAI_17_), .B(n3870), .S(n3692), .Z(n4098) );
  INV_X1 U32190 ( .A(n4110), .ZN(n4076) );
  INV_X1 U32200 ( .A(n4098), .ZN(n4092) );
  INV_X1 U32210 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2496) );
  NAND2_X1 U32220 ( .A1(n2497), .A2(n2496), .ZN(n2498) );
  NAND2_X1 U32230 ( .A1(n2506), .A2(n2498), .ZN(n3592) );
  OR2_X1 U32240 ( .A1(n3592), .A2(n2058), .ZN(n2502) );
  NAND2_X1 U32250 ( .A1(n2628), .A2(REG2_REG_18__SCAN_IN), .ZN(n2501) );
  NAND2_X1 U32260 ( .A1(n3704), .A2(REG0_REG_18__SCAN_IN), .ZN(n2500) );
  NAND2_X1 U32270 ( .A1(n2337), .A2(REG1_REG_18__SCAN_IN), .ZN(n2499) );
  NAND4_X1 U32280 ( .A1(n2502), .A2(n2501), .A3(n2500), .A4(n2499), .ZN(n3802)
         );
  INV_X1 U32290 ( .A(n2511), .ZN(n2504) );
  NAND2_X1 U32300 ( .A1(n2504), .A2(IR_REG_31__SCAN_IN), .ZN(n2505) );
  XNOR2_X1 U32310 ( .A(n2505), .B(IR_REG_18__SCAN_IN), .ZN(n4447) );
  MUX2_X1 U32320 ( .A(DATAI_18_), .B(n4447), .S(n3692), .Z(n4079) );
  NAND2_X1 U32330 ( .A1(n4093), .A2(n4079), .ZN(n4053) );
  INV_X1 U32340 ( .A(n4079), .ZN(n3272) );
  NAND2_X1 U32350 ( .A1(n3802), .A2(n3272), .ZN(n4054) );
  INV_X1 U32360 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4247) );
  AOI22_X1 U32370 ( .A1(n2628), .A2(REG2_REG_19__SCAN_IN), .B1(n3704), .B2(
        REG0_REG_19__SCAN_IN), .ZN(n2509) );
  NAND2_X1 U32380 ( .A1(n2506), .A2(n4649), .ZN(n2507) );
  NAND2_X1 U32390 ( .A1(n2527), .A2(n2507), .ZN(n3421) );
  OR2_X1 U32400 ( .A1(n3421), .A2(n2058), .ZN(n2508) );
  OAI211_X1 U32410 ( .C1(n2059), .C2(n4247), .A(n2509), .B(n2508), .ZN(n4074)
         );
  MUX2_X1 U32420 ( .A(DATAI_19_), .B(n2894), .S(n3692), .Z(n3420) );
  NAND2_X1 U32430 ( .A1(n2099), .A2(n3420), .ZN(n2515) );
  NAND2_X1 U32440 ( .A1(n4049), .A2(n2515), .ZN(n2517) );
  INV_X1 U32450 ( .A(n2099), .ZN(n3547) );
  NAND2_X1 U32460 ( .A1(n3547), .A2(n4064), .ZN(n2516) );
  NAND2_X1 U32470 ( .A1(n2517), .A2(n2516), .ZN(n4027) );
  XNOR2_X1 U32480 ( .A(n2527), .B(REG3_REG_20__SCAN_IN), .ZN(n4041) );
  NAND2_X1 U32490 ( .A1(n4041), .A2(n2589), .ZN(n2522) );
  INV_X1 U32500 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4243) );
  NAND2_X1 U32510 ( .A1(n2628), .A2(REG2_REG_20__SCAN_IN), .ZN(n2519) );
  NAND2_X1 U32520 ( .A1(n3704), .A2(REG0_REG_20__SCAN_IN), .ZN(n2518) );
  OAI211_X1 U32530 ( .C1(n4243), .C2(n2059), .A(n2519), .B(n2518), .ZN(n2520)
         );
  INV_X1 U32540 ( .A(n2520), .ZN(n2521) );
  INV_X1 U32550 ( .A(DATAI_20_), .ZN(n2523) );
  NAND2_X1 U32560 ( .A1(n4059), .A2(n4032), .ZN(n3747) );
  NAND2_X1 U32570 ( .A1(n4027), .A2(n3747), .ZN(n2524) );
  OR2_X1 U32580 ( .A1(n4059), .A2(n4032), .ZN(n3748) );
  NAND2_X1 U32590 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n2525) );
  INV_X1 U32600 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3546) );
  INV_X1 U32610 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2526) );
  OAI21_X1 U32620 ( .B1(n2527), .B2(n3546), .A(n2526), .ZN(n2528) );
  AND2_X1 U32630 ( .A1(n2537), .A2(n2528), .ZN(n4020) );
  NAND2_X1 U32640 ( .A1(n4020), .A2(n2589), .ZN(n2533) );
  INV_X1 U32650 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4672) );
  NAND2_X1 U32660 ( .A1(n2628), .A2(REG2_REG_21__SCAN_IN), .ZN(n2530) );
  NAND2_X1 U32670 ( .A1(n3704), .A2(REG0_REG_21__SCAN_IN), .ZN(n2529) );
  OAI211_X1 U32680 ( .C1(n4672), .C2(n2059), .A(n2530), .B(n2529), .ZN(n2531)
         );
  INV_X1 U32690 ( .A(n2531), .ZN(n2532) );
  INV_X1 U32700 ( .A(DATAI_21_), .ZN(n2534) );
  NAND2_X1 U32710 ( .A1(n4001), .A2(n3446), .ZN(n2535) );
  INV_X1 U32720 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4523) );
  NAND2_X1 U32730 ( .A1(n2537), .A2(n4523), .ZN(n2538) );
  AND2_X1 U32740 ( .A1(n2549), .A2(n2538), .ZN(n4006) );
  NAND2_X1 U32750 ( .A1(n4006), .A2(n2589), .ZN(n2544) );
  INV_X1 U32760 ( .A(REG1_REG_22__SCAN_IN), .ZN(n2541) );
  NAND2_X1 U32770 ( .A1(n2628), .A2(REG2_REG_22__SCAN_IN), .ZN(n2540) );
  NAND2_X1 U32780 ( .A1(n3704), .A2(REG0_REG_22__SCAN_IN), .ZN(n2539) );
  OAI211_X1 U32790 ( .C1(n2541), .C2(n2609), .A(n2540), .B(n2539), .ZN(n2542)
         );
  INV_X1 U32800 ( .A(n2542), .ZN(n2543) );
  INV_X1 U32810 ( .A(DATAI_22_), .ZN(n2545) );
  INV_X1 U32820 ( .A(n4007), .ZN(n3564) );
  NAND2_X1 U32830 ( .A1(n3800), .A2(n3564), .ZN(n2663) );
  NAND2_X1 U32840 ( .A1(n3800), .A2(n4007), .ZN(n2546) );
  NAND2_X1 U32850 ( .A1(n3996), .A2(n2546), .ZN(n3974) );
  INV_X1 U32860 ( .A(n2549), .ZN(n2547) );
  INV_X1 U32870 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2548) );
  NAND2_X1 U32880 ( .A1(n2549), .A2(n2548), .ZN(n2550) );
  NAND2_X1 U32890 ( .A1(n2560), .A2(n2550), .ZN(n3401) );
  OR2_X1 U32900 ( .A1(n3401), .A2(n2058), .ZN(n2555) );
  INV_X1 U32910 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4662) );
  NAND2_X1 U32920 ( .A1(n2628), .A2(REG2_REG_23__SCAN_IN), .ZN(n2552) );
  NAND2_X1 U32930 ( .A1(n3704), .A2(REG0_REG_23__SCAN_IN), .ZN(n2551) );
  OAI211_X1 U32940 ( .C1(n4662), .C2(n2609), .A(n2552), .B(n2551), .ZN(n2553)
         );
  INV_X1 U32950 ( .A(n2553), .ZN(n2554) );
  INV_X1 U32960 ( .A(DATAI_23_), .ZN(n2556) );
  INV_X1 U32970 ( .A(n3988), .ZN(n3983) );
  NAND2_X1 U32980 ( .A1(n4706), .A2(n3983), .ZN(n2557) );
  NAND2_X1 U32990 ( .A1(n3974), .A2(n2557), .ZN(n2559) );
  NAND2_X1 U33000 ( .A1(n4000), .A2(n3988), .ZN(n2558) );
  NAND2_X1 U33010 ( .A1(n2559), .A2(n2558), .ZN(n3958) );
  INV_X1 U33020 ( .A(n3958), .ZN(n2567) );
  NAND2_X1 U33030 ( .A1(n2560), .A2(n3512), .ZN(n2561) );
  NAND2_X1 U33040 ( .A1(n3969), .A2(n2589), .ZN(n2566) );
  INV_X1 U33050 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4228) );
  NAND2_X1 U33060 ( .A1(n2628), .A2(REG2_REG_24__SCAN_IN), .ZN(n2563) );
  NAND2_X1 U33070 ( .A1(n3704), .A2(REG0_REG_24__SCAN_IN), .ZN(n2562) );
  OAI211_X1 U33080 ( .C1(n4228), .C2(n2059), .A(n2563), .B(n2562), .ZN(n2564)
         );
  INV_X1 U33090 ( .A(n2564), .ZN(n2565) );
  INV_X1 U33100 ( .A(n3692), .ZN(n3708) );
  NAND2_X1 U33110 ( .A1(n2567), .A2(n2267), .ZN(n2569) );
  NAND2_X1 U33120 ( .A1(n3945), .A2(n3968), .ZN(n2568) );
  NAND2_X1 U33130 ( .A1(n2569), .A2(n2568), .ZN(n3939) );
  INV_X1 U33140 ( .A(n2571), .ZN(n2570) );
  INV_X1 U33150 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3469) );
  NAND2_X1 U33160 ( .A1(n2571), .A2(n3469), .ZN(n2572) );
  NAND2_X1 U33170 ( .A1(n2581), .A2(n2572), .ZN(n3468) );
  INV_X1 U33180 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4671) );
  NAND2_X1 U33190 ( .A1(n2628), .A2(REG2_REG_25__SCAN_IN), .ZN(n2574) );
  NAND2_X1 U33200 ( .A1(n3704), .A2(REG0_REG_25__SCAN_IN), .ZN(n2573) );
  OAI211_X1 U33210 ( .C1(n4671), .C2(n2059), .A(n2574), .B(n2573), .ZN(n2575)
         );
  INV_X1 U33220 ( .A(n2575), .ZN(n2576) );
  INV_X1 U33230 ( .A(DATAI_25_), .ZN(n2578) );
  NOR2_X1 U33240 ( .A1(n3964), .A2(n3950), .ZN(n2580) );
  NAND2_X1 U33250 ( .A1(n3964), .A2(n3950), .ZN(n2579) );
  INV_X1 U33260 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3612) );
  NAND2_X1 U33270 ( .A1(n2581), .A2(n3612), .ZN(n2582) );
  NAND2_X1 U33280 ( .A1(n3934), .A2(n2589), .ZN(n2587) );
  INV_X1 U33290 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4680) );
  NAND2_X1 U33300 ( .A1(n2628), .A2(REG2_REG_26__SCAN_IN), .ZN(n2584) );
  NAND2_X1 U33310 ( .A1(n2337), .A2(REG1_REG_26__SCAN_IN), .ZN(n2583) );
  OAI211_X1 U33320 ( .C1(n2590), .C2(n4680), .A(n2584), .B(n2583), .ZN(n2585)
         );
  INV_X1 U33330 ( .A(n2585), .ZN(n2586) );
  INV_X1 U33340 ( .A(DATAI_26_), .ZN(n2588) );
  NOR2_X1 U33350 ( .A1(n3909), .A2(n3932), .ZN(n3902) );
  XNOR2_X1 U33360 ( .A(n2603), .B(REG3_REG_27__SCAN_IN), .ZN(n3916) );
  NAND2_X1 U33370 ( .A1(n3916), .A2(n2589), .ZN(n2596) );
  INV_X1 U33380 ( .A(REG1_REG_27__SCAN_IN), .ZN(n2593) );
  NAND2_X1 U33390 ( .A1(n2628), .A2(REG2_REG_27__SCAN_IN), .ZN(n2592) );
  INV_X1 U33400 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4544) );
  OR2_X1 U33410 ( .A1(n2590), .A2(n4544), .ZN(n2591) );
  OAI211_X1 U33420 ( .C1(n2593), .C2(n2609), .A(n2592), .B(n2591), .ZN(n2594)
         );
  INV_X1 U33430 ( .A(n2594), .ZN(n2595) );
  INV_X1 U33440 ( .A(DATAI_27_), .ZN(n2597) );
  AND2_X1 U33450 ( .A1(n3927), .A2(n3915), .ZN(n2601) );
  OR2_X1 U33460 ( .A1(n3902), .A2(n2601), .ZN(n2598) );
  OR2_X1 U33470 ( .A1(n3927), .A2(n3915), .ZN(n2599) );
  NAND2_X1 U33480 ( .A1(n3909), .A2(n3932), .ZN(n3903) );
  AND2_X1 U33490 ( .A1(n2599), .A2(n3903), .ZN(n2600) );
  INV_X1 U33500 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3380) );
  INV_X1 U33510 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2602) );
  OAI21_X1 U33520 ( .B1(n2603), .B2(n3380), .A(n2602), .ZN(n2606) );
  INV_X1 U3353 ( .A(n2603), .ZN(n2605) );
  AND2_X1 U33540 ( .A1(REG3_REG_28__SCAN_IN), .A2(REG3_REG_27__SCAN_IN), .ZN(
        n2604) );
  NAND2_X1 U3355 ( .A1(n2605), .A2(n2604), .ZN(n3881) );
  NAND2_X1 U3356 ( .A1(n2606), .A2(n3881), .ZN(n3349) );
  OR2_X1 U3357 ( .A1(n3349), .A2(n2058), .ZN(n2613) );
  INV_X1 U3358 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2610) );
  NAND2_X1 U3359 ( .A1(n2628), .A2(REG2_REG_28__SCAN_IN), .ZN(n2608) );
  NAND2_X1 U3360 ( .A1(n3704), .A2(REG0_REG_28__SCAN_IN), .ZN(n2607) );
  OAI211_X1 U3361 ( .C1(n2610), .C2(n2609), .A(n2608), .B(n2607), .ZN(n2611)
         );
  INV_X1 U3362 ( .A(n2611), .ZN(n2612) );
  NAND2_X1 U3363 ( .A1(n3708), .A2(DATAI_28_), .ZN(n3341) );
  INV_X1 U3364 ( .A(n3341), .ZN(n3892) );
  AND2_X1 U3365 ( .A1(n3381), .A2(n3892), .ZN(n3698) );
  NAND2_X1 U3366 ( .A1(n3911), .A2(n3341), .ZN(n3882) );
  NAND2_X1 U3367 ( .A1(n3883), .A2(n3882), .ZN(n3893) );
  NAND2_X1 U3368 ( .A1(n2615), .A2(n2614), .ZN(n2617) );
  NAND2_X1 U3369 ( .A1(n2617), .A2(IR_REG_31__SCAN_IN), .ZN(n2616) );
  MUX2_X1 U3370 ( .A(IR_REG_31__SCAN_IN), .B(n2616), .S(IR_REG_21__SCAN_IN), 
        .Z(n2620) );
  XNOR2_X1 U3371 ( .A(n2895), .B(n2635), .ZN(n2626) );
  AND2_X1 U3372 ( .A1(n2707), .A2(n2894), .ZN(n4452) );
  NAND2_X1 U3373 ( .A1(n2071), .A2(IR_REG_31__SCAN_IN), .ZN(n2627) );
  NAND2_X1 U3374 ( .A1(n3794), .A2(n3786), .ZN(n2847) );
  OR2_X1 U3375 ( .A1(n3881), .A2(n2058), .ZN(n2634) );
  INV_X1 U3376 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2631) );
  NAND2_X1 U3377 ( .A1(n2628), .A2(REG2_REG_29__SCAN_IN), .ZN(n2630) );
  NAND2_X1 U3378 ( .A1(n3704), .A2(REG0_REG_29__SCAN_IN), .ZN(n2629) );
  OAI211_X1 U3379 ( .C1(n2631), .C2(n2059), .A(n2630), .B(n2629), .ZN(n2632)
         );
  INV_X1 U3380 ( .A(n2632), .ZN(n2633) );
  INV_X1 U3381 ( .A(n2707), .ZN(n4346) );
  OAI22_X1 U3382 ( .A1(n3710), .A2(n4127), .B1(n3341), .B2(n4198), .ZN(n2667)
         );
  INV_X1 U3383 ( .A(n2825), .ZN(n2953) );
  NAND2_X1 U3384 ( .A1(n2953), .A2(n2855), .ZN(n2889) );
  NAND2_X1 U3385 ( .A1(n2919), .A2(n3638), .ZN(n2637) );
  NAND2_X1 U3386 ( .A1(n2637), .A2(n3734), .ZN(n2921) );
  NAND2_X1 U3387 ( .A1(n2921), .A2(n2638), .ZN(n2904) );
  NAND2_X1 U3388 ( .A1(n2975), .A2(n2997), .ZN(n3643) );
  NAND2_X1 U3389 ( .A1(n3524), .A2(n2910), .ZN(n3640) );
  INV_X1 U3390 ( .A(n3644), .ZN(n2639) );
  AND2_X1 U3391 ( .A1(n3809), .A2(n3187), .ZN(n3030) );
  NAND2_X1 U3392 ( .A1(n3020), .A2(n3490), .ZN(n3662) );
  OAI21_X1 U3393 ( .B1(n3032), .B2(n3030), .A(n3662), .ZN(n3016) );
  INV_X1 U3394 ( .A(n3603), .ZN(n2640) );
  NAND2_X1 U3395 ( .A1(n3808), .A2(n2640), .ZN(n3660) );
  NAND2_X1 U3396 ( .A1(n3016), .A2(n3660), .ZN(n2642) );
  INV_X1 U3397 ( .A(n3808), .ZN(n2641) );
  NAND2_X1 U3398 ( .A1(n2641), .A2(n3603), .ZN(n3649) );
  NAND2_X1 U3399 ( .A1(n2642), .A2(n3649), .ZN(n3053) );
  INV_X1 U3400 ( .A(n2643), .ZN(n2644) );
  OR2_X1 U3401 ( .A1(n3053), .A2(n2644), .ZN(n2645) );
  NAND2_X1 U3402 ( .A1(n2645), .A2(n3652), .ZN(n3067) );
  NAND2_X1 U3403 ( .A1(n3089), .A2(n3431), .ZN(n3653) );
  NAND2_X1 U3404 ( .A1(n3806), .A2(n3207), .ZN(n3651) );
  AND2_X1 U3405 ( .A1(n3805), .A2(n3093), .ZN(n3670) );
  NAND2_X1 U3406 ( .A1(n3068), .A2(n3535), .ZN(n3654) );
  NAND2_X1 U3407 ( .A1(n3804), .A2(n3220), .ZN(n3673) );
  NAND2_X1 U3408 ( .A1(n3099), .A2(n3673), .ZN(n2646) );
  NAND2_X1 U3409 ( .A1(n3149), .A2(n3409), .ZN(n3671) );
  NAND2_X1 U3410 ( .A1(n2646), .A2(n3671), .ZN(n3161) );
  NAND2_X1 U3411 ( .A1(n3580), .A2(n3232), .ZN(n4166) );
  NAND2_X1 U3412 ( .A1(n3803), .A2(n4183), .ZN(n2647) );
  NAND2_X1 U3413 ( .A1(n4166), .A2(n2647), .ZN(n2649) );
  INV_X1 U3414 ( .A(n3160), .ZN(n2648) );
  NOR2_X1 U3415 ( .A1(n2649), .A2(n2648), .ZN(n3674) );
  NAND2_X1 U3416 ( .A1(n3161), .A2(n3674), .ZN(n2653) );
  NAND2_X1 U3417 ( .A1(n4177), .A2(n3457), .ZN(n4168) );
  NAND2_X1 U3418 ( .A1(n3158), .A2(n4168), .ZN(n2652) );
  INV_X1 U3419 ( .A(n2649), .ZN(n2651) );
  NOR2_X1 U3420 ( .A1(n3803), .A2(n4183), .ZN(n2650) );
  AOI21_X1 U3421 ( .B1(n2652), .B2(n2651), .A(n2650), .ZN(n3676) );
  NAND2_X1 U3422 ( .A1(n2653), .A2(n3676), .ZN(n4147) );
  INV_X1 U3423 ( .A(n4144), .ZN(n4148) );
  NAND2_X1 U3424 ( .A1(n4147), .A2(n4148), .ZN(n4146) );
  NAND2_X1 U3425 ( .A1(n2654), .A2(n3626), .ZN(n3677) );
  NAND2_X1 U3426 ( .A1(n4149), .A2(n2100), .ZN(n3659) );
  NAND2_X1 U3427 ( .A1(n3677), .A2(n3659), .ZN(n4125) );
  INV_X1 U3428 ( .A(n4124), .ZN(n2655) );
  NOR2_X1 U3429 ( .A1(n4125), .A2(n2655), .ZN(n2656) );
  NAND2_X1 U3430 ( .A1(n4146), .A2(n2656), .ZN(n2657) );
  INV_X1 U3431 ( .A(n4108), .ZN(n3728) );
  NAND2_X1 U3432 ( .A1(n4074), .A2(n4064), .ZN(n2658) );
  AND2_X1 U3433 ( .A1(n2658), .A2(n4054), .ZN(n2661) );
  NAND2_X1 U3434 ( .A1(n4110), .A2(n4092), .ZN(n4050) );
  NAND2_X1 U3435 ( .A1(n2661), .A2(n4050), .ZN(n3757) );
  NAND2_X1 U3436 ( .A1(n4076), .A2(n4098), .ZN(n4051) );
  NAND2_X1 U3437 ( .A1(n4053), .A2(n4051), .ZN(n2660) );
  NOR2_X1 U3438 ( .A1(n4074), .A2(n4064), .ZN(n2659) );
  AOI21_X1 U3439 ( .B1(n2661), .B2(n2660), .A(n2659), .ZN(n4028) );
  OR2_X1 U3440 ( .A1(n4059), .A2(n4040), .ZN(n2662) );
  AND2_X1 U3441 ( .A1(n4028), .A2(n2662), .ZN(n3763) );
  AND2_X1 U3442 ( .A1(n4059), .A2(n4040), .ZN(n3761) );
  AOI21_X1 U3443 ( .B1(n4029), .B2(n3763), .A(n3761), .ZN(n4014) );
  NAND2_X1 U3444 ( .A1(n4034), .A2(n3446), .ZN(n3975) );
  NAND2_X1 U3445 ( .A1(n3979), .A2(n3975), .ZN(n3766) );
  AND2_X1 U3446 ( .A1(n4001), .A2(n4019), .ZN(n3720) );
  OAI21_X1 U3447 ( .B1(n4706), .B2(n3988), .A(n2663), .ZN(n3687) );
  AOI21_X1 U3448 ( .B1(n3720), .B2(n3979), .A(n3687), .ZN(n3764) );
  OAI21_X1 U3449 ( .B1(n4014), .B2(n3766), .A(n3764), .ZN(n3960) );
  INV_X1 U3450 ( .A(n3968), .ZN(n2664) );
  NAND2_X1 U3451 ( .A1(n3945), .A2(n2664), .ZN(n3746) );
  NAND2_X1 U3452 ( .A1(n4706), .A2(n3988), .ZN(n3959) );
  AND2_X1 U3453 ( .A1(n3746), .A2(n3959), .ZN(n3768) );
  NAND2_X1 U3454 ( .A1(n3960), .A2(n3768), .ZN(n3941) );
  INV_X1 U3455 ( .A(n3950), .ZN(n3944) );
  NAND2_X1 U3456 ( .A1(n3964), .A2(n3944), .ZN(n3719) );
  NAND2_X1 U3457 ( .A1(n3985), .A2(n3968), .ZN(n3940) );
  AND2_X1 U34580 ( .A1(n3719), .A2(n3940), .ZN(n3776) );
  NAND2_X1 U34590 ( .A1(n3941), .A2(n3776), .ZN(n3923) );
  NOR2_X1 U3460 ( .A1(n3947), .A2(n3932), .ZN(n3717) );
  NOR2_X1 U3461 ( .A1(n3964), .A2(n3944), .ZN(n3718) );
  NOR2_X1 U3462 ( .A1(n3717), .A2(n3718), .ZN(n3772) );
  AOI21_X1 U3463 ( .B1(n3923), .B2(n3772), .A(n3716), .ZN(n3906) );
  XNOR2_X1 U3464 ( .A(n3927), .B(n3915), .ZN(n3907) );
  INV_X1 U3465 ( .A(n3915), .ZN(n3908) );
  NOR2_X1 U3466 ( .A1(n3927), .A2(n3908), .ZN(n3697) );
  AOI21_X1 U34670 ( .B1(n3906), .B2(n3907), .A(n3697), .ZN(n3885) );
  NAND2_X1 U3468 ( .A1(n3794), .A2(n2894), .ZN(n2666) );
  NAND2_X1 U34690 ( .A1(n4346), .A2(n3786), .ZN(n2665) );
  INV_X1 U3470 ( .A(n2668), .ZN(n2669) );
  NAND2_X1 U34710 ( .A1(n2669), .A2(IR_REG_31__SCAN_IN), .ZN(n2670) );
  MUX2_X1 U3472 ( .A(IR_REG_31__SCAN_IN), .B(n2670), .S(IR_REG_25__SCAN_IN), 
        .Z(n2672) );
  INV_X1 U34730 ( .A(n2671), .ZN(n2677) );
  NAND2_X1 U3474 ( .A1(n2718), .A2(B_REG_SCAN_IN), .ZN(n2676) );
  NAND2_X1 U34750 ( .A1(n2686), .A2(n2685), .ZN(n2684) );
  INV_X1 U3476 ( .A(n2683), .ZN(n2727) );
  MUX2_X1 U34770 ( .A(n2676), .B(B_REG_SCAN_IN), .S(n2727), .Z(n2681) );
  NAND2_X1 U3478 ( .A1(n2677), .A2(IR_REG_31__SCAN_IN), .ZN(n2680) );
  INV_X1 U34790 ( .A(n2703), .ZN(n4345) );
  NAND2_X1 U3480 ( .A1(n2703), .A2(n2718), .ZN(n2840) );
  OAI21_X1 U34810 ( .B1(n2839), .B2(D_REG_1__SCAN_IN), .A(n2840), .ZN(n2702)
         );
  OR2_X1 U3482 ( .A1(n2686), .A2(n2685), .ZN(n2687) );
  NAND2_X1 U34830 ( .A1(n4489), .A2(n2688), .ZN(n2853) );
  AND2_X1 U3484 ( .A1(n2707), .A2(n3876), .ZN(n2845) );
  OR2_X1 U34850 ( .A1(n2847), .A2(n2845), .ZN(n2880) );
  NAND2_X1 U3486 ( .A1(n2853), .A2(n2880), .ZN(n2689) );
  NOR2_X1 U34870 ( .A1(n2858), .A2(n2689), .ZN(n2701) );
  NOR4_X1 U3488 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n2693) );
  NOR4_X1 U34890 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2692) );
  NOR4_X1 U3490 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2691) );
  NOR4_X1 U34910 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_22__SCAN_IN), .ZN(n2690) );
  NAND4_X1 U3492 ( .A1(n2693), .A2(n2692), .A3(n2691), .A4(n2690), .ZN(n2699)
         );
  NOR2_X1 U34930 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_8__SCAN_IN), .ZN(n2697) );
  NOR4_X1 U3494 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2696) );
  NOR4_X1 U34950 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2695) );
  NOR4_X1 U3496 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2694) );
  NAND4_X1 U34970 ( .A1(n2697), .A2(n2696), .A3(n2695), .A4(n2694), .ZN(n2698)
         );
  NOR2_X1 U3498 ( .A1(n2699), .A2(n2698), .ZN(n2837) );
  OR2_X1 U34990 ( .A1(n2839), .A2(n2837), .ZN(n2700) );
  NAND2_X1 U3500 ( .A1(n2683), .A2(n2703), .ZN(n2732) );
  INV_X1 U35010 ( .A(n2881), .ZN(n2705) );
  MUX2_X1 U3502 ( .A(REG1_REG_28__SCAN_IN), .B(n2711), .S(n4519), .Z(n2706) );
  INV_X1 U35030 ( .A(n2706), .ZN(n2709) );
  NOR2_X1 U3504 ( .A1(n2943), .A2(n2855), .ZN(n2885) );
  NAND2_X1 U35050 ( .A1(n3989), .A2(n3968), .ZN(n3967) );
  OAI21_X1 U35060 ( .B1(n3914), .B2(n3341), .A(n2063), .ZN(n3362) );
  NAND2_X1 U35070 ( .A1(n2709), .A2(n2265), .ZN(U3546) );
  NAND2_X1 U35080 ( .A1(n2079), .A2(n2264), .ZN(U3514) );
  INV_X1 U35090 ( .A(n4464), .ZN(n2712) );
  INV_X1 U35100 ( .A(DATAI_3_), .ZN(n2713) );
  MUX2_X1 U35110 ( .A(n2791), .B(n2713), .S(U3149), .Z(n2714) );
  INV_X1 U35120 ( .A(n2714), .ZN(U3349) );
  INV_X1 U35130 ( .A(DATAI_13_), .ZN(n4558) );
  NAND2_X1 U35140 ( .A1(n3841), .A2(STATE_REG_SCAN_IN), .ZN(n2715) );
  OAI21_X1 U35150 ( .B1(STATE_REG_SCAN_IN), .B2(n4558), .A(n2715), .ZN(U3339)
         );
  INV_X1 U35160 ( .A(DATAI_6_), .ZN(n2716) );
  INV_X1 U35170 ( .A(n2777), .ZN(n2765) );
  MUX2_X1 U35180 ( .A(n2716), .B(n2765), .S(STATE_REG_SCAN_IN), .Z(n2717) );
  INV_X1 U35190 ( .A(n2717), .ZN(U3346) );
  INV_X1 U35200 ( .A(n2718), .ZN(n2719) );
  NAND2_X1 U35210 ( .A1(n2719), .A2(STATE_REG_SCAN_IN), .ZN(n2720) );
  OAI21_X1 U35220 ( .B1(STATE_REG_SCAN_IN), .B2(n2578), .A(n2720), .ZN(U3327)
         );
  INV_X1 U35230 ( .A(DATAI_9_), .ZN(n2721) );
  INV_X1 U35240 ( .A(n3131), .ZN(n3120) );
  MUX2_X1 U35250 ( .A(n2721), .B(n3120), .S(STATE_REG_SCAN_IN), .Z(n2722) );
  INV_X1 U35260 ( .A(n2722), .ZN(U3343) );
  NAND2_X1 U35270 ( .A1(n3786), .A2(STATE_REG_SCAN_IN), .ZN(n2723) );
  OAI21_X1 U35280 ( .B1(STATE_REG_SCAN_IN), .B2(n2534), .A(n2723), .ZN(U3331)
         );
  INV_X1 U35290 ( .A(DATAI_19_), .ZN(n2724) );
  MUX2_X1 U35300 ( .A(n3876), .B(n2724), .S(U3149), .Z(n2725) );
  INV_X1 U35310 ( .A(n2725), .ZN(U3333) );
  NAND2_X1 U35320 ( .A1(n3794), .A2(STATE_REG_SCAN_IN), .ZN(n2726) );
  OAI21_X1 U35330 ( .B1(STATE_REG_SCAN_IN), .B2(n2545), .A(n2726), .ZN(U3330)
         );
  INV_X1 U35340 ( .A(DATAI_24_), .ZN(n2729) );
  NAND2_X1 U35350 ( .A1(n2727), .A2(STATE_REG_SCAN_IN), .ZN(n2728) );
  OAI21_X1 U35360 ( .B1(STATE_REG_SCAN_IN), .B2(n2729), .A(n2728), .ZN(U3328)
         );
  INV_X1 U35370 ( .A(D_REG_1__SCAN_IN), .ZN(n2731) );
  INV_X1 U35380 ( .A(n2840), .ZN(n2730) );
  AOI22_X1 U35390 ( .A1(n4462), .A2(n2731), .B1(n2730), .B2(n4464), .ZN(U3459)
         );
  INV_X1 U35400 ( .A(D_REG_0__SCAN_IN), .ZN(n4542) );
  INV_X1 U35410 ( .A(n2732), .ZN(n2733) );
  AOI22_X1 U35420 ( .A1(n4462), .A2(n4542), .B1(n2733), .B2(n4464), .ZN(U3458)
         );
  OR2_X1 U35430 ( .A1(n2982), .A2(U3149), .ZN(n3797) );
  NAND2_X1 U35440 ( .A1(n2858), .A2(n3797), .ZN(n2748) );
  INV_X1 U35450 ( .A(n2847), .ZN(n2734) );
  AOI21_X1 U35460 ( .B1(n2734), .B2(n2982), .A(n3692), .ZN(n2747) );
  INV_X1 U35470 ( .A(n2747), .ZN(n2735) );
  NOR2_X1 U35480 ( .A1(n4425), .A2(U4043), .ZN(U3148) );
  INV_X1 U35490 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n4521) );
  NAND2_X1 U35500 ( .A1(n3491), .A2(U4043), .ZN(n2736) );
  OAI21_X1 U35510 ( .B1(U4043), .B2(n4521), .A(n2736), .ZN(U3554) );
  INV_X1 U35520 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n4660) );
  NAND2_X1 U35530 ( .A1(n3580), .A2(U4043), .ZN(n2737) );
  OAI21_X1 U35540 ( .B1(U4043), .B2(n4660), .A(n2737), .ZN(U3562) );
  INV_X1 U35550 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n4678) );
  NAND2_X1 U35560 ( .A1(n3458), .A2(U4043), .ZN(n2738) );
  OAI21_X1 U35570 ( .B1(U4043), .B2(n4678), .A(n2738), .ZN(U3561) );
  INV_X1 U35580 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n2740) );
  NAND2_X1 U35590 ( .A1(n4174), .A2(U4043), .ZN(n2739) );
  OAI21_X1 U35600 ( .B1(U4043), .B2(n2740), .A(n2739), .ZN(U3564) );
  INV_X1 U35610 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n2742) );
  NAND2_X1 U35620 ( .A1(n3524), .A2(U4043), .ZN(n2741) );
  OAI21_X1 U35630 ( .B1(U4043), .B2(n2742), .A(n2741), .ZN(U3553) );
  INV_X1 U35640 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n4651) );
  NAND2_X1 U35650 ( .A1(n2825), .A2(U4043), .ZN(n2743) );
  OAI21_X1 U35660 ( .B1(U4043), .B2(n4651), .A(n2743), .ZN(U3550) );
  MUX2_X1 U35670 ( .A(n2959), .B(REG2_REG_2__SCAN_IN), .S(n4352), .Z(n3827) );
  NOR2_X1 U35680 ( .A1(n3828), .A2(n3827), .ZN(n3826) );
  AOI21_X1 U35690 ( .B1(REG2_REG_2__SCAN_IN), .B2(n4352), .A(n3826), .ZN(n2744) );
  INV_X1 U35700 ( .A(n4351), .ZN(n2758) );
  XNOR2_X1 U35710 ( .A(n2746), .B(n2758), .ZN(n2820) );
  AOI22_X1 U35720 ( .A1(n2820), .A2(REG2_REG_4__SCAN_IN), .B1(n4351), .B2(
        n2746), .ZN(n2795) );
  MUX2_X1 U35730 ( .A(n3037), .B(REG2_REG_5__SCAN_IN), .S(n4350), .Z(n2794) );
  NOR2_X1 U35740 ( .A1(n2795), .A2(n2794), .ZN(n2793) );
  XNOR2_X1 U35750 ( .A(n2778), .B(REG2_REG_6__SCAN_IN), .ZN(n2769) );
  NAND2_X1 U35760 ( .A1(n2748), .A2(n2747), .ZN(n4369) );
  NOR2_X1 U35770 ( .A1(n2750), .A2(n2749), .ZN(n4367) );
  NAND2_X1 U35780 ( .A1(n4354), .A2(n4367), .ZN(n3792) );
  XNOR2_X1 U35790 ( .A(n4352), .B(n2929), .ZN(n3824) );
  AND2_X1 U35800 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2751) );
  NAND2_X1 U35810 ( .A1(n4353), .A2(REG1_REG_1__SCAN_IN), .ZN(n2752) );
  OAI211_X1 U3582 ( .C1(n4353), .C2(REG1_REG_1__SCAN_IN), .A(n2751), .B(n2752), 
        .ZN(n3818) );
  NAND2_X1 U3583 ( .A1(n3818), .A2(n2752), .ZN(n3823) );
  NAND2_X1 U3584 ( .A1(n3824), .A2(n3823), .ZN(n2754) );
  NAND2_X1 U3585 ( .A1(n4352), .A2(REG1_REG_2__SCAN_IN), .ZN(n2753) );
  XNOR2_X1 U3586 ( .A(n2756), .B(n2791), .ZN(n2786) );
  NAND2_X1 U3587 ( .A1(n2756), .A2(n2755), .ZN(n2757) );
  NAND2_X1 U3588 ( .A1(n2759), .A2(n4351), .ZN(n2760) );
  NAND2_X1 U3589 ( .A1(n2761), .A2(n2760), .ZN(n2797) );
  MUX2_X1 U3590 ( .A(REG1_REG_5__SCAN_IN), .B(n2762), .S(n4350), .Z(n2798) );
  NAND2_X1 U3591 ( .A1(n2797), .A2(n2798), .ZN(n2796) );
  NAND2_X1 U3592 ( .A1(n4350), .A2(REG1_REG_5__SCAN_IN), .ZN(n2763) );
  XNOR2_X1 U3593 ( .A(n2771), .B(n2765), .ZN(n2770) );
  XOR2_X1 U3594 ( .A(REG1_REG_6__SCAN_IN), .B(n2770), .Z(n2767) );
  AND2_X1 U3595 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3602) );
  AOI21_X1 U3596 ( .B1(n4425), .B2(ADDR_REG_6__SCAN_IN), .A(n3602), .ZN(n2764)
         );
  OAI21_X1 U3597 ( .B1(n4438), .B2(n2765), .A(n2764), .ZN(n2766) );
  AOI21_X1 U3598 ( .B1(n4435), .B2(n2767), .A(n2766), .ZN(n2768) );
  OAI21_X1 U3599 ( .B1(n2769), .B2(n4440), .A(n2768), .ZN(U3246) );
  MUX2_X1 U3600 ( .A(n2807), .B(REG1_REG_7__SCAN_IN), .S(n4349), .Z(n2774) );
  NAND2_X1 U3601 ( .A1(n2770), .A2(REG1_REG_6__SCAN_IN), .ZN(n2773) );
  NAND2_X1 U3602 ( .A1(n2771), .A2(n2777), .ZN(n2772) );
  XOR2_X1 U3603 ( .A(n2774), .B(n2806), .Z(n2785) );
  INV_X1 U3604 ( .A(n2775), .ZN(n2776) );
  INV_X1 U3605 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3060) );
  MUX2_X1 U3606 ( .A(n3060), .B(REG2_REG_7__SCAN_IN), .S(n4349), .Z(n2779) );
  AOI21_X1 U3607 ( .B1(n2780), .B2(n2779), .A(n4440), .ZN(n2783) );
  INV_X1 U3608 ( .A(n4349), .ZN(n2808) );
  AND2_X1 U3609 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3370) );
  AOI21_X1 U3610 ( .B1(n4425), .B2(ADDR_REG_7__SCAN_IN), .A(n3370), .ZN(n2781)
         );
  OAI21_X1 U3611 ( .B1(n4438), .B2(n2808), .A(n2781), .ZN(n2782) );
  AOI21_X1 U3612 ( .B1(n2783), .B2(n2804), .A(n2782), .ZN(n2784) );
  OAI21_X1 U3613 ( .B1(n4444), .B2(n2785), .A(n2784), .ZN(U3247) );
  XOR2_X1 U3614 ( .A(n2786), .B(REG1_REG_3__SCAN_IN), .Z(n2788) );
  AOI22_X1 U3615 ( .A1(n4435), .A2(n2788), .B1(n4433), .B2(n2787), .ZN(n2790)
         );
  INV_X1 U3616 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2911) );
  NOR2_X1 U3617 ( .A1(STATE_REG_SCAN_IN), .A2(n2911), .ZN(n2996) );
  AOI21_X1 U3618 ( .B1(n4425), .B2(ADDR_REG_3__SCAN_IN), .A(n2996), .ZN(n2789)
         );
  OAI211_X1 U3619 ( .C1(n2791), .C2(n4438), .A(n2790), .B(n2789), .ZN(U3243)
         );
  INV_X1 U3620 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4677) );
  NAND2_X1 U3621 ( .A1(n2099), .A2(U4043), .ZN(n2792) );
  OAI21_X1 U3622 ( .B1(U4043), .B2(n4677), .A(n2792), .ZN(U3569) );
  AOI211_X1 U3623 ( .C1(n2795), .C2(n2794), .A(n4440), .B(n2793), .ZN(n2803)
         );
  INV_X1 U3624 ( .A(n4350), .ZN(n2801) );
  OAI211_X1 U3625 ( .C1(n2798), .C2(n2797), .A(n4435), .B(n2796), .ZN(n2800)
         );
  AND2_X1 U3626 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3489) );
  AOI21_X1 U3627 ( .B1(n4425), .B2(ADDR_REG_5__SCAN_IN), .A(n3489), .ZN(n2799)
         );
  OAI211_X1 U3628 ( .C1(n4438), .C2(n2801), .A(n2800), .B(n2799), .ZN(n2802)
         );
  OR2_X1 U3629 ( .A1(n2803), .A2(n2802), .ZN(U3245) );
  OAI21_X1 U3630 ( .B1(n3060), .B2(n2808), .A(n2804), .ZN(n2865) );
  INV_X1 U3631 ( .A(n4348), .ZN(n2812) );
  XNOR2_X1 U3632 ( .A(n2865), .B(n2812), .ZN(n2866) );
  INV_X1 U3633 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3074) );
  XNOR2_X1 U3634 ( .A(n2866), .B(n3074), .ZN(n2815) );
  AND2_X1 U3635 ( .A1(n4349), .A2(REG1_REG_7__SCAN_IN), .ZN(n2805) );
  NAND2_X1 U3636 ( .A1(n2808), .A2(n2807), .ZN(n2809) );
  AOI211_X1 U3637 ( .C1(n2309), .C2(n2810), .A(n4444), .B(n2871), .ZN(n2814)
         );
  AND2_X1 U3638 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3430) );
  AOI21_X1 U3639 ( .B1(n4425), .B2(ADDR_REG_8__SCAN_IN), .A(n3430), .ZN(n2811)
         );
  OAI21_X1 U3640 ( .B1(n4438), .B2(n2812), .A(n2811), .ZN(n2813) );
  AOI211_X1 U3641 ( .C1(n2815), .C2(n4433), .A(n2814), .B(n2813), .ZN(n2816)
         );
  INV_X1 U3642 ( .A(n2816), .ZN(U3248) );
  INV_X1 U3643 ( .A(n2855), .ZN(n2886) );
  NAND2_X1 U3644 ( .A1(n2825), .A2(n2886), .ZN(n3637) );
  INV_X1 U3645 ( .A(n3736), .ZN(n4457) );
  INV_X1 U3646 ( .A(n2708), .ZN(n2846) );
  NOR2_X1 U3647 ( .A1(n2886), .A2(n2846), .ZN(n4455) );
  INV_X1 U3648 ( .A(n4182), .ZN(n3146) );
  NOR2_X1 U3649 ( .A1(n3146), .A2(n4179), .ZN(n2818) );
  INV_X1 U3650 ( .A(n2817), .ZN(n2948) );
  OAI22_X1 U3651 ( .A1(n3736), .A2(n2818), .B1(n2817), .B2(n4127), .ZN(n4453)
         );
  AOI211_X1 U3652 ( .C1(n4489), .C2(n4457), .A(n4455), .B(n4453), .ZN(n4475)
         );
  NAND2_X1 U3653 ( .A1(n4517), .A2(REG1_REG_0__SCAN_IN), .ZN(n2819) );
  OAI21_X1 U3654 ( .B1(n4475), .B2(n4517), .A(n2819), .ZN(U3518) );
  XNOR2_X1 U3655 ( .A(n2820), .B(REG2_REG_4__SCAN_IN), .ZN(n2836) );
  NAND2_X1 U3656 ( .A1(n2055), .A2(n2825), .ZN(n2824) );
  INV_X1 U3657 ( .A(n2821), .ZN(n2822) );
  AOI22_X1 U3658 ( .A1(n3331), .A2(n2855), .B1(n2822), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2823) );
  NAND2_X1 U3659 ( .A1(n2824), .A2(n2823), .ZN(n2941) );
  INV_X4 U3660 ( .A(n3188), .ZN(n3287) );
  INV_X2 U3661 ( .A(n3311), .ZN(n3300) );
  AOI22_X1 U3662 ( .A1(n2825), .A2(n3287), .B1(n3300), .B2(n2855), .ZN(n2938)
         );
  INV_X1 U3663 ( .A(REG1_REG_0__SCAN_IN), .ZN(n3816) );
  NAND2_X1 U3664 ( .A1(n2938), .A2(n2826), .ZN(n2940) );
  XOR2_X1 U3665 ( .A(n2941), .B(n2940), .Z(n2861) );
  NOR3_X1 U3666 ( .A1(n2861), .A2(n4367), .A3(n2852), .ZN(n2830) );
  NAND2_X1 U3667 ( .A1(n4367), .A2(n4460), .ZN(n2827) );
  AND2_X1 U3668 ( .A1(n2827), .A2(n4354), .ZN(n4368) );
  INV_X1 U3669 ( .A(IR_REG_0__SCAN_IN), .ZN(n4525) );
  NOR2_X1 U3670 ( .A1(n4525), .A2(n4460), .ZN(n3813) );
  INV_X1 U3671 ( .A(n3813), .ZN(n2828) );
  OAI22_X1 U3672 ( .A1(n4368), .A2(IR_REG_0__SCAN_IN), .B1(n2828), .B2(n3792), 
        .ZN(n2829) );
  OR3_X1 U3673 ( .A1(n2830), .A2(n3801), .A3(n2829), .ZN(n3833) );
  XOR2_X1 U3674 ( .A(n2831), .B(REG1_REG_4__SCAN_IN), .Z(n2834) );
  INV_X1 U3675 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4648) );
  INV_X1 U3676 ( .A(n4425), .ZN(n4451) );
  INV_X1 U3677 ( .A(n4438), .ZN(n4448) );
  NAND2_X1 U3678 ( .A1(n4448), .A2(n4351), .ZN(n2832) );
  NAND2_X1 U3679 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3521) );
  OAI211_X1 U3680 ( .C1(n4648), .C2(n4451), .A(n2832), .B(n3521), .ZN(n2833)
         );
  AOI21_X1 U3681 ( .B1(n4435), .B2(n2834), .A(n2833), .ZN(n2835) );
  OAI211_X1 U3682 ( .C1(n2836), .C2(n4440), .A(n3833), .B(n2835), .ZN(U3244)
         );
  AND2_X1 U3683 ( .A1(n2837), .A2(D_REG_1__SCAN_IN), .ZN(n2838) );
  OR2_X1 U3684 ( .A1(n2839), .A2(n2838), .ZN(n2841) );
  NAND2_X1 U3685 ( .A1(n2841), .A2(n2840), .ZN(n2879) );
  NAND2_X1 U3686 ( .A1(n3794), .A2(n3876), .ZN(n2937) );
  INV_X1 U3687 ( .A(n2937), .ZN(n2842) );
  NAND2_X1 U3688 ( .A1(n4464), .A2(n2842), .ZN(n2843) );
  INV_X1 U3689 ( .A(n3793), .ZN(n2844) );
  NAND2_X1 U3690 ( .A1(n2856), .A2(n2844), .ZN(n2985) );
  INV_X1 U3691 ( .A(n2985), .ZN(n2851) );
  OR2_X1 U3692 ( .A1(n2846), .A2(n2845), .ZN(n2848) );
  NAND2_X1 U3693 ( .A1(n2848), .A2(n2847), .ZN(n2857) );
  NAND2_X1 U3694 ( .A1(n2857), .A2(n4198), .ZN(n2849) );
  NAND2_X1 U3695 ( .A1(n2856), .A2(n2849), .ZN(n2850) );
  NAND2_X1 U3696 ( .A1(n2850), .A2(n2880), .ZN(n2984) );
  NOR3_X1 U3697 ( .A1(n2851), .A2(n2984), .A3(n2858), .ZN(n2977) );
  NOR2_X1 U3698 ( .A1(n2856), .A2(n3793), .ZN(n2951) );
  NAND2_X1 U3699 ( .A1(n2882), .A2(n4207), .ZN(n2854) );
  AOI22_X1 U3700 ( .A1(n3629), .A2(n2948), .B1(n2855), .B2(n3579), .ZN(n2863)
         );
  INV_X1 U3701 ( .A(n2856), .ZN(n2860) );
  NOR2_X1 U3702 ( .A1(n2858), .A2(n2857), .ZN(n2859) );
  NAND2_X1 U3703 ( .A1(n2861), .A2(n3623), .ZN(n2862) );
  OAI211_X1 U3704 ( .C1(n2977), .C2(n2864), .A(n2863), .B(n2862), .ZN(U3229)
         );
  AOI22_X1 U3705 ( .A1(n2866), .A2(REG2_REG_8__SCAN_IN), .B1(n4348), .B2(n2865), .ZN(n2868) );
  INV_X1 U3706 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3121) );
  MUX2_X1 U3707 ( .A(n3121), .B(REG2_REG_9__SCAN_IN), .S(n3131), .Z(n2867) );
  AOI211_X1 U3708 ( .C1(n2868), .C2(n2867), .A(n4440), .B(n3119), .ZN(n2869)
         );
  INV_X1 U3709 ( .A(n2869), .ZN(n2878) );
  NOR2_X1 U3710 ( .A1(STATE_REG_SCAN_IN), .A2(n2401), .ZN(n3534) );
  INV_X1 U3711 ( .A(n2870), .ZN(n2872) );
  MUX2_X1 U3712 ( .A(n2873), .B(REG1_REG_9__SCAN_IN), .S(n3131), .Z(n2874) );
  AOI211_X1 U3713 ( .C1(n2875), .C2(n2874), .A(n3130), .B(n4444), .ZN(n2876)
         );
  AOI211_X1 U3714 ( .C1(n4425), .C2(ADDR_REG_9__SCAN_IN), .A(n3534), .B(n2876), 
        .ZN(n2877) );
  OAI211_X1 U3715 ( .C1(n4438), .C2(n3120), .A(n2878), .B(n2877), .ZN(U3249)
         );
  INV_X1 U3716 ( .A(n2879), .ZN(n2883) );
  NAND4_X1 U3717 ( .A1(n2883), .A2(n2882), .A3(n2881), .A4(n2880), .ZN(n2884)
         );
  NAND2_X2 U3718 ( .A1(n2884), .A2(n4187), .ZN(n4357) );
  AND2_X1 U3719 ( .A1(n4357), .A2(n3876), .ZN(n4082) );
  INV_X1 U3720 ( .A(n2885), .ZN(n2926) );
  OAI21_X1 U3721 ( .B1(n2886), .B2(n2952), .A(n2926), .ZN(n4476) );
  XNOR2_X1 U3722 ( .A(n2887), .B(n2888), .ZN(n4477) );
  OAI21_X1 U3723 ( .B1(n2133), .B2(n2132), .A(n2919), .ZN(n2892) );
  AOI22_X1 U3724 ( .A1(n3810), .A2(n4173), .B1(n4207), .B2(n2943), .ZN(n2890)
         );
  OAI21_X1 U3725 ( .B1(n2953), .B2(n4176), .A(n2890), .ZN(n2891) );
  AOI21_X1 U3726 ( .B1(n2892), .B2(n4179), .A(n2891), .ZN(n2893) );
  OAI21_X1 U3727 ( .B1(n4477), .B2(n4182), .A(n2893), .ZN(n4479) );
  NAND2_X1 U3728 ( .A1(n2895), .A2(n2894), .ZN(n3022) );
  INV_X1 U3729 ( .A(n3022), .ZN(n2896) );
  NAND2_X1 U3730 ( .A1(n4357), .A2(n2896), .ZN(n4194) );
  INV_X2 U3731 ( .A(n4357), .ZN(n4361) );
  AOI22_X1 U3732 ( .A1(n4361), .A2(REG2_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4456), .ZN(n2897) );
  OAI21_X1 U3733 ( .B1(n4477), .B2(n4194), .A(n2897), .ZN(n2898) );
  AOI21_X1 U3734 ( .B1(n4357), .B2(n4479), .A(n2898), .ZN(n2899) );
  OAI21_X1 U3735 ( .B1(n4138), .B2(n4476), .A(n2899), .ZN(U3289) );
  NAND2_X1 U3736 ( .A1(n2900), .A2(n2901), .ZN(n2902) );
  XNOR2_X1 U3737 ( .A(n2902), .B(n3733), .ZN(n4483) );
  OAI21_X1 U3738 ( .B1(n3733), .B2(n2904), .A(n2903), .ZN(n2908) );
  AOI22_X1 U3739 ( .A1(n3491), .A2(n4173), .B1(n4207), .B2(n2997), .ZN(n2906)
         );
  OAI21_X1 U3740 ( .B1(n2905), .B2(n4176), .A(n2906), .ZN(n2907) );
  AOI21_X1 U3741 ( .B1(n2908), .B2(n4179), .A(n2907), .ZN(n2909) );
  OAI21_X1 U3742 ( .B1(n4483), .B2(n4182), .A(n2909), .ZN(n4485) );
  INV_X1 U3743 ( .A(n4485), .ZN(n2916) );
  INV_X1 U3744 ( .A(n4194), .ZN(n4458) );
  INV_X1 U3745 ( .A(n4483), .ZN(n2914) );
  OAI21_X1 U3746 ( .B1(n2925), .B2(n2910), .A(n3001), .ZN(n4481) );
  AOI22_X1 U3747 ( .A1(n4361), .A2(REG2_REG_3__SCAN_IN), .B1(n4456), .B2(n2911), .ZN(n2912) );
  OAI21_X1 U3748 ( .B1(n4138), .B2(n4481), .A(n2912), .ZN(n2913) );
  AOI21_X1 U3749 ( .B1(n4458), .B2(n2914), .A(n2913), .ZN(n2915) );
  OAI21_X1 U3750 ( .B1(n2916), .B2(n4361), .A(n2915), .ZN(U3287) );
  OAI21_X1 U3751 ( .B1(n2917), .B2(n2636), .A(n2900), .ZN(n2960) );
  INV_X1 U3752 ( .A(n2960), .ZN(n2924) );
  AOI22_X1 U3753 ( .A1(n3524), .A2(n4173), .B1(n2965), .B2(n4207), .ZN(n2918)
         );
  OAI21_X1 U3754 ( .B1(n2817), .B2(n4176), .A(n2918), .ZN(n2923) );
  NAND3_X1 U3755 ( .A1(n2636), .A2(n3638), .A3(n2919), .ZN(n2920) );
  AOI21_X1 U3756 ( .B1(n2921), .B2(n2920), .A(n4132), .ZN(n2922) );
  AOI211_X1 U3757 ( .C1(n3146), .C2(n2960), .A(n2923), .B(n2922), .ZN(n2958)
         );
  OAI21_X1 U3758 ( .B1(n2924), .B2(n4482), .A(n2958), .ZN(n2934) );
  INV_X1 U3759 ( .A(n2925), .ZN(n2928) );
  NAND2_X1 U3760 ( .A1(n2926), .A2(n2965), .ZN(n2927) );
  NAND2_X1 U3761 ( .A1(n2928), .A2(n2927), .ZN(n2963) );
  OAI22_X1 U3762 ( .A1(n4281), .A2(n2963), .B1(n4519), .B2(n2929), .ZN(n2930)
         );
  AOI21_X1 U3763 ( .B1(n2934), .B2(n4519), .A(n2930), .ZN(n2931) );
  INV_X1 U3764 ( .A(n2931), .ZN(U3520) );
  INV_X1 U3765 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2932) );
  OAI22_X1 U3766 ( .A1(n4341), .A2(n2963), .B1(n4511), .B2(n2932), .ZN(n2933)
         );
  AOI21_X1 U3767 ( .B1(n2934), .B2(n4511), .A(n2933), .ZN(n2935) );
  INV_X1 U3768 ( .A(n2935), .ZN(U3471) );
  NAND2_X4 U3769 ( .A1(n2937), .A2(n2936), .ZN(n3343) );
  AND2_X1 U3770 ( .A1(n2938), .A2(n3334), .ZN(n2939) );
  NAND2_X1 U3771 ( .A1(n2942), .A2(n3287), .ZN(n2945) );
  NOR2_X1 U3772 ( .A1(n3188), .A2(n2952), .ZN(n2947) );
  AOI21_X1 U3773 ( .B1(n2057), .B2(n2948), .A(n2947), .ZN(n2968) );
  AOI211_X1 U3774 ( .C1(n2950), .C2(n2949), .A(n3619), .B(n2971), .ZN(n2957)
         );
  INV_X1 U3775 ( .A(n3579), .ZN(n3565) );
  OAI22_X1 U3776 ( .A1(n3567), .A2(n2953), .B1(n3565), .B2(n2952), .ZN(n2956)
         );
  OAI22_X1 U3777 ( .A1(n2977), .A2(n2954), .B1(n2905), .B2(n3566), .ZN(n2955)
         );
  OR3_X1 U3778 ( .A1(n2957), .A2(n2956), .A3(n2955), .ZN(U3219) );
  MUX2_X1 U3779 ( .A(n2959), .B(n2958), .S(n4357), .Z(n2962) );
  AOI22_X1 U3780 ( .A1(n2960), .A2(n4458), .B1(REG3_REG_2__SCAN_IN), .B2(n4456), .ZN(n2961) );
  OAI211_X1 U3781 ( .C1(n4138), .C2(n2963), .A(n2962), .B(n2961), .ZN(U3288)
         );
  AOI22_X1 U3782 ( .A1(n3810), .A2(n3331), .B1(n2965), .B2(n2061), .ZN(n2964)
         );
  XNOR2_X1 U3783 ( .A(n2964), .B(n3343), .ZN(n2987) );
  AOI22_X1 U3784 ( .A1(n2056), .A2(n3810), .B1(n3299), .B2(n2965), .ZN(n2988)
         );
  XNOR2_X1 U3785 ( .A(n2987), .B(n2966), .ZN(n2973) );
  INV_X1 U3786 ( .A(n2967), .ZN(n2970) );
  INV_X1 U3787 ( .A(n2968), .ZN(n2969) );
  NOR2_X1 U3788 ( .A1(n2971), .A2(n2066), .ZN(n2972) );
  NAND2_X1 U3789 ( .A1(n2972), .A2(n2973), .ZN(n2990) );
  OAI21_X1 U3790 ( .B1(n2973), .B2(n2972), .A(n2990), .ZN(n2980) );
  OAI22_X1 U3791 ( .A1(n3567), .A2(n2817), .B1(n3565), .B2(n2974), .ZN(n2979)
         );
  OAI22_X1 U3792 ( .A1(n2977), .A2(n2976), .B1(n2975), .B2(n3566), .ZN(n2978)
         );
  AOI211_X1 U3793 ( .C1(n2980), .C2(n3623), .A(n2979), .B(n2978), .ZN(n2981)
         );
  INV_X1 U3794 ( .A(n2981), .ZN(U3234) );
  NAND2_X1 U3795 ( .A1(n2821), .A2(n2982), .ZN(n2983) );
  OAI21_X1 U3796 ( .B1(n2984), .B2(n2983), .A(STATE_REG_SCAN_IN), .ZN(n2986)
         );
  INV_X1 U3797 ( .A(n3631), .ZN(n3000) );
  NAND2_X1 U3798 ( .A1(n3524), .A2(n3287), .ZN(n2992) );
  NAND2_X1 U3799 ( .A1(n3300), .A2(n2997), .ZN(n2991) );
  AOI22_X1 U3800 ( .A1(n2056), .A2(n3524), .B1(n3299), .B2(n2997), .ZN(n3174)
         );
  XNOR2_X1 U3801 ( .A(n3173), .B(n3174), .ZN(n3176) );
  XNOR2_X1 U3802 ( .A(n3177), .B(n3176), .ZN(n2994) );
  NAND2_X1 U3803 ( .A1(n2994), .A2(n3623), .ZN(n2999) );
  INV_X1 U3804 ( .A(n3491), .ZN(n3034) );
  OAI22_X1 U3805 ( .A1(n3567), .A2(n2905), .B1(n3034), .B2(n3566), .ZN(n2995)
         );
  AOI211_X1 U3806 ( .C1(n2997), .C2(n3579), .A(n2996), .B(n2995), .ZN(n2998)
         );
  OAI211_X1 U3807 ( .C1(REG3_REG_3__SCAN_IN), .C2(n3000), .A(n2999), .B(n2998), 
        .ZN(U3215) );
  INV_X1 U3808 ( .A(n4496), .ZN(n4506) );
  AOI211_X1 U3809 ( .C1(n3523), .C2(n3001), .A(n4506), .B(n3038), .ZN(n4488)
         );
  NOR2_X1 U3810 ( .A1(n4187), .A2(n3525), .ZN(n3012) );
  XNOR2_X1 U3811 ( .A(n3002), .B(n3735), .ZN(n3010) );
  NAND2_X1 U3812 ( .A1(n3004), .A2(n3735), .ZN(n3005) );
  NAND2_X1 U3813 ( .A1(n3006), .A2(n3005), .ZN(n3013) );
  AOI22_X1 U3814 ( .A1(n3524), .A2(n4130), .B1(n3523), .B2(n4207), .ZN(n3008)
         );
  NAND2_X1 U3815 ( .A1(n3809), .A2(n4173), .ZN(n3007) );
  OAI211_X1 U3816 ( .C1(n3013), .C2(n4182), .A(n3008), .B(n3007), .ZN(n3009)
         );
  AOI21_X1 U3817 ( .B1(n3010), .B2(n4179), .A(n3009), .ZN(n3011) );
  INV_X1 U3818 ( .A(n3011), .ZN(n4487) );
  AOI211_X1 U3819 ( .C1(n4488), .C2(n3876), .A(n3012), .B(n4487), .ZN(n3015)
         );
  INV_X1 U3820 ( .A(n3013), .ZN(n4490) );
  AOI22_X1 U3821 ( .A1(n4490), .A2(n4458), .B1(REG2_REG_4__SCAN_IN), .B2(n4361), .ZN(n3014) );
  OAI21_X1 U3822 ( .B1(n3015), .B2(n4361), .A(n3014), .ZN(U3286) );
  AND2_X1 U3823 ( .A1(n3649), .A2(n3660), .ZN(n3732) );
  XNOR2_X1 U3824 ( .A(n3016), .B(n3732), .ZN(n3017) );
  NAND2_X1 U3825 ( .A1(n3017), .A2(n4179), .ZN(n3019) );
  AOI22_X1 U3826 ( .A1(n3807), .A2(n4173), .B1(n3603), .B2(n4207), .ZN(n3018)
         );
  OAI211_X1 U3827 ( .C1(n3020), .C2(n4176), .A(n3019), .B(n3018), .ZN(n3045)
         );
  INV_X1 U3828 ( .A(n3045), .ZN(n3029) );
  XOR2_X1 U3829 ( .A(n3732), .B(n3021), .Z(n3046) );
  NAND2_X1 U3830 ( .A1(n4182), .A2(n3022), .ZN(n3023) );
  NAND2_X1 U3831 ( .A1(n3039), .A2(n3603), .ZN(n3024) );
  NAND2_X1 U3832 ( .A1(n3058), .A2(n3024), .ZN(n3049) );
  INV_X1 U3833 ( .A(n3025), .ZN(n3604) );
  AOI22_X1 U3834 ( .A1(n4361), .A2(REG2_REG_6__SCAN_IN), .B1(n3604), .B2(n4456), .ZN(n3026) );
  OAI21_X1 U3835 ( .B1(n4138), .B2(n3049), .A(n3026), .ZN(n3027) );
  AOI21_X1 U3836 ( .B1(n3046), .B2(n3897), .A(n3027), .ZN(n3028) );
  OAI21_X1 U3837 ( .B1(n3029), .B2(n4361), .A(n3028), .ZN(U3284) );
  INV_X1 U3838 ( .A(n3030), .ZN(n3646) );
  XOR2_X1 U3839 ( .A(n3031), .B(n3723), .Z(n4491) );
  XOR2_X1 U3840 ( .A(n3723), .B(n3032), .Z(n3036) );
  AOI22_X1 U3841 ( .A1(n3808), .A2(n4173), .B1(n4207), .B2(n3490), .ZN(n3033)
         );
  OAI21_X1 U3842 ( .B1(n3034), .B2(n4176), .A(n3033), .ZN(n3035) );
  AOI21_X1 U3843 ( .B1(n3036), .B2(n4179), .A(n3035), .ZN(n4492) );
  MUX2_X1 U3844 ( .A(n4492), .B(n3037), .S(n4361), .Z(n3044) );
  INV_X1 U3845 ( .A(n3038), .ZN(n3041) );
  INV_X1 U3846 ( .A(n3039), .ZN(n3040) );
  AOI21_X1 U3847 ( .B1(n3490), .B2(n3041), .A(n3040), .ZN(n4495) );
  INV_X1 U3848 ( .A(n3042), .ZN(n3492) );
  AOI22_X1 U3849 ( .A1(n4495), .A2(n4362), .B1(n3492), .B2(n4456), .ZN(n3043)
         );
  OAI211_X1 U3850 ( .C1(n4141), .C2(n4491), .A(n3044), .B(n3043), .ZN(U3285)
         );
  AOI21_X1 U3851 ( .B1(n3046), .B2(n4508), .A(n3045), .ZN(n3052) );
  OAI22_X1 U3852 ( .A1(n3049), .A2(n4341), .B1(n4511), .B2(n2373), .ZN(n3047)
         );
  INV_X1 U3853 ( .A(n3047), .ZN(n3048) );
  OAI21_X1 U3854 ( .B1(n3052), .B2(n4510), .A(n3048), .ZN(U3479) );
  OAI22_X1 U3855 ( .A1(n3049), .A2(n4281), .B1(n4519), .B2(n2377), .ZN(n3050)
         );
  INV_X1 U3856 ( .A(n3050), .ZN(n3051) );
  OAI21_X1 U3857 ( .B1(n3052), .B2(n4517), .A(n3051), .ZN(U3524) );
  INV_X1 U3858 ( .A(n3061), .ZN(n3730) );
  XNOR2_X1 U3859 ( .A(n3053), .B(n3730), .ZN(n3057) );
  NAND2_X1 U3860 ( .A1(n3808), .A2(n4130), .ZN(n3055) );
  NAND2_X1 U3861 ( .A1(n3806), .A2(n4173), .ZN(n3054) );
  OAI211_X1 U3862 ( .C1(n4198), .C2(n3200), .A(n3055), .B(n3054), .ZN(n3056)
         );
  AOI21_X1 U3863 ( .B1(n3057), .B2(n4179), .A(n3056), .ZN(n4503) );
  AOI21_X1 U3864 ( .B1(n3058), .B2(n3371), .A(n4506), .ZN(n3059) );
  NAND2_X1 U3865 ( .A1(n3059), .A2(n3073), .ZN(n4502) );
  INV_X1 U3866 ( .A(n4502), .ZN(n3065) );
  OAI22_X1 U3867 ( .A1(n4357), .A2(n3060), .B1(n3372), .B2(n4187), .ZN(n3064)
         );
  NOR2_X1 U3868 ( .A1(n3062), .A2(n3061), .ZN(n4500) );
  NOR3_X1 U3869 ( .A1(n4500), .A2(n4498), .A3(n4141), .ZN(n3063) );
  AOI211_X1 U3870 ( .C1(n4082), .C2(n3065), .A(n3064), .B(n3063), .ZN(n3066)
         );
  OAI21_X1 U3871 ( .B1(n4361), .B2(n4503), .A(n3066), .ZN(U3283) );
  AND2_X1 U3872 ( .A1(n3653), .A2(n3651), .ZN(n3729) );
  XNOR2_X1 U3873 ( .A(n3067), .B(n3729), .ZN(n3071) );
  OAI22_X1 U3874 ( .A1(n3068), .A2(n4127), .B1(n3207), .B2(n4198), .ZN(n3069)
         );
  AOI21_X1 U3875 ( .B1(n4130), .B2(n3807), .A(n3069), .ZN(n3070) );
  OAI21_X1 U3876 ( .B1(n3071), .B2(n4132), .A(n3070), .ZN(n3079) );
  INV_X1 U3877 ( .A(n3079), .ZN(n3078) );
  XOR2_X1 U3878 ( .A(n3729), .B(n3072), .Z(n3080) );
  NAND2_X1 U3879 ( .A1(n3080), .A2(n3897), .ZN(n3077) );
  AOI21_X1 U3880 ( .B1(n3431), .B2(n3073), .A(n3094), .ZN(n3083) );
  OAI22_X1 U3881 ( .A1(n4357), .A2(n3074), .B1(n3432), .B2(n4187), .ZN(n3075)
         );
  AOI21_X1 U3882 ( .B1(n3083), .B2(n4362), .A(n3075), .ZN(n3076) );
  OAI211_X1 U3883 ( .C1(n4361), .C2(n3078), .A(n3077), .B(n3076), .ZN(U3282)
         );
  AOI21_X1 U3884 ( .B1(n3080), .B2(n4508), .A(n3079), .ZN(n3085) );
  INV_X1 U3885 ( .A(n4341), .ZN(n4282) );
  NOR2_X1 U3886 ( .A1(n4511), .A2(n2308), .ZN(n3081) );
  AOI21_X1 U3887 ( .B1(n3083), .B2(n4282), .A(n3081), .ZN(n3082) );
  OAI21_X1 U3888 ( .B1(n3085), .B2(n4510), .A(n3082), .ZN(U3483) );
  INV_X1 U3889 ( .A(n4281), .ZN(n4195) );
  AOI22_X1 U3890 ( .A1(n3083), .A2(n4195), .B1(n4517), .B2(REG1_REG_8__SCAN_IN), .ZN(n3084) );
  OAI21_X1 U3891 ( .B1(n3085), .B2(n4517), .A(n3084), .ZN(U3526) );
  INV_X1 U3892 ( .A(n3670), .ZN(n3086) );
  XOR2_X1 U3893 ( .A(n3724), .B(n3087), .Z(n3091) );
  AOI22_X1 U3894 ( .A1(n3804), .A2(n4173), .B1(n4207), .B2(n3535), .ZN(n3088)
         );
  OAI21_X1 U3895 ( .B1(n3089), .B2(n4176), .A(n3088), .ZN(n3090) );
  AOI21_X1 U3896 ( .B1(n3091), .B2(n4179), .A(n3090), .ZN(n4504) );
  XOR2_X1 U3897 ( .A(n3724), .B(n3092), .Z(n4509) );
  OAI21_X1 U3898 ( .B1(n3094), .B2(n3093), .A(n3105), .ZN(n4505) );
  INV_X1 U3899 ( .A(n3095), .ZN(n3536) );
  AOI22_X1 U3900 ( .A1(n4361), .A2(REG2_REG_9__SCAN_IN), .B1(n3536), .B2(n4456), .ZN(n3096) );
  OAI21_X1 U3901 ( .B1(n4505), .B2(n4138), .A(n3096), .ZN(n3097) );
  AOI21_X1 U3902 ( .B1(n4509), .B2(n3897), .A(n3097), .ZN(n3098) );
  OAI21_X1 U3903 ( .B1(n4361), .B2(n4504), .A(n3098), .ZN(U3281) );
  AND2_X1 U3904 ( .A1(n3671), .A2(n3673), .ZN(n3727) );
  XOR2_X1 U3905 ( .A(n3727), .B(n3099), .Z(n3102) );
  OAI22_X1 U3906 ( .A1(n3227), .A2(n4127), .B1(n4198), .B2(n3220), .ZN(n3100)
         );
  AOI21_X1 U3907 ( .B1(n4130), .B2(n3805), .A(n3100), .ZN(n3101) );
  OAI21_X1 U3908 ( .B1(n3102), .B2(n4132), .A(n3101), .ZN(n3111) );
  INV_X1 U3909 ( .A(n3111), .ZN(n3110) );
  XOR2_X1 U3910 ( .A(n3103), .B(n3727), .Z(n3112) );
  NAND2_X1 U3911 ( .A1(n3112), .A2(n3897), .ZN(n3109) );
  INV_X1 U3912 ( .A(n3104), .ZN(n3153) );
  AOI21_X1 U3913 ( .B1(n3409), .B2(n3105), .A(n3153), .ZN(n3116) );
  OAI22_X1 U3914 ( .A1(n4357), .A2(n3106), .B1(n3410), .B2(n4187), .ZN(n3107)
         );
  AOI21_X1 U3915 ( .B1(n3116), .B2(n4362), .A(n3107), .ZN(n3108) );
  OAI211_X1 U3916 ( .C1(n4361), .C2(n3110), .A(n3109), .B(n3108), .ZN(U3280)
         );
  AOI21_X1 U3917 ( .B1(n3112), .B2(n4508), .A(n3111), .ZN(n3118) );
  AOI22_X1 U3918 ( .A1(n3116), .A2(n4195), .B1(n4517), .B2(
        REG1_REG_10__SCAN_IN), .ZN(n3113) );
  OAI21_X1 U3919 ( .B1(n3118), .B2(n4517), .A(n3113), .ZN(U3528) );
  INV_X1 U3920 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3114) );
  NOR2_X1 U3921 ( .A1(n4511), .A2(n3114), .ZN(n3115) );
  AOI21_X1 U3922 ( .B1(n3116), .B2(n4282), .A(n3115), .ZN(n3117) );
  OAI21_X1 U3923 ( .B1(n3118), .B2(n4510), .A(n3117), .ZN(U3487) );
  NAND2_X1 U3924 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4470), .ZN(n3124) );
  INV_X1 U3925 ( .A(n4470), .ZN(n4394) );
  AOI22_X1 U3926 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4470), .B1(n4394), .B2(
        n2415), .ZN(n4391) );
  NAND2_X1 U3927 ( .A1(n4472), .A2(n3122), .ZN(n3123) );
  INV_X1 U3928 ( .A(n4472), .ZN(n4383) );
  NAND2_X1 U3929 ( .A1(n3134), .A2(n3125), .ZN(n3126) );
  AND2_X1 U3930 ( .A1(n3841), .A2(REG2_REG_13__SCAN_IN), .ZN(n3842) );
  AOI21_X1 U3931 ( .B1(n4189), .B2(n2119), .A(n3842), .ZN(n3128) );
  AOI21_X1 U3932 ( .B1(n3128), .B2(n3843), .A(n4440), .ZN(n3127) );
  OAI21_X1 U3933 ( .B1(n3843), .B2(n3128), .A(n3127), .ZN(n3142) );
  NOR2_X1 U3934 ( .A1(STATE_REG_SCAN_IN), .A2(n3129), .ZN(n3556) );
  NOR2_X1 U3935 ( .A1(n3132), .A2(n4383), .ZN(n3133) );
  INV_X1 U3936 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4376) );
  AOI22_X1 U3937 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4394), .B1(n4470), .B2(
        n4279), .ZN(n4385) );
  INV_X1 U3938 ( .A(n3134), .ZN(n4469) );
  NOR2_X1 U3939 ( .A1(n3135), .A2(n4469), .ZN(n3136) );
  NOR2_X1 U3940 ( .A1(n3136), .A2(n4395), .ZN(n3139) );
  NAND2_X1 U3941 ( .A1(n3841), .A2(REG1_REG_13__SCAN_IN), .ZN(n3834) );
  OAI21_X1 U3942 ( .B1(n3841), .B2(REG1_REG_13__SCAN_IN), .A(n3834), .ZN(n3138) );
  INV_X1 U3943 ( .A(n3835), .ZN(n3137) );
  AOI211_X1 U3944 ( .C1(n3139), .C2(n3138), .A(n3137), .B(n4444), .ZN(n3140)
         );
  AOI211_X1 U3945 ( .C1(n4425), .C2(ADDR_REG_13__SCAN_IN), .A(n3556), .B(n3140), .ZN(n3141) );
  OAI211_X1 U3946 ( .C1(n4438), .C2(n2119), .A(n3142), .B(n3141), .ZN(U3253)
         );
  INV_X1 U3947 ( .A(n3144), .ZN(n3731) );
  XNOR2_X1 U3948 ( .A(n3161), .B(n3731), .ZN(n3151) );
  OAI21_X1 U3949 ( .B1(n3145), .B2(n3144), .A(n3143), .ZN(n4278) );
  NAND2_X1 U3950 ( .A1(n4278), .A2(n3146), .ZN(n3148) );
  AOI22_X1 U3951 ( .A1(n3580), .A2(n4173), .B1(n4207), .B2(n3578), .ZN(n3147)
         );
  OAI211_X1 U3952 ( .C1(n3149), .C2(n4176), .A(n3148), .B(n3147), .ZN(n3150)
         );
  AOI21_X1 U3953 ( .B1(n3151), .B2(n4179), .A(n3150), .ZN(n4276) );
  INV_X1 U3954 ( .A(n3166), .ZN(n3152) );
  OAI21_X1 U3955 ( .B1(n3153), .B2(n3226), .A(n3152), .ZN(n4342) );
  INV_X1 U3956 ( .A(n3154), .ZN(n3581) );
  AOI22_X1 U3957 ( .A1(n4361), .A2(REG2_REG_11__SCAN_IN), .B1(n3581), .B2(
        n4456), .ZN(n3155) );
  OAI21_X1 U3958 ( .B1(n4342), .B2(n4138), .A(n3155), .ZN(n3156) );
  AOI21_X1 U3959 ( .B1(n4278), .B2(n4458), .A(n3156), .ZN(n3157) );
  OAI21_X1 U3960 ( .B1(n4276), .B2(n4361), .A(n3157), .ZN(U3279) );
  NAND2_X1 U3961 ( .A1(n4168), .A2(n4166), .ZN(n3725) );
  INV_X1 U3962 ( .A(n3158), .ZN(n3159) );
  AOI21_X1 U3963 ( .B1(n3161), .B2(n3160), .A(n3159), .ZN(n4169) );
  XOR2_X1 U3964 ( .A(n3725), .B(n4169), .Z(n3164) );
  OAI22_X1 U3965 ( .A1(n4151), .A2(n4127), .B1(n4198), .B2(n3232), .ZN(n3162)
         );
  AOI21_X1 U3966 ( .B1(n4130), .B2(n3458), .A(n3162), .ZN(n3163) );
  OAI21_X1 U3967 ( .B1(n3164), .B2(n4132), .A(n3163), .ZN(n4273) );
  INV_X1 U3968 ( .A(n4273), .ZN(n3172) );
  XNOR2_X1 U3969 ( .A(n3165), .B(n3725), .ZN(n4274) );
  NOR2_X1 U3970 ( .A1(n3166), .A2(n3232), .ZN(n3167) );
  OR2_X1 U3971 ( .A1(n4184), .A2(n3167), .ZN(n4337) );
  INV_X1 U3972 ( .A(n3168), .ZN(n3459) );
  AOI22_X1 U3973 ( .A1(n4361), .A2(REG2_REG_12__SCAN_IN), .B1(n3459), .B2(
        n4456), .ZN(n3169) );
  OAI21_X1 U3974 ( .B1(n4337), .B2(n4138), .A(n3169), .ZN(n3170) );
  AOI21_X1 U3975 ( .B1(n4274), .B2(n3897), .A(n3170), .ZN(n3171) );
  OAI21_X1 U3976 ( .B1(n4361), .B2(n3172), .A(n3171), .ZN(U3278) );
  INV_X1 U3977 ( .A(n3173), .ZN(n3175) );
  NAND2_X1 U3978 ( .A1(n3491), .A2(n3287), .ZN(n3179) );
  NAND2_X1 U3979 ( .A1(n2061), .A2(n3523), .ZN(n3178) );
  NAND2_X1 U3980 ( .A1(n3179), .A2(n3178), .ZN(n3180) );
  XNOR2_X1 U3981 ( .A(n3180), .B(n3343), .ZN(n3183) );
  NOR2_X1 U3982 ( .A1(n3188), .A2(n3181), .ZN(n3182) );
  AOI21_X1 U3983 ( .B1(n2056), .B2(n3491), .A(n3182), .ZN(n3184) );
  XNOR2_X1 U3984 ( .A(n3183), .B(n3184), .ZN(n3519) );
  NAND2_X1 U3985 ( .A1(n3520), .A2(n3519), .ZN(n3518) );
  NAND2_X1 U3986 ( .A1(n3518), .A2(n3186), .ZN(n3488) );
  NOR2_X1 U3987 ( .A1(n3188), .A2(n3187), .ZN(n3189) );
  AOI21_X1 U3988 ( .B1(n2056), .B2(n3809), .A(n3189), .ZN(n3192) );
  AOI22_X1 U3989 ( .A1(n3809), .A2(n3287), .B1(n3300), .B2(n3490), .ZN(n3190)
         );
  XNOR2_X1 U3990 ( .A(n3190), .B(n3343), .ZN(n3191) );
  XOR2_X1 U3991 ( .A(n3192), .B(n3191), .Z(n3487) );
  NAND2_X1 U3992 ( .A1(n3488), .A2(n3487), .ZN(n3486) );
  INV_X1 U3993 ( .A(n3191), .ZN(n3194) );
  NAND2_X1 U3994 ( .A1(n3194), .A2(n3193), .ZN(n3195) );
  NAND2_X1 U3995 ( .A1(n3486), .A2(n3195), .ZN(n3600) );
  AOI22_X1 U3996 ( .A1(n2056), .A2(n3808), .B1(n3299), .B2(n3603), .ZN(n3597)
         );
  INV_X1 U3997 ( .A(n3597), .ZN(n3196) );
  AOI22_X1 U3998 ( .A1(n3808), .A2(n3287), .B1(n3300), .B2(n3603), .ZN(n3197)
         );
  XNOR2_X1 U3999 ( .A(n3197), .B(n3343), .ZN(n3598) );
  INV_X1 U4000 ( .A(n3598), .ZN(n3198) );
  AOI22_X1 U4001 ( .A1(n3807), .A2(n3287), .B1(n3300), .B2(n3371), .ZN(n3199)
         );
  XNOR2_X1 U4002 ( .A(n3199), .B(n3343), .ZN(n3202) );
  NOR2_X1 U4003 ( .A1(n3342), .A2(n3200), .ZN(n3201) );
  AOI21_X1 U4004 ( .B1(n2056), .B2(n3807), .A(n3201), .ZN(n3203) );
  XNOR2_X1 U4005 ( .A(n3202), .B(n3203), .ZN(n3367) );
  NAND2_X1 U4006 ( .A1(n3806), .A2(n3287), .ZN(n3205) );
  NAND2_X1 U4007 ( .A1(n2061), .A2(n3431), .ZN(n3204) );
  NAND2_X1 U4008 ( .A1(n3205), .A2(n3204), .ZN(n3206) );
  XNOR2_X1 U4009 ( .A(n3206), .B(n3334), .ZN(n3210) );
  NOR2_X1 U4010 ( .A1(n3342), .A2(n3207), .ZN(n3208) );
  AOI21_X1 U4011 ( .B1(n2056), .B2(n3806), .A(n3208), .ZN(n3209) );
  NAND2_X1 U4012 ( .A1(n3210), .A2(n3209), .ZN(n3427) );
  NAND2_X1 U4013 ( .A1(n3805), .A2(n3287), .ZN(n3212) );
  NAND2_X1 U4014 ( .A1(n3300), .A2(n3535), .ZN(n3211) );
  NAND2_X1 U4015 ( .A1(n3212), .A2(n3211), .ZN(n3213) );
  XNOR2_X1 U4016 ( .A(n3213), .B(n3343), .ZN(n3214) );
  AOI22_X1 U4017 ( .A1(n2056), .A2(n3805), .B1(n3299), .B2(n3535), .ZN(n3215)
         );
  XNOR2_X1 U4018 ( .A(n3214), .B(n3215), .ZN(n3532) );
  INV_X1 U4019 ( .A(n3214), .ZN(n3216) );
  NAND2_X1 U4020 ( .A1(n3804), .A2(n3287), .ZN(n3218) );
  NAND2_X1 U4021 ( .A1(n2061), .A2(n3409), .ZN(n3217) );
  NAND2_X1 U4022 ( .A1(n3218), .A2(n3217), .ZN(n3219) );
  XNOR2_X1 U4023 ( .A(n3219), .B(n3343), .ZN(n3222) );
  NOR2_X1 U4024 ( .A1(n3342), .A2(n3220), .ZN(n3221) );
  AOI21_X1 U4025 ( .B1(n2056), .B2(n3804), .A(n3221), .ZN(n3223) );
  XNOR2_X1 U4026 ( .A(n3222), .B(n3223), .ZN(n3407) );
  NAND2_X1 U4027 ( .A1(n3408), .A2(n3407), .ZN(n3406) );
  NAND2_X1 U4028 ( .A1(n3406), .A2(n3225), .ZN(n3572) );
  OAI22_X1 U4029 ( .A1(n3227), .A2(n3340), .B1(n3342), .B2(n3226), .ZN(n3573)
         );
  AOI22_X1 U4030 ( .A1(n3458), .A2(n3287), .B1(n2061), .B2(n3578), .ZN(n3228)
         );
  XOR2_X1 U4031 ( .A(n3343), .B(n3228), .Z(n3574) );
  NAND2_X1 U4032 ( .A1(n3580), .A2(n3287), .ZN(n3230) );
  NAND2_X1 U4033 ( .A1(n2061), .A2(n3457), .ZN(n3229) );
  NAND2_X1 U4034 ( .A1(n3230), .A2(n3229), .ZN(n3231) );
  XNOR2_X1 U4035 ( .A(n3231), .B(n3334), .ZN(n3235) );
  NOR2_X1 U4036 ( .A1(n3342), .A2(n3232), .ZN(n3233) );
  AOI21_X1 U4037 ( .B1(n2056), .B2(n3580), .A(n3233), .ZN(n3234) );
  NOR2_X1 U4038 ( .A1(n3235), .A2(n3234), .ZN(n3451) );
  NAND2_X1 U4039 ( .A1(n3235), .A2(n3234), .ZN(n3452) );
  INV_X1 U4040 ( .A(n3554), .ZN(n3239) );
  AOI22_X1 U4041 ( .A1(n3803), .A2(n3287), .B1(n3300), .B2(n4172), .ZN(n3236)
         );
  XNOR2_X1 U4042 ( .A(n3236), .B(n3343), .ZN(n3237) );
  AOI22_X1 U40430 ( .A1(n2056), .A2(n3803), .B1(n3299), .B2(n4172), .ZN(n3552)
         );
  AOI21_X1 U4044 ( .B1(n3239), .B2(n2215), .A(n3238), .ZN(n3388) );
  NAND2_X1 U4045 ( .A1(n4174), .A2(n3287), .ZN(n3241) );
  NAND2_X1 U4046 ( .A1(n2061), .A2(n4155), .ZN(n3240) );
  NAND2_X1 U4047 ( .A1(n3241), .A2(n3240), .ZN(n3242) );
  XNOR2_X1 U4048 ( .A(n3242), .B(n3343), .ZN(n3245) );
  NAND2_X1 U4049 ( .A1(n2056), .A2(n4174), .ZN(n3244) );
  NAND2_X1 U4050 ( .A1(n3299), .A2(n4155), .ZN(n3243) );
  NAND2_X1 U4051 ( .A1(n3244), .A2(n3243), .ZN(n3246) );
  NAND2_X1 U4052 ( .A1(n3245), .A2(n3246), .ZN(n3386) );
  NAND2_X1 U4053 ( .A1(n3388), .A2(n3386), .ZN(n3249) );
  INV_X1 U4054 ( .A(n3245), .ZN(n3248) );
  INV_X1 U4055 ( .A(n3246), .ZN(n3247) );
  NAND2_X1 U4056 ( .A1(n3248), .A2(n3247), .ZN(n3387) );
  NAND2_X1 U4057 ( .A1(n3249), .A2(n3387), .ZN(n3261) );
  AOI22_X1 U4058 ( .A1(n4149), .A2(n3287), .B1(n3300), .B2(n3626), .ZN(n3250)
         );
  XNOR2_X1 U4059 ( .A(n3250), .B(n3343), .ZN(n3262) );
  NAND2_X1 U4060 ( .A1(n2056), .A2(n4149), .ZN(n3252) );
  NAND2_X1 U4061 ( .A1(n3299), .A2(n3626), .ZN(n3251) );
  NAND2_X1 U4062 ( .A1(n3252), .A2(n3251), .ZN(n3621) );
  NAND2_X1 U4063 ( .A1(n4095), .A2(n3331), .ZN(n3254) );
  NAND2_X1 U4064 ( .A1(n2061), .A2(n3480), .ZN(n3253) );
  NAND2_X1 U4065 ( .A1(n3254), .A2(n3253), .ZN(n3255) );
  XNOR2_X1 U4066 ( .A(n3255), .B(n3334), .ZN(n3258) );
  INV_X1 U4067 ( .A(n3258), .ZN(n3260) );
  NOR2_X1 U4068 ( .A1(n3342), .A2(n4118), .ZN(n3256) );
  AOI21_X1 U4069 ( .B1(n2056), .B2(n4095), .A(n3256), .ZN(n3257) );
  INV_X1 U4070 ( .A(n3257), .ZN(n3259) );
  AND2_X1 U4071 ( .A1(n3258), .A2(n3257), .ZN(n3264) );
  AOI21_X1 U4072 ( .B1(n3260), .B2(n3259), .A(n3264), .ZN(n3477) );
  INV_X1 U4073 ( .A(n3262), .ZN(n3263) );
  NAND2_X1 U4074 ( .A1(n4110), .A2(n3331), .ZN(n3266) );
  NAND2_X1 U4075 ( .A1(n3300), .A2(n4098), .ZN(n3265) );
  NAND2_X1 U4076 ( .A1(n3266), .A2(n3265), .ZN(n3267) );
  XNOR2_X1 U4077 ( .A(n3267), .B(n3343), .ZN(n3271) );
  NAND2_X1 U4078 ( .A1(n2056), .A2(n4110), .ZN(n3269) );
  NAND2_X1 U4079 ( .A1(n3299), .A2(n4098), .ZN(n3268) );
  NAND2_X1 U4080 ( .A1(n3269), .A2(n3268), .ZN(n3270) );
  NAND2_X1 U4081 ( .A1(n3271), .A2(n3270), .ZN(n3497) );
  NOR2_X1 U4082 ( .A1(n3271), .A2(n3270), .ZN(n3499) );
  OAI22_X1 U4083 ( .A1(n4093), .A2(n3340), .B1(n3342), .B2(n3272), .ZN(n3586)
         );
  AOI22_X1 U4084 ( .A1(n3802), .A2(n3287), .B1(n3300), .B2(n4079), .ZN(n3273)
         );
  XOR2_X1 U4085 ( .A(n3343), .B(n3273), .Z(n3587) );
  NAND2_X1 U4086 ( .A1(n2099), .A2(n3331), .ZN(n3275) );
  NAND2_X1 U4087 ( .A1(n2061), .A2(n3420), .ZN(n3274) );
  NAND2_X1 U4088 ( .A1(n3275), .A2(n3274), .ZN(n3276) );
  XNOR2_X1 U4089 ( .A(n3276), .B(n3334), .ZN(n3279) );
  NOR2_X1 U4090 ( .A1(n3342), .A2(n4064), .ZN(n3277) );
  AOI21_X1 U4091 ( .B1(n2099), .B2(n2056), .A(n3277), .ZN(n3278) );
  NAND2_X1 U4092 ( .A1(n3279), .A2(n3278), .ZN(n3280) );
  OAI21_X1 U4093 ( .B1(n3279), .B2(n3278), .A(n3280), .ZN(n3417) );
  NAND2_X1 U4094 ( .A1(n4059), .A2(n3287), .ZN(n3282) );
  NAND2_X1 U4095 ( .A1(n2061), .A2(n4032), .ZN(n3281) );
  NAND2_X1 U4096 ( .A1(n3282), .A2(n3281), .ZN(n3283) );
  XNOR2_X1 U4097 ( .A(n3283), .B(n3334), .ZN(n3286) );
  NOR2_X1 U4098 ( .A1(n3342), .A2(n4040), .ZN(n3284) );
  AOI21_X1 U4099 ( .B1(n4059), .B2(n2056), .A(n3284), .ZN(n3285) );
  OR2_X1 U4100 ( .A1(n3286), .A2(n3285), .ZN(n3542) );
  NAND2_X1 U4101 ( .A1(n3441), .A2(n3542), .ZN(n3541) );
  NAND2_X1 U4102 ( .A1(n3286), .A2(n3285), .ZN(n3544) );
  NAND2_X1 U4103 ( .A1(n3541), .A2(n3544), .ZN(n3445) );
  NAND2_X1 U4104 ( .A1(n4001), .A2(n3287), .ZN(n3289) );
  NAND2_X1 U4105 ( .A1(n2061), .A2(n3446), .ZN(n3288) );
  NAND2_X1 U4106 ( .A1(n3289), .A2(n3288), .ZN(n3290) );
  XNOR2_X1 U4107 ( .A(n3290), .B(n3334), .ZN(n3292) );
  NOR2_X1 U4108 ( .A1(n3342), .A2(n4019), .ZN(n3291) );
  AOI21_X1 U4109 ( .B1(n4001), .B2(n2056), .A(n3291), .ZN(n3293) );
  AND2_X1 U4110 ( .A1(n3292), .A2(n3293), .ZN(n3438) );
  INV_X1 U4111 ( .A(n3292), .ZN(n3295) );
  INV_X1 U4112 ( .A(n3293), .ZN(n3294) );
  NAND2_X1 U4113 ( .A1(n3295), .A2(n3294), .ZN(n3439) );
  NAND2_X1 U4114 ( .A1(n3800), .A2(n3331), .ZN(n3297) );
  NAND2_X1 U4115 ( .A1(n3300), .A2(n4007), .ZN(n3296) );
  NAND2_X1 U4116 ( .A1(n3297), .A2(n3296), .ZN(n3298) );
  XNOR2_X1 U4117 ( .A(n3298), .B(n3343), .ZN(n3306) );
  INV_X1 U4118 ( .A(n3800), .ZN(n4015) );
  OAI22_X1 U4119 ( .A1(n4015), .A2(n3340), .B1(n3342), .B2(n3564), .ZN(n3305)
         );
  XNOR2_X1 U4120 ( .A(n3306), .B(n3305), .ZN(n3563) );
  NAND2_X1 U4121 ( .A1(n4000), .A2(n3331), .ZN(n3302) );
  NAND2_X1 U4122 ( .A1(n3300), .A2(n3988), .ZN(n3301) );
  NAND2_X1 U4123 ( .A1(n3302), .A2(n3301), .ZN(n3303) );
  XNOR2_X1 U4124 ( .A(n3303), .B(n3334), .ZN(n3309) );
  NOR2_X1 U4125 ( .A1(n3342), .A2(n3983), .ZN(n3304) );
  AOI21_X1 U4126 ( .B1(n4000), .B2(n2057), .A(n3304), .ZN(n3308) );
  XNOR2_X1 U4127 ( .A(n3309), .B(n3308), .ZN(n3397) );
  NOR2_X1 U4128 ( .A1(n3306), .A2(n3305), .ZN(n3398) );
  NOR2_X1 U4129 ( .A1(n3397), .A2(n3398), .ZN(n3307) );
  OR2_X1 U4130 ( .A1(n3309), .A2(n3308), .ZN(n3313) );
  NOR2_X1 U4131 ( .A1(n3342), .A2(n3968), .ZN(n3310) );
  AOI21_X1 U4132 ( .B1(n3985), .B2(n2056), .A(n3310), .ZN(n3314) );
  OAI22_X1 U4133 ( .A1(n3945), .A2(n3342), .B1(n3311), .B2(n3968), .ZN(n3312)
         );
  XNOR2_X1 U4134 ( .A(n3312), .B(n3343), .ZN(n3511) );
  NAND2_X1 U4135 ( .A1(n3508), .A2(n3511), .ZN(n3317) );
  NAND2_X1 U4136 ( .A1(n3399), .A2(n3313), .ZN(n3316) );
  INV_X1 U4137 ( .A(n3314), .ZN(n3315) );
  NAND2_X1 U4138 ( .A1(n3316), .A2(n3315), .ZN(n3509) );
  NAND2_X1 U4139 ( .A1(n3964), .A2(n3331), .ZN(n3319) );
  NAND2_X1 U4140 ( .A1(n2061), .A2(n3950), .ZN(n3318) );
  NAND2_X1 U4141 ( .A1(n3319), .A2(n3318), .ZN(n3320) );
  XNOR2_X1 U4142 ( .A(n3320), .B(n3334), .ZN(n3323) );
  NOR2_X1 U4143 ( .A1(n3342), .A2(n3944), .ZN(n3321) );
  AOI21_X1 U4144 ( .B1(n3964), .B2(n2056), .A(n3321), .ZN(n3322) );
  NAND2_X1 U4145 ( .A1(n3323), .A2(n3322), .ZN(n3464) );
  OR2_X1 U4146 ( .A1(n3323), .A2(n3322), .ZN(n3465) );
  NAND2_X1 U4147 ( .A1(n3947), .A2(n3331), .ZN(n3325) );
  NAND2_X1 U4148 ( .A1(n3300), .A2(n3926), .ZN(n3324) );
  NAND2_X1 U4149 ( .A1(n3325), .A2(n3324), .ZN(n3326) );
  XNOR2_X1 U4150 ( .A(n3326), .B(n3334), .ZN(n3330) );
  NOR2_X1 U4151 ( .A1(n3342), .A2(n3932), .ZN(n3327) );
  AOI21_X1 U4152 ( .B1(n3947), .B2(n2057), .A(n3327), .ZN(n3329) );
  NOR2_X1 U4153 ( .A1(n3330), .A2(n3329), .ZN(n3609) );
  NAND2_X1 U4154 ( .A1(n3927), .A2(n3331), .ZN(n3333) );
  NAND2_X1 U4155 ( .A1(n2061), .A2(n3915), .ZN(n3332) );
  NAND2_X1 U4156 ( .A1(n3333), .A2(n3332), .ZN(n3335) );
  XNOR2_X1 U4157 ( .A(n3335), .B(n3334), .ZN(n3338) );
  NOR2_X1 U4158 ( .A1(n3342), .A2(n3908), .ZN(n3336) );
  AOI21_X1 U4159 ( .B1(n3927), .B2(n2057), .A(n3336), .ZN(n3337) );
  XNOR2_X1 U4160 ( .A(n3338), .B(n3337), .ZN(n3379) );
  OAI21_X1 U4161 ( .B1(n3378), .B2(n3379), .A(n3339), .ZN(n3348) );
  OAI22_X1 U4162 ( .A1(n3381), .A2(n3340), .B1(n3342), .B2(n3341), .ZN(n3346)
         );
  OAI22_X1 U4163 ( .A1(n3381), .A2(n3342), .B1(n3311), .B2(n3341), .ZN(n3344)
         );
  XNOR2_X1 U4164 ( .A(n3344), .B(n3343), .ZN(n3345) );
  XOR2_X1 U4165 ( .A(n3346), .B(n3345), .Z(n3347) );
  XNOR2_X1 U4166 ( .A(n3348), .B(n3347), .ZN(n3354) );
  INV_X1 U4167 ( .A(n3349), .ZN(n3360) );
  NAND2_X1 U4168 ( .A1(n3927), .A2(n3628), .ZN(n3351) );
  AOI22_X1 U4169 ( .A1(n3627), .A2(n3892), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3350) );
  OAI211_X1 U4170 ( .C1(n3710), .C2(n3566), .A(n3351), .B(n3350), .ZN(n3352)
         );
  AOI21_X1 U4171 ( .B1(n3360), .B2(n3631), .A(n3352), .ZN(n3353) );
  OAI21_X1 U4172 ( .B1(n3354), .B2(n3619), .A(n3353), .ZN(U3217) );
  INV_X1 U4173 ( .A(n3355), .ZN(n3358) );
  NAND3_X1 U4174 ( .A1(IR_REG_31__SCAN_IN), .A2(STATE_REG_SCAN_IN), .A3(n2286), 
        .ZN(n3357) );
  INV_X1 U4175 ( .A(DATAI_31_), .ZN(n3356) );
  OAI22_X1 U4176 ( .A1(n3358), .A2(n3357), .B1(STATE_REG_SCAN_IN), .B2(n3356), 
        .ZN(U3321) );
  INV_X1 U4177 ( .A(n3359), .ZN(n3364) );
  AOI22_X1 U4178 ( .A1(n3360), .A2(n4456), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4361), .ZN(n3361) );
  OAI21_X1 U4179 ( .B1(n3362), .B2(n4138), .A(n3361), .ZN(n3363) );
  AOI21_X1 U4180 ( .B1(n3364), .B2(n4357), .A(n3363), .ZN(n3365) );
  OAI21_X1 U4181 ( .B1(n3366), .B2(n4141), .A(n3365), .ZN(U3262) );
  XOR2_X1 U4182 ( .A(n3368), .B(n3367), .Z(n3369) );
  NAND2_X1 U4183 ( .A1(n3369), .A2(n3623), .ZN(n3377) );
  AOI21_X1 U4184 ( .B1(n3579), .B2(n3371), .A(n3370), .ZN(n3376) );
  AOI22_X1 U4185 ( .A1(n3629), .A2(n3806), .B1(n3628), .B2(n3808), .ZN(n3375)
         );
  INV_X1 U4186 ( .A(n3372), .ZN(n3373) );
  NAND2_X1 U4187 ( .A1(n3631), .A2(n3373), .ZN(n3374) );
  NAND4_X1 U4188 ( .A1(n3377), .A2(n3376), .A3(n3375), .A4(n3374), .ZN(U3210)
         );
  XNOR2_X1 U4189 ( .A(n3378), .B(n3379), .ZN(n3385) );
  OAI22_X1 U4190 ( .A1(n3565), .A2(n3908), .B1(STATE_REG_SCAN_IN), .B2(n3380), 
        .ZN(n3383) );
  OAI22_X1 U4191 ( .A1(n3381), .A2(n3566), .B1(n3909), .B2(n3567), .ZN(n3382)
         );
  AOI211_X1 U4192 ( .C1(n3916), .C2(n3631), .A(n3383), .B(n3382), .ZN(n3384)
         );
  OAI21_X1 U4193 ( .B1(n3385), .B2(n3619), .A(n3384), .ZN(U3211) );
  NAND2_X1 U4194 ( .A1(n3387), .A2(n3386), .ZN(n3389) );
  XOR2_X1 U4195 ( .A(n3389), .B(n3388), .Z(n3390) );
  NAND2_X1 U4196 ( .A1(n3390), .A2(n3623), .ZN(n3396) );
  NAND2_X1 U4197 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4411) );
  INV_X1 U4198 ( .A(n4411), .ZN(n3391) );
  AOI21_X1 U4199 ( .B1(n3627), .B2(n4155), .A(n3391), .ZN(n3395) );
  AOI22_X1 U4200 ( .A1(n3629), .A2(n4149), .B1(n3628), .B2(n3803), .ZN(n3394)
         );
  INV_X1 U4201 ( .A(n4158), .ZN(n3392) );
  NAND2_X1 U4202 ( .A1(n3631), .A2(n3392), .ZN(n3393) );
  NAND4_X1 U4203 ( .A1(n3396), .A2(n3395), .A3(n3394), .A4(n3393), .ZN(U3212)
         );
  OAI21_X1 U4204 ( .B1(n2072), .B2(n3398), .A(n3397), .ZN(n3400) );
  NAND3_X1 U4205 ( .A1(n3400), .A2(n3623), .A3(n3399), .ZN(n3405) );
  AOI22_X1 U4206 ( .A1(n3579), .A2(n3988), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3404) );
  AOI22_X1 U4207 ( .A1(n3629), .A2(n3985), .B1(n3628), .B2(n3800), .ZN(n3403)
         );
  INV_X1 U4208 ( .A(n3401), .ZN(n3991) );
  NAND2_X1 U4209 ( .A1(n3631), .A2(n3991), .ZN(n3402) );
  NAND4_X1 U4210 ( .A1(n3405), .A2(n3404), .A3(n3403), .A4(n3402), .ZN(U3213)
         );
  OAI211_X1 U4211 ( .C1(n3408), .C2(n3407), .A(n3406), .B(n3623), .ZN(n3415)
         );
  AND2_X1 U4212 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4377) );
  AOI21_X1 U4213 ( .B1(n3627), .B2(n3409), .A(n4377), .ZN(n3414) );
  AOI22_X1 U4214 ( .A1(n3629), .A2(n3458), .B1(n3628), .B2(n3805), .ZN(n3413)
         );
  INV_X1 U4215 ( .A(n3410), .ZN(n3411) );
  NAND2_X1 U4216 ( .A1(n3631), .A2(n3411), .ZN(n3412) );
  NAND4_X1 U4217 ( .A1(n3415), .A2(n3414), .A3(n3413), .A4(n3412), .ZN(U3214)
         );
  AOI21_X1 U4218 ( .B1(n3417), .B2(n3416), .A(n2077), .ZN(n3418) );
  OR2_X1 U4219 ( .A1(n3418), .A2(n3619), .ZN(n3425) );
  NAND2_X1 U4220 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3875) );
  INV_X1 U4221 ( .A(n3875), .ZN(n3419) );
  AOI21_X1 U4222 ( .B1(n3627), .B2(n3420), .A(n3419), .ZN(n3424) );
  AOI22_X1 U4223 ( .A1(n3629), .A2(n4059), .B1(n3628), .B2(n3802), .ZN(n3423)
         );
  INV_X1 U4224 ( .A(n3421), .ZN(n4066) );
  NAND2_X1 U4225 ( .A1(n3631), .A2(n4066), .ZN(n3422) );
  NAND4_X1 U4226 ( .A1(n3425), .A2(n3424), .A3(n3423), .A4(n3422), .ZN(U3216)
         );
  NAND2_X1 U4227 ( .A1(n2096), .A2(n3427), .ZN(n3428) );
  XNOR2_X1 U4228 ( .A(n3426), .B(n3428), .ZN(n3429) );
  NAND2_X1 U4229 ( .A1(n3429), .A2(n3623), .ZN(n3437) );
  AOI21_X1 U4230 ( .B1(n3579), .B2(n3431), .A(n3430), .ZN(n3436) );
  AOI22_X1 U4231 ( .A1(n3629), .A2(n3805), .B1(n3628), .B2(n3807), .ZN(n3435)
         );
  INV_X1 U4232 ( .A(n3432), .ZN(n3433) );
  NAND2_X1 U4233 ( .A1(n3631), .A2(n3433), .ZN(n3434) );
  NAND4_X1 U4234 ( .A1(n3437), .A2(n3436), .A3(n3435), .A4(n3434), .ZN(U3218)
         );
  INV_X1 U4235 ( .A(n3438), .ZN(n3440) );
  NAND2_X1 U4236 ( .A1(n3440), .A2(n3439), .ZN(n3444) );
  INV_X1 U4237 ( .A(n3544), .ZN(n3442) );
  OAI211_X1 U4238 ( .C1(n3441), .C2(n3442), .A(n3542), .B(n3444), .ZN(n3443)
         );
  OAI211_X1 U4239 ( .C1(n3445), .C2(n3444), .A(n3623), .B(n3443), .ZN(n3450)
         );
  AOI22_X1 U4240 ( .A1(n3627), .A2(n3446), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3449) );
  AOI22_X1 U4241 ( .A1(n3629), .A2(n3800), .B1(n3628), .B2(n4059), .ZN(n3448)
         );
  NAND2_X1 U4242 ( .A1(n3631), .A2(n4020), .ZN(n3447) );
  NAND4_X1 U4243 ( .A1(n3450), .A2(n3449), .A3(n3448), .A4(n3447), .ZN(U3220)
         );
  INV_X1 U4244 ( .A(n3451), .ZN(n3453) );
  NAND2_X1 U4245 ( .A1(n3453), .A2(n3452), .ZN(n3454) );
  XNOR2_X1 U4246 ( .A(n3455), .B(n3454), .ZN(n3456) );
  NAND2_X1 U4247 ( .A1(n3456), .A2(n3623), .ZN(n3463) );
  AND2_X1 U4248 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4397) );
  AOI21_X1 U4249 ( .B1(n3627), .B2(n3457), .A(n4397), .ZN(n3462) );
  AOI22_X1 U4250 ( .A1(n3629), .A2(n3803), .B1(n3628), .B2(n3458), .ZN(n3461)
         );
  NAND2_X1 U4251 ( .A1(n3631), .A2(n3459), .ZN(n3460) );
  NAND4_X1 U4252 ( .A1(n3463), .A2(n3462), .A3(n3461), .A4(n3460), .ZN(U3221)
         );
  NAND2_X1 U4253 ( .A1(n3465), .A2(n3464), .ZN(n3467) );
  XOR2_X1 U4254 ( .A(n3467), .B(n3466), .Z(n3473) );
  INV_X1 U4255 ( .A(n3468), .ZN(n3953) );
  OAI22_X1 U4256 ( .A1(n3565), .A2(n3944), .B1(STATE_REG_SCAN_IN), .B2(n3469), 
        .ZN(n3471) );
  OAI22_X1 U4257 ( .A1(n3909), .A2(n3566), .B1(n3945), .B2(n3567), .ZN(n3470)
         );
  AOI211_X1 U4258 ( .C1(n3953), .C2(n3631), .A(n3471), .B(n3470), .ZN(n3472)
         );
  OAI21_X1 U4259 ( .B1(n3473), .B2(n3619), .A(n3472), .ZN(U3222) );
  INV_X1 U4260 ( .A(n3474), .ZN(n3476) );
  OAI21_X1 U4261 ( .B1(n3476), .B2(n3621), .A(n3475), .ZN(n3478) );
  XNOR2_X1 U4262 ( .A(n3478), .B(n3477), .ZN(n3479) );
  NAND2_X1 U4263 ( .A1(n3479), .A2(n3623), .ZN(n3485) );
  AND2_X1 U4264 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4414) );
  AOI21_X1 U4265 ( .B1(n3627), .B2(n3480), .A(n4414), .ZN(n3484) );
  AOI22_X1 U4266 ( .A1(n3629), .A2(n4110), .B1(n3628), .B2(n4149), .ZN(n3483)
         );
  INV_X1 U4267 ( .A(n4115), .ZN(n3481) );
  NAND2_X1 U4268 ( .A1(n3631), .A2(n3481), .ZN(n3482) );
  NAND4_X1 U4269 ( .A1(n3485), .A2(n3484), .A3(n3483), .A4(n3482), .ZN(U3223)
         );
  OAI211_X1 U4270 ( .C1(n3488), .C2(n3487), .A(n3486), .B(n3623), .ZN(n3496)
         );
  AOI21_X1 U4271 ( .B1(n3627), .B2(n3490), .A(n3489), .ZN(n3495) );
  AOI22_X1 U4272 ( .A1(n3629), .A2(n3808), .B1(n3628), .B2(n3491), .ZN(n3494)
         );
  NAND2_X1 U4273 ( .A1(n3631), .A2(n3492), .ZN(n3493) );
  NAND4_X1 U4274 ( .A1(n3496), .A2(n3495), .A3(n3494), .A4(n3493), .ZN(U3224)
         );
  INV_X1 U4275 ( .A(n3497), .ZN(n3498) );
  NOR2_X1 U4276 ( .A1(n3499), .A2(n3498), .ZN(n3500) );
  XNOR2_X1 U4277 ( .A(n3501), .B(n3500), .ZN(n3502) );
  NAND2_X1 U4278 ( .A1(n3502), .A2(n3623), .ZN(n3507) );
  NOR2_X1 U4279 ( .A1(STATE_REG_SCAN_IN), .A2(n4556), .ZN(n4424) );
  AOI21_X1 U4280 ( .B1(n3579), .B2(n4098), .A(n4424), .ZN(n3506) );
  AOI22_X1 U4281 ( .A1(n3629), .A2(n3802), .B1(n3628), .B2(n4095), .ZN(n3505)
         );
  INV_X1 U4282 ( .A(n3503), .ZN(n4101) );
  NAND2_X1 U4283 ( .A1(n3631), .A2(n4101), .ZN(n3504) );
  NAND4_X1 U4284 ( .A1(n3507), .A2(n3506), .A3(n3505), .A4(n3504), .ZN(U3225)
         );
  NAND2_X1 U4285 ( .A1(n3509), .A2(n3508), .ZN(n3510) );
  XOR2_X1 U4286 ( .A(n3511), .B(n3510), .Z(n3517) );
  OAI22_X1 U4287 ( .A1(n3565), .A2(n3968), .B1(STATE_REG_SCAN_IN), .B2(n3512), 
        .ZN(n3515) );
  INV_X1 U4288 ( .A(n3964), .ZN(n3513) );
  OAI22_X1 U4289 ( .A1(n3513), .A2(n3566), .B1(n4706), .B2(n3567), .ZN(n3514)
         );
  AOI211_X1 U4290 ( .C1(n3969), .C2(n3631), .A(n3515), .B(n3514), .ZN(n3516)
         );
  OAI21_X1 U4291 ( .B1(n3517), .B2(n3619), .A(n3516), .ZN(U3226) );
  OAI211_X1 U4292 ( .C1(n3520), .C2(n3519), .A(n3518), .B(n3623), .ZN(n3530)
         );
  INV_X1 U4293 ( .A(n3521), .ZN(n3522) );
  AOI21_X1 U4294 ( .B1(n3579), .B2(n3523), .A(n3522), .ZN(n3529) );
  AOI22_X1 U4295 ( .A1(n3629), .A2(n3809), .B1(n3628), .B2(n3524), .ZN(n3528)
         );
  INV_X1 U4296 ( .A(n3525), .ZN(n3526) );
  NAND2_X1 U4297 ( .A1(n3631), .A2(n3526), .ZN(n3527) );
  NAND4_X1 U4298 ( .A1(n3530), .A2(n3529), .A3(n3528), .A4(n3527), .ZN(U3227)
         );
  XNOR2_X1 U4299 ( .A(n3531), .B(n3532), .ZN(n3533) );
  NAND2_X1 U4300 ( .A1(n3533), .A2(n3623), .ZN(n3540) );
  AOI21_X1 U4301 ( .B1(n3579), .B2(n3535), .A(n3534), .ZN(n3539) );
  AOI22_X1 U4302 ( .A1(n3629), .A2(n3804), .B1(n3628), .B2(n3806), .ZN(n3538)
         );
  NAND2_X1 U4303 ( .A1(n3631), .A2(n3536), .ZN(n3537) );
  NAND4_X1 U4304 ( .A1(n3540), .A2(n3539), .A3(n3538), .A4(n3537), .ZN(U3228)
         );
  INV_X1 U4305 ( .A(n3541), .ZN(n3545) );
  AOI21_X1 U4306 ( .B1(n3542), .B2(n3544), .A(n3441), .ZN(n3543) );
  AOI21_X1 U4307 ( .B1(n3545), .B2(n3544), .A(n3543), .ZN(n3551) );
  OAI22_X1 U4308 ( .A1(n3565), .A2(n4040), .B1(STATE_REG_SCAN_IN), .B2(n3546), 
        .ZN(n3549) );
  OAI22_X1 U4309 ( .A1(n3567), .A2(n3547), .B1(n4034), .B2(n3566), .ZN(n3548)
         );
  AOI211_X1 U4310 ( .C1(n4041), .C2(n3631), .A(n3549), .B(n3548), .ZN(n3550)
         );
  OAI21_X1 U4311 ( .B1(n3551), .B2(n3619), .A(n3550), .ZN(U3230) );
  XNOR2_X1 U4312 ( .A(n2215), .B(n3552), .ZN(n3553) );
  XNOR2_X1 U4313 ( .A(n3554), .B(n3553), .ZN(n3555) );
  NAND2_X1 U4314 ( .A1(n3555), .A2(n3623), .ZN(n3561) );
  AOI21_X1 U4315 ( .B1(n3579), .B2(n4172), .A(n3556), .ZN(n3560) );
  AOI22_X1 U4316 ( .A1(n3629), .A2(n4174), .B1(n3628), .B2(n3580), .ZN(n3559)
         );
  INV_X1 U4317 ( .A(n4188), .ZN(n3557) );
  NAND2_X1 U4318 ( .A1(n3631), .A2(n3557), .ZN(n3558) );
  NAND4_X1 U4319 ( .A1(n3561), .A2(n3560), .A3(n3559), .A4(n3558), .ZN(U3231)
         );
  AOI21_X1 U4320 ( .B1(n3563), .B2(n3562), .A(n2072), .ZN(n3571) );
  OAI22_X1 U4321 ( .A1(n3565), .A2(n3564), .B1(STATE_REG_SCAN_IN), .B2(n4523), 
        .ZN(n3569) );
  OAI22_X1 U4322 ( .A1(n3567), .A2(n4034), .B1(n4706), .B2(n3566), .ZN(n3568)
         );
  AOI211_X1 U4323 ( .C1(n4006), .C2(n3631), .A(n3569), .B(n3568), .ZN(n3570)
         );
  OAI21_X1 U4324 ( .B1(n3571), .B2(n3619), .A(n3570), .ZN(U3232) );
  XNOR2_X1 U4325 ( .A(n3574), .B(n3573), .ZN(n3575) );
  XNOR2_X1 U4326 ( .A(n3572), .B(n3575), .ZN(n3576) );
  NAND2_X1 U4327 ( .A1(n3576), .A2(n3623), .ZN(n3585) );
  NOR2_X1 U4328 ( .A1(STATE_REG_SCAN_IN), .A2(n3577), .ZN(n4387) );
  AOI21_X1 U4329 ( .B1(n3579), .B2(n3578), .A(n4387), .ZN(n3584) );
  AOI22_X1 U4330 ( .A1(n3629), .A2(n3580), .B1(n3628), .B2(n3804), .ZN(n3583)
         );
  NAND2_X1 U4331 ( .A1(n3631), .A2(n3581), .ZN(n3582) );
  NAND4_X1 U4332 ( .A1(n3585), .A2(n3584), .A3(n3583), .A4(n3582), .ZN(U3233)
         );
  XNOR2_X1 U4333 ( .A(n3587), .B(n3586), .ZN(n3588) );
  XNOR2_X1 U4334 ( .A(n3589), .B(n3588), .ZN(n3590) );
  NAND2_X1 U4335 ( .A1(n3590), .A2(n3623), .ZN(n3596) );
  NAND2_X1 U4336 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4449) );
  INV_X1 U4337 ( .A(n4449), .ZN(n3591) );
  AOI21_X1 U4338 ( .B1(n3627), .B2(n4079), .A(n3591), .ZN(n3595) );
  AOI22_X1 U4339 ( .A1(n3629), .A2(n2099), .B1(n3628), .B2(n4110), .ZN(n3594)
         );
  INV_X1 U4340 ( .A(n3592), .ZN(n4083) );
  NAND2_X1 U4341 ( .A1(n3631), .A2(n4083), .ZN(n3593) );
  NAND4_X1 U4342 ( .A1(n3596), .A2(n3595), .A3(n3594), .A4(n3593), .ZN(U3235)
         );
  XNOR2_X1 U4343 ( .A(n3598), .B(n3597), .ZN(n3599) );
  XNOR2_X1 U4344 ( .A(n3600), .B(n3599), .ZN(n3601) );
  NAND2_X1 U4345 ( .A1(n3601), .A2(n3623), .ZN(n3608) );
  AOI21_X1 U4346 ( .B1(n3627), .B2(n3603), .A(n3602), .ZN(n3607) );
  AOI22_X1 U4347 ( .A1(n3629), .A2(n3807), .B1(n3628), .B2(n3809), .ZN(n3606)
         );
  NAND2_X1 U4348 ( .A1(n3631), .A2(n3604), .ZN(n3605) );
  NAND4_X1 U4349 ( .A1(n3608), .A2(n3607), .A3(n3606), .A4(n3605), .ZN(U3236)
         );
  NOR2_X1 U4350 ( .A1(n3609), .A2(n2087), .ZN(n3610) );
  XNOR2_X1 U4351 ( .A(n3611), .B(n3610), .ZN(n3620) );
  NAND2_X1 U4352 ( .A1(n3964), .A2(n3628), .ZN(n3615) );
  NOR2_X1 U4353 ( .A1(n3612), .A2(STATE_REG_SCAN_IN), .ZN(n3613) );
  AOI21_X1 U4354 ( .B1(n3627), .B2(n3926), .A(n3613), .ZN(n3614) );
  NAND2_X1 U4355 ( .A1(n3615), .A2(n3614), .ZN(n3616) );
  AOI21_X1 U4356 ( .B1(n3927), .B2(n3629), .A(n3616), .ZN(n3618) );
  NAND2_X1 U4357 ( .A1(n3934), .A2(n3631), .ZN(n3617) );
  OAI211_X1 U4358 ( .C1(n3620), .C2(n3619), .A(n3618), .B(n3617), .ZN(U3237)
         );
  NAND2_X1 U4359 ( .A1(n3474), .A2(n3475), .ZN(n3622) );
  XNOR2_X1 U4360 ( .A(n3622), .B(n3621), .ZN(n3624) );
  NAND2_X1 U4361 ( .A1(n3624), .A2(n3623), .ZN(n3635) );
  NOR2_X1 U4362 ( .A1(STATE_REG_SCAN_IN), .A2(n3625), .ZN(n3853) );
  AOI21_X1 U4363 ( .B1(n3627), .B2(n3626), .A(n3853), .ZN(n3634) );
  AOI22_X1 U4364 ( .A1(n3629), .A2(n4095), .B1(n3628), .B2(n4174), .ZN(n3633)
         );
  INV_X1 U4365 ( .A(n3630), .ZN(n4136) );
  NAND2_X1 U4366 ( .A1(n3631), .A2(n4136), .ZN(n3632) );
  NAND4_X1 U4367 ( .A1(n3635), .A2(n3634), .A3(n3633), .A4(n3632), .ZN(U3238)
         );
  OAI211_X1 U4368 ( .C1(n2132), .C2(n3786), .A(n3637), .B(n3636), .ZN(n3639)
         );
  NAND3_X1 U4369 ( .A1(n3639), .A2(n2638), .A3(n3638), .ZN(n3642) );
  NAND3_X1 U4370 ( .A1(n3642), .A2(n3641), .A3(n3640), .ZN(n3645) );
  NAND3_X1 U4371 ( .A1(n3645), .A2(n3644), .A3(n3643), .ZN(n3648) );
  NAND4_X1 U4372 ( .A1(n3648), .A2(n3647), .A3(n3646), .A4(n3660), .ZN(n3650)
         );
  NAND3_X1 U4373 ( .A1(n3650), .A2(n3730), .A3(n3649), .ZN(n3657) );
  AND2_X1 U4374 ( .A1(n3652), .A2(n3651), .ZN(n3661) );
  INV_X1 U4375 ( .A(n3653), .ZN(n3656) );
  INV_X1 U4376 ( .A(n3654), .ZN(n3655) );
  AOI211_X1 U4377 ( .C1(n3657), .C2(n3661), .A(n3656), .B(n3655), .ZN(n3669)
         );
  NAND2_X1 U4378 ( .A1(n3659), .A2(n3658), .ZN(n3668) );
  INV_X1 U4379 ( .A(n3660), .ZN(n3664) );
  INV_X1 U4380 ( .A(n3661), .ZN(n3663) );
  NOR3_X1 U4381 ( .A1(n3664), .A2(n3663), .A3(n3662), .ZN(n3666) );
  INV_X1 U4382 ( .A(n3671), .ZN(n3665) );
  NAND2_X1 U4383 ( .A1(n3668), .A2(n3677), .ZN(n3755) );
  OAI21_X1 U4384 ( .B1(n3666), .B2(n3665), .A(n3755), .ZN(n3667) );
  OAI21_X1 U4385 ( .B1(n3669), .B2(n3668), .A(n3667), .ZN(n3675) );
  NAND2_X1 U4386 ( .A1(n3671), .A2(n3670), .ZN(n3672) );
  NAND4_X1 U4387 ( .A1(n3675), .A2(n3674), .A3(n3673), .A4(n3672), .ZN(n3681)
         );
  INV_X1 U4388 ( .A(n3676), .ZN(n3678) );
  NAND2_X1 U4389 ( .A1(n4124), .A2(n3677), .ZN(n3756) );
  OAI21_X1 U4390 ( .B1(n3678), .B2(n3756), .A(n3755), .ZN(n3680) );
  AOI21_X1 U4391 ( .B1(n3681), .B2(n3680), .A(n2130), .ZN(n3684) );
  INV_X1 U4392 ( .A(n3759), .ZN(n3683) );
  INV_X1 U4393 ( .A(n3757), .ZN(n3682) );
  OAI21_X1 U4394 ( .B1(n3684), .B2(n3683), .A(n3682), .ZN(n3685) );
  AOI211_X1 U4395 ( .C1(n3685), .C2(n3763), .A(n3761), .B(n3720), .ZN(n3686)
         );
  NOR2_X1 U4396 ( .A1(n3686), .A2(n3766), .ZN(n3688) );
  OAI21_X1 U4397 ( .B1(n3688), .B2(n3687), .A(n3768), .ZN(n3689) );
  NAND2_X1 U4398 ( .A1(n3776), .A2(n3689), .ZN(n3696) );
  INV_X1 U4399 ( .A(n3927), .ZN(n3690) );
  NOR2_X1 U4400 ( .A1(n3690), .A2(n3915), .ZN(n3695) );
  INV_X1 U4401 ( .A(n3710), .ZN(n3799) );
  INV_X1 U4402 ( .A(DATAI_29_), .ZN(n3691) );
  INV_X1 U4403 ( .A(n3898), .ZN(n3693) );
  NAND2_X1 U4404 ( .A1(n3799), .A2(n3693), .ZN(n3745) );
  NAND2_X1 U4405 ( .A1(n3745), .A2(n3882), .ZN(n3711) );
  NOR2_X1 U4406 ( .A1(n3716), .A2(n3711), .ZN(n3778) );
  INV_X1 U4407 ( .A(n3778), .ZN(n3694) );
  AOI211_X1 U4408 ( .C1(n3772), .C2(n3696), .A(n3695), .B(n3694), .ZN(n3712)
         );
  NOR2_X1 U4409 ( .A1(n3698), .A2(n3697), .ZN(n3769) );
  INV_X1 U4410 ( .A(REG1_REG_30__SCAN_IN), .ZN(n3702) );
  NAND2_X1 U4411 ( .A1(n3704), .A2(REG0_REG_30__SCAN_IN), .ZN(n3701) );
  INV_X1 U4412 ( .A(REG2_REG_30__SCAN_IN), .ZN(n3699) );
  OR2_X1 U4413 ( .A1(n2060), .A2(n3699), .ZN(n3700) );
  OAI211_X1 U4414 ( .C1(n2059), .C2(n3702), .A(n3701), .B(n3700), .ZN(n3887)
         );
  NAND2_X1 U4415 ( .A1(n3708), .A2(DATAI_30_), .ZN(n4203) );
  OR2_X1 U4416 ( .A1(n3887), .A2(n4203), .ZN(n3709) );
  INV_X1 U4417 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3707) );
  INV_X1 U4418 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3703) );
  OR2_X1 U4419 ( .A1(n2060), .A2(n3703), .ZN(n3706) );
  NAND2_X1 U4420 ( .A1(n3704), .A2(REG0_REG_31__SCAN_IN), .ZN(n3705) );
  OAI211_X1 U4421 ( .C1(n2609), .C2(n3707), .A(n3706), .B(n3705), .ZN(n4197)
         );
  NAND2_X1 U4422 ( .A1(n3708), .A2(DATAI_31_), .ZN(n4199) );
  NAND2_X1 U4423 ( .A1(n4197), .A2(n4199), .ZN(n3713) );
  AND2_X1 U4424 ( .A1(n3709), .A2(n3713), .ZN(n3770) );
  NAND2_X1 U4425 ( .A1(n3710), .A2(n3898), .ZN(n3771) );
  OAI211_X1 U4426 ( .C1(n3769), .C2(n3711), .A(n3770), .B(n3771), .ZN(n3777)
         );
  OR2_X1 U4427 ( .A1(n3712), .A2(n3777), .ZN(n3715) );
  OR2_X1 U4428 ( .A1(n4197), .A2(n4199), .ZN(n3779) );
  NAND2_X1 U4429 ( .A1(n3887), .A2(n4203), .ZN(n3780) );
  NAND2_X1 U4430 ( .A1(n3779), .A2(n3780), .ZN(n3721) );
  NAND2_X1 U4431 ( .A1(n3721), .A2(n3713), .ZN(n3714) );
  NAND2_X1 U4432 ( .A1(n3715), .A2(n3714), .ZN(n3790) );
  NOR2_X1 U4433 ( .A1(n3717), .A2(n3716), .ZN(n3925) );
  INV_X1 U4434 ( .A(n3925), .ZN(n3752) );
  INV_X1 U4435 ( .A(n3718), .ZN(n3922) );
  NAND2_X1 U4436 ( .A1(n3922), .A2(n3719), .ZN(n3943) );
  INV_X1 U4437 ( .A(n3943), .ZN(n3744) );
  XNOR2_X1 U4438 ( .A(n3803), .B(n4172), .ZN(n4170) );
  INV_X1 U4439 ( .A(n3720), .ZN(n3977) );
  NAND2_X1 U4440 ( .A1(n3977), .A2(n3975), .ZN(n4013) );
  INV_X1 U4441 ( .A(n3721), .ZN(n3722) );
  NAND4_X1 U4442 ( .A1(n3724), .A2(n3723), .A3(n3722), .A4(n3770), .ZN(n3726)
         );
  NAND2_X1 U4443 ( .A1(n4051), .A2(n4050), .ZN(n4091) );
  NOR4_X1 U4444 ( .A1(n4013), .A2(n3726), .A3(n4091), .A4(n3725), .ZN(n3743)
         );
  NAND3_X1 U4445 ( .A1(n3978), .A2(n3728), .A3(n3727), .ZN(n3741) );
  NAND4_X1 U4446 ( .A1(n4072), .A2(n3731), .A3(n3730), .A4(n3729), .ZN(n3740)
         );
  NAND4_X1 U4447 ( .A1(n3735), .A2(n3734), .A3(n3733), .A4(n3732), .ZN(n3739)
         );
  INV_X1 U4448 ( .A(n4125), .ZN(n3737) );
  NAND4_X1 U4449 ( .A1(n4148), .A2(n2133), .A3(n3737), .A4(n3736), .ZN(n3738)
         );
  NOR4_X1 U4450 ( .A1(n3741), .A2(n3740), .A3(n3739), .A4(n3738), .ZN(n3742)
         );
  NAND4_X1 U4451 ( .A1(n3744), .A2(n4170), .A3(n3743), .A4(n3742), .ZN(n3751)
         );
  NAND2_X1 U4452 ( .A1(n3745), .A2(n3771), .ZN(n3895) );
  NAND2_X1 U4453 ( .A1(n3746), .A2(n3940), .ZN(n3961) );
  INV_X1 U4454 ( .A(n3961), .ZN(n3749) );
  XNOR2_X1 U4455 ( .A(n4000), .B(n3988), .ZN(n3980) );
  XNOR2_X1 U4456 ( .A(n2099), .B(n4064), .ZN(n4048) );
  INV_X1 U4457 ( .A(n4048), .ZN(n4056) );
  NAND2_X1 U4458 ( .A1(n3748), .A2(n3747), .ZN(n4030) );
  NAND4_X1 U4459 ( .A1(n3749), .A2(n3980), .A3(n4056), .A4(n4030), .ZN(n3750)
         );
  NOR4_X1 U4460 ( .A1(n3752), .A2(n3751), .A3(n3895), .A4(n3750), .ZN(n3754)
         );
  INV_X1 U4461 ( .A(n3893), .ZN(n3753) );
  NAND3_X1 U4462 ( .A1(n3754), .A2(n3753), .A3(n3907), .ZN(n3788) );
  INV_X1 U4463 ( .A(n4203), .ZN(n4208) );
  OAI21_X1 U4464 ( .B1(n4147), .B2(n3756), .A(n3755), .ZN(n3758) );
  AOI211_X1 U4465 ( .C1(n3759), .C2(n3758), .A(n2130), .B(n3757), .ZN(n3760)
         );
  INV_X1 U4466 ( .A(n3760), .ZN(n3762) );
  AOI21_X1 U4467 ( .B1(n3763), .B2(n3762), .A(n3761), .ZN(n3765) );
  OAI21_X1 U4468 ( .B1(n3766), .B2(n3765), .A(n3764), .ZN(n3767) );
  NAND2_X1 U4469 ( .A1(n3768), .A2(n3767), .ZN(n3775) );
  NAND3_X1 U4470 ( .A1(n3771), .A2(n3770), .A3(n3769), .ZN(n3774) );
  INV_X1 U4471 ( .A(n3772), .ZN(n3773) );
  AOI211_X1 U4472 ( .C1(n3776), .C2(n3775), .A(n3774), .B(n3773), .ZN(n3784)
         );
  AOI21_X1 U4473 ( .B1(n3907), .B2(n3778), .A(n3777), .ZN(n3783) );
  INV_X1 U4474 ( .A(n3779), .ZN(n3782) );
  NOR2_X1 U4475 ( .A1(n3780), .A2(n4199), .ZN(n3781) );
  NOR4_X1 U4476 ( .A1(n3784), .A2(n3783), .A3(n3782), .A4(n3781), .ZN(n3785)
         );
  AOI21_X1 U4477 ( .B1(n4208), .B2(n4199), .A(n3785), .ZN(n3787) );
  MUX2_X1 U4478 ( .A(n3788), .B(n3787), .S(n3786), .Z(n3789) );
  MUX2_X1 U4479 ( .A(n3790), .B(n3789), .S(n4346), .Z(n3791) );
  XNOR2_X1 U4480 ( .A(n3791), .B(n3876), .ZN(n3798) );
  NOR2_X1 U4481 ( .A1(n3793), .A2(n3792), .ZN(n3796) );
  OAI21_X1 U4482 ( .B1(n3797), .B2(n3794), .A(B_REG_SCAN_IN), .ZN(n3795) );
  OAI22_X1 U4483 ( .A1(n3798), .A2(n3797), .B1(n3796), .B2(n3795), .ZN(U3239)
         );
  MUX2_X1 U4484 ( .A(DATAO_REG_31__SCAN_IN), .B(n4197), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4485 ( .A(DATAO_REG_30__SCAN_IN), .B(n3887), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4486 ( .A(DATAO_REG_29__SCAN_IN), .B(n3799), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4487 ( .A(DATAO_REG_28__SCAN_IN), .B(n3911), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4488 ( .A(DATAO_REG_27__SCAN_IN), .B(n3927), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4489 ( .A(DATAO_REG_26__SCAN_IN), .B(n3947), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4490 ( .A(DATAO_REG_25__SCAN_IN), .B(n3964), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4491 ( .A(n3985), .B(DATAO_REG_24__SCAN_IN), .S(n3801), .Z(U3574)
         );
  MUX2_X1 U4492 ( .A(DATAO_REG_22__SCAN_IN), .B(n3800), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4493 ( .A(n4001), .B(DATAO_REG_21__SCAN_IN), .S(n3801), .Z(U3571)
         );
  MUX2_X1 U4494 ( .A(n4059), .B(DATAO_REG_20__SCAN_IN), .S(n3801), .Z(U3570)
         );
  MUX2_X1 U4495 ( .A(DATAO_REG_18__SCAN_IN), .B(n3802), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4496 ( .A(DATAO_REG_17__SCAN_IN), .B(n4110), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4497 ( .A(DATAO_REG_16__SCAN_IN), .B(n4095), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4498 ( .A(DATAO_REG_15__SCAN_IN), .B(n4149), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4499 ( .A(DATAO_REG_13__SCAN_IN), .B(n3803), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4500 ( .A(DATAO_REG_10__SCAN_IN), .B(n3804), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4501 ( .A(DATAO_REG_9__SCAN_IN), .B(n3805), .S(U4043), .Z(U3559) );
  MUX2_X1 U4502 ( .A(DATAO_REG_8__SCAN_IN), .B(n3806), .S(U4043), .Z(U3558) );
  MUX2_X1 U4503 ( .A(DATAO_REG_7__SCAN_IN), .B(n3807), .S(U4043), .Z(U3557) );
  MUX2_X1 U4504 ( .A(DATAO_REG_6__SCAN_IN), .B(n3808), .S(U4043), .Z(U3556) );
  MUX2_X1 U4505 ( .A(DATAO_REG_5__SCAN_IN), .B(n3809), .S(U4043), .Z(U3555) );
  MUX2_X1 U4506 ( .A(DATAO_REG_2__SCAN_IN), .B(n3810), .S(U4043), .Z(U3552) );
  MUX2_X1 U4507 ( .A(DATAO_REG_1__SCAN_IN), .B(n2948), .S(U4043), .Z(U3551) );
  INV_X1 U4508 ( .A(n3811), .ZN(n3812) );
  OAI211_X1 U4509 ( .C1(n3814), .C2(n3813), .A(n4433), .B(n3812), .ZN(n3822)
         );
  MUX2_X1 U4510 ( .A(n2332), .B(REG1_REG_1__SCAN_IN), .S(n4353), .Z(n3815) );
  OAI21_X1 U4511 ( .B1(n4525), .B2(n3816), .A(n3815), .ZN(n3817) );
  NAND3_X1 U4512 ( .A1(n4435), .A2(n3818), .A3(n3817), .ZN(n3821) );
  NAND2_X1 U4513 ( .A1(n4448), .A2(n4353), .ZN(n3820) );
  AOI22_X1 U4514 ( .A1(n4425), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3819) );
  NAND4_X1 U4515 ( .A1(n3822), .A2(n3821), .A3(n3820), .A4(n3819), .ZN(U3241)
         );
  AOI22_X1 U4516 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4425), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3832) );
  XNOR2_X1 U4517 ( .A(n3824), .B(n3823), .ZN(n3825) );
  NOR2_X1 U4518 ( .A1(n4444), .A2(n3825), .ZN(n3830) );
  AOI211_X1 U4519 ( .C1(n3828), .C2(n3827), .A(n3826), .B(n4440), .ZN(n3829)
         );
  AOI211_X1 U4520 ( .C1(n4448), .C2(n4352), .A(n3830), .B(n3829), .ZN(n3831)
         );
  NAND3_X1 U4521 ( .A1(n3833), .A2(n3832), .A3(n3831), .ZN(U3242) );
  INV_X1 U4522 ( .A(n4347), .ZN(n3856) );
  NAND2_X1 U4523 ( .A1(n4347), .A2(REG1_REG_15__SCAN_IN), .ZN(n3857) );
  OAI21_X1 U4524 ( .B1(n4347), .B2(REG1_REG_15__SCAN_IN), .A(n3857), .ZN(n3839) );
  NOR2_X1 U4525 ( .A1(n2080), .A2(n2192), .ZN(n3836) );
  INV_X1 U4526 ( .A(n3858), .ZN(n3837) );
  AOI21_X1 U4527 ( .B1(n3839), .B2(n3838), .A(n3837), .ZN(n3840) );
  NAND2_X1 U4528 ( .A1(n4435), .A2(n3840), .ZN(n3855) );
  NOR2_X1 U4529 ( .A1(n2192), .A2(n3844), .ZN(n3845) );
  NAND2_X1 U4530 ( .A1(n3856), .A2(REG2_REG_15__SCAN_IN), .ZN(n3848) );
  INV_X1 U4531 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3846) );
  NAND2_X1 U4532 ( .A1(n4347), .A2(n3846), .ZN(n3847) );
  AND2_X1 U4533 ( .A1(n3848), .A2(n3847), .ZN(n3850) );
  INV_X1 U4534 ( .A(n3867), .ZN(n3849) );
  AOI211_X1 U4535 ( .C1(n3851), .C2(n3850), .A(n3849), .B(n4440), .ZN(n3852)
         );
  AOI211_X1 U4536 ( .C1(n4425), .C2(ADDR_REG_15__SCAN_IN), .A(n3853), .B(n3852), .ZN(n3854) );
  OAI211_X1 U4537 ( .C1(n4438), .C2(n3856), .A(n3855), .B(n3854), .ZN(U3255)
         );
  INV_X1 U4538 ( .A(n3870), .ZN(n4466) );
  AOI22_X1 U4539 ( .A1(n3870), .A2(REG1_REG_17__SCAN_IN), .B1(n4254), .B2(
        n4466), .ZN(n4428) );
  NAND2_X1 U4540 ( .A1(n3859), .A2(n4468), .ZN(n3860) );
  NAND2_X1 U4541 ( .A1(n4417), .A2(n4416), .ZN(n4415) );
  NAND2_X1 U4542 ( .A1(n3860), .A2(n4415), .ZN(n4427) );
  NAND2_X1 U4543 ( .A1(n4428), .A2(n4427), .ZN(n4426) );
  NAND2_X1 U4544 ( .A1(n4447), .A2(REG1_REG_18__SCAN_IN), .ZN(n3862) );
  OR2_X1 U4545 ( .A1(n4447), .A2(REG1_REG_18__SCAN_IN), .ZN(n3861) );
  NAND2_X1 U4546 ( .A1(n3862), .A2(n3861), .ZN(n4445) );
  NAND2_X1 U4547 ( .A1(n4443), .A2(n3862), .ZN(n3864) );
  XNOR2_X1 U4548 ( .A(n3876), .B(REG1_REG_19__SCAN_IN), .ZN(n3863) );
  XNOR2_X1 U4549 ( .A(n3864), .B(n3863), .ZN(n3880) );
  NOR2_X1 U4550 ( .A1(n3870), .A2(REG2_REG_17__SCAN_IN), .ZN(n3865) );
  AOI21_X1 U4551 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3870), .A(n3865), .ZN(n4431) );
  NAND2_X1 U4552 ( .A1(n4347), .A2(REG2_REG_15__SCAN_IN), .ZN(n3866) );
  NAND2_X1 U4553 ( .A1(n3868), .A2(n4468), .ZN(n3869) );
  XNOR2_X1 U4554 ( .A(n4447), .B(REG2_REG_18__SCAN_IN), .ZN(n4441) );
  AOI21_X1 U4555 ( .B1(n4447), .B2(REG2_REG_18__SCAN_IN), .A(n4439), .ZN(n3873) );
  INV_X1 U4556 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3871) );
  MUX2_X1 U4557 ( .A(n3871), .B(REG2_REG_19__SCAN_IN), .S(n3876), .Z(n3872) );
  XNOR2_X1 U4558 ( .A(n3873), .B(n3872), .ZN(n3878) );
  NAND2_X1 U4559 ( .A1(n4425), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3874) );
  OAI211_X1 U4560 ( .C1(n4438), .C2(n3876), .A(n3875), .B(n3874), .ZN(n3877)
         );
  AOI21_X1 U4561 ( .B1(n3878), .B2(n4433), .A(n3877), .ZN(n3879) );
  OAI21_X1 U4562 ( .B1(n3880), .B2(n4444), .A(n3879), .ZN(U3259) );
  INV_X1 U4563 ( .A(n3881), .ZN(n3891) );
  INV_X1 U4564 ( .A(n3882), .ZN(n3884) );
  OAI21_X1 U4565 ( .B1(n3885), .B2(n3884), .A(n3883), .ZN(n3886) );
  XNOR2_X1 U4566 ( .A(n3886), .B(n3895), .ZN(n3890) );
  AOI21_X1 U4567 ( .B1(B_REG_SCAN_IN), .B2(n4367), .A(n4127), .ZN(n4196) );
  AOI22_X1 U4568 ( .A1(n3887), .A2(n4196), .B1(n4207), .B2(n3898), .ZN(n3889)
         );
  NAND2_X1 U4569 ( .A1(n3911), .A2(n4130), .ZN(n3888) );
  OAI211_X1 U4570 ( .C1(n3890), .C2(n4132), .A(n3889), .B(n3888), .ZN(n4211)
         );
  AOI21_X1 U4571 ( .B1(n3891), .B2(n4456), .A(n4211), .ZN(n3901) );
  AOI22_X1 U4572 ( .A1(n3894), .A2(n3893), .B1(n3892), .B2(n3911), .ZN(n3896)
         );
  XNOR2_X1 U4573 ( .A(n3896), .B(n3895), .ZN(n4210) );
  NAND2_X1 U4574 ( .A1(n4210), .A2(n3897), .ZN(n3900) );
  AOI22_X1 U4575 ( .A1(n4212), .A2(n4362), .B1(REG2_REG_29__SCAN_IN), .B2(
        n4361), .ZN(n3899) );
  OAI211_X1 U4576 ( .C1(n4361), .C2(n3901), .A(n3900), .B(n3899), .ZN(U3354)
         );
  NAND2_X1 U4577 ( .A1(n3904), .A2(n3903), .ZN(n3905) );
  XNOR2_X1 U4578 ( .A(n3905), .B(n3907), .ZN(n4218) );
  XOR2_X1 U4579 ( .A(n3907), .B(n3906), .Z(n3913) );
  OAI22_X1 U4580 ( .A1(n3909), .A2(n4176), .B1(n3908), .B2(n4198), .ZN(n3910)
         );
  AOI21_X1 U4581 ( .B1(n4173), .B2(n3911), .A(n3910), .ZN(n3912) );
  OAI21_X1 U4582 ( .B1(n3913), .B2(n4132), .A(n3912), .ZN(n4215) );
  AOI21_X1 U4583 ( .B1(n3915), .B2(n3931), .A(n3914), .ZN(n4216) );
  INV_X1 U4584 ( .A(n4216), .ZN(n3918) );
  AOI22_X1 U4585 ( .A1(n3916), .A2(n4456), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4361), .ZN(n3917) );
  OAI21_X1 U4586 ( .B1(n3918), .B2(n4138), .A(n3917), .ZN(n3919) );
  AOI21_X1 U4587 ( .B1(n4215), .B2(n4357), .A(n3919), .ZN(n3920) );
  OAI21_X1 U4588 ( .B1(n4218), .B2(n4141), .A(n3920), .ZN(U3263) );
  XNOR2_X1 U4589 ( .A(n3921), .B(n3925), .ZN(n4220) );
  INV_X1 U4590 ( .A(n4220), .ZN(n3938) );
  NAND2_X1 U4591 ( .A1(n3923), .A2(n3922), .ZN(n3924) );
  XOR2_X1 U4592 ( .A(n3925), .B(n3924), .Z(n3930) );
  AOI22_X1 U4593 ( .A1(n3964), .A2(n4130), .B1(n3926), .B2(n4207), .ZN(n3929)
         );
  NAND2_X1 U4594 ( .A1(n3927), .A2(n4173), .ZN(n3928) );
  OAI211_X1 U4595 ( .C1(n3930), .C2(n4132), .A(n3929), .B(n3928), .ZN(n4219)
         );
  INV_X1 U4596 ( .A(n3952), .ZN(n3933) );
  OAI21_X1 U4597 ( .B1(n3933), .B2(n3932), .A(n3931), .ZN(n4290) );
  AOI22_X1 U4598 ( .A1(n3934), .A2(n4456), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4361), .ZN(n3935) );
  OAI21_X1 U4599 ( .B1(n4290), .B2(n4138), .A(n3935), .ZN(n3936) );
  AOI21_X1 U4600 ( .B1(n4219), .B2(n4357), .A(n3936), .ZN(n3937) );
  OAI21_X1 U4601 ( .B1(n3938), .B2(n4141), .A(n3937), .ZN(U3264) );
  XNOR2_X1 U4602 ( .A(n3939), .B(n3943), .ZN(n4224) );
  INV_X1 U4603 ( .A(n4224), .ZN(n3957) );
  NAND2_X1 U4604 ( .A1(n3941), .A2(n3940), .ZN(n3942) );
  XOR2_X1 U4605 ( .A(n3943), .B(n3942), .Z(n3949) );
  OAI22_X1 U4606 ( .A1(n3945), .A2(n4176), .B1(n3944), .B2(n4198), .ZN(n3946)
         );
  AOI21_X1 U4607 ( .B1(n4173), .B2(n3947), .A(n3946), .ZN(n3948) );
  OAI21_X1 U4608 ( .B1(n3949), .B2(n4132), .A(n3948), .ZN(n4223) );
  NAND2_X1 U4609 ( .A1(n3967), .A2(n3950), .ZN(n3951) );
  NAND2_X1 U4610 ( .A1(n3952), .A2(n3951), .ZN(n4294) );
  AOI22_X1 U4611 ( .A1(n3953), .A2(n4456), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4361), .ZN(n3954) );
  OAI21_X1 U4612 ( .B1(n4294), .B2(n4138), .A(n3954), .ZN(n3955) );
  AOI21_X1 U4613 ( .B1(n4223), .B2(n4357), .A(n3955), .ZN(n3956) );
  OAI21_X1 U4614 ( .B1(n3957), .B2(n4141), .A(n3956), .ZN(U3265) );
  XOR2_X1 U4615 ( .A(n3961), .B(n3958), .Z(n4227) );
  INV_X1 U4616 ( .A(n4227), .ZN(n3973) );
  NAND2_X1 U4617 ( .A1(n3960), .A2(n3959), .ZN(n3962) );
  XNOR2_X1 U4618 ( .A(n3962), .B(n3961), .ZN(n3966) );
  OAI22_X1 U4619 ( .A1(n4706), .A2(n4176), .B1(n4198), .B2(n3968), .ZN(n3963)
         );
  AOI21_X1 U4620 ( .B1(n4173), .B2(n3964), .A(n3963), .ZN(n3965) );
  OAI21_X1 U4621 ( .B1(n3966), .B2(n4132), .A(n3965), .ZN(n4226) );
  OAI21_X1 U4622 ( .B1(n3989), .B2(n3968), .A(n3967), .ZN(n4298) );
  AOI22_X1 U4623 ( .A1(n4361), .A2(REG2_REG_24__SCAN_IN), .B1(n3969), .B2(
        n4456), .ZN(n3970) );
  OAI21_X1 U4624 ( .B1(n4298), .B2(n4138), .A(n3970), .ZN(n3971) );
  AOI21_X1 U4625 ( .B1(n4226), .B2(n4357), .A(n3971), .ZN(n3972) );
  OAI21_X1 U4626 ( .B1(n3973), .B2(n4141), .A(n3972), .ZN(U3266) );
  XNOR2_X1 U4627 ( .A(n3974), .B(n3980), .ZN(n4231) );
  INV_X1 U4628 ( .A(n4231), .ZN(n3995) );
  INV_X1 U4629 ( .A(n3975), .ZN(n3976) );
  AOI21_X1 U4630 ( .B1(n4014), .B2(n3977), .A(n3976), .ZN(n3999) );
  OAI21_X1 U4631 ( .B1(n3999), .B2(n3998), .A(n3979), .ZN(n3982) );
  INV_X1 U4632 ( .A(n3980), .ZN(n3981) );
  XNOR2_X1 U4633 ( .A(n3982), .B(n3981), .ZN(n3987) );
  OAI22_X1 U4634 ( .A1(n4015), .A2(n4176), .B1(n4198), .B2(n3983), .ZN(n3984)
         );
  AOI21_X1 U4635 ( .B1(n4173), .B2(n3985), .A(n3984), .ZN(n3986) );
  OAI21_X1 U4636 ( .B1(n3987), .B2(n4132), .A(n3986), .ZN(n4230) );
  AND2_X1 U4637 ( .A1(n2062), .A2(n3988), .ZN(n3990) );
  OR2_X1 U4638 ( .A1(n3990), .A2(n3989), .ZN(n4302) );
  AOI22_X1 U4639 ( .A1(n4361), .A2(REG2_REG_23__SCAN_IN), .B1(n3991), .B2(
        n4456), .ZN(n3992) );
  OAI21_X1 U4640 ( .B1(n4302), .B2(n4138), .A(n3992), .ZN(n3993) );
  AOI21_X1 U4641 ( .B1(n4230), .B2(n4357), .A(n3993), .ZN(n3994) );
  OAI21_X1 U4642 ( .B1(n3995), .B2(n4141), .A(n3994), .ZN(U3267) );
  OAI21_X1 U4643 ( .B1(n3997), .B2(n3998), .A(n3996), .ZN(n4236) );
  XNOR2_X1 U4644 ( .A(n3999), .B(n3998), .ZN(n4005) );
  NAND2_X1 U4645 ( .A1(n4000), .A2(n4173), .ZN(n4003) );
  AOI22_X1 U4646 ( .A1(n4001), .A2(n4130), .B1(n4007), .B2(n4207), .ZN(n4002)
         );
  NAND2_X1 U4647 ( .A1(n4003), .A2(n4002), .ZN(n4004) );
  AOI21_X1 U4648 ( .B1(n4005), .B2(n4179), .A(n4004), .ZN(n4235) );
  AOI22_X1 U4649 ( .A1(n4361), .A2(REG2_REG_22__SCAN_IN), .B1(n4006), .B2(
        n4456), .ZN(n4009) );
  NAND2_X1 U4650 ( .A1(n2073), .A2(n4007), .ZN(n4233) );
  NAND3_X1 U4651 ( .A1(n2062), .A2(n4362), .A3(n4233), .ZN(n4008) );
  OAI211_X1 U4652 ( .C1(n4235), .C2(n4361), .A(n4009), .B(n4008), .ZN(n4010)
         );
  INV_X1 U4653 ( .A(n4010), .ZN(n4011) );
  OAI21_X1 U4654 ( .B1(n4236), .B2(n4141), .A(n4011), .ZN(U3268) );
  XNOR2_X1 U4655 ( .A(n4012), .B(n4013), .ZN(n4238) );
  INV_X1 U4656 ( .A(n4238), .ZN(n4026) );
  XNOR2_X1 U4657 ( .A(n4014), .B(n4013), .ZN(n4018) );
  OAI22_X1 U4658 ( .A1(n4015), .A2(n4127), .B1(n4198), .B2(n4019), .ZN(n4016)
         );
  AOI21_X1 U4659 ( .B1(n4130), .B2(n4059), .A(n4016), .ZN(n4017) );
  OAI21_X1 U4660 ( .B1(n4018), .B2(n4132), .A(n4017), .ZN(n4237) );
  OAI21_X1 U4661 ( .B1(n4038), .B2(n4019), .A(n2073), .ZN(n4307) );
  NOR2_X1 U4662 ( .A1(n4307), .A2(n4138), .ZN(n4024) );
  INV_X1 U4663 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4022) );
  INV_X1 U4664 ( .A(n4020), .ZN(n4021) );
  OAI22_X1 U4665 ( .A1(n4357), .A2(n4022), .B1(n4021), .B2(n4187), .ZN(n4023)
         );
  AOI211_X1 U4666 ( .C1(n4237), .C2(n4357), .A(n4024), .B(n4023), .ZN(n4025)
         );
  OAI21_X1 U4667 ( .B1(n4026), .B2(n4141), .A(n4025), .ZN(U3269) );
  XNOR2_X1 U4668 ( .A(n4027), .B(n4030), .ZN(n4240) );
  NAND2_X1 U4669 ( .A1(n4029), .A2(n4028), .ZN(n4031) );
  XNOR2_X1 U4670 ( .A(n4031), .B(n4030), .ZN(n4036) );
  AOI22_X1 U4671 ( .A1(n2099), .A2(n4130), .B1(n4032), .B2(n4207), .ZN(n4033)
         );
  OAI21_X1 U4672 ( .B1(n4034), .B2(n4127), .A(n4033), .ZN(n4035) );
  AOI21_X1 U4673 ( .B1(n4036), .B2(n4179), .A(n4035), .ZN(n4037) );
  OAI21_X1 U4674 ( .B1(n4240), .B2(n4182), .A(n4037), .ZN(n4241) );
  NAND2_X1 U4675 ( .A1(n4241), .A2(n4357), .ZN(n4047) );
  INV_X1 U4676 ( .A(n4038), .ZN(n4039) );
  OAI21_X1 U4677 ( .B1(n4062), .B2(n4040), .A(n4039), .ZN(n4311) );
  INV_X1 U4678 ( .A(n4311), .ZN(n4045) );
  INV_X1 U4679 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4043) );
  INV_X1 U4680 ( .A(n4041), .ZN(n4042) );
  OAI22_X1 U4681 ( .A1(n4357), .A2(n4043), .B1(n4042), .B2(n4187), .ZN(n4044)
         );
  AOI21_X1 U4682 ( .B1(n4045), .B2(n4362), .A(n4044), .ZN(n4046) );
  OAI211_X1 U4683 ( .C1(n4240), .C2(n4194), .A(n4047), .B(n4046), .ZN(U3270)
         );
  XNOR2_X1 U4684 ( .A(n4049), .B(n4048), .ZN(n4246) );
  INV_X1 U4685 ( .A(n4246), .ZN(n4070) );
  INV_X1 U4686 ( .A(n4050), .ZN(n4052) );
  OAI21_X1 U4687 ( .B1(n4090), .B2(n4052), .A(n4051), .ZN(n4073) );
  INV_X1 U4688 ( .A(n4053), .ZN(n4055) );
  OAI21_X1 U4689 ( .B1(n4073), .B2(n4055), .A(n4054), .ZN(n4057) );
  XNOR2_X1 U4690 ( .A(n4057), .B(n4056), .ZN(n4061) );
  OAI22_X1 U4691 ( .A1(n4093), .A2(n4176), .B1(n4064), .B2(n4198), .ZN(n4058)
         );
  AOI21_X1 U4692 ( .B1(n4173), .B2(n4059), .A(n4058), .ZN(n4060) );
  OAI21_X1 U4693 ( .B1(n4061), .B2(n4132), .A(n4060), .ZN(n4245) );
  INV_X1 U4694 ( .A(n4080), .ZN(n4065) );
  INV_X1 U4695 ( .A(n4062), .ZN(n4063) );
  OAI21_X1 U4696 ( .B1(n4065), .B2(n4064), .A(n4063), .ZN(n4315) );
  AOI22_X1 U4697 ( .A1(n4361), .A2(REG2_REG_19__SCAN_IN), .B1(n4066), .B2(
        n4456), .ZN(n4067) );
  OAI21_X1 U4698 ( .B1(n4315), .B2(n4138), .A(n4067), .ZN(n4068) );
  AOI21_X1 U4699 ( .B1(n4245), .B2(n4357), .A(n4068), .ZN(n4069) );
  OAI21_X1 U4700 ( .B1(n4070), .B2(n4141), .A(n4069), .ZN(U3271) );
  AOI21_X1 U4701 ( .B1(n4072), .B2(n4071), .A(n2093), .ZN(n4251) );
  XNOR2_X1 U4702 ( .A(n4073), .B(n4072), .ZN(n4078) );
  AOI22_X1 U4703 ( .A1(n2099), .A2(n4173), .B1(n4207), .B2(n4079), .ZN(n4075)
         );
  OAI21_X1 U4704 ( .B1(n4076), .B2(n4176), .A(n4075), .ZN(n4077) );
  AOI21_X1 U4705 ( .B1(n4078), .B2(n4179), .A(n4077), .ZN(n4250) );
  INV_X1 U4706 ( .A(n4250), .ZN(n4087) );
  AOI21_X1 U4707 ( .B1(n4100), .B2(n4079), .A(n4506), .ZN(n4081) );
  NAND2_X1 U4708 ( .A1(n4081), .A2(n4080), .ZN(n4249) );
  INV_X1 U4709 ( .A(n4082), .ZN(n4085) );
  AOI22_X1 U4710 ( .A1(n4361), .A2(REG2_REG_18__SCAN_IN), .B1(n4083), .B2(
        n4456), .ZN(n4084) );
  OAI21_X1 U4711 ( .B1(n4249), .B2(n4085), .A(n4084), .ZN(n4086) );
  AOI21_X1 U4712 ( .B1(n4087), .B2(n4357), .A(n4086), .ZN(n4088) );
  OAI21_X1 U4713 ( .B1(n4251), .B2(n4141), .A(n4088), .ZN(U3272) );
  XOR2_X1 U4714 ( .A(n4091), .B(n4089), .Z(n4253) );
  INV_X1 U4715 ( .A(n4253), .ZN(n4105) );
  XOR2_X1 U4716 ( .A(n4091), .B(n4090), .Z(n4097) );
  OAI22_X1 U4717 ( .A1(n4093), .A2(n4127), .B1(n4092), .B2(n4198), .ZN(n4094)
         );
  AOI21_X1 U4718 ( .B1(n4130), .B2(n4095), .A(n4094), .ZN(n4096) );
  OAI21_X1 U4719 ( .B1(n4097), .B2(n4132), .A(n4096), .ZN(n4252) );
  NAND2_X1 U4720 ( .A1(n4256), .A2(n4098), .ZN(n4099) );
  NAND2_X1 U4721 ( .A1(n4100), .A2(n4099), .ZN(n4320) );
  AOI22_X1 U4722 ( .A1(n4361), .A2(REG2_REG_17__SCAN_IN), .B1(n4101), .B2(
        n4456), .ZN(n4102) );
  OAI21_X1 U4723 ( .B1(n4320), .B2(n4138), .A(n4102), .ZN(n4103) );
  AOI21_X1 U4724 ( .B1(n4252), .B2(n4357), .A(n4103), .ZN(n4104) );
  OAI21_X1 U4725 ( .B1(n4105), .B2(n4141), .A(n4104), .ZN(U3273) );
  OAI21_X1 U4726 ( .B1(n4107), .B2(n4108), .A(n4106), .ZN(n4260) );
  XNOR2_X1 U4727 ( .A(n4109), .B(n4108), .ZN(n4114) );
  NAND2_X1 U4728 ( .A1(n4149), .A2(n4130), .ZN(n4112) );
  NAND2_X1 U4729 ( .A1(n4110), .A2(n4173), .ZN(n4111) );
  OAI211_X1 U4730 ( .C1(n4198), .C2(n4118), .A(n4112), .B(n4111), .ZN(n4113)
         );
  AOI21_X1 U4731 ( .B1(n4114), .B2(n4179), .A(n4113), .ZN(n4259) );
  OAI22_X1 U4732 ( .A1(n4357), .A2(n4116), .B1(n4115), .B2(n4187), .ZN(n4117)
         );
  INV_X1 U4733 ( .A(n4117), .ZN(n4120) );
  OR2_X1 U4734 ( .A1(n4134), .A2(n4118), .ZN(n4257) );
  NAND3_X1 U4735 ( .A1(n4256), .A2(n4257), .A3(n4362), .ZN(n4119) );
  OAI211_X1 U4736 ( .C1(n4259), .C2(n4361), .A(n4120), .B(n4119), .ZN(n4121)
         );
  INV_X1 U4737 ( .A(n4121), .ZN(n4122) );
  OAI21_X1 U4738 ( .B1(n4260), .B2(n4141), .A(n4122), .ZN(U3274) );
  XNOR2_X1 U4739 ( .A(n4123), .B(n4125), .ZN(n4262) );
  INV_X1 U4740 ( .A(n4262), .ZN(n4142) );
  NAND2_X1 U4741 ( .A1(n4146), .A2(n4124), .ZN(n4126) );
  XNOR2_X1 U4742 ( .A(n4126), .B(n4125), .ZN(n4133) );
  OAI22_X1 U4743 ( .A1(n4128), .A2(n4127), .B1(n4198), .B2(n2100), .ZN(n4129)
         );
  AOI21_X1 U4744 ( .B1(n4130), .B2(n4174), .A(n4129), .ZN(n4131) );
  OAI21_X1 U4745 ( .B1(n4133), .B2(n4132), .A(n4131), .ZN(n4261) );
  INV_X1 U4746 ( .A(n4157), .ZN(n4135) );
  OAI21_X1 U4747 ( .B1(n4135), .B2(n2100), .A(n2101), .ZN(n4325) );
  AOI22_X1 U4748 ( .A1(n4361), .A2(REG2_REG_15__SCAN_IN), .B1(n4136), .B2(
        n4456), .ZN(n4137) );
  OAI21_X1 U4749 ( .B1(n4325), .B2(n4138), .A(n4137), .ZN(n4139) );
  AOI21_X1 U4750 ( .B1(n4261), .B2(n4357), .A(n4139), .ZN(n4140) );
  OAI21_X1 U4751 ( .B1(n4142), .B2(n4141), .A(n4140), .ZN(U3275) );
  OAI21_X1 U4752 ( .B1(n4145), .B2(n4144), .A(n4143), .ZN(n4266) );
  INV_X1 U4753 ( .A(n4266), .ZN(n4164) );
  OAI21_X1 U4754 ( .B1(n4148), .B2(n4147), .A(n4146), .ZN(n4153) );
  AOI22_X1 U4755 ( .A1(n4149), .A2(n4173), .B1(n4207), .B2(n4155), .ZN(n4150)
         );
  OAI21_X1 U4756 ( .B1(n4151), .B2(n4176), .A(n4150), .ZN(n4152) );
  AOI21_X1 U4757 ( .B1(n4153), .B2(n4179), .A(n4152), .ZN(n4154) );
  OAI21_X1 U4758 ( .B1(n4164), .B2(n4182), .A(n4154), .ZN(n4265) );
  NAND2_X1 U4759 ( .A1(n4265), .A2(n4357), .ZN(n4163) );
  NAND2_X1 U4760 ( .A1(n4186), .A2(n4155), .ZN(n4156) );
  NAND2_X1 U4761 ( .A1(n4157), .A2(n4156), .ZN(n4329) );
  INV_X1 U4762 ( .A(n4329), .ZN(n4161) );
  OAI22_X1 U4763 ( .A1(n4357), .A2(n4159), .B1(n4158), .B2(n4187), .ZN(n4160)
         );
  AOI21_X1 U4764 ( .B1(n4161), .B2(n4362), .A(n4160), .ZN(n4162) );
  OAI211_X1 U4765 ( .C1(n4164), .C2(n4194), .A(n4163), .B(n4162), .ZN(U3276)
         );
  XNOR2_X1 U4766 ( .A(n4165), .B(n4170), .ZN(n4268) );
  INV_X1 U4767 ( .A(n4166), .ZN(n4167) );
  AOI21_X1 U4768 ( .B1(n4169), .B2(n4168), .A(n4167), .ZN(n4171) );
  XNOR2_X1 U4769 ( .A(n4171), .B(n4170), .ZN(n4180) );
  AOI22_X1 U4770 ( .A1(n4174), .A2(n4173), .B1(n4207), .B2(n4172), .ZN(n4175)
         );
  OAI21_X1 U4771 ( .B1(n4177), .B2(n4176), .A(n4175), .ZN(n4178) );
  AOI21_X1 U4772 ( .B1(n4180), .B2(n4179), .A(n4178), .ZN(n4181) );
  OAI21_X1 U4773 ( .B1(n4268), .B2(n4182), .A(n4181), .ZN(n4269) );
  NAND2_X1 U4774 ( .A1(n4269), .A2(n4357), .ZN(n4193) );
  OR2_X1 U4775 ( .A1(n4184), .A2(n4183), .ZN(n4185) );
  NAND2_X1 U4776 ( .A1(n4186), .A2(n4185), .ZN(n4333) );
  INV_X1 U4777 ( .A(n4333), .ZN(n4191) );
  OAI22_X1 U4778 ( .A1(n4357), .A2(n4189), .B1(n4188), .B2(n4187), .ZN(n4190)
         );
  AOI21_X1 U4779 ( .B1(n4191), .B2(n4362), .A(n4190), .ZN(n4192) );
  OAI211_X1 U4780 ( .C1(n4268), .C2(n4194), .A(n4193), .B(n4192), .ZN(U3277)
         );
  NAND2_X1 U4781 ( .A1(n4204), .A2(n4203), .ZN(n4202) );
  XNOR2_X1 U4782 ( .A(n4202), .B(n4199), .ZN(n4358) );
  NAND2_X1 U4783 ( .A1(n4358), .A2(n4195), .ZN(n4201) );
  NAND2_X1 U4784 ( .A1(n4197), .A2(n4196), .ZN(n4205) );
  OAI21_X1 U4785 ( .B1(n4199), .B2(n4198), .A(n4205), .ZN(n4356) );
  NAND2_X1 U4786 ( .A1(n4519), .A2(n4356), .ZN(n4200) );
  OAI211_X1 U4787 ( .C1(n4519), .C2(n3707), .A(n4201), .B(n4200), .ZN(U3549)
         );
  OAI21_X1 U4788 ( .B1(n4204), .B2(n4203), .A(n4202), .ZN(n4360) );
  INV_X1 U4789 ( .A(n4205), .ZN(n4206) );
  AOI21_X1 U4790 ( .B1(n4208), .B2(n4207), .A(n4206), .ZN(n4365) );
  MUX2_X1 U4791 ( .A(n3702), .B(n4365), .S(n4519), .Z(n4209) );
  OAI21_X1 U4792 ( .B1(n4360), .B2(n4281), .A(n4209), .ZN(U3548) );
  NAND2_X1 U4793 ( .A1(n4210), .A2(n4508), .ZN(n4214) );
  AOI21_X1 U4794 ( .B1(n4496), .B2(n4212), .A(n4211), .ZN(n4213) );
  NAND2_X1 U4795 ( .A1(n4214), .A2(n4213), .ZN(n4286) );
  MUX2_X1 U4796 ( .A(REG1_REG_29__SCAN_IN), .B(n4286), .S(n4519), .Z(U3547) );
  AOI21_X1 U4797 ( .B1(n4496), .B2(n4216), .A(n4215), .ZN(n4217) );
  OAI21_X1 U4798 ( .B1(n4218), .B2(n4499), .A(n4217), .ZN(n4287) );
  MUX2_X1 U4799 ( .A(REG1_REG_27__SCAN_IN), .B(n4287), .S(n4519), .Z(U3545) );
  INV_X1 U4800 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4221) );
  AOI21_X1 U4801 ( .B1(n4220), .B2(n4508), .A(n4219), .ZN(n4288) );
  MUX2_X1 U4802 ( .A(n4221), .B(n4288), .S(n4519), .Z(n4222) );
  OAI21_X1 U4803 ( .B1(n4281), .B2(n4290), .A(n4222), .ZN(U3544) );
  AOI21_X1 U4804 ( .B1(n4224), .B2(n4508), .A(n4223), .ZN(n4291) );
  MUX2_X1 U4805 ( .A(n4671), .B(n4291), .S(n4519), .Z(n4225) );
  OAI21_X1 U4806 ( .B1(n4281), .B2(n4294), .A(n4225), .ZN(U3543) );
  AOI21_X1 U4807 ( .B1(n4227), .B2(n4508), .A(n4226), .ZN(n4295) );
  MUX2_X1 U4808 ( .A(n4228), .B(n4295), .S(n4519), .Z(n4229) );
  OAI21_X1 U4809 ( .B1(n4281), .B2(n4298), .A(n4229), .ZN(U3542) );
  AOI21_X1 U4810 ( .B1(n4231), .B2(n4508), .A(n4230), .ZN(n4299) );
  MUX2_X1 U4811 ( .A(n4662), .B(n4299), .S(n4519), .Z(n4232) );
  OAI21_X1 U4812 ( .B1(n4281), .B2(n4302), .A(n4232), .ZN(U3541) );
  NAND3_X1 U4813 ( .A1(n2062), .A2(n4496), .A3(n4233), .ZN(n4234) );
  OAI211_X1 U4814 ( .C1(n4236), .C2(n4499), .A(n4235), .B(n4234), .ZN(n4303)
         );
  MUX2_X1 U4815 ( .A(REG1_REG_22__SCAN_IN), .B(n4303), .S(n4519), .Z(U3540) );
  AOI21_X1 U4816 ( .B1(n4238), .B2(n4508), .A(n4237), .ZN(n4304) );
  MUX2_X1 U4817 ( .A(n4672), .B(n4304), .S(n4519), .Z(n4239) );
  OAI21_X1 U4818 ( .B1(n4281), .B2(n4307), .A(n4239), .ZN(U3539) );
  INV_X1 U4819 ( .A(n4240), .ZN(n4242) );
  AOI21_X1 U4820 ( .B1(n4489), .B2(n4242), .A(n4241), .ZN(n4308) );
  MUX2_X1 U4821 ( .A(n4243), .B(n4308), .S(n4519), .Z(n4244) );
  OAI21_X1 U4822 ( .B1(n4281), .B2(n4311), .A(n4244), .ZN(U3538) );
  AOI21_X1 U4823 ( .B1(n4246), .B2(n4508), .A(n4245), .ZN(n4312) );
  MUX2_X1 U4824 ( .A(n4247), .B(n4312), .S(n4519), .Z(n4248) );
  OAI21_X1 U4825 ( .B1(n4281), .B2(n4315), .A(n4248), .ZN(U3537) );
  OAI211_X1 U4826 ( .C1(n4251), .C2(n4499), .A(n4250), .B(n4249), .ZN(n4316)
         );
  MUX2_X1 U4827 ( .A(REG1_REG_18__SCAN_IN), .B(n4316), .S(n4519), .Z(U3536) );
  AOI21_X1 U4828 ( .B1(n4253), .B2(n4508), .A(n4252), .ZN(n4317) );
  MUX2_X1 U4829 ( .A(n4254), .B(n4317), .S(n4519), .Z(n4255) );
  OAI21_X1 U4830 ( .B1(n4281), .B2(n4320), .A(n4255), .ZN(U3535) );
  NAND3_X1 U4831 ( .A1(n4257), .A2(n4496), .A3(n4256), .ZN(n4258) );
  OAI211_X1 U4832 ( .C1(n4260), .C2(n4499), .A(n4259), .B(n4258), .ZN(n4321)
         );
  MUX2_X1 U4833 ( .A(REG1_REG_16__SCAN_IN), .B(n4321), .S(n4519), .Z(U3534) );
  AOI21_X1 U4834 ( .B1(n4262), .B2(n4508), .A(n4261), .ZN(n4322) );
  MUX2_X1 U4835 ( .A(n4263), .B(n4322), .S(n4519), .Z(n4264) );
  OAI21_X1 U4836 ( .B1(n4281), .B2(n4325), .A(n4264), .ZN(U3533) );
  AOI21_X1 U4837 ( .B1(n4489), .B2(n4266), .A(n4265), .ZN(n4326) );
  MUX2_X1 U4838 ( .A(n4405), .B(n4326), .S(n4519), .Z(n4267) );
  OAI21_X1 U4839 ( .B1(n4281), .B2(n4329), .A(n4267), .ZN(U3532) );
  INV_X1 U4840 ( .A(n4268), .ZN(n4270) );
  AOI21_X1 U4841 ( .B1(n4489), .B2(n4270), .A(n4269), .ZN(n4330) );
  MUX2_X1 U4842 ( .A(n4271), .B(n4330), .S(n4519), .Z(n4272) );
  OAI21_X1 U4843 ( .B1(n4281), .B2(n4333), .A(n4272), .ZN(U3531) );
  AOI21_X1 U4844 ( .B1(n4274), .B2(n4508), .A(n4273), .ZN(n4334) );
  MUX2_X1 U4845 ( .A(n4536), .B(n4334), .S(n4519), .Z(n4275) );
  OAI21_X1 U4846 ( .B1(n4281), .B2(n4337), .A(n4275), .ZN(U3530) );
  INV_X1 U4847 ( .A(n4276), .ZN(n4277) );
  AOI21_X1 U4848 ( .B1(n4489), .B2(n4278), .A(n4277), .ZN(n4338) );
  MUX2_X1 U4849 ( .A(n4279), .B(n4338), .S(n4519), .Z(n4280) );
  OAI21_X1 U4850 ( .B1(n4281), .B2(n4342), .A(n4280), .ZN(U3529) );
  INV_X1 U4851 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4545) );
  NAND2_X1 U4852 ( .A1(n4358), .A2(n4282), .ZN(n4284) );
  NAND2_X1 U4853 ( .A1(n4511), .A2(n4356), .ZN(n4283) );
  OAI211_X1 U4854 ( .C1(n4511), .C2(n4545), .A(n4284), .B(n4283), .ZN(U3517)
         );
  INV_X1 U4855 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4645) );
  MUX2_X1 U4856 ( .A(n4645), .B(n4365), .S(n4511), .Z(n4285) );
  OAI21_X1 U4857 ( .B1(n4360), .B2(n4341), .A(n4285), .ZN(U3516) );
  MUX2_X1 U4858 ( .A(REG0_REG_29__SCAN_IN), .B(n4286), .S(n4511), .Z(U3515) );
  MUX2_X1 U4859 ( .A(REG0_REG_27__SCAN_IN), .B(n4287), .S(n4511), .Z(U3513) );
  MUX2_X1 U4860 ( .A(n4680), .B(n4288), .S(n4511), .Z(n4289) );
  OAI21_X1 U4861 ( .B1(n4290), .B2(n4341), .A(n4289), .ZN(U3512) );
  INV_X1 U4862 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4292) );
  MUX2_X1 U4863 ( .A(n4292), .B(n4291), .S(n4511), .Z(n4293) );
  OAI21_X1 U4864 ( .B1(n4294), .B2(n4341), .A(n4293), .ZN(U3511) );
  INV_X1 U4865 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4296) );
  MUX2_X1 U4866 ( .A(n4296), .B(n4295), .S(n4511), .Z(n4297) );
  OAI21_X1 U4867 ( .B1(n4298), .B2(n4341), .A(n4297), .ZN(U3510) );
  INV_X1 U4868 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4300) );
  MUX2_X1 U4869 ( .A(n4300), .B(n4299), .S(n4511), .Z(n4301) );
  OAI21_X1 U4870 ( .B1(n4302), .B2(n4341), .A(n4301), .ZN(U3509) );
  MUX2_X1 U4871 ( .A(REG0_REG_22__SCAN_IN), .B(n4303), .S(n4511), .Z(U3508) );
  INV_X1 U4872 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4305) );
  MUX2_X1 U4873 ( .A(n4305), .B(n4304), .S(n4511), .Z(n4306) );
  OAI21_X1 U4874 ( .B1(n4307), .B2(n4341), .A(n4306), .ZN(U3507) );
  INV_X1 U4875 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4309) );
  MUX2_X1 U4876 ( .A(n4309), .B(n4308), .S(n4511), .Z(n4310) );
  OAI21_X1 U4877 ( .B1(n4311), .B2(n4341), .A(n4310), .ZN(U3506) );
  INV_X1 U4878 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4313) );
  MUX2_X1 U4879 ( .A(n4313), .B(n4312), .S(n4511), .Z(n4314) );
  OAI21_X1 U4880 ( .B1(n4315), .B2(n4341), .A(n4314), .ZN(U3505) );
  MUX2_X1 U4881 ( .A(REG0_REG_18__SCAN_IN), .B(n4316), .S(n4511), .Z(U3503) );
  MUX2_X1 U4882 ( .A(n4318), .B(n4317), .S(n4511), .Z(n4319) );
  OAI21_X1 U4883 ( .B1(n4320), .B2(n4341), .A(n4319), .ZN(U3501) );
  MUX2_X1 U4884 ( .A(REG0_REG_16__SCAN_IN), .B(n4321), .S(n4511), .Z(U3499) );
  MUX2_X1 U4885 ( .A(n4323), .B(n4322), .S(n4511), .Z(n4324) );
  OAI21_X1 U4886 ( .B1(n4325), .B2(n4341), .A(n4324), .ZN(U3497) );
  INV_X1 U4887 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4327) );
  MUX2_X1 U4888 ( .A(n4327), .B(n4326), .S(n4511), .Z(n4328) );
  OAI21_X1 U4889 ( .B1(n4329), .B2(n4341), .A(n4328), .ZN(U3495) );
  INV_X1 U4890 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4331) );
  MUX2_X1 U4891 ( .A(n4331), .B(n4330), .S(n4511), .Z(n4332) );
  OAI21_X1 U4892 ( .B1(n4333), .B2(n4341), .A(n4332), .ZN(U3493) );
  MUX2_X1 U4893 ( .A(n4335), .B(n4334), .S(n4511), .Z(n4336) );
  OAI21_X1 U4894 ( .B1(n4337), .B2(n4341), .A(n4336), .ZN(U3491) );
  INV_X1 U4895 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4339) );
  MUX2_X1 U4896 ( .A(n4339), .B(n4338), .S(n4511), .Z(n4340) );
  OAI21_X1 U4897 ( .B1(n4342), .B2(n4341), .A(n4340), .ZN(U3489) );
  MUX2_X1 U4898 ( .A(DATAI_30_), .B(n4343), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4899 ( .A(DATAI_29_), .B(n4344), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U4900 ( .A(DATAI_27_), .B(n4367), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U4901 ( .A(n4345), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U4902 ( .A(DATAI_20_), .B(n4346), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4903 ( .A(DATAI_18_), .B(n4447), .S(STATE_REG_SCAN_IN), .Z(U3334)
         );
  MUX2_X1 U4904 ( .A(n4347), .B(DATAI_15_), .S(U3149), .Z(U3337) );
  MUX2_X1 U4905 ( .A(DATAI_8_), .B(n4348), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U4906 ( .A(n4349), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4907 ( .A(DATAI_5_), .B(n4350), .S(STATE_REG_SCAN_IN), .Z(U3347) );
  MUX2_X1 U4908 ( .A(n4351), .B(DATAI_4_), .S(U3149), .Z(U3348) );
  MUX2_X1 U4909 ( .A(n4352), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4910 ( .A(n4353), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  OAI22_X1 U4911 ( .A1(U3149), .A2(n4354), .B1(DATAI_28_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4355) );
  INV_X1 U4912 ( .A(n4355), .ZN(U3324) );
  AOI22_X1 U4913 ( .A1(n4358), .A2(n4362), .B1(n4357), .B2(n4356), .ZN(n4359)
         );
  OAI21_X1 U4914 ( .B1(n4357), .B2(n3703), .A(n4359), .ZN(U3260) );
  INV_X1 U4915 ( .A(n4360), .ZN(n4363) );
  AOI22_X1 U4916 ( .A1(n4363), .A2(n4362), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4361), .ZN(n4364) );
  OAI21_X1 U4917 ( .B1(n4361), .B2(n4365), .A(n4364), .ZN(U3261) );
  INV_X1 U4918 ( .A(n4369), .ZN(n4366) );
  OAI211_X1 U4919 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4367), .A(n4366), .B(n4368), 
        .ZN(n4373) );
  OAI22_X1 U4920 ( .A1(n4369), .A2(n4368), .B1(n4444), .B2(REG1_REG_0__SCAN_IN), .ZN(n4370) );
  INV_X1 U4921 ( .A(n4370), .ZN(n4372) );
  AOI22_X1 U4922 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4425), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4371) );
  OAI221_X1 U4923 ( .B1(IR_REG_0__SCAN_IN), .B2(n4373), .C1(n4525), .C2(n4372), 
        .A(n4371), .ZN(U3240) );
  AOI211_X1 U4924 ( .C1(n4376), .C2(n4375), .A(n4374), .B(n4444), .ZN(n4378)
         );
  AOI211_X1 U4925 ( .C1(n4425), .C2(ADDR_REG_10__SCAN_IN), .A(n4378), .B(n4377), .ZN(n4382) );
  OAI211_X1 U4926 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4380), .A(n4433), .B(n4379), .ZN(n4381) );
  OAI211_X1 U4927 ( .C1(n4438), .C2(n4383), .A(n4382), .B(n4381), .ZN(U3250)
         );
  AOI211_X1 U4928 ( .C1(n4386), .C2(n4385), .A(n4384), .B(n4444), .ZN(n4388)
         );
  AOI211_X1 U4929 ( .C1(n4425), .C2(ADDR_REG_11__SCAN_IN), .A(n4388), .B(n4387), .ZN(n4393) );
  OAI211_X1 U4930 ( .C1(n4391), .C2(n4390), .A(n4433), .B(n4389), .ZN(n4392)
         );
  OAI211_X1 U4931 ( .C1(n4438), .C2(n4394), .A(n4393), .B(n4392), .ZN(U3251)
         );
  AOI211_X1 U4932 ( .C1(n4536), .C2(n4396), .A(n4395), .B(n4444), .ZN(n4398)
         );
  AOI211_X1 U4933 ( .C1(n4425), .C2(ADDR_REG_12__SCAN_IN), .A(n4398), .B(n4397), .ZN(n4402) );
  OAI211_X1 U4934 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4400), .A(n4433), .B(n4399), .ZN(n4401) );
  OAI211_X1 U4935 ( .C1(n4438), .C2(n4469), .A(n4402), .B(n4401), .ZN(U3252)
         );
  NAND2_X1 U4936 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4425), .ZN(n4413) );
  AOI211_X1 U4937 ( .C1(n4405), .C2(n4404), .A(n4403), .B(n4444), .ZN(n4409)
         );
  AOI211_X1 U4938 ( .C1(n4159), .C2(n4407), .A(n4406), .B(n4440), .ZN(n4408)
         );
  AOI211_X1 U4939 ( .C1(n4448), .C2(n4410), .A(n4409), .B(n4408), .ZN(n4412)
         );
  NAND3_X1 U4940 ( .A1(n4413), .A2(n4412), .A3(n4411), .ZN(U3254) );
  AOI21_X1 U4941 ( .B1(n4425), .B2(ADDR_REG_16__SCAN_IN), .A(n4414), .ZN(n4423) );
  OAI21_X1 U4942 ( .B1(n4417), .B2(n4416), .A(n4415), .ZN(n4421) );
  OAI21_X1 U4943 ( .B1(n4419), .B2(n4116), .A(n4418), .ZN(n4420) );
  AOI22_X1 U4944 ( .A1(n4435), .A2(n4421), .B1(n4433), .B2(n4420), .ZN(n4422)
         );
  OAI211_X1 U4945 ( .C1(n4468), .C2(n4438), .A(n4423), .B(n4422), .ZN(U3256)
         );
  AOI21_X1 U4946 ( .B1(n4425), .B2(ADDR_REG_17__SCAN_IN), .A(n4424), .ZN(n4437) );
  OAI21_X1 U4947 ( .B1(n4428), .B2(n4427), .A(n4426), .ZN(n4434) );
  OAI21_X1 U4948 ( .B1(n4431), .B2(n4430), .A(n4429), .ZN(n4432) );
  AOI22_X1 U4949 ( .A1(n4435), .A2(n4434), .B1(n4433), .B2(n4432), .ZN(n4436)
         );
  OAI211_X1 U4950 ( .C1(n4466), .C2(n4438), .A(n4437), .B(n4436), .ZN(U3257)
         );
  INV_X1 U4951 ( .A(ADDR_REG_18__SCAN_IN), .ZN(n4450) );
  INV_X1 U4952 ( .A(n4452), .ZN(n4454) );
  AOI21_X1 U4953 ( .B1(n4455), .B2(n4454), .A(n4453), .ZN(n4461) );
  AOI22_X1 U4954 ( .A1(n4458), .A2(n4457), .B1(REG3_REG_0__SCAN_IN), .B2(n4456), .ZN(n4459) );
  OAI221_X1 U4955 ( .B1(n4361), .B2(n4461), .C1(n4357), .C2(n4460), .A(n4459), 
        .ZN(U3290) );
  AND2_X1 U4956 ( .A1(D_REG_31__SCAN_IN), .A2(n4462), .ZN(U3291) );
  AND2_X1 U4957 ( .A1(D_REG_30__SCAN_IN), .A2(n4462), .ZN(U3292) );
  INV_X1 U4958 ( .A(D_REG_29__SCAN_IN), .ZN(n4689) );
  NOR2_X1 U4959 ( .A1(n4463), .A2(n4689), .ZN(U3293) );
  INV_X1 U4960 ( .A(D_REG_28__SCAN_IN), .ZN(n4688) );
  NOR2_X1 U4961 ( .A1(n4463), .A2(n4688), .ZN(U3294) );
  AND2_X1 U4962 ( .A1(D_REG_27__SCAN_IN), .A2(n4462), .ZN(U3295) );
  AND2_X1 U4963 ( .A1(D_REG_26__SCAN_IN), .A2(n4462), .ZN(U3296) );
  INV_X1 U4964 ( .A(D_REG_25__SCAN_IN), .ZN(n4686) );
  NOR2_X1 U4965 ( .A1(n4463), .A2(n4686), .ZN(U3297) );
  AND2_X1 U4966 ( .A1(D_REG_24__SCAN_IN), .A2(n4462), .ZN(U3298) );
  AND2_X1 U4967 ( .A1(D_REG_23__SCAN_IN), .A2(n4462), .ZN(U3299) );
  AND2_X1 U4968 ( .A1(D_REG_22__SCAN_IN), .A2(n4462), .ZN(U3300) );
  AND2_X1 U4969 ( .A1(D_REG_21__SCAN_IN), .A2(n4462), .ZN(U3301) );
  AND2_X1 U4970 ( .A1(D_REG_20__SCAN_IN), .A2(n4462), .ZN(U3302) );
  AND2_X1 U4971 ( .A1(D_REG_19__SCAN_IN), .A2(n4462), .ZN(U3303) );
  AND2_X1 U4972 ( .A1(D_REG_18__SCAN_IN), .A2(n4462), .ZN(U3304) );
  INV_X1 U4973 ( .A(D_REG_17__SCAN_IN), .ZN(n4693) );
  NOR2_X1 U4974 ( .A1(n4463), .A2(n4693), .ZN(U3305) );
  INV_X1 U4975 ( .A(D_REG_16__SCAN_IN), .ZN(n4646) );
  NOR2_X1 U4976 ( .A1(n4463), .A2(n4646), .ZN(U3306) );
  AND2_X1 U4977 ( .A1(D_REG_15__SCAN_IN), .A2(n4462), .ZN(U3307) );
  AND2_X1 U4978 ( .A1(D_REG_14__SCAN_IN), .A2(n4462), .ZN(U3308) );
  AND2_X1 U4979 ( .A1(D_REG_13__SCAN_IN), .A2(n4462), .ZN(U3309) );
  AND2_X1 U4980 ( .A1(D_REG_12__SCAN_IN), .A2(n4462), .ZN(U3310) );
  AND2_X1 U4981 ( .A1(D_REG_11__SCAN_IN), .A2(n4462), .ZN(U3311) );
  AND2_X1 U4982 ( .A1(D_REG_10__SCAN_IN), .A2(n4462), .ZN(U3312) );
  INV_X1 U4983 ( .A(D_REG_9__SCAN_IN), .ZN(n4657) );
  NOR2_X1 U4984 ( .A1(n4463), .A2(n4657), .ZN(U3313) );
  INV_X1 U4985 ( .A(D_REG_8__SCAN_IN), .ZN(n4663) );
  NOR2_X1 U4986 ( .A1(n4463), .A2(n4663), .ZN(U3314) );
  AND2_X1 U4987 ( .A1(D_REG_7__SCAN_IN), .A2(n4462), .ZN(U3315) );
  AND2_X1 U4988 ( .A1(D_REG_6__SCAN_IN), .A2(n4462), .ZN(U3316) );
  INV_X1 U4989 ( .A(D_REG_5__SCAN_IN), .ZN(n4675) );
  NOR2_X1 U4990 ( .A1(n4463), .A2(n4675), .ZN(U3317) );
  AND2_X1 U4991 ( .A1(n4462), .A2(D_REG_4__SCAN_IN), .ZN(U3318) );
  AND2_X1 U4992 ( .A1(D_REG_3__SCAN_IN), .A2(n4462), .ZN(U3319) );
  INV_X1 U4993 ( .A(D_REG_2__SCAN_IN), .ZN(n4674) );
  NOR2_X1 U4994 ( .A1(n4463), .A2(n4674), .ZN(U3320) );
  AOI21_X1 U4995 ( .B1(U3149), .B2(n2556), .A(n4464), .ZN(U3329) );
  INV_X1 U4996 ( .A(DATAI_17_), .ZN(n4465) );
  AOI22_X1 U4997 ( .A1(STATE_REG_SCAN_IN), .A2(n4466), .B1(n4465), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U4998 ( .A(DATAI_16_), .ZN(n4467) );
  AOI22_X1 U4999 ( .A1(STATE_REG_SCAN_IN), .A2(n4468), .B1(n4467), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5000 ( .A(DATAI_14_), .ZN(n4658) );
  AOI22_X1 U5001 ( .A1(STATE_REG_SCAN_IN), .A2(n2192), .B1(n4658), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5002 ( .A(DATAI_12_), .ZN(n4691) );
  AOI22_X1 U5003 ( .A1(STATE_REG_SCAN_IN), .A2(n4469), .B1(n4691), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5004 ( .A1(U3149), .A2(n4470), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4471) );
  INV_X1 U5005 ( .A(n4471), .ZN(U3341) );
  OAI22_X1 U5006 ( .A1(U3149), .A2(n4472), .B1(DATAI_10_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4473) );
  INV_X1 U5007 ( .A(n4473), .ZN(U3342) );
  OAI22_X1 U5008 ( .A1(U3149), .A2(IR_REG_0__SCAN_IN), .B1(DATAI_0_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4474) );
  INV_X1 U5009 ( .A(n4474), .ZN(U3352) );
  AOI22_X1 U5010 ( .A1(n4511), .A2(n4475), .B1(n2339), .B2(n4510), .ZN(U3467)
         );
  OAI22_X1 U5011 ( .A1(n4477), .A2(n4482), .B1(n4506), .B2(n4476), .ZN(n4478)
         );
  NOR2_X1 U5012 ( .A1(n4479), .A2(n4478), .ZN(n4512) );
  INV_X1 U5013 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4480) );
  AOI22_X1 U5014 ( .A1(n4511), .A2(n4512), .B1(n4480), .B2(n4510), .ZN(U3469)
         );
  OAI22_X1 U5015 ( .A1(n4483), .A2(n4482), .B1(n4506), .B2(n4481), .ZN(n4484)
         );
  NOR2_X1 U5016 ( .A1(n4485), .A2(n4484), .ZN(n4513) );
  INV_X1 U5017 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4486) );
  AOI22_X1 U5018 ( .A1(n4511), .A2(n4513), .B1(n4486), .B2(n4510), .ZN(U3473)
         );
  AOI211_X1 U5019 ( .C1(n4490), .C2(n4489), .A(n4488), .B(n4487), .ZN(n4514)
         );
  AOI22_X1 U5020 ( .A1(n4511), .A2(n4514), .B1(n2350), .B2(n4510), .ZN(U3475)
         );
  NOR2_X1 U5021 ( .A1(n4491), .A2(n4499), .ZN(n4494) );
  INV_X1 U5022 ( .A(n4492), .ZN(n4493) );
  AOI211_X1 U5023 ( .C1(n4496), .C2(n4495), .A(n4494), .B(n4493), .ZN(n4515)
         );
  INV_X1 U5024 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4497) );
  AOI22_X1 U5025 ( .A1(n4511), .A2(n4515), .B1(n4497), .B2(n4510), .ZN(U3477)
         );
  OR3_X1 U5026 ( .A1(n4500), .A2(n4499), .A3(n4498), .ZN(n4501) );
  AND3_X1 U5027 ( .A1(n4503), .A2(n4502), .A3(n4501), .ZN(n4516) );
  AOI22_X1 U5028 ( .A1(n4511), .A2(n4516), .B1(n2386), .B2(n4510), .ZN(U3481)
         );
  OAI21_X1 U5029 ( .B1(n4506), .B2(n4505), .A(n4504), .ZN(n4507) );
  AOI21_X1 U5030 ( .B1(n4509), .B2(n4508), .A(n4507), .ZN(n4518) );
  AOI22_X1 U5031 ( .A1(n4511), .A2(n4518), .B1(n2400), .B2(n4510), .ZN(U3485)
         );
  AOI22_X1 U5032 ( .A1(n4519), .A2(n4512), .B1(n2332), .B2(n4517), .ZN(U3519)
         );
  AOI22_X1 U5033 ( .A1(n4519), .A2(n4513), .B1(n2321), .B2(n4517), .ZN(U3521)
         );
  AOI22_X1 U5034 ( .A1(n4519), .A2(n4514), .B1(n2352), .B2(n4517), .ZN(U3522)
         );
  AOI22_X1 U5035 ( .A1(n4519), .A2(n4515), .B1(n2762), .B2(n4517), .ZN(U3523)
         );
  AOI22_X1 U5036 ( .A1(n4519), .A2(n4516), .B1(n2807), .B2(n4517), .ZN(U3525)
         );
  AOI22_X1 U5037 ( .A1(n4519), .A2(n4518), .B1(n2873), .B2(n4517), .ZN(U3527)
         );
  AOI22_X1 U5038 ( .A1(n2401), .A2(keyinput104), .B1(keyinput67), .B2(n4521), 
        .ZN(n4520) );
  OAI221_X1 U5039 ( .B1(n2401), .B2(keyinput104), .C1(n4521), .C2(keyinput67), 
        .A(n4520), .ZN(n4531) );
  AOI22_X1 U5040 ( .A1(n4663), .A2(keyinput118), .B1(keyinput84), .B2(n4523), 
        .ZN(n4522) );
  OAI221_X1 U5041 ( .B1(n4663), .B2(keyinput118), .C1(n4523), .C2(keyinput84), 
        .A(n4522), .ZN(n4530) );
  AOI22_X1 U5042 ( .A1(n4678), .A2(keyinput86), .B1(n4525), .B2(keyinput97), 
        .ZN(n4524) );
  OAI221_X1 U5043 ( .B1(n4678), .B2(keyinput86), .C1(n4525), .C2(keyinput97), 
        .A(n4524), .ZN(n4529) );
  INV_X1 U5044 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n4527) );
  AOI22_X1 U5045 ( .A1(n4527), .A2(keyinput72), .B1(keyinput82), .B2(n4677), 
        .ZN(n4526) );
  OAI221_X1 U5046 ( .B1(n4527), .B2(keyinput72), .C1(n4677), .C2(keyinput82), 
        .A(n4526), .ZN(n4528) );
  NOR4_X1 U5047 ( .A1(n4531), .A2(n4530), .A3(n4529), .A4(n4528), .ZN(n4568)
         );
  AOI22_X1 U5048 ( .A1(n4648), .A2(keyinput77), .B1(n3703), .B2(keyinput75), 
        .ZN(n4532) );
  OAI221_X1 U5049 ( .B1(n4648), .B2(keyinput77), .C1(n3703), .C2(keyinput75), 
        .A(n4532), .ZN(n4540) );
  AOI22_X1 U5050 ( .A1(n4189), .A2(keyinput96), .B1(keyinput73), .B2(n3074), 
        .ZN(n4533) );
  OAI221_X1 U5051 ( .B1(n4189), .B2(keyinput96), .C1(n3074), .C2(keyinput73), 
        .A(n4533), .ZN(n4539) );
  AOI22_X1 U5052 ( .A1(n4671), .A2(keyinput78), .B1(keyinput115), .B2(n4662), 
        .ZN(n4534) );
  OAI221_X1 U5053 ( .B1(n4671), .B2(keyinput78), .C1(n4662), .C2(keyinput115), 
        .A(n4534), .ZN(n4538) );
  AOI22_X1 U5054 ( .A1(n4536), .A2(keyinput94), .B1(n4672), .B2(keyinput79), 
        .ZN(n4535) );
  OAI221_X1 U5055 ( .B1(n4536), .B2(keyinput94), .C1(n4672), .C2(keyinput79), 
        .A(n4535), .ZN(n4537) );
  NOR4_X1 U5056 ( .A1(n4540), .A2(n4539), .A3(n4538), .A4(n4537), .ZN(n4567)
         );
  AOI22_X1 U5057 ( .A1(n4674), .A2(keyinput107), .B1(keyinput98), .B2(n4542), 
        .ZN(n4541) );
  OAI221_X1 U5058 ( .B1(n4674), .B2(keyinput107), .C1(n4542), .C2(keyinput98), 
        .A(n4541), .ZN(n4551) );
  AOI22_X1 U5059 ( .A1(n4545), .A2(keyinput88), .B1(n4544), .B2(keyinput64), 
        .ZN(n4543) );
  OAI221_X1 U5060 ( .B1(n4545), .B2(keyinput88), .C1(n4544), .C2(keyinput64), 
        .A(n4543), .ZN(n4550) );
  AOI22_X1 U5061 ( .A1(n4693), .A2(keyinput109), .B1(n4646), .B2(keyinput100), 
        .ZN(n4546) );
  OAI221_X1 U5062 ( .B1(n4693), .B2(keyinput109), .C1(n4646), .C2(keyinput100), 
        .A(n4546), .ZN(n4549) );
  AOI22_X1 U5063 ( .A1(n2282), .A2(keyinput116), .B1(keyinput89), .B2(n4686), 
        .ZN(n4547) );
  OAI221_X1 U5064 ( .B1(n2282), .B2(keyinput116), .C1(n4686), .C2(keyinput89), 
        .A(n4547), .ZN(n4548) );
  NOR4_X1 U5065 ( .A1(n4551), .A2(n4550), .A3(n4549), .A4(n4548), .ZN(n4566)
         );
  INV_X1 U5066 ( .A(DATAI_7_), .ZN(n4554) );
  INV_X1 U5067 ( .A(DATAI_8_), .ZN(n4553) );
  AOI22_X1 U5068 ( .A1(n4554), .A2(keyinput105), .B1(n4553), .B2(keyinput121), 
        .ZN(n4552) );
  OAI221_X1 U5069 ( .B1(n4554), .B2(keyinput105), .C1(n4553), .C2(keyinput121), 
        .A(n4552), .ZN(n4564) );
  AOI22_X1 U5070 ( .A1(n4556), .A2(keyinput106), .B1(keyinput74), .B2(n2954), 
        .ZN(n4555) );
  OAI221_X1 U5071 ( .B1(n4556), .B2(keyinput106), .C1(n2954), .C2(keyinput74), 
        .A(n4555), .ZN(n4563) );
  AOI22_X1 U5072 ( .A1(n4558), .A2(keyinput85), .B1(n2556), .B2(keyinput70), 
        .ZN(n4557) );
  OAI221_X1 U5073 ( .B1(n4558), .B2(keyinput85), .C1(n2556), .C2(keyinput70), 
        .A(n4557), .ZN(n4562) );
  XNOR2_X1 U5074 ( .A(IR_REG_16__SCAN_IN), .B(keyinput66), .ZN(n4560) );
  XNOR2_X1 U5075 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput122), .ZN(n4559) );
  NAND2_X1 U5076 ( .A1(n4560), .A2(n4559), .ZN(n4561) );
  NOR4_X1 U5077 ( .A1(n4564), .A2(n4563), .A3(n4562), .A4(n4561), .ZN(n4565)
         );
  AND4_X1 U5078 ( .A1(n4568), .A2(n4567), .A3(n4566), .A4(n4565), .ZN(n4705)
         );
  OAI22_X1 U5079 ( .A1(IR_REG_30__SCAN_IN), .A2(keyinput95), .B1(keyinput123), 
        .B2(ADDR_REG_19__SCAN_IN), .ZN(n4569) );
  AOI221_X1 U5080 ( .B1(IR_REG_30__SCAN_IN), .B2(keyinput95), .C1(
        ADDR_REG_19__SCAN_IN), .C2(keyinput123), .A(n4569), .ZN(n4576) );
  OAI22_X1 U5081 ( .A1(D_REG_9__SCAN_IN), .A2(keyinput68), .B1(
        REG3_REG_19__SCAN_IN), .B2(keyinput69), .ZN(n4570) );
  AOI221_X1 U5082 ( .B1(D_REG_9__SCAN_IN), .B2(keyinput68), .C1(keyinput69), 
        .C2(REG3_REG_19__SCAN_IN), .A(n4570), .ZN(n4575) );
  OAI22_X1 U5083 ( .A1(DATAO_REG_14__SCAN_IN), .A2(keyinput119), .B1(
        DATAO_REG_12__SCAN_IN), .B2(keyinput114), .ZN(n4571) );
  AOI221_X1 U5084 ( .B1(DATAO_REG_14__SCAN_IN), .B2(keyinput119), .C1(
        keyinput114), .C2(DATAO_REG_12__SCAN_IN), .A(n4571), .ZN(n4574) );
  OAI22_X1 U5085 ( .A1(DATAO_REG_3__SCAN_IN), .A2(keyinput124), .B1(
        DATAO_REG_0__SCAN_IN), .B2(keyinput65), .ZN(n4572) );
  AOI221_X1 U5086 ( .B1(DATAO_REG_3__SCAN_IN), .B2(keyinput124), .C1(
        keyinput65), .C2(DATAO_REG_0__SCAN_IN), .A(n4572), .ZN(n4573) );
  NAND4_X1 U5087 ( .A1(n4576), .A2(n4575), .A3(n4574), .A4(n4573), .ZN(n4604)
         );
  OAI22_X1 U5088 ( .A1(REG1_REG_7__SCAN_IN), .A2(keyinput120), .B1(keyinput111), .B2(ADDR_REG_18__SCAN_IN), .ZN(n4577) );
  AOI221_X1 U5089 ( .B1(REG1_REG_7__SCAN_IN), .B2(keyinput120), .C1(
        ADDR_REG_18__SCAN_IN), .C2(keyinput111), .A(n4577), .ZN(n4584) );
  OAI22_X1 U5090 ( .A1(REG2_REG_1__SCAN_IN), .A2(keyinput125), .B1(
        ADDR_REG_5__SCAN_IN), .B2(keyinput126), .ZN(n4578) );
  AOI221_X1 U5091 ( .B1(REG2_REG_1__SCAN_IN), .B2(keyinput125), .C1(
        keyinput126), .C2(ADDR_REG_5__SCAN_IN), .A(n4578), .ZN(n4583) );
  OAI22_X1 U5092 ( .A1(IR_REG_29__SCAN_IN), .A2(keyinput127), .B1(keyinput99), 
        .B2(REG1_REG_27__SCAN_IN), .ZN(n4579) );
  AOI221_X1 U5093 ( .B1(IR_REG_29__SCAN_IN), .B2(keyinput127), .C1(
        REG1_REG_27__SCAN_IN), .C2(keyinput99), .A(n4579), .ZN(n4582) );
  OAI22_X1 U5094 ( .A1(REG1_REG_5__SCAN_IN), .A2(keyinput83), .B1(
        REG1_REG_31__SCAN_IN), .B2(keyinput80), .ZN(n4580) );
  AOI221_X1 U5095 ( .B1(REG1_REG_5__SCAN_IN), .B2(keyinput83), .C1(keyinput80), 
        .C2(REG1_REG_31__SCAN_IN), .A(n4580), .ZN(n4581) );
  NAND4_X1 U5096 ( .A1(n4584), .A2(n4583), .A3(n4582), .A4(n4581), .ZN(n4603)
         );
  OAI22_X1 U5097 ( .A1(D_REG_28__SCAN_IN), .A2(keyinput93), .B1(
        REG0_REG_30__SCAN_IN), .B2(keyinput112), .ZN(n4585) );
  AOI221_X1 U5098 ( .B1(D_REG_28__SCAN_IN), .B2(keyinput93), .C1(keyinput112), 
        .C2(REG0_REG_30__SCAN_IN), .A(n4585), .ZN(n4592) );
  OAI22_X1 U5099 ( .A1(D_REG_29__SCAN_IN), .A2(keyinput81), .B1(keyinput110), 
        .B2(REG0_REG_12__SCAN_IN), .ZN(n4586) );
  AOI221_X1 U5100 ( .B1(D_REG_29__SCAN_IN), .B2(keyinput81), .C1(
        REG0_REG_12__SCAN_IN), .C2(keyinput110), .A(n4586), .ZN(n4591) );
  OAI22_X1 U5101 ( .A1(n4022), .A2(keyinput101), .B1(keyinput90), .B2(
        D_REG_5__SCAN_IN), .ZN(n4587) );
  AOI221_X1 U5102 ( .B1(n4022), .B2(keyinput101), .C1(D_REG_5__SCAN_IN), .C2(
        keyinput90), .A(n4587), .ZN(n4590) );
  OAI22_X1 U5103 ( .A1(D_REG_4__SCAN_IN), .A2(keyinput87), .B1(keyinput71), 
        .B2(REG0_REG_26__SCAN_IN), .ZN(n4588) );
  AOI221_X1 U5104 ( .B1(D_REG_4__SCAN_IN), .B2(keyinput87), .C1(
        REG0_REG_26__SCAN_IN), .C2(keyinput71), .A(n4588), .ZN(n4589) );
  NAND4_X1 U5105 ( .A1(n4592), .A2(n4591), .A3(n4590), .A4(n4589), .ZN(n4602)
         );
  OAI22_X1 U5106 ( .A1(IR_REG_5__SCAN_IN), .A2(keyinput91), .B1(DATAI_14_), 
        .B2(keyinput117), .ZN(n4593) );
  AOI221_X1 U5107 ( .B1(IR_REG_5__SCAN_IN), .B2(keyinput91), .C1(keyinput117), 
        .C2(DATAI_14_), .A(n4593), .ZN(n4600) );
  OAI22_X1 U5108 ( .A1(IR_REG_12__SCAN_IN), .A2(keyinput108), .B1(
        IR_REG_4__SCAN_IN), .B2(keyinput76), .ZN(n4594) );
  AOI221_X1 U5109 ( .B1(IR_REG_12__SCAN_IN), .B2(keyinput108), .C1(keyinput76), 
        .C2(IR_REG_4__SCAN_IN), .A(n4594), .ZN(n4599) );
  OAI22_X1 U5110 ( .A1(DATAI_12_), .A2(keyinput103), .B1(REG0_REG_0__SCAN_IN), 
        .B2(keyinput92), .ZN(n4595) );
  AOI221_X1 U5111 ( .B1(DATAI_12_), .B2(keyinput103), .C1(keyinput92), .C2(
        REG0_REG_0__SCAN_IN), .A(n4595), .ZN(n4598) );
  OAI22_X1 U5112 ( .A1(STATE_REG_SCAN_IN), .A2(keyinput102), .B1(keyinput113), 
        .B2(DATAI_16_), .ZN(n4596) );
  AOI221_X1 U5113 ( .B1(STATE_REG_SCAN_IN), .B2(keyinput102), .C1(DATAI_16_), 
        .C2(keyinput113), .A(n4596), .ZN(n4597) );
  NAND4_X1 U5114 ( .A1(n4600), .A2(n4599), .A3(n4598), .A4(n4597), .ZN(n4601)
         );
  NOR4_X1 U5115 ( .A1(n4604), .A2(n4603), .A3(n4602), .A4(n4601), .ZN(n4704)
         );
  AOI22_X1 U5116 ( .A1(REG0_REG_0__SCAN_IN), .A2(keyinput28), .B1(
        REG3_REG_10__SCAN_IN), .B2(keyinput58), .ZN(n4605) );
  OAI221_X1 U5117 ( .B1(REG0_REG_0__SCAN_IN), .B2(keyinput28), .C1(
        REG3_REG_10__SCAN_IN), .C2(keyinput58), .A(n4605), .ZN(n4612) );
  AOI22_X1 U5118 ( .A1(REG0_REG_12__SCAN_IN), .A2(keyinput46), .B1(
        REG3_REG_17__SCAN_IN), .B2(keyinput42), .ZN(n4606) );
  OAI221_X1 U5119 ( .B1(REG0_REG_12__SCAN_IN), .B2(keyinput46), .C1(
        REG3_REG_17__SCAN_IN), .C2(keyinput42), .A(n4606), .ZN(n4611) );
  AOI22_X1 U5120 ( .A1(REG1_REG_31__SCAN_IN), .A2(keyinput16), .B1(
        REG0_REG_31__SCAN_IN), .B2(keyinput24), .ZN(n4607) );
  OAI221_X1 U5121 ( .B1(REG1_REG_31__SCAN_IN), .B2(keyinput16), .C1(
        REG0_REG_31__SCAN_IN), .C2(keyinput24), .A(n4607), .ZN(n4610) );
  AOI22_X1 U5122 ( .A1(DATAO_REG_3__SCAN_IN), .A2(keyinput60), .B1(
        IR_REG_12__SCAN_IN), .B2(keyinput44), .ZN(n4608) );
  OAI221_X1 U5123 ( .B1(DATAO_REG_3__SCAN_IN), .B2(keyinput60), .C1(
        IR_REG_12__SCAN_IN), .C2(keyinput44), .A(n4608), .ZN(n4609) );
  NOR4_X1 U5124 ( .A1(n4612), .A2(n4611), .A3(n4610), .A4(n4609), .ZN(n4641)
         );
  AOI22_X1 U5125 ( .A1(REG1_REG_7__SCAN_IN), .A2(keyinput56), .B1(
        REG3_REG_9__SCAN_IN), .B2(keyinput40), .ZN(n4613) );
  OAI221_X1 U5126 ( .B1(REG1_REG_7__SCAN_IN), .B2(keyinput56), .C1(
        REG3_REG_9__SCAN_IN), .C2(keyinput40), .A(n4613), .ZN(n4620) );
  AOI22_X1 U5127 ( .A1(REG0_REG_27__SCAN_IN), .A2(keyinput0), .B1(
        REG3_REG_22__SCAN_IN), .B2(keyinput20), .ZN(n4614) );
  OAI221_X1 U5128 ( .B1(REG0_REG_27__SCAN_IN), .B2(keyinput0), .C1(
        REG3_REG_22__SCAN_IN), .C2(keyinput20), .A(n4614), .ZN(n4619) );
  AOI22_X1 U5129 ( .A1(ADDR_REG_0__SCAN_IN), .A2(keyinput8), .B1(
        IR_REG_0__SCAN_IN), .B2(keyinput33), .ZN(n4615) );
  OAI221_X1 U5130 ( .B1(ADDR_REG_0__SCAN_IN), .B2(keyinput8), .C1(
        IR_REG_0__SCAN_IN), .C2(keyinput33), .A(n4615), .ZN(n4618) );
  AOI22_X1 U5131 ( .A1(DATAI_7_), .A2(keyinput41), .B1(IR_REG_4__SCAN_IN), 
        .B2(keyinput12), .ZN(n4616) );
  OAI221_X1 U5132 ( .B1(DATAI_7_), .B2(keyinput41), .C1(IR_REG_4__SCAN_IN), 
        .C2(keyinput12), .A(n4616), .ZN(n4617) );
  NOR4_X1 U5133 ( .A1(n4620), .A2(n4619), .A3(n4618), .A4(n4617), .ZN(n4640)
         );
  AOI22_X1 U5134 ( .A1(DATAI_13_), .A2(keyinput21), .B1(DATAI_16_), .B2(
        keyinput49), .ZN(n4621) );
  OAI221_X1 U5135 ( .B1(DATAI_13_), .B2(keyinput21), .C1(DATAI_16_), .C2(
        keyinput49), .A(n4621), .ZN(n4628) );
  AOI22_X1 U5136 ( .A1(DATAO_REG_14__SCAN_IN), .A2(keyinput55), .B1(DATAI_8_), 
        .B2(keyinput57), .ZN(n4622) );
  OAI221_X1 U5137 ( .B1(DATAO_REG_14__SCAN_IN), .B2(keyinput55), .C1(DATAI_8_), 
        .C2(keyinput57), .A(n4622), .ZN(n4627) );
  AOI22_X1 U5138 ( .A1(ADDR_REG_18__SCAN_IN), .A2(keyinput47), .B1(
        REG1_REG_27__SCAN_IN), .B2(keyinput35), .ZN(n4623) );
  OAI221_X1 U5139 ( .B1(ADDR_REG_18__SCAN_IN), .B2(keyinput47), .C1(
        REG1_REG_27__SCAN_IN), .C2(keyinput35), .A(n4623), .ZN(n4626) );
  AOI22_X1 U5140 ( .A1(REG2_REG_31__SCAN_IN), .A2(keyinput11), .B1(
        IR_REG_5__SCAN_IN), .B2(keyinput27), .ZN(n4624) );
  OAI221_X1 U5141 ( .B1(REG2_REG_31__SCAN_IN), .B2(keyinput11), .C1(
        IR_REG_5__SCAN_IN), .C2(keyinput27), .A(n4624), .ZN(n4625) );
  NOR4_X1 U5142 ( .A1(n4628), .A2(n4627), .A3(n4626), .A4(n4625), .ZN(n4639)
         );
  AOI22_X1 U5143 ( .A1(DATAO_REG_4__SCAN_IN), .A2(keyinput3), .B1(
        D_REG_4__SCAN_IN), .B2(keyinput23), .ZN(n4629) );
  OAI221_X1 U5144 ( .B1(DATAO_REG_4__SCAN_IN), .B2(keyinput3), .C1(
        D_REG_4__SCAN_IN), .C2(keyinput23), .A(n4629), .ZN(n4637) );
  AOI22_X1 U5145 ( .A1(DATAI_23_), .A2(keyinput6), .B1(STATE_REG_SCAN_IN), 
        .B2(keyinput38), .ZN(n4630) );
  OAI221_X1 U5146 ( .B1(DATAI_23_), .B2(keyinput6), .C1(STATE_REG_SCAN_IN), 
        .C2(keyinput38), .A(n4630), .ZN(n4636) );
  AOI22_X1 U5147 ( .A1(REG1_REG_12__SCAN_IN), .A2(keyinput30), .B1(
        IR_REG_16__SCAN_IN), .B2(keyinput2), .ZN(n4631) );
  OAI221_X1 U5148 ( .B1(REG1_REG_12__SCAN_IN), .B2(keyinput30), .C1(
        IR_REG_16__SCAN_IN), .C2(keyinput2), .A(n4631), .ZN(n4635) );
  INV_X1 U5149 ( .A(ADDR_REG_19__SCAN_IN), .ZN(n4633) );
  AOI22_X1 U5150 ( .A1(D_REG_0__SCAN_IN), .A2(keyinput34), .B1(n4633), .B2(
        keyinput59), .ZN(n4632) );
  OAI221_X1 U5151 ( .B1(D_REG_0__SCAN_IN), .B2(keyinput34), .C1(n4633), .C2(
        keyinput59), .A(n4632), .ZN(n4634) );
  NOR4_X1 U5152 ( .A1(n4637), .A2(n4636), .A3(n4635), .A4(n4634), .ZN(n4638)
         );
  NAND4_X1 U5153 ( .A1(n4641), .A2(n4640), .A3(n4639), .A4(n4638), .ZN(n4703)
         );
  INV_X1 U5154 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n4643) );
  AOI22_X1 U5155 ( .A1(n4643), .A2(keyinput62), .B1(n2282), .B2(keyinput52), 
        .ZN(n4642) );
  OAI221_X1 U5156 ( .B1(n4643), .B2(keyinput62), .C1(n2282), .C2(keyinput52), 
        .A(n4642), .ZN(n4655) );
  AOI22_X1 U5157 ( .A1(n4646), .A2(keyinput36), .B1(keyinput48), .B2(n4645), 
        .ZN(n4644) );
  OAI221_X1 U5158 ( .B1(n4646), .B2(keyinput36), .C1(n4645), .C2(keyinput48), 
        .A(n4644), .ZN(n4654) );
  AOI22_X1 U5159 ( .A1(n4649), .A2(keyinput5), .B1(keyinput13), .B2(n4648), 
        .ZN(n4647) );
  OAI221_X1 U5160 ( .B1(n4649), .B2(keyinput5), .C1(n4648), .C2(keyinput13), 
        .A(n4647), .ZN(n4653) );
  AOI22_X1 U5161 ( .A1(n4651), .A2(keyinput1), .B1(n3074), .B2(keyinput9), 
        .ZN(n4650) );
  OAI221_X1 U5162 ( .B1(n4651), .B2(keyinput1), .C1(n3074), .C2(keyinput9), 
        .A(n4650), .ZN(n4652) );
  NOR4_X1 U5163 ( .A1(n4655), .A2(n4654), .A3(n4653), .A4(n4652), .ZN(n4701)
         );
  AOI22_X1 U5164 ( .A1(n4658), .A2(keyinput53), .B1(n4657), .B2(keyinput4), 
        .ZN(n4656) );
  OAI221_X1 U5165 ( .B1(n4658), .B2(keyinput53), .C1(n4657), .C2(keyinput4), 
        .A(n4656), .ZN(n4669) );
  AOI22_X1 U5166 ( .A1(n2257), .A2(keyinput63), .B1(keyinput50), .B2(n4660), 
        .ZN(n4659) );
  OAI221_X1 U5167 ( .B1(n2257), .B2(keyinput63), .C1(n4660), .C2(keyinput50), 
        .A(n4659), .ZN(n4668) );
  AOI22_X1 U5168 ( .A1(n4663), .A2(keyinput54), .B1(keyinput51), .B2(n4662), 
        .ZN(n4661) );
  OAI221_X1 U5169 ( .B1(n4663), .B2(keyinput54), .C1(n4662), .C2(keyinput51), 
        .A(n4661), .ZN(n4667) );
  XNOR2_X1 U5170 ( .A(REG2_REG_1__SCAN_IN), .B(keyinput61), .ZN(n4665) );
  XNOR2_X1 U5171 ( .A(keyinput32), .B(REG2_REG_13__SCAN_IN), .ZN(n4664) );
  NAND2_X1 U5172 ( .A1(n4665), .A2(n4664), .ZN(n4666) );
  NOR4_X1 U5173 ( .A1(n4669), .A2(n4668), .A3(n4667), .A4(n4666), .ZN(n4700)
         );
  AOI22_X1 U5174 ( .A1(n4672), .A2(keyinput15), .B1(n4671), .B2(keyinput14), 
        .ZN(n4670) );
  OAI221_X1 U5175 ( .B1(n4672), .B2(keyinput15), .C1(n4671), .C2(keyinput14), 
        .A(n4670), .ZN(n4684) );
  AOI22_X1 U5176 ( .A1(n4675), .A2(keyinput26), .B1(keyinput43), .B2(n4674), 
        .ZN(n4673) );
  OAI221_X1 U5177 ( .B1(n4675), .B2(keyinput26), .C1(n4674), .C2(keyinput43), 
        .A(n4673), .ZN(n4683) );
  AOI22_X1 U5178 ( .A1(n4678), .A2(keyinput22), .B1(n4677), .B2(keyinput18), 
        .ZN(n4676) );
  OAI221_X1 U5179 ( .B1(n4678), .B2(keyinput22), .C1(n4677), .C2(keyinput18), 
        .A(n4676), .ZN(n4682) );
  AOI22_X1 U5180 ( .A1(n4680), .A2(keyinput7), .B1(n2286), .B2(keyinput31), 
        .ZN(n4679) );
  OAI221_X1 U5181 ( .B1(n4680), .B2(keyinput7), .C1(n2286), .C2(keyinput31), 
        .A(n4679), .ZN(n4681) );
  NOR4_X1 U5182 ( .A1(n4684), .A2(n4683), .A3(n4682), .A4(n4681), .ZN(n4699)
         );
  AOI22_X1 U5183 ( .A1(n4686), .A2(keyinput25), .B1(keyinput37), .B2(n4022), 
        .ZN(n4685) );
  OAI221_X1 U5184 ( .B1(n4686), .B2(keyinput25), .C1(n4022), .C2(keyinput37), 
        .A(n4685), .ZN(n4697) );
  AOI22_X1 U5185 ( .A1(n4689), .A2(keyinput17), .B1(keyinput29), .B2(n4688), 
        .ZN(n4687) );
  OAI221_X1 U5186 ( .B1(n4689), .B2(keyinput17), .C1(n4688), .C2(keyinput29), 
        .A(n4687), .ZN(n4696) );
  AOI22_X1 U5187 ( .A1(n2762), .A2(keyinput19), .B1(n4691), .B2(keyinput39), 
        .ZN(n4690) );
  OAI221_X1 U5188 ( .B1(n2762), .B2(keyinput19), .C1(n4691), .C2(keyinput39), 
        .A(n4690), .ZN(n4695) );
  AOI22_X1 U5189 ( .A1(n4693), .A2(keyinput45), .B1(keyinput10), .B2(n2954), 
        .ZN(n4692) );
  OAI221_X1 U5190 ( .B1(n4693), .B2(keyinput45), .C1(n2954), .C2(keyinput10), 
        .A(n4692), .ZN(n4694) );
  NOR4_X1 U5191 ( .A1(n4697), .A2(n4696), .A3(n4695), .A4(n4694), .ZN(n4698)
         );
  NAND4_X1 U5192 ( .A1(n4701), .A2(n4700), .A3(n4699), .A4(n4698), .ZN(n4702)
         );
  AOI211_X1 U5193 ( .C1(n4705), .C2(n4704), .A(n4703), .B(n4702), .ZN(n4710)
         );
  NAND2_X1 U5194 ( .A1(n4706), .A2(U4043), .ZN(n4707) );
  OAI21_X1 U5195 ( .B1(U4043), .B2(DATAO_REG_23__SCAN_IN), .A(n4707), .ZN(
        n4709) );
  XNOR2_X1 U5196 ( .A(n4710), .B(n4709), .ZN(U3573) );
  CLKBUF_X3 U2302 ( .A(n2342), .Z(n2058) );
endmodule

