

module b15_C_SARLock_k_128_1 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024;

  OAI221_X1 U3559 ( .B1(n6830), .B2(keyinput82), .C1(n6829), .C2(
        W_R_N_REG_SCAN_IN), .A(n6828), .ZN(n6835) );
  INV_X2 U3560 ( .A(n5206), .ZN(n6039) );
  CLKBUF_X2 U3561 ( .A(n3866), .Z(n5456) );
  BUF_X1 U3562 ( .A(n5658), .Z(n3112) );
  INV_X2 U3563 ( .A(n3538), .ZN(n3795) );
  AND4_X1 U3564 ( .A1(n3146), .A2(n3145), .A3(n3144), .A4(n3143), .ZN(n3162)
         );
  AND4_X1 U3565 ( .A1(n3158), .A2(n3157), .A3(n3156), .A4(n3155), .ZN(n3159)
         );
  BUF_X2 U3566 ( .A(n3496), .Z(n4949) );
  CLKBUF_X2 U3567 ( .A(n3269), .Z(n5619) );
  CLKBUF_X2 U3568 ( .A(n3249), .Z(n5634) );
  AND2_X1 U3569 ( .A1(n5808), .A2(n3705), .ZN(n3267) );
  AND2_X1 U3570 ( .A1(n5808), .A2(n3704), .ZN(n3517) );
  AND2_X2 U3571 ( .A1(n3128), .A2(n5800), .ZN(n3501) );
  AND2_X2 U3572 ( .A1(n3399), .A2(n3705), .ZN(n3518) );
  AOI22_X1 U3573 ( .A1(n4048), .A2(keyinput70), .B1(keyinput88), .B2(n6912), 
        .ZN(n6911) );
  AOI22_X1 U3574 ( .A1(n6859), .A2(keyinput108), .B1(keyinput118), .B2(n6858), 
        .ZN(n6857) );
  AOI22_X1 U3575 ( .A1(n6830), .A2(keyinput82), .B1(W_R_N_REG_SCAN_IN), .B2(
        n6829), .ZN(n6828) );
  AND2_X1 U3576 ( .A1(n3354), .A2(n3397), .ZN(n3378) );
  OAI221_X1 U3577 ( .B1(n4048), .B2(keyinput70), .C1(n6912), .C2(keyinput88), 
        .A(n6911), .ZN(n6920) );
  OAI221_X1 U3578 ( .B1(n6859), .B2(keyinput108), .C1(n6858), .C2(keyinput118), 
        .A(n6857), .ZN(n6868) );
  OAI22_X1 U3579 ( .A1(n4334), .A2(keyinput7), .B1(n6795), .B2(keyinput44), 
        .ZN(n6794) );
  NAND2_X2 U3580 ( .A1(n3646), .A2(n3370), .ZN(n4155) );
  OAI22_X1 U3581 ( .A1(n6131), .A2(n5646), .B1(n5005), .B2(n6795), .ZN(n4660)
         );
  AOI221_X1 U3582 ( .B1(n4334), .B2(keyinput7), .C1(keyinput44), .C2(n6795), 
        .A(n6794), .ZN(n6808) );
  OR2_X1 U3583 ( .A1(n5436), .A2(n5435), .ZN(n5485) );
  NAND4_X2 U3584 ( .A1(n3162), .A2(n3161), .A3(n3160), .A4(n3159), .ZN(n3645)
         );
  OR2_X1 U3585 ( .A1(n5271), .A2(n5270), .ZN(n5403) );
  NOR2_X4 U3586 ( .A1(n3352), .A2(n3301), .ZN(n3350) );
  BUF_X2 U3587 ( .A(n3743), .Z(n5946) );
  NAND2_X1 U3589 ( .A1(n3799), .A2(n3645), .ZN(n5658) );
  INV_X2 U3590 ( .A(n3808), .ZN(n5679) );
  INV_X1 U3591 ( .A(n3516), .ZN(n4496) );
  CLKBUF_X2 U3592 ( .A(n5619), .Z(n5692) );
  CLKBUF_X2 U3593 ( .A(n3501), .Z(n3607) );
  CLKBUF_X2 U3594 ( .A(n3270), .Z(n3608) );
  CLKBUF_X2 U3595 ( .A(n3517), .Z(n5689) );
  INV_X2 U3596 ( .A(n3248), .ZN(n3516) );
  CLKBUF_X2 U3597 ( .A(n3495), .Z(n5682) );
  AND2_X1 U3598 ( .A1(n5243), .A2(n5242), .ZN(n6317) );
  OR2_X1 U3599 ( .A1(n5241), .A2(n5195), .ZN(n5205) );
  NAND2_X1 U3600 ( .A1(n4891), .A2(n4890), .ZN(n5241) );
  AND2_X1 U3601 ( .A1(n5212), .A2(n5596), .ZN(n5213) );
  NAND2_X2 U3602 ( .A1(n4463), .A2(n4462), .ZN(n5209) );
  AND2_X1 U3604 ( .A1(n3871), .A2(n3870), .ZN(n3982) );
  AND2_X1 U3605 ( .A1(n3649), .A2(n5169), .ZN(n3589) );
  OR2_X1 U3606 ( .A1(n3353), .A2(n4155), .ZN(n3397) );
  NAND2_X1 U3607 ( .A1(n3345), .A2(n3344), .ZN(n3372) );
  AND2_X2 U3608 ( .A1(n3646), .A2(n3645), .ZN(n5457) );
  AND4_X1 U3609 ( .A1(n3127), .A2(n3126), .A3(n3125), .A4(n3124), .ZN(n3141)
         );
  INV_X1 U3610 ( .A(n3646), .ZN(n3790) );
  AND4_X1 U3611 ( .A1(n3281), .A2(n3280), .A3(n3279), .A4(n3278), .ZN(n3298)
         );
  AND4_X1 U3612 ( .A1(n3286), .A2(n3285), .A3(n3284), .A4(n3283), .ZN(n3297)
         );
  OR2_X2 U3613 ( .A1(n3172), .A2(n3171), .ZN(n3646) );
  AND4_X1 U3614 ( .A1(n3150), .A2(n3149), .A3(n3148), .A4(n3147), .ZN(n3161)
         );
  AND4_X1 U3615 ( .A1(n3154), .A2(n3153), .A3(n3152), .A4(n3151), .ZN(n3160)
         );
  BUF_X2 U3616 ( .A(n3267), .Z(n5080) );
  INV_X2 U3617 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3214) );
  OR2_X1 U3618 ( .A1(n5241), .A2(n5240), .ZN(n5243) );
  XNOR2_X1 U3619 ( .A(n3467), .B(n3466), .ZN(n3494) );
  INV_X2 U3620 ( .A(n3725), .ZN(n6080) );
  AND2_X4 U3621 ( .A1(n3133), .A2(n3707), .ZN(n3270) );
  AND2_X4 U3622 ( .A1(n3133), .A2(n3705), .ZN(n3241) );
  NOR2_X2 U3623 ( .A1(n5316), .A2(n5315), .ZN(n5317) );
  OR2_X2 U3624 ( .A1(n5042), .A2(n5041), .ZN(n5316) );
  XNOR2_X2 U3625 ( .A(n4000), .B(n6413), .ZN(n3999) );
  OAI21_X2 U3626 ( .B1(n3953), .B2(n4460), .A(n3742), .ZN(n4000) );
  BUF_X4 U3627 ( .A(n4155), .Z(n5659) );
  OAI21_X2 U3628 ( .B1(n5667), .B2(n5666), .A(n5772), .ZN(n5846) );
  AOI211_X2 U3629 ( .C1(n5841), .C2(REIP_REG_29__SCAN_IN), .A(n5675), .B(n5674), .ZN(n5676) );
  INV_X1 U3630 ( .A(n6238), .ZN(n3111) );
  OR3_X4 U3631 ( .A1(n6234), .A2(n5188), .A3(n5806), .ZN(n6238) );
  NAND2_X1 U3632 ( .A1(n4068), .A2(n6580), .ZN(n3620) );
  INV_X1 U3633 ( .A(n3300), .ZN(n3322) );
  NAND2_X1 U3634 ( .A1(n4148), .A2(n4147), .ZN(n4463) );
  AND2_X1 U3635 ( .A1(n4782), .A2(n4783), .ZN(n4971) );
  AND2_X1 U3636 ( .A1(n4909), .A2(n4882), .ZN(n4783) );
  INV_X1 U3637 ( .A(n4146), .ZN(n4446) );
  NAND2_X1 U3638 ( .A1(n3387), .A2(n3386), .ZN(n3673) );
  OR2_X1 U3639 ( .A1(n3363), .A2(n3423), .ZN(n3387) );
  NOR2_X1 U3640 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n3773), .ZN(n4261) );
  INV_X1 U3641 ( .A(n5792), .ZN(n5188) );
  OR2_X1 U3642 ( .A1(n6234), .A2(n6814), .ZN(n5817) );
  NAND2_X1 U3643 ( .A1(n3995), .A2(n3865), .ZN(n3983) );
  NAND2_X1 U3644 ( .A1(n5092), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5267)
         );
  NAND2_X1 U3645 ( .A1(n4488), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4503)
         );
  OR2_X1 U3646 ( .A1(n3643), .A2(n6587), .ZN(n3739) );
  AND4_X1 U3647 ( .A1(n3132), .A2(n3131), .A3(n3130), .A4(n3129), .ZN(n3140)
         );
  AND2_X1 U3648 ( .A1(n3419), .A2(n3418), .ZN(n3727) );
  AND2_X1 U3649 ( .A1(n5946), .A2(n4237), .ZN(n4352) );
  INV_X1 U3650 ( .A(n5031), .ZN(n5372) );
  CLKBUF_X1 U3651 ( .A(n5118), .Z(n6445) );
  NAND2_X1 U3652 ( .A1(n3262), .A2(n4787), .ZN(n3300) );
  OR2_X1 U3653 ( .A1(n3843), .A2(n3842), .ZN(n4150) );
  NAND2_X1 U3654 ( .A1(n3816), .A2(n3817), .ZN(n3843) );
  INV_X1 U3655 ( .A(n3819), .ZN(n3816) );
  OR2_X1 U3656 ( .A1(n5240), .A2(n5194), .ZN(n5195) );
  NOR2_X1 U3657 ( .A1(n3388), .A2(n3746), .ZN(n3358) );
  INV_X1 U3658 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5471) );
  OR2_X1 U3659 ( .A1(n5192), .A2(n3115), .ZN(n5240) );
  INV_X1 U3660 ( .A(n4448), .ZN(n4460) );
  OR2_X1 U3661 ( .A1(n3508), .A2(n3507), .ZN(n4464) );
  OAI21_X1 U3662 ( .B1(n6080), .B2(n3341), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3360) );
  OAI21_X1 U3663 ( .B1(n3534), .B2(n3355), .A(n3539), .ZN(n3341) );
  AND2_X1 U3664 ( .A1(n3551), .A2(n3550), .ZN(n3626) );
  OR2_X1 U3665 ( .A1(n3395), .A2(n3379), .ZN(n3465) );
  AOI21_X1 U3666 ( .B1(n6582), .B2(n3735), .A(n5807), .ZN(n3773) );
  OR2_X1 U3667 ( .A1(n3739), .A2(n3534), .ZN(n3313) );
  NOR2_X1 U3668 ( .A1(n5070), .A2(n4860), .ZN(n5017) );
  OR2_X1 U3669 ( .A1(n5267), .A2(n5885), .ZN(n5385) );
  AND2_X1 U3670 ( .A1(n5095), .A2(n5094), .ZN(n5096) );
  OR2_X1 U3671 ( .A1(n5519), .A2(n5703), .ZN(n5094) );
  AND2_X1 U3672 ( .A1(n4971), .A2(n4970), .ZN(n4972) );
  NOR2_X1 U3673 ( .A1(n4629), .A2(n5425), .ZN(n4596) );
  NAND2_X1 U3674 ( .A1(n4596), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4963)
         );
  NAND2_X1 U3675 ( .A1(n4630), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4629)
         );
  NAND2_X1 U3676 ( .A1(n4659), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4777)
         );
  NOR2_X1 U3677 ( .A1(n6795), .A2(n4757), .ZN(n4659) );
  NAND2_X1 U3678 ( .A1(n4704), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4673)
         );
  NOR2_X1 U3679 ( .A1(n6912), .A2(n4673), .ZN(n4758) );
  NOR2_X1 U3680 ( .A1(n6858), .A2(n4720), .ZN(n4704) );
  NAND2_X1 U3681 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n4725), .ZN(n4720)
         );
  NAND2_X1 U3682 ( .A1(n4508), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4578)
         );
  INV_X1 U3683 ( .A(n4503), .ZN(n4508) );
  AOI21_X1 U3684 ( .B1(n4491), .B2(n4754), .A(n4490), .ZN(n4870) );
  CLKBUF_X1 U3685 ( .A(n4830), .Z(n4868) );
  NOR2_X1 U3686 ( .A1(n4210), .A2(n6195), .ZN(n4488) );
  INV_X1 U3687 ( .A(n3845), .ZN(n3846) );
  NAND2_X1 U3688 ( .A1(n3846), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4210)
         );
  NAND2_X1 U3689 ( .A1(n3821), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3845)
         );
  NAND2_X1 U3690 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3695) );
  NAND2_X1 U3691 ( .A1(n5832), .A2(n5831), .ZN(n5834) );
  AND2_X1 U3692 ( .A1(n5573), .A2(n5574), .ZN(n5832) );
  NOR2_X1 U3693 ( .A1(n5463), .A2(n5462), .ZN(n5573) );
  AND2_X1 U3694 ( .A1(n6039), .A2(n6974), .ZN(n5547) );
  OR2_X1 U3695 ( .A1(n5162), .A2(n5161), .ZN(n5463) );
  AND2_X1 U3696 ( .A1(n5017), .A2(n5016), .ZN(n5063) );
  NAND2_X1 U3697 ( .A1(n5063), .A2(n5062), .ZN(n5162) );
  INV_X1 U3698 ( .A(n5929), .ZN(n5936) );
  OR2_X1 U3699 ( .A1(n5515), .A2(n5420), .ZN(n5422) );
  NAND2_X1 U3700 ( .A1(n5102), .A2(n4840), .ZN(n4916) );
  AND2_X1 U3701 ( .A1(n5538), .A2(n5196), .ZN(n5494) );
  NAND2_X1 U3702 ( .A1(n5024), .A2(n5023), .ZN(n5042) );
  NAND2_X1 U3703 ( .A1(n4472), .A2(n4471), .ZN(n4479) );
  INV_X1 U3704 ( .A(n4794), .ZN(n4472) );
  NAND2_X1 U3705 ( .A1(n4458), .A2(n4457), .ZN(n4888) );
  INV_X1 U3706 ( .A(n3982), .ZN(n3872) );
  AND2_X1 U3707 ( .A1(n3541), .A2(n3488), .ZN(n4164) );
  NAND2_X1 U3708 ( .A1(n3494), .A2(n6580), .ZN(n3551) );
  XNOR2_X1 U3709 ( .A(n3623), .B(n3622), .ZN(n3631) );
  NAND2_X1 U3710 ( .A1(n3620), .A2(n3619), .ZN(n3623) );
  NAND2_X1 U3711 ( .A1(n3631), .A2(n3632), .ZN(n3692) );
  OR2_X2 U3712 ( .A1(n3692), .A2(n3943), .ZN(n3819) );
  INV_X1 U3713 ( .A(n5801), .ZN(n3472) );
  INV_X1 U3714 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3119) );
  NAND2_X1 U3715 ( .A1(n3674), .A2(n3673), .ZN(n3723) );
  INV_X1 U3716 ( .A(n5946), .ZN(n4230) );
  AND2_X1 U3717 ( .A1(n6667), .A2(n3942), .ZN(n6490) );
  AND4_X1 U3718 ( .A1(n3290), .A2(n3289), .A3(n3288), .A4(n3287), .ZN(n3296)
         );
  INV_X1 U3719 ( .A(n5111), .ZN(n4237) );
  OR3_X1 U3720 ( .A1(n6826), .A2(STATE2_REG_0__SCAN_IN), .A3(n3773), .ZN(n3925) );
  NAND2_X1 U3721 ( .A1(n3236), .A2(n3235), .ZN(n3643) );
  CLKBUF_X1 U3722 ( .A(n5703), .Z(n5646) );
  INV_X1 U3723 ( .A(n6220), .ZN(n6235) );
  OR2_X1 U3724 ( .A1(n5817), .A2(n5175), .ZN(n6209) );
  INV_X1 U3725 ( .A(n6199), .ZN(n6190) );
  CLKBUF_X1 U3726 ( .A(n3702), .Z(n5469) );
  INV_X1 U3727 ( .A(n6175), .ZN(n6231) );
  AND2_X1 U3728 ( .A1(n5796), .A2(n3596), .ZN(n6248) );
  AND2_X1 U3729 ( .A1(n5796), .A2(n4789), .ZN(n6251) );
  XNOR2_X1 U3730 ( .A(n5171), .B(n5818), .ZN(n5792) );
  AND2_X1 U3731 ( .A1(n5037), .A2(n4928), .ZN(n5031) );
  NAND2_X1 U3732 ( .A1(n6339), .A2(n6362), .ZN(n6355) );
  INV_X1 U3733 ( .A(n6339), .ZN(n6363) );
  INV_X1 U3734 ( .A(n6405), .ZN(n6428) );
  INV_X1 U3735 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3118) );
  OR2_X1 U3736 ( .A1(n3781), .A2(n5111), .ZN(n4525) );
  OAI21_X1 U3737 ( .B1(n4406), .B2(n6826), .A(n4405), .ZN(n4430) );
  INV_X1 U3738 ( .A(n4434), .ZN(n4399) );
  INV_X1 U3739 ( .A(n5155), .ZN(n5113) );
  INV_X1 U3740 ( .A(n4346), .ZN(n4339) );
  NOR2_X1 U3741 ( .A1(n4189), .A2(n4237), .ZN(n4346) );
  AND2_X1 U3742 ( .A1(n3889), .A2(n4237), .ZN(n4054) );
  NAND2_X1 U3743 ( .A1(n3359), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3363) );
  NOR2_X1 U3744 ( .A1(n5864), .A2(n5516), .ZN(n5548) );
  AND2_X2 U3745 ( .A1(n3704), .A2(n3399), .ZN(n3255) );
  INV_X2 U3746 ( .A(n5901), .ZN(n6360) );
  NAND2_X1 U3747 ( .A1(n5209), .A2(n6930), .ZN(n3113) );
  AND2_X1 U3748 ( .A1(n5723), .A2(n5722), .ZN(n3114) );
  NOR2_X1 U3749 ( .A1(n5209), .A2(n6385), .ZN(n3115) );
  OR2_X1 U3750 ( .A1(n5774), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3116)
         );
  OR2_X1 U3751 ( .A1(n5774), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3117)
         );
  INV_X1 U3752 ( .A(n5209), .ZN(n5206) );
  INV_X1 U3753 ( .A(n3576), .ZN(n3345) );
  OAI21_X1 U3754 ( .B1(n3472), .B2(n3759), .A(n5176), .ZN(n3347) );
  OAI21_X1 U3755 ( .B1(n3350), .B2(n3349), .A(n3348), .ZN(n3351) );
  AND2_X1 U3756 ( .A1(n3538), .A2(n3852), .ZN(n3344) );
  NAND2_X1 U3757 ( .A1(n5185), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3189) );
  INV_X1 U3758 ( .A(n3255), .ZN(n3502) );
  NOR2_X1 U3759 ( .A1(n3857), .A2(n4155), .ZN(n3866) );
  CLKBUF_X3 U3760 ( .A(n3249), .Z(n5683) );
  INV_X1 U3761 ( .A(n4795), .ZN(n4471) );
  INV_X1 U3762 ( .A(n4150), .ZN(n4148) );
  INV_X1 U3763 ( .A(n3189), .ZN(n3190) );
  INV_X1 U3764 ( .A(n3465), .ZN(n3466) );
  OR2_X1 U3765 ( .A1(n5185), .A2(n6580), .ZN(n3567) );
  INV_X1 U3766 ( .A(n4777), .ZN(n4579) );
  OR2_X1 U3767 ( .A1(n4578), .A2(n6163), .ZN(n4724) );
  AND2_X1 U3768 ( .A1(n3113), .A2(n5494), .ZN(n5437) );
  AND2_X1 U3769 ( .A1(n3646), .A2(n3747), .ZN(n4448) );
  INV_X1 U3770 ( .A(n3983), .ZN(n3873) );
  AND4_X1 U3771 ( .A1(n3138), .A2(n3137), .A3(n3136), .A4(n3135), .ZN(n3139)
         );
  NAND2_X1 U3772 ( .A1(n3587), .A2(n3567), .ZN(n4443) );
  INV_X1 U3773 ( .A(n5456), .ZN(n5662) );
  OR2_X1 U3774 ( .A1(n3538), .A2(n6580), .ZN(n3587) );
  AND2_X1 U3775 ( .A1(n3585), .A2(n4787), .ZN(n3571) );
  OR2_X1 U3776 ( .A1(n5705), .A2(n6842), .ZN(n5171) );
  NAND2_X1 U3777 ( .A1(n5612), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5705)
         );
  AND2_X1 U3778 ( .A1(n5091), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5092)
         );
  AND2_X1 U3779 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n4579), .ZN(n4630)
         );
  NOR2_X1 U3780 ( .A1(n6830), .A2(n4724), .ZN(n4725) );
  XNOR2_X1 U3781 ( .A(n4463), .B(n4447), .ZN(n4491) );
  INV_X1 U3782 ( .A(n5457), .ZN(n5773) );
  AND2_X1 U3783 ( .A1(n6039), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5725)
         );
  AND2_X1 U3784 ( .A1(n5486), .A2(n5208), .ZN(n5492) );
  NAND2_X1 U3785 ( .A1(n3873), .A2(n3872), .ZN(n3989) );
  NAND2_X1 U3786 ( .A1(n3365), .A2(n3364), .ZN(n3467) );
  NAND2_X1 U3787 ( .A1(n3702), .A2(n6580), .ZN(n3691) );
  XNOR2_X1 U3788 ( .A(n3723), .B(n5114), .ZN(n3702) );
  AND4_X1 U3789 ( .A1(n3294), .A2(n3293), .A3(n3292), .A4(n3291), .ZN(n3295)
         );
  OR2_X1 U3790 ( .A1(n3233), .A2(n3232), .ZN(n3236) );
  AOI21_X1 U3791 ( .B1(n5821), .B2(n6656), .A(n5721), .ZN(n5722) );
  OR2_X1 U3792 ( .A1(n4963), .A2(n5900), .ZN(n4965) );
  OR2_X1 U3793 ( .A1(n6209), .A2(n5332), .ZN(n5352) );
  INV_X1 U3794 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6195) );
  OR2_X1 U3795 ( .A1(n6234), .A2(n6826), .ZN(n6220) );
  AND2_X1 U3796 ( .A1(n3340), .A2(n3799), .ZN(n3649) );
  OR2_X1 U3797 ( .A1(n5385), .A2(n6910), .ZN(n5647) );
  NAND2_X1 U3798 ( .A1(n4979), .A2(n4972), .ZN(n5008) );
  NAND2_X1 U3799 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n4758), .ZN(n4757)
         );
  AND2_X1 U3800 ( .A1(n4921), .A2(n4920), .ZN(n5106) );
  AND2_X1 U3801 ( .A1(n5201), .A2(n5200), .ZN(n5242) );
  NOR2_X1 U3802 ( .A1(n3831), .A2(n3830), .ZN(n4009) );
  NAND2_X1 U3803 ( .A1(n5863), .A2(n5725), .ZN(n5877) );
  OR2_X1 U3804 ( .A1(n5211), .A2(n5210), .ZN(n5596) );
  OR2_X1 U3805 ( .A1(n3739), .A2(n3483), .ZN(n3484) );
  NAND2_X1 U3806 ( .A1(n3467), .A2(n3465), .ZN(n3552) );
  OR2_X1 U3807 ( .A1(n3781), .A2(n4237), .ZN(n4114) );
  NAND2_X1 U3808 ( .A1(n3952), .A2(n4352), .ZN(n4432) );
  AND2_X1 U3809 ( .A1(n3691), .A2(n3690), .ZN(n3943) );
  INV_X1 U3810 ( .A(n5283), .ZN(n5325) );
  NAND2_X1 U3811 ( .A1(n3679), .A2(n3678), .ZN(n5114) );
  NAND2_X1 U3812 ( .A1(n3313), .A2(n5960), .ZN(n6686) );
  NOR2_X1 U3813 ( .A1(n4965), .A2(n4964), .ZN(n5091) );
  NOR2_X1 U3814 ( .A1(n6917), .A2(n6120), .ZN(n6111) );
  NOR2_X1 U3815 ( .A1(n6628), .A2(n5352), .ZN(n6156) );
  NAND2_X1 U3816 ( .A1(n4162), .A2(n4161), .ZN(n4794) );
  NOR2_X1 U3817 ( .A1(n6686), .A2(n5168), .ZN(n6234) );
  MUX2_X1 U3818 ( .A(n5710), .B(n5659), .S(n5834), .Z(n5712) );
  NOR2_X1 U3819 ( .A1(n4063), .A2(n3881), .ZN(n4162) );
  NAND2_X1 U3820 ( .A1(n3112), .A2(n5659), .ZN(n5774) );
  NAND2_X1 U3821 ( .A1(n5097), .A2(n5096), .ZN(n5271) );
  INV_X1 U3822 ( .A(n5796), .ZN(n6250) );
  INV_X1 U3823 ( .A(n6285), .ZN(n3460) );
  INV_X1 U3824 ( .A(n3645), .ZN(n3785) );
  INV_X1 U3825 ( .A(n6313), .ZN(n6698) );
  NOR2_X1 U3826 ( .A1(n5403), .A2(n5404), .ZN(n5830) );
  AND2_X1 U3827 ( .A1(n4912), .A2(n4911), .ZN(n6008) );
  AND2_X1 U3828 ( .A1(n5049), .A2(n4933), .ZN(n6249) );
  AND2_X1 U3829 ( .A1(n5107), .A2(n5038), .ZN(n6320) );
  INV_X1 U3830 ( .A(n6355), .ZN(n6332) );
  NOR2_X1 U3831 ( .A1(n5558), .A2(n5559), .ZN(n5580) );
  AND2_X1 U3832 ( .A1(n6052), .A2(n5231), .ZN(n5929) );
  AND2_X1 U3833 ( .A1(n5507), .A2(n5221), .ZN(n6052) );
  NOR2_X1 U3834 ( .A1(n5225), .A2(n6372), .ZN(n5507) );
  AND2_X1 U3835 ( .A1(n3541), .A2(n3540), .ZN(n6405) );
  NAND2_X1 U3836 ( .A1(n3485), .A2(n3484), .ZN(n3541) );
  INV_X1 U3837 ( .A(n6406), .ZN(n6434) );
  INV_X1 U3838 ( .A(n6416), .ZN(n5222) );
  INV_X1 U3839 ( .A(n4261), .ZN(n4310) );
  INV_X1 U3840 ( .A(n6581), .ZN(n5807) );
  INV_X1 U3841 ( .A(n4525), .ZN(n4561) );
  NOR2_X1 U3842 ( .A1(n4238), .A2(n4237), .ZN(n4434) );
  NOR2_X1 U3843 ( .A1(n4238), .A2(n5111), .ZN(n5155) );
  AND2_X1 U3844 ( .A1(n5950), .A2(n3943), .ZN(n5112) );
  AND2_X1 U3845 ( .A1(n4190), .A2(n4237), .ZN(n5283) );
  AND2_X1 U3846 ( .A1(n5277), .A2(n6445), .ZN(n5286) );
  INV_X1 U3847 ( .A(n6539), .ZN(n6542) );
  OR2_X1 U3848 ( .A1(n3643), .A2(n6826), .ZN(n6581) );
  INV_X1 U3849 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6580) );
  OR2_X1 U3850 ( .A1(n5817), .A2(n5187), .ZN(n6175) );
  OR2_X1 U3851 ( .A1(n6234), .A2(n5172), .ZN(n6199) );
  OR2_X1 U3852 ( .A1(n5817), .A2(n5177), .ZN(n6243) );
  INV_X1 U3853 ( .A(n6320), .ZN(n5358) );
  NAND2_X1 U3854 ( .A1(n6298), .A2(n3595), .ZN(n5796) );
  NOR2_X1 U3855 ( .A1(n3460), .A2(n6689), .ZN(n6280) );
  NAND2_X1 U3856 ( .A1(n3459), .A2(n3475), .ZN(n6285) );
  NAND2_X1 U3857 ( .A1(n3316), .A2(n3315), .ZN(n6298) );
  NAND2_X1 U3858 ( .A1(n6323), .A2(n3767), .ZN(n6339) );
  OR2_X1 U3859 ( .A1(n3739), .A2(n6566), .ZN(n6323) );
  INV_X1 U3860 ( .A(n6055), .ZN(n6372) );
  INV_X1 U3861 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6927) );
  INV_X1 U3862 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n6872) );
  AND2_X1 U3863 ( .A1(n4021), .A2(n4020), .ZN(n4060) );
  NOR2_X1 U3864 ( .A1(n4312), .A2(n4311), .ZN(n4351) );
  NOR2_X1 U3865 ( .A1(n4359), .A2(n4358), .ZN(n4397) );
  INV_X1 U3866 ( .A(n3939), .ZN(n3933) );
  INV_X1 U3867 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4181) );
  AOI22_X1 U3868 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n4181), .B1(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6872), .ZN(n3200) );
  NAND2_X1 U3869 ( .A1(n6927), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3183) );
  INV_X1 U3870 ( .A(n3183), .ZN(n3199) );
  XOR2_X1 U3871 ( .A(n3200), .B(n3199), .Z(n3305) );
  NAND2_X1 U3872 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n3305), .ZN(n3198) );
  INV_X2 U3873 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3468) );
  AND2_X2 U3874 ( .A1(n3468), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3133)
         );
  AND2_X2 U3875 ( .A1(n3214), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3128)
         );
  AND2_X2 U3876 ( .A1(n3133), .A2(n3128), .ZN(n3248) );
  NAND2_X1 U3877 ( .A1(n4496), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3123) );
  AND2_X2 U3878 ( .A1(n3118), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5808)
         );
  AND2_X2 U3879 ( .A1(n5808), .A2(n3128), .ZN(n3249) );
  NAND2_X1 U3880 ( .A1(n5683), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3122) );
  AND2_X2 U3881 ( .A1(n3119), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3707)
         );
  AND2_X2 U3882 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3399) );
  AND2_X2 U3883 ( .A1(n3707), .A2(n3399), .ZN(n3511) );
  NAND2_X1 U3884 ( .A1(n3511), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3121)
         );
  NOR2_X4 U3885 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3704) );
  NAND2_X1 U3886 ( .A1(n3517), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3120) );
  AND2_X2 U3888 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3705) );
  NAND2_X1 U3889 ( .A1(n5080), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3127)
         );
  AND2_X2 U3890 ( .A1(n3133), .A2(n3704), .ZN(n3254) );
  NAND2_X1 U3891 ( .A1(n5679), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3126) );
  NOR2_X4 U3892 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5800) );
  AND2_X2 U3893 ( .A1(n3707), .A2(n5800), .ZN(n3268) );
  BUF_X2 U3894 ( .A(n3268), .Z(n4728) );
  NAND2_X1 U3895 ( .A1(n4728), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3125) );
  AND2_X2 U3896 ( .A1(n3128), .A2(n3399), .ZN(n3269) );
  NAND2_X1 U3897 ( .A1(n5619), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3124) );
  AND2_X2 U3898 ( .A1(n5808), .A2(n3707), .ZN(n3510) );
  NAND2_X1 U3899 ( .A1(n3510), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3132) );
  NAND2_X1 U3900 ( .A1(n3270), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3131)
         );
  NAND2_X1 U3901 ( .A1(n3501), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3130) );
  INV_X1 U3902 ( .A(n3502), .ZN(n3282) );
  NAND2_X1 U3903 ( .A1(n3282), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3129) );
  INV_X1 U3904 ( .A(n3241), .ZN(n3134) );
  NAND2_X1 U3905 ( .A1(n3241), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3138)
         );
  AND2_X2 U3906 ( .A1(n5800), .A2(n3705), .ZN(n3496) );
  NAND2_X1 U3907 ( .A1(n4949), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3137)
         );
  AND2_X2 U3908 ( .A1(n3704), .A2(n5800), .ZN(n3495) );
  NAND2_X1 U3909 ( .A1(n3495), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3136) );
  NAND2_X1 U3910 ( .A1(n3518), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3135)
         );
  NAND4_X4 U3911 ( .A1(n3142), .A2(n3141), .A3(n3140), .A4(n3139), .ZN(n3538)
         );
  NAND2_X1 U3912 ( .A1(n3511), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3146)
         );
  NAND2_X1 U3913 ( .A1(n5634), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3145) );
  NAND2_X1 U3914 ( .A1(n3254), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3144) );
  NAND2_X1 U3915 ( .A1(n3518), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3143)
         );
  NAND2_X1 U3916 ( .A1(n3268), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3150) );
  NAND2_X1 U3917 ( .A1(n3510), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3149) );
  NAND2_X1 U3918 ( .A1(n3241), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3148)
         );
  NAND2_X1 U3919 ( .A1(n3255), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3147) );
  NAND2_X1 U3920 ( .A1(n5080), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3154)
         );
  NAND2_X1 U3921 ( .A1(n3270), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3153)
         );
  NAND2_X1 U3922 ( .A1(n3269), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3152) );
  NAND2_X1 U3923 ( .A1(n3501), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3151) );
  NAND2_X1 U3924 ( .A1(n3517), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3158) );
  NAND2_X1 U3925 ( .A1(n3248), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3157) );
  NAND2_X1 U3926 ( .A1(n4949), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3156)
         );
  NAND2_X1 U3927 ( .A1(n3495), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3155) );
  CLKBUF_X3 U3928 ( .A(n3645), .Z(n5185) );
  AOI22_X1 U3929 ( .A1(n3248), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3166) );
  AOI22_X1 U3930 ( .A1(n3511), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3517), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3165) );
  AOI22_X1 U3931 ( .A1(n3495), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3496), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3164) );
  AOI22_X1 U3932 ( .A1(n3241), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3163) );
  NAND4_X1 U3933 ( .A1(n3166), .A2(n3165), .A3(n3164), .A4(n3163), .ZN(n3172)
         );
  AOI22_X1 U3934 ( .A1(n3267), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3170) );
  AOI22_X1 U3935 ( .A1(n3268), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3169) );
  AOI22_X1 U3936 ( .A1(n3510), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3501), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3168) );
  AOI22_X1 U3937 ( .A1(n3270), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3255), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3167) );
  NAND4_X1 U3938 ( .A1(n3170), .A2(n3169), .A3(n3168), .A4(n3167), .ZN(n3171)
         );
  AOI22_X1 U3939 ( .A1(n3248), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3517), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3176) );
  AOI22_X1 U3940 ( .A1(n3511), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3241), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3175) );
  AOI22_X1 U3941 ( .A1(n3510), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3174) );
  AOI22_X1 U3942 ( .A1(n3501), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3255), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3173) );
  NAND4_X1 U3943 ( .A1(n3176), .A2(n3175), .A3(n3174), .A4(n3173), .ZN(n3182)
         );
  AOI22_X1 U3944 ( .A1(n3270), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3180) );
  AOI22_X1 U3945 ( .A1(n3267), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3179) );
  AOI22_X1 U3946 ( .A1(n3249), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3495), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3178) );
  AOI22_X1 U3947 ( .A1(n3254), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3496), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3177) );
  NAND4_X1 U3948 ( .A1(n3180), .A2(n3179), .A3(n3178), .A4(n3177), .ZN(n3181)
         );
  OR2_X2 U3949 ( .A1(n3182), .A2(n3181), .ZN(n3747) );
  INV_X2 U3950 ( .A(n3747), .ZN(n4788) );
  AOI21_X1 U3951 ( .B1(n4443), .B2(n3646), .A(n4788), .ZN(n3197) );
  NAND2_X1 U3952 ( .A1(n3197), .A2(n3198), .ZN(n3187) );
  NAND2_X1 U3953 ( .A1(n3795), .A2(n3747), .ZN(n3353) );
  OAI21_X1 U3954 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6927), .A(n3183), 
        .ZN(n3184) );
  INV_X1 U3955 ( .A(n3184), .ZN(n3188) );
  AOI21_X1 U3956 ( .B1(n3353), .B2(n3188), .A(n3189), .ZN(n3185) );
  AOI21_X1 U3957 ( .B1(n4788), .B2(n5185), .A(n3646), .ZN(n3206) );
  OR2_X1 U3958 ( .A1(n3185), .A2(n3206), .ZN(n3186) );
  NAND2_X1 U3959 ( .A1(n3187), .A2(n3186), .ZN(n3192) );
  INV_X1 U3960 ( .A(n3192), .ZN(n3195) );
  INV_X1 U3961 ( .A(n3305), .ZN(n3194) );
  NAND2_X1 U3962 ( .A1(n4443), .A2(n3188), .ZN(n3191) );
  AND2_X4 U3963 ( .A1(n3190), .A2(n3538), .ZN(n4146) );
  NAND2_X1 U3964 ( .A1(n4146), .A2(n4448), .ZN(n3231) );
  OAI21_X1 U3965 ( .B1(n3192), .B2(n3191), .A(n3231), .ZN(n3193) );
  OAI21_X1 U3966 ( .B1(n3195), .B2(n3194), .A(n3193), .ZN(n3196) );
  OAI21_X1 U3967 ( .B1(n3198), .B2(n3197), .A(n3196), .ZN(n3205) );
  NAND2_X1 U3968 ( .A1(n3200), .A2(n3199), .ZN(n3201) );
  OAI21_X1 U3969 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6872), .A(n3201), 
        .ZN(n3211) );
  INV_X1 U3970 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3423) );
  XNOR2_X1 U3971 ( .A(n3423), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3209)
         );
  XNOR2_X1 U3972 ( .A(n3211), .B(n3209), .ZN(n3304) );
  INV_X1 U3973 ( .A(n3206), .ZN(n3203) );
  NAND2_X1 U3974 ( .A1(n4443), .A2(n3304), .ZN(n3202) );
  OAI211_X1 U3975 ( .C1(n4446), .C2(n3304), .A(n3203), .B(n3202), .ZN(n3204)
         );
  NAND2_X1 U3976 ( .A1(n3205), .A2(n3204), .ZN(n3208) );
  NAND3_X1 U3977 ( .A1(n3206), .A2(n4443), .A3(n3304), .ZN(n3207) );
  NAND2_X1 U3978 ( .A1(n3208), .A2(n3207), .ZN(n3226) );
  INV_X1 U3979 ( .A(n3209), .ZN(n3210) );
  NAND2_X1 U3980 ( .A1(n3211), .A2(n3210), .ZN(n3213) );
  INV_X1 U3981 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6560) );
  NAND2_X1 U3982 ( .A1(n6560), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3212) );
  NAND2_X1 U3983 ( .A1(n3213), .A2(n3212), .ZN(n3218) );
  XNOR2_X1 U3984 ( .A(n3214), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3216)
         );
  XNOR2_X1 U3985 ( .A(n3218), .B(n3216), .ZN(n3303) );
  INV_X1 U3986 ( .A(n3303), .ZN(n3215) );
  NAND2_X1 U3987 ( .A1(n3215), .A2(n4446), .ZN(n3225) );
  INV_X1 U3988 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U3989 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6083), .ZN(n3229) );
  NOR2_X1 U3990 ( .A1(n4460), .A2(n3229), .ZN(n3222) );
  INV_X1 U3991 ( .A(n3216), .ZN(n3217) );
  NAND2_X1 U3992 ( .A1(n3218), .A2(n3217), .ZN(n3220) );
  INV_X1 U3993 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6674) );
  NAND2_X1 U3994 ( .A1(n6674), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3219) );
  NAND2_X1 U3995 ( .A1(n3220), .A2(n3219), .ZN(n3230) );
  INV_X1 U3996 ( .A(n3230), .ZN(n3221) );
  AOI22_X1 U3997 ( .A1(n3222), .A2(n3221), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6580), .ZN(n3223) );
  OAI21_X1 U3998 ( .B1(n3231), .B2(n3303), .A(n3223), .ZN(n3224) );
  AOI21_X1 U3999 ( .B1(n3226), .B2(n3225), .A(n3224), .ZN(n3233) );
  INV_X1 U4000 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6438) );
  AND2_X1 U4001 ( .A1(n6438), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3227)
         );
  OR2_X1 U4002 ( .A1(n3230), .A2(n3227), .ZN(n3228) );
  NAND2_X1 U4003 ( .A1(n3228), .A2(n3229), .ZN(n3306) );
  OR2_X1 U4004 ( .A1(n3230), .A2(n3229), .ZN(n3302) );
  OAI22_X1 U4005 ( .A1(n3231), .A2(n3306), .B1(n3302), .B2(n4146), .ZN(n3232)
         );
  INV_X1 U4006 ( .A(n3306), .ZN(n3234) );
  NAND2_X1 U4007 ( .A1(n3234), .A2(n4443), .ZN(n3235) );
  INV_X1 U4008 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5806) );
  AND2_X1 U4009 ( .A1(n5806), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3586) );
  NAND2_X1 U4010 ( .A1(n3586), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6587) );
  AOI22_X1 U4011 ( .A1(n3267), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3240) );
  AOI22_X1 U4012 ( .A1(n3268), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3239) );
  AOI22_X1 U4013 ( .A1(n3510), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3501), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3238) );
  AOI22_X1 U4014 ( .A1(n3270), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3255), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3237) );
  NAND4_X1 U4015 ( .A1(n3240), .A2(n3239), .A3(n3238), .A4(n3237), .ZN(n3247)
         );
  AOI22_X1 U4016 ( .A1(n3248), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3245) );
  AOI22_X1 U4017 ( .A1(n3511), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3517), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3244) );
  AOI22_X1 U4018 ( .A1(n3495), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3496), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3243) );
  AOI22_X1 U4019 ( .A1(n3241), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3242) );
  NAND4_X1 U4020 ( .A1(n3245), .A2(n3244), .A3(n3243), .A4(n3242), .ZN(n3246)
         );
  OR2_X2 U4021 ( .A1(n3247), .A2(n3246), .ZN(n3585) );
  NAND2_X1 U4022 ( .A1(n4788), .A2(n3585), .ZN(n3262) );
  AOI22_X1 U4023 ( .A1(n3248), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U4024 ( .A1(n3511), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3517), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3252) );
  AOI22_X1 U4025 ( .A1(n3495), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3496), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3251) );
  AOI22_X1 U4026 ( .A1(n3241), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3250) );
  NAND4_X1 U4027 ( .A1(n3253), .A2(n3252), .A3(n3251), .A4(n3250), .ZN(n3261)
         );
  AOI22_X1 U4029 ( .A1(n5681), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3259) );
  AOI22_X1 U4030 ( .A1(n4728), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5619), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3258) );
  AOI22_X1 U4031 ( .A1(n3510), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3501), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4032 ( .A1(n3270), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3255), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3256) );
  NAND4_X1 U4033 ( .A1(n3259), .A2(n3258), .A3(n3257), .A4(n3256), .ZN(n3260)
         );
  OR2_X2 U4034 ( .A1(n3261), .A2(n3260), .ZN(n4787) );
  AOI22_X1 U4035 ( .A1(n4496), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n5634), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3266) );
  AOI22_X1 U4036 ( .A1(n3511), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3517), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3265) );
  AOI22_X1 U4037 ( .A1(n3495), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4949), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3264) );
  AOI22_X1 U4038 ( .A1(n3241), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3263) );
  NAND4_X1 U4039 ( .A1(n3266), .A2(n3265), .A3(n3264), .A4(n3263), .ZN(n3276)
         );
  BUF_X2 U4040 ( .A(n3267), .Z(n5620) );
  AOI22_X1 U4041 ( .A1(n5620), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3254), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3274) );
  BUF_X4 U4042 ( .A(n3268), .Z(n5680) );
  AOI22_X1 U4043 ( .A1(n5680), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5619), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3273) );
  AOI22_X1 U4044 ( .A1(n3510), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3501), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3272) );
  AOI22_X1 U4045 ( .A1(n3270), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3255), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3271) );
  NAND4_X1 U4046 ( .A1(n3274), .A2(n3273), .A3(n3272), .A4(n3271), .ZN(n3275)
         );
  OR2_X2 U4047 ( .A1(n3276), .A2(n3275), .ZN(n3370) );
  INV_X2 U4048 ( .A(n3585), .ZN(n3919) );
  NAND2_X2 U4049 ( .A1(n3919), .A2(n3747), .ZN(n5801) );
  NAND2_X1 U4050 ( .A1(n5801), .A2(n3538), .ZN(n3277) );
  NAND3_X1 U4051 ( .A1(n3322), .A2(n3370), .A3(n3277), .ZN(n3375) );
  NAND2_X1 U4052 ( .A1(n4496), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3281) );
  NAND2_X1 U4053 ( .A1(n5634), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3280) );
  NAND2_X1 U4054 ( .A1(n3254), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3279) );
  NAND2_X1 U4055 ( .A1(n3511), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3278)
         );
  NAND2_X1 U4056 ( .A1(n3510), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3286) );
  NAND2_X1 U4057 ( .A1(n3270), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3285)
         );
  NAND2_X1 U4058 ( .A1(n4728), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3284) );
  NAND2_X1 U4059 ( .A1(n3282), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3283) );
  NAND2_X1 U4060 ( .A1(n3517), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3290) );
  NAND2_X1 U4061 ( .A1(n3241), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3289)
         );
  NAND2_X1 U4062 ( .A1(n3495), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3288) );
  NAND2_X1 U4063 ( .A1(n4949), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3287)
         );
  NAND2_X1 U4064 ( .A1(n5080), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3294)
         );
  NAND2_X1 U4065 ( .A1(n3501), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3293) );
  NAND2_X1 U4066 ( .A1(n5619), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3292) );
  NAND2_X1 U4067 ( .A1(n3518), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3291)
         );
  AND4_X2 U4068 ( .A1(n3298), .A2(n3297), .A3(n3296), .A4(n3295), .ZN(n3852)
         );
  NAND2_X1 U4069 ( .A1(n4788), .A2(n3852), .ZN(n3346) );
  OR2_X2 U4070 ( .A1(n3375), .A2(n3346), .ZN(n3481) );
  INV_X2 U4071 ( .A(n3481), .ZN(n3408) );
  NAND2_X2 U4072 ( .A1(n3408), .A2(n5185), .ZN(n3534) );
  NOR2_X1 U4073 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5118) );
  NAND2_X1 U4074 ( .A1(n6445), .A2(n5806), .ZN(n3299) );
  NAND2_X1 U4075 ( .A1(n3313), .A2(n3299), .ZN(n5959) );
  OR2_X2 U4076 ( .A1(n3300), .A2(n3538), .ZN(n3352) );
  NAND2_X1 U4077 ( .A1(n3919), .A2(n4787), .ZN(n3576) );
  INV_X2 U4078 ( .A(n3852), .ZN(n3474) );
  NAND2_X1 U4079 ( .A1(n3576), .A2(n3474), .ZN(n3301) );
  NOR2_X1 U4080 ( .A1(n3370), .A2(n5185), .ZN(n3373) );
  NAND2_X2 U4081 ( .A1(n3350), .A2(n3373), .ZN(n3400) );
  NAND4_X1 U4082 ( .A1(n3305), .A2(n3304), .A3(n3303), .A4(n3302), .ZN(n3307)
         );
  NAND2_X1 U4083 ( .A1(n3307), .A2(n3306), .ZN(n3413) );
  NOR2_X1 U4084 ( .A1(n3400), .A2(n3413), .ZN(n3319) );
  INV_X1 U4085 ( .A(n6587), .ZN(n3590) );
  NAND2_X1 U4086 ( .A1(n3319), .A2(n3590), .ZN(n5960) );
  INV_X1 U4087 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n3308) );
  NAND2_X1 U4088 ( .A1(n5960), .A2(n3308), .ZN(n3311) );
  AND2_X2 U4089 ( .A1(n3790), .A2(n3645), .ZN(n5182) );
  NAND2_X1 U4090 ( .A1(n3785), .A2(n3646), .ZN(n5176) );
  INV_X1 U4091 ( .A(n5176), .ZN(n3309) );
  OR2_X1 U4092 ( .A1(n5182), .A2(n3309), .ZN(n3320) );
  NAND2_X1 U4093 ( .A1(n6686), .A2(n3320), .ZN(n3310) );
  OAI21_X1 U4094 ( .B1(n5959), .B2(n3311), .A(n3310), .ZN(n3312) );
  INV_X1 U4095 ( .A(n3312), .ZN(U3474) );
  NAND2_X1 U4096 ( .A1(n3408), .A2(n5182), .ZN(n6576) );
  OR2_X1 U4097 ( .A1(n3739), .A2(n6576), .ZN(n6313) );
  INV_X1 U4098 ( .A(EAX_REG_15__SCAN_IN), .ZN(n3318) );
  INV_X1 U4099 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n3317) );
  INV_X1 U4100 ( .A(n3313), .ZN(n3316) );
  INV_X1 U4101 ( .A(n5182), .ZN(n6691) );
  NAND2_X1 U4102 ( .A1(n6691), .A2(READY_N), .ZN(n3314) );
  AND2_X1 U4103 ( .A1(n3316), .A2(n3314), .ZN(n3429) );
  INV_X1 U4104 ( .A(READY_N), .ZN(n6688) );
  AND2_X1 U4105 ( .A1(n3646), .A2(n6688), .ZN(n3315) );
  INV_X1 U4106 ( .A(DATAI_15_), .ZN(n6766) );
  OAI222_X1 U4107 ( .A1(n6313), .A2(n3318), .B1(n3317), .B2(n3429), .C1(n6298), 
        .C2(n6766), .ZN(U2954) );
  INV_X1 U4108 ( .A(n3643), .ZN(n3410) );
  NOR2_X1 U4109 ( .A1(n5185), .A2(n3646), .ZN(n5169) );
  INV_X1 U4110 ( .A(n3534), .ZN(n3330) );
  OAI22_X1 U4111 ( .A1(n3410), .A2(n5169), .B1(n3330), .B2(n3319), .ZN(n6086)
         );
  INV_X1 U4112 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6602) );
  XNOR2_X1 U4113 ( .A(n6602), .B(STATE_REG_2__SCAN_IN), .ZN(n3339) );
  INV_X1 U4114 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6603) );
  NAND2_X1 U4115 ( .A1(n3339), .A2(n6603), .ZN(n6601) );
  AOI21_X1 U4116 ( .B1(n3320), .B2(n6601), .A(READY_N), .ZN(n6690) );
  NOR2_X1 U4117 ( .A1(n6086), .A2(n6690), .ZN(n6565) );
  OR2_X1 U4118 ( .A1(n6565), .A2(n6587), .ZN(n6092) );
  INV_X1 U4119 ( .A(n6092), .ZN(n3337) );
  INV_X1 U4120 ( .A(MORE_REG_SCAN_IN), .ZN(n3336) );
  OR2_X1 U4121 ( .A1(n5801), .A2(n3538), .ZN(n3321) );
  NAND2_X1 U4122 ( .A1(n3322), .A2(n3321), .ZN(n3388) );
  NAND2_X1 U4123 ( .A1(n3852), .A2(n3370), .ZN(n3746) );
  NAND2_X1 U4124 ( .A1(n5801), .A2(n3785), .ZN(n3323) );
  AND2_X1 U4125 ( .A1(n3358), .A2(n3323), .ZN(n3329) );
  NAND2_X1 U4126 ( .A1(n4448), .A2(n3919), .ZN(n3325) );
  OAI211_X1 U4127 ( .C1(n3352), .C2(n3472), .A(n5185), .B(n3325), .ZN(n3393)
         );
  NAND2_X1 U4128 ( .A1(n3329), .A2(n3393), .ZN(n3324) );
  NAND2_X1 U4129 ( .A1(n3324), .A2(n3400), .ZN(n3477) );
  OR2_X1 U4130 ( .A1(n5176), .A2(n3474), .ZN(n3415) );
  INV_X1 U4131 ( .A(n3325), .ZN(n3326) );
  AND2_X1 U4132 ( .A1(n3415), .A2(n3326), .ZN(n3327) );
  NAND2_X1 U4133 ( .A1(n3477), .A2(n3327), .ZN(n3641) );
  INV_X1 U4134 ( .A(n3641), .ZN(n3489) );
  NAND2_X1 U4135 ( .A1(n3329), .A2(n5169), .ZN(n3593) );
  INV_X1 U4136 ( .A(n3593), .ZN(n3412) );
  INV_X1 U4137 ( .A(n3353), .ZN(n3328) );
  NAND2_X1 U4138 ( .A1(n3329), .A2(n3328), .ZN(n6566) );
  INV_X1 U4139 ( .A(n6566), .ZN(n3331) );
  NOR3_X1 U4140 ( .A1(n3412), .A2(n3331), .A3(n3330), .ZN(n3333) );
  INV_X1 U4141 ( .A(n3413), .ZN(n3332) );
  OAI22_X1 U4142 ( .A1(n3410), .A2(n3333), .B1(n3332), .B2(n3400), .ZN(n3334)
         );
  AOI21_X1 U4143 ( .B1(n3410), .B2(n3489), .A(n3334), .ZN(n6567) );
  OR2_X1 U4144 ( .A1(n6092), .A2(n6567), .ZN(n3335) );
  OAI21_X1 U4145 ( .B1(n3337), .B2(n3336), .A(n3335), .ZN(U3471) );
  NOR2_X1 U4146 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6079) );
  NAND2_X1 U4147 ( .A1(n6079), .A2(n6580), .ZN(n3766) );
  INV_X1 U4148 ( .A(n3766), .ZN(n3677) );
  XNOR2_X1 U4149 ( .A(n6927), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5282)
         );
  INV_X1 U4150 ( .A(n3586), .ZN(n3676) );
  AND2_X1 U4151 ( .A1(n3676), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3338)
         );
  AOI21_X1 U4152 ( .B1(n3677), .B2(n5282), .A(n3338), .ZN(n3361) );
  INV_X1 U4153 ( .A(n3361), .ZN(n3343) );
  OR2_X2 U4154 ( .A1(n3400), .A2(n3646), .ZN(n3725) );
  NOR2_X1 U4155 ( .A1(n3646), .A2(n3339), .ZN(n3355) );
  INV_X1 U4156 ( .A(n3346), .ZN(n3340) );
  INV_X1 U4157 ( .A(n3370), .ZN(n3799) );
  NAND2_X1 U4158 ( .A1(n3589), .A2(n3571), .ZN(n3539) );
  INV_X1 U4159 ( .A(n3360), .ZN(n3342) );
  OAI21_X1 U4160 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n3343), .A(n3342), 
        .ZN(n3362) );
  INV_X2 U4161 ( .A(n3571), .ZN(n4786) );
  OAI211_X1 U4162 ( .C1(n3346), .C2(n4786), .A(n3372), .B(n3785), .ZN(n3349)
         );
  NAND2_X1 U4163 ( .A1(n3785), .A2(n3370), .ZN(n3759) );
  INV_X1 U4164 ( .A(n3347), .ZN(n3348) );
  INV_X1 U4165 ( .A(n3351), .ZN(n3366) );
  NAND2_X1 U4166 ( .A1(n3352), .A2(n5182), .ZN(n3354) );
  INV_X1 U4167 ( .A(n3355), .ZN(n3356) );
  AOI22_X1 U4168 ( .A1(n4146), .A2(n5801), .B1(n3356), .B2(n4788), .ZN(n3357)
         );
  NAND4_X1 U4169 ( .A1(n3366), .A2(n3378), .A3(n3358), .A4(n3357), .ZN(n3359)
         );
  OAI211_X1 U4170 ( .C1(n3363), .C2(n6872), .A(n3361), .B(n3360), .ZN(n3381)
         );
  NAND2_X1 U4171 ( .A1(n3362), .A2(n3381), .ZN(n3553) );
  INV_X1 U4172 ( .A(n3553), .ZN(n3380) );
  OR2_X2 U4173 ( .A1(n3363), .A2(n3468), .ZN(n3365) );
  MUX2_X1 U4174 ( .A(n3586), .B(n3766), .S(n6927), .Z(n3364) );
  INV_X1 U4175 ( .A(n3366), .ZN(n3367) );
  NAND2_X1 U4176 ( .A1(n4448), .A2(n3795), .ZN(n3487) );
  NAND2_X1 U4177 ( .A1(n3367), .A2(n3487), .ZN(n3369) );
  NAND2_X1 U4178 ( .A1(n3474), .A2(n5185), .ZN(n3368) );
  NAND2_X1 U4179 ( .A1(n3369), .A2(n3368), .ZN(n3395) );
  NAND2_X1 U4180 ( .A1(n5801), .A2(n3370), .ZN(n3371) );
  NAND2_X1 U4181 ( .A1(n6079), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6588) );
  AOI21_X1 U4182 ( .B1(n3371), .B2(n5182), .A(n6588), .ZN(n3377) );
  INV_X1 U4183 ( .A(n3372), .ZN(n3374) );
  NAND2_X1 U4184 ( .A1(n3374), .A2(n3373), .ZN(n3714) );
  NAND2_X1 U4185 ( .A1(n3375), .A2(n3646), .ZN(n3376) );
  NAND4_X1 U4186 ( .A1(n3378), .A2(n3377), .A3(n3714), .A4(n3376), .ZN(n3379)
         );
  NAND2_X1 U4187 ( .A1(n3380), .A2(n3552), .ZN(n3382) );
  NAND2_X1 U4188 ( .A1(n3382), .A2(n3381), .ZN(n3672) );
  AND2_X1 U4189 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3383) );
  NAND2_X1 U4190 ( .A1(n3383), .A2(n6560), .ZN(n6486) );
  INV_X1 U4191 ( .A(n3383), .ZN(n3384) );
  NAND2_X1 U4192 ( .A1(n3384), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3385) );
  NAND2_X1 U4193 ( .A1(n6486), .A2(n3385), .ZN(n4023) );
  AOI22_X1 U4194 ( .A1(n3677), .A2(n4023), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3676), .ZN(n3386) );
  XNOR2_X2 U4195 ( .A(n3672), .B(n3673), .ZN(n4068) );
  INV_X1 U4196 ( .A(n4068), .ZN(n5951) );
  INV_X1 U4197 ( .A(n4155), .ZN(n5769) );
  AOI22_X1 U4198 ( .A1(n3388), .A2(n5769), .B1(n3474), .B2(n4786), .ZN(n3392)
         );
  INV_X1 U4199 ( .A(n5774), .ZN(n3389) );
  NAND2_X1 U4200 ( .A1(n3389), .A2(n3415), .ZN(n3390) );
  NAND2_X1 U4201 ( .A1(n3390), .A2(n3746), .ZN(n3391) );
  NAND3_X1 U4202 ( .A1(n3393), .A2(n3392), .A3(n3391), .ZN(n3394) );
  NOR2_X1 U4203 ( .A1(n3395), .A2(n3394), .ZN(n3486) );
  INV_X1 U4204 ( .A(n3589), .ZN(n3396) );
  AND4_X1 U4205 ( .A1(n3725), .A2(n3397), .A3(n3481), .A4(n3396), .ZN(n3398)
         );
  AND2_X1 U4206 ( .A1(n3486), .A2(n3398), .ZN(n5805) );
  NAND2_X1 U4207 ( .A1(n3641), .A2(n3593), .ZN(n3717) );
  XNOR2_X1 U4208 ( .A(n3399), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3403)
         );
  NOR2_X1 U4209 ( .A1(n3400), .A2(n3790), .ZN(n5803) );
  INV_X1 U4210 ( .A(n5803), .ZN(n3457) );
  XNOR2_X1 U4211 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3401) );
  OAI22_X1 U4212 ( .A1(n3457), .A2(n3401), .B1(n3714), .B2(n3403), .ZN(n3402)
         );
  AOI21_X1 U4213 ( .B1(n3717), .B2(n3403), .A(n3402), .ZN(n3404) );
  OAI21_X1 U4214 ( .B1(n5951), .B2(n5805), .A(n3404), .ZN(n3701) );
  INV_X1 U4215 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6431) );
  INV_X1 U4216 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n6859) );
  AOI22_X1 U4217 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6859), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n3858), .ZN(n5810) );
  NOR3_X1 U4218 ( .A1(n5806), .A2(n6431), .A3(n5810), .ZN(n3406) );
  INV_X1 U4219 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6826) );
  INV_X1 U4220 ( .A(n3399), .ZN(n3422) );
  NOR3_X1 U4221 ( .A1(n6581), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n3422), 
        .ZN(n3405) );
  AOI211_X1 U4222 ( .C1(n3701), .C2(n6079), .A(n3406), .B(n3405), .ZN(n3425)
         );
  NAND2_X1 U4223 ( .A1(n3790), .A2(n6601), .ZN(n5174) );
  NAND2_X1 U4224 ( .A1(n5174), .A2(n6688), .ZN(n3480) );
  AOI21_X1 U4225 ( .B1(n3534), .B2(n6601), .A(n3480), .ZN(n3407) );
  OAI21_X1 U4226 ( .B1(n5803), .B2(n3408), .A(n3407), .ZN(n3409) );
  INV_X1 U4227 ( .A(n3409), .ZN(n3411) );
  OAI21_X1 U4228 ( .B1(n3412), .B2(n3411), .A(n3410), .ZN(n3419) );
  NOR2_X1 U4229 ( .A1(READY_N), .A2(n3413), .ZN(n3473) );
  INV_X1 U4230 ( .A(n3473), .ZN(n3414) );
  NOR2_X1 U4231 ( .A1(n3725), .A2(n3414), .ZN(n3591) );
  NAND2_X1 U4232 ( .A1(n3477), .A2(n3415), .ZN(n3416) );
  OR2_X1 U4233 ( .A1(n3591), .A2(n3416), .ZN(n3417) );
  AOI21_X1 U4234 ( .B1(n3643), .B2(n3489), .A(n3417), .ZN(n3418) );
  OR2_X1 U4235 ( .A1(n3727), .A2(n6587), .ZN(n3421) );
  NAND2_X1 U4236 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n3735) );
  NOR2_X1 U4237 ( .A1(n6580), .A2(n3735), .ZN(n3733) );
  NAND2_X1 U4238 ( .A1(FLUSH_REG_SCAN_IN), .A2(n3733), .ZN(n3420) );
  AND2_X1 U4239 ( .A1(n3421), .A2(n3420), .ZN(n6078) );
  OAI21_X1 U4240 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6826), .A(n6078), .ZN(
        n6084) );
  INV_X1 U4241 ( .A(n6084), .ZN(n5812) );
  AOI21_X1 U4242 ( .B1(n5807), .B2(n3422), .A(n5812), .ZN(n3424) );
  OAI22_X1 U4243 ( .A1(n3425), .A2(n5812), .B1(n3424), .B2(n3423), .ZN(U3459)
         );
  AOI22_X1 U4244 ( .A1(n6699), .A2(UWORD_REG_8__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n3426) );
  INV_X1 U4245 ( .A(n6298), .ZN(n6305) );
  NAND2_X1 U4246 ( .A1(n6305), .A2(DATAI_8_), .ZN(n3448) );
  NAND2_X1 U4247 ( .A1(n3426), .A2(n3448), .ZN(U2932) );
  AOI22_X1 U4248 ( .A1(n6699), .A2(UWORD_REG_7__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n3427) );
  INV_X1 U4249 ( .A(DATAI_7_), .ZN(n3780) );
  OR2_X1 U4250 ( .A1(n6298), .A2(n3780), .ZN(n3432) );
  NAND2_X1 U4251 ( .A1(n3427), .A2(n3432), .ZN(U2931) );
  AOI22_X1 U4252 ( .A1(n6699), .A2(LWORD_REG_3__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_3__SCAN_IN), .ZN(n3428) );
  NAND2_X1 U4253 ( .A1(n6305), .A2(DATAI_3_), .ZN(n3435) );
  NAND2_X1 U4254 ( .A1(n3428), .A2(n3435), .ZN(U2942) );
  INV_X2 U4255 ( .A(n3429), .ZN(n6699) );
  AOI22_X1 U4256 ( .A1(n6699), .A2(LWORD_REG_13__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n3430) );
  NAND2_X1 U4257 ( .A1(n6305), .A2(DATAI_13_), .ZN(n3453) );
  NAND2_X1 U4258 ( .A1(n3430), .A2(n3453), .ZN(U2952) );
  AOI22_X1 U4259 ( .A1(n6699), .A2(LWORD_REG_2__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n3431) );
  NAND2_X1 U4260 ( .A1(n6305), .A2(DATAI_2_), .ZN(n3443) );
  NAND2_X1 U4261 ( .A1(n3431), .A2(n3443), .ZN(U2941) );
  AOI22_X1 U4262 ( .A1(n6699), .A2(LWORD_REG_7__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n3433) );
  NAND2_X1 U4263 ( .A1(n3433), .A2(n3432), .ZN(U2946) );
  AOI22_X1 U4264 ( .A1(n6699), .A2(UWORD_REG_5__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n3434) );
  INV_X1 U4265 ( .A(DATAI_5_), .ZN(n3926) );
  OR2_X1 U4266 ( .A1(n6298), .A2(n3926), .ZN(n3438) );
  NAND2_X1 U4267 ( .A1(n3434), .A2(n3438), .ZN(U2929) );
  AOI22_X1 U4268 ( .A1(n6699), .A2(UWORD_REG_3__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n3436) );
  NAND2_X1 U4269 ( .A1(n3436), .A2(n3435), .ZN(U2927) );
  AOI22_X1 U4270 ( .A1(n6699), .A2(UWORD_REG_4__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n3437) );
  NAND2_X1 U4271 ( .A1(n6305), .A2(DATAI_4_), .ZN(n3445) );
  NAND2_X1 U4272 ( .A1(n3437), .A2(n3445), .ZN(U2928) );
  AOI22_X1 U4273 ( .A1(n6699), .A2(LWORD_REG_5__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n3439) );
  NAND2_X1 U4274 ( .A1(n3439), .A2(n3438), .ZN(U2944) );
  AOI22_X1 U4275 ( .A1(n6699), .A2(UWORD_REG_6__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n3440) );
  OR2_X1 U4276 ( .A1(n6298), .A2(n4227), .ZN(n3441) );
  NAND2_X1 U4277 ( .A1(n3440), .A2(n3441), .ZN(U2930) );
  AOI22_X1 U4278 ( .A1(n6699), .A2(LWORD_REG_6__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n3442) );
  NAND2_X1 U4279 ( .A1(n3442), .A2(n3441), .ZN(U2945) );
  AOI22_X1 U4280 ( .A1(n6699), .A2(UWORD_REG_2__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n3444) );
  NAND2_X1 U4281 ( .A1(n3444), .A2(n3443), .ZN(U2926) );
  AOI22_X1 U4282 ( .A1(n6699), .A2(LWORD_REG_4__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n3446) );
  NAND2_X1 U4283 ( .A1(n3446), .A2(n3445), .ZN(U2943) );
  AOI22_X1 U4284 ( .A1(n6699), .A2(UWORD_REG_0__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n3447) );
  NAND2_X1 U4285 ( .A1(n6305), .A2(DATAI_0_), .ZN(n3451) );
  NAND2_X1 U4286 ( .A1(n3447), .A2(n3451), .ZN(U2924) );
  AOI22_X1 U4287 ( .A1(n6699), .A2(LWORD_REG_8__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n3449) );
  NAND2_X1 U4288 ( .A1(n3449), .A2(n3448), .ZN(U2947) );
  AOI22_X1 U4289 ( .A1(n6699), .A2(LWORD_REG_1__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n3450) );
  NAND2_X1 U4290 ( .A1(n6305), .A2(DATAI_1_), .ZN(n3455) );
  NAND2_X1 U4291 ( .A1(n3450), .A2(n3455), .ZN(U2940) );
  AOI22_X1 U4292 ( .A1(n6699), .A2(LWORD_REG_0__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_0__SCAN_IN), .ZN(n3452) );
  NAND2_X1 U4293 ( .A1(n3452), .A2(n3451), .ZN(U2939) );
  AOI22_X1 U4294 ( .A1(n6699), .A2(UWORD_REG_13__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n3454) );
  NAND2_X1 U4295 ( .A1(n3454), .A2(n3453), .ZN(U2937) );
  AOI22_X1 U4296 ( .A1(n6699), .A2(UWORD_REG_1__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n3456) );
  NAND2_X1 U4297 ( .A1(n3456), .A2(n3455), .ZN(U2925) );
  INV_X1 U4298 ( .A(EAX_REG_22__SCAN_IN), .ZN(n3462) );
  OR2_X1 U4299 ( .A1(n3739), .A2(n3457), .ZN(n3458) );
  NAND2_X1 U4300 ( .A1(n6313), .A2(n3458), .ZN(n3459) );
  INV_X1 U4301 ( .A(n6601), .ZN(n3475) );
  OR2_X1 U4302 ( .A1(n6285), .A2(n3785), .ZN(n6254) );
  NOR2_X1 U4303 ( .A1(n3735), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6277) );
  INV_X1 U4304 ( .A(n6277), .ZN(n6573) );
  INV_X1 U4305 ( .A(n6573), .ZN(n6689) );
  AOI22_X1 U4306 ( .A1(n6689), .A2(UWORD_REG_6__SCAN_IN), .B1(n6280), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n3461) );
  OAI21_X1 U4307 ( .B1(n3462), .B2(n6254), .A(n3461), .ZN(U2901) );
  INV_X1 U4308 ( .A(EAX_REG_19__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4309 ( .A1(n6689), .A2(UWORD_REG_3__SCAN_IN), .B1(n6280), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n3463) );
  OAI21_X1 U4310 ( .B1(n3464), .B2(n6254), .A(n3463), .ZN(U2904) );
  NAND2_X1 U4311 ( .A1(n5803), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6552) );
  INV_X1 U4312 ( .A(n6079), .ZN(n5956) );
  AOI21_X1 U4313 ( .B1(n5807), .B2(n3468), .A(n5812), .ZN(n5811) );
  INV_X1 U4314 ( .A(n5811), .ZN(n3470) );
  INV_X1 U4315 ( .A(n5805), .ZN(n3703) );
  AOI22_X1 U4316 ( .A1(n3110), .A2(n3703), .B1(n3472), .B2(n3468), .ZN(n6553)
         );
  OAI22_X1 U4317 ( .A1(n6553), .A2(n5956), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n5806), .ZN(n3469) );
  OAI22_X1 U4318 ( .A1(n3470), .A2(n3469), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6084), .ZN(n3471) );
  OAI21_X1 U4319 ( .B1(n6552), .B2(n5956), .A(n3471), .ZN(U3461) );
  NAND3_X1 U4320 ( .A1(n3643), .A2(n3472), .A3(n3646), .ZN(n3478) );
  OAI211_X1 U4321 ( .C1(n3790), .C2(n3475), .A(n3474), .B(n3473), .ZN(n3476)
         );
  NAND3_X1 U4322 ( .A1(n3478), .A2(n3477), .A3(n3476), .ZN(n3479) );
  NAND2_X1 U4323 ( .A1(n3479), .A2(n3590), .ZN(n3485) );
  OAI211_X1 U4324 ( .C1(n3481), .C2(n3480), .A(n5185), .B(n4786), .ZN(n3482)
         );
  NAND2_X1 U4325 ( .A1(n3482), .A2(n3852), .ZN(n3483) );
  OAI211_X1 U4326 ( .C1(n3487), .C2(n3759), .A(n3486), .B(n3714), .ZN(n3488)
         );
  INV_X1 U4327 ( .A(n4164), .ZN(n3490) );
  NAND2_X1 U4328 ( .A1(n3541), .A2(n3489), .ZN(n6416) );
  AND2_X1 U4329 ( .A1(n3490), .A2(n6416), .ZN(n6059) );
  NAND2_X1 U4330 ( .A1(n4164), .A2(n6431), .ZN(n3493) );
  INV_X1 U4331 ( .A(n3541), .ZN(n3491) );
  OR2_X1 U4332 ( .A1(n3766), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6426) );
  NAND2_X1 U4333 ( .A1(n3491), .A2(n6426), .ZN(n3492) );
  AND2_X1 U4334 ( .A1(n3493), .A2(n3492), .ZN(n5223) );
  INV_X1 U4335 ( .A(n5223), .ZN(n4469) );
  AOI21_X1 U4336 ( .B1(n5222), .B2(n6431), .A(n4469), .ZN(n6437) );
  NAND2_X1 U4337 ( .A1(n3541), .A2(n5803), .ZN(n6430) );
  AOI22_X1 U4338 ( .A1(n6059), .A2(n6431), .B1(n6437), .B2(n6430), .ZN(n3547)
         );
  INV_X1 U4339 ( .A(n3516), .ZN(n4995) );
  AOI22_X1 U4340 ( .A1(n4995), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5683), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3500) );
  AOI22_X1 U4341 ( .A1(n3241), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n5629), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3499) );
  AOI22_X1 U4342 ( .A1(n5680), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5692), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3498) );
  AOI22_X1 U4344 ( .A1(n5682), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3497) );
  NAND4_X1 U4345 ( .A1(n3500), .A2(n3499), .A3(n3498), .A4(n3497), .ZN(n3508)
         );
  AOI22_X1 U4346 ( .A1(n5691), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3506) );
  AOI22_X1 U4347 ( .A1(n5688), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3501), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3505) );
  BUF_X1 U4348 ( .A(n3518), .Z(n5635) );
  AOI22_X1 U4349 ( .A1(n5681), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3504) );
  AOI22_X1 U4350 ( .A1(n3608), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3503) );
  NAND4_X1 U4351 ( .A1(n3506), .A2(n3505), .A3(n3504), .A4(n3503), .ZN(n3507)
         );
  INV_X1 U4352 ( .A(n4464), .ZN(n3509) );
  NOR2_X1 U4353 ( .A1(n3509), .A2(n3587), .ZN(n4459) );
  NOR2_X1 U4354 ( .A1(n3587), .A2(n4464), .ZN(n3566) );
  AOI22_X1 U4355 ( .A1(n3241), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n5629), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4356 ( .A1(n5681), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3514) );
  BUF_X1 U4357 ( .A(n3510), .Z(n5688) );
  AOI22_X1 U4358 ( .A1(n5688), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3501), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3513) );
  BUF_X1 U4359 ( .A(n3511), .Z(n5691) );
  AOI22_X1 U4360 ( .A1(n5691), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3512) );
  NAND4_X1 U4361 ( .A1(n3515), .A2(n3514), .A3(n3513), .A4(n3512), .ZN(n3524)
         );
  AOI22_X1 U4362 ( .A1(n4995), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5683), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U4363 ( .A1(n5689), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n5682), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3521) );
  AOI22_X1 U4364 ( .A1(n3608), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3520) );
  AOI22_X1 U4365 ( .A1(n5692), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3519) );
  NAND4_X1 U4366 ( .A1(n3522), .A2(n3521), .A3(n3520), .A4(n3519), .ZN(n3523)
         );
  OR2_X1 U4367 ( .A1(n3524), .A2(n3523), .ZN(n3744) );
  MUX2_X1 U4368 ( .A(n4459), .B(n3566), .S(n3744), .Z(n3549) );
  INV_X1 U4369 ( .A(n3549), .ZN(n3527) );
  INV_X1 U4370 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4048) );
  AOI21_X1 U4371 ( .B1(n3785), .B2(n3744), .A(n6580), .ZN(n3526) );
  NAND2_X1 U4372 ( .A1(n3795), .A2(n4464), .ZN(n3525) );
  OAI211_X1 U4373 ( .C1(n4446), .C2(n4048), .A(n3526), .B(n3525), .ZN(n3548)
         );
  XNOR2_X1 U4374 ( .A(n3527), .B(n3548), .ZN(n3528) );
  NAND2_X1 U4375 ( .A1(n3551), .A2(n3528), .ZN(n5111) );
  OR2_X1 U4376 ( .A1(n5111), .A2(n4460), .ZN(n3531) );
  OAI21_X1 U4377 ( .B1(n6691), .B2(n3744), .A(n3759), .ZN(n3529) );
  INV_X1 U4378 ( .A(n3529), .ZN(n3530) );
  NAND2_X1 U4379 ( .A1(n3531), .A2(n3530), .ZN(n3532) );
  NAND2_X1 U4380 ( .A1(n3532), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3753)
         );
  OAI21_X1 U4381 ( .B1(n3532), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n3753), 
        .ZN(n6357) );
  NAND2_X1 U4382 ( .A1(n3593), .A2(n3725), .ZN(n3536) );
  OR2_X1 U4383 ( .A1(n3539), .A2(n3795), .ZN(n3533) );
  OAI211_X1 U4384 ( .C1(n3534), .C2(n3790), .A(n6566), .B(n3533), .ZN(n3535)
         );
  OR2_X1 U4385 ( .A1(n3536), .A2(n3535), .ZN(n3537) );
  NAND2_X1 U4386 ( .A1(n3541), .A2(n3537), .ZN(n6406) );
  NOR2_X1 U4387 ( .A1(n6357), .A2(n6406), .ZN(n3546) );
  OAI21_X1 U4388 ( .B1(n3539), .B2(n3538), .A(n6576), .ZN(n3540) );
  NAND2_X1 U4389 ( .A1(n5658), .A2(EBX_REG_0__SCAN_IN), .ZN(n3543) );
  INV_X1 U4390 ( .A(EBX_REG_0__SCAN_IN), .ZN(n7001) );
  NAND2_X1 U4391 ( .A1(n4155), .A2(n7001), .ZN(n3542) );
  NAND2_X1 U4392 ( .A1(n3543), .A2(n3542), .ZN(n3864) );
  OAI21_X1 U4393 ( .B1(n5774), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n3864), 
        .ZN(n5178) );
  INV_X1 U4394 ( .A(REIP_REG_0__SCAN_IN), .ZN(n3544) );
  OR2_X1 U4395 ( .A1(n6426), .A2(n3544), .ZN(n6365) );
  OAI21_X1 U4396 ( .B1(n6428), .B2(n5178), .A(n6365), .ZN(n3545) );
  OR3_X1 U4397 ( .A1(n3547), .A2(n3546), .A3(n3545), .ZN(U3018) );
  AOI21_X1 U4398 ( .B1(n3549), .B2(n3548), .A(n4459), .ZN(n3550) );
  XNOR2_X2 U4399 ( .A(n3553), .B(n3552), .ZN(n5948) );
  OR2_X2 U4400 ( .A1(n5948), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3565) );
  INV_X1 U4401 ( .A(n3587), .ZN(n3648) );
  AOI22_X1 U4402 ( .A1(n5683), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3557) );
  AOI22_X1 U4403 ( .A1(n5688), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3556) );
  AOI22_X1 U4404 ( .A1(n5691), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5682), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3555) );
  INV_X1 U4405 ( .A(n3254), .ZN(n3808) );
  AOI22_X1 U4406 ( .A1(n5679), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3554) );
  NAND4_X1 U4407 ( .A1(n3557), .A2(n3556), .A3(n3555), .A4(n3554), .ZN(n3563)
         );
  INV_X1 U4408 ( .A(n3134), .ZN(n4729) );
  AOI22_X1 U4409 ( .A1(n4995), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4729), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4410 ( .A1(n5680), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3501), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4411 ( .A1(n5692), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U4412 ( .A1(n3608), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3558) );
  NAND4_X1 U4413 ( .A1(n3561), .A2(n3560), .A3(n3559), .A4(n3558), .ZN(n3562)
         );
  OR2_X1 U4414 ( .A1(n3563), .A2(n3562), .ZN(n3745) );
  NAND2_X1 U4415 ( .A1(n3648), .A2(n3745), .ZN(n3564) );
  NAND2_X2 U4416 ( .A1(n3565), .A2(n3564), .ZN(n3628) );
  XNOR2_X2 U4417 ( .A(n3626), .B(n3628), .ZN(n3625) );
  INV_X1 U4418 ( .A(n3625), .ZN(n3570) );
  INV_X1 U4419 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4033) );
  INV_X1 U4420 ( .A(n3566), .ZN(n3569) );
  INV_X1 U4421 ( .A(n3567), .ZN(n3621) );
  NAND2_X1 U4422 ( .A1(n3621), .A2(n3745), .ZN(n3568) );
  OAI211_X1 U4423 ( .C1(n4446), .C2(n4033), .A(n3569), .B(n3568), .ZN(n3624)
         );
  XNOR2_X1 U4424 ( .A(n3570), .B(n3624), .ZN(n3743) );
  INV_X2 U4425 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6814) );
  NOR2_X2 U4426 ( .A1(n3585), .A2(n6814), .ZN(n4754) );
  NAND2_X1 U4427 ( .A1(n3743), .A2(n4754), .ZN(n3575) );
  OR2_X1 U4428 ( .A1(n4787), .A2(n6814), .ZN(n4692) );
  INV_X2 U4429 ( .A(n4692), .ZN(n5785) );
  AOI22_X1 U4430 ( .A1(n5785), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6814), .ZN(n3573) );
  AND2_X1 U4431 ( .A1(n3571), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3694) );
  NAND2_X1 U4432 ( .A1(n3694), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3572) );
  AND2_X1 U4433 ( .A1(n3573), .A2(n3572), .ZN(n3574) );
  NAND2_X1 U4434 ( .A1(n3575), .A2(n3574), .ZN(n3584) );
  NAND2_X1 U4435 ( .A1(n5111), .A2(n3345), .ZN(n3598) );
  NAND2_X1 U4436 ( .A1(n3110), .A2(n4754), .ZN(n3580) );
  AOI22_X1 U4437 ( .A1(n5785), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6814), .ZN(n3578) );
  NAND2_X1 U4438 ( .A1(n3694), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3577) );
  AND2_X1 U4439 ( .A1(n3578), .A2(n3577), .ZN(n3579) );
  NAND2_X1 U4440 ( .A1(n3580), .A2(n3579), .ZN(n3600) );
  AND2_X1 U4441 ( .A1(n3600), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3581) );
  NAND2_X1 U4442 ( .A1(n3598), .A2(n3581), .ZN(n3599) );
  INV_X1 U4443 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6091) );
  NAND2_X1 U4444 ( .A1(n6814), .A2(n6091), .ZN(n5703) );
  OR2_X1 U4445 ( .A1(n3600), .A2(n5646), .ZN(n3582) );
  NAND2_X1 U4446 ( .A1(n3599), .A2(n3582), .ZN(n3583) );
  NAND2_X1 U4447 ( .A1(n3584), .A2(n3583), .ZN(n3637) );
  OAI21_X1 U4448 ( .B1(n3584), .B2(n3583), .A(n3637), .ZN(n6230) );
  INV_X1 U4449 ( .A(n4787), .ZN(n5797) );
  NAND3_X1 U4450 ( .A1(n5797), .A2(n3586), .A3(n3585), .ZN(n3644) );
  NOR2_X1 U4451 ( .A1(n3644), .A2(n3587), .ZN(n3588) );
  AOI22_X1 U4452 ( .A1(n3591), .A2(n3590), .B1(n3589), .B2(n3588), .ZN(n3592)
         );
  OAI21_X1 U4453 ( .B1(n3739), .B2(n3593), .A(n3592), .ZN(n3594) );
  INV_X1 U4454 ( .A(n3594), .ZN(n3595) );
  NAND2_X1 U4455 ( .A1(n5801), .A2(n4787), .ZN(n3596) );
  INV_X2 U4456 ( .A(n6248), .ZN(n5862) );
  INV_X1 U4457 ( .A(n3596), .ZN(n3597) );
  NAND2_X1 U4458 ( .A1(n5796), .A2(n3597), .ZN(n5109) );
  INV_X1 U4459 ( .A(DATAI_1_), .ZN(n3791) );
  INV_X1 U4460 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6282) );
  OAI222_X1 U4461 ( .A1(n6230), .A2(n5862), .B1(n5109), .B2(n3791), .C1(n5796), 
        .C2(n6282), .ZN(U2890) );
  AND2_X1 U4462 ( .A1(n3598), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3601) );
  OAI21_X1 U4463 ( .B1(n3601), .B2(n3600), .A(n3599), .ZN(n6356) );
  INV_X1 U4464 ( .A(DATAI_0_), .ZN(n3786) );
  INV_X1 U4465 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6938) );
  OAI222_X1 U4466 ( .A1(n6356), .A2(n5862), .B1(n5109), .B2(n3786), .C1(n5796), 
        .C2(n6938), .ZN(U2891) );
  NAND2_X1 U4467 ( .A1(n3694), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3606) );
  OAI21_X1 U4468 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3695), .ZN(n6347) );
  INV_X1 U4469 ( .A(n6347), .ZN(n3603) );
  AND2_X1 U4470 ( .A1(n6814), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5784) );
  INV_X1 U4471 ( .A(n5784), .ZN(n5005) );
  INV_X1 U4472 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3602) );
  OAI22_X1 U4473 ( .A1(n5646), .A2(n3603), .B1(n5005), .B2(n3602), .ZN(n3604)
         );
  AOI21_X1 U4474 ( .B1(n5785), .B2(EAX_REG_2__SCAN_IN), .A(n3604), .ZN(n3605)
         );
  AND2_X1 U4475 ( .A1(n3606), .A2(n3605), .ZN(n3638) );
  OR2_X1 U4476 ( .A1(n3637), .A2(n3638), .ZN(n3634) );
  AOI22_X1 U4477 ( .A1(n5681), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5629), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3612) );
  AOI22_X1 U4478 ( .A1(n4728), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5692), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4479 ( .A1(n5688), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3607), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3610) );
  INV_X1 U4480 ( .A(n3502), .ZN(n4709) );
  AOI22_X1 U4481 ( .A1(n3608), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3609) );
  NAND4_X1 U4482 ( .A1(n3612), .A2(n3611), .A3(n3610), .A4(n3609), .ZN(n3618)
         );
  AOI22_X1 U4483 ( .A1(n4995), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5683), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4484 ( .A1(n5691), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4485 ( .A1(n5682), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4486 ( .A1(n4729), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3613) );
  NAND4_X1 U4487 ( .A1(n3616), .A2(n3615), .A3(n3614), .A4(n3613), .ZN(n3617)
         );
  OR2_X1 U4488 ( .A1(n3618), .A2(n3617), .ZN(n3740) );
  NAND2_X1 U4489 ( .A1(n3648), .A2(n3740), .ZN(n3619) );
  AOI22_X1 U4490 ( .A1(n4146), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3621), 
        .B2(n3740), .ZN(n3622) );
  NAND2_X1 U4491 ( .A1(n3625), .A2(n3624), .ZN(n3630) );
  INV_X1 U4492 ( .A(n3626), .ZN(n3627) );
  NAND2_X1 U4493 ( .A1(n3628), .A2(n3627), .ZN(n3629) );
  NAND2_X1 U4494 ( .A1(n3630), .A2(n3629), .ZN(n3632) );
  OR2_X1 U4495 ( .A1(n3632), .A2(n3631), .ZN(n3633) );
  AND2_X2 U4496 ( .A1(n3692), .A2(n3633), .ZN(n5950) );
  AOI21_X1 U4497 ( .B1(n5950), .B2(n4754), .A(n5784), .ZN(n3639) );
  NAND2_X1 U4498 ( .A1(n3634), .A2(n3639), .ZN(n3636) );
  NAND2_X1 U4499 ( .A1(n3637), .A2(n3638), .ZN(n3635) );
  NAND2_X1 U4500 ( .A1(n3636), .A2(n3635), .ZN(n3830) );
  NAND3_X1 U4501 ( .A1(n3639), .A2(n3638), .A3(n3637), .ZN(n3640) );
  AND2_X1 U4502 ( .A1(n3830), .A2(n3640), .ZN(n6344) );
  INV_X1 U4503 ( .A(n6344), .ZN(n3987) );
  INV_X1 U4504 ( .A(DATAI_2_), .ZN(n3853) );
  INV_X1 U4505 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6279) );
  OAI222_X1 U4506 ( .A1(n3987), .A2(n5862), .B1(n5109), .B2(n3853), .C1(n5796), 
        .C2(n6279), .ZN(U2889) );
  NOR2_X1 U4507 ( .A1(n3641), .A2(n6587), .ZN(n3642) );
  NAND2_X1 U4508 ( .A1(n3643), .A2(n3642), .ZN(n3651) );
  INV_X1 U4509 ( .A(n3644), .ZN(n3647) );
  NAND4_X1 U4510 ( .A1(n3649), .A2(n3648), .A3(n3647), .A4(n5457), .ZN(n3650)
         );
  NAND2_X2 U4511 ( .A1(n3651), .A2(n3650), .ZN(n5848) );
  NAND2_X1 U4512 ( .A1(n5848), .A2(n5797), .ZN(n5852) );
  AND2_X1 U4513 ( .A1(n5848), .A2(n4787), .ZN(n5104) );
  INV_X2 U4514 ( .A(n5104), .ZN(n5850) );
  OAI222_X1 U4515 ( .A1(n5178), .A2(n5852), .B1(n5848), .B2(n7001), .C1(n6356), 
        .C2(n5850), .ZN(U2859) );
  INV_X1 U4516 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6937) );
  AOI22_X1 U4517 ( .A1(n6689), .A2(UWORD_REG_14__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n3652) );
  OAI21_X1 U4518 ( .B1(n6937), .B2(n6254), .A(n3652), .ZN(U2893) );
  INV_X1 U4519 ( .A(EAX_REG_16__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4520 ( .A1(n6689), .A2(UWORD_REG_0__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n3653) );
  OAI21_X1 U4521 ( .B1(n3654), .B2(n6254), .A(n3653), .ZN(U2907) );
  INV_X1 U4522 ( .A(EAX_REG_17__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4523 ( .A1(n6689), .A2(UWORD_REG_1__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n3655) );
  OAI21_X1 U4524 ( .B1(n3656), .B2(n6254), .A(n3655), .ZN(U2906) );
  INV_X1 U4525 ( .A(EAX_REG_18__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4526 ( .A1(n6689), .A2(UWORD_REG_2__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n3657) );
  OAI21_X1 U4527 ( .B1(n3658), .B2(n6254), .A(n3657), .ZN(U2905) );
  INV_X1 U4528 ( .A(EAX_REG_21__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4529 ( .A1(n6689), .A2(UWORD_REG_5__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n3659) );
  OAI21_X1 U4530 ( .B1(n3660), .B2(n6254), .A(n3659), .ZN(U2902) );
  INV_X1 U4531 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6289) );
  AOI22_X1 U4532 ( .A1(n6689), .A2(UWORD_REG_9__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n3661) );
  OAI21_X1 U4533 ( .B1(n6289), .B2(n6254), .A(n3661), .ZN(U2898) );
  INV_X1 U4534 ( .A(EAX_REG_27__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4535 ( .A1(n6689), .A2(UWORD_REG_11__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n3662) );
  OAI21_X1 U4536 ( .B1(n3663), .B2(n6254), .A(n3662), .ZN(U2896) );
  INV_X1 U4537 ( .A(EAX_REG_29__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4538 ( .A1(n6689), .A2(UWORD_REG_13__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n3664) );
  OAI21_X1 U4539 ( .B1(n3665), .B2(n6254), .A(n3664), .ZN(U2894) );
  INV_X1 U4540 ( .A(EAX_REG_20__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4541 ( .A1(n6689), .A2(UWORD_REG_4__SCAN_IN), .B1(
        DATAO_REG_20__SCAN_IN), .B2(n6283), .ZN(n3666) );
  OAI21_X1 U4542 ( .B1(n3667), .B2(n6254), .A(n3666), .ZN(U2903) );
  INV_X1 U4543 ( .A(EAX_REG_23__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4544 ( .A1(n6689), .A2(UWORD_REG_7__SCAN_IN), .B1(
        DATAO_REG_23__SCAN_IN), .B2(n6283), .ZN(n3668) );
  OAI21_X1 U4545 ( .B1(n3669), .B2(n6254), .A(n3668), .ZN(U2900) );
  INV_X1 U4546 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6810) );
  AOI22_X1 U4547 ( .A1(n6689), .A2(UWORD_REG_10__SCAN_IN), .B1(
        DATAO_REG_26__SCAN_IN), .B2(n6283), .ZN(n3670) );
  OAI21_X1 U4548 ( .B1(n6810), .B2(n6254), .A(n3670), .ZN(U2897) );
  INV_X1 U4549 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6296) );
  AOI22_X1 U4550 ( .A1(n6689), .A2(UWORD_REG_12__SCAN_IN), .B1(
        DATAO_REG_28__SCAN_IN), .B2(n6283), .ZN(n3671) );
  OAI21_X1 U4551 ( .B1(n6296), .B2(n6254), .A(n3671), .ZN(U2895) );
  INV_X1 U4552 ( .A(n3672), .ZN(n3674) );
  OR2_X1 U4553 ( .A1(n3363), .A2(n3214), .ZN(n3679) );
  NAND3_X1 U4554 ( .A1(n6674), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6447) );
  INV_X1 U4555 ( .A(n6447), .ZN(n6446) );
  NAND2_X1 U4556 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6446), .ZN(n6439) );
  NAND2_X1 U4557 ( .A1(n6674), .A2(n6439), .ZN(n3675) );
  NAND3_X1 U4558 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4260) );
  INV_X1 U4559 ( .A(n4260), .ZN(n3891) );
  NAND2_X1 U4560 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3891), .ZN(n3937) );
  AND2_X1 U4561 ( .A1(n3675), .A2(n3937), .ZN(n4308) );
  AOI22_X1 U4562 ( .A1(n3677), .A2(n4308), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3676), .ZN(n3678) );
  AOI22_X1 U4563 ( .A1(n5681), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n5629), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4564 ( .A1(n5680), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5692), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4565 ( .A1(n5688), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3607), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4566 ( .A1(n3608), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3680) );
  NAND4_X1 U4567 ( .A1(n3683), .A2(n3682), .A3(n3681), .A4(n3680), .ZN(n3689)
         );
  AOI22_X1 U4568 ( .A1(n4995), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5634), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4569 ( .A1(n5691), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4570 ( .A1(n5682), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4571 ( .A1(n4729), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3684) );
  NAND4_X1 U4572 ( .A1(n3687), .A2(n3686), .A3(n3685), .A4(n3684), .ZN(n3688)
         );
  OR2_X1 U4573 ( .A1(n3689), .A2(n3688), .ZN(n3741) );
  AOI22_X1 U4574 ( .A1(n4146), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4443), 
        .B2(n3741), .ZN(n3690) );
  NAND2_X1 U4575 ( .A1(n3692), .A2(n3943), .ZN(n3693) );
  AND2_X2 U4576 ( .A1(n3819), .A2(n3693), .ZN(n6667) );
  INV_X1 U4577 ( .A(n3694), .ZN(n3824) );
  INV_X1 U4578 ( .A(n5703), .ZN(n5706) );
  INV_X1 U4579 ( .A(n3695), .ZN(n3697) );
  NOR2_X2 U4580 ( .A1(n3695), .A2(n5471), .ZN(n3821) );
  INV_X1 U4581 ( .A(n3821), .ZN(n3696) );
  OAI21_X1 U4582 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3697), .A(n3696), 
        .ZN(n5470) );
  AOI22_X1 U4583 ( .A1(n5706), .A2(n5470), .B1(n5784), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3699) );
  NAND2_X1 U4584 ( .A1(n5785), .A2(EAX_REG_3__SCAN_IN), .ZN(n3698) );
  OAI211_X1 U4585 ( .C1(n3824), .C2(n3214), .A(n3699), .B(n3698), .ZN(n3700)
         );
  AOI21_X1 U4586 ( .B1(n6667), .B2(n4754), .A(n3700), .ZN(n3829) );
  NOR2_X1 U4587 ( .A1(n3830), .A2(n3829), .ZN(n4008) );
  AOI21_X1 U4588 ( .B1(n3829), .B2(n3830), .A(n4008), .ZN(n5482) );
  INV_X1 U4589 ( .A(n5482), .ZN(n3992) );
  INV_X1 U4590 ( .A(DATAI_3_), .ZN(n3800) );
  INV_X1 U4591 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6276) );
  OAI222_X1 U4592 ( .A1(n3992), .A2(n5862), .B1(n5109), .B2(n3800), .C1(n5796), 
        .C2(n6276), .ZN(U2888) );
  NOR2_X1 U4593 ( .A1(n5806), .A2(FLUSH_REG_SCAN_IN), .ZN(n3726) );
  INV_X1 U4594 ( .A(n3726), .ZN(n3722) );
  INV_X1 U4595 ( .A(n3705), .ZN(n3721) );
  MUX2_X1 U4596 ( .A(n3701), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(n3727), 
        .Z(n6559) );
  NAND2_X1 U4597 ( .A1(n5469), .A2(n3703), .ZN(n3719) );
  MUX2_X1 U4598 ( .A(n3704), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n3399), 
        .Z(n3706) );
  NOR2_X1 U4599 ( .A1(n3706), .A2(n3705), .ZN(n3716) );
  INV_X1 U4600 ( .A(n3707), .ZN(n3708) );
  OAI21_X1 U4601 ( .B1(n3399), .B2(n3214), .A(n3708), .ZN(n3709) );
  NOR2_X1 U4602 ( .A1(n3709), .A2(n5692), .ZN(n5955) );
  NAND2_X1 U4603 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3710) );
  INV_X1 U4604 ( .A(n3710), .ZN(n3711) );
  MUX2_X1 U4605 ( .A(n3711), .B(n3710), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n3712) );
  NAND2_X1 U4606 ( .A1(n5803), .A2(n3712), .ZN(n3713) );
  OAI21_X1 U4607 ( .B1(n5955), .B2(n3714), .A(n3713), .ZN(n3715) );
  AOI21_X1 U4608 ( .B1(n3717), .B2(n3716), .A(n3715), .ZN(n3718) );
  NAND2_X1 U4609 ( .A1(n3719), .A2(n3718), .ZN(n5954) );
  INV_X1 U4610 ( .A(n3727), .ZN(n6555) );
  MUX2_X1 U4611 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5954), .S(n6555), 
        .Z(n6561) );
  NAND3_X1 U4612 ( .A1(n6559), .A2(n6561), .A3(n5806), .ZN(n3720) );
  OAI21_X1 U4613 ( .B1(n3722), .B2(n3721), .A(n3720), .ZN(n6571) );
  INV_X1 U4614 ( .A(n6571), .ZN(n3732) );
  INV_X1 U4615 ( .A(n5114), .ZN(n4231) );
  OR2_X1 U4616 ( .A1(n3723), .A2(n4231), .ZN(n3724) );
  XNOR2_X1 U4617 ( .A(n3724), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6226)
         );
  NAND3_X1 U4618 ( .A1(n6226), .A2(n6080), .A3(n5806), .ZN(n3730) );
  AOI21_X1 U4619 ( .B1(n3727), .B2(n5806), .A(n3726), .ZN(n3728) );
  OR2_X1 U4620 ( .A1(n3728), .A2(n6083), .ZN(n3729) );
  NAND2_X1 U4621 ( .A1(n3730), .A2(n3729), .ZN(n6570) );
  INV_X1 U4622 ( .A(n6570), .ZN(n3731) );
  OAI21_X1 U4623 ( .B1(n3732), .B2(n5800), .A(n3731), .ZN(n3736) );
  NOR2_X1 U4624 ( .A1(n3736), .A2(FLUSH_REG_SCAN_IN), .ZN(n3734) );
  INV_X1 U4625 ( .A(n3733), .ZN(n6664) );
  NOR2_X1 U4626 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6692) );
  INV_X1 U4627 ( .A(n6692), .ZN(n6582) );
  OAI21_X1 U4628 ( .B1(n3734), .B2(n6664), .A(n4310), .ZN(n6675) );
  NOR2_X1 U4629 ( .A1(n3736), .A2(n3735), .ZN(n6579) );
  INV_X1 U4630 ( .A(n5118), .ZN(n6492) );
  INV_X1 U4631 ( .A(n3110), .ZN(n5179) );
  AND2_X1 U4632 ( .A1(n6826), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6670) );
  OAI22_X1 U4633 ( .A1(n5111), .A2(n6492), .B1(n5179), .B2(n6670), .ZN(n3737)
         );
  OAI21_X1 U4634 ( .B1(n6579), .B2(n3737), .A(n6675), .ZN(n3738) );
  OAI21_X1 U4635 ( .B1(n6675), .B2(n6927), .A(n3738), .ZN(U3465) );
  INV_X2 U4636 ( .A(n6667), .ZN(n3953) );
  NAND2_X1 U4637 ( .A1(n3744), .A2(n3745), .ZN(n3757) );
  INV_X1 U4638 ( .A(n3740), .ZN(n3758) );
  NAND2_X1 U4639 ( .A1(n3757), .A2(n3758), .ZN(n3756) );
  NAND2_X1 U4640 ( .A1(n3756), .A2(n3741), .ZN(n4127) );
  OAI211_X1 U4641 ( .C1(n3741), .C2(n3756), .A(n4127), .B(n5182), .ZN(n3742)
         );
  NAND2_X1 U4642 ( .A1(n5946), .A2(n4448), .ZN(n3752) );
  OAI21_X1 U4643 ( .B1(n3745), .B2(n3744), .A(n3757), .ZN(n3749) );
  INV_X1 U4644 ( .A(n3746), .ZN(n3748) );
  OAI211_X1 U4645 ( .C1(n3749), .C2(n6691), .A(n3748), .B(n3747), .ZN(n3750)
         );
  INV_X1 U4646 ( .A(n3750), .ZN(n3751) );
  NAND2_X1 U4647 ( .A1(n3752), .A2(n3751), .ZN(n6350) );
  XNOR2_X1 U4648 ( .A(n3753), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6349)
         );
  NAND2_X1 U4649 ( .A1(n6350), .A2(n6349), .ZN(n6348) );
  INV_X1 U4650 ( .A(n3753), .ZN(n3754) );
  NAND2_X1 U4651 ( .A1(n3754), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3755)
         );
  NAND2_X1 U4652 ( .A1(n6348), .A2(n3755), .ZN(n6342) );
  INV_X1 U4653 ( .A(n5950), .ZN(n3942) );
  OAI21_X1 U4654 ( .B1(n3758), .B2(n3757), .A(n3756), .ZN(n3761) );
  INV_X1 U4655 ( .A(n3759), .ZN(n3760) );
  AOI21_X1 U4656 ( .B1(n3761), .B2(n5182), .A(n3760), .ZN(n3762) );
  OAI21_X1 U4657 ( .B1(n3942), .B2(n4460), .A(n3762), .ZN(n6341) );
  OAI21_X1 U4658 ( .B1(n6342), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .A(n6341), 
        .ZN(n3764) );
  NAND2_X1 U4659 ( .A1(n6342), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3763)
         );
  NAND2_X1 U4660 ( .A1(n3764), .A2(n3763), .ZN(n3998) );
  XNOR2_X1 U4661 ( .A(n3999), .B(n3998), .ZN(n6407) );
  NAND3_X1 U4662 ( .A1(n6580), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6593) );
  INV_X1 U4663 ( .A(n6593), .ZN(n3765) );
  NAND2_X1 U4664 ( .A1(n3765), .A2(n6445), .ZN(n5901) );
  NAND2_X1 U4665 ( .A1(n6492), .A2(n3766), .ZN(n6687) );
  NAND2_X1 U4666 ( .A1(n6687), .A2(n6580), .ZN(n3767) );
  NAND2_X1 U4667 ( .A1(n6580), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3769) );
  NAND2_X1 U4668 ( .A1(n6091), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3768) );
  NAND2_X1 U4669 ( .A1(n3769), .A2(n3768), .ZN(n6362) );
  INV_X1 U4670 ( .A(n6426), .ZN(n6379) );
  AOI22_X1 U4671 ( .A1(n6363), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n6379), 
        .B2(REIP_REG_3__SCAN_IN), .ZN(n3770) );
  OAI21_X1 U4672 ( .B1(n5470), .B2(n6355), .A(n3770), .ZN(n3771) );
  AOI21_X1 U4673 ( .B1(n5482), .B2(n6360), .A(n3771), .ZN(n3772) );
  OAI21_X1 U4674 ( .B1(n6323), .B2(n6407), .A(n3772), .ZN(U2983) );
  NAND3_X1 U4675 ( .A1(n6674), .A2(n6560), .A3(n4181), .ZN(n4015) );
  OR2_X1 U4676 ( .A1(n6927), .A2(n4015), .ZN(n4119) );
  NOR2_X1 U4677 ( .A1(n3925), .A2(n5797), .ZN(n6544) );
  INV_X1 U4678 ( .A(n6544), .ZN(n5143) );
  INV_X1 U4679 ( .A(n5948), .ZN(n6233) );
  OR2_X1 U4680 ( .A1(n4068), .A2(n6233), .ZN(n4304) );
  NOR2_X1 U4681 ( .A1(n5469), .A2(n4304), .ZN(n4022) );
  NAND2_X1 U4682 ( .A1(n4022), .A2(n3110), .ZN(n3774) );
  NAND2_X1 U4683 ( .A1(n3774), .A2(n4119), .ZN(n3777) );
  NOR2_X1 U4684 ( .A1(n5950), .A2(n5946), .ZN(n3775) );
  NAND2_X1 U4685 ( .A1(n3953), .A2(n3775), .ZN(n3781) );
  OAI21_X1 U4686 ( .B1(n3781), .B2(n6091), .A(n5118), .ZN(n3779) );
  AOI21_X1 U4687 ( .B1(n6927), .B2(STATE2_REG_3__SCAN_IN), .A(n4310), .ZN(
        n6494) );
  NAND2_X1 U4688 ( .A1(n6492), .A2(n4015), .ZN(n3776) );
  OAI211_X1 U4689 ( .C1(n3777), .C2(n3779), .A(n6494), .B(n3776), .ZN(n4113)
         );
  NAND2_X1 U4690 ( .A1(n4113), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3784) );
  INV_X1 U4691 ( .A(n3777), .ZN(n3778) );
  OAI22_X1 U4692 ( .A1(n3779), .A2(n3778), .B1(n4015), .B2(n6814), .ZN(n4116)
         );
  NOR2_X1 U4693 ( .A1(n3780), .A2(n4310), .ZN(n6546) );
  NAND2_X1 U4694 ( .A1(n6360), .A2(DATAI_31_), .ZN(n6485) );
  NAND2_X1 U4695 ( .A1(n6360), .A2(DATAI_23_), .ZN(n6551) );
  OAI22_X1 U4696 ( .A1(n6485), .A2(n4114), .B1(n4525), .B2(n6551), .ZN(n3782)
         );
  AOI21_X1 U4697 ( .B1(n4116), .B2(n6546), .A(n3782), .ZN(n3783) );
  OAI211_X1 U4698 ( .C1(n4119), .C2(n5143), .A(n3784), .B(n3783), .ZN(U3035)
         );
  NOR2_X1 U4699 ( .A1(n3925), .A2(n3785), .ZN(n6488) );
  INV_X1 U4700 ( .A(n6488), .ZN(n5135) );
  NAND2_X1 U4701 ( .A1(n4113), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3789) );
  NOR2_X1 U4702 ( .A1(n3786), .A2(n4310), .ZN(n6499) );
  NAND2_X1 U4703 ( .A1(n6360), .A2(DATAI_24_), .ZN(n6502) );
  NAND2_X1 U4704 ( .A1(n6360), .A2(DATAI_16_), .ZN(n6452) );
  OAI22_X1 U4705 ( .A1(n6502), .A2(n4114), .B1(n4525), .B2(n6452), .ZN(n3787)
         );
  AOI21_X1 U4706 ( .B1(n4116), .B2(n6499), .A(n3787), .ZN(n3788) );
  OAI211_X1 U4707 ( .C1(n5135), .C2(n4119), .A(n3789), .B(n3788), .ZN(U3028)
         );
  NOR2_X1 U4708 ( .A1(n3925), .A2(n3790), .ZN(n6504) );
  INV_X1 U4709 ( .A(n6504), .ZN(n5158) );
  NAND2_X1 U4710 ( .A1(n4113), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3794) );
  NOR2_X1 U4711 ( .A1(n3791), .A2(n4310), .ZN(n6505) );
  NAND2_X1 U4712 ( .A1(n6360), .A2(DATAI_25_), .ZN(n6508) );
  NAND2_X1 U4713 ( .A1(n6360), .A2(DATAI_17_), .ZN(n6456) );
  OAI22_X1 U4714 ( .A1(n6508), .A2(n4114), .B1(n4525), .B2(n6456), .ZN(n3792)
         );
  AOI21_X1 U4715 ( .B1(n4116), .B2(n6505), .A(n3792), .ZN(n3793) );
  OAI211_X1 U4716 ( .C1(n4119), .C2(n5158), .A(n3794), .B(n3793), .ZN(U3029)
         );
  NOR2_X1 U4717 ( .A1(n3925), .A2(n3795), .ZN(n6522) );
  INV_X1 U4718 ( .A(n6522), .ZN(n5127) );
  NAND2_X1 U4719 ( .A1(n4113), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3798) );
  INV_X1 U4720 ( .A(DATAI_4_), .ZN(n4098) );
  NOR2_X1 U4721 ( .A1(n4098), .A2(n4310), .ZN(n6523) );
  NAND2_X1 U4722 ( .A1(n6360), .A2(DATAI_28_), .ZN(n6466) );
  NAND2_X1 U4723 ( .A1(n6360), .A2(DATAI_20_), .ZN(n6526) );
  OAI22_X1 U4724 ( .A1(n6466), .A2(n4114), .B1(n4525), .B2(n6526), .ZN(n3796)
         );
  AOI21_X1 U4725 ( .B1(n4116), .B2(n6523), .A(n3796), .ZN(n3797) );
  OAI211_X1 U4726 ( .C1(n4119), .C2(n5127), .A(n3798), .B(n3797), .ZN(U3032)
         );
  NOR2_X1 U4727 ( .A1(n3925), .A2(n3799), .ZN(n6516) );
  INV_X1 U4728 ( .A(n6516), .ZN(n5139) );
  NAND2_X1 U4729 ( .A1(n4113), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3803) );
  NOR2_X1 U4730 ( .A1(n3800), .A2(n4310), .ZN(n6517) );
  NAND2_X1 U4731 ( .A1(n6360), .A2(DATAI_27_), .ZN(n6462) );
  NAND2_X1 U4732 ( .A1(n6360), .A2(DATAI_19_), .ZN(n6520) );
  OAI22_X1 U4733 ( .A1(n6462), .A2(n4114), .B1(n4525), .B2(n6520), .ZN(n3801)
         );
  AOI21_X1 U4734 ( .B1(n4116), .B2(n6517), .A(n3801), .ZN(n3802) );
  OAI211_X1 U4735 ( .C1(n4119), .C2(n5139), .A(n3803), .B(n3802), .ZN(U3031)
         );
  INV_X1 U4736 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U4737 ( .A1(n4995), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4738 ( .A1(n5688), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4729), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4739 ( .A1(n5691), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4740 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n3607), .B1(n4709), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3804) );
  NAND4_X1 U4741 ( .A1(n3807), .A2(n3806), .A3(n3805), .A4(n3804), .ZN(n3814)
         );
  AOI22_X1 U4742 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3608), .B1(n5680), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4743 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n5620), .B1(n5692), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4744 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n5634), .B1(n5682), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3810) );
  INV_X1 U4745 ( .A(n3808), .ZN(n5629) );
  AOI22_X1 U4746 ( .A1(n5629), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3809) );
  NAND4_X1 U4747 ( .A1(n3812), .A2(n3811), .A3(n3810), .A4(n3809), .ZN(n3813)
         );
  OR2_X1 U4748 ( .A1(n3814), .A2(n3813), .ZN(n4125) );
  NAND2_X1 U4749 ( .A1(n4443), .A2(n4125), .ZN(n3815) );
  OAI21_X1 U4750 ( .B1(n4446), .B2(n4044), .A(n3815), .ZN(n3817) );
  INV_X1 U4751 ( .A(n3817), .ZN(n3818) );
  NAND2_X1 U4752 ( .A1(n3819), .A2(n3818), .ZN(n3820) );
  NAND2_X1 U4753 ( .A1(n3843), .A2(n3820), .ZN(n4003) );
  INV_X1 U4754 ( .A(n4754), .ZN(n4507) );
  NOR2_X1 U4755 ( .A1(n4003), .A2(n4507), .ZN(n3828) );
  OAI21_X1 U4756 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3821), .A(n3845), 
        .ZN(n6221) );
  OAI21_X1 U4757 ( .B1(n6091), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6814), 
        .ZN(n3823) );
  NAND2_X1 U4758 ( .A1(n5785), .A2(EAX_REG_4__SCAN_IN), .ZN(n3822) );
  OAI211_X1 U4759 ( .C1(n3824), .C2(n6083), .A(n3823), .B(n3822), .ZN(n3825)
         );
  OAI21_X1 U4760 ( .B1(n5646), .B2(n6221), .A(n3825), .ZN(n3826) );
  INV_X1 U4761 ( .A(n3826), .ZN(n3827) );
  NOR2_X1 U4762 ( .A1(n3828), .A2(n3827), .ZN(n4011) );
  OR2_X2 U4763 ( .A1(n4011), .A2(n3829), .ZN(n3831) );
  AOI22_X1 U4764 ( .A1(n5681), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n5629), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4765 ( .A1(n5680), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5692), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4766 ( .A1(n5688), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3607), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4767 ( .A1(n3608), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3832) );
  NAND4_X1 U4768 ( .A1(n3835), .A2(n3834), .A3(n3833), .A4(n3832), .ZN(n3841)
         );
  AOI22_X1 U4769 ( .A1(n4995), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n5683), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4770 ( .A1(n5691), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4771 ( .A1(n5682), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4772 ( .A1(n4729), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3836) );
  NAND4_X1 U4773 ( .A1(n3839), .A2(n3838), .A3(n3837), .A4(n3836), .ZN(n3840)
         );
  OR2_X1 U4774 ( .A1(n3841), .A2(n3840), .ZN(n4128) );
  AOI22_X1 U4775 ( .A1(n4146), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4443), 
        .B2(n4128), .ZN(n3842) );
  NAND2_X1 U4776 ( .A1(n3843), .A2(n3842), .ZN(n3844) );
  NAND2_X1 U4777 ( .A1(n4150), .A2(n3844), .ZN(n4131) );
  OAI21_X1 U4778 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3846), .A(n4210), 
        .ZN(n6331) );
  AOI22_X1 U4779 ( .A1(n5706), .A2(n6331), .B1(n5784), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3848) );
  NAND2_X1 U4780 ( .A1(n5785), .A2(EAX_REG_5__SCAN_IN), .ZN(n3847) );
  OAI211_X1 U4781 ( .C1(n4131), .C2(n4507), .A(n3848), .B(n3847), .ZN(n3849)
         );
  NAND2_X1 U4782 ( .A1(n4009), .A2(n3849), .ZN(n4217) );
  OR2_X1 U4783 ( .A1(n4009), .A2(n3849), .ZN(n3850) );
  AND2_X1 U4784 ( .A1(n4217), .A2(n3850), .ZN(n6334) );
  INV_X1 U4785 ( .A(n6334), .ZN(n3884) );
  INV_X1 U4786 ( .A(n5109), .ZN(n5039) );
  AOI22_X1 U4787 ( .A1(n5039), .A2(DATAI_5_), .B1(EAX_REG_5__SCAN_IN), .B2(
        n6250), .ZN(n3851) );
  OAI21_X1 U4788 ( .B1(n3884), .B2(n5862), .A(n3851), .ZN(U2886) );
  NOR2_X1 U4789 ( .A1(n3925), .A2(n3852), .ZN(n6510) );
  INV_X1 U4790 ( .A(n6510), .ZN(n5131) );
  NAND2_X1 U4791 ( .A1(n4113), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3856) );
  NOR2_X1 U4792 ( .A1(n3853), .A2(n4310), .ZN(n6511) );
  AND2_X1 U4793 ( .A1(n6360), .A2(DATAI_26_), .ZN(n6509) );
  INV_X1 U4794 ( .A(n6509), .ZN(n5311) );
  NAND2_X1 U4795 ( .A1(n6360), .A2(DATAI_18_), .ZN(n6514) );
  OAI22_X1 U4796 ( .A1(n5311), .A2(n4114), .B1(n4525), .B2(n6514), .ZN(n3854)
         );
  AOI21_X1 U4797 ( .B1(n4116), .B2(n6511), .A(n3854), .ZN(n3855) );
  OAI211_X1 U4798 ( .C1(n4119), .C2(n5131), .A(n3856), .B(n3855), .ZN(U3030)
         );
  INV_X1 U4799 ( .A(EBX_REG_5__SCAN_IN), .ZN(n3883) );
  INV_X1 U4800 ( .A(n5457), .ZN(n3857) );
  INV_X1 U4801 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3859) );
  NAND2_X1 U4802 ( .A1(n3866), .A2(n3859), .ZN(n3863) );
  INV_X1 U4803 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3858) );
  NAND2_X1 U4804 ( .A1(n5658), .A2(n3858), .ZN(n3861) );
  NAND2_X1 U4805 ( .A1(n5457), .A2(n3859), .ZN(n3860) );
  NAND3_X1 U4806 ( .A1(n3861), .A2(n5659), .A3(n3860), .ZN(n3862) );
  NAND2_X1 U4807 ( .A1(n3863), .A2(n3862), .ZN(n3865) );
  XNOR2_X1 U4808 ( .A(n3865), .B(n3864), .ZN(n3993) );
  NAND2_X1 U4809 ( .A1(n3993), .A2(n5457), .ZN(n3995) );
  INV_X1 U4810 ( .A(EBX_REG_2__SCAN_IN), .ZN(n7007) );
  NAND2_X1 U4811 ( .A1(n5456), .A2(n7007), .ZN(n3871) );
  INV_X1 U4812 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3867) );
  NAND2_X1 U4813 ( .A1(n3112), .A2(n3867), .ZN(n3869) );
  NAND2_X1 U4814 ( .A1(n5457), .A2(n7007), .ZN(n3868) );
  NAND3_X1 U4815 ( .A1(n3869), .A2(n5659), .A3(n3868), .ZN(n3870) );
  NAND2_X1 U4816 ( .A1(n5457), .A2(n5659), .ZN(n5569) );
  MUX2_X1 U4817 ( .A(n5569), .B(n5659), .S(EBX_REG_3__SCAN_IN), .Z(n3874) );
  OAI21_X1 U4818 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n5774), .A(n3874), 
        .ZN(n3988) );
  OR2_X2 U4819 ( .A1(n3989), .A2(n3988), .ZN(n4063) );
  INV_X1 U4820 ( .A(n4063), .ZN(n3879) );
  MUX2_X1 U4821 ( .A(n5662), .B(n3112), .S(EBX_REG_4__SCAN_IN), .Z(n3877) );
  INV_X1 U4822 ( .A(n3112), .ZN(n4856) );
  NAND2_X1 U4823 ( .A1(n4856), .A2(n5773), .ZN(n5059) );
  NAND2_X1 U4824 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n5773), .ZN(n3875)
         );
  AND2_X1 U4825 ( .A1(n5059), .A2(n3875), .ZN(n3876) );
  NAND2_X1 U4826 ( .A1(n3877), .A2(n3876), .ZN(n4062) );
  MUX2_X1 U4827 ( .A(n5569), .B(n4155), .S(EBX_REG_5__SCAN_IN), .Z(n3878) );
  AND2_X1 U4828 ( .A1(n3878), .A2(n3117), .ZN(n3880) );
  AOI21_X1 U4829 ( .B1(n3879), .B2(n4062), .A(n3880), .ZN(n3882) );
  NAND2_X1 U4830 ( .A1(n3880), .A2(n4062), .ZN(n3881) );
  OR2_X1 U4831 ( .A1(n3882), .A2(n4162), .ZN(n6205) );
  OAI222_X1 U4832 ( .A1(n3884), .A2(n5850), .B1(n5848), .B2(n3883), .C1(n5852), 
        .C2(n6205), .ZN(U2854) );
  NAND2_X1 U4833 ( .A1(n5469), .A2(n3110), .ZN(n4182) );
  NAND2_X1 U4834 ( .A1(n4068), .A2(n6233), .ZN(n5115) );
  OR2_X1 U4835 ( .A1(n4182), .A2(n5115), .ZN(n3885) );
  AND2_X1 U4836 ( .A1(n3885), .A2(n3937), .ZN(n3890) );
  INV_X1 U4837 ( .A(n3943), .ZN(n3886) );
  NAND2_X1 U4838 ( .A1(n5950), .A2(n3886), .ZN(n3941) );
  NOR2_X1 U4839 ( .A1(n3941), .A2(n4230), .ZN(n3889) );
  AND2_X1 U4840 ( .A1(n5118), .A2(n6091), .ZN(n6666) );
  INV_X1 U4841 ( .A(n6666), .ZN(n4526) );
  OAI21_X1 U4842 ( .B1(n3889), .B2(n5901), .A(n4526), .ZN(n3887) );
  AOI22_X1 U4843 ( .A1(n3890), .A2(n3887), .B1(n4260), .B2(n6492), .ZN(n3888)
         );
  NAND2_X1 U4844 ( .A1(n6494), .A2(n3888), .ZN(n3939) );
  INV_X1 U4845 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3898) );
  INV_X1 U4846 ( .A(n3937), .ZN(n3930) );
  NAND2_X1 U4847 ( .A1(n3889), .A2(n5111), .ZN(n4292) );
  INV_X1 U4848 ( .A(n6526), .ZN(n6463) );
  NAND2_X1 U4849 ( .A1(n4054), .A2(n6463), .ZN(n3895) );
  OR2_X1 U4850 ( .A1(n3890), .A2(n6492), .ZN(n3893) );
  NAND2_X1 U4851 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n3891), .ZN(n3892) );
  NAND2_X1 U4852 ( .A1(n3893), .A2(n3892), .ZN(n3934) );
  NAND2_X1 U4853 ( .A1(n3934), .A2(n6523), .ZN(n3894) );
  OAI211_X1 U4854 ( .C1(n4292), .C2(n6466), .A(n3895), .B(n3894), .ZN(n3896)
         );
  AOI21_X1 U4855 ( .B1(n3930), .B2(n6522), .A(n3896), .ZN(n3897) );
  OAI21_X1 U4856 ( .B1(n3933), .B2(n3898), .A(n3897), .ZN(U3144) );
  INV_X1 U4857 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3903) );
  INV_X1 U4858 ( .A(n6514), .ZN(n5309) );
  NAND2_X1 U4859 ( .A1(n4054), .A2(n5309), .ZN(n3900) );
  NAND2_X1 U4860 ( .A1(n3934), .A2(n6511), .ZN(n3899) );
  OAI211_X1 U4861 ( .C1(n4292), .C2(n5311), .A(n3900), .B(n3899), .ZN(n3901)
         );
  AOI21_X1 U4862 ( .B1(n3930), .B2(n6510), .A(n3901), .ZN(n3902) );
  OAI21_X1 U4863 ( .B1(n3933), .B2(n3903), .A(n3902), .ZN(U3142) );
  INV_X1 U4864 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3908) );
  INV_X1 U4865 ( .A(n6551), .ZN(n6478) );
  NAND2_X1 U4866 ( .A1(n4054), .A2(n6478), .ZN(n3905) );
  NAND2_X1 U4867 ( .A1(n3934), .A2(n6546), .ZN(n3904) );
  OAI211_X1 U4868 ( .C1(n4292), .C2(n6485), .A(n3905), .B(n3904), .ZN(n3906)
         );
  AOI21_X1 U4869 ( .B1(n3930), .B2(n6544), .A(n3906), .ZN(n3907) );
  OAI21_X1 U4870 ( .B1(n3933), .B2(n3908), .A(n3907), .ZN(U3147) );
  INV_X1 U4871 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3913) );
  INV_X1 U4872 ( .A(n6456), .ZN(n6503) );
  NAND2_X1 U4873 ( .A1(n4054), .A2(n6503), .ZN(n3910) );
  NAND2_X1 U4874 ( .A1(n3934), .A2(n6505), .ZN(n3909) );
  OAI211_X1 U4875 ( .C1(n4292), .C2(n6508), .A(n3910), .B(n3909), .ZN(n3911)
         );
  AOI21_X1 U4876 ( .B1(n3930), .B2(n6504), .A(n3911), .ZN(n3912) );
  OAI21_X1 U4877 ( .B1(n3933), .B2(n3913), .A(n3912), .ZN(U3141) );
  INV_X1 U4878 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3918) );
  INV_X1 U4879 ( .A(n6520), .ZN(n6459) );
  NAND2_X1 U4880 ( .A1(n4054), .A2(n6459), .ZN(n3915) );
  NAND2_X1 U4881 ( .A1(n3934), .A2(n6517), .ZN(n3914) );
  OAI211_X1 U4882 ( .C1(n4292), .C2(n6462), .A(n3915), .B(n3914), .ZN(n3916)
         );
  AOI21_X1 U4883 ( .B1(n3930), .B2(n6516), .A(n3916), .ZN(n3917) );
  OAI21_X1 U4884 ( .B1(n3933), .B2(n3918), .A(n3917), .ZN(U3143) );
  INV_X1 U4885 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3924) );
  NOR2_X1 U4886 ( .A1(n3925), .A2(n3919), .ZN(n6535) );
  NAND2_X1 U4887 ( .A1(n6360), .A2(DATAI_30_), .ZN(n6540) );
  NAND2_X1 U4888 ( .A1(n6360), .A2(DATAI_22_), .ZN(n6476) );
  INV_X1 U4889 ( .A(n6476), .ZN(n6533) );
  NAND2_X1 U4890 ( .A1(n4054), .A2(n6533), .ZN(n3921) );
  NOR2_X1 U4891 ( .A1(n4227), .A2(n4310), .ZN(n6536) );
  NAND2_X1 U4892 ( .A1(n3934), .A2(n6536), .ZN(n3920) );
  OAI211_X1 U4893 ( .C1(n4292), .C2(n6540), .A(n3921), .B(n3920), .ZN(n3922)
         );
  AOI21_X1 U4894 ( .B1(n3930), .B2(n6535), .A(n3922), .ZN(n3923) );
  OAI21_X1 U4895 ( .B1(n3933), .B2(n3924), .A(n3923), .ZN(U3146) );
  INV_X1 U4896 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3932) );
  NOR2_X1 U4897 ( .A1(n3925), .A2(n4788), .ZN(n6528) );
  NAND2_X1 U4898 ( .A1(n6360), .A2(DATAI_29_), .ZN(n6470) );
  NAND2_X1 U4899 ( .A1(n6360), .A2(DATAI_21_), .ZN(n6532) );
  INV_X1 U4900 ( .A(n6532), .ZN(n6467) );
  NAND2_X1 U4901 ( .A1(n4054), .A2(n6467), .ZN(n3928) );
  NOR2_X1 U4902 ( .A1(n3926), .A2(n4310), .ZN(n6529) );
  NAND2_X1 U4903 ( .A1(n3934), .A2(n6529), .ZN(n3927) );
  OAI211_X1 U4904 ( .C1(n4292), .C2(n6470), .A(n3928), .B(n3927), .ZN(n3929)
         );
  AOI21_X1 U4905 ( .B1(n3930), .B2(n6528), .A(n3929), .ZN(n3931) );
  OAI21_X1 U4906 ( .B1(n3933), .B2(n3932), .A(n3931), .ZN(U3145) );
  INV_X1 U4907 ( .A(n6452), .ZN(n6487) );
  AOI22_X1 U4908 ( .A1(n4054), .A2(n6487), .B1(n6499), .B2(n3934), .ZN(n3936)
         );
  OR2_X1 U4909 ( .A1(n4292), .A2(n6502), .ZN(n3935) );
  OAI211_X1 U4910 ( .C1(n5135), .C2(n3937), .A(n3936), .B(n3935), .ZN(n3938)
         );
  AOI21_X1 U4911 ( .B1(n3939), .B2(INSTQUEUE_REG_15__0__SCAN_IN), .A(n3938), 
        .ZN(n3940) );
  INV_X1 U4912 ( .A(n3940), .ZN(U3140) );
  NOR2_X1 U4913 ( .A1(n3941), .A2(n5946), .ZN(n4066) );
  INV_X1 U4914 ( .A(n4066), .ZN(n4067) );
  INV_X1 U4915 ( .A(n6490), .ZN(n3944) );
  AND2_X1 U4916 ( .A1(n5946), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6489) );
  NAND2_X1 U4917 ( .A1(n5112), .A2(n6489), .ZN(n6441) );
  NAND3_X1 U4918 ( .A1(n4067), .A2(n3944), .A3(n6441), .ZN(n3945) );
  NAND2_X1 U4919 ( .A1(n3945), .A2(n6445), .ZN(n6669) );
  INV_X1 U4920 ( .A(n6489), .ZN(n5945) );
  OAI21_X1 U4921 ( .B1(n5950), .B2(n5945), .A(n6445), .ZN(n3946) );
  NAND2_X1 U4922 ( .A1(n6669), .A2(n3946), .ZN(n3950) );
  OR2_X1 U4923 ( .A1(n4068), .A2(n5948), .ZN(n5278) );
  NOR2_X1 U4924 ( .A1(n5469), .A2(n5278), .ZN(n4535) );
  NOR2_X1 U4925 ( .A1(n6486), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3978)
         );
  AOI21_X1 U4926 ( .B1(n4535), .B2(n3110), .A(n3978), .ZN(n3949) );
  INV_X1 U4927 ( .A(n3949), .ZN(n3948) );
  NAND3_X1 U4928 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6674), .A3(n6560), .ZN(n4524) );
  INV_X1 U4929 ( .A(n4524), .ZN(n3947) );
  AOI22_X1 U4930 ( .A1(n3950), .A2(n3948), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3947), .ZN(n3981) );
  INV_X1 U4931 ( .A(n6499), .ZN(n5292) );
  AOI22_X1 U4932 ( .A1(n3950), .A2(n3949), .B1(n4524), .B2(n6492), .ZN(n3951)
         );
  NAND2_X1 U4933 ( .A1(n6494), .A2(n3951), .ZN(n3976) );
  NAND2_X1 U4934 ( .A1(n3976), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3957) );
  NOR2_X1 U4935 ( .A1(n6667), .A2(n5950), .ZN(n3952) );
  NOR3_X1 U4936 ( .A1(n5950), .A2(n4230), .A3(n4237), .ZN(n3954) );
  NAND2_X1 U4937 ( .A1(n3954), .A2(n3953), .ZN(n4559) );
  OAI22_X1 U4938 ( .A1(n6452), .A2(n4432), .B1(n4559), .B2(n6502), .ZN(n3955)
         );
  AOI21_X1 U4939 ( .B1(n6488), .B2(n3978), .A(n3955), .ZN(n3956) );
  OAI211_X1 U4940 ( .C1(n3981), .C2(n5292), .A(n3957), .B(n3956), .ZN(U3044)
         );
  INV_X1 U4941 ( .A(n6536), .ZN(n5329) );
  NAND2_X1 U4942 ( .A1(n3976), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3960) );
  OAI22_X1 U4943 ( .A1(n6476), .A2(n4432), .B1(n4559), .B2(n6540), .ZN(n3958)
         );
  AOI21_X1 U4944 ( .B1(n6535), .B2(n3978), .A(n3958), .ZN(n3959) );
  OAI211_X1 U4945 ( .C1(n3981), .C2(n5329), .A(n3960), .B(n3959), .ZN(U3050)
         );
  INV_X1 U4946 ( .A(n6505), .ZN(n5296) );
  NAND2_X1 U4947 ( .A1(n3976), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3963) );
  OAI22_X1 U4948 ( .A1(n6456), .A2(n4432), .B1(n4559), .B2(n6508), .ZN(n3961)
         );
  AOI21_X1 U4949 ( .B1(n6504), .B2(n3978), .A(n3961), .ZN(n3962) );
  OAI211_X1 U4950 ( .C1(n3981), .C2(n5296), .A(n3963), .B(n3962), .ZN(U3045)
         );
  INV_X1 U4951 ( .A(n6517), .ZN(n5304) );
  NAND2_X1 U4952 ( .A1(n3976), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3966) );
  OAI22_X1 U4953 ( .A1(n6520), .A2(n4432), .B1(n4559), .B2(n6462), .ZN(n3964)
         );
  AOI21_X1 U4954 ( .B1(n6516), .B2(n3978), .A(n3964), .ZN(n3965) );
  OAI211_X1 U4955 ( .C1(n3981), .C2(n5304), .A(n3966), .B(n3965), .ZN(U3047)
         );
  INV_X1 U4956 ( .A(n6511), .ZN(n5314) );
  NAND2_X1 U4957 ( .A1(n3976), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3969) );
  OAI22_X1 U4958 ( .A1(n6514), .A2(n4432), .B1(n4559), .B2(n5311), .ZN(n3967)
         );
  AOI21_X1 U4959 ( .B1(n6510), .B2(n3978), .A(n3967), .ZN(n3968) );
  OAI211_X1 U4960 ( .C1(n3981), .C2(n5314), .A(n3969), .B(n3968), .ZN(U3046)
         );
  INV_X1 U4961 ( .A(n6546), .ZN(n5300) );
  NAND2_X1 U4962 ( .A1(n3976), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3972) );
  OAI22_X1 U4963 ( .A1(n6551), .A2(n4432), .B1(n4559), .B2(n6485), .ZN(n3970)
         );
  AOI21_X1 U4964 ( .B1(n6544), .B2(n3978), .A(n3970), .ZN(n3971) );
  OAI211_X1 U4965 ( .C1(n3981), .C2(n5300), .A(n3972), .B(n3971), .ZN(U3051)
         );
  INV_X1 U4966 ( .A(n6529), .ZN(n5322) );
  NAND2_X1 U4967 ( .A1(n3976), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3975) );
  OAI22_X1 U4968 ( .A1(n6532), .A2(n4432), .B1(n4559), .B2(n6470), .ZN(n3973)
         );
  AOI21_X1 U4969 ( .B1(n6528), .B2(n3978), .A(n3973), .ZN(n3974) );
  OAI211_X1 U4970 ( .C1(n3981), .C2(n5322), .A(n3975), .B(n3974), .ZN(U3049)
         );
  INV_X1 U4971 ( .A(n6523), .ZN(n5308) );
  NAND2_X1 U4972 ( .A1(n3976), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3980) );
  OAI22_X1 U4973 ( .A1(n6526), .A2(n4432), .B1(n4559), .B2(n6466), .ZN(n3977)
         );
  AOI21_X1 U4974 ( .B1(n6522), .B2(n3978), .A(n3977), .ZN(n3979) );
  OAI211_X1 U4975 ( .C1(n3981), .C2(n5308), .A(n3980), .B(n3979), .ZN(U3048)
         );
  INV_X1 U4976 ( .A(n5852), .ZN(n5045) );
  NAND2_X1 U4977 ( .A1(n3983), .A2(n3982), .ZN(n3984) );
  NAND2_X1 U4978 ( .A1(n3989), .A2(n3984), .ZN(n6419) );
  INV_X1 U4979 ( .A(n6419), .ZN(n3985) );
  INV_X1 U4980 ( .A(n5848), .ZN(n5044) );
  AOI22_X1 U4981 ( .A1(n5045), .A2(n3985), .B1(n5044), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n3986) );
  OAI21_X1 U4982 ( .B1(n3987), .B2(n5850), .A(n3986), .ZN(U2857) );
  NAND2_X1 U4983 ( .A1(n3989), .A2(n3988), .ZN(n3990) );
  AND2_X1 U4984 ( .A1(n4063), .A2(n3990), .ZN(n6404) );
  AOI22_X1 U4985 ( .A1(n5045), .A2(n6404), .B1(n5044), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n3991) );
  OAI21_X1 U4986 ( .B1(n3992), .B2(n5850), .A(n3991), .ZN(U2856) );
  OR2_X1 U4987 ( .A1(n3993), .A2(n5457), .ZN(n3994) );
  AND2_X1 U4988 ( .A1(n3995), .A2(n3994), .ZN(n6427) );
  INV_X1 U4989 ( .A(n6427), .ZN(n3996) );
  AOI22_X1 U4990 ( .A1(n5045), .A2(n3996), .B1(n5044), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n3997) );
  OAI21_X1 U4991 ( .B1(n6230), .B2(n5850), .A(n3997), .ZN(U2858) );
  NAND2_X1 U4992 ( .A1(n3999), .A2(n3998), .ZN(n4002) );
  NAND2_X1 U4993 ( .A1(n4000), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4001)
         );
  NAND2_X1 U4994 ( .A1(n4002), .A2(n4001), .ZN(n4121) );
  OR2_X1 U4995 ( .A1(n4003), .A2(n4460), .ZN(n4006) );
  XNOR2_X1 U4996 ( .A(n4127), .B(n4125), .ZN(n4004) );
  NAND2_X1 U4997 ( .A1(n4004), .A2(n5182), .ZN(n4005) );
  NAND2_X1 U4998 ( .A1(n4006), .A2(n4005), .ZN(n4122) );
  INV_X1 U4999 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4007) );
  XNOR2_X1 U5000 ( .A(n4122), .B(n4007), .ZN(n4120) );
  XNOR2_X1 U5001 ( .A(n4121), .B(n4120), .ZN(n6397) );
  INV_X1 U5002 ( .A(n4008), .ZN(n4010) );
  AOI21_X1 U5003 ( .B1(n4011), .B2(n4010), .A(n4009), .ZN(n4061) );
  INV_X1 U5004 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6617) );
  NOR2_X1 U5005 ( .A1(n6426), .A2(n6617), .ZN(n6395) );
  AOI21_X1 U5006 ( .B1(n6363), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6395), 
        .ZN(n4012) );
  OAI21_X1 U5007 ( .B1(n6221), .B2(n6355), .A(n4012), .ZN(n4013) );
  AOI21_X1 U5008 ( .B1(n4061), .B2(n6360), .A(n4013), .ZN(n4014) );
  OAI21_X1 U5009 ( .B1(n6323), .B2(n6397), .A(n4014), .ZN(U2982) );
  NOR2_X1 U5010 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4015), .ZN(n4057)
         );
  INV_X1 U5011 ( .A(n4057), .ZN(n4016) );
  AND2_X1 U5012 ( .A1(n4023), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4531) );
  NOR2_X1 U5013 ( .A1(n4308), .A2(n5282), .ZN(n4407) );
  OAI21_X1 U5014 ( .B1(n4407), .B2(n6814), .A(n4261), .ZN(n4402) );
  AOI211_X1 U5015 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4016), .A(n4531), .B(
        n4402), .ZN(n4021) );
  INV_X1 U5016 ( .A(n4114), .ZN(n4017) );
  OAI21_X1 U5017 ( .B1(n4017), .B2(n4054), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4019) );
  INV_X1 U5018 ( .A(n4022), .ZN(n4018) );
  NAND3_X1 U5019 ( .A1(n4019), .A2(n6445), .A3(n4018), .ZN(n4020) );
  INV_X1 U5020 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4029) );
  INV_X1 U5021 ( .A(n6462), .ZN(n6515) );
  NAND2_X1 U5022 ( .A1(n4022), .A2(n5118), .ZN(n4025) );
  NOR2_X1 U5023 ( .A1(n4023), .A2(n6814), .ZN(n4403) );
  NAND2_X1 U5024 ( .A1(n4403), .A2(n4407), .ZN(n4024) );
  NAND2_X1 U5025 ( .A1(n4025), .A2(n4024), .ZN(n4053) );
  AOI22_X1 U5026 ( .A1(n4054), .A2(n6515), .B1(n6517), .B2(n4053), .ZN(n4026)
         );
  OAI21_X1 U5027 ( .B1(n6520), .B2(n4114), .A(n4026), .ZN(n4027) );
  AOI21_X1 U5028 ( .B1(n6516), .B2(n4057), .A(n4027), .ZN(n4028) );
  OAI21_X1 U5029 ( .B1(n4060), .B2(n4029), .A(n4028), .ZN(U3023) );
  INV_X1 U5030 ( .A(n6508), .ZN(n6453) );
  AOI22_X1 U5031 ( .A1(n4054), .A2(n6453), .B1(n6505), .B2(n4053), .ZN(n4030)
         );
  OAI21_X1 U5032 ( .B1(n6456), .B2(n4114), .A(n4030), .ZN(n4031) );
  AOI21_X1 U5033 ( .B1(n6504), .B2(n4057), .A(n4031), .ZN(n4032) );
  OAI21_X1 U5034 ( .B1(n4060), .B2(n4033), .A(n4032), .ZN(U3021) );
  INV_X1 U5035 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4445) );
  INV_X1 U5036 ( .A(n6485), .ZN(n6541) );
  AOI22_X1 U5037 ( .A1(n4054), .A2(n6541), .B1(n6546), .B2(n4053), .ZN(n4034)
         );
  OAI21_X1 U5038 ( .B1(n6551), .B2(n4114), .A(n4034), .ZN(n4035) );
  AOI21_X1 U5039 ( .B1(n6544), .B2(n4057), .A(n4035), .ZN(n4036) );
  OAI21_X1 U5040 ( .B1(n4060), .B2(n4445), .A(n4036), .ZN(U3027) );
  INV_X1 U5041 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4040) );
  INV_X1 U5042 ( .A(n6470), .ZN(n6527) );
  AOI22_X1 U5043 ( .A1(n4054), .A2(n6527), .B1(n6529), .B2(n4053), .ZN(n4037)
         );
  OAI21_X1 U5044 ( .B1(n6532), .B2(n4114), .A(n4037), .ZN(n4038) );
  AOI21_X1 U5045 ( .B1(n6528), .B2(n4057), .A(n4038), .ZN(n4039) );
  OAI21_X1 U5046 ( .B1(n4060), .B2(n4040), .A(n4039), .ZN(U3025) );
  INV_X1 U5047 ( .A(n6466), .ZN(n6521) );
  AOI22_X1 U5048 ( .A1(n4054), .A2(n6521), .B1(n6523), .B2(n4053), .ZN(n4041)
         );
  OAI21_X1 U5049 ( .B1(n6526), .B2(n4114), .A(n4041), .ZN(n4042) );
  AOI21_X1 U5050 ( .B1(n6522), .B2(n4057), .A(n4042), .ZN(n4043) );
  OAI21_X1 U5051 ( .B1(n4060), .B2(n4044), .A(n4043), .ZN(U3024) );
  INV_X1 U5052 ( .A(n6502), .ZN(n6440) );
  AOI22_X1 U5053 ( .A1(n4054), .A2(n6440), .B1(n6499), .B2(n4053), .ZN(n4045)
         );
  OAI21_X1 U5054 ( .B1(n6452), .B2(n4114), .A(n4045), .ZN(n4046) );
  AOI21_X1 U5055 ( .B1(n6488), .B2(n4057), .A(n4046), .ZN(n4047) );
  OAI21_X1 U5056 ( .B1(n4060), .B2(n4048), .A(n4047), .ZN(U3020) );
  INV_X1 U5057 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4052) );
  INV_X1 U5058 ( .A(n6540), .ZN(n6471) );
  AOI22_X1 U5059 ( .A1(n4054), .A2(n6471), .B1(n6536), .B2(n4053), .ZN(n4049)
         );
  OAI21_X1 U5060 ( .B1(n6476), .B2(n4114), .A(n4049), .ZN(n4050) );
  AOI21_X1 U5061 ( .B1(n6535), .B2(n4057), .A(n4050), .ZN(n4051) );
  OAI21_X1 U5062 ( .B1(n4060), .B2(n4052), .A(n4051), .ZN(U3026) );
  INV_X1 U5063 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U5064 ( .A1(n4054), .A2(n6509), .B1(n6511), .B2(n4053), .ZN(n4055)
         );
  OAI21_X1 U5065 ( .B1(n6514), .B2(n4114), .A(n4055), .ZN(n4056) );
  AOI21_X1 U5066 ( .B1(n6510), .B2(n4057), .A(n4056), .ZN(n4058) );
  OAI21_X1 U5067 ( .B1(n4060), .B2(n4059), .A(n4058), .ZN(U3022) );
  INV_X1 U5068 ( .A(n4061), .ZN(n6223) );
  XNOR2_X1 U5069 ( .A(n4063), .B(n4062), .ZN(n6396) );
  AOI22_X1 U5070 ( .A1(n5045), .A2(n6396), .B1(EBX_REG_4__SCAN_IN), .B2(n5044), 
        .ZN(n4064) );
  OAI21_X1 U5071 ( .B1(n6223), .B2(n5850), .A(n4064), .ZN(U2855) );
  NAND2_X1 U5072 ( .A1(n4181), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4229) );
  OR2_X1 U5073 ( .A1(n6674), .A2(n4229), .ZN(n4356) );
  NAND3_X1 U5074 ( .A1(n4066), .A2(n6445), .A3(STATEBS16_REG_SCAN_IN), .ZN(
        n4065) );
  INV_X1 U5075 ( .A(n6494), .ZN(n4184) );
  AOI21_X1 U5076 ( .B1(n4356), .B2(n4065), .A(n4184), .ZN(n4109) );
  INV_X1 U5077 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4077) );
  NOR2_X1 U5078 ( .A1(n6927), .A2(n4356), .ZN(n4106) );
  NAND2_X1 U5079 ( .A1(n4066), .A2(n4237), .ZN(n4267) );
  NOR2_X2 U5080 ( .A1(n4067), .A2(n4237), .ZN(n4391) );
  INV_X1 U5081 ( .A(n4182), .ZN(n4069) );
  AND2_X1 U5082 ( .A1(n4068), .A2(n5948), .ZN(n4355) );
  AND2_X1 U5083 ( .A1(n4355), .A2(n6445), .ZN(n4408) );
  NAND2_X1 U5084 ( .A1(n4069), .A2(n4408), .ZN(n4073) );
  NAND2_X1 U5085 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4070) );
  NOR2_X1 U5086 ( .A1(n4070), .A2(n4229), .ZN(n4071) );
  AOI21_X1 U5087 ( .B1(n6445), .B2(n4106), .A(n4071), .ZN(n4072) );
  NAND2_X1 U5088 ( .A1(n4073), .A2(n4072), .ZN(n4103) );
  AOI22_X1 U5089 ( .A1(n4391), .A2(n6453), .B1(n6505), .B2(n4103), .ZN(n4074)
         );
  OAI21_X1 U5090 ( .B1(n6456), .B2(n4267), .A(n4074), .ZN(n4075) );
  AOI21_X1 U5091 ( .B1(n6504), .B2(n4106), .A(n4075), .ZN(n4076) );
  OAI21_X1 U5092 ( .B1(n4109), .B2(n4077), .A(n4076), .ZN(U3125) );
  INV_X1 U5093 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U5094 ( .A1(n4391), .A2(n6541), .B1(n6546), .B2(n4103), .ZN(n4078)
         );
  OAI21_X1 U5095 ( .B1(n6551), .B2(n4267), .A(n4078), .ZN(n4079) );
  AOI21_X1 U5096 ( .B1(n6544), .B2(n4106), .A(n4079), .ZN(n4080) );
  OAI21_X1 U5097 ( .B1(n4109), .B2(n4081), .A(n4080), .ZN(U3131) );
  INV_X1 U5098 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U5099 ( .A1(n4391), .A2(n6515), .B1(n6517), .B2(n4103), .ZN(n4082)
         );
  OAI21_X1 U5100 ( .B1(n6520), .B2(n4267), .A(n4082), .ZN(n4083) );
  AOI21_X1 U5101 ( .B1(n6516), .B2(n4106), .A(n4083), .ZN(n4084) );
  OAI21_X1 U5102 ( .B1(n4109), .B2(n4085), .A(n4084), .ZN(U3127) );
  INV_X1 U5103 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U5104 ( .A1(n4391), .A2(n6440), .B1(n6499), .B2(n4103), .ZN(n4086)
         );
  OAI21_X1 U5105 ( .B1(n6452), .B2(n4267), .A(n4086), .ZN(n4087) );
  AOI21_X1 U5106 ( .B1(n6488), .B2(n4106), .A(n4087), .ZN(n4088) );
  OAI21_X1 U5107 ( .B1(n4109), .B2(n4089), .A(n4088), .ZN(U3124) );
  INV_X1 U5108 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4093) );
  AOI22_X1 U5109 ( .A1(n4391), .A2(n6509), .B1(n6511), .B2(n4103), .ZN(n4090)
         );
  OAI21_X1 U5110 ( .B1(n6514), .B2(n4267), .A(n4090), .ZN(n4091) );
  AOI21_X1 U5111 ( .B1(n6510), .B2(n4106), .A(n4091), .ZN(n4092) );
  OAI21_X1 U5112 ( .B1(n4109), .B2(n4093), .A(n4092), .ZN(U3126) );
  INV_X1 U5113 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4097) );
  AOI22_X1 U5114 ( .A1(n4391), .A2(n6521), .B1(n6523), .B2(n4103), .ZN(n4094)
         );
  OAI21_X1 U5115 ( .B1(n6526), .B2(n4267), .A(n4094), .ZN(n4095) );
  AOI21_X1 U5116 ( .B1(n6522), .B2(n4106), .A(n4095), .ZN(n4096) );
  OAI21_X1 U5117 ( .B1(n4109), .B2(n4097), .A(n4096), .ZN(U3128) );
  INV_X1 U5118 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6274) );
  OAI222_X1 U5119 ( .A1(n6223), .A2(n5862), .B1(n5109), .B2(n4098), .C1(n6274), 
        .C2(n5796), .ZN(U2887) );
  INV_X1 U5120 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5121 ( .A1(n4391), .A2(n6527), .B1(n6529), .B2(n4103), .ZN(n4099)
         );
  OAI21_X1 U5122 ( .B1(n6532), .B2(n4267), .A(n4099), .ZN(n4100) );
  AOI21_X1 U5123 ( .B1(n6528), .B2(n4106), .A(n4100), .ZN(n4101) );
  OAI21_X1 U5124 ( .B1(n4109), .B2(n4102), .A(n4101), .ZN(U3129) );
  INV_X1 U5125 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U5126 ( .A1(n4391), .A2(n6471), .B1(n6536), .B2(n4103), .ZN(n4104)
         );
  OAI21_X1 U5127 ( .B1(n6476), .B2(n4267), .A(n4104), .ZN(n4105) );
  AOI21_X1 U5128 ( .B1(n6535), .B2(n4106), .A(n4105), .ZN(n4107) );
  OAI21_X1 U5129 ( .B1(n4109), .B2(n4108), .A(n4107), .ZN(U3130) );
  INV_X1 U5130 ( .A(n6528), .ZN(n5151) );
  NAND2_X1 U5131 ( .A1(n4113), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4112) );
  OAI22_X1 U5132 ( .A1(n6470), .A2(n4114), .B1(n4525), .B2(n6532), .ZN(n4110)
         );
  AOI21_X1 U5133 ( .B1(n4116), .B2(n6529), .A(n4110), .ZN(n4111) );
  OAI211_X1 U5134 ( .C1(n4119), .C2(n5151), .A(n4112), .B(n4111), .ZN(U3033)
         );
  INV_X1 U5135 ( .A(n6535), .ZN(n5147) );
  NAND2_X1 U5136 ( .A1(n4113), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4118) );
  OAI22_X1 U5137 ( .A1(n6540), .A2(n4114), .B1(n4525), .B2(n6476), .ZN(n4115)
         );
  AOI21_X1 U5138 ( .B1(n4116), .B2(n6536), .A(n4115), .ZN(n4117) );
  OAI211_X1 U5139 ( .C1(n4119), .C2(n5147), .A(n4118), .B(n4117), .ZN(U3034)
         );
  NAND2_X1 U5140 ( .A1(n4121), .A2(n4120), .ZN(n4124) );
  NAND2_X1 U5141 ( .A1(n4122), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4123)
         );
  NAND2_X1 U5142 ( .A1(n4124), .A2(n4123), .ZN(n4170) );
  INV_X1 U5143 ( .A(n4125), .ZN(n4126) );
  NOR2_X1 U5144 ( .A1(n4127), .A2(n4126), .ZN(n4129) );
  NAND2_X1 U5145 ( .A1(n4129), .A2(n4128), .ZN(n4449) );
  OAI211_X1 U5146 ( .C1(n4129), .C2(n4128), .A(n4449), .B(n5182), .ZN(n4130)
         );
  OAI21_X1 U5147 ( .B1(n4131), .B2(n4460), .A(n4130), .ZN(n4133) );
  INV_X1 U5148 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4132) );
  XNOR2_X1 U5149 ( .A(n4133), .B(n4132), .ZN(n4171) );
  NAND2_X1 U5150 ( .A1(n4170), .A2(n4171), .ZN(n4135) );
  NAND2_X1 U5151 ( .A1(n4133), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4134)
         );
  NAND2_X1 U5152 ( .A1(n4135), .A2(n4134), .ZN(n4439) );
  AOI22_X1 U5153 ( .A1(n5691), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4139) );
  AOI22_X1 U5154 ( .A1(n5680), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5692), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U5155 ( .A1(n5688), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3607), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4137) );
  AOI22_X1 U5156 ( .A1(n5679), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4136) );
  NAND4_X1 U5157 ( .A1(n4139), .A2(n4138), .A3(n4137), .A4(n4136), .ZN(n4145)
         );
  AOI22_X1 U5158 ( .A1(n4995), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5634), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4143) );
  AOI22_X1 U5159 ( .A1(n4729), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4142) );
  AOI22_X1 U5160 ( .A1(n5682), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4141) );
  AOI22_X1 U5161 ( .A1(n3608), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4140) );
  NAND4_X1 U5162 ( .A1(n4143), .A2(n4142), .A3(n4141), .A4(n4140), .ZN(n4144)
         );
  OR2_X1 U5163 ( .A1(n4145), .A2(n4144), .ZN(n4450) );
  AOI22_X1 U5164 ( .A1(n4146), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4443), 
        .B2(n4450), .ZN(n4149) );
  INV_X1 U5165 ( .A(n4149), .ZN(n4147) );
  NAND2_X1 U5166 ( .A1(n4150), .A2(n4149), .ZN(n4215) );
  NAND3_X1 U5167 ( .A1(n4463), .A2(n4448), .A3(n4215), .ZN(n4153) );
  XNOR2_X1 U5168 ( .A(n4449), .B(n4450), .ZN(n4151) );
  NAND2_X1 U5169 ( .A1(n4151), .A2(n5182), .ZN(n4152) );
  NAND2_X1 U5170 ( .A1(n4153), .A2(n4152), .ZN(n4440) );
  INV_X1 U5171 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4154) );
  XNOR2_X1 U5172 ( .A(n4440), .B(n4154), .ZN(n4438) );
  XNOR2_X1 U5173 ( .A(n4439), .B(n4438), .ZN(n4223) );
  NAND2_X1 U5174 ( .A1(n6059), .A2(n6430), .ZN(n6374) );
  INV_X1 U5175 ( .A(n6374), .ZN(n6429) );
  OAI21_X1 U5176 ( .B1(n3858), .B2(n6431), .A(n3867), .ZN(n6418) );
  INV_X1 U5177 ( .A(n6418), .ZN(n5219) );
  NAND2_X1 U5178 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6394) );
  NOR3_X1 U5179 ( .A1(n5219), .A2(n4132), .A3(n6394), .ZN(n4165) );
  NAND2_X1 U5180 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5226) );
  INV_X1 U5181 ( .A(n6430), .ZN(n6062) );
  NOR2_X1 U5182 ( .A1(n6062), .A2(n4164), .ZN(n5229) );
  INV_X1 U5183 ( .A(n5229), .ZN(n5411) );
  AOI21_X1 U5184 ( .B1(n5226), .B2(n5411), .A(n4469), .ZN(n6424) );
  OAI21_X1 U5185 ( .B1(n6429), .B2(n4165), .A(n6424), .ZN(n4172) );
  INV_X1 U5186 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4156) );
  NAND2_X1 U5187 ( .A1(n5456), .A2(n4156), .ZN(n4160) );
  NAND2_X1 U5188 ( .A1(n3112), .A2(n4154), .ZN(n4158) );
  NAND2_X1 U5189 ( .A1(n5457), .A2(n4156), .ZN(n4157) );
  NAND3_X1 U5190 ( .A1(n4158), .A2(n5659), .A3(n4157), .ZN(n4159) );
  NAND2_X1 U5191 ( .A1(n4160), .A2(n4159), .ZN(n4161) );
  OR2_X1 U5192 ( .A1(n4162), .A2(n4161), .ZN(n4163) );
  NAND2_X1 U5193 ( .A1(n4794), .A2(n4163), .ZN(n6204) );
  NAND2_X1 U5194 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n4164), .ZN(n6063)
         );
  NAND2_X1 U5195 ( .A1(n6430), .A2(n6063), .ZN(n6415) );
  NAND3_X1 U5196 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_2__SCAN_IN), .A3(n6415), .ZN(n5220) );
  NAND2_X1 U5197 ( .A1(n6416), .A2(n5220), .ZN(n4482) );
  NAND3_X1 U5198 ( .A1(n4165), .A2(n4154), .A3(n4482), .ZN(n4167) );
  INV_X1 U5199 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6621) );
  NOR2_X1 U5200 ( .A1(n6426), .A2(n6621), .ZN(n4219) );
  INV_X1 U5201 ( .A(n4219), .ZN(n4166) );
  OAI211_X1 U5202 ( .C1(n6428), .C2(n6204), .A(n4167), .B(n4166), .ZN(n4168)
         );
  AOI21_X1 U5203 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n4172), .A(n4168), 
        .ZN(n4169) );
  OAI21_X1 U5204 ( .B1(n4223), .B2(n6406), .A(n4169), .ZN(U3012) );
  XOR2_X1 U5205 ( .A(n4171), .B(n4170), .Z(n6335) );
  NOR3_X1 U5206 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6394), .A3(n5220), 
        .ZN(n4179) );
  INV_X1 U5207 ( .A(n4172), .ZN(n4177) );
  NOR2_X1 U5208 ( .A1(n5219), .A2(n6394), .ZN(n4173) );
  AOI21_X1 U5209 ( .B1(n5222), .B2(n4173), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n4176) );
  INV_X1 U5210 ( .A(n6205), .ZN(n4174) );
  INV_X1 U5211 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6619) );
  NOR2_X1 U5212 ( .A1(n6426), .A2(n6619), .ZN(n6336) );
  AOI21_X1 U5213 ( .B1(n6405), .B2(n4174), .A(n6336), .ZN(n4175) );
  OAI21_X1 U5214 ( .B1(n4177), .B2(n4176), .A(n4175), .ZN(n4178) );
  AOI211_X1 U5215 ( .C1(n6335), .C2(n6434), .A(n4179), .B(n4178), .ZN(n4180)
         );
  INV_X1 U5216 ( .A(n4180), .ZN(U3013) );
  NAND3_X1 U5217 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6560), .A3(n4181), .ZN(n4307) );
  OR2_X1 U5218 ( .A1(n6927), .A2(n4307), .ZN(n4209) );
  NAND2_X1 U5219 ( .A1(n6490), .A2(n4230), .ZN(n4189) );
  OAI21_X1 U5220 ( .B1(n4189), .B2(n6091), .A(n5118), .ZN(n4187) );
  OR2_X1 U5221 ( .A1(n4304), .A2(n4182), .ZN(n4183) );
  AND2_X1 U5222 ( .A1(n4183), .A2(n4209), .ZN(n4188) );
  INV_X1 U5223 ( .A(n4188), .ZN(n4186) );
  AOI21_X1 U5224 ( .B1(n6492), .B2(n4307), .A(n4184), .ZN(n4185) );
  OAI21_X1 U5225 ( .B1(n4187), .B2(n4186), .A(n4185), .ZN(n4206) );
  OAI22_X1 U5226 ( .A1(n4188), .A2(n4187), .B1(n6814), .B2(n4307), .ZN(n4205)
         );
  AOI22_X1 U5227 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4206), .B1(n6517), 
        .B2(n4205), .ZN(n4192) );
  INV_X1 U5228 ( .A(n4189), .ZN(n4190) );
  AOI22_X1 U5229 ( .A1(n6515), .A2(n4346), .B1(n5283), .B2(n6459), .ZN(n4191)
         );
  OAI211_X1 U5230 ( .C1(n5139), .C2(n4209), .A(n4192), .B(n4191), .ZN(U3095)
         );
  AOI22_X1 U5231 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4206), .B1(n6523), 
        .B2(n4205), .ZN(n4194) );
  AOI22_X1 U5232 ( .A1(n6521), .A2(n4346), .B1(n5283), .B2(n6463), .ZN(n4193)
         );
  OAI211_X1 U5233 ( .C1(n5127), .C2(n4209), .A(n4194), .B(n4193), .ZN(U3096)
         );
  AOI22_X1 U5234 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4206), .B1(n6536), 
        .B2(n4205), .ZN(n4196) );
  AOI22_X1 U5235 ( .A1(n6471), .A2(n4346), .B1(n5283), .B2(n6533), .ZN(n4195)
         );
  OAI211_X1 U5236 ( .C1(n5147), .C2(n4209), .A(n4196), .B(n4195), .ZN(U3098)
         );
  AOI22_X1 U5237 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4206), .B1(n6505), 
        .B2(n4205), .ZN(n4198) );
  AOI22_X1 U5238 ( .A1(n6453), .A2(n4346), .B1(n5283), .B2(n6503), .ZN(n4197)
         );
  OAI211_X1 U5239 ( .C1(n5158), .C2(n4209), .A(n4198), .B(n4197), .ZN(U3093)
         );
  AOI22_X1 U5240 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4206), .B1(n6499), 
        .B2(n4205), .ZN(n4200) );
  AOI22_X1 U5241 ( .A1(n6440), .A2(n4346), .B1(n5283), .B2(n6487), .ZN(n4199)
         );
  OAI211_X1 U5242 ( .C1(n5135), .C2(n4209), .A(n4200), .B(n4199), .ZN(U3092)
         );
  AOI22_X1 U5243 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4206), .B1(n6511), 
        .B2(n4205), .ZN(n4202) );
  AOI22_X1 U5244 ( .A1(n6509), .A2(n4346), .B1(n5283), .B2(n5309), .ZN(n4201)
         );
  OAI211_X1 U5245 ( .C1(n5131), .C2(n4209), .A(n4202), .B(n4201), .ZN(U3094)
         );
  AOI22_X1 U5246 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4206), .B1(n6529), 
        .B2(n4205), .ZN(n4204) );
  AOI22_X1 U5247 ( .A1(n6527), .A2(n4346), .B1(n5283), .B2(n6467), .ZN(n4203)
         );
  OAI211_X1 U5248 ( .C1(n5151), .C2(n4209), .A(n4204), .B(n4203), .ZN(U3097)
         );
  AOI22_X1 U5249 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4206), .B1(n6546), 
        .B2(n4205), .ZN(n4208) );
  AOI22_X1 U5250 ( .A1(n6541), .A2(n4346), .B1(n5283), .B2(n6478), .ZN(n4207)
         );
  OAI211_X1 U5251 ( .C1(n5143), .C2(n4209), .A(n4208), .B(n4207), .ZN(U3099)
         );
  INV_X1 U5252 ( .A(n4210), .ZN(n4212) );
  INV_X1 U5253 ( .A(n4488), .ZN(n4211) );
  OAI21_X1 U5254 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n4212), .A(n4211), 
        .ZN(n6198) );
  INV_X1 U5255 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4228) );
  OAI22_X1 U5256 ( .A1(n4692), .A2(n4228), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6195), .ZN(n4213) );
  MUX2_X1 U5257 ( .A(n6198), .B(n4213), .S(n5646), .Z(n4214) );
  AOI21_X1 U5258 ( .B1(n4215), .B2(n4754), .A(n4214), .ZN(n4218) );
  OR2_X2 U5259 ( .A1(n4217), .A2(n4218), .ZN(n4869) );
  INV_X1 U5260 ( .A(n4869), .ZN(n4216) );
  AOI21_X1 U5261 ( .B1(n4218), .B2(n4217), .A(n4216), .ZN(n4224) );
  AOI21_X1 U5262 ( .B1(n6363), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n4219), 
        .ZN(n4220) );
  OAI21_X1 U5263 ( .B1(n6198), .B2(n6355), .A(n4220), .ZN(n4221) );
  AOI21_X1 U5264 ( .B1(n4224), .B2(n6360), .A(n4221), .ZN(n4222) );
  OAI21_X1 U5265 ( .B1(n6323), .B2(n4223), .A(n4222), .ZN(U2980) );
  INV_X1 U5266 ( .A(n4224), .ZN(n6200) );
  INV_X1 U5267 ( .A(n6204), .ZN(n4225) );
  AOI22_X1 U5268 ( .A1(n5045), .A2(n4225), .B1(n5044), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4226) );
  OAI21_X1 U5269 ( .B1(n6200), .B2(n5850), .A(n4226), .ZN(U2853) );
  INV_X1 U5270 ( .A(DATAI_6_), .ZN(n4227) );
  OAI222_X1 U5271 ( .A1(n6200), .A2(n5862), .B1(n5796), .B2(n4228), .C1(n5109), 
        .C2(n4227), .ZN(U2885) );
  OR2_X1 U5272 ( .A1(n4229), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4398)
         );
  NOR2_X1 U5273 ( .A1(n6927), .A2(n4398), .ZN(n4232) );
  INV_X1 U5274 ( .A(n4232), .ZN(n4303) );
  NAND2_X1 U5275 ( .A1(n5112), .A2(n4230), .ZN(n4238) );
  AOI21_X1 U5276 ( .B1(n4238), .B2(n5118), .A(n6666), .ZN(n4236) );
  INV_X1 U5277 ( .A(n4236), .ZN(n4233) );
  AND2_X1 U5278 ( .A1(n4355), .A2(n4231), .ZN(n4400) );
  AOI21_X1 U5279 ( .B1(n4400), .B2(n3110), .A(n4232), .ZN(n4235) );
  AOI22_X1 U5280 ( .A1(n4233), .A2(n4235), .B1(n4398), .B2(n6492), .ZN(n4234)
         );
  NAND2_X1 U5281 ( .A1(n6494), .A2(n4234), .ZN(n4298) );
  NAND2_X1 U5282 ( .A1(n4298), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4241) );
  OAI22_X1 U5283 ( .A1(n4236), .A2(n4235), .B1(n4398), .B2(n6814), .ZN(n4300)
         );
  OAI22_X1 U5284 ( .A1(n5113), .A2(n6551), .B1(n4399), .B2(n6485), .ZN(n4239)
         );
  AOI21_X1 U5285 ( .B1(n6546), .B2(n4300), .A(n4239), .ZN(n4240) );
  OAI211_X1 U5286 ( .C1(n4303), .C2(n5143), .A(n4241), .B(n4240), .ZN(U3067)
         );
  NAND2_X1 U5287 ( .A1(n4298), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4244) );
  OAI22_X1 U5288 ( .A1(n5113), .A2(n6476), .B1(n4399), .B2(n6540), .ZN(n4242)
         );
  AOI21_X1 U5289 ( .B1(n6536), .B2(n4300), .A(n4242), .ZN(n4243) );
  OAI211_X1 U5290 ( .C1(n4303), .C2(n5147), .A(n4244), .B(n4243), .ZN(U3066)
         );
  NAND2_X1 U5291 ( .A1(n4298), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4247) );
  OAI22_X1 U5292 ( .A1(n5113), .A2(n6532), .B1(n4399), .B2(n6470), .ZN(n4245)
         );
  AOI21_X1 U5293 ( .B1(n6529), .B2(n4300), .A(n4245), .ZN(n4246) );
  OAI211_X1 U5294 ( .C1(n4303), .C2(n5151), .A(n4247), .B(n4246), .ZN(U3065)
         );
  NAND2_X1 U5295 ( .A1(n4298), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4250) );
  OAI22_X1 U5296 ( .A1(n5113), .A2(n6514), .B1(n4399), .B2(n5311), .ZN(n4248)
         );
  AOI21_X1 U5297 ( .B1(n6511), .B2(n4300), .A(n4248), .ZN(n4249) );
  OAI211_X1 U5298 ( .C1(n4303), .C2(n5131), .A(n4250), .B(n4249), .ZN(U3062)
         );
  NAND2_X1 U5299 ( .A1(n4298), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4253) );
  OAI22_X1 U5300 ( .A1(n5113), .A2(n6456), .B1(n4399), .B2(n6508), .ZN(n4251)
         );
  AOI21_X1 U5301 ( .B1(n6505), .B2(n4300), .A(n4251), .ZN(n4252) );
  OAI211_X1 U5302 ( .C1(n4303), .C2(n5158), .A(n4253), .B(n4252), .ZN(U3061)
         );
  NAND2_X1 U5303 ( .A1(n4298), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4256) );
  OAI22_X1 U5304 ( .A1(n5113), .A2(n6526), .B1(n4399), .B2(n6466), .ZN(n4254)
         );
  AOI21_X1 U5305 ( .B1(n6523), .B2(n4300), .A(n4254), .ZN(n4255) );
  OAI211_X1 U5306 ( .C1(n4303), .C2(n5127), .A(n4256), .B(n4255), .ZN(U3064)
         );
  NAND2_X1 U5307 ( .A1(n4298), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4259) );
  OAI22_X1 U5308 ( .A1(n5113), .A2(n6520), .B1(n4399), .B2(n6462), .ZN(n4257)
         );
  AOI21_X1 U5309 ( .B1(n6517), .B2(n4300), .A(n4257), .ZN(n4258) );
  OAI211_X1 U5310 ( .C1(n4303), .C2(n5139), .A(n4259), .B(n4258), .ZN(U3063)
         );
  NOR2_X1 U5311 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4260), .ZN(n4262)
         );
  INV_X1 U5312 ( .A(n4262), .ZN(n4297) );
  AOI21_X1 U5313 ( .B1(n4267), .B2(n4292), .A(n6091), .ZN(n4266) );
  NAND2_X1 U5314 ( .A1(n5118), .A2(n5115), .ZN(n4265) );
  OAI21_X1 U5315 ( .B1(n5282), .B2(n6814), .A(n4261), .ZN(n4530) );
  NOR2_X1 U5316 ( .A1(n4403), .A2(n4530), .ZN(n5119) );
  OAI21_X1 U5317 ( .B1(n6826), .B2(n4262), .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n4263) );
  INV_X1 U5318 ( .A(n4263), .ZN(n4264) );
  OAI211_X1 U5319 ( .C1(n4266), .C2(n4265), .A(n5119), .B(n4264), .ZN(n4290)
         );
  NAND2_X1 U5320 ( .A1(n4290), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4271)
         );
  INV_X1 U5321 ( .A(n4267), .ZN(n4294) );
  NOR2_X1 U5322 ( .A1(n5115), .A2(n6492), .ZN(n5123) );
  INV_X1 U5323 ( .A(n4531), .ZN(n5121) );
  NOR2_X1 U5324 ( .A1(n5121), .A2(n6674), .ZN(n4268) );
  AOI22_X1 U5325 ( .A1(n5123), .A2(n5469), .B1(n5282), .B2(n4268), .ZN(n4291)
         );
  OAI22_X1 U5326 ( .A1(n4292), .A2(n6526), .B1(n4291), .B2(n5308), .ZN(n4269)
         );
  AOI21_X1 U5327 ( .B1(n6521), .B2(n4294), .A(n4269), .ZN(n4270) );
  OAI211_X1 U5328 ( .C1(n4297), .C2(n5127), .A(n4271), .B(n4270), .ZN(U3136)
         );
  NAND2_X1 U5329 ( .A1(n4290), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4274)
         );
  OAI22_X1 U5330 ( .A1(n4292), .A2(n6514), .B1(n4291), .B2(n5314), .ZN(n4272)
         );
  AOI21_X1 U5331 ( .B1(n6509), .B2(n4294), .A(n4272), .ZN(n4273) );
  OAI211_X1 U5332 ( .C1(n4297), .C2(n5131), .A(n4274), .B(n4273), .ZN(U3134)
         );
  NAND2_X1 U5333 ( .A1(n4290), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4277)
         );
  OAI22_X1 U5334 ( .A1(n4292), .A2(n6476), .B1(n4291), .B2(n5329), .ZN(n4275)
         );
  AOI21_X1 U5335 ( .B1(n6471), .B2(n4294), .A(n4275), .ZN(n4276) );
  OAI211_X1 U5336 ( .C1(n4297), .C2(n5147), .A(n4277), .B(n4276), .ZN(U3138)
         );
  NAND2_X1 U5337 ( .A1(n4290), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4280)
         );
  OAI22_X1 U5338 ( .A1(n4292), .A2(n6452), .B1(n4291), .B2(n5292), .ZN(n4278)
         );
  AOI21_X1 U5339 ( .B1(n6440), .B2(n4294), .A(n4278), .ZN(n4279) );
  OAI211_X1 U5340 ( .C1(n5135), .C2(n4297), .A(n4280), .B(n4279), .ZN(U3132)
         );
  NAND2_X1 U5341 ( .A1(n4290), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4283)
         );
  OAI22_X1 U5342 ( .A1(n4292), .A2(n6532), .B1(n4291), .B2(n5322), .ZN(n4281)
         );
  AOI21_X1 U5343 ( .B1(n6527), .B2(n4294), .A(n4281), .ZN(n4282) );
  OAI211_X1 U5344 ( .C1(n4297), .C2(n5151), .A(n4283), .B(n4282), .ZN(U3137)
         );
  NAND2_X1 U5345 ( .A1(n4290), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4286)
         );
  OAI22_X1 U5346 ( .A1(n4292), .A2(n6551), .B1(n4291), .B2(n5300), .ZN(n4284)
         );
  AOI21_X1 U5347 ( .B1(n6541), .B2(n4294), .A(n4284), .ZN(n4285) );
  OAI211_X1 U5348 ( .C1(n4297), .C2(n5143), .A(n4286), .B(n4285), .ZN(U3139)
         );
  NAND2_X1 U5349 ( .A1(n4290), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4289)
         );
  OAI22_X1 U5350 ( .A1(n4292), .A2(n6456), .B1(n4291), .B2(n5296), .ZN(n4287)
         );
  AOI21_X1 U5351 ( .B1(n6453), .B2(n4294), .A(n4287), .ZN(n4288) );
  OAI211_X1 U5352 ( .C1(n4297), .C2(n5158), .A(n4289), .B(n4288), .ZN(U3133)
         );
  NAND2_X1 U5353 ( .A1(n4290), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4296)
         );
  OAI22_X1 U5354 ( .A1(n4292), .A2(n6520), .B1(n4291), .B2(n5304), .ZN(n4293)
         );
  AOI21_X1 U5355 ( .B1(n6515), .B2(n4294), .A(n4293), .ZN(n4295) );
  OAI211_X1 U5356 ( .C1(n4297), .C2(n5139), .A(n4296), .B(n4295), .ZN(U3135)
         );
  NAND2_X1 U5357 ( .A1(n4298), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4302) );
  OAI22_X1 U5358 ( .A1(n6502), .A2(n4399), .B1(n5113), .B2(n6452), .ZN(n4299)
         );
  AOI21_X1 U5359 ( .B1(n6499), .B2(n4300), .A(n4299), .ZN(n4301) );
  OAI211_X1 U5360 ( .C1(n5135), .C2(n4303), .A(n4302), .B(n4301), .ZN(U3060)
         );
  NAND2_X1 U5361 ( .A1(n5112), .A2(n4352), .ZN(n6475) );
  AOI21_X1 U5362 ( .B1(n4339), .B2(n6475), .A(n6091), .ZN(n4306) );
  INV_X1 U5363 ( .A(n4304), .ZN(n4305) );
  AND2_X1 U5364 ( .A1(n4305), .A2(n5469), .ZN(n4314) );
  NOR3_X1 U5365 ( .A1(n4306), .A2(n4314), .A3(n6492), .ZN(n4312) );
  NOR2_X1 U5366 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4307), .ZN(n4347)
         );
  INV_X1 U5367 ( .A(n4308), .ZN(n4309) );
  OR2_X1 U5368 ( .A1(n4309), .A2(n5282), .ZN(n4360) );
  AOI21_X1 U5369 ( .B1(n4360), .B2(STATE2_REG_2__SCAN_IN), .A(n4310), .ZN(
        n4357) );
  OAI211_X1 U5370 ( .C1(n6826), .C2(n4347), .A(n5121), .B(n4357), .ZN(n4311)
         );
  INV_X1 U5371 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4318) );
  INV_X1 U5372 ( .A(n4360), .ZN(n4313) );
  AOI22_X1 U5373 ( .A1(n4314), .A2(n6445), .B1(n4403), .B2(n4313), .ZN(n4344)
         );
  OAI22_X1 U5374 ( .A1(n6475), .A2(n6508), .B1(n4344), .B2(n5296), .ZN(n4316)
         );
  NOR2_X1 U5375 ( .A1(n4339), .A2(n6456), .ZN(n4315) );
  AOI211_X1 U5376 ( .C1(n4347), .C2(n6504), .A(n4316), .B(n4315), .ZN(n4317)
         );
  OAI21_X1 U5377 ( .B1(n4351), .B2(n4318), .A(n4317), .ZN(U3085) );
  INV_X1 U5378 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4322) );
  OAI22_X1 U5379 ( .A1(n6475), .A2(n6466), .B1(n4344), .B2(n5308), .ZN(n4320)
         );
  NOR2_X1 U5380 ( .A1(n4339), .A2(n6526), .ZN(n4319) );
  AOI211_X1 U5381 ( .C1(n4347), .C2(n6522), .A(n4320), .B(n4319), .ZN(n4321)
         );
  OAI21_X1 U5382 ( .B1(n4351), .B2(n4322), .A(n4321), .ZN(U3088) );
  INV_X1 U5383 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4326) );
  OAI22_X1 U5384 ( .A1(n6475), .A2(n6470), .B1(n4344), .B2(n5322), .ZN(n4324)
         );
  NOR2_X1 U5385 ( .A1(n4339), .A2(n6532), .ZN(n4323) );
  AOI211_X1 U5386 ( .C1(n4347), .C2(n6528), .A(n4324), .B(n4323), .ZN(n4325)
         );
  OAI21_X1 U5387 ( .B1(n4351), .B2(n4326), .A(n4325), .ZN(U3089) );
  INV_X1 U5388 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4330) );
  OAI22_X1 U5389 ( .A1(n6475), .A2(n6540), .B1(n4344), .B2(n5329), .ZN(n4328)
         );
  NOR2_X1 U5390 ( .A1(n4339), .A2(n6476), .ZN(n4327) );
  AOI211_X1 U5391 ( .C1(n4347), .C2(n6535), .A(n4328), .B(n4327), .ZN(n4329)
         );
  OAI21_X1 U5392 ( .B1(n4351), .B2(n4330), .A(n4329), .ZN(U3090) );
  INV_X1 U5393 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4334) );
  OAI22_X1 U5394 ( .A1(n6475), .A2(n6485), .B1(n4344), .B2(n5300), .ZN(n4332)
         );
  NOR2_X1 U5395 ( .A1(n4339), .A2(n6551), .ZN(n4331) );
  AOI211_X1 U5396 ( .C1(n4347), .C2(n6544), .A(n4332), .B(n4331), .ZN(n4333)
         );
  OAI21_X1 U5397 ( .B1(n4351), .B2(n4334), .A(n4333), .ZN(U3091) );
  INV_X1 U5398 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4338) );
  OAI22_X1 U5399 ( .A1(n6475), .A2(n5311), .B1(n4344), .B2(n5314), .ZN(n4336)
         );
  NOR2_X1 U5400 ( .A1(n4339), .A2(n6514), .ZN(n4335) );
  AOI211_X1 U5401 ( .C1(n4347), .C2(n6510), .A(n4336), .B(n4335), .ZN(n4337)
         );
  OAI21_X1 U5402 ( .B1(n4351), .B2(n4338), .A(n4337), .ZN(U3086) );
  INV_X1 U5403 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4343) );
  OAI22_X1 U5404 ( .A1(n6475), .A2(n6462), .B1(n4344), .B2(n5304), .ZN(n4341)
         );
  NOR2_X1 U5405 ( .A1(n4339), .A2(n6520), .ZN(n4340) );
  AOI211_X1 U5406 ( .C1(n4347), .C2(n6516), .A(n4341), .B(n4340), .ZN(n4342)
         );
  OAI21_X1 U5407 ( .B1(n4351), .B2(n4343), .A(n4342), .ZN(U3087) );
  INV_X1 U5408 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4350) );
  OAI22_X1 U5409 ( .A1(n6475), .A2(n6502), .B1(n4344), .B2(n5292), .ZN(n4345)
         );
  AOI21_X1 U5410 ( .B1(n4346), .B2(n6487), .A(n4345), .ZN(n4349) );
  NAND2_X1 U5411 ( .A1(n6488), .A2(n4347), .ZN(n4348) );
  OAI211_X1 U5412 ( .C1(n4351), .C2(n4350), .A(n4349), .B(n4348), .ZN(U3084)
         );
  INV_X1 U5413 ( .A(n4391), .ZN(n4353) );
  NAND2_X1 U5414 ( .A1(n6490), .A2(n4352), .ZN(n6550) );
  AOI21_X1 U5415 ( .B1(n4353), .B2(n6550), .A(n6091), .ZN(n4354) );
  AOI211_X1 U5416 ( .C1(n4355), .C2(n5114), .A(n6492), .B(n4354), .ZN(n4359)
         );
  NOR2_X1 U5417 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4356), .ZN(n4394)
         );
  INV_X1 U5418 ( .A(n4403), .ZN(n5280) );
  OAI211_X1 U5419 ( .C1(n6826), .C2(n4394), .A(n5280), .B(n4357), .ZN(n4358)
         );
  INV_X1 U5420 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4365) );
  INV_X1 U5421 ( .A(n4408), .ZN(n4361) );
  INV_X1 U5422 ( .A(n5469), .ZN(n6671) );
  OAI22_X1 U5423 ( .A1(n4361), .A2(n6671), .B1(n4360), .B2(n5121), .ZN(n4390)
         );
  AOI22_X1 U5424 ( .A1(n4391), .A2(n6533), .B1(n6536), .B2(n4390), .ZN(n4362)
         );
  OAI21_X1 U5425 ( .B1(n6540), .B2(n6550), .A(n4362), .ZN(n4363) );
  AOI21_X1 U5426 ( .B1(n6535), .B2(n4394), .A(n4363), .ZN(n4364) );
  OAI21_X1 U5427 ( .B1(n4397), .B2(n4365), .A(n4364), .ZN(U3122) );
  INV_X1 U5428 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4369) );
  AOI22_X1 U5429 ( .A1(n4391), .A2(n6459), .B1(n6517), .B2(n4390), .ZN(n4366)
         );
  OAI21_X1 U5430 ( .B1(n6462), .B2(n6550), .A(n4366), .ZN(n4367) );
  AOI21_X1 U5431 ( .B1(n6516), .B2(n4394), .A(n4367), .ZN(n4368) );
  OAI21_X1 U5432 ( .B1(n4397), .B2(n4369), .A(n4368), .ZN(U3119) );
  INV_X1 U5433 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4373) );
  AOI22_X1 U5434 ( .A1(n4391), .A2(n5309), .B1(n6511), .B2(n4390), .ZN(n4370)
         );
  OAI21_X1 U5435 ( .B1(n5311), .B2(n6550), .A(n4370), .ZN(n4371) );
  AOI21_X1 U5436 ( .B1(n6510), .B2(n4394), .A(n4371), .ZN(n4372) );
  OAI21_X1 U5437 ( .B1(n4397), .B2(n4373), .A(n4372), .ZN(U3118) );
  INV_X1 U5438 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4377) );
  AOI22_X1 U5439 ( .A1(n4391), .A2(n6463), .B1(n6523), .B2(n4390), .ZN(n4374)
         );
  OAI21_X1 U5440 ( .B1(n6466), .B2(n6550), .A(n4374), .ZN(n4375) );
  AOI21_X1 U5441 ( .B1(n6522), .B2(n4394), .A(n4375), .ZN(n4376) );
  OAI21_X1 U5442 ( .B1(n4397), .B2(n4377), .A(n4376), .ZN(U3120) );
  INV_X1 U5443 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4381) );
  AOI22_X1 U5444 ( .A1(n4391), .A2(n6467), .B1(n6529), .B2(n4390), .ZN(n4378)
         );
  OAI21_X1 U5445 ( .B1(n6470), .B2(n6550), .A(n4378), .ZN(n4379) );
  AOI21_X1 U5446 ( .B1(n6528), .B2(n4394), .A(n4379), .ZN(n4380) );
  OAI21_X1 U5447 ( .B1(n4397), .B2(n4381), .A(n4380), .ZN(U3121) );
  INV_X1 U5448 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4385) );
  AOI22_X1 U5449 ( .A1(n4391), .A2(n6487), .B1(n6499), .B2(n4390), .ZN(n4382)
         );
  OAI21_X1 U5450 ( .B1(n6502), .B2(n6550), .A(n4382), .ZN(n4383) );
  AOI21_X1 U5451 ( .B1(n6488), .B2(n4394), .A(n4383), .ZN(n4384) );
  OAI21_X1 U5452 ( .B1(n4397), .B2(n4385), .A(n4384), .ZN(U3116) );
  INV_X1 U5453 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4389) );
  AOI22_X1 U5454 ( .A1(n4391), .A2(n6478), .B1(n6546), .B2(n4390), .ZN(n4386)
         );
  OAI21_X1 U5455 ( .B1(n6485), .B2(n6550), .A(n4386), .ZN(n4387) );
  AOI21_X1 U5456 ( .B1(n6544), .B2(n4394), .A(n4387), .ZN(n4388) );
  OAI21_X1 U5457 ( .B1(n4397), .B2(n4389), .A(n4388), .ZN(U3123) );
  INV_X1 U5458 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4396) );
  AOI22_X1 U5459 ( .A1(n4391), .A2(n6503), .B1(n6505), .B2(n4390), .ZN(n4392)
         );
  OAI21_X1 U5460 ( .B1(n6508), .B2(n6550), .A(n4392), .ZN(n4393) );
  AOI21_X1 U5461 ( .B1(n6504), .B2(n4394), .A(n4393), .ZN(n4395) );
  OAI21_X1 U5462 ( .B1(n4397), .B2(n4396), .A(n4395), .ZN(U3117) );
  NOR2_X1 U5463 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4398), .ZN(n4406)
         );
  INV_X1 U5464 ( .A(n4406), .ZN(n4437) );
  AOI21_X1 U5465 ( .B1(n4399), .B2(n4432), .A(n6091), .ZN(n4401) );
  NOR2_X1 U5466 ( .A1(n4401), .A2(n4400), .ZN(n4404) );
  AOI211_X1 U5467 ( .C1(n6445), .C2(n4404), .A(n4403), .B(n4402), .ZN(n4405)
         );
  NAND2_X1 U5468 ( .A1(n4430), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4411) );
  AOI22_X1 U5469 ( .A1(n4408), .A2(n6671), .B1(n4531), .B2(n4407), .ZN(n4431)
         );
  OAI22_X1 U5470 ( .A1(n4432), .A2(n6466), .B1(n4431), .B2(n5308), .ZN(n4409)
         );
  AOI21_X1 U5471 ( .B1(n6463), .B2(n4434), .A(n4409), .ZN(n4410) );
  OAI211_X1 U5472 ( .C1(n4437), .C2(n5127), .A(n4411), .B(n4410), .ZN(U3056)
         );
  NAND2_X1 U5473 ( .A1(n4430), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4414) );
  OAI22_X1 U5474 ( .A1(n4432), .A2(n6485), .B1(n4431), .B2(n5300), .ZN(n4412)
         );
  AOI21_X1 U5475 ( .B1(n6478), .B2(n4434), .A(n4412), .ZN(n4413) );
  OAI211_X1 U5476 ( .C1(n4437), .C2(n5143), .A(n4414), .B(n4413), .ZN(U3059)
         );
  NAND2_X1 U5477 ( .A1(n4430), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4417) );
  OAI22_X1 U5478 ( .A1(n4432), .A2(n6540), .B1(n4431), .B2(n5329), .ZN(n4415)
         );
  AOI21_X1 U5479 ( .B1(n6533), .B2(n4434), .A(n4415), .ZN(n4416) );
  OAI211_X1 U5480 ( .C1(n4437), .C2(n5147), .A(n4417), .B(n4416), .ZN(U3058)
         );
  NAND2_X1 U5481 ( .A1(n4430), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4420) );
  OAI22_X1 U5482 ( .A1(n4432), .A2(n6462), .B1(n4431), .B2(n5304), .ZN(n4418)
         );
  AOI21_X1 U5483 ( .B1(n6459), .B2(n4434), .A(n4418), .ZN(n4419) );
  OAI211_X1 U5484 ( .C1(n4437), .C2(n5139), .A(n4420), .B(n4419), .ZN(U3055)
         );
  NAND2_X1 U5485 ( .A1(n4430), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4423) );
  OAI22_X1 U5486 ( .A1(n4432), .A2(n6470), .B1(n4431), .B2(n5322), .ZN(n4421)
         );
  AOI21_X1 U5487 ( .B1(n6467), .B2(n4434), .A(n4421), .ZN(n4422) );
  OAI211_X1 U5488 ( .C1(n4437), .C2(n5151), .A(n4423), .B(n4422), .ZN(U3057)
         );
  NAND2_X1 U5489 ( .A1(n4430), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4426) );
  OAI22_X1 U5490 ( .A1(n4432), .A2(n5311), .B1(n4431), .B2(n5314), .ZN(n4424)
         );
  AOI21_X1 U5491 ( .B1(n5309), .B2(n4434), .A(n4424), .ZN(n4425) );
  OAI211_X1 U5492 ( .C1(n4437), .C2(n5131), .A(n4426), .B(n4425), .ZN(U3054)
         );
  NAND2_X1 U5493 ( .A1(n4430), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4429) );
  OAI22_X1 U5494 ( .A1(n4432), .A2(n6502), .B1(n4431), .B2(n5292), .ZN(n4427)
         );
  AOI21_X1 U5495 ( .B1(n6487), .B2(n4434), .A(n4427), .ZN(n4428) );
  OAI211_X1 U5496 ( .C1(n5135), .C2(n4437), .A(n4429), .B(n4428), .ZN(U3052)
         );
  NAND2_X1 U5497 ( .A1(n4430), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4436) );
  OAI22_X1 U5498 ( .A1(n4432), .A2(n6508), .B1(n4431), .B2(n5296), .ZN(n4433)
         );
  AOI21_X1 U5499 ( .B1(n6503), .B2(n4434), .A(n4433), .ZN(n4435) );
  OAI211_X1 U5500 ( .C1(n4437), .C2(n5158), .A(n4436), .B(n4435), .ZN(U3053)
         );
  NAND2_X1 U5501 ( .A1(n4439), .A2(n4438), .ZN(n4442) );
  NAND2_X1 U5502 ( .A1(n4440), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4441)
         );
  NAND2_X1 U5503 ( .A1(n4442), .A2(n4441), .ZN(n4792) );
  NAND2_X1 U5504 ( .A1(n4443), .A2(n4464), .ZN(n4444) );
  OAI21_X1 U5505 ( .B1(n4446), .B2(n4445), .A(n4444), .ZN(n4447) );
  NAND2_X1 U5506 ( .A1(n4491), .A2(n4448), .ZN(n4454) );
  INV_X1 U5507 ( .A(n4449), .ZN(n4451) );
  NAND2_X1 U5508 ( .A1(n4451), .A2(n4450), .ZN(n4466) );
  XNOR2_X1 U5509 ( .A(n4466), .B(n4464), .ZN(n4452) );
  NAND2_X1 U5510 ( .A1(n4452), .A2(n5182), .ZN(n4453) );
  NAND2_X1 U5511 ( .A1(n4454), .A2(n4453), .ZN(n4456) );
  INV_X1 U5512 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4455) );
  XNOR2_X1 U5513 ( .A(n4456), .B(n4455), .ZN(n4793) );
  NAND2_X1 U5514 ( .A1(n4792), .A2(n4793), .ZN(n4458) );
  NAND2_X1 U5515 ( .A1(n4456), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4457)
         );
  INV_X1 U5516 ( .A(n4459), .ZN(n4461) );
  NOR2_X1 U5517 ( .A1(n4461), .A2(n4460), .ZN(n4462) );
  NAND2_X1 U5518 ( .A1(n5182), .A2(n4464), .ZN(n4465) );
  OR2_X1 U5519 ( .A1(n4466), .A2(n4465), .ZN(n4467) );
  NAND2_X1 U5520 ( .A1(n5209), .A2(n4467), .ZN(n4889) );
  INV_X1 U5521 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4473) );
  XNOR2_X1 U5522 ( .A(n4889), .B(n4473), .ZN(n4887) );
  XNOR2_X1 U5523 ( .A(n4888), .B(n4887), .ZN(n4867) );
  NOR3_X1 U5524 ( .A1(n4132), .A2(n4154), .A3(n6394), .ZN(n5218) );
  OR2_X1 U5525 ( .A1(n6416), .A2(n6418), .ZN(n4468) );
  AND2_X1 U5526 ( .A1(n6424), .A2(n4468), .ZN(n6414) );
  NOR2_X1 U5527 ( .A1(n4469), .A2(n6374), .ZN(n5412) );
  AOI21_X1 U5528 ( .B1(n5218), .B2(n6414), .A(n5412), .ZN(n6373) );
  MUX2_X1 U5529 ( .A(n5569), .B(n5659), .S(EBX_REG_7__SCAN_IN), .Z(n4470) );
  NAND2_X1 U5530 ( .A1(n3116), .A2(n4470), .ZN(n4795) );
  INV_X1 U5531 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U5532 ( .A1(n5456), .A2(n6176), .ZN(n4477) );
  NAND2_X1 U5533 ( .A1(n3112), .A2(n4473), .ZN(n4475) );
  NAND2_X1 U5534 ( .A1(n5457), .A2(n6176), .ZN(n4474) );
  NAND3_X1 U5535 ( .A1(n4475), .A2(n5659), .A3(n4474), .ZN(n4476) );
  AND2_X1 U5536 ( .A1(n4477), .A2(n4476), .ZN(n4478) );
  AND2_X1 U5537 ( .A1(n4479), .A2(n4478), .ZN(n4480) );
  NOR2_X2 U5538 ( .A1(n4479), .A2(n4478), .ZN(n4825) );
  OR2_X1 U5539 ( .A1(n4480), .A2(n4825), .ZN(n6174) );
  INV_X1 U5540 ( .A(REIP_REG_8__SCAN_IN), .ZN(n4481) );
  OAI22_X1 U5541 ( .A1(n6428), .A2(n6174), .B1(n4481), .B2(n6426), .ZN(n4486)
         );
  INV_X1 U5542 ( .A(n5218), .ZN(n4483) );
  NAND2_X1 U5543 ( .A1(n6418), .A2(n4482), .ZN(n6410) );
  NOR2_X1 U5544 ( .A1(n4483), .A2(n6410), .ZN(n6376) );
  NAND2_X1 U5545 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6375) );
  OAI211_X1 U5546 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6376), .B(n6375), .ZN(n4484) );
  INV_X1 U5547 ( .A(n4484), .ZN(n4485) );
  AOI211_X1 U5548 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n6373), .A(n4486), 
        .B(n4485), .ZN(n4487) );
  OAI21_X1 U5549 ( .B1(n6406), .B2(n4867), .A(n4487), .ZN(U3010) );
  INV_X1 U5550 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4873) );
  OAI21_X1 U5551 ( .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n4488), .A(n4503), 
        .ZN(n6324) );
  AOI22_X1 U5552 ( .A1(n5706), .A2(n6324), .B1(n5784), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4489) );
  OAI21_X1 U5553 ( .B1(n4692), .B2(n4873), .A(n4489), .ZN(n4490) );
  NOR2_X2 U5554 ( .A1(n4869), .A2(n4870), .ZN(n4830) );
  AOI22_X1 U5555 ( .A1(n5629), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n5619), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4495) );
  AOI22_X1 U5556 ( .A1(n3510), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4494) );
  AOI22_X1 U5557 ( .A1(n3270), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3607), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4493) );
  AOI22_X1 U5558 ( .A1(n5683), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4492) );
  NAND4_X1 U5559 ( .A1(n4495), .A2(n4494), .A3(n4493), .A4(n4492), .ZN(n4502)
         );
  AOI22_X1 U5560 ( .A1(n4496), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4500) );
  AOI22_X1 U5561 ( .A1(n3511), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5682), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4499) );
  AOI22_X1 U5562 ( .A1(n5681), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4498) );
  AOI22_X1 U5563 ( .A1(n4729), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4497) );
  NAND4_X1 U5564 ( .A1(n4500), .A2(n4499), .A3(n4498), .A4(n4497), .ZN(n4501)
         );
  NOR2_X1 U5565 ( .A1(n4502), .A2(n4501), .ZN(n4506) );
  XNOR2_X1 U5566 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n4508), .ZN(n6178) );
  AOI22_X1 U5567 ( .A1(n5706), .A2(n6178), .B1(n5784), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4505) );
  NAND2_X1 U5568 ( .A1(n5785), .A2(EAX_REG_8__SCAN_IN), .ZN(n4504) );
  OAI211_X1 U5569 ( .C1(n4507), .C2(n4506), .A(n4505), .B(n4504), .ZN(n4829)
         );
  AND2_X4 U5570 ( .A1(n4830), .A2(n4829), .ZN(n4979) );
  INV_X1 U5571 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6163) );
  XOR2_X1 U5572 ( .A(n6163), .B(n4578), .Z(n6170) );
  AOI22_X1 U5573 ( .A1(n4995), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5683), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4512) );
  AOI22_X1 U5574 ( .A1(n5688), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4511) );
  AOI22_X1 U5575 ( .A1(n3608), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3607), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4510) );
  AOI22_X1 U5576 ( .A1(n5691), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5682), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4509) );
  NAND4_X1 U5577 ( .A1(n4512), .A2(n4511), .A3(n4510), .A4(n4509), .ZN(n4518)
         );
  AOI22_X1 U5578 ( .A1(n5681), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5679), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4516) );
  AOI22_X1 U5579 ( .A1(n5689), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4515) );
  AOI22_X1 U5580 ( .A1(n5692), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4514) );
  AOI22_X1 U5581 ( .A1(n4729), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4513) );
  NAND4_X1 U5582 ( .A1(n4516), .A2(n4515), .A3(n4514), .A4(n4513), .ZN(n4517)
         );
  OR2_X1 U5583 ( .A1(n4518), .A2(n4517), .ZN(n4519) );
  AOI22_X1 U5584 ( .A1(n4754), .A2(n4519), .B1(n5784), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4521) );
  NAND2_X1 U5585 ( .A1(n5785), .A2(EAX_REG_9__SCAN_IN), .ZN(n4520) );
  OAI211_X1 U5586 ( .C1(n6170), .C2(n5646), .A(n4521), .B(n4520), .ZN(n4919)
         );
  NAND2_X1 U5587 ( .A1(n4979), .A2(n4919), .ZN(n5035) );
  OR2_X1 U5588 ( .A1(n4979), .A2(n4919), .ZN(n4522) );
  NAND2_X1 U5589 ( .A1(n5035), .A2(n4522), .ZN(n6167) );
  AOI22_X1 U5590 ( .A1(n5039), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n6250), .ZN(n4523) );
  OAI21_X1 U5591 ( .B1(n6167), .B2(n5862), .A(n4523), .ZN(U2882) );
  NOR2_X1 U5592 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4524), .ZN(n4532)
         );
  INV_X1 U5593 ( .A(n4532), .ZN(n4564) );
  INV_X1 U5594 ( .A(n4559), .ZN(n4527) );
  OAI21_X1 U5595 ( .B1(n4561), .B2(n4527), .A(n4526), .ZN(n4529) );
  INV_X1 U5596 ( .A(n4535), .ZN(n4528) );
  AOI21_X1 U5597 ( .B1(n4529), .B2(n4528), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4533) );
  NOR2_X1 U5598 ( .A1(n4531), .A2(n4530), .ZN(n5288) );
  OAI21_X1 U5599 ( .B1(n4533), .B2(n4532), .A(n5288), .ZN(n4557) );
  NAND2_X1 U5600 ( .A1(n4557), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4538) );
  NOR2_X1 U5601 ( .A1(n5280), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4534)
         );
  AOI22_X1 U5602 ( .A1(n4535), .A2(n5118), .B1(n5282), .B2(n4534), .ZN(n4558)
         );
  OAI22_X1 U5603 ( .A1(n4559), .A2(n6514), .B1(n4558), .B2(n5314), .ZN(n4536)
         );
  AOI21_X1 U5604 ( .B1(n6509), .B2(n4561), .A(n4536), .ZN(n4537) );
  OAI211_X1 U5605 ( .C1(n4564), .C2(n5131), .A(n4538), .B(n4537), .ZN(U3038)
         );
  NAND2_X1 U5606 ( .A1(n4557), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4541) );
  OAI22_X1 U5607 ( .A1(n4559), .A2(n6456), .B1(n4558), .B2(n5296), .ZN(n4539)
         );
  AOI21_X1 U5608 ( .B1(n6453), .B2(n4561), .A(n4539), .ZN(n4540) );
  OAI211_X1 U5609 ( .C1(n4564), .C2(n5158), .A(n4541), .B(n4540), .ZN(U3037)
         );
  NAND2_X1 U5610 ( .A1(n4557), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4544) );
  OAI22_X1 U5611 ( .A1(n4559), .A2(n6551), .B1(n4558), .B2(n5300), .ZN(n4542)
         );
  AOI21_X1 U5612 ( .B1(n6541), .B2(n4561), .A(n4542), .ZN(n4543) );
  OAI211_X1 U5613 ( .C1(n4564), .C2(n5143), .A(n4544), .B(n4543), .ZN(U3043)
         );
  NAND2_X1 U5614 ( .A1(n4557), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4547) );
  OAI22_X1 U5615 ( .A1(n4559), .A2(n6532), .B1(n4558), .B2(n5322), .ZN(n4545)
         );
  AOI21_X1 U5616 ( .B1(n6527), .B2(n4561), .A(n4545), .ZN(n4546) );
  OAI211_X1 U5617 ( .C1(n4564), .C2(n5151), .A(n4547), .B(n4546), .ZN(U3041)
         );
  NAND2_X1 U5618 ( .A1(n4557), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4550) );
  OAI22_X1 U5619 ( .A1(n4559), .A2(n6476), .B1(n4558), .B2(n5329), .ZN(n4548)
         );
  AOI21_X1 U5620 ( .B1(n6471), .B2(n4561), .A(n4548), .ZN(n4549) );
  OAI211_X1 U5621 ( .C1(n4564), .C2(n5147), .A(n4550), .B(n4549), .ZN(U3042)
         );
  NAND2_X1 U5622 ( .A1(n4557), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4553) );
  OAI22_X1 U5623 ( .A1(n4559), .A2(n6452), .B1(n4558), .B2(n5292), .ZN(n4551)
         );
  AOI21_X1 U5624 ( .B1(n6440), .B2(n4561), .A(n4551), .ZN(n4552) );
  OAI211_X1 U5625 ( .C1(n5135), .C2(n4564), .A(n4553), .B(n4552), .ZN(U3036)
         );
  NAND2_X1 U5626 ( .A1(n4557), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4556) );
  OAI22_X1 U5627 ( .A1(n4559), .A2(n6526), .B1(n4558), .B2(n5308), .ZN(n4554)
         );
  AOI21_X1 U5628 ( .B1(n6521), .B2(n4561), .A(n4554), .ZN(n4555) );
  OAI211_X1 U5629 ( .C1(n4564), .C2(n5127), .A(n4556), .B(n4555), .ZN(U3040)
         );
  NAND2_X1 U5630 ( .A1(n4557), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4563) );
  OAI22_X1 U5631 ( .A1(n4559), .A2(n6520), .B1(n4558), .B2(n5304), .ZN(n4560)
         );
  AOI21_X1 U5632 ( .B1(n6515), .B2(n4561), .A(n4560), .ZN(n4562) );
  OAI211_X1 U5633 ( .C1(n4564), .C2(n5139), .A(n4563), .B(n4562), .ZN(U3039)
         );
  OR2_X1 U5634 ( .A1(n5801), .A2(n6580), .ZN(n5650) );
  AOI22_X1 U5635 ( .A1(n4995), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5683), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5636 ( .A1(n5691), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4567) );
  AOI22_X1 U5637 ( .A1(n5682), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4566) );
  AOI22_X1 U5638 ( .A1(n3241), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4565) );
  NAND4_X1 U5639 ( .A1(n4568), .A2(n4567), .A3(n4566), .A4(n4565), .ZN(n4574)
         );
  AOI22_X1 U5640 ( .A1(n5681), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n5679), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4572) );
  AOI22_X1 U5641 ( .A1(n5680), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5692), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4571) );
  AOI22_X1 U5642 ( .A1(n5688), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3607), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4570) );
  AOI22_X1 U5643 ( .A1(n3270), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4569) );
  NAND4_X1 U5644 ( .A1(n4572), .A2(n4571), .A3(n4570), .A4(n4569), .ZN(n4573)
         );
  NOR2_X1 U5645 ( .A1(n4574), .A2(n4573), .ZN(n4577) );
  INV_X1 U5646 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5900) );
  AOI21_X1 U5647 ( .B1(n5900), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4575) );
  AOI21_X1 U5648 ( .B1(n5785), .B2(EAX_REG_22__SCAN_IN), .A(n4575), .ZN(n4576)
         );
  OAI21_X1 U5649 ( .B1(n5650), .B2(n4577), .A(n4576), .ZN(n4581) );
  INV_X1 U5650 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6795) );
  INV_X1 U5651 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6912) );
  INV_X1 U5652 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6858) );
  INV_X1 U5653 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6830) );
  INV_X1 U5654 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5425) );
  XNOR2_X1 U5655 ( .A(n4963), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5993)
         );
  NAND2_X1 U5656 ( .A1(n5993), .A2(n5706), .ZN(n4580) );
  NAND2_X1 U5657 ( .A1(n4581), .A2(n4580), .ZN(n4784) );
  INV_X1 U5658 ( .A(n4784), .ZN(n4782) );
  AOI22_X1 U5659 ( .A1(n4995), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5634), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4585) );
  AOI22_X1 U5660 ( .A1(n4729), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n5629), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4584) );
  AOI22_X1 U5661 ( .A1(n3608), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5680), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4583) );
  AOI22_X1 U5662 ( .A1(n5689), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n5682), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4582) );
  NAND4_X1 U5663 ( .A1(n4585), .A2(n4584), .A3(n4583), .A4(n4582), .ZN(n4591)
         );
  AOI22_X1 U5664 ( .A1(n3510), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5692), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4589) );
  AOI22_X1 U5665 ( .A1(n3511), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4949), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4588) );
  AOI22_X1 U5666 ( .A1(n3607), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4587) );
  AOI22_X1 U5667 ( .A1(n5620), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4586) );
  NAND4_X1 U5668 ( .A1(n4589), .A2(n4588), .A3(n4587), .A4(n4586), .ZN(n4590)
         );
  NOR2_X1 U5669 ( .A1(n4591), .A2(n4590), .ZN(n4595) );
  NAND2_X1 U5670 ( .A1(n6814), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4592)
         );
  NAND2_X1 U5671 ( .A1(n5646), .A2(n4592), .ZN(n4593) );
  AOI21_X1 U5672 ( .B1(n5785), .B2(EAX_REG_21__SCAN_IN), .A(n4593), .ZN(n4594)
         );
  OAI21_X1 U5673 ( .B1(n5650), .B2(n4595), .A(n4594), .ZN(n4599) );
  OR2_X1 U5674 ( .A1(n4596), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4597)
         );
  NAND2_X1 U5675 ( .A1(n4963), .A2(n4597), .ZN(n6004) );
  OR2_X1 U5676 ( .A1(n6004), .A2(n5646), .ZN(n4598) );
  AND2_X1 U5677 ( .A1(n4599), .A2(n4598), .ZN(n4909) );
  AOI22_X1 U5678 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4729), .B1(n5080), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4603) );
  AOI22_X1 U5679 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n5680), .B1(n5692), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4602) );
  AOI22_X1 U5680 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3608), .B1(n3607), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4601) );
  AOI22_X1 U5681 ( .A1(n5689), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4949), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4600) );
  NAND4_X1 U5682 ( .A1(n4603), .A2(n4602), .A3(n4601), .A4(n4600), .ZN(n4609)
         );
  AOI22_X1 U5683 ( .A1(n3248), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5683), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4607) );
  AOI22_X1 U5684 ( .A1(n3511), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n5682), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4606) );
  AOI22_X1 U5685 ( .A1(n3510), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4605) );
  AOI22_X1 U5686 ( .A1(n5629), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4604) );
  NAND4_X1 U5687 ( .A1(n4607), .A2(n4606), .A3(n4605), .A4(n4604), .ZN(n4608)
         );
  NOR2_X1 U5688 ( .A1(n4609), .A2(n4608), .ZN(n4612) );
  OAI21_X1 U5689 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5425), .A(n5646), .ZN(
        n4610) );
  AOI21_X1 U5690 ( .B1(n5785), .B2(EAX_REG_20__SCAN_IN), .A(n4610), .ZN(n4611)
         );
  OAI21_X1 U5691 ( .B1(n5650), .B2(n4612), .A(n4611), .ZN(n4614) );
  XNOR2_X1 U5692 ( .A(n4629), .B(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6020)
         );
  NAND2_X1 U5693 ( .A1(n6020), .A2(n5706), .ZN(n4613) );
  AND2_X1 U5694 ( .A1(n4614), .A2(n4613), .ZN(n4884) );
  AOI22_X1 U5695 ( .A1(n4496), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4618) );
  AOI22_X1 U5696 ( .A1(n3510), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4729), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4617) );
  AOI22_X1 U5697 ( .A1(n5682), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4949), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4616) );
  AOI22_X1 U5698 ( .A1(n3608), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4615) );
  NAND4_X1 U5699 ( .A1(n4618), .A2(n4617), .A3(n4616), .A4(n4615), .ZN(n4624)
         );
  AOI22_X1 U5700 ( .A1(n5683), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5691), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4622) );
  AOI22_X1 U5701 ( .A1(n5620), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n5692), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4621) );
  AOI22_X1 U5702 ( .A1(n4728), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3607), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4620) );
  AOI22_X1 U5703 ( .A1(n5629), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4619) );
  NAND4_X1 U5704 ( .A1(n4622), .A2(n4621), .A3(n4620), .A4(n4619), .ZN(n4623)
         );
  NOR2_X1 U5705 ( .A1(n4624), .A2(n4623), .ZN(n4628) );
  NAND2_X1 U5706 ( .A1(n6814), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4625)
         );
  NAND2_X1 U5707 ( .A1(n5646), .A2(n4625), .ZN(n4626) );
  AOI21_X1 U5708 ( .B1(n5785), .B2(EAX_REG_19__SCAN_IN), .A(n4626), .ZN(n4627)
         );
  OAI21_X1 U5709 ( .B1(n5650), .B2(n4628), .A(n4627), .ZN(n4632) );
  OAI21_X1 U5710 ( .B1(n4630), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n4629), 
        .ZN(n6026) );
  OR2_X1 U5711 ( .A1(n6026), .A2(n5646), .ZN(n4631) );
  NAND2_X1 U5712 ( .A1(n4632), .A2(n4631), .ZN(n4981) );
  INV_X1 U5713 ( .A(n4981), .ZN(n4781) );
  AOI22_X1 U5714 ( .A1(n4995), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5683), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4636) );
  AOI22_X1 U5715 ( .A1(n5688), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4635) );
  AOI22_X1 U5716 ( .A1(n5691), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4949), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4634) );
  AOI22_X1 U5717 ( .A1(n3608), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4633) );
  NAND4_X1 U5718 ( .A1(n4636), .A2(n4635), .A3(n4634), .A4(n4633), .ZN(n4642)
         );
  AOI22_X1 U5719 ( .A1(n5620), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n5679), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4640) );
  AOI22_X1 U5720 ( .A1(n5692), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3607), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4639) );
  AOI22_X1 U5721 ( .A1(n5689), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5682), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4638) );
  AOI22_X1 U5722 ( .A1(n4729), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4637) );
  NAND4_X1 U5723 ( .A1(n4640), .A2(n4639), .A3(n4638), .A4(n4637), .ZN(n4641)
         );
  NOR2_X1 U5724 ( .A1(n4642), .A2(n4641), .ZN(n4646) );
  NAND2_X1 U5725 ( .A1(n6814), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4643)
         );
  NAND2_X1 U5726 ( .A1(n5646), .A2(n4643), .ZN(n4644) );
  AOI21_X1 U5727 ( .B1(n5785), .B2(EAX_REG_17__SCAN_IN), .A(n4644), .ZN(n4645)
         );
  OAI21_X1 U5728 ( .B1(n5650), .B2(n4646), .A(n4645), .ZN(n4648) );
  OAI21_X1 U5729 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n4659), .A(n4777), 
        .ZN(n6127) );
  OR2_X1 U5730 ( .A1(n5646), .A2(n6127), .ZN(n4647) );
  AND2_X1 U5731 ( .A1(n4648), .A2(n4647), .ZN(n4931) );
  AOI22_X1 U5732 ( .A1(n4995), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4652) );
  AOI22_X1 U5733 ( .A1(n3608), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4651) );
  AOI22_X1 U5734 ( .A1(n5691), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5682), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4650) );
  AOI22_X1 U5735 ( .A1(n4949), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4649) );
  NAND4_X1 U5736 ( .A1(n4652), .A2(n4651), .A3(n4650), .A4(n4649), .ZN(n4658)
         );
  AOI22_X1 U5737 ( .A1(n5683), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4729), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4656) );
  AOI22_X1 U5738 ( .A1(n5688), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5680), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4655) );
  AOI22_X1 U5739 ( .A1(n5679), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5692), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4654) );
  AOI22_X1 U5740 ( .A1(n3607), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4653) );
  NAND4_X1 U5741 ( .A1(n4656), .A2(n4655), .A3(n4654), .A4(n4653), .ZN(n4657)
         );
  NOR2_X1 U5742 ( .A1(n4658), .A2(n4657), .ZN(n4662) );
  AOI21_X1 U5743 ( .B1(n6795), .B2(n4757), .A(n4659), .ZN(n6131) );
  AOI21_X1 U5744 ( .B1(n5785), .B2(EAX_REG_16__SCAN_IN), .A(n4660), .ZN(n4661)
         );
  OAI21_X1 U5745 ( .B1(n5650), .B2(n4662), .A(n4661), .ZN(n4878) );
  AOI22_X1 U5746 ( .A1(n4995), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4666) );
  AOI22_X1 U5747 ( .A1(n3608), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5692), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4665) );
  AOI22_X1 U5748 ( .A1(n5691), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4664) );
  AOI22_X1 U5749 ( .A1(n5620), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4663) );
  NAND4_X1 U5750 ( .A1(n4666), .A2(n4665), .A3(n4664), .A4(n4663), .ZN(n4672)
         );
  AOI22_X1 U5751 ( .A1(n4729), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n5629), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4670) );
  AOI22_X1 U5752 ( .A1(n5688), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4728), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4669) );
  AOI22_X1 U5753 ( .A1(n5683), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5682), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4668) );
  AOI22_X1 U5754 ( .A1(n3607), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4667) );
  NAND4_X1 U5755 ( .A1(n4670), .A2(n4669), .A3(n4668), .A4(n4667), .ZN(n4671)
         );
  OAI21_X1 U5756 ( .B1(n4672), .B2(n4671), .A(n4754), .ZN(n4678) );
  NAND2_X1 U5757 ( .A1(n5785), .A2(EAX_REG_14__SCAN_IN), .ZN(n4677) );
  INV_X1 U5758 ( .A(n4673), .ZN(n4675) );
  INV_X1 U5759 ( .A(n4758), .ZN(n4674) );
  OAI21_X1 U5760 ( .B1(PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n4675), .A(n4674), 
        .ZN(n5542) );
  AOI22_X1 U5761 ( .A1(n5706), .A2(n5542), .B1(n5784), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4676) );
  AND3_X1 U5762 ( .A1(n4678), .A2(n4677), .A3(n4676), .ZN(n4803) );
  INV_X1 U5763 ( .A(n4803), .ZN(n4745) );
  INV_X1 U5764 ( .A(EAX_REG_13__SCAN_IN), .ZN(n4926) );
  AOI22_X1 U5765 ( .A1(n4995), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5691), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4682) );
  AOI22_X1 U5766 ( .A1(n5629), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n5680), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4681) );
  AOI22_X1 U5767 ( .A1(n4729), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4680) );
  AOI22_X1 U5768 ( .A1(n5688), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4679) );
  NAND4_X1 U5769 ( .A1(n4682), .A2(n4681), .A3(n4680), .A4(n4679), .ZN(n4688)
         );
  AOI22_X1 U5770 ( .A1(n5683), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4686) );
  AOI22_X1 U5771 ( .A1(n5620), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5692), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4685) );
  AOI22_X1 U5772 ( .A1(n3608), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3607), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4684) );
  AOI22_X1 U5773 ( .A1(n5682), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4683) );
  NAND4_X1 U5774 ( .A1(n4686), .A2(n4685), .A3(n4684), .A4(n4683), .ZN(n4687)
         );
  OAI21_X1 U5775 ( .B1(n4688), .B2(n4687), .A(n4754), .ZN(n4691) );
  XOR2_X1 U5776 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n4704), .Z(n6152) );
  INV_X1 U5777 ( .A(n6152), .ZN(n4689) );
  AOI22_X1 U5778 ( .A1(n5706), .A2(n4689), .B1(n5784), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4690) );
  OAI211_X1 U5779 ( .C1(n4692), .C2(n4926), .A(n4691), .B(n4690), .ZN(n4922)
         );
  INV_X1 U5780 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5110) );
  OAI22_X1 U5781 ( .A1(n4692), .A2(n5110), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6858), .ZN(n4693) );
  NAND2_X1 U5782 ( .A1(n4693), .A2(n5646), .ZN(n4708) );
  AOI22_X1 U5783 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n4729), .B1(n5679), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4697) );
  AOI22_X1 U5784 ( .A1(n4728), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5692), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4696) );
  AOI22_X1 U5785 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3608), .B1(n3607), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4695) );
  AOI22_X1 U5786 ( .A1(n5691), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4694) );
  NAND4_X1 U5787 ( .A1(n4697), .A2(n4696), .A3(n4695), .A4(n4694), .ZN(n4703)
         );
  AOI22_X1 U5788 ( .A1(n4995), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5683), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4701) );
  AOI22_X1 U5789 ( .A1(n5689), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n5682), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4700) );
  AOI22_X1 U5790 ( .A1(n5688), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4699) );
  AOI22_X1 U5791 ( .A1(n5681), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4698) );
  NAND4_X1 U5792 ( .A1(n4701), .A2(n4700), .A3(n4699), .A4(n4698), .ZN(n4702)
         );
  OR2_X1 U5793 ( .A1(n4703), .A2(n4702), .ZN(n4706) );
  AOI21_X1 U5794 ( .B1(n6858), .B2(n4720), .A(n4704), .ZN(n5348) );
  NOR2_X1 U5795 ( .A1(n5348), .A2(n5646), .ZN(n4705) );
  AOI21_X1 U5796 ( .B1(n4754), .B2(n4706), .A(n4705), .ZN(n4707) );
  AND2_X1 U5797 ( .A1(n4708), .A2(n4707), .ZN(n5108) );
  AOI22_X1 U5798 ( .A1(n5683), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4713) );
  AOI22_X1 U5799 ( .A1(n5680), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5692), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4712) );
  AOI22_X1 U5800 ( .A1(n4729), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4711) );
  AOI22_X1 U5801 ( .A1(n3608), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4710) );
  NAND4_X1 U5802 ( .A1(n4713), .A2(n4712), .A3(n4711), .A4(n4710), .ZN(n4719)
         );
  AOI22_X1 U5803 ( .A1(n4995), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5691), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4717) );
  AOI22_X1 U5804 ( .A1(n5620), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5679), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4716) );
  AOI22_X1 U5805 ( .A1(n5688), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3607), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4715) );
  AOI22_X1 U5806 ( .A1(n5682), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4714) );
  NAND4_X1 U5807 ( .A1(n4717), .A2(n4716), .A3(n4715), .A4(n4714), .ZN(n4718)
         );
  OAI21_X1 U5808 ( .B1(n4719), .B2(n4718), .A(n4754), .ZN(n4723) );
  NAND2_X1 U5809 ( .A1(n5785), .A2(EAX_REG_11__SCAN_IN), .ZN(n4722) );
  OAI21_X1 U5810 ( .B1(PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n4725), .A(n4720), 
        .ZN(n6318) );
  AOI22_X1 U5811 ( .A1(n5706), .A2(n6318), .B1(n5784), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4721) );
  AND3_X1 U5812 ( .A1(n4723), .A2(n4722), .A3(n4721), .ZN(n5036) );
  NAND2_X1 U5813 ( .A1(n4724), .A2(n6830), .ZN(n4727) );
  INV_X1 U5814 ( .A(n4725), .ZN(n4726) );
  NAND2_X1 U5815 ( .A1(n4727), .A2(n4726), .ZN(n5359) );
  AOI22_X1 U5816 ( .A1(n4995), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5691), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4733) );
  AOI22_X1 U5817 ( .A1(n5620), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5629), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4732) );
  AOI22_X1 U5818 ( .A1(n4728), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3501), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4731) );
  AOI22_X1 U5819 ( .A1(n4729), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n5682), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4730) );
  NAND4_X1 U5820 ( .A1(n4733), .A2(n4732), .A3(n4731), .A4(n4730), .ZN(n4739)
         );
  AOI22_X1 U5821 ( .A1(n5683), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4737) );
  AOI22_X1 U5822 ( .A1(n5688), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5692), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4736) );
  AOI22_X1 U5823 ( .A1(n4949), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4735) );
  AOI22_X1 U5824 ( .A1(n3608), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4734) );
  NAND4_X1 U5825 ( .A1(n4737), .A2(n4736), .A3(n4735), .A4(n4734), .ZN(n4738)
         );
  OAI21_X1 U5826 ( .B1(n4739), .B2(n4738), .A(n4754), .ZN(n4742) );
  NAND2_X1 U5827 ( .A1(n5785), .A2(EAX_REG_10__SCAN_IN), .ZN(n4741) );
  NAND2_X1 U5828 ( .A1(n5784), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4740)
         );
  NAND3_X1 U5829 ( .A1(n4742), .A2(n4741), .A3(n4740), .ZN(n4743) );
  AOI21_X1 U5830 ( .B1(n5706), .B2(n5359), .A(n4743), .ZN(n4927) );
  OR2_X1 U5831 ( .A1(n5036), .A2(n4927), .ZN(n5034) );
  NOR2_X1 U5832 ( .A1(n5108), .A2(n5034), .ZN(n4920) );
  AND2_X1 U5833 ( .A1(n4922), .A2(n4920), .ZN(n4744) );
  AND2_X1 U5834 ( .A1(n4744), .A2(n4919), .ZN(n4802) );
  AND2_X1 U5835 ( .A1(n4745), .A2(n4802), .ZN(n4801) );
  AOI22_X1 U5836 ( .A1(n5634), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5691), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4749) );
  AOI22_X1 U5837 ( .A1(n3608), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5680), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4748) );
  AOI22_X1 U5838 ( .A1(n5629), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n5619), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4747) );
  AOI22_X1 U5839 ( .A1(n4729), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n5682), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4746) );
  NAND4_X1 U5840 ( .A1(n4749), .A2(n4748), .A3(n4747), .A4(n4746), .ZN(n4756)
         );
  AOI22_X1 U5841 ( .A1(n4995), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4753) );
  AOI22_X1 U5842 ( .A1(n5688), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5080), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4752) );
  AOI22_X1 U5843 ( .A1(n4949), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4751) );
  AOI22_X1 U5844 ( .A1(n3607), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4750) );
  NAND4_X1 U5845 ( .A1(n4753), .A2(n4752), .A3(n4751), .A4(n4750), .ZN(n4755)
         );
  OAI21_X1 U5846 ( .B1(n4756), .B2(n4755), .A(n4754), .ZN(n4761) );
  NAND2_X1 U5847 ( .A1(n5785), .A2(EAX_REG_15__SCAN_IN), .ZN(n4760) );
  OAI21_X1 U5848 ( .B1(PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n4758), .A(n4757), 
        .ZN(n6143) );
  AOI22_X1 U5849 ( .A1(n5706), .A2(n6143), .B1(n5784), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4759) );
  AND3_X1 U5850 ( .A1(n4761), .A2(n4760), .A3(n4759), .ZN(n4898) );
  INV_X1 U5851 ( .A(n4898), .ZN(n4762) );
  AND2_X1 U5852 ( .A1(n4801), .A2(n4762), .ZN(n4875) );
  AND2_X1 U5853 ( .A1(n4878), .A2(n4875), .ZN(n4876) );
  AND2_X1 U5854 ( .A1(n4931), .A2(n4876), .ZN(n4930) );
  AOI22_X1 U5855 ( .A1(n5620), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n5629), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4766) );
  AOI22_X1 U5856 ( .A1(n5680), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5619), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4765) );
  AOI22_X1 U5857 ( .A1(n5688), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3607), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4764) );
  AOI22_X1 U5858 ( .A1(n3608), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4763) );
  NAND4_X1 U5859 ( .A1(n4766), .A2(n4765), .A3(n4764), .A4(n4763), .ZN(n4772)
         );
  AOI22_X1 U5860 ( .A1(n4995), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5634), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4770) );
  AOI22_X1 U5861 ( .A1(n5691), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4769) );
  AOI22_X1 U5862 ( .A1(n5682), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4768) );
  AOI22_X1 U5863 ( .A1(n4729), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4767) );
  NAND4_X1 U5864 ( .A1(n4770), .A2(n4769), .A3(n4768), .A4(n4767), .ZN(n4771)
         );
  NOR2_X1 U5865 ( .A1(n4772), .A2(n4771), .ZN(n4776) );
  INV_X1 U5866 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4773) );
  AOI21_X1 U5867 ( .B1(n4773), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4774) );
  AOI21_X1 U5868 ( .B1(n5785), .B2(EAX_REG_18__SCAN_IN), .A(n4774), .ZN(n4775)
         );
  OAI21_X1 U5869 ( .B1(n5650), .B2(n4776), .A(n4775), .ZN(n4779) );
  XNOR2_X1 U5870 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4777), .ZN(n6115)
         );
  NAND2_X1 U5871 ( .A1(n5706), .A2(n6115), .ZN(n4778) );
  NAND2_X1 U5872 ( .A1(n4779), .A2(n4778), .ZN(n5050) );
  INV_X1 U5873 ( .A(n5050), .ZN(n4780) );
  AND2_X1 U5874 ( .A1(n4930), .A2(n4780), .ZN(n4978) );
  AND2_X1 U5875 ( .A1(n4781), .A2(n4978), .ZN(n4881) );
  AND2_X1 U5876 ( .A1(n4884), .A2(n4881), .ZN(n4882) );
  NAND2_X1 U5877 ( .A1(n4979), .A2(n4971), .ZN(n4974) );
  NAND2_X1 U5878 ( .A1(n4979), .A2(n4783), .ZN(n4912) );
  NAND2_X1 U5879 ( .A1(n4912), .A2(n4784), .ZN(n4785) );
  NAND2_X1 U5880 ( .A1(n4974), .A2(n4785), .ZN(n6000) );
  NOR2_X2 U5881 ( .A1(n6250), .A2(n4786), .ZN(n6247) );
  AOI22_X1 U5882 ( .A1(n6247), .A2(DATAI_22_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n6250), .ZN(n4791) );
  AND2_X1 U5883 ( .A1(n4788), .A2(n4787), .ZN(n4789) );
  NAND2_X1 U5884 ( .A1(n6251), .A2(DATAI_6_), .ZN(n4790) );
  OAI211_X1 U5885 ( .C1(n6000), .C2(n5862), .A(n4791), .B(n4790), .ZN(U2869)
         );
  INV_X1 U5886 ( .A(n6376), .ZN(n4800) );
  XOR2_X1 U5887 ( .A(n4793), .B(n4792), .Z(n6327) );
  NAND2_X1 U5888 ( .A1(n6327), .A2(n6434), .ZN(n4799) );
  XOR2_X1 U5889 ( .A(n4795), .B(n4794), .Z(n6186) );
  INV_X1 U5890 ( .A(n6186), .ZN(n4871) );
  INV_X1 U5891 ( .A(REIP_REG_7__SCAN_IN), .ZN(n4796) );
  OR2_X1 U5892 ( .A1(n6426), .A2(n4796), .ZN(n6328) );
  OAI21_X1 U5893 ( .B1(n4871), .B2(n6428), .A(n6328), .ZN(n4797) );
  AOI21_X1 U5894 ( .B1(n6373), .B2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n4797), 
        .ZN(n4798) );
  OAI211_X1 U5895 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n4800), .A(n4799), 
        .B(n4798), .ZN(U3011) );
  NAND2_X1 U5896 ( .A1(n4979), .A2(n4801), .ZN(n4897) );
  NAND2_X1 U5897 ( .A1(n4979), .A2(n4802), .ZN(n4924) );
  NAND2_X1 U5898 ( .A1(n4924), .A2(n4803), .ZN(n4804) );
  NAND2_X1 U5899 ( .A1(n4897), .A2(n4804), .ZN(n5546) );
  AOI22_X1 U5900 ( .A1(n5039), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n6250), .ZN(n4805) );
  OAI21_X1 U5901 ( .B1(n5546), .B2(n5862), .A(n4805), .ZN(U2877) );
  MUX2_X1 U5902 ( .A(n5662), .B(n3112), .S(EBX_REG_14__SCAN_IN), .Z(n4808) );
  NAND2_X1 U5903 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5773), .ZN(n4806) );
  AND2_X1 U5904 ( .A1(n5059), .A2(n4806), .ZN(n4807) );
  NAND2_X1 U5905 ( .A1(n4808), .A2(n4807), .ZN(n4900) );
  MUX2_X1 U5906 ( .A(n5569), .B(n5659), .S(EBX_REG_9__SCAN_IN), .Z(n4809) );
  INV_X1 U5907 ( .A(n4809), .ZN(n4811) );
  NOR2_X1 U5908 ( .A1(n5774), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4810)
         );
  NOR2_X1 U5909 ( .A1(n4811), .A2(n4810), .ZN(n4824) );
  AND2_X2 U5910 ( .A1(n4825), .A2(n4824), .ZN(n5024) );
  MUX2_X1 U5911 ( .A(n5662), .B(n3112), .S(EBX_REG_10__SCAN_IN), .Z(n4814) );
  NAND2_X1 U5912 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n5773), .ZN(n4812) );
  AND2_X1 U5913 ( .A1(n5059), .A2(n4812), .ZN(n4813) );
  NAND2_X1 U5914 ( .A1(n4814), .A2(n4813), .ZN(n5023) );
  NAND2_X1 U5915 ( .A1(n5659), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4815) );
  OAI211_X1 U5916 ( .C1(n5773), .C2(EBX_REG_11__SCAN_IN), .A(n3112), .B(n4815), 
        .ZN(n4816) );
  OAI21_X1 U5917 ( .B1(n5569), .B2(EBX_REG_11__SCAN_IN), .A(n4816), .ZN(n5041)
         );
  MUX2_X1 U5918 ( .A(n5456), .B(n4856), .S(EBX_REG_12__SCAN_IN), .Z(n4819) );
  NAND2_X1 U5919 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n5773), .ZN(n4817) );
  NAND2_X1 U5920 ( .A1(n5059), .A2(n4817), .ZN(n4818) );
  NOR2_X1 U5921 ( .A1(n4819), .A2(n4818), .ZN(n5315) );
  INV_X1 U5922 ( .A(n5569), .ZN(n5012) );
  INV_X1 U5923 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U5924 ( .A1(n5012), .A2(n6150), .ZN(n4822) );
  NAND2_X1 U5925 ( .A1(n4155), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4820) );
  OAI211_X1 U5926 ( .C1(n5773), .C2(EBX_REG_13__SCAN_IN), .A(n3112), .B(n4820), 
        .ZN(n4821) );
  AND2_X1 U5927 ( .A1(n4822), .A2(n4821), .ZN(n5100) );
  AND2_X2 U5928 ( .A1(n5317), .A2(n5100), .ZN(n5102) );
  XOR2_X1 U5929 ( .A(n4900), .B(n5102), .Z(n6057) );
  AOI22_X1 U5930 ( .A1(n6057), .A2(n5045), .B1(EBX_REG_14__SCAN_IN), .B2(n5044), .ZN(n4823) );
  OAI21_X1 U5931 ( .B1(n5546), .B2(n5850), .A(n4823), .ZN(U2845) );
  INV_X1 U5932 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4828) );
  INV_X1 U5933 ( .A(n4824), .ZN(n4827) );
  INV_X1 U5934 ( .A(n4825), .ZN(n4826) );
  AOI21_X1 U5935 ( .B1(n4827), .B2(n4826), .A(n5024), .ZN(n6161) );
  INV_X1 U5936 ( .A(n6161), .ZN(n6387) );
  OAI222_X1 U5937 ( .A1(n6167), .A2(n5850), .B1(n5848), .B2(n4828), .C1(n6387), 
        .C2(n5852), .ZN(U2850) );
  INV_X1 U5938 ( .A(n4829), .ZN(n4832) );
  INV_X1 U5939 ( .A(n4868), .ZN(n4831) );
  AOI21_X1 U5940 ( .B1(n4832), .B2(n4831), .A(n4979), .ZN(n6180) );
  INV_X1 U5941 ( .A(n6180), .ZN(n4834) );
  AOI22_X1 U5942 ( .A1(n5039), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n6250), .ZN(n4833) );
  OAI21_X1 U5943 ( .B1(n4834), .B2(n5862), .A(n4833), .ZN(U2883) );
  OAI22_X1 U5944 ( .A1(n6174), .A2(n5852), .B1(n6176), .B2(n5848), .ZN(n4835)
         );
  AOI21_X1 U5945 ( .B1(n6180), .B2(n5104), .A(n4835), .ZN(n4836) );
  INV_X1 U5946 ( .A(n4836), .ZN(U2851) );
  INV_X1 U5947 ( .A(EBX_REG_22__SCAN_IN), .ZN(n4863) );
  INV_X1 U5948 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U5949 ( .A1(n5012), .A2(n6140), .ZN(n4839) );
  NAND2_X1 U5950 ( .A1(n5659), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4837) );
  OAI211_X1 U5951 ( .C1(n5773), .C2(EBX_REG_15__SCAN_IN), .A(n3112), .B(n4837), 
        .ZN(n4838) );
  AND2_X1 U5952 ( .A1(n4839), .A2(n4838), .ZN(n4899) );
  AND2_X1 U5953 ( .A1(n4900), .A2(n4899), .ZN(n4840) );
  MUX2_X1 U5954 ( .A(n5456), .B(n4856), .S(EBX_REG_16__SCAN_IN), .Z(n4842) );
  INV_X1 U5955 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5448) );
  OAI21_X1 U5956 ( .B1(n5457), .B2(n5448), .A(n5059), .ZN(n4841) );
  NOR2_X1 U5957 ( .A1(n4842), .A2(n4841), .ZN(n4915) );
  OR2_X2 U5958 ( .A1(n4916), .A2(n4915), .ZN(n4935) );
  INV_X1 U5959 ( .A(EBX_REG_19__SCAN_IN), .ZN(n4986) );
  NAND2_X1 U5960 ( .A1(n5456), .A2(n4986), .ZN(n4846) );
  INV_X1 U5961 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U5962 ( .A1(n3112), .A2(n5431), .ZN(n4844) );
  NAND2_X1 U5963 ( .A1(n5457), .A2(n4986), .ZN(n4843) );
  NAND3_X1 U5964 ( .A1(n4844), .A2(n5659), .A3(n4843), .ZN(n4845) );
  AND2_X1 U5965 ( .A1(n4846), .A2(n4845), .ZN(n4985) );
  NAND2_X1 U5966 ( .A1(n5659), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4847) );
  OAI211_X1 U5967 ( .C1(n5773), .C2(EBX_REG_17__SCAN_IN), .A(n3112), .B(n4847), 
        .ZN(n4848) );
  OAI21_X1 U5968 ( .B1(n5569), .B2(EBX_REG_17__SCAN_IN), .A(n4848), .ZN(n4934)
         );
  OR2_X1 U5969 ( .A1(n4985), .A2(n4934), .ZN(n4849) );
  NOR2_X2 U5970 ( .A1(n4935), .A2(n4849), .ZN(n4904) );
  AND2_X1 U5971 ( .A1(n5773), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4850)
         );
  AOI21_X1 U5972 ( .B1(n5774), .B2(EBX_REG_18__SCAN_IN), .A(n4850), .ZN(n4905)
         );
  INV_X1 U5973 ( .A(n4905), .ZN(n4851) );
  AND2_X1 U5974 ( .A1(n4851), .A2(n5659), .ZN(n4982) );
  AND2_X1 U5975 ( .A1(n4905), .A2(n5769), .ZN(n4983) );
  OR2_X1 U5976 ( .A1(n5774), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4853)
         );
  INV_X1 U5977 ( .A(EBX_REG_20__SCAN_IN), .ZN(n4908) );
  NAND2_X1 U5978 ( .A1(n5457), .A2(n4908), .ZN(n4852) );
  NAND2_X1 U5979 ( .A1(n4853), .A2(n4852), .ZN(n4906) );
  MUX2_X1 U5980 ( .A(n4982), .B(n4983), .S(n4906), .Z(n4854) );
  NAND2_X1 U5981 ( .A1(n4904), .A2(n4854), .ZN(n5068) );
  MUX2_X1 U5982 ( .A(n5569), .B(n5659), .S(EBX_REG_21__SCAN_IN), .Z(n4855) );
  OAI21_X1 U5983 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5774), .A(n4855), 
        .ZN(n5067) );
  OR2_X2 U5984 ( .A1(n5068), .A2(n5067), .ZN(n5070) );
  MUX2_X1 U5985 ( .A(n5456), .B(n4856), .S(EBX_REG_22__SCAN_IN), .Z(n4859) );
  NAND2_X1 U5986 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n5773), .ZN(n4857) );
  NAND2_X1 U5987 ( .A1(n5059), .A2(n4857), .ZN(n4858) );
  NOR2_X1 U5988 ( .A1(n4859), .A2(n4858), .ZN(n4860) );
  INV_X1 U5989 ( .A(n5017), .ZN(n4862) );
  NAND2_X1 U5990 ( .A1(n5070), .A2(n4860), .ZN(n4861) );
  NAND2_X1 U5991 ( .A1(n4862), .A2(n4861), .ZN(n6003) );
  OAI222_X1 U5992 ( .A1(n5850), .A2(n6000), .B1(n5848), .B2(n4863), .C1(n6003), 
        .C2(n5852), .ZN(U2837) );
  AOI22_X1 U5993 ( .A1(n6363), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6379), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n4864) );
  OAI21_X1 U5994 ( .B1(n6178), .B2(n6355), .A(n4864), .ZN(n4865) );
  AOI21_X1 U5995 ( .B1(n6180), .B2(n6360), .A(n4865), .ZN(n4866) );
  OAI21_X1 U5996 ( .B1(n6323), .B2(n4867), .A(n4866), .ZN(U2978) );
  AOI21_X1 U5997 ( .B1(n4870), .B2(n4869), .A(n4868), .ZN(n6326) );
  INV_X1 U5998 ( .A(n6326), .ZN(n4874) );
  INV_X1 U5999 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4872) );
  OAI222_X1 U6000 ( .A1(n4874), .A2(n5850), .B1(n5848), .B2(n4872), .C1(n5852), 
        .C2(n4871), .ZN(U2852) );
  OAI222_X1 U6001 ( .A1(n4874), .A2(n5862), .B1(n5796), .B2(n4873), .C1(n5109), 
        .C2(n3780), .ZN(U2884) );
  AND2_X1 U6002 ( .A1(n4979), .A2(n4875), .ZN(n4896) );
  AND2_X1 U6003 ( .A1(n4979), .A2(n4876), .ZN(n4932) );
  INV_X1 U6004 ( .A(n4932), .ZN(n4877) );
  OAI21_X1 U6005 ( .B1(n4896), .B2(n4878), .A(n4877), .ZN(n6129) );
  AOI22_X1 U6006 ( .A1(n6247), .A2(DATAI_16_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n6250), .ZN(n4880) );
  NAND2_X1 U6007 ( .A1(n6251), .A2(DATAI_0_), .ZN(n4879) );
  OAI211_X1 U6008 ( .C1(n6129), .C2(n5862), .A(n4880), .B(n4879), .ZN(U2875)
         );
  AND2_X1 U6009 ( .A1(n4979), .A2(n4881), .ZN(n4980) );
  AND2_X1 U6010 ( .A1(n4979), .A2(n4882), .ZN(n4910) );
  INV_X1 U6011 ( .A(n4910), .ZN(n4883) );
  OAI21_X1 U6012 ( .B1(n4884), .B2(n4980), .A(n4883), .ZN(n6014) );
  AOI22_X1 U6013 ( .A1(n6247), .A2(DATAI_20_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n6250), .ZN(n4886) );
  NAND2_X1 U6014 ( .A1(n6251), .A2(DATAI_4_), .ZN(n4885) );
  OAI211_X1 U6015 ( .C1(n6014), .C2(n5862), .A(n4886), .B(n4885), .ZN(U2871)
         );
  NAND2_X1 U6016 ( .A1(n4888), .A2(n4887), .ZN(n4891) );
  NAND2_X1 U6017 ( .A1(n4889), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4890)
         );
  INV_X1 U6018 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6392) );
  XNOR2_X1 U6019 ( .A(n6039), .B(n6392), .ZN(n4892) );
  XNOR2_X1 U6020 ( .A(n5241), .B(n4892), .ZN(n6390) );
  INV_X1 U6021 ( .A(n6323), .ZN(n6358) );
  NAND2_X1 U6022 ( .A1(n6390), .A2(n6358), .ZN(n4895) );
  INV_X1 U6023 ( .A(REIP_REG_9__SCAN_IN), .ZN(n5368) );
  OAI22_X1 U6024 ( .A1(n6339), .A2(n6163), .B1(n6426), .B2(n5368), .ZN(n4893)
         );
  AOI21_X1 U6025 ( .B1(n6332), .B2(n6170), .A(n4893), .ZN(n4894) );
  OAI211_X1 U6026 ( .C1(n5901), .C2(n6167), .A(n4895), .B(n4894), .ZN(U2977)
         );
  AOI21_X1 U6027 ( .B1(n4898), .B2(n4897), .A(n4896), .ZN(n6145) );
  INV_X1 U6028 ( .A(n6145), .ZN(n5073) );
  INV_X1 U6029 ( .A(n4916), .ZN(n4902) );
  AOI21_X1 U6030 ( .B1(n5102), .B2(n4900), .A(n4899), .ZN(n4901) );
  NOR2_X1 U6031 ( .A1(n4902), .A2(n4901), .ZN(n6139) );
  AOI22_X1 U6032 ( .A1(n6139), .A2(n5045), .B1(n5044), .B2(EBX_REG_15__SCAN_IN), .ZN(n4903) );
  OAI21_X1 U6033 ( .B1(n5073), .B2(n5850), .A(n4903), .ZN(U2844) );
  MUX2_X1 U6034 ( .A(n5659), .B(n4905), .S(n4904), .Z(n4907) );
  XNOR2_X1 U6035 ( .A(n4907), .B(n4906), .ZN(n6015) );
  OAI222_X1 U6036 ( .A1(n6014), .A2(n5850), .B1(n5852), .B2(n6015), .C1(n4908), 
        .C2(n5848), .ZN(U2839) );
  OR2_X1 U6037 ( .A1(n4910), .A2(n4909), .ZN(n4911) );
  INV_X1 U6038 ( .A(n6008), .ZN(n5071) );
  AOI22_X1 U6039 ( .A1(n6247), .A2(DATAI_21_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n6250), .ZN(n4914) );
  NAND2_X1 U6040 ( .A1(n6251), .A2(DATAI_5_), .ZN(n4913) );
  OAI211_X1 U6041 ( .C1(n5071), .C2(n5862), .A(n4914), .B(n4913), .ZN(U2870)
         );
  NAND2_X1 U6042 ( .A1(n4916), .A2(n4915), .ZN(n4917) );
  NAND2_X1 U6043 ( .A1(n4935), .A2(n4917), .ZN(n6128) );
  INV_X1 U6044 ( .A(EBX_REG_16__SCAN_IN), .ZN(n4918) );
  OAI222_X1 U6045 ( .A1(n6128), .A2(n5852), .B1(n5848), .B2(n4918), .C1(n5850), 
        .C2(n6129), .ZN(U2843) );
  AND2_X1 U6046 ( .A1(n4979), .A2(n4919), .ZN(n4921) );
  OR2_X1 U6047 ( .A1(n5106), .A2(n4922), .ZN(n4923) );
  NAND2_X1 U6048 ( .A1(n4924), .A2(n4923), .ZN(n5491) );
  INV_X1 U6049 ( .A(DATAI_13_), .ZN(n4925) );
  OAI222_X1 U6050 ( .A1(n5491), .A2(n5862), .B1(n5796), .B2(n4926), .C1(n4925), 
        .C2(n5109), .ZN(U2878) );
  OR2_X1 U6051 ( .A1(n5035), .A2(n4927), .ZN(n5037) );
  NAND2_X1 U6052 ( .A1(n5035), .A2(n4927), .ZN(n4928) );
  AOI22_X1 U6053 ( .A1(n5039), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n6250), .ZN(n4929) );
  OAI21_X1 U6054 ( .B1(n5372), .B2(n5862), .A(n4929), .ZN(U2881) );
  INV_X1 U6055 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6909) );
  NAND2_X1 U6056 ( .A1(n4979), .A2(n4930), .ZN(n5049) );
  OR2_X1 U6057 ( .A1(n4932), .A2(n4931), .ZN(n4933) );
  NAND2_X1 U6058 ( .A1(n6249), .A2(n5104), .ZN(n4938) );
  OR2_X1 U6059 ( .A1(n4935), .A2(n4934), .ZN(n5053) );
  NAND2_X1 U6060 ( .A1(n4935), .A2(n4934), .ZN(n4936) );
  AND2_X1 U6061 ( .A1(n5053), .A2(n4936), .ZN(n6124) );
  NAND2_X1 U6062 ( .A1(n6124), .A2(n5045), .ZN(n4937) );
  OAI211_X1 U6063 ( .C1(n6909), .C2(n5848), .A(n4938), .B(n4937), .ZN(U2842)
         );
  AOI22_X1 U6064 ( .A1(n4995), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4942) );
  AOI22_X1 U6065 ( .A1(n3510), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5680), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4941) );
  AOI22_X1 U6066 ( .A1(n5629), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n5619), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4940) );
  AOI22_X1 U6067 ( .A1(n4729), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n5682), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4939) );
  NAND4_X1 U6068 ( .A1(n4942), .A2(n4941), .A3(n4940), .A4(n4939), .ZN(n4948)
         );
  AOI22_X1 U6069 ( .A1(n5683), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3511), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4946) );
  AOI22_X1 U6070 ( .A1(n5620), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3607), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4945) );
  AOI22_X1 U6071 ( .A1(n4949), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4944) );
  AOI22_X1 U6072 ( .A1(n3608), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4943) );
  NAND4_X1 U6073 ( .A1(n4946), .A2(n4945), .A3(n4944), .A4(n4943), .ZN(n4947)
         );
  NOR2_X1 U6074 ( .A1(n4948), .A2(n4947), .ZN(n4989) );
  AOI22_X1 U6075 ( .A1(n3248), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5683), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4953) );
  AOI22_X1 U6076 ( .A1(n5691), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4952) );
  AOI22_X1 U6077 ( .A1(n5682), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4949), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4951) );
  AOI22_X1 U6078 ( .A1(n4729), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4950) );
  NAND4_X1 U6079 ( .A1(n4953), .A2(n4952), .A3(n4951), .A4(n4950), .ZN(n4959)
         );
  AOI22_X1 U6080 ( .A1(n5620), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n5629), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4957) );
  AOI22_X1 U6081 ( .A1(n5680), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5692), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4956) );
  AOI22_X1 U6082 ( .A1(n5688), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3607), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4955) );
  AOI22_X1 U6083 ( .A1(n3608), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4954) );
  NAND4_X1 U6084 ( .A1(n4957), .A2(n4956), .A3(n4955), .A4(n4954), .ZN(n4958)
         );
  NOR2_X1 U6085 ( .A1(n4959), .A2(n4958), .ZN(n4990) );
  XNOR2_X1 U6086 ( .A(n4989), .B(n4990), .ZN(n4962) );
  INV_X1 U6087 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4964) );
  OAI21_X1 U6088 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4964), .A(n5646), .ZN(
        n4960) );
  AOI21_X1 U6089 ( .B1(n5785), .B2(EAX_REG_23__SCAN_IN), .A(n4960), .ZN(n4961)
         );
  OAI21_X1 U6090 ( .B1(n4962), .B2(n5650), .A(n4961), .ZN(n4969) );
  AND2_X1 U6091 ( .A1(n4965), .A2(n4964), .ZN(n4966) );
  OR2_X1 U6092 ( .A1(n4966), .A2(n5091), .ZN(n5991) );
  INV_X1 U6093 ( .A(n5991), .ZN(n4967) );
  NAND2_X1 U6094 ( .A1(n4967), .A2(n5706), .ZN(n4968) );
  NAND2_X1 U6095 ( .A1(n4969), .A2(n4968), .ZN(n4975) );
  INV_X1 U6096 ( .A(n4975), .ZN(n4970) );
  INV_X1 U6097 ( .A(n5008), .ZN(n4973) );
  AOI21_X1 U6098 ( .B1(n4975), .B2(n4974), .A(n4973), .ZN(n5988) );
  INV_X1 U6099 ( .A(n5988), .ZN(n5022) );
  AOI22_X1 U6100 ( .A1(n6247), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6250), .ZN(n4977) );
  NAND2_X1 U6101 ( .A1(n6251), .A2(DATAI_7_), .ZN(n4976) );
  OAI211_X1 U6102 ( .C1(n5022), .C2(n5862), .A(n4977), .B(n4976), .ZN(U2868)
         );
  NAND2_X1 U6103 ( .A1(n4979), .A2(n4978), .ZN(n5047) );
  AOI21_X1 U6104 ( .B1(n4981), .B2(n5047), .A(n4980), .ZN(n6035) );
  INV_X1 U6105 ( .A(n5053), .ZN(n4984) );
  OR2_X1 U6106 ( .A1(n4983), .A2(n4982), .ZN(n5051) );
  NAND2_X1 U6107 ( .A1(n4984), .A2(n5051), .ZN(n5055) );
  XNOR2_X1 U6108 ( .A(n5055), .B(n4985), .ZN(n6030) );
  OAI22_X1 U6109 ( .A1(n6030), .A2(n5852), .B1(n4986), .B2(n5848), .ZN(n4987)
         );
  AOI21_X1 U6110 ( .B1(n6035), .B2(n5104), .A(n4987), .ZN(n4988) );
  INV_X1 U6111 ( .A(n4988), .ZN(U2840) );
  NOR2_X1 U6112 ( .A1(n4990), .A2(n4989), .ZN(n5075) );
  AOI22_X1 U6113 ( .A1(n5080), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n5629), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4994) );
  AOI22_X1 U6114 ( .A1(n5680), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5692), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4993) );
  AOI22_X1 U6115 ( .A1(n3510), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3607), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4992) );
  AOI22_X1 U6116 ( .A1(n3608), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4991) );
  NAND4_X1 U6117 ( .A1(n4994), .A2(n4993), .A3(n4992), .A4(n4991), .ZN(n5001)
         );
  AOI22_X1 U6118 ( .A1(n4995), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5683), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4999) );
  AOI22_X1 U6119 ( .A1(n3511), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4998) );
  AOI22_X1 U6120 ( .A1(n5682), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4997) );
  AOI22_X1 U6121 ( .A1(n4729), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4996) );
  NAND4_X1 U6122 ( .A1(n4999), .A2(n4998), .A3(n4997), .A4(n4996), .ZN(n5000)
         );
  OR2_X1 U6123 ( .A1(n5001), .A2(n5000), .ZN(n5074) );
  INV_X1 U6124 ( .A(n5074), .ZN(n5002) );
  XNOR2_X1 U6125 ( .A(n5075), .B(n5002), .ZN(n5007) );
  INV_X1 U6126 ( .A(n5650), .ZN(n5701) );
  INV_X1 U6127 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5976) );
  XNOR2_X1 U6128 ( .A(n5091), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5975)
         );
  NAND2_X1 U6129 ( .A1(n5975), .A2(n5706), .ZN(n5004) );
  NAND2_X1 U6130 ( .A1(n5785), .A2(EAX_REG_24__SCAN_IN), .ZN(n5003) );
  OAI211_X1 U6131 ( .C1(n5976), .C2(n5005), .A(n5004), .B(n5003), .ZN(n5006)
         );
  AOI21_X1 U6132 ( .B1(n5007), .B2(n5701), .A(n5006), .ZN(n5009) );
  NOR2_X2 U6133 ( .A1(n5008), .A2(n5009), .ZN(n5097) );
  AOI21_X1 U6134 ( .B1(n5009), .B2(n5008), .A(n5097), .ZN(n5974) );
  INV_X1 U6135 ( .A(n5974), .ZN(n5066) );
  AOI22_X1 U6136 ( .A1(n6247), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6250), .ZN(n5011) );
  NAND2_X1 U6137 ( .A1(n6251), .A2(DATAI_8_), .ZN(n5010) );
  OAI211_X1 U6138 ( .C1(n5066), .C2(n5862), .A(n5011), .B(n5010), .ZN(U2867)
         );
  INV_X1 U6139 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5019) );
  NAND2_X1 U6140 ( .A1(n5012), .A2(n5019), .ZN(n5015) );
  NAND2_X1 U6141 ( .A1(n5659), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5013) );
  OAI211_X1 U6142 ( .C1(n5773), .C2(EBX_REG_23__SCAN_IN), .A(n3112), .B(n5013), 
        .ZN(n5014) );
  AND2_X1 U6143 ( .A1(n5015), .A2(n5014), .ZN(n5016) );
  NOR2_X1 U6144 ( .A1(n5017), .A2(n5016), .ZN(n5018) );
  OR2_X1 U6145 ( .A1(n5063), .A2(n5018), .ZN(n5984) );
  OAI22_X1 U6146 ( .A1(n5984), .A2(n5852), .B1(n5019), .B2(n5848), .ZN(n5020)
         );
  INV_X1 U6147 ( .A(n5020), .ZN(n5021) );
  OAI21_X1 U6148 ( .B1(n5022), .B2(n5850), .A(n5021), .ZN(U2836) );
  OR2_X1 U6149 ( .A1(n5024), .A2(n5023), .ZN(n5025) );
  NAND2_X1 U6150 ( .A1(n5042), .A2(n5025), .ZN(n6381) );
  INV_X1 U6151 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6845) );
  OAI222_X1 U6152 ( .A1(n6381), .A2(n5852), .B1(n5848), .B2(n6845), .C1(n5850), 
        .C2(n5372), .ZN(U2849) );
  NOR2_X1 U6153 ( .A1(n5209), .A2(n6392), .ZN(n5192) );
  OR2_X1 U6154 ( .A1(n5241), .A2(n5192), .ZN(n5026) );
  NAND2_X1 U6155 ( .A1(n5209), .A2(n6392), .ZN(n5200) );
  NAND2_X1 U6156 ( .A1(n5026), .A2(n5200), .ZN(n5028) );
  INV_X1 U6157 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6385) );
  AND2_X1 U6158 ( .A1(n5209), .A2(n6385), .ZN(n5199) );
  NOR2_X1 U6159 ( .A1(n3115), .A2(n5199), .ZN(n5027) );
  XNOR2_X1 U6160 ( .A(n5028), .B(n5027), .ZN(n6383) );
  INV_X1 U6161 ( .A(n6383), .ZN(n5033) );
  AOI22_X1 U6162 ( .A1(n6363), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6379), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5029) );
  OAI21_X1 U6163 ( .B1(n5359), .B2(n6355), .A(n5029), .ZN(n5030) );
  AOI21_X1 U6164 ( .B1(n5031), .B2(n6360), .A(n5030), .ZN(n5032) );
  OAI21_X1 U6165 ( .B1(n5033), .B2(n6323), .A(n5032), .ZN(U2976) );
  OR2_X1 U6166 ( .A1(n5035), .A2(n5034), .ZN(n5107) );
  NAND2_X1 U6167 ( .A1(n5037), .A2(n5036), .ZN(n5038) );
  AOI22_X1 U6168 ( .A1(n5039), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n6250), .ZN(n5040) );
  OAI21_X1 U6169 ( .B1(n5358), .B2(n5862), .A(n5040), .ZN(U2880) );
  NAND2_X1 U6170 ( .A1(n5042), .A2(n5041), .ZN(n5043) );
  AND2_X1 U6171 ( .A1(n5316), .A2(n5043), .ZN(n6368) );
  AOI22_X1 U6172 ( .A1(n6368), .A2(n5045), .B1(n5044), .B2(EBX_REG_11__SCAN_IN), .ZN(n5046) );
  OAI21_X1 U6173 ( .B1(n5358), .B2(n5850), .A(n5046), .ZN(U2848) );
  INV_X1 U6174 ( .A(n5047), .ZN(n5048) );
  AOI21_X1 U6175 ( .B1(n5050), .B2(n5049), .A(n5048), .ZN(n6244) );
  INV_X1 U6176 ( .A(n6244), .ZN(n5057) );
  INV_X1 U6177 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5056) );
  INV_X1 U6178 ( .A(n5051), .ZN(n5052) );
  NAND2_X1 U6179 ( .A1(n5053), .A2(n5052), .ZN(n5054) );
  NAND2_X1 U6180 ( .A1(n5055), .A2(n5054), .ZN(n6118) );
  OAI222_X1 U6181 ( .A1(n5850), .A2(n5057), .B1(n5848), .B2(n5056), .C1(n6118), 
        .C2(n5852), .ZN(U2841) );
  INV_X1 U6182 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5065) );
  MUX2_X1 U6183 ( .A(n5662), .B(n3112), .S(EBX_REG_24__SCAN_IN), .Z(n5061) );
  NAND2_X1 U6184 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n5773), .ZN(n5058) );
  AND2_X1 U6185 ( .A1(n5059), .A2(n5058), .ZN(n5060) );
  NAND2_X1 U6186 ( .A1(n5061), .A2(n5060), .ZN(n5062) );
  OR2_X1 U6187 ( .A1(n5063), .A2(n5062), .ZN(n5064) );
  NAND2_X1 U6188 ( .A1(n5162), .A2(n5064), .ZN(n5983) );
  OAI222_X1 U6189 ( .A1(n5850), .A2(n5066), .B1(n5848), .B2(n5065), .C1(n5983), 
        .C2(n5852), .ZN(U2835) );
  NAND2_X1 U6190 ( .A1(n5068), .A2(n5067), .ZN(n5069) );
  NAND2_X1 U6191 ( .A1(n5070), .A2(n5069), .ZN(n6006) );
  INV_X1 U6192 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5072) );
  OAI222_X1 U6193 ( .A1(n5852), .A2(n6006), .B1(n5848), .B2(n5072), .C1(n5850), 
        .C2(n5071), .ZN(U2838) );
  OAI222_X1 U6194 ( .A1(n5109), .A2(n6766), .B1(n5796), .B2(n3318), .C1(n5862), 
        .C2(n5073), .ZN(U2876) );
  NAND2_X1 U6195 ( .A1(n5075), .A2(n5074), .ZN(n5251) );
  AOI22_X1 U6196 ( .A1(n5680), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5692), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n5079) );
  AOI22_X1 U6197 ( .A1(n5688), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3607), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5078) );
  AOI22_X1 U6198 ( .A1(n5689), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5077) );
  AOI22_X1 U6199 ( .A1(n3241), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5076) );
  NAND4_X1 U6200 ( .A1(n5079), .A2(n5078), .A3(n5077), .A4(n5076), .ZN(n5086)
         );
  AOI22_X1 U6201 ( .A1(n4995), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5683), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n5084) );
  AOI22_X1 U6202 ( .A1(n5080), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n5629), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5083) );
  AOI22_X1 U6203 ( .A1(n3511), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5682), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5082) );
  AOI22_X1 U6204 ( .A1(n3270), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n5081) );
  NAND4_X1 U6205 ( .A1(n5084), .A2(n5083), .A3(n5082), .A4(n5081), .ZN(n5085)
         );
  NOR2_X1 U6206 ( .A1(n5086), .A2(n5085), .ZN(n5252) );
  XNOR2_X1 U6207 ( .A(n5251), .B(n5252), .ZN(n5090) );
  NAND2_X1 U6208 ( .A1(n6814), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5087)
         );
  NAND2_X1 U6209 ( .A1(n5703), .A2(n5087), .ZN(n5088) );
  AOI21_X1 U6210 ( .B1(n5785), .B2(EAX_REG_25__SCAN_IN), .A(n5088), .ZN(n5089)
         );
  OAI21_X1 U6211 ( .B1(n5090), .B2(n5650), .A(n5089), .ZN(n5095) );
  OR2_X1 U6212 ( .A1(n5092), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5093)
         );
  NAND2_X1 U6213 ( .A1(n5267), .A2(n5093), .ZN(n5519) );
  OAI21_X1 U6214 ( .B1(n5097), .B2(n5096), .A(n5271), .ZN(n5517) );
  AOI22_X1 U6215 ( .A1(n6247), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6250), .ZN(n5099) );
  NAND2_X1 U6216 ( .A1(n6251), .A2(DATAI_9_), .ZN(n5098) );
  OAI211_X1 U6217 ( .C1(n5517), .C2(n5862), .A(n5099), .B(n5098), .ZN(U2866)
         );
  INV_X1 U6218 ( .A(n5491), .ZN(n6153) );
  NOR2_X1 U6219 ( .A1(n5317), .A2(n5100), .ZN(n5101) );
  OR2_X1 U6220 ( .A1(n5102), .A2(n5101), .ZN(n6149) );
  OAI22_X1 U6221 ( .A1(n6149), .A2(n5852), .B1(n6150), .B2(n5848), .ZN(n5103)
         );
  AOI21_X1 U6222 ( .B1(n6153), .B2(n5104), .A(n5103), .ZN(n5105) );
  INV_X1 U6223 ( .A(n5105), .ZN(U2846) );
  AOI21_X1 U6224 ( .B1(n5108), .B2(n5107), .A(n5106), .ZN(n5248) );
  INV_X1 U6225 ( .A(n5248), .ZN(n5351) );
  INV_X1 U6226 ( .A(DATAI_12_), .ZN(n6293) );
  OAI222_X1 U6227 ( .A1(n5351), .A2(n5862), .B1(n5796), .B2(n5110), .C1(n6293), 
        .C2(n5109), .ZN(U2879) );
  NAND2_X1 U6228 ( .A1(n6927), .A2(n6446), .ZN(n5159) );
  AND2_X1 U6229 ( .A1(n5946), .A2(n5111), .ZN(n5276) );
  NAND2_X1 U6230 ( .A1(n5112), .A2(n5276), .ZN(n6484) );
  AOI21_X1 U6231 ( .B1(n5113), .B2(n6484), .A(n6091), .ZN(n5116) );
  NOR2_X1 U6232 ( .A1(n5115), .A2(n5114), .ZN(n6442) );
  NOR2_X1 U6233 ( .A1(n5116), .A2(n6442), .ZN(n5117) );
  AOI22_X1 U6234 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5159), .B1(n5118), .B2(
        n5117), .ZN(n5120) );
  NAND3_X1 U6235 ( .A1(n6674), .A2(n5120), .A3(n5119), .ZN(n5152) );
  NAND2_X1 U6236 ( .A1(n5152), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5126) );
  NOR2_X1 U6237 ( .A1(n5121), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5122)
         );
  AOI22_X1 U6238 ( .A1(n5123), .A2(n6671), .B1(n5282), .B2(n5122), .ZN(n5153)
         );
  OAI22_X1 U6239 ( .A1(n6484), .A2(n6526), .B1(n5153), .B2(n5308), .ZN(n5124)
         );
  AOI21_X1 U6240 ( .B1(n5155), .B2(n6521), .A(n5124), .ZN(n5125) );
  OAI211_X1 U6241 ( .C1(n5159), .C2(n5127), .A(n5126), .B(n5125), .ZN(U3072)
         );
  NAND2_X1 U6242 ( .A1(n5152), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5130) );
  OAI22_X1 U6243 ( .A1(n6484), .A2(n6514), .B1(n5153), .B2(n5314), .ZN(n5128)
         );
  AOI21_X1 U6244 ( .B1(n5155), .B2(n6509), .A(n5128), .ZN(n5129) );
  OAI211_X1 U6245 ( .C1(n5159), .C2(n5131), .A(n5130), .B(n5129), .ZN(U3070)
         );
  NAND2_X1 U6246 ( .A1(n5152), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5134) );
  OAI22_X1 U6247 ( .A1(n6484), .A2(n6452), .B1(n5153), .B2(n5292), .ZN(n5132)
         );
  AOI21_X1 U6248 ( .B1(n6440), .B2(n5155), .A(n5132), .ZN(n5133) );
  OAI211_X1 U6249 ( .C1(n5135), .C2(n5159), .A(n5134), .B(n5133), .ZN(U3068)
         );
  NAND2_X1 U6250 ( .A1(n5152), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5138) );
  OAI22_X1 U6251 ( .A1(n6484), .A2(n6520), .B1(n5153), .B2(n5304), .ZN(n5136)
         );
  AOI21_X1 U6252 ( .B1(n5155), .B2(n6515), .A(n5136), .ZN(n5137) );
  OAI211_X1 U6253 ( .C1(n5159), .C2(n5139), .A(n5138), .B(n5137), .ZN(U3071)
         );
  NAND2_X1 U6254 ( .A1(n5152), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5142) );
  OAI22_X1 U6255 ( .A1(n6484), .A2(n6551), .B1(n5153), .B2(n5300), .ZN(n5140)
         );
  AOI21_X1 U6256 ( .B1(n5155), .B2(n6541), .A(n5140), .ZN(n5141) );
  OAI211_X1 U6257 ( .C1(n5159), .C2(n5143), .A(n5142), .B(n5141), .ZN(U3075)
         );
  NAND2_X1 U6258 ( .A1(n5152), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5146) );
  OAI22_X1 U6259 ( .A1(n6484), .A2(n6476), .B1(n5153), .B2(n5329), .ZN(n5144)
         );
  AOI21_X1 U6260 ( .B1(n5155), .B2(n6471), .A(n5144), .ZN(n5145) );
  OAI211_X1 U6261 ( .C1(n5159), .C2(n5147), .A(n5146), .B(n5145), .ZN(U3074)
         );
  NAND2_X1 U6262 ( .A1(n5152), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5150) );
  OAI22_X1 U6263 ( .A1(n6484), .A2(n6532), .B1(n5153), .B2(n5322), .ZN(n5148)
         );
  AOI21_X1 U6264 ( .B1(n5155), .B2(n6527), .A(n5148), .ZN(n5149) );
  OAI211_X1 U6265 ( .C1(n5159), .C2(n5151), .A(n5150), .B(n5149), .ZN(U3073)
         );
  NAND2_X1 U6266 ( .A1(n5152), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5157) );
  OAI22_X1 U6267 ( .A1(n6484), .A2(n6456), .B1(n5153), .B2(n5296), .ZN(n5154)
         );
  AOI21_X1 U6268 ( .B1(n5155), .B2(n6453), .A(n5154), .ZN(n5156) );
  OAI211_X1 U6269 ( .C1(n5159), .C2(n5158), .A(n5157), .B(n5156), .ZN(U3069)
         );
  INV_X1 U6270 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5165) );
  INV_X1 U6271 ( .A(n5162), .ZN(n5164) );
  MUX2_X1 U6272 ( .A(n5569), .B(n5659), .S(EBX_REG_25__SCAN_IN), .Z(n5160) );
  OAI21_X1 U6273 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5774), .A(n5160), 
        .ZN(n5161) );
  INV_X1 U6274 ( .A(n5161), .ZN(n5163) );
  OAI21_X1 U6275 ( .B1(n5164), .B2(n5163), .A(n5463), .ZN(n5532) );
  OAI222_X1 U6276 ( .A1(n5517), .A2(n5850), .B1(n5848), .B2(n5165), .C1(n5532), 
        .C2(n5852), .ZN(U2834) );
  NOR3_X1 U6277 ( .A1(n6580), .A2(n6826), .A3(n6582), .ZN(n6578) );
  NOR3_X1 U6278 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5806), .A3(n5646), .ZN(
        n6589) );
  INV_X1 U6279 ( .A(n6589), .ZN(n5166) );
  NAND2_X1 U6280 ( .A1(n6426), .A2(n5166), .ZN(n5167) );
  OR2_X1 U6281 ( .A1(n6578), .A2(n5167), .ZN(n5168) );
  INV_X1 U6282 ( .A(n5169), .ZN(n5170) );
  OR2_X1 U6283 ( .A1(n5817), .A2(n5170), .ZN(n5173) );
  INV_X1 U6284 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5885) );
  INV_X1 U6285 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6910) );
  INV_X1 U6286 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5870) );
  NOR2_X2 U6287 ( .A1(n5647), .A2(n5870), .ZN(n5612) );
  INV_X1 U6288 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6842) );
  INV_X1 U6289 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U6290 ( .A1(n5188), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U6291 ( .A1(n5173), .A2(n6199), .ZN(n6240) );
  INV_X1 U6292 ( .A(n6240), .ZN(n6222) );
  NOR2_X1 U6293 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5183) );
  NAND3_X1 U6294 ( .A1(n5174), .A2(n5183), .A3(n5185), .ZN(n5175) );
  INV_X1 U6295 ( .A(n6234), .ZN(n6191) );
  NAND2_X1 U6296 ( .A1(n6209), .A2(n6191), .ZN(n6110) );
  NOR2_X1 U6297 ( .A1(n5817), .A2(n5176), .ZN(n6232) );
  INV_X1 U6298 ( .A(n6232), .ZN(n5339) );
  INV_X1 U6299 ( .A(n5183), .ZN(n5181) );
  NAND3_X1 U6300 ( .A1(n5457), .A2(EBX_REG_31__SCAN_IN), .A3(n5181), .ZN(n5177) );
  OAI22_X1 U6301 ( .A1(n5339), .A2(n5179), .B1(n6243), .B2(n5178), .ZN(n5180)
         );
  AOI21_X1 U6302 ( .B1(REIP_REG_0__SCAN_IN), .B2(n6110), .A(n5180), .ZN(n5191)
         );
  OR2_X1 U6303 ( .A1(n6601), .A2(n5181), .ZN(n6577) );
  AND2_X1 U6304 ( .A1(n5182), .A2(n6577), .ZN(n5815) );
  NOR2_X1 U6305 ( .A1(n5183), .A2(EBX_REG_31__SCAN_IN), .ZN(n5184) );
  AND2_X1 U6306 ( .A1(n5185), .A2(n5184), .ZN(n5186) );
  NOR2_X1 U6307 ( .A1(n5815), .A2(n5186), .ZN(n5187) );
  INV_X1 U6308 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n6926) );
  AOI21_X1 U6309 ( .B1(n6220), .B2(n6238), .A(n6926), .ZN(n5189) );
  AOI21_X1 U6310 ( .B1(n6231), .B2(EBX_REG_0__SCAN_IN), .A(n5189), .ZN(n5190)
         );
  OAI211_X1 U6311 ( .C1(n6222), .C2(n6356), .A(n5191), .B(n5190), .ZN(U2827)
         );
  INV_X1 U6312 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6058) );
  NOR2_X1 U6313 ( .A1(n5209), .A2(n6058), .ZN(n5435) );
  INV_X1 U6314 ( .A(n5435), .ZN(n5193) );
  INV_X1 U6315 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6861) );
  OR2_X1 U6316 ( .A1(n5209), .A2(n6861), .ZN(n6315) );
  NAND2_X1 U6317 ( .A1(n5193), .A2(n6315), .ZN(n5194) );
  NAND2_X1 U6318 ( .A1(n5209), .A2(n6058), .ZN(n5484) );
  INV_X1 U6319 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U6320 ( .A1(n5209), .A2(n6076), .ZN(n5538) );
  INV_X1 U6321 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6865) );
  NAND2_X1 U6322 ( .A1(n5209), .A2(n6865), .ZN(n5196) );
  INV_X1 U6323 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6930) );
  NAND2_X1 U6324 ( .A1(n5209), .A2(n5448), .ZN(n5440) );
  AND2_X1 U6325 ( .A1(n3113), .A2(n5440), .ZN(n5197) );
  AND2_X1 U6326 ( .A1(n5494), .A2(n5197), .ZN(n5198) );
  AND2_X1 U6327 ( .A1(n5484), .A2(n5198), .ZN(n5203) );
  NAND2_X1 U6328 ( .A1(n5209), .A2(n6861), .ZN(n6314) );
  INV_X1 U6329 ( .A(n5199), .ZN(n5201) );
  AND2_X1 U6330 ( .A1(n6314), .A2(n5242), .ZN(n5202) );
  AND2_X1 U6331 ( .A1(n5203), .A2(n5202), .ZN(n5204) );
  NAND2_X1 U6332 ( .A1(n5205), .A2(n5204), .ZN(n5597) );
  INV_X1 U6333 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U6334 ( .A1(n5448), .A2(n6051), .ZN(n5598) );
  NOR2_X1 U6335 ( .A1(n5598), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5207)
         );
  OR2_X1 U6336 ( .A1(n6039), .A2(n5207), .ZN(n5212) );
  INV_X1 U6337 ( .A(n5437), .ZN(n5211) );
  XNOR2_X1 U6338 ( .A(n5209), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5486)
         );
  OR2_X1 U6339 ( .A1(n5209), .A2(n6865), .ZN(n5208) );
  OR2_X1 U6340 ( .A1(n5209), .A2(n6930), .ZN(n5496) );
  AND2_X1 U6341 ( .A1(n5492), .A2(n5496), .ZN(n5210) );
  NAND2_X1 U6342 ( .A1(n5597), .A2(n5213), .ZN(n5215) );
  NAND2_X1 U6343 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U6344 ( .A1(n6039), .A2(n5523), .ZN(n5214) );
  NAND2_X1 U6345 ( .A1(n5215), .A2(n5214), .ZN(n5515) );
  AND2_X1 U6346 ( .A1(n6039), .A2(n5431), .ZN(n5420) );
  INV_X1 U6347 ( .A(n5420), .ZN(n5216) );
  OR2_X1 U6348 ( .A1(n6039), .A2(n5431), .ZN(n5421) );
  NAND2_X1 U6349 ( .A1(n5216), .A2(n5421), .ZN(n5217) );
  XNOR2_X1 U6350 ( .A(n5515), .B(n5217), .ZN(n5239) );
  NAND3_X1 U6351 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n6070) );
  NOR2_X1 U6352 ( .A1(n6865), .A2(n6070), .ZN(n5446) );
  INV_X1 U6353 ( .A(n5446), .ZN(n5225) );
  INV_X1 U6354 ( .A(n6375), .ZN(n6377) );
  NAND4_X1 U6355 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n5218), .A4(n6377), .ZN(n5227)
         );
  NOR2_X1 U6356 ( .A1(n5219), .A2(n5227), .ZN(n5224) );
  NAND2_X1 U6357 ( .A1(n5222), .A2(n5224), .ZN(n6064) );
  OAI21_X1 U6358 ( .B1(n5227), .B2(n5220), .A(n6064), .ZN(n6055) );
  NAND2_X1 U6359 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5450) );
  INV_X1 U6360 ( .A(n5450), .ZN(n5221) );
  INV_X1 U6361 ( .A(n5523), .ZN(n5231) );
  NOR2_X1 U6362 ( .A1(n6415), .A2(n5222), .ZN(n5529) );
  OAI21_X1 U6363 ( .B1(n5224), .B2(n6416), .A(n5223), .ZN(n5409) );
  NOR2_X1 U6364 ( .A1(n5225), .A2(n5450), .ZN(n5228) );
  NOR2_X1 U6365 ( .A1(n5227), .A2(n5226), .ZN(n5408) );
  AOI222_X1 U6366 ( .A1(n5229), .A2(n5228), .B1(n5229), .B2(n6416), .C1(n5228), 
        .C2(n5408), .ZN(n5230) );
  NOR2_X1 U6367 ( .A1(n5409), .A2(n5230), .ZN(n6048) );
  OAI21_X1 U6368 ( .B1(n5231), .B2(n5529), .A(n6048), .ZN(n5608) );
  NAND2_X1 U6369 ( .A1(n5608), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5232) );
  NAND2_X1 U6370 ( .A1(n6379), .A2(REIP_REG_19__SCAN_IN), .ZN(n5236) );
  OAI211_X1 U6371 ( .C1(n6030), .C2(n6428), .A(n5232), .B(n5236), .ZN(n5233)
         );
  AOI21_X1 U6372 ( .B1(n5929), .B2(n5431), .A(n5233), .ZN(n5234) );
  OAI21_X1 U6373 ( .B1(n5239), .B2(n6406), .A(n5234), .ZN(U2999) );
  NAND2_X1 U6374 ( .A1(n6363), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5235)
         );
  OAI211_X1 U6375 ( .C1(n6355), .C2(n6026), .A(n5236), .B(n5235), .ZN(n5237)
         );
  AOI21_X1 U6376 ( .B1(n6035), .B2(n6360), .A(n5237), .ZN(n5238) );
  OAI21_X1 U6377 ( .B1(n5239), .B2(n6323), .A(n5238), .ZN(U2967) );
  NAND2_X1 U6378 ( .A1(n6317), .A2(n6314), .ZN(n5244) );
  NAND2_X1 U6379 ( .A1(n5244), .A2(n6315), .ZN(n5436) );
  INV_X1 U6380 ( .A(n5484), .ZN(n5245) );
  NOR2_X1 U6381 ( .A1(n5435), .A2(n5245), .ZN(n5246) );
  XNOR2_X1 U6382 ( .A(n5436), .B(n5246), .ZN(n5407) );
  NOR2_X1 U6383 ( .A1(n6426), .A2(n6878), .ZN(n5414) );
  NOR2_X1 U6384 ( .A1(n6339), .A2(n6858), .ZN(n5247) );
  AOI211_X1 U6385 ( .C1(n6332), .C2(n5348), .A(n5414), .B(n5247), .ZN(n5250)
         );
  NAND2_X1 U6386 ( .A1(n5248), .A2(n6360), .ZN(n5249) );
  OAI211_X1 U6387 ( .C1(n5407), .C2(n6323), .A(n5250), .B(n5249), .ZN(U2974)
         );
  INV_X1 U6388 ( .A(n5271), .ZN(n5273) );
  NOR2_X1 U6389 ( .A1(n5252), .A2(n5251), .ZN(n5398) );
  AOI22_X1 U6390 ( .A1(n5620), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n5679), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5256) );
  AOI22_X1 U6391 ( .A1(n5680), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5692), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n5255) );
  AOI22_X1 U6392 ( .A1(n5688), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3607), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5254) );
  AOI22_X1 U6393 ( .A1(n3270), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n5253) );
  NAND4_X1 U6394 ( .A1(n5256), .A2(n5255), .A3(n5254), .A4(n5253), .ZN(n5262)
         );
  AOI22_X1 U6395 ( .A1(n4995), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5683), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n5260) );
  AOI22_X1 U6396 ( .A1(n5691), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n5259) );
  AOI22_X1 U6397 ( .A1(n5682), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5258) );
  AOI22_X1 U6398 ( .A1(n3241), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5257) );
  NAND4_X1 U6399 ( .A1(n5260), .A2(n5259), .A3(n5258), .A4(n5257), .ZN(n5261)
         );
  OR2_X1 U6400 ( .A1(n5262), .A2(n5261), .ZN(n5397) );
  XNOR2_X1 U6401 ( .A(n5398), .B(n5397), .ZN(n5266) );
  NAND2_X1 U6402 ( .A1(n6814), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5263)
         );
  NAND2_X1 U6403 ( .A1(n5703), .A2(n5263), .ZN(n5264) );
  AOI21_X1 U6404 ( .B1(n5785), .B2(EAX_REG_26__SCAN_IN), .A(n5264), .ZN(n5265)
         );
  OAI21_X1 U6405 ( .B1(n5266), .B2(n5650), .A(n5265), .ZN(n5269) );
  XNOR2_X1 U6406 ( .A(n5267), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5962)
         );
  NAND2_X1 U6407 ( .A1(n5962), .A2(n5706), .ZN(n5268) );
  NAND2_X1 U6408 ( .A1(n5269), .A2(n5268), .ZN(n5270) );
  INV_X1 U6409 ( .A(n5270), .ZN(n5272) );
  OAI21_X1 U6410 ( .B1(n5273), .B2(n5272), .A(n5403), .ZN(n5967) );
  AOI22_X1 U6411 ( .A1(n6247), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6250), .ZN(n5275) );
  NAND2_X1 U6412 ( .A1(n6251), .A2(DATAI_10_), .ZN(n5274) );
  OAI211_X1 U6413 ( .C1(n5967), .C2(n5862), .A(n5275), .B(n5274), .ZN(U2865)
         );
  NAND2_X1 U6414 ( .A1(n6490), .A2(n5276), .ZN(n6539) );
  OAI21_X1 U6415 ( .B1(n5283), .B2(n6542), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5277) );
  INV_X1 U6416 ( .A(n5278), .ZN(n5279) );
  AND2_X1 U6417 ( .A1(n5279), .A2(n5469), .ZN(n6491) );
  NOR2_X1 U6418 ( .A1(n5280), .A2(n6674), .ZN(n5281) );
  AOI22_X1 U6419 ( .A1(n5286), .A2(n6491), .B1(n5282), .B2(n5281), .ZN(n5330)
         );
  NAND3_X1 U6420 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6560), .ZN(n6496) );
  NOR2_X1 U6421 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6496), .ZN(n5327)
         );
  INV_X1 U6422 ( .A(n6491), .ZN(n5285) );
  INV_X1 U6423 ( .A(n5327), .ZN(n5284) );
  AOI22_X1 U6424 ( .A1(n5286), .A2(n5285), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5284), .ZN(n5287) );
  OAI211_X1 U6425 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6814), .A(n5288), .B(n5287), .ZN(n5323) );
  AOI22_X1 U6426 ( .A1(n6542), .A2(n6487), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5323), .ZN(n5289) );
  OAI21_X1 U6427 ( .B1(n5325), .B2(n6502), .A(n5289), .ZN(n5290) );
  AOI21_X1 U6428 ( .B1(n6488), .B2(n5327), .A(n5290), .ZN(n5291) );
  OAI21_X1 U6429 ( .B1(n5330), .B2(n5292), .A(n5291), .ZN(U3100) );
  AOI22_X1 U6430 ( .A1(n6542), .A2(n6503), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5323), .ZN(n5293) );
  OAI21_X1 U6431 ( .B1(n5325), .B2(n6508), .A(n5293), .ZN(n5294) );
  AOI21_X1 U6432 ( .B1(n6504), .B2(n5327), .A(n5294), .ZN(n5295) );
  OAI21_X1 U6433 ( .B1(n5330), .B2(n5296), .A(n5295), .ZN(U3101) );
  AOI22_X1 U6434 ( .A1(n6542), .A2(n6478), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5323), .ZN(n5297) );
  OAI21_X1 U6435 ( .B1(n5325), .B2(n6485), .A(n5297), .ZN(n5298) );
  AOI21_X1 U6436 ( .B1(n6544), .B2(n5327), .A(n5298), .ZN(n5299) );
  OAI21_X1 U6437 ( .B1(n5330), .B2(n5300), .A(n5299), .ZN(U3107) );
  AOI22_X1 U6438 ( .A1(n6542), .A2(n6459), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5323), .ZN(n5301) );
  OAI21_X1 U6439 ( .B1(n5325), .B2(n6462), .A(n5301), .ZN(n5302) );
  AOI21_X1 U6440 ( .B1(n6516), .B2(n5327), .A(n5302), .ZN(n5303) );
  OAI21_X1 U6441 ( .B1(n5330), .B2(n5304), .A(n5303), .ZN(U3103) );
  AOI22_X1 U6442 ( .A1(n6542), .A2(n6463), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5323), .ZN(n5305) );
  OAI21_X1 U6443 ( .B1(n5325), .B2(n6466), .A(n5305), .ZN(n5306) );
  AOI21_X1 U6444 ( .B1(n6522), .B2(n5327), .A(n5306), .ZN(n5307) );
  OAI21_X1 U6445 ( .B1(n5330), .B2(n5308), .A(n5307), .ZN(U3104) );
  AOI22_X1 U6446 ( .A1(n6542), .A2(n5309), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5323), .ZN(n5310) );
  OAI21_X1 U6447 ( .B1(n5325), .B2(n5311), .A(n5310), .ZN(n5312) );
  AOI21_X1 U6448 ( .B1(n6510), .B2(n5327), .A(n5312), .ZN(n5313) );
  OAI21_X1 U6449 ( .B1(n5330), .B2(n5314), .A(n5313), .ZN(U3102) );
  AND2_X1 U6450 ( .A1(n5316), .A2(n5315), .ZN(n5318) );
  OR2_X1 U6451 ( .A1(n5318), .A2(n5317), .ZN(n5416) );
  INV_X1 U6452 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6856) );
  OAI222_X1 U6453 ( .A1(n5416), .A2(n5852), .B1(n5848), .B2(n6856), .C1(n5850), 
        .C2(n5351), .ZN(U2847) );
  AOI22_X1 U6454 ( .A1(n6542), .A2(n6467), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5323), .ZN(n5319) );
  OAI21_X1 U6455 ( .B1(n5325), .B2(n6470), .A(n5319), .ZN(n5320) );
  AOI21_X1 U6456 ( .B1(n6528), .B2(n5327), .A(n5320), .ZN(n5321) );
  OAI21_X1 U6457 ( .B1(n5330), .B2(n5322), .A(n5321), .ZN(U3105) );
  AOI22_X1 U6458 ( .A1(n6542), .A2(n6533), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5323), .ZN(n5324) );
  OAI21_X1 U6459 ( .B1(n5325), .B2(n6540), .A(n5324), .ZN(n5326) );
  AOI21_X1 U6460 ( .B1(n6535), .B2(n5327), .A(n5326), .ZN(n5328) );
  OAI21_X1 U6461 ( .B1(n5330), .B2(n5329), .A(n5328), .ZN(U3106) );
  INV_X1 U6462 ( .A(n5542), .ZN(n5336) );
  INV_X1 U6463 ( .A(n6243), .ZN(n6214) );
  AOI22_X1 U6464 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6231), .B1(n6214), .B2(n6057), .ZN(n5331) );
  NOR3_X2 U6465 ( .A1(n6492), .A2(STATE2_REG_1__SCAN_IN), .A3(n6234), .ZN(
        n6207) );
  INV_X1 U6466 ( .A(n6207), .ZN(n6218) );
  OAI211_X1 U6467 ( .C1(n6220), .C2(n6912), .A(n5331), .B(n6218), .ZN(n5335)
         );
  INV_X1 U6468 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6633) );
  INV_X1 U6469 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6628) );
  INV_X1 U6470 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6676) );
  INV_X1 U6471 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6614) );
  NOR3_X1 U6472 ( .A1(n6676), .A2(n5480), .A3(n6614), .ZN(n6215) );
  NAND2_X1 U6473 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6215), .ZN(n6208) );
  NOR2_X1 U6474 ( .A1(n6619), .A2(n6208), .ZN(n6192) );
  NAND2_X1 U6475 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6192), .ZN(n6185) );
  NOR2_X1 U6476 ( .A1(n4796), .A2(n6185), .ZN(n6173) );
  NAND2_X1 U6477 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6173), .ZN(n5366) );
  NOR2_X1 U6478 ( .A1(n5368), .A2(n5366), .ZN(n5360) );
  NAND2_X1 U6479 ( .A1(REIP_REG_10__SCAN_IN), .A2(n5360), .ZN(n5332) );
  NAND3_X1 U6480 ( .A1(n6156), .A2(REIP_REG_12__SCAN_IN), .A3(
        REIP_REG_13__SCAN_IN), .ZN(n6132) );
  INV_X1 U6481 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6878) );
  INV_X1 U6482 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6631) );
  NOR3_X1 U6483 ( .A1(n6633), .A2(n6878), .A3(n6631), .ZN(n5373) );
  NOR3_X1 U6484 ( .A1(n6234), .A2(n6628), .A3(n5332), .ZN(n5375) );
  INV_X1 U6485 ( .A(n6110), .ZN(n5567) );
  AOI21_X1 U6486 ( .B1(n5373), .B2(n5375), .A(n5567), .ZN(n6142) );
  INV_X1 U6487 ( .A(n6142), .ZN(n5333) );
  AOI21_X1 U6488 ( .B1(n6633), .B2(n6132), .A(n5333), .ZN(n5334) );
  AOI211_X1 U6489 ( .C1(n5994), .C2(n5336), .A(n5335), .B(n5334), .ZN(n5337)
         );
  OAI21_X1 U6490 ( .B1(n5546), .B2(n6199), .A(n5337), .ZN(U2813) );
  INV_X1 U6491 ( .A(n6209), .ZN(n6216) );
  NAND2_X1 U6492 ( .A1(n6216), .A2(n6676), .ZN(n6241) );
  INV_X1 U6493 ( .A(n6241), .ZN(n5338) );
  NOR3_X1 U6494 ( .A1(n5338), .A2(n6234), .A3(n6614), .ZN(n5345) );
  AOI21_X1 U6495 ( .B1(n6216), .B2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .ZN(n5344) );
  OAI22_X1 U6496 ( .A1(n3602), .A2(n6220), .B1(n6238), .B2(n6347), .ZN(n5341)
         );
  OAI22_X1 U6497 ( .A1(n5339), .A2(n5951), .B1(n6419), .B2(n6243), .ZN(n5340)
         );
  AOI211_X1 U6498 ( .C1(n6231), .C2(EBX_REG_2__SCAN_IN), .A(n5341), .B(n5340), 
        .ZN(n5343) );
  NAND2_X1 U6499 ( .A1(n6344), .A2(n6240), .ZN(n5342) );
  OAI211_X1 U6500 ( .C1(n5345), .C2(n5344), .A(n5343), .B(n5342), .ZN(U2825)
         );
  NOR2_X1 U6501 ( .A1(n5567), .A2(n5375), .ZN(n6155) );
  AND2_X1 U6502 ( .A1(n6878), .A2(n6156), .ZN(n6154) );
  AOI22_X1 U6503 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6231), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6235), .ZN(n5346) );
  OAI211_X1 U6504 ( .C1(n5416), .C2(n6243), .A(n5346), .B(n6218), .ZN(n5347)
         );
  AOI211_X1 U6505 ( .C1(n6155), .C2(REIP_REG_12__SCAN_IN), .A(n6154), .B(n5347), .ZN(n5350) );
  NAND2_X1 U6506 ( .A1(n5994), .A2(n5348), .ZN(n5349) );
  OAI211_X1 U6507 ( .C1(n5351), .C2(n6199), .A(n5350), .B(n5349), .ZN(U2815)
         );
  NAND2_X1 U6508 ( .A1(n6628), .A2(n5352), .ZN(n5356) );
  INV_X1 U6509 ( .A(EBX_REG_11__SCAN_IN), .ZN(n7004) );
  INV_X1 U6510 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6970) );
  OAI22_X1 U6511 ( .A1(n7004), .A2(n6175), .B1(n6970), .B2(n6220), .ZN(n5355)
         );
  NAND2_X1 U6512 ( .A1(n6214), .A2(n6368), .ZN(n5353) );
  OAI211_X1 U6513 ( .C1(n6318), .C2(n6238), .A(n5353), .B(n6218), .ZN(n5354)
         );
  AOI211_X1 U6514 ( .C1(n6155), .C2(n5356), .A(n5355), .B(n5354), .ZN(n5357)
         );
  OAI21_X1 U6515 ( .B1(n5358), .B2(n6199), .A(n5357), .ZN(U2816) );
  INV_X1 U6516 ( .A(n5359), .ZN(n5364) );
  INV_X1 U6517 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6626) );
  NAND3_X1 U6518 ( .A1(n6216), .A2(n6626), .A3(n5360), .ZN(n5361) );
  OAI211_X1 U6519 ( .C1(n6220), .C2(n6830), .A(n6218), .B(n5361), .ZN(n5363)
         );
  OAI22_X1 U6520 ( .A1(n6845), .A2(n6175), .B1(n6243), .B2(n6381), .ZN(n5362)
         );
  AOI211_X1 U6521 ( .C1(n5994), .C2(n5364), .A(n5363), .B(n5362), .ZN(n5371)
         );
  OR2_X1 U6522 ( .A1(n6234), .A2(n5366), .ZN(n5365) );
  NAND2_X1 U6523 ( .A1(n6110), .A2(n5365), .ZN(n6183) );
  INV_X1 U6524 ( .A(n6183), .ZN(n6169) );
  INV_X1 U6525 ( .A(n5366), .ZN(n5367) );
  NAND2_X1 U6526 ( .A1(n5368), .A2(n5367), .ZN(n5369) );
  NOR2_X1 U6527 ( .A1(n6209), .A2(n5369), .ZN(n6165) );
  OAI21_X1 U6528 ( .B1(n6169), .B2(n6165), .A(REIP_REG_10__SCAN_IN), .ZN(n5370) );
  OAI211_X1 U6529 ( .C1(n5372), .C2(n6199), .A(n5371), .B(n5370), .ZN(U2817)
         );
  INV_X1 U6530 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6896) );
  INV_X1 U6531 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6639) );
  INV_X1 U6532 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6917) );
  INV_X1 U6533 ( .A(n5373), .ZN(n5374) );
  NAND2_X1 U6534 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n6133) );
  NOR2_X1 U6535 ( .A1(n5374), .A2(n6133), .ZN(n5376) );
  NAND2_X1 U6536 ( .A1(n6156), .A2(n5376), .ZN(n6120) );
  NAND2_X1 U6537 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6111), .ZN(n6027) );
  NOR2_X1 U6538 ( .A1(n6639), .A2(n6027), .ZN(n6019) );
  NAND2_X1 U6539 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6019), .ZN(n5992) );
  NAND3_X1 U6540 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5378) );
  NOR2_X1 U6541 ( .A1(n5992), .A2(n5378), .ZN(n5673) );
  AND2_X1 U6542 ( .A1(n6896), .A2(n5673), .ZN(n5980) );
  INV_X1 U6543 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6113) );
  NAND3_X1 U6544 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5376), .A3(n5375), .ZN(
        n6109) );
  NOR3_X1 U6545 ( .A1(n6639), .A2(n6113), .A3(n6109), .ZN(n5377) );
  AOI21_X1 U6546 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5377), .A(n5567), .ZN(n6018) );
  AOI21_X1 U6547 ( .B1(n5378), .B2(n6110), .A(n6018), .ZN(n5986) );
  INV_X1 U6548 ( .A(n5986), .ZN(n5379) );
  OAI21_X1 U6549 ( .B1(n5980), .B2(n5379), .A(REIP_REG_25__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U6550 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5673), .ZN(n5964) );
  OAI22_X1 U6551 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5964), .B1(n5519), .B2(
        n6238), .ZN(n5382) );
  AOI22_X1 U6552 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6231), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6235), .ZN(n5380) );
  OAI21_X1 U6553 ( .B1(n5532), .B2(n6243), .A(n5380), .ZN(n5381) );
  NOR2_X1 U6554 ( .A1(n5382), .A2(n5381), .ZN(n5383) );
  OAI211_X1 U6555 ( .C1(n5517), .C2(n6199), .A(n5384), .B(n5383), .ZN(U2802)
         );
  NAND2_X1 U6556 ( .A1(n5385), .A2(n6910), .ZN(n5386) );
  NAND2_X1 U6557 ( .A1(n5647), .A2(n5386), .ZN(n5880) );
  AOI22_X1 U6558 ( .A1(n5634), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5390) );
  AOI22_X1 U6559 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n5629), .B1(n3241), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5389) );
  AOI22_X1 U6560 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n5680), .B1(n3607), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5388) );
  AOI22_X1 U6561 ( .A1(n3511), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n5682), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5387) );
  NAND4_X1 U6562 ( .A1(n5390), .A2(n5389), .A3(n5388), .A4(n5387), .ZN(n5396)
         );
  AOI22_X1 U6563 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3510), .B1(n5692), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n5394) );
  AOI22_X1 U6564 ( .A1(n3248), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5393) );
  AOI22_X1 U6565 ( .A1(n3270), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4709), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n5392) );
  AOI22_X1 U6566 ( .A1(n5620), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5391) );
  NAND4_X1 U6567 ( .A1(n5394), .A2(n5393), .A3(n5392), .A4(n5391), .ZN(n5395)
         );
  NOR2_X1 U6568 ( .A1(n5396), .A2(n5395), .ZN(n5628) );
  NAND2_X1 U6569 ( .A1(n5398), .A2(n5397), .ZN(n5627) );
  XNOR2_X1 U6570 ( .A(n5628), .B(n5627), .ZN(n5401) );
  OAI21_X1 U6571 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6910), .A(n5703), .ZN(
        n5399) );
  AOI21_X1 U6572 ( .B1(n5785), .B2(EAX_REG_27__SCAN_IN), .A(n5399), .ZN(n5400)
         );
  OAI21_X1 U6573 ( .B1(n5401), .B2(n5650), .A(n5400), .ZN(n5402) );
  OAI21_X1 U6574 ( .B1(n5646), .B2(n5880), .A(n5402), .ZN(n5404) );
  AOI21_X1 U6575 ( .B1(n5404), .B2(n5403), .A(n5830), .ZN(n5882) );
  INV_X1 U6576 ( .A(n5882), .ZN(n5851) );
  AOI22_X1 U6577 ( .A1(n6247), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6250), .ZN(n5406) );
  NAND2_X1 U6578 ( .A1(n6251), .A2(DATAI_11_), .ZN(n5405) );
  OAI211_X1 U6579 ( .C1(n5851), .C2(n5862), .A(n5406), .B(n5405), .ZN(U2864)
         );
  NOR2_X1 U6580 ( .A1(n5407), .A2(n6406), .ZN(n5419) );
  INV_X1 U6581 ( .A(n5408), .ZN(n5410) );
  AOI21_X1 U6582 ( .B1(n5411), .B2(n5410), .A(n5409), .ZN(n6371) );
  AOI211_X1 U6583 ( .C1(INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n6371), .A(n5412), .B(n6058), .ZN(n5418) );
  NOR3_X1 U6584 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6372), .A3(n6861), 
        .ZN(n5413) );
  NOR2_X1 U6585 ( .A1(n5414), .A2(n5413), .ZN(n5415) );
  OAI21_X1 U6586 ( .B1(n5416), .B2(n6428), .A(n5415), .ZN(n5417) );
  OR3_X1 U6587 ( .A1(n5419), .A2(n5418), .A3(n5417), .ZN(U3006) );
  NAND2_X1 U6588 ( .A1(n5422), .A2(n5421), .ZN(n5424) );
  XNOR2_X1 U6589 ( .A(n5209), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5423)
         );
  NAND2_X1 U6590 ( .A1(n5424), .A2(n5423), .ZN(n5892) );
  OAI21_X1 U6591 ( .B1(n5424), .B2(n5423), .A(n5892), .ZN(n5434) );
  NAND2_X1 U6592 ( .A1(n6379), .A2(REIP_REG_20__SCAN_IN), .ZN(n5429) );
  OAI21_X1 U6593 ( .B1(n6339), .B2(n5425), .A(n5429), .ZN(n5427) );
  NOR2_X1 U6594 ( .A1(n6014), .A2(n5901), .ZN(n5426) );
  AOI211_X1 U6595 ( .C1(n6332), .C2(n6020), .A(n5427), .B(n5426), .ZN(n5428)
         );
  OAI21_X1 U6596 ( .B1(n6323), .B2(n5434), .A(n5428), .ZN(U2966) );
  OAI21_X1 U6597 ( .B1(n6015), .B2(n6428), .A(n5429), .ZN(n5430) );
  AOI21_X1 U6598 ( .B1(n5608), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5430), 
        .ZN(n5433) );
  INV_X1 U6599 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U6600 ( .A1(n5556), .A2(n5431), .ZN(n5512) );
  AND2_X1 U6601 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5513) );
  INV_X1 U6602 ( .A(n5513), .ZN(n5935) );
  NAND3_X1 U6603 ( .A1(n5929), .A2(n5512), .A3(n5935), .ZN(n5432) );
  OAI211_X1 U6604 ( .C1(n5434), .C2(n6406), .A(n5433), .B(n5432), .ZN(U2998)
         );
  AND2_X1 U6605 ( .A1(n5484), .A2(n5437), .ZN(n5438) );
  NAND2_X1 U6606 ( .A1(n5485), .A2(n5438), .ZN(n5439) );
  NAND2_X1 U6607 ( .A1(n5439), .A2(n5596), .ZN(n5594) );
  NOR2_X1 U6608 ( .A1(n6039), .A2(n5448), .ZN(n6041) );
  INV_X1 U6609 ( .A(n5440), .ZN(n5441) );
  NOR2_X1 U6610 ( .A1(n6041), .A2(n5441), .ZN(n5442) );
  XNOR2_X1 U6611 ( .A(n5594), .B(n5442), .ZN(n5455) );
  NAND2_X1 U6612 ( .A1(n6379), .A2(REIP_REG_16__SCAN_IN), .ZN(n5452) );
  OAI21_X1 U6613 ( .B1(n6339), .B2(n6795), .A(n5452), .ZN(n5444) );
  NOR2_X1 U6614 ( .A1(n6129), .A2(n5901), .ZN(n5443) );
  AOI211_X1 U6615 ( .C1(n6332), .C2(n6131), .A(n5444), .B(n5443), .ZN(n5445)
         );
  OAI21_X1 U6616 ( .B1(n5455), .B2(n6323), .A(n5445), .ZN(U2970) );
  OAI21_X1 U6617 ( .B1(n5446), .B2(n6429), .A(n6371), .ZN(n5506) );
  INV_X1 U6618 ( .A(n5507), .ZN(n5447) );
  AOI21_X1 U6619 ( .B1(n6930), .B2(n5448), .A(n5447), .ZN(n5449) );
  NAND2_X1 U6620 ( .A1(n5450), .A2(n5449), .ZN(n5451) );
  OAI211_X1 U6621 ( .C1(n6128), .C2(n6428), .A(n5452), .B(n5451), .ZN(n5453)
         );
  AOI21_X1 U6622 ( .B1(n5506), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5453), 
        .ZN(n5454) );
  OAI21_X1 U6623 ( .B1(n5455), .B2(n6406), .A(n5454), .ZN(U3002) );
  INV_X1 U6624 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U6625 ( .A1(n5456), .A2(n5973), .ZN(n5461) );
  INV_X1 U6626 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6775) );
  NAND2_X1 U6627 ( .A1(n3112), .A2(n6775), .ZN(n5459) );
  NAND2_X1 U6628 ( .A1(n5457), .A2(n5973), .ZN(n5458) );
  NAND3_X1 U6629 ( .A1(n5459), .A2(n5659), .A3(n5458), .ZN(n5460) );
  AND2_X1 U6630 ( .A1(n5461), .A2(n5460), .ZN(n5462) );
  AND2_X1 U6631 ( .A1(n5463), .A2(n5462), .ZN(n5464) );
  OR2_X1 U6632 ( .A1(n5464), .A2(n5573), .ZN(n5966) );
  OAI22_X1 U6633 ( .A1(n5966), .A2(n5852), .B1(n5973), .B2(n5848), .ZN(n5465)
         );
  INV_X1 U6634 ( .A(n5465), .ZN(n5466) );
  OAI21_X1 U6635 ( .B1(n5967), .B2(n5850), .A(n5466), .ZN(U2833) );
  INV_X1 U6636 ( .A(REIP_REG_3__SCAN_IN), .ZN(n5480) );
  INV_X1 U6637 ( .A(n6215), .ZN(n5467) );
  OR2_X1 U6638 ( .A1(n6234), .A2(n5467), .ZN(n5468) );
  NAND2_X1 U6639 ( .A1(n6110), .A2(n5468), .ZN(n6229) );
  AOI22_X1 U6640 ( .A1(n6232), .A2(n5469), .B1(n6231), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n5479) );
  INV_X1 U6641 ( .A(n6404), .ZN(n5476) );
  OAI22_X1 U6642 ( .A1(n5471), .A2(n6220), .B1(n6238), .B2(n5470), .ZN(n5472)
         );
  INV_X1 U6643 ( .A(n5472), .ZN(n5475) );
  NOR3_X1 U6644 ( .A1(n6614), .A2(n6215), .A3(n6676), .ZN(n5473) );
  NAND2_X1 U6645 ( .A1(n6216), .A2(n5473), .ZN(n5474) );
  OAI211_X1 U6646 ( .C1(n5476), .C2(n6243), .A(n5475), .B(n5474), .ZN(n5477)
         );
  INV_X1 U6647 ( .A(n5477), .ZN(n5478) );
  OAI211_X1 U6648 ( .C1(n5480), .C2(n6229), .A(n5479), .B(n5478), .ZN(n5481)
         );
  AOI21_X1 U6649 ( .B1(n5482), .B2(n6240), .A(n5481), .ZN(n5483) );
  INV_X1 U6650 ( .A(n5483), .ZN(U2824) );
  NAND2_X1 U6651 ( .A1(n5485), .A2(n5484), .ZN(n5493) );
  NAND2_X1 U6652 ( .A1(n5493), .A2(n5486), .ZN(n5539) );
  OAI21_X1 U6653 ( .B1(n5493), .B2(n5486), .A(n5539), .ZN(n6074) );
  NAND2_X1 U6654 ( .A1(n6074), .A2(n6358), .ZN(n5490) );
  INV_X1 U6655 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5487) );
  OAI22_X1 U6656 ( .A1(n6339), .A2(n5487), .B1(n6426), .B2(n6631), .ZN(n5488)
         );
  AOI21_X1 U6657 ( .B1(n6332), .B2(n6152), .A(n5488), .ZN(n5489) );
  OAI211_X1 U6658 ( .C1(n5901), .C2(n5491), .A(n5490), .B(n5489), .ZN(U2973)
         );
  NAND2_X1 U6659 ( .A1(n5493), .A2(n5492), .ZN(n5495) );
  NAND2_X1 U6660 ( .A1(n5495), .A2(n5494), .ZN(n5498) );
  NAND2_X1 U6661 ( .A1(n3113), .A2(n5496), .ZN(n5497) );
  XNOR2_X1 U6662 ( .A(n5498), .B(n5497), .ZN(n5510) );
  INV_X1 U6663 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5499) );
  NOR2_X1 U6664 ( .A1(n6426), .A2(n5499), .ZN(n5505) );
  AOI21_X1 U6665 ( .B1(n6363), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5505), 
        .ZN(n5500) );
  OAI21_X1 U6666 ( .B1(n6143), .B2(n6355), .A(n5500), .ZN(n5501) );
  AOI21_X1 U6667 ( .B1(n6145), .B2(n6360), .A(n5501), .ZN(n5502) );
  OAI21_X1 U6668 ( .B1(n5510), .B2(n6323), .A(n5502), .ZN(U2971) );
  INV_X1 U6669 ( .A(n6139), .ZN(n5503) );
  NOR2_X1 U6670 ( .A1(n5503), .A2(n6428), .ZN(n5504) );
  AOI211_X1 U6671 ( .C1(n5506), .C2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5505), .B(n5504), .ZN(n5509) );
  NAND2_X1 U6672 ( .A1(n5507), .A2(n6930), .ZN(n5508) );
  OAI211_X1 U6673 ( .C1(n5510), .C2(n6406), .A(n5509), .B(n5508), .ZN(U3003)
         );
  OR4_X1 U6674 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .A3(INSTADDRPOINTER_REG_22__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5511) );
  OAI21_X1 U6675 ( .B1(n5512), .B2(n5511), .A(n5206), .ZN(n5514) );
  AND2_X1 U6676 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5525) );
  AND2_X1 U6677 ( .A1(n5513), .A2(n5525), .ZN(n5928) );
  AND2_X1 U6678 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5528) );
  NAND2_X1 U6679 ( .A1(n5928), .A2(n5528), .ZN(n5733) );
  AOI22_X2 U6680 ( .A1(n5515), .A2(n5514), .B1(n5209), .B2(n5733), .ZN(n5864)
         );
  XOR2_X1 U6681 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(n6039), .Z(n5516) );
  AOI21_X1 U6682 ( .B1(n5864), .B2(n5516), .A(n5548), .ZN(n5537) );
  INV_X1 U6683 ( .A(n5517), .ZN(n5521) );
  INV_X1 U6684 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5965) );
  OR2_X1 U6685 ( .A1(n6426), .A2(n5965), .ZN(n5531) );
  NAND2_X1 U6686 ( .A1(n6363), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5518)
         );
  OAI211_X1 U6687 ( .C1(n6355), .C2(n5519), .A(n5531), .B(n5518), .ZN(n5520)
         );
  AOI21_X1 U6688 ( .B1(n5521), .B2(n6360), .A(n5520), .ZN(n5522) );
  OAI21_X1 U6689 ( .B1(n5537), .B2(n6323), .A(n5522), .ZN(U2961) );
  OAI21_X1 U6690 ( .B1(n5935), .B2(n5523), .A(n6374), .ZN(n5524) );
  NAND2_X1 U6691 ( .A1(n6048), .A2(n5524), .ZN(n5940) );
  INV_X1 U6692 ( .A(n5525), .ZN(n5526) );
  AND2_X1 U6693 ( .A1(n6374), .A2(n5526), .ZN(n5527) );
  OR2_X1 U6694 ( .A1(n5940), .A2(n5527), .ZN(n5926) );
  NOR2_X1 U6695 ( .A1(n5529), .A2(n5528), .ZN(n5530) );
  NOR2_X1 U6696 ( .A1(n5926), .A2(n5530), .ZN(n5756) );
  INV_X1 U6697 ( .A(n5756), .ZN(n5554) );
  OAI21_X1 U6698 ( .B1(n5532), .B2(n6428), .A(n5531), .ZN(n5535) );
  INV_X1 U6699 ( .A(n5733), .ZN(n5533) );
  NAND2_X1 U6700 ( .A1(n5929), .A2(n5533), .ZN(n5551) );
  NOR2_X1 U6701 ( .A1(n5551), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5534)
         );
  AOI211_X1 U6702 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n5554), .A(n5535), .B(n5534), .ZN(n5536) );
  OAI21_X1 U6703 ( .B1(n5537), .B2(n6406), .A(n5536), .ZN(U2993) );
  NAND2_X1 U6704 ( .A1(n5539), .A2(n5538), .ZN(n5541) );
  XNOR2_X1 U6705 ( .A(n6039), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5540)
         );
  XNOR2_X1 U6706 ( .A(n5541), .B(n5540), .ZN(n6066) );
  NAND2_X1 U6707 ( .A1(n6066), .A2(n6358), .ZN(n5545) );
  NOR2_X1 U6708 ( .A1(n6426), .A2(n6633), .ZN(n6056) );
  NOR2_X1 U6709 ( .A1(n6355), .A2(n5542), .ZN(n5543) );
  AOI211_X1 U6710 ( .C1(n6363), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6056), 
        .B(n5543), .ZN(n5544) );
  OAI211_X1 U6711 ( .C1(n5901), .C2(n5546), .A(n5545), .B(n5544), .ZN(U2972)
         );
  INV_X1 U6712 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6974) );
  NOR2_X2 U6713 ( .A1(n5548), .A2(n5547), .ZN(n5863) );
  XNOR2_X1 U6714 ( .A(n6039), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5549)
         );
  XNOR2_X1 U6715 ( .A(n5863), .B(n5549), .ZN(n5889) );
  NAND2_X1 U6716 ( .A1(n6379), .A2(REIP_REG_26__SCAN_IN), .ZN(n5884) );
  OAI21_X1 U6717 ( .B1(n5966), .B2(n6428), .A(n5884), .ZN(n5553) );
  NAND2_X1 U6718 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5734) );
  INV_X1 U6719 ( .A(n5734), .ZN(n5550) );
  NOR2_X1 U6720 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5865) );
  NOR3_X1 U6721 ( .A1(n5551), .A2(n5550), .A3(n5865), .ZN(n5552) );
  AOI211_X1 U6722 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5554), .A(n5553), .B(n5552), .ZN(n5555) );
  OAI21_X1 U6723 ( .B1(n5889), .B2(n6406), .A(n5555), .ZN(U2992) );
  INV_X1 U6724 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5934) );
  XNOR2_X1 U6725 ( .A(n6039), .B(n5934), .ZN(n5559) );
  OR2_X1 U6726 ( .A1(n5209), .A2(n5556), .ZN(n5557) );
  NAND2_X1 U6727 ( .A1(n5892), .A2(n5557), .ZN(n5558) );
  AOI21_X1 U6728 ( .B1(n5559), .B2(n5558), .A(n5580), .ZN(n5566) );
  NAND2_X1 U6729 ( .A1(n6379), .A2(REIP_REG_21__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U6730 ( .A1(n6363), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5560)
         );
  OAI211_X1 U6731 ( .C1(n6355), .C2(n6004), .A(n5563), .B(n5560), .ZN(n5561)
         );
  AOI21_X1 U6732 ( .B1(n6008), .B2(n6360), .A(n5561), .ZN(n5562) );
  OAI21_X1 U6733 ( .B1(n5566), .B2(n6323), .A(n5562), .ZN(U2965) );
  OAI21_X1 U6734 ( .B1(n6006), .B2(n6428), .A(n5563), .ZN(n5564) );
  NOR3_X1 U6735 ( .A1(n5936), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n5935), 
        .ZN(n5941) );
  AOI211_X1 U6736 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5940), .A(n5564), .B(n5941), .ZN(n5565) );
  OAI21_X1 U6737 ( .B1(n5566), .B2(n6406), .A(n5565), .ZN(U2997) );
  INV_X1 U6738 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6647) );
  NAND3_X1 U6739 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5671) );
  INV_X1 U6740 ( .A(n5671), .ZN(n5568) );
  OAI21_X1 U6741 ( .B1(n5568), .B2(n5567), .A(n5986), .ZN(n5970) );
  NOR2_X1 U6742 ( .A1(n6647), .A2(n5970), .ZN(n5656) );
  AOI21_X1 U6743 ( .B1(n5673), .B2(n5568), .A(REIP_REG_27__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U6744 ( .A1(n5882), .A2(n6190), .ZN(n5578) );
  OAI22_X1 U6745 ( .A1(n6910), .A2(n6220), .B1(n6238), .B2(n5880), .ZN(n5576)
         );
  MUX2_X1 U6746 ( .A(n5569), .B(n5659), .S(EBX_REG_27__SCAN_IN), .Z(n5570) );
  OAI21_X1 U6747 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5774), .A(n5570), 
        .ZN(n5571) );
  INV_X1 U6748 ( .A(n5571), .ZN(n5574) );
  INV_X1 U6749 ( .A(n5832), .ZN(n5572) );
  OAI21_X1 U6750 ( .B1(n5574), .B2(n5573), .A(n5572), .ZN(n5916) );
  NOR2_X1 U6751 ( .A1(n5916), .A2(n6243), .ZN(n5575) );
  AOI211_X1 U6752 ( .C1(n6231), .C2(EBX_REG_27__SCAN_IN), .A(n5576), .B(n5575), 
        .ZN(n5577) );
  OAI211_X1 U6753 ( .C1(n5656), .C2(n5579), .A(n5578), .B(n5577), .ZN(U2800)
         );
  NOR2_X1 U6754 ( .A1(n5209), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5897)
         );
  NAND2_X1 U6755 ( .A1(n5580), .A2(n5897), .ZN(n5890) );
  INV_X1 U6756 ( .A(n5580), .ZN(n5581) );
  OAI21_X1 U6757 ( .B1(n5206), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5581), 
        .ZN(n5899) );
  NAND3_X1 U6758 ( .A1(n6039), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5582) );
  OAI22_X1 U6759 ( .A1(n5890), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5899), .B2(n5582), .ZN(n5583) );
  XNOR2_X1 U6760 ( .A(n5583), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5593)
         );
  INV_X1 U6761 ( .A(n5983), .ZN(n5587) );
  NOR2_X1 U6762 ( .A1(n6426), .A2(n6896), .ZN(n5589) );
  NAND3_X1 U6763 ( .A1(n5929), .A2(n5928), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5585) );
  INV_X1 U6764 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5584) );
  AOI21_X1 U6765 ( .B1(n5585), .B2(n5584), .A(n5756), .ZN(n5586) );
  AOI211_X1 U6766 ( .C1(n6405), .C2(n5587), .A(n5589), .B(n5586), .ZN(n5588)
         );
  OAI21_X1 U6767 ( .B1(n5593), .B2(n6406), .A(n5588), .ZN(U2994) );
  AOI21_X1 U6768 ( .B1(n6363), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5589), 
        .ZN(n5590) );
  OAI21_X1 U6769 ( .B1(n5975), .B2(n6355), .A(n5590), .ZN(n5591) );
  AOI21_X1 U6770 ( .B1(n5974), .B2(n6360), .A(n5591), .ZN(n5592) );
  OAI21_X1 U6771 ( .B1(n5593), .B2(n6323), .A(n5592), .ZN(U2962) );
  OR2_X1 U6772 ( .A1(n5594), .A2(n5598), .ZN(n5595) );
  MUX2_X1 U6773 ( .A(n5595), .B(n6051), .S(n6039), .Z(n6044) );
  AND2_X1 U6774 ( .A1(n5597), .A2(n5596), .ZN(n6038) );
  AND2_X1 U6775 ( .A1(n6038), .A2(n5598), .ZN(n5599) );
  NOR2_X1 U6776 ( .A1(n6044), .A2(n5599), .ZN(n5600) );
  XNOR2_X1 U6777 ( .A(n5600), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5611)
         );
  INV_X1 U6778 ( .A(n6115), .ZN(n5602) );
  NAND2_X1 U6779 ( .A1(n6363), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5601)
         );
  NAND2_X1 U6780 ( .A1(n6379), .A2(REIP_REG_18__SCAN_IN), .ZN(n5606) );
  OAI211_X1 U6781 ( .C1(n6355), .C2(n5602), .A(n5601), .B(n5606), .ZN(n5603)
         );
  AOI21_X1 U6782 ( .B1(n6244), .B2(n6360), .A(n5603), .ZN(n5604) );
  OAI21_X1 U6783 ( .B1(n5611), .B2(n6323), .A(n5604), .ZN(U2968) );
  INV_X1 U6784 ( .A(n6052), .ZN(n5605) );
  INV_X1 U6785 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6783) );
  OAI21_X1 U6786 ( .B1(n5605), .B2(n6051), .A(n6783), .ZN(n5609) );
  OAI21_X1 U6787 ( .B1(n6118), .B2(n6428), .A(n5606), .ZN(n5607) );
  AOI21_X1 U6788 ( .B1(n5609), .B2(n5608), .A(n5607), .ZN(n5610) );
  OAI21_X1 U6789 ( .B1(n5611), .B2(n6406), .A(n5610), .ZN(U3000) );
  INV_X1 U6790 ( .A(n5612), .ZN(n5613) );
  INV_X1 U6791 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U6792 ( .A1(n5613), .A2(n5668), .ZN(n5614) );
  NAND2_X1 U6793 ( .A1(n5705), .A2(n5614), .ZN(n5728) );
  AOI22_X1 U6794 ( .A1(n5683), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5618) );
  AOI22_X1 U6795 ( .A1(n3510), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5680), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5617) );
  AOI22_X1 U6796 ( .A1(n5629), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5682), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5616) );
  AOI22_X1 U6797 ( .A1(n3270), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3255), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n5615) );
  NAND4_X1 U6798 ( .A1(n5618), .A2(n5617), .A3(n5616), .A4(n5615), .ZN(n5626)
         );
  AOI22_X1 U6799 ( .A1(n3248), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3511), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5624) );
  AOI22_X1 U6800 ( .A1(n5619), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3607), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5623) );
  AOI22_X1 U6801 ( .A1(n4729), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5622) );
  AOI22_X1 U6802 ( .A1(n5620), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5621) );
  NAND4_X1 U6803 ( .A1(n5624), .A2(n5623), .A3(n5622), .A4(n5621), .ZN(n5625)
         );
  NOR2_X1 U6804 ( .A1(n5626), .A2(n5625), .ZN(n5678) );
  NOR2_X1 U6805 ( .A1(n5628), .A2(n5627), .ZN(n5649) );
  AOI22_X1 U6806 ( .A1(n5681), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n5629), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5633) );
  AOI22_X1 U6807 ( .A1(n5680), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5692), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n5632) );
  AOI22_X1 U6808 ( .A1(n5688), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3607), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5631) );
  AOI22_X1 U6809 ( .A1(n3270), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n5630) );
  NAND4_X1 U6810 ( .A1(n5633), .A2(n5632), .A3(n5631), .A4(n5630), .ZN(n5641)
         );
  AOI22_X1 U6811 ( .A1(n3248), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5634), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n5639) );
  AOI22_X1 U6812 ( .A1(n5691), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n5638) );
  AOI22_X1 U6813 ( .A1(n5682), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5637) );
  AOI22_X1 U6814 ( .A1(n3241), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5635), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5636) );
  NAND4_X1 U6815 ( .A1(n5639), .A2(n5638), .A3(n5637), .A4(n5636), .ZN(n5640)
         );
  OR2_X1 U6816 ( .A1(n5641), .A2(n5640), .ZN(n5648) );
  NAND2_X1 U6817 ( .A1(n5649), .A2(n5648), .ZN(n5677) );
  XNOR2_X1 U6818 ( .A(n5678), .B(n5677), .ZN(n5644) );
  AOI21_X1 U6819 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6814), .A(n5706), 
        .ZN(n5643) );
  NAND2_X1 U6820 ( .A1(n5785), .A2(EAX_REG_29__SCAN_IN), .ZN(n5642) );
  OAI211_X1 U6821 ( .C1(n5644), .C2(n5650), .A(n5643), .B(n5642), .ZN(n5645)
         );
  OAI21_X1 U6822 ( .B1(n5646), .B2(n5728), .A(n5645), .ZN(n5655) );
  XNOR2_X1 U6823 ( .A(n5647), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5872)
         );
  OAI21_X1 U6824 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5870), .A(n5703), .ZN(
        n5653) );
  XNOR2_X1 U6825 ( .A(n5649), .B(n5648), .ZN(n5651) );
  NOR2_X1 U6826 ( .A1(n5651), .A2(n5650), .ZN(n5652) );
  AOI211_X1 U6827 ( .C1(n5785), .C2(EAX_REG_28__SCAN_IN), .A(n5653), .B(n5652), 
        .ZN(n5654) );
  AOI21_X1 U6828 ( .B1(n5706), .B2(n5872), .A(n5654), .ZN(n5829) );
  NAND2_X1 U6829 ( .A1(n5830), .A2(n5829), .ZN(n5828) );
  NOR2_X2 U6830 ( .A1(n5828), .A2(n5655), .ZN(n5787) );
  AOI21_X1 U6831 ( .B1(n5655), .B2(n5828), .A(n5787), .ZN(n5730) );
  INV_X1 U6832 ( .A(n5730), .ZN(n5859) );
  NAND2_X1 U6833 ( .A1(n5656), .A2(REIP_REG_28__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U6834 ( .A1(n5657), .A2(n6110), .ZN(n5717) );
  INV_X1 U6835 ( .A(n5717), .ZN(n5841) );
  INV_X1 U6836 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6875) );
  NAND2_X1 U6837 ( .A1(n3112), .A2(n6875), .ZN(n5660) );
  OAI211_X1 U6838 ( .C1(EBX_REG_28__SCAN_IN), .C2(n5773), .A(n5660), .B(n5659), 
        .ZN(n5661) );
  OAI21_X1 U6839 ( .B1(n5662), .B2(EBX_REG_28__SCAN_IN), .A(n5661), .ZN(n5831)
         );
  INV_X1 U6840 ( .A(n5834), .ZN(n5667) );
  OAI22_X1 U6841 ( .A1(n5774), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n5773), .ZN(n5710) );
  NAND2_X1 U6842 ( .A1(n5710), .A2(n5659), .ZN(n5664) );
  INV_X1 U6843 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5847) );
  NOR2_X1 U6844 ( .A1(n5659), .A2(n5847), .ZN(n5768) );
  INV_X1 U6845 ( .A(n5768), .ZN(n5663) );
  NAND2_X1 U6846 ( .A1(n5664), .A2(n5663), .ZN(n5665) );
  INV_X1 U6847 ( .A(n5665), .ZN(n5666) );
  OR2_X2 U6848 ( .A1(n5834), .A2(n5665), .ZN(n5772) );
  OAI22_X1 U6849 ( .A1(n5668), .A2(n6220), .B1(n6238), .B2(n5728), .ZN(n5669)
         );
  AOI21_X1 U6850 ( .B1(EBX_REG_29__SCAN_IN), .B2(n6231), .A(n5669), .ZN(n5670)
         );
  OAI21_X1 U6851 ( .B1(n5846), .B2(n6243), .A(n5670), .ZN(n5675) );
  NOR2_X1 U6852 ( .A1(n5671), .A2(n6647), .ZN(n5672) );
  NAND2_X1 U6853 ( .A1(n5673), .A2(n5672), .ZN(n5838) );
  INV_X1 U6854 ( .A(REIP_REG_28__SCAN_IN), .ZN(n5869) );
  NOR3_X1 U6855 ( .A1(n5838), .A2(REIP_REG_29__SCAN_IN), .A3(n5869), .ZN(n5674) );
  OAI21_X1 U6856 ( .B1(n5859), .B2(n6199), .A(n5676), .ZN(U2798) );
  NOR2_X1 U6857 ( .A1(n5678), .A2(n5677), .ZN(n5700) );
  AOI22_X1 U6858 ( .A1(n3241), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5679), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5687) );
  AOI22_X1 U6859 ( .A1(n5681), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n5680), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5686) );
  AOI22_X1 U6860 ( .A1(n5683), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5682), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5685) );
  AOI22_X1 U6861 ( .A1(n3607), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3255), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5684) );
  NAND4_X1 U6862 ( .A1(n5687), .A2(n5686), .A3(n5685), .A4(n5684), .ZN(n5698)
         );
  AOI22_X1 U6863 ( .A1(n5688), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5696) );
  AOI22_X1 U6864 ( .A1(n3248), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5689), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5695) );
  AOI22_X1 U6865 ( .A1(n5691), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n5690), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5694) );
  AOI22_X1 U6866 ( .A1(n5692), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3518), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5693) );
  NAND4_X1 U6867 ( .A1(n5696), .A2(n5695), .A3(n5694), .A4(n5693), .ZN(n5697)
         );
  NOR2_X1 U6868 ( .A1(n5698), .A2(n5697), .ZN(n5699) );
  XNOR2_X1 U6869 ( .A(n5700), .B(n5699), .ZN(n5702) );
  NAND2_X1 U6870 ( .A1(n5702), .A2(n5701), .ZN(n5709) );
  OAI21_X1 U6871 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6842), .A(n5703), .ZN(
        n5704) );
  AOI21_X1 U6872 ( .B1(n5785), .B2(EAX_REG_30__SCAN_IN), .A(n5704), .ZN(n5708)
         );
  XNOR2_X1 U6873 ( .A(n5705), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5746)
         );
  AND2_X1 U6874 ( .A1(n5746), .A2(n5706), .ZN(n5707) );
  AOI21_X1 U6875 ( .B1(n5709), .B2(n5708), .A(n5707), .ZN(n5786) );
  XOR2_X1 U6876 ( .A(n5786), .B(n5787), .Z(n5749) );
  INV_X1 U6877 ( .A(n5749), .ZN(n5856) );
  AND2_X1 U6878 ( .A1(n5773), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5711)
         );
  AOI21_X1 U6879 ( .B1(n5774), .B2(EBX_REG_30__SCAN_IN), .A(n5711), .ZN(n5771)
         );
  XNOR2_X1 U6880 ( .A(n5712), .B(n5771), .ZN(n5751) );
  OR2_X1 U6881 ( .A1(n5751), .A2(n6243), .ZN(n5723) );
  NAND2_X1 U6882 ( .A1(REIP_REG_29__SCAN_IN), .A2(REIP_REG_28__SCAN_IN), .ZN(
        n5713) );
  NOR2_X1 U6883 ( .A1(n5838), .A2(n5713), .ZN(n5821) );
  INV_X1 U6884 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6656) );
  INV_X1 U6885 ( .A(n5746), .ZN(n5714) );
  OAI22_X1 U6886 ( .A1(n6842), .A2(n6220), .B1(n6238), .B2(n5714), .ZN(n5715)
         );
  INV_X1 U6887 ( .A(n5715), .ZN(n5720) );
  NAND2_X1 U6888 ( .A1(n6231), .A2(EBX_REG_30__SCAN_IN), .ZN(n5719) );
  INV_X1 U6889 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6998) );
  NAND2_X1 U6890 ( .A1(n6216), .A2(n6998), .ZN(n5716) );
  NAND2_X1 U6891 ( .A1(n5717), .A2(n5716), .ZN(n5823) );
  NAND2_X1 U6892 ( .A1(n5823), .A2(REIP_REG_30__SCAN_IN), .ZN(n5718) );
  NAND3_X1 U6893 ( .A1(n5720), .A2(n5719), .A3(n5718), .ZN(n5721) );
  OAI21_X1 U6894 ( .B1(n5856), .B2(n6199), .A(n3114), .ZN(U2797) );
  INV_X1 U6895 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5724) );
  OAI222_X1 U6896 ( .A1(n5850), .A2(n5856), .B1(n5852), .B2(n5751), .C1(n5724), 
        .C2(n5848), .ZN(U2829) );
  NAND2_X1 U6897 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5908) );
  NOR2_X2 U6898 ( .A1(n5877), .A2(n5908), .ZN(n5766) );
  INV_X1 U6899 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6943) );
  NAND2_X1 U6900 ( .A1(n6943), .A2(n6875), .ZN(n5909) );
  OR3_X1 U6901 ( .A1(n6039), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n5909), 
        .ZN(n5762) );
  NOR2_X1 U6902 ( .A1(n5863), .A2(n5762), .ZN(n5744) );
  NOR2_X1 U6903 ( .A1(n5766), .A2(n5744), .ZN(n5726) );
  XOR2_X1 U6904 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .B(n5726), .Z(n5743) );
  OR2_X1 U6905 ( .A1(n6426), .A2(n6998), .ZN(n5732) );
  NAND2_X1 U6906 ( .A1(n6363), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5727)
         );
  OAI211_X1 U6907 ( .C1(n6355), .C2(n5728), .A(n5732), .B(n5727), .ZN(n5729)
         );
  AOI21_X1 U6908 ( .B1(n5730), .B2(n6360), .A(n5729), .ZN(n5731) );
  OAI21_X1 U6909 ( .B1(n5743), .B2(n6323), .A(n5731), .ZN(U2957) );
  INV_X1 U6910 ( .A(n5846), .ZN(n5741) );
  INV_X1 U6911 ( .A(n5732), .ZN(n5740) );
  NOR3_X1 U6912 ( .A1(n5936), .A2(n5733), .A3(n5734), .ZN(n5920) );
  INV_X1 U6913 ( .A(n5908), .ZN(n5752) );
  AOI21_X1 U6914 ( .B1(n5920), .B2(n5752), .A(INSTADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n5738) );
  NAND2_X1 U6915 ( .A1(n6374), .A2(n5734), .ZN(n5735) );
  AND2_X1 U6916 ( .A1(n5756), .A2(n5735), .ZN(n5912) );
  INV_X1 U6917 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5736) );
  AOI21_X1 U6918 ( .B1(n6374), .B2(n5908), .A(n5736), .ZN(n5737) );
  AND2_X1 U6919 ( .A1(n5912), .A2(n5737), .ZN(n5755) );
  NOR2_X1 U6920 ( .A1(n5738), .A2(n5755), .ZN(n5739) );
  AOI211_X1 U6921 ( .C1(n6405), .C2(n5741), .A(n5740), .B(n5739), .ZN(n5742)
         );
  OAI21_X1 U6922 ( .B1(n5743), .B2(n6406), .A(n5742), .ZN(U2989) );
  MUX2_X1 U6923 ( .A(n5744), .B(n5766), .S(INSTADDRPOINTER_REG_29__SCAN_IN), 
        .Z(n5745) );
  XNOR2_X1 U6924 ( .A(n5745), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5761)
         );
  NAND2_X1 U6925 ( .A1(n6332), .A2(n5746), .ZN(n5747) );
  NAND2_X1 U6926 ( .A1(n6379), .A2(REIP_REG_30__SCAN_IN), .ZN(n5753) );
  OAI211_X1 U6927 ( .C1(n6842), .C2(n6339), .A(n5747), .B(n5753), .ZN(n5748)
         );
  AOI21_X1 U6928 ( .B1(n5749), .B2(n6360), .A(n5748), .ZN(n5750) );
  OAI21_X1 U6929 ( .B1(n5761), .B2(n6323), .A(n5750), .ZN(U2956) );
  INV_X1 U6930 ( .A(n5751), .ZN(n5759) );
  INV_X1 U6931 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6993) );
  NAND4_X1 U6932 ( .A1(n5920), .A2(n5752), .A3(INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n6993), .ZN(n5754) );
  NAND2_X1 U6933 ( .A1(n5754), .A2(n5753), .ZN(n5758) );
  AOI211_X1 U6934 ( .C1(n6429), .C2(n5756), .A(n6993), .B(n5755), .ZN(n5757)
         );
  AOI211_X1 U6935 ( .C1(n6405), .C2(n5759), .A(n5758), .B(n5757), .ZN(n5760)
         );
  OAI21_X1 U6936 ( .B1(n5761), .B2(n6406), .A(n5760), .ZN(U2988) );
  NAND2_X1 U6937 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5777) );
  INV_X1 U6938 ( .A(n5777), .ZN(n5765) );
  INV_X1 U6939 ( .A(n5548), .ZN(n5763) );
  NOR4_X1 U6940 ( .A1(n5763), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A4(n5762), .ZN(n5764) );
  AOI21_X1 U6941 ( .B1(n5766), .B2(n5765), .A(n5764), .ZN(n5767) );
  XOR2_X1 U6942 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .B(n5767), .Z(n5795) );
  AOI21_X1 U6943 ( .B1(n5834), .B2(n5769), .A(n5768), .ZN(n5770) );
  OAI21_X1 U6944 ( .B1(n5772), .B2(n5771), .A(n5770), .ZN(n5776) );
  OAI22_X1 U6945 ( .A1(n5774), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n5773), .ZN(n5775) );
  XNOR2_X1 U6946 ( .A(n5776), .B(n5775), .ZN(n5843) );
  NOR2_X1 U6947 ( .A1(n5908), .A2(n5777), .ZN(n5779) );
  INV_X1 U6948 ( .A(n5779), .ZN(n5778) );
  INV_X1 U6949 ( .A(n5912), .ZN(n5919) );
  AOI21_X1 U6950 ( .B1(n6374), .B2(n5778), .A(n5919), .ZN(n5781) );
  INV_X1 U6951 ( .A(REIP_REG_31__SCAN_IN), .ZN(n5820) );
  OR2_X1 U6952 ( .A1(n6426), .A2(n5820), .ZN(n5791) );
  NAND3_X1 U6953 ( .A1(n5920), .A2(n5779), .A3(n6859), .ZN(n5780) );
  OAI211_X1 U6954 ( .C1(n5781), .C2(n6859), .A(n5791), .B(n5780), .ZN(n5782)
         );
  AOI21_X1 U6955 ( .B1(n5843), .B2(n6405), .A(n5782), .ZN(n5783) );
  OAI21_X1 U6956 ( .B1(n5795), .B2(n6406), .A(n5783), .ZN(U2987) );
  AOI22_X1 U6957 ( .A1(n5785), .A2(EAX_REG_31__SCAN_IN), .B1(n5784), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U6958 ( .A1(n5787), .A2(n5786), .ZN(n5788) );
  XOR2_X1 U6959 ( .A(n5789), .B(n5788), .Z(n5814) );
  NAND2_X1 U6960 ( .A1(n6363), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5790)
         );
  OAI211_X1 U6961 ( .C1(n6355), .C2(n5792), .A(n5791), .B(n5790), .ZN(n5793)
         );
  AOI21_X1 U6962 ( .B1(n5814), .B2(n6360), .A(n5793), .ZN(n5794) );
  OAI21_X1 U6963 ( .B1(n5795), .B2(n6323), .A(n5794), .ZN(U2955) );
  NAND3_X1 U6964 ( .A1(n5814), .A2(n5797), .A3(n5796), .ZN(n5799) );
  AOI22_X1 U6965 ( .A1(n6247), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6250), .ZN(n5798) );
  NAND2_X1 U6966 ( .A1(n5799), .A2(n5798), .ZN(U2860) );
  NOR3_X1 U6967 ( .A1(n5801), .A2(n3399), .A3(n5800), .ZN(n5802) );
  AOI21_X1 U6968 ( .B1(n5803), .B2(n6872), .A(n5802), .ZN(n5804) );
  OAI21_X1 U6969 ( .B1(n5948), .B2(n5805), .A(n5804), .ZN(n6554) );
  NOR2_X1 U6970 ( .A1(n5806), .A2(n6431), .ZN(n5809) );
  AOI222_X1 U6971 ( .A1(n6554), .A2(n6079), .B1(n5810), .B2(n5809), .C1(n5808), 
        .C2(n5807), .ZN(n5813) );
  OAI22_X1 U6972 ( .A1(n5813), .A2(n5812), .B1(n5811), .B2(n6872), .ZN(U3460)
         );
  NAND2_X1 U6973 ( .A1(n5814), .A2(n6190), .ZN(n5827) );
  NAND2_X1 U6974 ( .A1(n5815), .A2(EBX_REG_31__SCAN_IN), .ZN(n5816) );
  OAI22_X1 U6975 ( .A1(n5818), .A2(n6220), .B1(n5817), .B2(n5816), .ZN(n5819)
         );
  AOI21_X1 U6976 ( .B1(n5843), .B2(n6214), .A(n5819), .ZN(n5826) );
  NAND3_X1 U6977 ( .A1(n5821), .A2(REIP_REG_30__SCAN_IN), .A3(n5820), .ZN(
        n5825) );
  NOR2_X1 U6978 ( .A1(n6209), .A2(REIP_REG_30__SCAN_IN), .ZN(n5822) );
  OAI21_X1 U6979 ( .B1(n5823), .B2(n5822), .A(REIP_REG_31__SCAN_IN), .ZN(n5824) );
  NAND4_X1 U6980 ( .A1(n5827), .A2(n5826), .A3(n5825), .A4(n5824), .ZN(U2796)
         );
  OAI21_X1 U6981 ( .B1(n5830), .B2(n5829), .A(n5828), .ZN(n5875) );
  OR2_X1 U6982 ( .A1(n5832), .A2(n5831), .ZN(n5833) );
  NAND2_X1 U6983 ( .A1(n5834), .A2(n5833), .ZN(n5905) );
  INV_X1 U6984 ( .A(n5872), .ZN(n5835) );
  OAI22_X1 U6985 ( .A1(n5870), .A2(n6220), .B1(n6238), .B2(n5835), .ZN(n5836)
         );
  AOI21_X1 U6986 ( .B1(n6231), .B2(EBX_REG_28__SCAN_IN), .A(n5836), .ZN(n5837)
         );
  OAI21_X1 U6987 ( .B1(n5905), .B2(n6243), .A(n5837), .ZN(n5840) );
  NOR2_X1 U6988 ( .A1(n5838), .A2(REIP_REG_28__SCAN_IN), .ZN(n5839) );
  AOI211_X1 U6989 ( .C1(n5841), .C2(REIP_REG_28__SCAN_IN), .A(n5840), .B(n5839), .ZN(n5842) );
  OAI21_X1 U6990 ( .B1(n5875), .B2(n6199), .A(n5842), .ZN(U2799) );
  INV_X1 U6991 ( .A(n5843), .ZN(n5845) );
  INV_X1 U6992 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5844) );
  OAI22_X1 U6993 ( .A1(n5845), .A2(n5852), .B1(n5848), .B2(n5844), .ZN(U2828)
         );
  OAI222_X1 U6994 ( .A1(n5850), .A2(n5859), .B1(n5848), .B2(n5847), .C1(n5846), 
        .C2(n5852), .ZN(U2830) );
  INV_X1 U6995 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5849) );
  OAI222_X1 U6996 ( .A1(n5849), .A2(n5848), .B1(n5852), .B2(n5905), .C1(n5875), 
        .C2(n5850), .ZN(U2831) );
  INV_X1 U6997 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5853) );
  OAI222_X1 U6998 ( .A1(n5853), .A2(n5848), .B1(n5852), .B2(n5916), .C1(n5851), 
        .C2(n5850), .ZN(U2832) );
  AOI22_X1 U6999 ( .A1(n6247), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6250), .ZN(n5855) );
  NAND2_X1 U7000 ( .A1(n6251), .A2(DATAI_14_), .ZN(n5854) );
  OAI211_X1 U7001 ( .C1(n5856), .C2(n5862), .A(n5855), .B(n5854), .ZN(U2861)
         );
  AOI22_X1 U7002 ( .A1(n6247), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6250), .ZN(n5858) );
  NAND2_X1 U7003 ( .A1(n6251), .A2(DATAI_13_), .ZN(n5857) );
  OAI211_X1 U7004 ( .C1(n5859), .C2(n5862), .A(n5858), .B(n5857), .ZN(U2862)
         );
  AOI22_X1 U7005 ( .A1(n6247), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6250), .ZN(n5861) );
  NAND2_X1 U7006 ( .A1(n6251), .A2(DATAI_12_), .ZN(n5860) );
  OAI211_X1 U7007 ( .C1(n5875), .C2(n5862), .A(n5861), .B(n5860), .ZN(U2863)
         );
  NAND3_X1 U7008 ( .A1(n5863), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n6039), .ZN(n5867) );
  INV_X1 U7009 ( .A(n5864), .ZN(n5866) );
  NAND3_X1 U7010 ( .A1(n5866), .A2(n5206), .A3(n5865), .ZN(n5876) );
  AOI22_X1 U7011 ( .A1(n5867), .A2(n5876), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n6775), .ZN(n5868) );
  XNOR2_X1 U7012 ( .A(n5868), .B(n6875), .ZN(n5914) );
  NAND2_X1 U7013 ( .A1(n5914), .A2(n6358), .ZN(n5874) );
  NOR2_X1 U7014 ( .A1(n6426), .A2(n5869), .ZN(n5906) );
  NOR2_X1 U7015 ( .A1(n6339), .A2(n5870), .ZN(n5871) );
  AOI211_X1 U7016 ( .C1(n6332), .C2(n5872), .A(n5906), .B(n5871), .ZN(n5873)
         );
  OAI211_X1 U7017 ( .C1(n5901), .C2(n5875), .A(n5874), .B(n5873), .ZN(U2958)
         );
  NAND2_X1 U7018 ( .A1(n5877), .A2(n5876), .ZN(n5878) );
  XNOR2_X1 U7019 ( .A(n5878), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5923)
         );
  NOR2_X1 U7020 ( .A1(n6426), .A2(n6647), .ZN(n5918) );
  AOI21_X1 U7021 ( .B1(n6363), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5918), 
        .ZN(n5879) );
  OAI21_X1 U7022 ( .B1(n5880), .B2(n6355), .A(n5879), .ZN(n5881) );
  AOI21_X1 U7023 ( .B1(n5882), .B2(n6360), .A(n5881), .ZN(n5883) );
  OAI21_X1 U7024 ( .B1(n5923), .B2(n6323), .A(n5883), .ZN(U2959) );
  OAI21_X1 U7025 ( .B1(n6339), .B2(n5885), .A(n5884), .ZN(n5887) );
  NOR2_X1 U7026 ( .A1(n5967), .A2(n5901), .ZN(n5886) );
  AOI211_X1 U7027 ( .C1(n6332), .C2(n5962), .A(n5887), .B(n5886), .ZN(n5888)
         );
  OAI21_X1 U7028 ( .B1(n6323), .B2(n5889), .A(n5888), .ZN(U2960) );
  INV_X1 U7029 ( .A(n5928), .ZN(n5891) );
  OAI21_X1 U7030 ( .B1(n5892), .B2(n5891), .A(n5890), .ZN(n5893) );
  XNOR2_X1 U7031 ( .A(n5893), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5932)
         );
  NAND2_X1 U7032 ( .A1(n6379), .A2(REIP_REG_23__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7033 ( .A1(n6363), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5894)
         );
  OAI211_X1 U7034 ( .C1(n6355), .C2(n5991), .A(n5924), .B(n5894), .ZN(n5895)
         );
  AOI21_X1 U7035 ( .B1(n5988), .B2(n6360), .A(n5895), .ZN(n5896) );
  OAI21_X1 U7036 ( .B1(n5932), .B2(n6323), .A(n5896), .ZN(U2963) );
  AOI21_X1 U7037 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n6039), .A(n5897), 
        .ZN(n5898) );
  XNOR2_X1 U7038 ( .A(n5899), .B(n5898), .ZN(n5944) );
  NAND2_X1 U7039 ( .A1(n6379), .A2(REIP_REG_22__SCAN_IN), .ZN(n5933) );
  OAI21_X1 U7040 ( .B1(n6339), .B2(n5900), .A(n5933), .ZN(n5903) );
  NOR2_X1 U7041 ( .A1(n6000), .A2(n5901), .ZN(n5902) );
  AOI211_X1 U7042 ( .C1(n6332), .C2(n5993), .A(n5903), .B(n5902), .ZN(n5904)
         );
  OAI21_X1 U7043 ( .B1(n5944), .B2(n6323), .A(n5904), .ZN(U2964) );
  INV_X1 U7044 ( .A(n5905), .ZN(n5907) );
  AOI21_X1 U7045 ( .B1(n5907), .B2(n6405), .A(n5906), .ZN(n5911) );
  NAND3_X1 U7046 ( .A1(n5920), .A2(n5909), .A3(n5908), .ZN(n5910) );
  OAI211_X1 U7047 ( .C1(n5912), .C2(n6875), .A(n5911), .B(n5910), .ZN(n5913)
         );
  AOI21_X1 U7048 ( .B1(n5914), .B2(n6434), .A(n5913), .ZN(n5915) );
  INV_X1 U7049 ( .A(n5915), .ZN(U2990) );
  NOR2_X1 U7050 ( .A1(n5916), .A2(n6428), .ZN(n5917) );
  AOI211_X1 U7051 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5919), .A(n5918), .B(n5917), .ZN(n5922) );
  NAND2_X1 U7052 ( .A1(n5920), .A2(n6943), .ZN(n5921) );
  OAI211_X1 U7053 ( .C1(n5923), .C2(n6406), .A(n5922), .B(n5921), .ZN(U2991)
         );
  OAI21_X1 U7054 ( .B1(n5984), .B2(n6428), .A(n5924), .ZN(n5925) );
  AOI21_X1 U7055 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5926), .A(n5925), 
        .ZN(n5931) );
  INV_X1 U7056 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5927) );
  NAND3_X1 U7057 ( .A1(n5929), .A2(n5928), .A3(n5927), .ZN(n5930) );
  OAI211_X1 U7058 ( .C1(n5932), .C2(n6406), .A(n5931), .B(n5930), .ZN(U2995)
         );
  INV_X1 U7059 ( .A(n6003), .ZN(n5939) );
  INV_X1 U7060 ( .A(n5933), .ZN(n5938) );
  NOR4_X1 U7061 ( .A1(n5936), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n5935), 
        .A4(n5934), .ZN(n5937) );
  AOI211_X1 U7062 ( .C1(n6405), .C2(n5939), .A(n5938), .B(n5937), .ZN(n5943)
         );
  OAI21_X1 U7063 ( .B1(n5941), .B2(n5940), .A(INSTADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n5942) );
  OAI211_X1 U7064 ( .C1(n5944), .C2(n6406), .A(n5943), .B(n5942), .ZN(U2996)
         );
  OAI211_X1 U7065 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n5946), .A(n5945), .B(
        n6445), .ZN(n5947) );
  OAI21_X1 U7066 ( .B1(n6670), .B2(n5948), .A(n5947), .ZN(n5949) );
  MUX2_X1 U7067 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5949), .S(n6675), 
        .Z(U3464) );
  XNOR2_X1 U7068 ( .A(n5950), .B(n6489), .ZN(n5952) );
  OAI22_X1 U7069 ( .A1(n5952), .A2(n6492), .B1(n5951), .B2(n6670), .ZN(n5953)
         );
  MUX2_X1 U7070 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5953), .S(n6675), 
        .Z(U3463) );
  INV_X1 U7071 ( .A(n5954), .ZN(n5957) );
  OAI22_X1 U7072 ( .A1(n5957), .A2(n5956), .B1(n5955), .B2(n6581), .ZN(n5958)
         );
  MUX2_X1 U7073 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5958), .S(n6084), 
        .Z(U3456) );
  AND2_X1 U7074 ( .A1(DATAO_REG_31__SCAN_IN), .A2(n6280), .ZN(U2892) );
  AOI21_X1 U7075 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n5960), .A(n5959), .ZN(
        n5961) );
  INV_X1 U7076 ( .A(n5961), .ZN(U2788) );
  AOI22_X1 U7077 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n6235), .B1(n5962), 
        .B2(n5994), .ZN(n5972) );
  INV_X1 U7078 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5963) );
  OAI21_X1 U7079 ( .B1(n5965), .B2(n5964), .A(n5963), .ZN(n5969) );
  OAI22_X1 U7080 ( .A1(n5967), .A2(n6199), .B1(n5966), .B2(n6243), .ZN(n5968)
         );
  AOI21_X1 U7081 ( .B1(n5970), .B2(n5969), .A(n5968), .ZN(n5971) );
  OAI211_X1 U7082 ( .C1(n5973), .C2(n6175), .A(n5972), .B(n5971), .ZN(U2801)
         );
  NAND2_X1 U7083 ( .A1(n5974), .A2(n6190), .ZN(n5979) );
  OAI22_X1 U7084 ( .A1(n5976), .A2(n6220), .B1(n6238), .B2(n5975), .ZN(n5977)
         );
  AOI21_X1 U7085 ( .B1(EBX_REG_24__SCAN_IN), .B2(n6231), .A(n5977), .ZN(n5978)
         );
  OAI211_X1 U7086 ( .C1(n5986), .C2(n6896), .A(n5979), .B(n5978), .ZN(n5981)
         );
  NOR2_X1 U7087 ( .A1(n5981), .A2(n5980), .ZN(n5982) );
  OAI21_X1 U7088 ( .B1(n5983), .B2(n6243), .A(n5982), .ZN(U2803) );
  AOI22_X1 U7089 ( .A1(EBX_REG_23__SCAN_IN), .A2(n6231), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6235), .ZN(n5990) );
  INV_X1 U7090 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6880) );
  NOR2_X1 U7091 ( .A1(n6880), .A2(n5992), .ZN(n5998) );
  AOI21_X1 U7092 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5998), .A(
        REIP_REG_23__SCAN_IN), .ZN(n5985) );
  OAI22_X1 U7093 ( .A1(n5986), .A2(n5985), .B1(n5984), .B2(n6243), .ZN(n5987)
         );
  AOI21_X1 U7094 ( .B1(n5988), .B2(n6190), .A(n5987), .ZN(n5989) );
  OAI211_X1 U7095 ( .C1(n5991), .C2(n6238), .A(n5990), .B(n5989), .ZN(U2804)
         );
  NOR2_X1 U7096 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5992), .ZN(n6009) );
  INV_X1 U7097 ( .A(REIP_REG_22__SCAN_IN), .ZN(n5997) );
  INV_X1 U7098 ( .A(n6238), .ZN(n5994) );
  AOI22_X1 U7099 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n6235), .B1(n3111), 
        .B2(n5993), .ZN(n5995) );
  OAI21_X1 U7100 ( .B1(n4863), .B2(n6175), .A(n5995), .ZN(n5996) );
  AOI21_X1 U7101 ( .B1(n5998), .B2(n5997), .A(n5996), .ZN(n5999) );
  OAI21_X1 U7102 ( .B1(n6000), .B2(n6199), .A(n5999), .ZN(n6001) );
  AOI221_X1 U7103 ( .B1(n6018), .B2(REIP_REG_22__SCAN_IN), .C1(n6009), .C2(
        REIP_REG_22__SCAN_IN), .A(n6001), .ZN(n6002) );
  OAI21_X1 U7104 ( .B1(n6003), .B2(n6243), .A(n6002), .ZN(U2805) );
  INV_X1 U7105 ( .A(n6004), .ZN(n6005) );
  AOI22_X1 U7106 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6231), .B1(n6005), .B2(n5994), .ZN(n6013) );
  AOI22_X1 U7107 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n6235), .B1(
        REIP_REG_21__SCAN_IN), .B2(n6018), .ZN(n6012) );
  NOR2_X1 U7108 ( .A1(n6006), .A2(n6243), .ZN(n6007) );
  AOI21_X1 U7109 ( .B1(n6008), .B2(n6190), .A(n6007), .ZN(n6011) );
  INV_X1 U7110 ( .A(n6009), .ZN(n6010) );
  NAND4_X1 U7111 ( .A1(n6013), .A2(n6012), .A3(n6011), .A4(n6010), .ZN(U2806)
         );
  AOI22_X1 U7112 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6231), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6235), .ZN(n6024) );
  INV_X1 U7113 ( .A(n6014), .ZN(n6017) );
  INV_X1 U7114 ( .A(n6015), .ZN(n6016) );
  AOI22_X1 U7115 ( .A1(n6017), .A2(n6190), .B1(n6214), .B2(n6016), .ZN(n6023)
         );
  OAI21_X1 U7116 ( .B1(REIP_REG_20__SCAN_IN), .B2(n6019), .A(n6018), .ZN(n6022) );
  NAND2_X1 U7117 ( .A1(n6020), .A2(n5994), .ZN(n6021) );
  NAND4_X1 U7118 ( .A1(n6024), .A2(n6023), .A3(n6022), .A4(n6021), .ZN(U2807)
         );
  AOI22_X1 U7119 ( .A1(n6111), .A2(n6113), .B1(n6110), .B2(n6109), .ZN(n6034)
         );
  AOI21_X1 U7120 ( .B1(n6235), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6207), 
        .ZN(n6025) );
  INV_X1 U7121 ( .A(n6025), .ZN(n6029) );
  OAI22_X1 U7122 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6027), .B1(n6026), .B2(
        n6238), .ZN(n6028) );
  AOI211_X1 U7123 ( .C1(EBX_REG_19__SCAN_IN), .C2(n6231), .A(n6029), .B(n6028), 
        .ZN(n6033) );
  INV_X1 U7124 ( .A(n6030), .ZN(n6031) );
  AOI22_X1 U7125 ( .A1(n6035), .A2(n6190), .B1(n6214), .B2(n6031), .ZN(n6032)
         );
  OAI211_X1 U7126 ( .C1(n6034), .C2(n6639), .A(n6033), .B(n6032), .ZN(U2808)
         );
  AOI22_X1 U7127 ( .A1(n6035), .A2(n6248), .B1(n6247), .B2(DATAI_19_), .ZN(
        n6037) );
  AOI22_X1 U7128 ( .A1(n6251), .A2(DATAI_3_), .B1(n6250), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7129 ( .A1(n6037), .A2(n6036), .ZN(U2872) );
  AOI22_X1 U7130 ( .A1(n6379), .A2(REIP_REG_17__SCAN_IN), .B1(n6363), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6046) );
  INV_X1 U7131 ( .A(n6038), .ZN(n6043) );
  XNOR2_X1 U7132 ( .A(n6039), .B(n6051), .ZN(n6040) );
  OAI21_X1 U7133 ( .B1(n6043), .B2(n6041), .A(n6040), .ZN(n6042) );
  OAI21_X1 U7134 ( .B1(n6044), .B2(n6043), .A(n6042), .ZN(n6047) );
  AOI22_X1 U7135 ( .A1(n6047), .A2(n6358), .B1(n6360), .B2(n6249), .ZN(n6045)
         );
  OAI211_X1 U7136 ( .C1(n6355), .C2(n6127), .A(n6046), .B(n6045), .ZN(U2969)
         );
  AOI22_X1 U7137 ( .A1(n6047), .A2(n6434), .B1(n6405), .B2(n6124), .ZN(n6054)
         );
  INV_X1 U7138 ( .A(n6048), .ZN(n6050) );
  NOR2_X1 U7139 ( .A1(n6426), .A2(n6917), .ZN(n6049) );
  AOI221_X1 U7140 ( .B1(n6052), .B2(n6051), .C1(n6050), .C2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A(n6049), .ZN(n6053) );
  NAND2_X1 U7141 ( .A1(n6054), .A2(n6053), .ZN(U3001) );
  NAND2_X1 U7142 ( .A1(n6865), .A2(n6055), .ZN(n6069) );
  AOI21_X1 U7143 ( .B1(n6057), .B2(n6405), .A(n6056), .ZN(n6068) );
  NAND3_X1 U7144 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n6076), .ZN(n6071) );
  NOR2_X1 U7145 ( .A1(n6861), .A2(n6058), .ZN(n6060) );
  OAI21_X1 U7146 ( .B1(n6060), .B2(n6059), .A(n6371), .ZN(n6061) );
  AOI21_X1 U7147 ( .B1(n6062), .B2(n6070), .A(n6061), .ZN(n6077) );
  OAI221_X1 U7148 ( .B1(n6071), .B2(n6064), .C1(n6071), .C2(n6063), .A(n6077), 
        .ZN(n6065) );
  AOI22_X1 U7149 ( .A1(n6066), .A2(n6434), .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n6065), .ZN(n6067) );
  OAI211_X1 U7150 ( .C1(n6070), .C2(n6069), .A(n6068), .B(n6067), .ZN(U3004)
         );
  NOR2_X1 U7151 ( .A1(n6372), .A2(n6071), .ZN(n6073) );
  OAI22_X1 U7152 ( .A1(n6149), .A2(n6428), .B1(n6631), .B2(n6426), .ZN(n6072)
         );
  AOI211_X1 U7153 ( .C1(n6074), .C2(n6434), .A(n6073), .B(n6072), .ZN(n6075)
         );
  OAI21_X1 U7154 ( .B1(n6077), .B2(n6076), .A(n6075), .ZN(U3005) );
  INV_X1 U7155 ( .A(n6078), .ZN(n6081) );
  NAND4_X1 U7156 ( .A1(n6081), .A2(n6080), .A3(n6079), .A4(n6226), .ZN(n6082)
         );
  OAI21_X1 U7157 ( .B1(n6084), .B2(n6083), .A(n6082), .ZN(U3455) );
  INV_X1 U7158 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6781) );
  AOI21_X1 U7159 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6781), .A(n6603), .ZN(n6089) );
  INV_X1 U7160 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6085) );
  NAND2_X1 U7161 ( .A1(n6603), .A2(STATE_REG_1__SCAN_IN), .ZN(n6697) );
  INV_X1 U7162 ( .A(n6697), .ZN(n6657) );
  AOI21_X1 U7163 ( .B1(n6089), .B2(n6085), .A(n6657), .ZN(U2789) );
  OAI21_X1 U7164 ( .B1(n6086), .B2(n6587), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6087) );
  OAI21_X1 U7165 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6588), .A(n6087), .ZN(
        U2790) );
  INV_X1 U7166 ( .A(n6657), .ZN(n6684) );
  NOR2_X1 U7167 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6090) );
  OAI21_X1 U7168 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6090), .A(n6697), .ZN(n6088)
         );
  OAI21_X1 U7169 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6684), .A(n6088), .ZN(
        U2791) );
  NOR2_X1 U7170 ( .A1(n6657), .A2(n6089), .ZN(n6663) );
  OAI21_X1 U7171 ( .B1(BS16_N), .B2(n6090), .A(n6663), .ZN(n6661) );
  OAI21_X1 U7172 ( .B1(n6663), .B2(n6091), .A(n6661), .ZN(U2792) );
  AOI21_X1 U7173 ( .B1(n6092), .B2(FLUSH_REG_SCAN_IN), .A(n6358), .ZN(n6093)
         );
  INV_X1 U7174 ( .A(n6093), .ZN(U2793) );
  NOR4_X1 U7175 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n6097) );
  NOR4_X1 U7176 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6096) );
  NOR4_X1 U7177 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_27__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6095) );
  NOR4_X1 U7178 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n6094) );
  NAND4_X1 U7179 ( .A1(n6097), .A2(n6096), .A3(n6095), .A4(n6094), .ZN(n6103)
         );
  NOR4_X1 U7180 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6101) );
  AOI211_X1 U7181 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_19__SCAN_IN), .B(
        DATAWIDTH_REG_28__SCAN_IN), .ZN(n6100) );
  NOR4_X1 U7182 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_10__SCAN_IN), .ZN(
        n6099) );
  NOR4_X1 U7183 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), .A3(DATAWIDTH_REG_4__SCAN_IN), .A4(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6098) );
  NAND4_X1 U7184 ( .A1(n6101), .A2(n6100), .A3(n6099), .A4(n6098), .ZN(n6102)
         );
  NOR2_X1 U7185 ( .A1(n6103), .A2(n6102), .ZN(n6680) );
  INV_X1 U7186 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6105) );
  NOR3_X1 U7187 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6106) );
  OAI21_X1 U7188 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6106), .A(n6680), .ZN(n6104)
         );
  OAI21_X1 U7189 ( .B1(n6680), .B2(n6105), .A(n6104), .ZN(U2794) );
  INV_X1 U7190 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6662) );
  AOI21_X1 U7191 ( .B1(n6676), .B2(n6662), .A(n6106), .ZN(n6108) );
  INV_X1 U7192 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6107) );
  INV_X1 U7193 ( .A(n6680), .ZN(n6682) );
  AOI22_X1 U7194 ( .A1(n6680), .A2(n6108), .B1(n6107), .B2(n6682), .ZN(U2795)
         );
  NAND2_X1 U7195 ( .A1(n6110), .A2(n6109), .ZN(n6119) );
  AOI22_X1 U7196 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6231), .B1(n6111), .B2(n6113), .ZN(n6112) );
  OAI21_X1 U7197 ( .B1(n6113), .B2(n6119), .A(n6112), .ZN(n6114) );
  AOI211_X1 U7198 ( .C1(n6235), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6207), 
        .B(n6114), .ZN(n6117) );
  AOI22_X1 U7199 ( .A1(n6244), .A2(n6190), .B1(n5994), .B2(n6115), .ZN(n6116)
         );
  OAI211_X1 U7200 ( .C1(n6243), .C2(n6118), .A(n6117), .B(n6116), .ZN(U2809)
         );
  AOI21_X1 U7201 ( .B1(n6917), .B2(n6120), .A(n6119), .ZN(n6123) );
  AOI22_X1 U7202 ( .A1(EBX_REG_17__SCAN_IN), .A2(n6231), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6235), .ZN(n6121) );
  INV_X1 U7203 ( .A(n6121), .ZN(n6122) );
  NOR3_X1 U7204 ( .A1(n6207), .A2(n6123), .A3(n6122), .ZN(n6126) );
  AOI22_X1 U7205 ( .A1(n6249), .A2(n6190), .B1(n6214), .B2(n6124), .ZN(n6125)
         );
  OAI211_X1 U7206 ( .C1(n6127), .C2(n6238), .A(n6126), .B(n6125), .ZN(U2810)
         );
  AOI21_X1 U7207 ( .B1(n6235), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6207), 
        .ZN(n6137) );
  AOI22_X1 U7208 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6231), .B1(
        REIP_REG_16__SCAN_IN), .B2(n6142), .ZN(n6136) );
  OAI22_X1 U7209 ( .A1(n6129), .A2(n6199), .B1(n6243), .B2(n6128), .ZN(n6130)
         );
  AOI21_X1 U7210 ( .B1(n6131), .B2(n5994), .A(n6130), .ZN(n6135) );
  NOR2_X1 U7211 ( .A1(n6633), .A2(n6132), .ZN(n6138) );
  OAI211_X1 U7212 ( .C1(REIP_REG_16__SCAN_IN), .C2(REIP_REG_15__SCAN_IN), .A(
        n6138), .B(n6133), .ZN(n6134) );
  NAND4_X1 U7213 ( .A1(n6137), .A2(n6136), .A3(n6135), .A4(n6134), .ZN(U2811)
         );
  AOI22_X1 U7214 ( .A1(n6214), .A2(n6139), .B1(n6138), .B2(n5499), .ZN(n6148)
         );
  INV_X1 U7215 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6946) );
  OAI22_X1 U7216 ( .A1(n6140), .A2(n6175), .B1(n6946), .B2(n6220), .ZN(n6141)
         );
  AOI211_X1 U7217 ( .C1(REIP_REG_15__SCAN_IN), .C2(n6142), .A(n6207), .B(n6141), .ZN(n6147) );
  INV_X1 U7218 ( .A(n6143), .ZN(n6144) );
  AOI22_X1 U7219 ( .A1(n6145), .A2(n6190), .B1(n5994), .B2(n6144), .ZN(n6146)
         );
  NAND3_X1 U7220 ( .A1(n6148), .A2(n6147), .A3(n6146), .ZN(U2812) );
  OAI22_X1 U7221 ( .A1(n6150), .A2(n6175), .B1(n6243), .B2(n6149), .ZN(n6151)
         );
  AOI211_X1 U7222 ( .C1(n6235), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6207), 
        .B(n6151), .ZN(n6160) );
  AOI22_X1 U7223 ( .A1(n6153), .A2(n6190), .B1(n5994), .B2(n6152), .ZN(n6159)
         );
  OAI21_X1 U7224 ( .B1(n6155), .B2(n6154), .A(REIP_REG_13__SCAN_IN), .ZN(n6158) );
  NAND3_X1 U7225 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6156), .A3(n6631), .ZN(
        n6157) );
  NAND4_X1 U7226 ( .A1(n6160), .A2(n6159), .A3(n6158), .A4(n6157), .ZN(U2814)
         );
  AOI22_X1 U7227 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6231), .B1(n6214), .B2(n6161), 
        .ZN(n6162) );
  OAI211_X1 U7228 ( .C1(n6220), .C2(n6163), .A(n6162), .B(n6218), .ZN(n6164)
         );
  NOR2_X1 U7229 ( .A1(n6165), .A2(n6164), .ZN(n6166) );
  OAI21_X1 U7230 ( .B1(n6167), .B2(n6199), .A(n6166), .ZN(n6168) );
  INV_X1 U7231 ( .A(n6168), .ZN(n6172) );
  AOI22_X1 U7232 ( .A1(n6170), .A2(n5994), .B1(REIP_REG_9__SCAN_IN), .B2(n6169), .ZN(n6171) );
  NAND2_X1 U7233 ( .A1(n6172), .A2(n6171), .ZN(U2818) );
  AOI21_X1 U7234 ( .B1(n6216), .B2(n6173), .A(REIP_REG_8__SCAN_IN), .ZN(n6184)
         );
  OAI22_X1 U7235 ( .A1(n6176), .A2(n6175), .B1(n6243), .B2(n6174), .ZN(n6177)
         );
  AOI211_X1 U7236 ( .C1(n6235), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6207), 
        .B(n6177), .ZN(n6182) );
  INV_X1 U7237 ( .A(n6178), .ZN(n6179) );
  AOI22_X1 U7238 ( .A1(n6180), .A2(n6190), .B1(n5994), .B2(n6179), .ZN(n6181)
         );
  OAI211_X1 U7239 ( .C1(n6184), .C2(n6183), .A(n6182), .B(n6181), .ZN(U2819)
         );
  NOR3_X1 U7240 ( .A1(n6209), .A2(REIP_REG_7__SCAN_IN), .A3(n6185), .ZN(n6189)
         );
  INV_X1 U7241 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6330) );
  AOI22_X1 U7242 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6231), .B1(n6214), .B2(n6186), 
        .ZN(n6187) );
  OAI211_X1 U7243 ( .C1(n6220), .C2(n6330), .A(n6187), .B(n6218), .ZN(n6188)
         );
  AOI211_X1 U7244 ( .C1(n6326), .C2(n6190), .A(n6189), .B(n6188), .ZN(n6194)
         );
  OAI21_X1 U7245 ( .B1(n6209), .B2(n6192), .A(n6191), .ZN(n6211) );
  AND3_X1 U7246 ( .A1(n6216), .A2(n6192), .A3(n6621), .ZN(n6197) );
  OAI21_X1 U7247 ( .B1(n6211), .B2(n6197), .A(REIP_REG_7__SCAN_IN), .ZN(n6193)
         );
  OAI211_X1 U7248 ( .C1(n6238), .C2(n6324), .A(n6194), .B(n6193), .ZN(U2820)
         );
  OAI21_X1 U7249 ( .B1(n6220), .B2(n6195), .A(n6218), .ZN(n6196) );
  AOI211_X1 U7250 ( .C1(n6231), .C2(EBX_REG_6__SCAN_IN), .A(n6197), .B(n6196), 
        .ZN(n6203) );
  OAI22_X1 U7251 ( .A1(n6200), .A2(n6199), .B1(n6198), .B2(n6238), .ZN(n6201)
         );
  AOI21_X1 U7252 ( .B1(REIP_REG_6__SCAN_IN), .B2(n6211), .A(n6201), .ZN(n6202)
         );
  OAI211_X1 U7253 ( .C1(n6243), .C2(n6204), .A(n6203), .B(n6202), .ZN(U2821)
         );
  INV_X1 U7254 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6340) );
  OAI22_X1 U7255 ( .A1(n6340), .A2(n6220), .B1(n6243), .B2(n6205), .ZN(n6206)
         );
  AOI211_X1 U7256 ( .C1(n6231), .C2(EBX_REG_5__SCAN_IN), .A(n6207), .B(n6206), 
        .ZN(n6213) );
  OAI21_X1 U7257 ( .B1(n6209), .B2(n6208), .A(n6619), .ZN(n6210) );
  AOI22_X1 U7258 ( .A1(n6334), .A2(n6240), .B1(n6211), .B2(n6210), .ZN(n6212)
         );
  OAI211_X1 U7259 ( .C1(n6331), .C2(n6238), .A(n6213), .B(n6212), .ZN(U2822)
         );
  AOI22_X1 U7260 ( .A1(EBX_REG_4__SCAN_IN), .A2(n6231), .B1(n6214), .B2(n6396), 
        .ZN(n6228) );
  INV_X1 U7261 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6219) );
  NAND3_X1 U7262 ( .A1(n6216), .A2(n6617), .A3(n6215), .ZN(n6217) );
  OAI211_X1 U7263 ( .C1(n6220), .C2(n6219), .A(n6218), .B(n6217), .ZN(n6225)
         );
  OAI22_X1 U7264 ( .A1(n6223), .A2(n6222), .B1(n6221), .B2(n6238), .ZN(n6224)
         );
  AOI211_X1 U7265 ( .C1(n6226), .C2(n6232), .A(n6225), .B(n6224), .ZN(n6227)
         );
  OAI211_X1 U7266 ( .C1(n6617), .C2(n6229), .A(n6228), .B(n6227), .ZN(U2823)
         );
  INV_X1 U7267 ( .A(n6230), .ZN(n6352) );
  AOI22_X1 U7268 ( .A1(n6233), .A2(n6232), .B1(n6231), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n6237) );
  AOI22_X1 U7269 ( .A1(n6235), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6234), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n6236) );
  OAI211_X1 U7270 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6238), .A(n6237), 
        .B(n6236), .ZN(n6239) );
  AOI21_X1 U7271 ( .B1(n6352), .B2(n6240), .A(n6239), .ZN(n6242) );
  OAI211_X1 U7272 ( .C1(n6427), .C2(n6243), .A(n6242), .B(n6241), .ZN(U2826)
         );
  AOI22_X1 U7273 ( .A1(n6244), .A2(n6248), .B1(n6247), .B2(DATAI_18_), .ZN(
        n6246) );
  AOI22_X1 U7274 ( .A1(n6251), .A2(DATAI_2_), .B1(n6250), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7275 ( .A1(n6246), .A2(n6245), .ZN(U2873) );
  AOI22_X1 U7276 ( .A1(n6249), .A2(n6248), .B1(n6247), .B2(DATAI_17_), .ZN(
        n6253) );
  AOI22_X1 U7277 ( .A1(n6251), .A2(DATAI_1_), .B1(n6250), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U7278 ( .A1(n6253), .A2(n6252), .ZN(U2874) );
  INV_X1 U7279 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n6924) );
  INV_X1 U7280 ( .A(n6254), .ZN(n6255) );
  AOI22_X1 U7281 ( .A1(n6283), .A2(DATAO_REG_24__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n6255), .ZN(n6256) );
  OAI21_X1 U7282 ( .B1(n6573), .B2(n6924), .A(n6256), .ZN(U2899) );
  AOI22_X1 U7283 ( .A1(n6689), .A2(LWORD_REG_15__SCAN_IN), .B1(
        DATAO_REG_15__SCAN_IN), .B2(n6283), .ZN(n6257) );
  OAI21_X1 U7284 ( .B1(n3318), .B2(n6285), .A(n6257), .ZN(U2908) );
  INV_X1 U7285 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6811) );
  AOI22_X1 U7286 ( .A1(n6689), .A2(LWORD_REG_14__SCAN_IN), .B1(n6280), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6258) );
  OAI21_X1 U7287 ( .B1(n6811), .B2(n6285), .A(n6258), .ZN(U2909) );
  AOI22_X1 U7288 ( .A1(n6689), .A2(LWORD_REG_13__SCAN_IN), .B1(n6280), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6259) );
  OAI21_X1 U7289 ( .B1(n4926), .B2(n6285), .A(n6259), .ZN(U2910) );
  AOI22_X1 U7290 ( .A1(n6689), .A2(LWORD_REG_12__SCAN_IN), .B1(n6280), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6260) );
  OAI21_X1 U7291 ( .B1(n5110), .B2(n6285), .A(n6260), .ZN(U2911) );
  INV_X1 U7292 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6262) );
  AOI22_X1 U7293 ( .A1(n6277), .A2(LWORD_REG_11__SCAN_IN), .B1(
        DATAO_REG_11__SCAN_IN), .B2(n6283), .ZN(n6261) );
  OAI21_X1 U7294 ( .B1(n6262), .B2(n6285), .A(n6261), .ZN(U2912) );
  INV_X1 U7295 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6264) );
  AOI22_X1 U7296 ( .A1(n6277), .A2(LWORD_REG_10__SCAN_IN), .B1(n6280), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6263) );
  OAI21_X1 U7297 ( .B1(n6264), .B2(n6285), .A(n6263), .ZN(U2913) );
  INV_X1 U7298 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6266) );
  AOI22_X1 U7299 ( .A1(n6277), .A2(LWORD_REG_9__SCAN_IN), .B1(n6280), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6265) );
  OAI21_X1 U7300 ( .B1(n6266), .B2(n6285), .A(n6265), .ZN(U2914) );
  INV_X1 U7301 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6268) );
  AOI22_X1 U7302 ( .A1(n6277), .A2(LWORD_REG_8__SCAN_IN), .B1(
        DATAO_REG_8__SCAN_IN), .B2(n6283), .ZN(n6267) );
  OAI21_X1 U7303 ( .B1(n6268), .B2(n6285), .A(n6267), .ZN(U2915) );
  AOI22_X1 U7304 ( .A1(n6277), .A2(LWORD_REG_7__SCAN_IN), .B1(
        DATAO_REG_7__SCAN_IN), .B2(n6283), .ZN(n6269) );
  OAI21_X1 U7305 ( .B1(n4873), .B2(n6285), .A(n6269), .ZN(U2916) );
  AOI22_X1 U7306 ( .A1(n6277), .A2(LWORD_REG_6__SCAN_IN), .B1(n6280), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6270) );
  OAI21_X1 U7307 ( .B1(n4228), .B2(n6285), .A(n6270), .ZN(U2917) );
  INV_X1 U7308 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6272) );
  AOI22_X1 U7309 ( .A1(n6277), .A2(LWORD_REG_5__SCAN_IN), .B1(
        DATAO_REG_5__SCAN_IN), .B2(n6283), .ZN(n6271) );
  OAI21_X1 U7310 ( .B1(n6272), .B2(n6285), .A(n6271), .ZN(U2918) );
  AOI22_X1 U7311 ( .A1(n6277), .A2(LWORD_REG_4__SCAN_IN), .B1(n6280), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6273) );
  OAI21_X1 U7312 ( .B1(n6274), .B2(n6285), .A(n6273), .ZN(U2919) );
  AOI22_X1 U7313 ( .A1(n6277), .A2(LWORD_REG_3__SCAN_IN), .B1(
        DATAO_REG_3__SCAN_IN), .B2(n6283), .ZN(n6275) );
  OAI21_X1 U7314 ( .B1(n6276), .B2(n6285), .A(n6275), .ZN(U2920) );
  AOI22_X1 U7315 ( .A1(n6277), .A2(LWORD_REG_2__SCAN_IN), .B1(
        DATAO_REG_2__SCAN_IN), .B2(n6283), .ZN(n6278) );
  OAI21_X1 U7316 ( .B1(n6279), .B2(n6285), .A(n6278), .ZN(U2921) );
  AOI22_X1 U7317 ( .A1(n6689), .A2(LWORD_REG_1__SCAN_IN), .B1(n6280), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6281) );
  OAI21_X1 U7318 ( .B1(n6282), .B2(n6285), .A(n6281), .ZN(U2922) );
  AOI22_X1 U7319 ( .A1(n6689), .A2(LWORD_REG_0__SCAN_IN), .B1(n6283), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6284) );
  OAI21_X1 U7320 ( .B1(n6938), .B2(n6285), .A(n6284), .ZN(U2923) );
  INV_X1 U7321 ( .A(DATAI_9_), .ZN(n6286) );
  OR2_X1 U7322 ( .A1(n6298), .A2(n6286), .ZN(n6301) );
  NAND2_X1 U7323 ( .A1(n6699), .A2(UWORD_REG_9__SCAN_IN), .ZN(n6287) );
  AND2_X1 U7324 ( .A1(n6301), .A2(n6287), .ZN(n6288) );
  OAI21_X1 U7325 ( .B1(n6289), .B2(n6313), .A(n6288), .ZN(U2933) );
  INV_X1 U7326 ( .A(DATAI_10_), .ZN(n6290) );
  OR2_X1 U7327 ( .A1(n6298), .A2(n6290), .ZN(n6303) );
  NAND2_X1 U7328 ( .A1(n6699), .A2(UWORD_REG_10__SCAN_IN), .ZN(n6291) );
  AND2_X1 U7329 ( .A1(n6303), .A2(n6291), .ZN(n6292) );
  OAI21_X1 U7330 ( .B1(n6810), .B2(n6313), .A(n6292), .ZN(U2934) );
  OR2_X1 U7331 ( .A1(n6298), .A2(n6293), .ZN(n6308) );
  NAND2_X1 U7332 ( .A1(n6699), .A2(UWORD_REG_12__SCAN_IN), .ZN(n6294) );
  AND2_X1 U7333 ( .A1(n6308), .A2(n6294), .ZN(n6295) );
  OAI21_X1 U7334 ( .B1(n6296), .B2(n6313), .A(n6295), .ZN(U2936) );
  INV_X1 U7335 ( .A(DATAI_14_), .ZN(n6297) );
  OR2_X1 U7336 ( .A1(n6298), .A2(n6297), .ZN(n6311) );
  NAND2_X1 U7337 ( .A1(n6699), .A2(UWORD_REG_14__SCAN_IN), .ZN(n6299) );
  AND2_X1 U7338 ( .A1(n6311), .A2(n6299), .ZN(n6300) );
  OAI21_X1 U7339 ( .B1(n6937), .B2(n6313), .A(n6300), .ZN(U2938) );
  AOI22_X1 U7340 ( .A1(n6699), .A2(LWORD_REG_9__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U7341 ( .A1(n6302), .A2(n6301), .ZN(U2948) );
  AOI22_X1 U7342 ( .A1(n6699), .A2(LWORD_REG_10__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n6304) );
  NAND2_X1 U7343 ( .A1(n6304), .A2(n6303), .ZN(U2949) );
  AOI22_X1 U7344 ( .A1(n6699), .A2(LWORD_REG_11__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U7345 ( .A1(n6305), .A2(DATAI_11_), .ZN(n6701) );
  NAND2_X1 U7346 ( .A1(n6306), .A2(n6701), .ZN(U2950) );
  NAND2_X1 U7347 ( .A1(n6699), .A2(LWORD_REG_12__SCAN_IN), .ZN(n6307) );
  AND2_X1 U7348 ( .A1(n6308), .A2(n6307), .ZN(n6309) );
  OAI21_X1 U7349 ( .B1(n5110), .B2(n6313), .A(n6309), .ZN(U2951) );
  NAND2_X1 U7350 ( .A1(n6699), .A2(LWORD_REG_14__SCAN_IN), .ZN(n6310) );
  AND2_X1 U7351 ( .A1(n6311), .A2(n6310), .ZN(n6312) );
  OAI21_X1 U7352 ( .B1(n6811), .B2(n6313), .A(n6312), .ZN(U2953) );
  AND2_X1 U7353 ( .A1(n6315), .A2(n6314), .ZN(n6316) );
  XNOR2_X1 U7354 ( .A(n6317), .B(n6316), .ZN(n6367) );
  AOI22_X1 U7355 ( .A1(n6379), .A2(REIP_REG_11__SCAN_IN), .B1(n6363), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6322) );
  NOR2_X1 U7356 ( .A1(n6355), .A2(n6318), .ZN(n6319) );
  AOI21_X1 U7357 ( .B1(n6320), .B2(n6360), .A(n6319), .ZN(n6321) );
  OAI211_X1 U7358 ( .C1(n6367), .C2(n6323), .A(n6322), .B(n6321), .ZN(U2975)
         );
  INV_X1 U7359 ( .A(n6324), .ZN(n6325) );
  AOI222_X1 U7360 ( .A1(n6327), .A2(n6358), .B1(n6326), .B2(n6360), .C1(n6325), 
        .C2(n6332), .ZN(n6329) );
  OAI211_X1 U7361 ( .C1(n6330), .C2(n6339), .A(n6329), .B(n6328), .ZN(U2979)
         );
  INV_X1 U7362 ( .A(n6331), .ZN(n6333) );
  AOI222_X1 U7363 ( .A1(n6335), .A2(n6358), .B1(n6360), .B2(n6334), .C1(n6333), 
        .C2(n6332), .ZN(n6338) );
  INV_X1 U7364 ( .A(n6336), .ZN(n6337) );
  OAI211_X1 U7365 ( .C1(n6340), .C2(n6339), .A(n6338), .B(n6337), .ZN(U2981)
         );
  AOI22_X1 U7366 ( .A1(n6379), .A2(REIP_REG_2__SCAN_IN), .B1(n6363), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6346) );
  XNOR2_X1 U7367 ( .A(n6341), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6343)
         );
  XNOR2_X1 U7368 ( .A(n6343), .B(n6342), .ZN(n6422) );
  AOI22_X1 U7369 ( .A1(n6422), .A2(n6358), .B1(n6344), .B2(n6360), .ZN(n6345)
         );
  OAI211_X1 U7370 ( .C1(n6355), .C2(n6347), .A(n6346), .B(n6345), .ZN(U2984)
         );
  AOI22_X1 U7371 ( .A1(n6379), .A2(REIP_REG_1__SCAN_IN), .B1(n6363), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6354) );
  OAI21_X1 U7372 ( .B1(n6350), .B2(n6349), .A(n6348), .ZN(n6351) );
  INV_X1 U7373 ( .A(n6351), .ZN(n6435) );
  AOI22_X1 U7374 ( .A1(n6360), .A2(n6352), .B1(n6435), .B2(n6358), .ZN(n6353)
         );
  OAI211_X1 U7375 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6355), .A(n6354), 
        .B(n6353), .ZN(U2985) );
  INV_X1 U7376 ( .A(n6356), .ZN(n6361) );
  INV_X1 U7377 ( .A(n6357), .ZN(n6359) );
  AOI22_X1 U7378 ( .A1(n6361), .A2(n6360), .B1(n6359), .B2(n6358), .ZN(n6366)
         );
  OAI21_X1 U7379 ( .B1(n6363), .B2(n6362), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6364) );
  NAND3_X1 U7380 ( .A1(n6366), .A2(n6365), .A3(n6364), .ZN(U2986) );
  INV_X1 U7381 ( .A(n6367), .ZN(n6369) );
  AOI222_X1 U7382 ( .A1(n6369), .A2(n6434), .B1(n6405), .B2(n6368), .C1(
        REIP_REG_11__SCAN_IN), .C2(n6379), .ZN(n6370) );
  OAI221_X1 U7383 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6372), .C1(
        n6861), .C2(n6371), .A(n6370), .ZN(U3007) );
  AOI21_X1 U7384 ( .B1(n6375), .B2(n6374), .A(n6373), .ZN(n6393) );
  NAND2_X1 U7385 ( .A1(n6377), .A2(n6376), .ZN(n6386) );
  AOI221_X1 U7386 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n6392), .C2(n6385), .A(n6386), 
        .ZN(n6378) );
  AOI21_X1 U7387 ( .B1(n6379), .B2(REIP_REG_10__SCAN_IN), .A(n6378), .ZN(n6380) );
  OAI21_X1 U7388 ( .B1(n6381), .B2(n6428), .A(n6380), .ZN(n6382) );
  AOI21_X1 U7389 ( .B1(n6383), .B2(n6434), .A(n6382), .ZN(n6384) );
  OAI21_X1 U7390 ( .B1(n6393), .B2(n6385), .A(n6384), .ZN(U3008) );
  NOR2_X1 U7391 ( .A1(n6386), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6389)
         );
  OAI22_X1 U7392 ( .A1(n6387), .A2(n6428), .B1(n5368), .B2(n6426), .ZN(n6388)
         );
  AOI211_X1 U7393 ( .C1(n6390), .C2(n6434), .A(n6389), .B(n6388), .ZN(n6391)
         );
  OAI21_X1 U7394 ( .B1(n6393), .B2(n6392), .A(n6391), .ZN(U3009) );
  OAI21_X1 U7395 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6394), .ZN(n6402) );
  AOI21_X1 U7396 ( .B1(n6405), .B2(n6396), .A(n6395), .ZN(n6399) );
  OR2_X1 U7397 ( .A1(n6397), .A2(n6406), .ZN(n6398) );
  OAI211_X1 U7398 ( .C1(n6414), .C2(n4007), .A(n6399), .B(n6398), .ZN(n6400)
         );
  INV_X1 U7399 ( .A(n6400), .ZN(n6401) );
  OAI21_X1 U7400 ( .B1(n6410), .B2(n6402), .A(n6401), .ZN(U3014) );
  INV_X1 U7401 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6413) );
  NOR2_X1 U7402 ( .A1(n6426), .A2(n5480), .ZN(n6403) );
  AOI21_X1 U7403 ( .B1(n6405), .B2(n6404), .A(n6403), .ZN(n6409) );
  OR2_X1 U7404 ( .A1(n6407), .A2(n6406), .ZN(n6408) );
  OAI211_X1 U7405 ( .C1(n6410), .C2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6409), 
        .B(n6408), .ZN(n6411) );
  INV_X1 U7406 ( .A(n6411), .ZN(n6412) );
  OAI21_X1 U7407 ( .B1(n6414), .B2(n6413), .A(n6412), .ZN(U3015) );
  NAND2_X1 U7408 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6415), .ZN(n6425)
         );
  NAND3_X1 U7409 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A3(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6417) );
  AOI21_X1 U7410 ( .B1(n6418), .B2(n6417), .A(n6416), .ZN(n6421) );
  OAI22_X1 U7411 ( .A1(n6428), .A2(n6419), .B1(n6614), .B2(n6426), .ZN(n6420)
         );
  AOI211_X1 U7412 ( .C1(n6422), .C2(n6434), .A(n6421), .B(n6420), .ZN(n6423)
         );
  OAI221_X1 U7413 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6425), .C1(n3867), .C2(n6424), .A(n6423), .ZN(U3016) );
  OAI22_X1 U7414 ( .A1(n6428), .A2(n6427), .B1(n6676), .B2(n6426), .ZN(n6433)
         );
  AOI211_X1 U7415 ( .C1(n6431), .C2(n6430), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .B(n6429), .ZN(n6432) );
  AOI211_X1 U7416 ( .C1(n6435), .C2(n6434), .A(n6433), .B(n6432), .ZN(n6436)
         );
  OAI21_X1 U7417 ( .B1(n6437), .B2(n3858), .A(n6436), .ZN(U3017) );
  NOR2_X1 U7418 ( .A1(n6438), .A2(n6675), .ZN(U3019) );
  INV_X1 U7419 ( .A(n6439), .ZN(n6479) );
  INV_X1 U7420 ( .A(n6484), .ZN(n6472) );
  AOI22_X1 U7421 ( .A1(n6488), .A2(n6479), .B1(n6440), .B2(n6472), .ZN(n6451)
         );
  NAND2_X1 U7422 ( .A1(n6441), .A2(n6445), .ZN(n6449) );
  INV_X1 U7423 ( .A(n6449), .ZN(n6443) );
  AOI21_X1 U7424 ( .B1(n6442), .B2(n3110), .A(n6479), .ZN(n6448) );
  NAND2_X1 U7425 ( .A1(n6443), .A2(n6448), .ZN(n6444) );
  OAI211_X1 U7426 ( .C1(n6446), .C2(n6445), .A(n6494), .B(n6444), .ZN(n6481)
         );
  OAI22_X1 U7427 ( .A1(n6449), .A2(n6448), .B1(n6447), .B2(n6814), .ZN(n6480)
         );
  AOI22_X1 U7428 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6481), .B1(n6499), 
        .B2(n6480), .ZN(n6450) );
  OAI211_X1 U7429 ( .C1(n6452), .C2(n6475), .A(n6451), .B(n6450), .ZN(U3076)
         );
  AOI22_X1 U7430 ( .A1(n6504), .A2(n6479), .B1(n6472), .B2(n6453), .ZN(n6455)
         );
  AOI22_X1 U7431 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6481), .B1(n6505), 
        .B2(n6480), .ZN(n6454) );
  OAI211_X1 U7432 ( .C1(n6456), .C2(n6475), .A(n6455), .B(n6454), .ZN(U3077)
         );
  AOI22_X1 U7433 ( .A1(n6510), .A2(n6479), .B1(n6472), .B2(n6509), .ZN(n6458)
         );
  AOI22_X1 U7434 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6481), .B1(n6511), 
        .B2(n6480), .ZN(n6457) );
  OAI211_X1 U7435 ( .C1(n6514), .C2(n6475), .A(n6458), .B(n6457), .ZN(U3078)
         );
  INV_X1 U7436 ( .A(n6475), .ZN(n6477) );
  AOI22_X1 U7437 ( .A1(n6516), .A2(n6479), .B1(n6459), .B2(n6477), .ZN(n6461)
         );
  AOI22_X1 U7438 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6481), .B1(n6517), 
        .B2(n6480), .ZN(n6460) );
  OAI211_X1 U7439 ( .C1(n6462), .C2(n6484), .A(n6461), .B(n6460), .ZN(U3079)
         );
  AOI22_X1 U7440 ( .A1(n6522), .A2(n6479), .B1(n6463), .B2(n6477), .ZN(n6465)
         );
  AOI22_X1 U7441 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6481), .B1(n6523), 
        .B2(n6480), .ZN(n6464) );
  OAI211_X1 U7442 ( .C1(n6466), .C2(n6484), .A(n6465), .B(n6464), .ZN(U3080)
         );
  AOI22_X1 U7443 ( .A1(n6528), .A2(n6479), .B1(n6467), .B2(n6477), .ZN(n6469)
         );
  AOI22_X1 U7444 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6481), .B1(n6529), 
        .B2(n6480), .ZN(n6468) );
  OAI211_X1 U7445 ( .C1(n6470), .C2(n6484), .A(n6469), .B(n6468), .ZN(U3081)
         );
  AOI22_X1 U7446 ( .A1(n6535), .A2(n6479), .B1(n6472), .B2(n6471), .ZN(n6474)
         );
  AOI22_X1 U7447 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6481), .B1(n6536), 
        .B2(n6480), .ZN(n6473) );
  OAI211_X1 U7448 ( .C1(n6476), .C2(n6475), .A(n6474), .B(n6473), .ZN(U3082)
         );
  AOI22_X1 U7449 ( .A1(n6544), .A2(n6479), .B1(n6478), .B2(n6477), .ZN(n6483)
         );
  AOI22_X1 U7450 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6481), .B1(n6546), 
        .B2(n6480), .ZN(n6482) );
  OAI211_X1 U7451 ( .C1(n6485), .C2(n6484), .A(n6483), .B(n6482), .ZN(U3083)
         );
  NOR2_X1 U7452 ( .A1(n6486), .A2(n6674), .ZN(n6543) );
  INV_X1 U7453 ( .A(n6550), .ZN(n6534) );
  AOI22_X1 U7454 ( .A1(n6488), .A2(n6543), .B1(n6534), .B2(n6487), .ZN(n6501)
         );
  AOI21_X1 U7455 ( .B1(n6490), .B2(n6489), .A(n6492), .ZN(n6495) );
  AOI21_X1 U7456 ( .B1(n6491), .B2(n3110), .A(n6543), .ZN(n6497) );
  AOI22_X1 U7457 ( .A1(n6495), .A2(n6497), .B1(n6496), .B2(n6492), .ZN(n6493)
         );
  NAND2_X1 U7458 ( .A1(n6494), .A2(n6493), .ZN(n6547) );
  INV_X1 U7459 ( .A(n6495), .ZN(n6498) );
  OAI22_X1 U7460 ( .A1(n6498), .A2(n6497), .B1(n6496), .B2(n6814), .ZN(n6545)
         );
  AOI22_X1 U7461 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6547), .B1(n6499), 
        .B2(n6545), .ZN(n6500) );
  OAI211_X1 U7462 ( .C1(n6502), .C2(n6539), .A(n6501), .B(n6500), .ZN(U3108)
         );
  AOI22_X1 U7463 ( .A1(n6504), .A2(n6543), .B1(n6534), .B2(n6503), .ZN(n6507)
         );
  AOI22_X1 U7464 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6547), .B1(n6505), 
        .B2(n6545), .ZN(n6506) );
  OAI211_X1 U7465 ( .C1(n6508), .C2(n6539), .A(n6507), .B(n6506), .ZN(U3109)
         );
  AOI22_X1 U7466 ( .A1(n6510), .A2(n6543), .B1(n6542), .B2(n6509), .ZN(n6513)
         );
  AOI22_X1 U7467 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6547), .B1(n6511), 
        .B2(n6545), .ZN(n6512) );
  OAI211_X1 U7468 ( .C1(n6514), .C2(n6550), .A(n6513), .B(n6512), .ZN(U3110)
         );
  AOI22_X1 U7469 ( .A1(n6516), .A2(n6543), .B1(n6542), .B2(n6515), .ZN(n6519)
         );
  AOI22_X1 U7470 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6547), .B1(n6517), 
        .B2(n6545), .ZN(n6518) );
  OAI211_X1 U7471 ( .C1(n6520), .C2(n6550), .A(n6519), .B(n6518), .ZN(U3111)
         );
  AOI22_X1 U7472 ( .A1(n6522), .A2(n6543), .B1(n6542), .B2(n6521), .ZN(n6525)
         );
  AOI22_X1 U7473 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6547), .B1(n6523), 
        .B2(n6545), .ZN(n6524) );
  OAI211_X1 U7474 ( .C1(n6526), .C2(n6550), .A(n6525), .B(n6524), .ZN(U3112)
         );
  AOI22_X1 U7475 ( .A1(n6528), .A2(n6543), .B1(n6542), .B2(n6527), .ZN(n6531)
         );
  AOI22_X1 U7476 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6547), .B1(n6529), 
        .B2(n6545), .ZN(n6530) );
  OAI211_X1 U7477 ( .C1(n6532), .C2(n6550), .A(n6531), .B(n6530), .ZN(U3113)
         );
  AOI22_X1 U7478 ( .A1(n6535), .A2(n6543), .B1(n6534), .B2(n6533), .ZN(n6538)
         );
  AOI22_X1 U7479 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6547), .B1(n6536), 
        .B2(n6545), .ZN(n6537) );
  OAI211_X1 U7480 ( .C1(n6540), .C2(n6539), .A(n6538), .B(n6537), .ZN(U3114)
         );
  AOI22_X1 U7481 ( .A1(n6544), .A2(n6543), .B1(n6542), .B2(n6541), .ZN(n6549)
         );
  AOI22_X1 U7482 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6547), .B1(n6546), 
        .B2(n6545), .ZN(n6548) );
  OAI211_X1 U7483 ( .C1(n6551), .C2(n6550), .A(n6549), .B(n6548), .ZN(U3115)
         );
  AND3_X1 U7484 ( .A1(n6553), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6552), 
        .ZN(n6557) );
  NAND2_X1 U7485 ( .A1(n6555), .A2(n6554), .ZN(n6556) );
  AOI222_X1 U7486 ( .A1(n6557), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n6557), .B2(n6556), .C1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n6556), 
        .ZN(n6558) );
  AOI222_X1 U7487 ( .A1(n6560), .A2(n6559), .B1(n6560), .B2(n6558), .C1(n6559), 
        .C2(n6558), .ZN(n6564) );
  INV_X1 U7488 ( .A(n6564), .ZN(n6562) );
  AOI21_X1 U7489 ( .B1(n6562), .B2(n6674), .A(n6561), .ZN(n6563) );
  AOI211_X1 U7490 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6564), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n6563), .ZN(n6572) );
  OAI21_X1 U7491 ( .B1(MORE_REG_SCAN_IN), .B2(FLUSH_REG_SCAN_IN), .A(n6565), 
        .ZN(n6568) );
  NAND3_X1 U7492 ( .A1(n6568), .A2(n6567), .A3(n6566), .ZN(n6569) );
  NOR4_X1 U7493 ( .A1(n6572), .A2(n6571), .A3(n6570), .A4(n6569), .ZN(n6585)
         );
  INV_X1 U7494 ( .A(n6585), .ZN(n6574) );
  OAI22_X1 U7495 ( .A1(n6574), .A2(n6587), .B1(n6688), .B2(n6573), .ZN(n6575)
         );
  OAI21_X1 U7496 ( .B1(n6577), .B2(n6576), .A(n6575), .ZN(n6665) );
  OAI21_X1 U7497 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6688), .A(n6665), .ZN(
        n6586) );
  AOI221_X1 U7498 ( .B1(n6579), .B2(STATE2_REG_0__SCAN_IN), .C1(n6586), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6578), .ZN(n6584) );
  OAI211_X1 U7499 ( .C1(n6582), .C2(n6581), .A(n6580), .B(n6665), .ZN(n6583)
         );
  OAI211_X1 U7500 ( .C1(n6585), .C2(n6587), .A(n6584), .B(n6583), .ZN(U3148)
         );
  OAI211_X1 U7501 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(STATE2_REG_1__SCAN_IN), .B(n6586), .ZN(n6592) );
  OAI21_X1 U7502 ( .B1(READY_N), .B2(n6588), .A(n6587), .ZN(n6590) );
  AOI21_X1 U7503 ( .B1(n6590), .B2(n6665), .A(n6589), .ZN(n6591) );
  NAND2_X1 U7504 ( .A1(n6592), .A2(n6591), .ZN(U3149) );
  OAI221_X1 U7505 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(n6688), .A(n6664), .ZN(n6594) );
  OAI21_X1 U7506 ( .B1(n6692), .B2(n6594), .A(n6593), .ZN(U3150) );
  INV_X1 U7507 ( .A(n6663), .ZN(n6595) );
  AND2_X1 U7508 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6595), .ZN(U3151) );
  AND2_X1 U7509 ( .A1(n6595), .A2(DATAWIDTH_REG_30__SCAN_IN), .ZN(U3152) );
  AND2_X1 U7510 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6595), .ZN(U3153) );
  INV_X1 U7511 ( .A(DATAWIDTH_REG_28__SCAN_IN), .ZN(n6798) );
  NOR2_X1 U7512 ( .A1(n6663), .A2(n6798), .ZN(U3154) );
  AND2_X1 U7513 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6595), .ZN(U3155) );
  AND2_X1 U7514 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6595), .ZN(U3156) );
  AND2_X1 U7515 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6595), .ZN(U3157) );
  AND2_X1 U7516 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6595), .ZN(U3158) );
  AND2_X1 U7517 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6595), .ZN(U3159) );
  AND2_X1 U7518 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6595), .ZN(U3160) );
  AND2_X1 U7519 ( .A1(n6595), .A2(DATAWIDTH_REG_21__SCAN_IN), .ZN(U3161) );
  AND2_X1 U7520 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6595), .ZN(U3162) );
  AND2_X1 U7521 ( .A1(n6595), .A2(DATAWIDTH_REG_19__SCAN_IN), .ZN(U3163) );
  AND2_X1 U7522 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6595), .ZN(U3164) );
  AND2_X1 U7523 ( .A1(n6595), .A2(DATAWIDTH_REG_17__SCAN_IN), .ZN(U3165) );
  AND2_X1 U7524 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6595), .ZN(U3166) );
  AND2_X1 U7525 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6595), .ZN(U3167) );
  AND2_X1 U7526 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6595), .ZN(U3168) );
  AND2_X1 U7527 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6595), .ZN(U3169) );
  AND2_X1 U7528 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6595), .ZN(U3170) );
  AND2_X1 U7529 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6595), .ZN(U3171) );
  AND2_X1 U7530 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6595), .ZN(U3172) );
  AND2_X1 U7531 ( .A1(n6595), .A2(DATAWIDTH_REG_9__SCAN_IN), .ZN(U3173) );
  AND2_X1 U7532 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6595), .ZN(U3174) );
  AND2_X1 U7533 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6595), .ZN(U3175) );
  AND2_X1 U7534 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6595), .ZN(U3176) );
  AND2_X1 U7535 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6595), .ZN(U3177) );
  AND2_X1 U7536 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6595), .ZN(U3178) );
  INV_X1 U7537 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6986) );
  NOR2_X1 U7538 ( .A1(n6663), .A2(n6986), .ZN(U3179) );
  AND2_X1 U7539 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6595), .ZN(U3180) );
  NOR2_X1 U7540 ( .A1(n6781), .A2(n6602), .ZN(n6605) );
  AOI22_X1 U7541 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6609) );
  AND2_X1 U7542 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6599) );
  INV_X1 U7543 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6597) );
  INV_X1 U7544 ( .A(NA_N), .ZN(n6606) );
  AOI221_X1 U7545 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6606), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6611) );
  AOI221_X1 U7546 ( .B1(n6599), .B2(n6697), .C1(n6597), .C2(n6684), .A(n6611), 
        .ZN(n6596) );
  OAI21_X1 U7547 ( .B1(n6605), .B2(n6609), .A(n6596), .ZN(U3181) );
  NOR2_X1 U7548 ( .A1(n6603), .A2(n6597), .ZN(n6607) );
  NAND2_X1 U7549 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6598) );
  OAI21_X1 U7550 ( .B1(n6607), .B2(n6599), .A(n6598), .ZN(n6600) );
  OAI211_X1 U7551 ( .C1(n6602), .C2(n6688), .A(n6601), .B(n6600), .ZN(U3182)
         );
  AOI221_X1 U7552 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6688), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6604) );
  AOI221_X1 U7553 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6604), .C2(HOLD), .A(n6603), .ZN(n6610) );
  AOI21_X1 U7554 ( .B1(n6607), .B2(n6606), .A(n6605), .ZN(n6608) );
  OAI22_X1 U7555 ( .A1(n6611), .A2(n6610), .B1(n6609), .B2(n6608), .ZN(U3183)
         );
  OR2_X1 U7556 ( .A1(n6697), .A2(STATE_REG_2__SCAN_IN), .ZN(n6651) );
  INV_X1 U7557 ( .A(n6651), .ZN(n6653) );
  NOR2_X2 U7558 ( .A1(n6781), .A2(n6697), .ZN(n6649) );
  AOI222_X1 U7559 ( .A1(n6653), .A2(REIP_REG_2__SCAN_IN), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6684), .C1(REIP_REG_1__SCAN_IN), .C2(
        n6649), .ZN(n6612) );
  INV_X1 U7560 ( .A(n6612), .ZN(U3184) );
  INV_X1 U7561 ( .A(n6649), .ZN(n6655) );
  AOI22_X1 U7562 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6684), .ZN(n6613) );
  OAI21_X1 U7563 ( .B1(n6614), .B2(n6655), .A(n6613), .ZN(U3185) );
  AOI22_X1 U7564 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6697), .ZN(n6615) );
  OAI21_X1 U7565 ( .B1(n5480), .B2(n6655), .A(n6615), .ZN(U3186) );
  AOI22_X1 U7566 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6697), .ZN(n6616) );
  OAI21_X1 U7567 ( .B1(n6617), .B2(n6655), .A(n6616), .ZN(U3187) );
  AOI22_X1 U7568 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6697), .ZN(n6618) );
  OAI21_X1 U7569 ( .B1(n6619), .B2(n6655), .A(n6618), .ZN(U3188) );
  AOI22_X1 U7570 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6697), .ZN(n6620) );
  OAI21_X1 U7571 ( .B1(n6621), .B2(n6655), .A(n6620), .ZN(U3189) );
  AOI22_X1 U7572 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6697), .ZN(n6622) );
  OAI21_X1 U7573 ( .B1(n4796), .B2(n6655), .A(n6622), .ZN(U3190) );
  AOI222_X1 U7574 ( .A1(n6649), .A2(REIP_REG_8__SCAN_IN), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6684), .C1(REIP_REG_9__SCAN_IN), .C2(
        n6653), .ZN(n6623) );
  INV_X1 U7575 ( .A(n6623), .ZN(U3191) );
  AOI222_X1 U7576 ( .A1(n6649), .A2(REIP_REG_9__SCAN_IN), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6684), .C1(REIP_REG_10__SCAN_IN), .C2(
        n6653), .ZN(n6624) );
  INV_X1 U7577 ( .A(n6624), .ZN(U3192) );
  AOI22_X1 U7578 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6697), .ZN(n6625) );
  OAI21_X1 U7579 ( .B1(n6626), .B2(n6655), .A(n6625), .ZN(U3193) );
  AOI22_X1 U7580 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6684), .ZN(n6627) );
  OAI21_X1 U7581 ( .B1(n6628), .B2(n6655), .A(n6627), .ZN(U3194) );
  AOI22_X1 U7582 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6697), .ZN(n6629) );
  OAI21_X1 U7583 ( .B1(n6878), .B2(n6655), .A(n6629), .ZN(U3195) );
  AOI22_X1 U7584 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6684), .ZN(n6630) );
  OAI21_X1 U7585 ( .B1(n6631), .B2(n6655), .A(n6630), .ZN(U3196) );
  AOI22_X1 U7586 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6684), .ZN(n6632) );
  OAI21_X1 U7587 ( .B1(n6633), .B2(n6655), .A(n6632), .ZN(U3197) );
  AOI22_X1 U7588 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6684), .ZN(n6634) );
  OAI21_X1 U7589 ( .B1(n5499), .B2(n6655), .A(n6634), .ZN(U3198) );
  AOI22_X1 U7590 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6649), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6684), .ZN(n6635) );
  OAI21_X1 U7591 ( .B1(n6917), .B2(n6651), .A(n6635), .ZN(U3199) );
  AOI22_X1 U7592 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6684), .ZN(n6636) );
  OAI21_X1 U7593 ( .B1(n6917), .B2(n6655), .A(n6636), .ZN(U3200) );
  AOI222_X1 U7594 ( .A1(n6649), .A2(REIP_REG_18__SCAN_IN), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6684), .C1(REIP_REG_19__SCAN_IN), .C2(
        n6653), .ZN(n6637) );
  INV_X1 U7595 ( .A(n6637), .ZN(U3201) );
  AOI22_X1 U7596 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6684), .ZN(n6638) );
  OAI21_X1 U7597 ( .B1(n6639), .B2(n6655), .A(n6638), .ZN(U3202) );
  AOI22_X1 U7598 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6649), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6697), .ZN(n6640) );
  OAI21_X1 U7599 ( .B1(n6880), .B2(n6651), .A(n6640), .ZN(U3203) );
  AOI222_X1 U7600 ( .A1(n6649), .A2(REIP_REG_21__SCAN_IN), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6684), .C1(REIP_REG_22__SCAN_IN), .C2(
        n6653), .ZN(n6641) );
  INV_X1 U7601 ( .A(n6641), .ZN(U3204) );
  INV_X1 U7602 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6932) );
  AOI22_X1 U7603 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6649), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6684), .ZN(n6642) );
  OAI21_X1 U7604 ( .B1(n6932), .B2(n6651), .A(n6642), .ZN(U3205) );
  AOI22_X1 U7605 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6649), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6684), .ZN(n6643) );
  OAI21_X1 U7606 ( .B1(n6896), .B2(n6651), .A(n6643), .ZN(U3206) );
  AOI222_X1 U7607 ( .A1(n6653), .A2(REIP_REG_25__SCAN_IN), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6684), .C1(REIP_REG_24__SCAN_IN), .C2(
        n6649), .ZN(n6644) );
  INV_X1 U7608 ( .A(n6644), .ZN(U3207) );
  AOI222_X1 U7609 ( .A1(n6649), .A2(REIP_REG_25__SCAN_IN), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6684), .C1(REIP_REG_26__SCAN_IN), .C2(
        n6653), .ZN(n6645) );
  INV_X1 U7610 ( .A(n6645), .ZN(U3208) );
  AOI22_X1 U7611 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6649), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6697), .ZN(n6646) );
  OAI21_X1 U7612 ( .B1(n6647), .B2(n6651), .A(n6646), .ZN(U3209) );
  AOI222_X1 U7613 ( .A1(n6649), .A2(REIP_REG_27__SCAN_IN), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6684), .C1(REIP_REG_28__SCAN_IN), .C2(
        n6653), .ZN(n6648) );
  INV_X1 U7614 ( .A(n6648), .ZN(U3210) );
  AOI22_X1 U7615 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6649), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6684), .ZN(n6650) );
  OAI21_X1 U7616 ( .B1(n6998), .B2(n6651), .A(n6650), .ZN(U3211) );
  AOI22_X1 U7617 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6684), .ZN(n6652) );
  OAI21_X1 U7618 ( .B1(n6998), .B2(n6655), .A(n6652), .ZN(U3212) );
  AOI22_X1 U7619 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6653), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6684), .ZN(n6654) );
  OAI21_X1 U7620 ( .B1(n6656), .B2(n6655), .A(n6654), .ZN(U3213) );
  OAI22_X1 U7621 ( .A1(n6697), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n6657), .ZN(n6658) );
  INV_X1 U7622 ( .A(n6658), .ZN(U3445) );
  MUX2_X1 U7623 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6697), .Z(U3446) );
  OAI22_X1 U7624 ( .A1(n6697), .A2(BYTEENABLE_REG_1__SCAN_IN), .B1(
        BE_N_REG_1__SCAN_IN), .B2(n6657), .ZN(n6659) );
  INV_X1 U7625 ( .A(n6659), .ZN(U3447) );
  MUX2_X1 U7626 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6697), .Z(U3448) );
  OAI21_X1 U7627 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6663), .A(n6661), .ZN(
        n6660) );
  INV_X1 U7628 ( .A(n6660), .ZN(U3451) );
  OAI21_X1 U7629 ( .B1(n6663), .B2(n6662), .A(n6661), .ZN(U3452) );
  OAI221_X1 U7630 ( .B1(n6826), .B2(STATE2_REG_0__SCAN_IN), .C1(n6826), .C2(
        n6665), .A(n6664), .ZN(U3453) );
  NAND2_X1 U7631 ( .A1(n6667), .A2(n6666), .ZN(n6668) );
  OAI211_X1 U7632 ( .C1(n6671), .C2(n6670), .A(n6669), .B(n6668), .ZN(n6672)
         );
  NAND2_X1 U7633 ( .A1(n6675), .A2(n6672), .ZN(n6673) );
  OAI21_X1 U7634 ( .B1(n6675), .B2(n6674), .A(n6673), .ZN(U3462) );
  AOI21_X1 U7635 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6677) );
  AOI22_X1 U7636 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6677), .B2(n6676), .ZN(n6679) );
  INV_X1 U7637 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6678) );
  AOI22_X1 U7638 ( .A1(n6680), .A2(n6679), .B1(n6678), .B2(n6682), .ZN(U3468)
         );
  INV_X1 U7639 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6683) );
  NOR2_X1 U7640 ( .A1(n6682), .A2(REIP_REG_1__SCAN_IN), .ZN(n6681) );
  AOI22_X1 U7641 ( .A1(n6683), .A2(n6682), .B1(n3544), .B2(n6681), .ZN(U3469)
         );
  INV_X1 U7642 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6685) );
  AOI22_X1 U7643 ( .A1(n6657), .A2(READREQUEST_REG_SCAN_IN), .B1(n6685), .B2(
        n6684), .ZN(U3470) );
  AOI211_X1 U7644 ( .C1(n6689), .C2(n6688), .A(n6687), .B(n6686), .ZN(n6696)
         );
  OAI211_X1 U7645 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6691), .A(n6690), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6693) );
  AOI21_X1 U7646 ( .B1(n6693), .B2(STATE2_REG_0__SCAN_IN), .A(n6692), .ZN(
        n6695) );
  NAND2_X1 U7647 ( .A1(n6696), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6694) );
  OAI21_X1 U7648 ( .B1(n6696), .B2(n6695), .A(n6694), .ZN(U3472) );
  MUX2_X1 U7649 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6697), .Z(U3473) );
  AOI22_X1 U7650 ( .A1(n6699), .A2(UWORD_REG_11__SCAN_IN), .B1(n6698), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n6700) );
  NAND2_X1 U7651 ( .A1(n6701), .A2(n6700), .ZN(n7024) );
  INV_X1 U7652 ( .A(keyinput18), .ZN(n6813) );
  NOR4_X1 U7653 ( .A1(keyinput48), .A2(keyinput83), .A3(keyinput1), .A4(
        keyinput8), .ZN(n6702) );
  NAND3_X1 U7654 ( .A1(keyinput112), .A2(keyinput7), .A3(n6702), .ZN(n6713) );
  INV_X1 U7655 ( .A(keyinput69), .ZN(n6704) );
  NAND4_X1 U7656 ( .A1(keyinput124), .A2(keyinput86), .A3(keyinput3), .A4(
        keyinput11), .ZN(n6703) );
  NOR3_X1 U7657 ( .A1(keyinput38), .A2(n6704), .A3(n6703), .ZN(n6711) );
  NOR2_X1 U7658 ( .A1(keyinput30), .A2(keyinput95), .ZN(n6705) );
  NAND3_X1 U7659 ( .A1(keyinput94), .A2(keyinput2), .A3(n6705), .ZN(n6709) );
  NAND4_X1 U7660 ( .A1(keyinput37), .A2(keyinput74), .A3(keyinput22), .A4(
        keyinput17), .ZN(n6708) );
  INV_X1 U7661 ( .A(keyinput65), .ZN(n6817) );
  NAND4_X1 U7662 ( .A1(keyinput52), .A2(keyinput110), .A3(keyinput99), .A4(
        n6817), .ZN(n6707) );
  NAND4_X1 U7663 ( .A1(keyinput44), .A2(keyinput33), .A3(keyinput87), .A4(
        keyinput114), .ZN(n6706) );
  NOR4_X1 U7664 ( .A1(n6709), .A2(n6708), .A3(n6707), .A4(n6706), .ZN(n6710)
         );
  NAND3_X1 U7665 ( .A1(keyinput105), .A2(n6711), .A3(n6710), .ZN(n6712) );
  NOR4_X1 U7666 ( .A1(keyinput51), .A2(n6813), .A3(n6713), .A4(n6712), .ZN(
        n6763) );
  NAND4_X1 U7667 ( .A1(keyinput64), .A2(keyinput60), .A3(keyinput96), .A4(
        keyinput13), .ZN(n6761) );
  INV_X1 U7668 ( .A(keyinput10), .ZN(n6714) );
  NAND4_X1 U7669 ( .A1(keyinput79), .A2(keyinput5), .A3(keyinput90), .A4(n6714), .ZN(n6760) );
  INV_X1 U7670 ( .A(keyinput73), .ZN(n6715) );
  NOR4_X1 U7671 ( .A1(keyinput49), .A2(keyinput111), .A3(keyinput23), .A4(
        n6715), .ZN(n6726) );
  NAND2_X1 U7672 ( .A1(keyinput122), .A2(keyinput77), .ZN(n6716) );
  NOR3_X1 U7673 ( .A1(keyinput118), .A2(keyinput108), .A3(n6716), .ZN(n6725)
         );
  NOR2_X1 U7674 ( .A1(keyinput63), .A2(keyinput82), .ZN(n6717) );
  NAND3_X1 U7675 ( .A1(keyinput28), .A2(keyinput50), .A3(n6717), .ZN(n6723) );
  INV_X1 U7676 ( .A(keyinput67), .ZN(n6718) );
  NAND4_X1 U7677 ( .A1(keyinput115), .A2(keyinput32), .A3(keyinput35), .A4(
        n6718), .ZN(n6722) );
  NAND4_X1 U7678 ( .A1(keyinput66), .A2(keyinput72), .A3(keyinput76), .A4(
        keyinput0), .ZN(n6721) );
  NOR2_X1 U7679 ( .A1(keyinput43), .A2(keyinput46), .ZN(n6719) );
  NAND3_X1 U7680 ( .A1(keyinput15), .A2(keyinput25), .A3(n6719), .ZN(n6720) );
  NOR4_X1 U7681 ( .A1(n6723), .A2(n6722), .A3(n6721), .A4(n6720), .ZN(n6724)
         );
  NAND3_X1 U7682 ( .A1(n6726), .A2(n6725), .A3(n6724), .ZN(n6759) );
  NAND2_X1 U7683 ( .A1(keyinput100), .A2(keyinput120), .ZN(n6727) );
  NOR3_X1 U7684 ( .A1(keyinput59), .A2(keyinput20), .A3(n6727), .ZN(n6729) );
  INV_X1 U7685 ( .A(keyinput109), .ZN(n6728) );
  NAND3_X1 U7686 ( .A1(keyinput75), .A2(n6729), .A3(n6728), .ZN(n6740) );
  NAND4_X1 U7687 ( .A1(keyinput126), .A2(keyinput62), .A3(keyinput61), .A4(
        keyinput45), .ZN(n6730) );
  NOR3_X1 U7688 ( .A1(keyinput41), .A2(keyinput103), .A3(n6730), .ZN(n6738) );
  INV_X1 U7689 ( .A(keyinput12), .ZN(n6916) );
  NAND4_X1 U7690 ( .A1(keyinput54), .A2(keyinput88), .A3(keyinput101), .A4(
        n6916), .ZN(n6735) );
  NOR2_X1 U7691 ( .A1(keyinput80), .A2(keyinput70), .ZN(n6731) );
  NAND3_X1 U7692 ( .A1(keyinput6), .A2(keyinput55), .A3(n6731), .ZN(n6734) );
  INV_X1 U7693 ( .A(keyinput58), .ZN(n6923) );
  NAND4_X1 U7694 ( .A1(keyinput117), .A2(keyinput53), .A3(keyinput47), .A4(
        n6923), .ZN(n6733) );
  NAND4_X1 U7695 ( .A1(keyinput42), .A2(keyinput9), .A3(keyinput21), .A4(
        keyinput113), .ZN(n6732) );
  NOR4_X1 U7696 ( .A1(n6735), .A2(n6734), .A3(n6733), .A4(n6732), .ZN(n6737)
         );
  INV_X1 U7697 ( .A(keyinput97), .ZN(n6736) );
  NAND4_X1 U7698 ( .A1(keyinput14), .A2(n6738), .A3(n6737), .A4(n6736), .ZN(
        n6739) );
  NOR4_X1 U7699 ( .A1(keyinput104), .A2(keyinput89), .A3(n6740), .A4(n6739), 
        .ZN(n6757) );
  INV_X1 U7700 ( .A(keyinput121), .ZN(n6741) );
  NOR4_X1 U7701 ( .A1(keyinput102), .A2(keyinput106), .A3(keyinput125), .A4(
        n6741), .ZN(n6756) );
  NAND2_X1 U7702 ( .A1(keyinput68), .A2(keyinput93), .ZN(n6742) );
  NOR3_X1 U7703 ( .A1(keyinput4), .A2(keyinput84), .A3(n6742), .ZN(n6755) );
  NAND2_X1 U7704 ( .A1(keyinput81), .A2(keyinput123), .ZN(n6743) );
  NOR3_X1 U7705 ( .A1(keyinput119), .A2(keyinput29), .A3(n6743), .ZN(n6744) );
  NAND3_X1 U7706 ( .A1(keyinput116), .A2(keyinput127), .A3(n6744), .ZN(n6753)
         );
  NAND2_X1 U7707 ( .A1(keyinput26), .A2(keyinput36), .ZN(n6745) );
  NOR3_X1 U7708 ( .A1(keyinput98), .A2(keyinput16), .A3(n6745), .ZN(n6751) );
  NAND2_X1 U7709 ( .A1(keyinput71), .A2(keyinput91), .ZN(n6746) );
  NOR3_X1 U7710 ( .A1(keyinput92), .A2(keyinput107), .A3(n6746), .ZN(n6750) );
  NOR4_X1 U7711 ( .A1(keyinput40), .A2(keyinput19), .A3(keyinput85), .A4(
        keyinput34), .ZN(n6749) );
  NAND2_X1 U7712 ( .A1(keyinput24), .A2(keyinput27), .ZN(n6747) );
  NOR3_X1 U7713 ( .A1(keyinput56), .A2(keyinput57), .A3(n6747), .ZN(n6748) );
  NAND4_X1 U7714 ( .A1(n6751), .A2(n6750), .A3(n6749), .A4(n6748), .ZN(n6752)
         );
  NOR4_X1 U7715 ( .A1(keyinput39), .A2(keyinput31), .A3(n6753), .A4(n6752), 
        .ZN(n6754) );
  NAND4_X1 U7716 ( .A1(n6757), .A2(n6756), .A3(n6755), .A4(n6754), .ZN(n6758)
         );
  NOR4_X1 U7717 ( .A1(n6761), .A2(n6760), .A3(n6759), .A4(n6758), .ZN(n6762)
         );
  AOI21_X1 U7718 ( .B1(n6763), .B2(n6762), .A(keyinput78), .ZN(n7022) );
  INV_X1 U7719 ( .A(keyinput78), .ZN(n6769) );
  XOR2_X1 U7720 ( .A(keyinput124), .B(DATAWIDTH_REG_19__SCAN_IN), .Z(n6768) );
  INV_X1 U7721 ( .A(DATAI_28_), .ZN(n6765) );
  AOI22_X1 U7722 ( .A1(n6766), .A2(keyinput86), .B1(n6765), .B2(keyinput38), 
        .ZN(n6764) );
  OAI221_X1 U7723 ( .B1(n6766), .B2(keyinput86), .C1(n6765), .C2(keyinput38), 
        .A(n6764), .ZN(n6767) );
  AOI211_X1 U7724 ( .C1(ADDRESS_REG_7__SCAN_IN), .C2(n6769), .A(n6768), .B(
        n6767), .ZN(n6793) );
  INV_X1 U7725 ( .A(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n6772) );
  INV_X1 U7726 ( .A(keyinput11), .ZN(n6771) );
  OAI22_X1 U7727 ( .A1(n6772), .A2(keyinput37), .B1(n6771), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6770) );
  AOI221_X1 U7728 ( .B1(n6772), .B2(keyinput37), .C1(DATAO_REG_3__SCAN_IN), 
        .C2(n6771), .A(n6770), .ZN(n6792) );
  INV_X1 U7729 ( .A(keyinput3), .ZN(n6774) );
  OAI22_X1 U7730 ( .A1(n6775), .A2(keyinput69), .B1(n6774), .B2(
        ADDRESS_REG_23__SCAN_IN), .ZN(n6773) );
  AOI221_X1 U7731 ( .B1(n6775), .B2(keyinput69), .C1(ADDRESS_REG_23__SCAN_IN), 
        .C2(n6774), .A(n6773), .ZN(n6791) );
  INV_X1 U7732 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6778) );
  INV_X1 U7733 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6777) );
  AOI22_X1 U7734 ( .A1(n6778), .A2(keyinput2), .B1(keyinput51), .B2(n6777), 
        .ZN(n6776) );
  OAI221_X1 U7735 ( .B1(n6778), .B2(keyinput2), .C1(n6777), .C2(keyinput51), 
        .A(n6776), .ZN(n6789) );
  INV_X1 U7736 ( .A(keyinput17), .ZN(n6780) );
  AOI22_X1 U7737 ( .A1(n6781), .A2(keyinput94), .B1(M_IO_N_REG_SCAN_IN), .B2(
        n6780), .ZN(n6779) );
  OAI221_X1 U7738 ( .B1(n6781), .B2(keyinput94), .C1(n6780), .C2(
        M_IO_N_REG_SCAN_IN), .A(n6779), .ZN(n6788) );
  AOI22_X1 U7739 ( .A1(n4381), .A2(keyinput95), .B1(keyinput30), .B2(n6783), 
        .ZN(n6782) );
  OAI221_X1 U7740 ( .B1(n4381), .B2(keyinput95), .C1(n6783), .C2(keyinput30), 
        .A(n6782), .ZN(n6787) );
  XNOR2_X1 U7741 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .B(keyinput74), .ZN(n6785)
         );
  XNOR2_X1 U7742 ( .A(keyinput22), .B(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n6784)
         );
  NAND2_X1 U7743 ( .A1(n6785), .A2(n6784), .ZN(n6786) );
  NOR4_X1 U7744 ( .A1(n6789), .A2(n6788), .A3(n6787), .A4(n6786), .ZN(n6790)
         );
  NAND4_X1 U7745 ( .A1(n6793), .A2(n6792), .A3(n6791), .A4(n6790), .ZN(n6893)
         );
  INV_X1 U7746 ( .A(keyinput112), .ZN(n6797) );
  OAI22_X1 U7747 ( .A1(keyinput8), .A2(n6798), .B1(n6797), .B2(
        BE_N_REG_3__SCAN_IN), .ZN(n6796) );
  AOI221_X1 U7748 ( .B1(n6798), .B2(keyinput8), .C1(n6797), .C2(
        BE_N_REG_3__SCAN_IN), .A(n6796), .ZN(n6807) );
  INV_X1 U7749 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n6801) );
  INV_X1 U7750 ( .A(keyinput110), .ZN(n6800) );
  OAI22_X1 U7751 ( .A1(n6801), .A2(keyinput87), .B1(n6800), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n6799) );
  AOI221_X1 U7752 ( .B1(n6801), .B2(keyinput87), .C1(UWORD_REG_14__SCAN_IN), 
        .C2(n6800), .A(n6799), .ZN(n6806) );
  INV_X1 U7753 ( .A(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n6804) );
  INV_X1 U7754 ( .A(keyinput114), .ZN(n6803) );
  OAI22_X1 U7755 ( .A1(n6804), .A2(keyinput33), .B1(n6803), .B2(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6802) );
  AOI221_X1 U7756 ( .B1(n6804), .B2(keyinput33), .C1(DATAWIDTH_REG_30__SCAN_IN), .C2(n6803), .A(n6802), .ZN(n6805) );
  NAND4_X1 U7757 ( .A1(n6808), .A2(n6807), .A3(n6806), .A4(n6805), .ZN(n6892)
         );
  OAI22_X1 U7758 ( .A1(n6811), .A2(keyinput83), .B1(n6810), .B2(keyinput1), 
        .ZN(n6809) );
  AOI221_X1 U7759 ( .B1(n6811), .B2(keyinput83), .C1(keyinput1), .C2(n6810), 
        .A(n6809), .ZN(n6823) );
  OAI22_X1 U7760 ( .A1(n6814), .A2(keyinput48), .B1(n6813), .B2(
        BYTEENABLE_REG_1__SCAN_IN), .ZN(n6812) );
  AOI221_X1 U7761 ( .B1(n6814), .B2(keyinput48), .C1(BYTEENABLE_REG_1__SCAN_IN), .C2(n6813), .A(n6812), .ZN(n6822) );
  INV_X1 U7762 ( .A(keyinput52), .ZN(n6816) );
  OAI22_X1 U7763 ( .A1(n5853), .A2(keyinput99), .B1(n6816), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n6815) );
  AOI221_X1 U7764 ( .B1(n5853), .B2(keyinput99), .C1(UWORD_REG_2__SCAN_IN), 
        .C2(n6816), .A(n6815), .ZN(n6821) );
  XNOR2_X1 U7765 ( .A(n6817), .B(ADDRESS_REG_20__SCAN_IN), .ZN(n6819) );
  XOR2_X1 U7766 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .B(keyinput5), .Z(n6818) );
  NOR2_X1 U7767 ( .A1(n6819), .A2(n6818), .ZN(n6820) );
  NAND4_X1 U7768 ( .A1(n6823), .A2(n6822), .A3(n6821), .A4(n6820), .ZN(n6891)
         );
  INV_X1 U7769 ( .A(keyinput35), .ZN(n6825) );
  AOI22_X1 U7770 ( .A1(n6826), .A2(keyinput28), .B1(LWORD_REG_7__SCAN_IN), 
        .B2(n6825), .ZN(n6824) );
  OAI221_X1 U7771 ( .B1(n6826), .B2(keyinput28), .C1(n6825), .C2(
        LWORD_REG_7__SCAN_IN), .A(n6824), .ZN(n6837) );
  AOI22_X1 U7772 ( .A1(n4925), .A2(keyinput115), .B1(n3318), .B2(keyinput67), 
        .ZN(n6827) );
  OAI221_X1 U7773 ( .B1(n4925), .B2(keyinput115), .C1(n3318), .C2(keyinput67), 
        .A(n6827), .ZN(n6836) );
  INV_X1 U7774 ( .A(keyinput43), .ZN(n6829) );
  INV_X1 U7775 ( .A(keyinput63), .ZN(n6833) );
  INV_X1 U7776 ( .A(keyinput50), .ZN(n6832) );
  AOI22_X1 U7777 ( .A1(n6833), .A2(DATAO_REG_28__SCAN_IN), .B1(
        UWORD_REG_3__SCAN_IN), .B2(n6832), .ZN(n6831) );
  OAI221_X1 U7778 ( .B1(n6833), .B2(DATAO_REG_28__SCAN_IN), .C1(n6832), .C2(
        UWORD_REG_3__SCAN_IN), .A(n6831), .ZN(n6834) );
  NOR4_X1 U7779 ( .A1(n6837), .A2(n6836), .A3(n6835), .A4(n6834), .ZN(n6889)
         );
  INV_X1 U7780 ( .A(keyinput90), .ZN(n6840) );
  INV_X1 U7781 ( .A(keyinput64), .ZN(n6839) );
  AOI22_X1 U7782 ( .A1(n6840), .A2(BE_N_REG_1__SCAN_IN), .B1(
        DATAWIDTH_REG_9__SCAN_IN), .B2(n6839), .ZN(n6838) );
  OAI221_X1 U7783 ( .B1(n6840), .B2(BE_N_REG_1__SCAN_IN), .C1(n6839), .C2(
        DATAWIDTH_REG_9__SCAN_IN), .A(n6838), .ZN(n6853) );
  INV_X1 U7784 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n6843) );
  AOI22_X1 U7785 ( .A1(n6843), .A2(keyinput79), .B1(keyinput10), .B2(n6842), 
        .ZN(n6841) );
  OAI221_X1 U7786 ( .B1(n6843), .B2(keyinput79), .C1(n6842), .C2(keyinput10), 
        .A(n6841), .ZN(n6852) );
  INV_X1 U7787 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n6846) );
  AOI22_X1 U7788 ( .A1(n6846), .A2(keyinput13), .B1(keyinput32), .B2(n6845), 
        .ZN(n6844) );
  OAI221_X1 U7789 ( .B1(n6846), .B2(keyinput13), .C1(n6845), .C2(keyinput32), 
        .A(n6844), .ZN(n6851) );
  INV_X1 U7790 ( .A(keyinput60), .ZN(n6849) );
  INV_X1 U7791 ( .A(keyinput96), .ZN(n6848) );
  AOI22_X1 U7792 ( .A1(n6849), .A2(DATAO_REG_11__SCAN_IN), .B1(
        DATAO_REG_8__SCAN_IN), .B2(n6848), .ZN(n6847) );
  OAI221_X1 U7793 ( .B1(n6849), .B2(DATAO_REG_11__SCAN_IN), .C1(n6848), .C2(
        DATAO_REG_8__SCAN_IN), .A(n6847), .ZN(n6850) );
  NOR4_X1 U7794 ( .A1(n6853), .A2(n6852), .A3(n6851), .A4(n6850), .ZN(n6888)
         );
  INV_X1 U7795 ( .A(keyinput122), .ZN(n6855) );
  AOI22_X1 U7796 ( .A1(n6856), .A2(keyinput73), .B1(ADDRESS_REG_8__SCAN_IN), 
        .B2(n6855), .ZN(n6854) );
  OAI221_X1 U7797 ( .B1(n6856), .B2(keyinput73), .C1(n6855), .C2(
        ADDRESS_REG_8__SCAN_IN), .A(n6854), .ZN(n6869) );
  INV_X1 U7798 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n6862) );
  AOI22_X1 U7799 ( .A1(n6862), .A2(keyinput23), .B1(keyinput97), .B2(n6861), 
        .ZN(n6860) );
  OAI221_X1 U7800 ( .B1(n6862), .B2(keyinput23), .C1(n6861), .C2(keyinput97), 
        .A(n6860), .ZN(n6867) );
  INV_X1 U7801 ( .A(DATAI_8_), .ZN(n6864) );
  AOI22_X1 U7802 ( .A1(n6865), .A2(keyinput111), .B1(keyinput49), .B2(n6864), 
        .ZN(n6863) );
  OAI221_X1 U7803 ( .B1(n6865), .B2(keyinput111), .C1(n6864), .C2(keyinput49), 
        .A(n6863), .ZN(n6866) );
  NOR4_X1 U7804 ( .A1(n6869), .A2(n6868), .A3(n6867), .A4(n6866), .ZN(n6887)
         );
  INV_X1 U7805 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6871) );
  AOI22_X1 U7806 ( .A1(n6872), .A2(keyinput46), .B1(keyinput66), .B2(n6871), 
        .ZN(n6870) );
  OAI221_X1 U7807 ( .B1(n6872), .B2(keyinput46), .C1(n6871), .C2(keyinput66), 
        .A(n6870), .ZN(n6885) );
  INV_X1 U7808 ( .A(keyinput25), .ZN(n6874) );
  AOI22_X1 U7809 ( .A1(n6875), .A2(keyinput15), .B1(DATAO_REG_26__SCAN_IN), 
        .B2(n6874), .ZN(n6873) );
  OAI221_X1 U7810 ( .B1(n6875), .B2(keyinput15), .C1(n6874), .C2(
        DATAO_REG_26__SCAN_IN), .A(n6873), .ZN(n6884) );
  INV_X1 U7811 ( .A(keyinput77), .ZN(n6877) );
  AOI22_X1 U7812 ( .A1(n6878), .A2(keyinput0), .B1(CODEFETCH_REG_SCAN_IN), 
        .B2(n6877), .ZN(n6876) );
  OAI221_X1 U7813 ( .B1(n6878), .B2(keyinput0), .C1(n6877), .C2(
        CODEFETCH_REG_SCAN_IN), .A(n6876), .ZN(n6883) );
  INV_X1 U7814 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n6881) );
  AOI22_X1 U7815 ( .A1(n6881), .A2(keyinput72), .B1(keyinput76), .B2(n6880), 
        .ZN(n6879) );
  OAI221_X1 U7816 ( .B1(n6881), .B2(keyinput72), .C1(n6880), .C2(keyinput76), 
        .A(n6879), .ZN(n6882) );
  NOR4_X1 U7817 ( .A1(n6885), .A2(n6884), .A3(n6883), .A4(n6882), .ZN(n6886)
         );
  NAND4_X1 U7818 ( .A1(n6889), .A2(n6888), .A3(n6887), .A4(n6886), .ZN(n6890)
         );
  NOR4_X1 U7819 ( .A1(n6893), .A2(n6892), .A3(n6891), .A4(n6890), .ZN(n7021)
         );
  INV_X1 U7820 ( .A(keyinput14), .ZN(n6895) );
  OAI22_X1 U7821 ( .A1(n6896), .A2(keyinput126), .B1(n6895), .B2(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n6894) );
  AOI221_X1 U7822 ( .B1(n6896), .B2(keyinput126), .C1(
        DATAWIDTH_REG_17__SCAN_IN), .C2(n6895), .A(n6894), .ZN(n6907) );
  INV_X1 U7823 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n6899) );
  INV_X1 U7824 ( .A(keyinput62), .ZN(n6898) );
  OAI22_X1 U7825 ( .A1(n6899), .A2(keyinput61), .B1(n6898), .B2(
        LWORD_REG_6__SCAN_IN), .ZN(n6897) );
  AOI221_X1 U7826 ( .B1(n6899), .B2(keyinput61), .C1(LWORD_REG_6__SCAN_IN), 
        .C2(n6898), .A(n6897), .ZN(n6906) );
  INV_X1 U7827 ( .A(keyinput45), .ZN(n6901) );
  OAI22_X1 U7828 ( .A1(n4322), .A2(keyinput41), .B1(n6901), .B2(
        ADDRESS_REG_29__SCAN_IN), .ZN(n6900) );
  AOI221_X1 U7829 ( .B1(n4322), .B2(keyinput41), .C1(ADDRESS_REG_29__SCAN_IN), 
        .C2(n6901), .A(n6900), .ZN(n6905) );
  INV_X1 U7830 ( .A(keyinput103), .ZN(n6903) );
  OAI22_X1 U7831 ( .A1(n5110), .A2(keyinput6), .B1(n6903), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6902) );
  AOI221_X1 U7832 ( .B1(n5110), .B2(keyinput6), .C1(DATAO_REG_7__SCAN_IN), 
        .C2(n6903), .A(n6902), .ZN(n6904) );
  NAND4_X1 U7833 ( .A1(n6907), .A2(n6906), .A3(n6905), .A4(n6904), .ZN(n7019)
         );
  AOI22_X1 U7834 ( .A1(n6910), .A2(keyinput80), .B1(n6909), .B2(keyinput55), 
        .ZN(n6908) );
  OAI221_X1 U7835 ( .B1(n6910), .B2(keyinput80), .C1(n6909), .C2(keyinput55), 
        .A(n6908), .ZN(n6921) );
  INV_X1 U7836 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n6914) );
  AOI22_X1 U7837 ( .A1(n6914), .A2(keyinput54), .B1(keyinput101), .B2(n4473), 
        .ZN(n6913) );
  OAI221_X1 U7838 ( .B1(n6914), .B2(keyinput54), .C1(n4473), .C2(keyinput101), 
        .A(n6913), .ZN(n6919) );
  AOI22_X1 U7839 ( .A1(n6917), .A2(keyinput42), .B1(DATAO_REG_20__SCAN_IN), 
        .B2(n6916), .ZN(n6915) );
  OAI221_X1 U7840 ( .B1(n6917), .B2(keyinput42), .C1(n6916), .C2(
        DATAO_REG_20__SCAN_IN), .A(n6915), .ZN(n6918) );
  NOR4_X1 U7841 ( .A1(n6921), .A2(n6920), .A3(n6919), .A4(n6918), .ZN(n6954)
         );
  OAI22_X1 U7842 ( .A1(keyinput117), .A2(n6924), .B1(n6923), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n6922) );
  AOI221_X1 U7843 ( .B1(n6924), .B2(keyinput117), .C1(n6923), .C2(
        UWORD_REG_11__SCAN_IN), .A(n6922), .ZN(n6953) );
  AOI22_X1 U7844 ( .A1(n6927), .A2(keyinput9), .B1(keyinput21), .B2(n6926), 
        .ZN(n6925) );
  OAI221_X1 U7845 ( .B1(n6927), .B2(keyinput9), .C1(n6926), .C2(keyinput21), 
        .A(n6925), .ZN(n6935) );
  INV_X1 U7846 ( .A(keyinput53), .ZN(n6929) );
  AOI22_X1 U7847 ( .A1(n6930), .A2(keyinput113), .B1(ADDRESS_REG_0__SCAN_IN), 
        .B2(n6929), .ZN(n6928) );
  OAI221_X1 U7848 ( .B1(n6930), .B2(keyinput113), .C1(n6929), .C2(
        ADDRESS_REG_0__SCAN_IN), .A(n6928), .ZN(n6934) );
  AOI22_X1 U7849 ( .A1(n4132), .A2(keyinput47), .B1(keyinput109), .B2(n6932), 
        .ZN(n6931) );
  OAI221_X1 U7850 ( .B1(n4132), .B2(keyinput47), .C1(n6932), .C2(keyinput109), 
        .A(n6931), .ZN(n6933) );
  NOR3_X1 U7851 ( .A1(n6935), .A2(n6934), .A3(n6933), .ZN(n6952) );
  AOI22_X1 U7852 ( .A1(n6938), .A2(keyinput75), .B1(n6937), .B2(keyinput104), 
        .ZN(n6936) );
  OAI221_X1 U7853 ( .B1(n6938), .B2(keyinput75), .C1(n6937), .C2(keyinput104), 
        .A(n6936), .ZN(n6950) );
  INV_X1 U7854 ( .A(keyinput89), .ZN(n6940) );
  AOI22_X1 U7855 ( .A1(n3544), .A2(keyinput59), .B1(LWORD_REG_14__SCAN_IN), 
        .B2(n6940), .ZN(n6939) );
  OAI221_X1 U7856 ( .B1(n3544), .B2(keyinput59), .C1(n6940), .C2(
        LWORD_REG_14__SCAN_IN), .A(n6939), .ZN(n6949) );
  INV_X1 U7857 ( .A(keyinput100), .ZN(n6942) );
  AOI22_X1 U7858 ( .A1(n6943), .A2(keyinput120), .B1(UWORD_REG_7__SCAN_IN), 
        .B2(n6942), .ZN(n6941) );
  OAI221_X1 U7859 ( .B1(n6943), .B2(keyinput120), .C1(n6942), .C2(
        UWORD_REG_7__SCAN_IN), .A(n6941), .ZN(n6948) );
  INV_X1 U7860 ( .A(keyinput93), .ZN(n6945) );
  AOI22_X1 U7861 ( .A1(n6946), .A2(keyinput20), .B1(ADDRESS_REG_24__SCAN_IN), 
        .B2(n6945), .ZN(n6944) );
  OAI221_X1 U7862 ( .B1(n6946), .B2(keyinput20), .C1(n6945), .C2(
        ADDRESS_REG_24__SCAN_IN), .A(n6944), .ZN(n6947) );
  NOR4_X1 U7863 ( .A1(n6950), .A2(n6949), .A3(n6948), .A4(n6947), .ZN(n6951)
         );
  NAND4_X1 U7864 ( .A1(n6954), .A2(n6953), .A3(n6952), .A4(n6951), .ZN(n7018)
         );
  INV_X1 U7865 ( .A(keyinput92), .ZN(n6956) );
  OAI22_X1 U7866 ( .A1(n4926), .A2(keyinput71), .B1(n6956), .B2(
        ADDRESS_REG_26__SCAN_IN), .ZN(n6955) );
  AOI221_X1 U7867 ( .B1(n4926), .B2(keyinput71), .C1(ADDRESS_REG_26__SCAN_IN), 
        .C2(n6956), .A(n6955), .ZN(n6968) );
  INV_X1 U7868 ( .A(keyinput98), .ZN(n6958) );
  OAI22_X1 U7869 ( .A1(n3918), .A2(keyinput107), .B1(n6958), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n6957) );
  AOI221_X1 U7870 ( .B1(n3918), .B2(keyinput107), .C1(UWORD_REG_9__SCAN_IN), 
        .C2(n6958), .A(n6957), .ZN(n6967) );
  INV_X1 U7871 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n6961) );
  INV_X1 U7872 ( .A(keyinput36), .ZN(n6960) );
  OAI22_X1 U7873 ( .A1(n6961), .A2(keyinput26), .B1(n6960), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6959) );
  AOI221_X1 U7874 ( .B1(n6961), .B2(keyinput26), .C1(DATAO_REG_15__SCAN_IN), 
        .C2(n6960), .A(n6959), .ZN(n6966) );
  INV_X1 U7875 ( .A(DATAI_26_), .ZN(n6964) );
  INV_X1 U7876 ( .A(DATAI_21_), .ZN(n6963) );
  OAI22_X1 U7877 ( .A1(n6964), .A2(keyinput16), .B1(n6963), .B2(keyinput119), 
        .ZN(n6962) );
  AOI221_X1 U7878 ( .B1(n6964), .B2(keyinput16), .C1(keyinput119), .C2(n6963), 
        .A(n6962), .ZN(n6965) );
  NAND4_X1 U7879 ( .A1(n6968), .A2(n6967), .A3(n6966), .A4(n6965), .ZN(n7017)
         );
  INV_X1 U7880 ( .A(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n6971) );
  AOI22_X1 U7881 ( .A1(n6971), .A2(keyinput125), .B1(keyinput91), .B2(n6970), 
        .ZN(n6969) );
  OAI221_X1 U7882 ( .B1(n6971), .B2(keyinput125), .C1(n6970), .C2(keyinput91), 
        .A(n6969), .ZN(n6983) );
  INV_X1 U7883 ( .A(keyinput84), .ZN(n6973) );
  AOI22_X1 U7884 ( .A1(n6974), .A2(keyinput4), .B1(DATAO_REG_5__SCAN_IN), .B2(
        n6973), .ZN(n6972) );
  OAI221_X1 U7885 ( .B1(n6974), .B2(keyinput4), .C1(n6973), .C2(
        DATAO_REG_5__SCAN_IN), .A(n6972), .ZN(n6982) );
  INV_X1 U7886 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n6976) );
  AOI22_X1 U7887 ( .A1(n3898), .A2(keyinput68), .B1(n6976), .B2(keyinput121), 
        .ZN(n6975) );
  OAI221_X1 U7888 ( .B1(n3898), .B2(keyinput68), .C1(n6976), .C2(keyinput121), 
        .A(n6975), .ZN(n6981) );
  INV_X1 U7889 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6977) );
  XOR2_X1 U7890 ( .A(n6977), .B(keyinput102), .Z(n6979) );
  XNOR2_X1 U7891 ( .A(INSTQUEUE_REG_9__6__SCAN_IN), .B(keyinput106), .ZN(n6978) );
  NAND2_X1 U7892 ( .A1(n6979), .A2(n6978), .ZN(n6980) );
  NOR4_X1 U7893 ( .A1(n6983), .A2(n6982), .A3(n6981), .A4(n6980), .ZN(n7015)
         );
  INV_X1 U7894 ( .A(keyinput39), .ZN(n6985) );
  OAI22_X1 U7895 ( .A1(keyinput123), .A2(n6986), .B1(n6985), .B2(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n6984) );
  AOI221_X1 U7896 ( .B1(n6986), .B2(keyinput123), .C1(n6985), .C2(
        DATAWIDTH_REG_21__SCAN_IN), .A(n6984), .ZN(n7014) );
  INV_X1 U7897 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n6988) );
  AOI22_X1 U7898 ( .A1(n5668), .A2(keyinput31), .B1(n6988), .B2(keyinput29), 
        .ZN(n6987) );
  OAI221_X1 U7899 ( .B1(n5668), .B2(keyinput31), .C1(n6988), .C2(keyinput29), 
        .A(n6987), .ZN(n6996) );
  INV_X1 U7900 ( .A(DATAI_24_), .ZN(n6990) );
  AOI22_X1 U7901 ( .A1(n4108), .A2(keyinput81), .B1(keyinput116), .B2(n6990), 
        .ZN(n6989) );
  OAI221_X1 U7902 ( .B1(n4108), .B2(keyinput81), .C1(n6990), .C2(keyinput116), 
        .A(n6989), .ZN(n6995) );
  INV_X1 U7903 ( .A(keyinput127), .ZN(n6992) );
  AOI22_X1 U7904 ( .A1(n6993), .A2(keyinput56), .B1(DATAO_REG_31__SCAN_IN), 
        .B2(n6992), .ZN(n6991) );
  OAI221_X1 U7905 ( .B1(n6993), .B2(keyinput56), .C1(n6992), .C2(
        DATAO_REG_31__SCAN_IN), .A(n6991), .ZN(n6994) );
  NOR3_X1 U7906 ( .A1(n6996), .A2(n6995), .A3(n6994), .ZN(n7013) );
  AOI22_X1 U7907 ( .A1(n4081), .A2(keyinput27), .B1(keyinput40), .B2(n6998), 
        .ZN(n6997) );
  OAI221_X1 U7908 ( .B1(n4081), .B2(keyinput27), .C1(n6998), .C2(keyinput40), 
        .A(n6997), .ZN(n7011) );
  INV_X1 U7909 ( .A(keyinput19), .ZN(n7000) );
  AOI22_X1 U7910 ( .A1(n7001), .A2(keyinput85), .B1(DATAO_REG_23__SCAN_IN), 
        .B2(n7000), .ZN(n6999) );
  OAI221_X1 U7911 ( .B1(n7001), .B2(keyinput85), .C1(n7000), .C2(
        DATAO_REG_23__SCAN_IN), .A(n6999), .ZN(n7010) );
  INV_X1 U7912 ( .A(keyinput24), .ZN(n7003) );
  AOI22_X1 U7913 ( .A1(n7004), .A2(keyinput34), .B1(DATAO_REG_2__SCAN_IN), 
        .B2(n7003), .ZN(n7002) );
  OAI221_X1 U7914 ( .B1(n7004), .B2(keyinput34), .C1(n7003), .C2(
        DATAO_REG_2__SCAN_IN), .A(n7002), .ZN(n7009) );
  INV_X1 U7915 ( .A(keyinput105), .ZN(n7006) );
  AOI22_X1 U7916 ( .A1(n7007), .A2(keyinput57), .B1(ADDRESS_REG_17__SCAN_IN), 
        .B2(n7006), .ZN(n7005) );
  OAI221_X1 U7917 ( .B1(n7007), .B2(keyinput57), .C1(n7006), .C2(
        ADDRESS_REG_17__SCAN_IN), .A(n7005), .ZN(n7008) );
  NOR4_X1 U7918 ( .A1(n7011), .A2(n7010), .A3(n7009), .A4(n7008), .ZN(n7012)
         );
  NAND4_X1 U7919 ( .A1(n7015), .A2(n7014), .A3(n7013), .A4(n7012), .ZN(n7016)
         );
  NOR4_X1 U7920 ( .A1(n7019), .A2(n7018), .A3(n7017), .A4(n7016), .ZN(n7020)
         );
  OAI211_X1 U7921 ( .C1(ADDRESS_REG_7__SCAN_IN), .C2(n7022), .A(n7021), .B(
        n7020), .ZN(n7023) );
  XNOR2_X1 U7922 ( .A(n7024), .B(n7023), .ZN(U2935) );
  AND4_X1 U3887 ( .A1(n3123), .A2(n3122), .A3(n3121), .A4(n3120), .ZN(n3142)
         );
  CLKBUF_X1 U3588 ( .A(n3496), .Z(n5690) );
  CLKBUF_X2 U3603 ( .A(n3267), .Z(n5681) );
  CLKBUF_X1 U4028 ( .A(n3494), .Z(n3110) );
  CLKBUF_X1 U4343 ( .A(n6280), .Z(n6283) );
endmodule

